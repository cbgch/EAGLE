//Key = 1100111101011100110111001111000011111011001011010001010001110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389;

XNOR2_X1 U766 ( .A(G107), .B(n1056), .ZN(G9) );
NAND3_X1 U767 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
XNOR2_X1 U768 ( .A(n1060), .B(KEYINPUT34), .ZN(n1059) );
NOR2_X1 U769 ( .A1(n1061), .A2(n1062), .ZN(G75) );
NOR4_X1 U770 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
XOR2_X1 U771 ( .A(n1067), .B(KEYINPUT4), .Z(n1066) );
NAND3_X1 U772 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
OR4_X1 U773 ( .A1(n1071), .A2(n1072), .A3(KEYINPUT40), .A4(n1073), .ZN(n1063) );
NOR2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
INV_X1 U775 ( .A(n1070), .ZN(n1075) );
NOR3_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1070) );
NOR2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR3_X1 U781 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1079) );
NOR2_X1 U782 ( .A1(n1090), .A2(n1089), .ZN(n1071) );
NOR2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U784 ( .A1(KEYINPUT32), .A2(n1093), .ZN(n1092) );
NOR4_X1 U785 ( .A1(n1077), .A2(n1094), .A3(n1082), .A4(n1078), .ZN(n1093) );
NOR3_X1 U786 ( .A1(n1078), .A2(n1095), .A3(n1082), .ZN(n1091) );
INV_X1 U787 ( .A(n1096), .ZN(n1082) );
NOR2_X1 U788 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NOR2_X1 U789 ( .A1(n1099), .A2(n1076), .ZN(n1098) );
INV_X1 U790 ( .A(n1100), .ZN(n1076) );
NOR2_X1 U791 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
INV_X1 U793 ( .A(n1105), .ZN(n1103) );
NOR2_X1 U794 ( .A1(n1106), .A2(n1077), .ZN(n1097) );
NOR2_X1 U795 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
AND2_X1 U796 ( .A1(n1058), .A2(KEYINPUT32), .ZN(n1107) );
NOR3_X1 U797 ( .A1(n1065), .A2(G952), .A3(n1073), .ZN(n1061) );
AND4_X1 U798 ( .A1(n1109), .A2(n1110), .A3(n1068), .A4(n1087), .ZN(n1073) );
XOR2_X1 U799 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U800 ( .A(KEYINPUT36), .B(KEYINPUT35), .Z(n1112) );
XOR2_X1 U801 ( .A(n1113), .B(G469), .Z(n1111) );
XOR2_X1 U802 ( .A(n1114), .B(KEYINPUT53), .Z(n1109) );
NAND4_X1 U803 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1114) );
NOR2_X1 U804 ( .A1(n1119), .A2(n1105), .ZN(n1118) );
XNOR2_X1 U805 ( .A(n1120), .B(KEYINPUT44), .ZN(n1119) );
NAND2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1116) );
XNOR2_X1 U807 ( .A(KEYINPUT3), .B(n1123), .ZN(n1121) );
NAND2_X1 U808 ( .A1(n1124), .A2(G475), .ZN(n1115) );
XNOR2_X1 U809 ( .A(KEYINPUT59), .B(n1123), .ZN(n1124) );
INV_X1 U810 ( .A(n1125), .ZN(n1065) );
XOR2_X1 U811 ( .A(n1126), .B(n1127), .Z(G72) );
XOR2_X1 U812 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR3_X1 U813 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
AND2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR2_X1 U817 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
INV_X1 U818 ( .A(KEYINPUT29), .ZN(n1139) );
NOR2_X1 U819 ( .A1(KEYINPUT29), .A2(n1133), .ZN(n1136) );
NOR2_X1 U820 ( .A1(n1140), .A2(n1138), .ZN(n1133) );
XNOR2_X1 U821 ( .A(n1141), .B(n1142), .ZN(n1138) );
XNOR2_X1 U822 ( .A(n1143), .B(n1144), .ZN(n1142) );
XNOR2_X1 U823 ( .A(G134), .B(G137), .ZN(n1141) );
INV_X1 U824 ( .A(KEYINPUT20), .ZN(n1140) );
NOR2_X1 U825 ( .A1(G900), .A2(n1145), .ZN(n1130) );
NAND3_X1 U826 ( .A1(G953), .A2(n1146), .A3(KEYINPUT1), .ZN(n1128) );
XOR2_X1 U827 ( .A(KEYINPUT62), .B(n1147), .Z(n1146) );
NOR2_X1 U828 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U829 ( .A1(n1145), .A2(n1150), .ZN(n1126) );
NAND2_X1 U830 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND2_X1 U831 ( .A1(n1153), .A2(n1154), .ZN(G69) );
NAND2_X1 U832 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
OR2_X1 U833 ( .A1(n1145), .A2(G224), .ZN(n1156) );
NAND3_X1 U834 ( .A1(G953), .A2(n1157), .A3(n1158), .ZN(n1153) );
INV_X1 U835 ( .A(n1155), .ZN(n1158) );
XNOR2_X1 U836 ( .A(n1159), .B(n1160), .ZN(n1155) );
NOR2_X1 U837 ( .A1(n1161), .A2(G953), .ZN(n1160) );
NOR2_X1 U838 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND3_X1 U839 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1159) );
INV_X1 U840 ( .A(n1167), .ZN(n1166) );
NAND2_X1 U841 ( .A1(G953), .A2(n1168), .ZN(n1164) );
NAND2_X1 U842 ( .A1(G898), .A2(G224), .ZN(n1157) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1170), .ZN(G66) );
XNOR2_X1 U844 ( .A(n1171), .B(n1172), .ZN(n1170) );
NOR2_X1 U845 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U846 ( .A1(n1169), .A2(n1175), .ZN(G63) );
XNOR2_X1 U847 ( .A(n1176), .B(n1177), .ZN(n1175) );
NOR2_X1 U848 ( .A1(n1178), .A2(n1174), .ZN(n1177) );
NOR2_X1 U849 ( .A1(n1169), .A2(n1179), .ZN(G60) );
XOR2_X1 U850 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U851 ( .A1(n1122), .A2(n1174), .ZN(n1181) );
NOR2_X1 U852 ( .A1(KEYINPUT41), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U853 ( .A(G104), .B(n1183), .ZN(G6) );
NOR2_X1 U854 ( .A1(n1169), .A2(n1184), .ZN(G57) );
XOR2_X1 U855 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U856 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NOR2_X1 U857 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
INV_X1 U858 ( .A(KEYINPUT25), .ZN(n1190) );
NOR2_X1 U859 ( .A1(KEYINPUT25), .A2(n1191), .ZN(n1187) );
NOR2_X1 U860 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U861 ( .A(n1194), .B(n1195), .Z(n1185) );
NOR2_X1 U862 ( .A1(n1196), .A2(n1174), .ZN(n1195) );
NAND2_X1 U863 ( .A1(n1197), .A2(n1198), .ZN(n1194) );
NOR2_X1 U864 ( .A1(n1169), .A2(n1199), .ZN(G54) );
XOR2_X1 U865 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U866 ( .A(KEYINPUT2), .B(n1202), .Z(n1201) );
NOR2_X1 U867 ( .A1(n1174), .A2(n1203), .ZN(n1202) );
XOR2_X1 U868 ( .A(KEYINPUT63), .B(G469), .Z(n1203) );
XOR2_X1 U869 ( .A(n1204), .B(n1205), .Z(n1200) );
NAND2_X1 U870 ( .A1(n1206), .A2(n1207), .ZN(n1204) );
NAND2_X1 U871 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U872 ( .A(KEYINPUT16), .B(n1210), .Z(n1206) );
NOR2_X1 U873 ( .A1(n1208), .A2(n1209), .ZN(n1210) );
NOR2_X1 U874 ( .A1(n1169), .A2(n1211), .ZN(G51) );
XOR2_X1 U875 ( .A(n1212), .B(n1213), .Z(n1211) );
NOR2_X1 U876 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U877 ( .A(KEYINPUT14), .B(n1216), .Z(n1215) );
NOR2_X1 U878 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U879 ( .A(n1219), .B(n1220), .Z(n1217) );
XOR2_X1 U880 ( .A(KEYINPUT45), .B(KEYINPUT18), .Z(n1220) );
NOR2_X1 U881 ( .A1(n1221), .A2(n1219), .ZN(n1214) );
XOR2_X1 U882 ( .A(n1222), .B(n1223), .Z(n1212) );
NOR3_X1 U883 ( .A1(n1174), .A2(n1224), .A3(n1225), .ZN(n1223) );
NAND2_X1 U884 ( .A1(G902), .A2(n1064), .ZN(n1174) );
NAND4_X1 U885 ( .A1(n1226), .A2(n1151), .A3(n1227), .A4(n1228), .ZN(n1064) );
XNOR2_X1 U886 ( .A(KEYINPUT11), .B(n1152), .ZN(n1228) );
INV_X1 U887 ( .A(n1163), .ZN(n1227) );
NAND4_X1 U888 ( .A1(n1229), .A2(n1183), .A3(n1230), .A4(n1231), .ZN(n1163) );
NAND3_X1 U889 ( .A1(n1057), .A2(n1060), .A3(n1108), .ZN(n1183) );
NAND3_X1 U890 ( .A1(n1058), .A2(n1060), .A3(n1057), .ZN(n1229) );
AND4_X1 U891 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1151) );
AND4_X1 U892 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
XOR2_X1 U893 ( .A(n1162), .B(KEYINPUT27), .Z(n1226) );
NAND4_X1 U894 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1162) );
NAND3_X1 U895 ( .A1(n1244), .A2(n1096), .A3(n1245), .ZN(n1241) );
NOR3_X1 U896 ( .A1(n1246), .A2(n1247), .A3(n1094), .ZN(n1245) );
INV_X1 U897 ( .A(n1058), .ZN(n1094) );
XOR2_X1 U898 ( .A(n1248), .B(KEYINPUT47), .Z(n1247) );
XNOR2_X1 U899 ( .A(n1084), .B(KEYINPUT7), .ZN(n1244) );
NAND2_X1 U900 ( .A1(n1084), .A2(n1249), .ZN(n1240) );
XNOR2_X1 U901 ( .A(KEYINPUT30), .B(n1250), .ZN(n1249) );
NOR2_X1 U902 ( .A1(n1145), .A2(G952), .ZN(n1169) );
XNOR2_X1 U903 ( .A(G146), .B(n1234), .ZN(G48) );
NAND2_X1 U904 ( .A1(n1251), .A2(n1108), .ZN(n1234) );
XNOR2_X1 U905 ( .A(n1252), .B(n1232), .ZN(G45) );
NAND4_X1 U906 ( .A1(n1253), .A2(n1084), .A3(n1120), .A4(n1254), .ZN(n1232) );
NAND2_X1 U907 ( .A1(KEYINPUT33), .A2(n1255), .ZN(n1252) );
XNOR2_X1 U908 ( .A(G140), .B(n1233), .ZN(G42) );
NAND4_X1 U909 ( .A1(n1256), .A2(n1108), .A3(n1117), .A4(n1068), .ZN(n1233) );
XOR2_X1 U910 ( .A(n1238), .B(n1257), .Z(G39) );
XNOR2_X1 U911 ( .A(G137), .B(KEYINPUT22), .ZN(n1257) );
NAND4_X1 U912 ( .A1(n1100), .A2(n1256), .A3(n1068), .A4(n1104), .ZN(n1238) );
XNOR2_X1 U913 ( .A(G134), .B(n1258), .ZN(G36) );
NAND2_X1 U914 ( .A1(KEYINPUT13), .A2(n1259), .ZN(n1258) );
INV_X1 U915 ( .A(n1237), .ZN(n1259) );
NAND3_X1 U916 ( .A1(n1068), .A2(n1058), .A3(n1253), .ZN(n1237) );
XNOR2_X1 U917 ( .A(G131), .B(n1236), .ZN(G33) );
NAND3_X1 U918 ( .A1(n1108), .A2(n1068), .A3(n1253), .ZN(n1236) );
AND3_X1 U919 ( .A1(n1069), .A2(n1260), .A3(n1102), .ZN(n1253) );
INV_X1 U920 ( .A(n1089), .ZN(n1068) );
NAND2_X1 U921 ( .A1(n1261), .A2(n1086), .ZN(n1089) );
INV_X1 U922 ( .A(n1085), .ZN(n1261) );
XNOR2_X1 U923 ( .A(G128), .B(n1152), .ZN(G30) );
NAND2_X1 U924 ( .A1(n1251), .A2(n1058), .ZN(n1152) );
AND3_X1 U925 ( .A1(n1084), .A2(n1104), .A3(n1256), .ZN(n1251) );
AND3_X1 U926 ( .A1(n1105), .A2(n1260), .A3(n1069), .ZN(n1256) );
XNOR2_X1 U927 ( .A(G101), .B(n1230), .ZN(G3) );
NAND3_X1 U928 ( .A1(n1102), .A2(n1057), .A3(n1100), .ZN(n1230) );
XNOR2_X1 U929 ( .A(G125), .B(n1239), .ZN(G27) );
NAND4_X1 U930 ( .A1(n1117), .A2(n1108), .A3(n1096), .A4(n1262), .ZN(n1239) );
AND3_X1 U931 ( .A1(n1084), .A2(n1260), .A3(n1105), .ZN(n1262) );
NAND2_X1 U932 ( .A1(n1263), .A2(n1078), .ZN(n1260) );
NAND4_X1 U933 ( .A1(G953), .A2(G902), .A3(n1264), .A4(n1149), .ZN(n1263) );
INV_X1 U934 ( .A(G900), .ZN(n1149) );
XOR2_X1 U935 ( .A(G122), .B(n1265), .Z(G24) );
NOR2_X1 U936 ( .A1(n1266), .A2(n1250), .ZN(n1265) );
NAND3_X1 U937 ( .A1(n1096), .A2(n1060), .A3(n1267), .ZN(n1250) );
AND3_X1 U938 ( .A1(n1120), .A2(n1248), .A3(n1254), .ZN(n1267) );
INV_X1 U939 ( .A(n1077), .ZN(n1060) );
NAND2_X1 U940 ( .A1(n1268), .A2(n1117), .ZN(n1077) );
XNOR2_X1 U941 ( .A(G119), .B(n1242), .ZN(G21) );
NAND4_X1 U942 ( .A1(n1269), .A2(n1100), .A3(n1105), .A4(n1104), .ZN(n1242) );
XNOR2_X1 U943 ( .A(G116), .B(n1270), .ZN(G18) );
NAND4_X1 U944 ( .A1(KEYINPUT19), .A2(n1269), .A3(n1102), .A4(n1058), .ZN(n1270) );
NOR2_X1 U945 ( .A1(n1254), .A2(n1271), .ZN(n1058) );
INV_X1 U946 ( .A(n1120), .ZN(n1271) );
XNOR2_X1 U947 ( .A(G113), .B(n1243), .ZN(G15) );
NAND3_X1 U948 ( .A1(n1108), .A2(n1102), .A3(n1269), .ZN(n1243) );
AND3_X1 U949 ( .A1(n1084), .A2(n1248), .A3(n1096), .ZN(n1269) );
NOR2_X1 U950 ( .A1(n1088), .A2(n1272), .ZN(n1096) );
INV_X1 U951 ( .A(n1087), .ZN(n1272) );
INV_X1 U952 ( .A(n1246), .ZN(n1102) );
NAND2_X1 U953 ( .A1(n1268), .A2(n1104), .ZN(n1246) );
XNOR2_X1 U954 ( .A(n1105), .B(KEYINPUT23), .ZN(n1268) );
NOR2_X1 U955 ( .A1(n1120), .A2(n1273), .ZN(n1108) );
INV_X1 U956 ( .A(n1254), .ZN(n1273) );
XNOR2_X1 U957 ( .A(G110), .B(n1231), .ZN(G12) );
NAND4_X1 U958 ( .A1(n1100), .A2(n1057), .A3(n1117), .A4(n1105), .ZN(n1231) );
XOR2_X1 U959 ( .A(n1274), .B(n1173), .Z(n1105) );
NAND2_X1 U960 ( .A1(G217), .A2(n1275), .ZN(n1173) );
NAND2_X1 U961 ( .A1(n1171), .A2(n1276), .ZN(n1274) );
XNOR2_X1 U962 ( .A(n1277), .B(n1278), .ZN(n1171) );
XOR2_X1 U963 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U964 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U965 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U966 ( .A(n1285), .B(KEYINPUT39), .Z(n1284) );
NAND2_X1 U967 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U968 ( .A(KEYINPUT58), .B(n1208), .ZN(n1286) );
NOR2_X1 U969 ( .A1(n1208), .A2(n1287), .ZN(n1283) );
NOR2_X1 U970 ( .A1(KEYINPUT56), .A2(n1288), .ZN(n1281) );
XNOR2_X1 U971 ( .A(G119), .B(G128), .ZN(n1288) );
XOR2_X1 U972 ( .A(n1289), .B(n1290), .Z(n1277) );
NOR2_X1 U973 ( .A1(KEYINPUT31), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U974 ( .A(n1292), .B(n1293), .ZN(n1291) );
INV_X1 U975 ( .A(G137), .ZN(n1293) );
NAND2_X1 U976 ( .A1(n1294), .A2(G221), .ZN(n1292) );
XNOR2_X1 U977 ( .A(G110), .B(KEYINPUT10), .ZN(n1289) );
INV_X1 U978 ( .A(n1104), .ZN(n1117) );
XOR2_X1 U979 ( .A(n1295), .B(n1196), .Z(n1104) );
INV_X1 U980 ( .A(G472), .ZN(n1196) );
NAND2_X1 U981 ( .A1(n1296), .A2(n1276), .ZN(n1295) );
XOR2_X1 U982 ( .A(n1297), .B(n1189), .Z(n1296) );
XNOR2_X1 U983 ( .A(n1298), .B(n1193), .ZN(n1189) );
XNOR2_X1 U984 ( .A(n1299), .B(n1300), .ZN(n1193) );
NOR2_X1 U985 ( .A1(n1301), .A2(n1302), .ZN(n1297) );
XNOR2_X1 U986 ( .A(KEYINPUT43), .B(n1198), .ZN(n1302) );
NAND4_X1 U987 ( .A1(G101), .A2(G210), .A3(n1303), .A4(n1145), .ZN(n1198) );
INV_X1 U988 ( .A(n1197), .ZN(n1301) );
NAND2_X1 U989 ( .A1(n1304), .A2(n1305), .ZN(n1197) );
NAND3_X1 U990 ( .A1(n1303), .A2(n1145), .A3(G210), .ZN(n1305) );
AND3_X1 U991 ( .A1(n1069), .A2(n1248), .A3(n1084), .ZN(n1057) );
INV_X1 U992 ( .A(n1266), .ZN(n1084) );
NAND2_X1 U993 ( .A1(n1085), .A2(n1086), .ZN(n1266) );
NAND2_X1 U994 ( .A1(G214), .A2(n1306), .ZN(n1086) );
XNOR2_X1 U995 ( .A(n1307), .B(n1308), .ZN(n1085) );
NOR2_X1 U996 ( .A1(n1224), .A2(n1225), .ZN(n1308) );
INV_X1 U997 ( .A(G210), .ZN(n1225) );
INV_X1 U998 ( .A(n1306), .ZN(n1224) );
NAND2_X1 U999 ( .A1(n1309), .A2(n1303), .ZN(n1306) );
NAND2_X1 U1000 ( .A1(n1310), .A2(n1276), .ZN(n1307) );
XOR2_X1 U1001 ( .A(n1311), .B(n1222), .Z(n1310) );
NAND3_X1 U1002 ( .A1(n1312), .A2(n1313), .A3(n1165), .ZN(n1222) );
OR2_X1 U1003 ( .A1(n1314), .A2(n1315), .ZN(n1165) );
NAND2_X1 U1004 ( .A1(n1316), .A2(n1317), .ZN(n1313) );
INV_X1 U1005 ( .A(KEYINPUT5), .ZN(n1317) );
XOR2_X1 U1006 ( .A(n1318), .B(n1315), .Z(n1316) );
NAND2_X1 U1007 ( .A1(KEYINPUT5), .A2(n1167), .ZN(n1312) );
NAND2_X1 U1008 ( .A1(n1319), .A2(n1320), .ZN(n1167) );
NAND3_X1 U1009 ( .A1(n1315), .A2(n1314), .A3(n1318), .ZN(n1320) );
NAND2_X1 U1010 ( .A1(n1298), .A2(n1321), .ZN(n1314) );
XNOR2_X1 U1011 ( .A(n1322), .B(n1323), .ZN(n1321) );
INV_X1 U1012 ( .A(n1192), .ZN(n1298) );
OR2_X1 U1013 ( .A1(n1318), .A2(n1315), .ZN(n1319) );
XNOR2_X1 U1014 ( .A(G122), .B(G110), .ZN(n1315) );
NAND2_X1 U1015 ( .A1(n1324), .A2(n1192), .ZN(n1318) );
XOR2_X1 U1016 ( .A(G113), .B(n1325), .Z(n1192) );
XOR2_X1 U1017 ( .A(G119), .B(G116), .Z(n1325) );
XOR2_X1 U1018 ( .A(n1322), .B(n1323), .Z(n1324) );
NAND2_X1 U1019 ( .A1(KEYINPUT6), .A2(n1304), .ZN(n1322) );
INV_X1 U1020 ( .A(G101), .ZN(n1304) );
NAND2_X1 U1021 ( .A1(n1326), .A2(n1327), .ZN(n1311) );
NAND2_X1 U1022 ( .A1(n1219), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1023 ( .A(KEYINPUT9), .B(n1329), .Z(n1326) );
NOR2_X1 U1024 ( .A1(n1219), .A2(n1328), .ZN(n1329) );
XNOR2_X1 U1025 ( .A(n1221), .B(KEYINPUT57), .ZN(n1328) );
INV_X1 U1026 ( .A(n1218), .ZN(n1221) );
NAND2_X1 U1027 ( .A1(G224), .A2(n1145), .ZN(n1218) );
XNOR2_X1 U1028 ( .A(n1299), .B(n1287), .ZN(n1219) );
INV_X1 U1029 ( .A(G125), .ZN(n1287) );
NAND2_X1 U1030 ( .A1(n1330), .A2(n1331), .ZN(n1299) );
NAND2_X1 U1031 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1032 ( .A(n1334), .B(KEYINPUT60), .Z(n1330) );
OR2_X1 U1033 ( .A1(n1333), .A2(n1332), .ZN(n1334) );
XOR2_X1 U1034 ( .A(n1335), .B(n1255), .Z(n1332) );
NAND2_X1 U1035 ( .A1(KEYINPUT42), .A2(n1279), .ZN(n1335) );
INV_X1 U1036 ( .A(G128), .ZN(n1333) );
NAND2_X1 U1037 ( .A1(n1078), .A2(n1336), .ZN(n1248) );
NAND4_X1 U1038 ( .A1(G953), .A2(G902), .A3(n1264), .A4(n1168), .ZN(n1336) );
INV_X1 U1039 ( .A(G898), .ZN(n1168) );
NAND3_X1 U1040 ( .A1(n1337), .A2(n1264), .A3(n1125), .ZN(n1078) );
XOR2_X1 U1041 ( .A(G953), .B(KEYINPUT61), .Z(n1125) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1264) );
XOR2_X1 U1043 ( .A(KEYINPUT52), .B(G952), .Z(n1337) );
AND2_X1 U1044 ( .A1(n1088), .A2(n1087), .ZN(n1069) );
NAND2_X1 U1045 ( .A1(G221), .A2(n1275), .ZN(n1087) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1309), .ZN(n1275) );
XNOR2_X1 U1047 ( .A(G902), .B(KEYINPUT28), .ZN(n1309) );
XOR2_X1 U1048 ( .A(n1338), .B(G469), .Z(n1088) );
NAND2_X1 U1049 ( .A1(KEYINPUT26), .A2(n1113), .ZN(n1338) );
NAND2_X1 U1050 ( .A1(n1339), .A2(n1276), .ZN(n1113) );
XOR2_X1 U1051 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1052 ( .A(KEYINPUT49), .B(n1209), .ZN(n1341) );
INV_X1 U1053 ( .A(G110), .ZN(n1209) );
XNOR2_X1 U1054 ( .A(n1205), .B(n1342), .ZN(n1340) );
NOR2_X1 U1055 ( .A1(KEYINPUT37), .A2(n1343), .ZN(n1342) );
XNOR2_X1 U1056 ( .A(n1344), .B(n1345), .ZN(n1205) );
XNOR2_X1 U1057 ( .A(n1300), .B(n1346), .ZN(n1345) );
XNOR2_X1 U1058 ( .A(G101), .B(n1347), .ZN(n1346) );
NOR2_X1 U1059 ( .A1(G953), .A2(n1148), .ZN(n1347) );
INV_X1 U1060 ( .A(G227), .ZN(n1148) );
XNOR2_X1 U1061 ( .A(n1348), .B(n1349), .ZN(n1300) );
NOR2_X1 U1062 ( .A1(KEYINPUT8), .A2(n1350), .ZN(n1349) );
NOR2_X1 U1063 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NOR2_X1 U1064 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NOR2_X1 U1065 ( .A1(n1355), .A2(KEYINPUT46), .ZN(n1353) );
NOR2_X1 U1066 ( .A1(KEYINPUT54), .A2(n1356), .ZN(n1355) );
INV_X1 U1067 ( .A(n1357), .ZN(n1356) );
NOR2_X1 U1068 ( .A1(n1358), .A2(n1357), .ZN(n1351) );
XOR2_X1 U1069 ( .A(G137), .B(KEYINPUT55), .Z(n1357) );
NOR2_X1 U1070 ( .A1(n1359), .A2(KEYINPUT54), .ZN(n1358) );
NOR2_X1 U1071 ( .A1(KEYINPUT46), .A2(G134), .ZN(n1359) );
XNOR2_X1 U1072 ( .A(G131), .B(KEYINPUT24), .ZN(n1348) );
XNOR2_X1 U1073 ( .A(n1323), .B(n1144), .ZN(n1344) );
XOR2_X1 U1074 ( .A(n1360), .B(n1279), .Z(n1144) );
XNOR2_X1 U1075 ( .A(G107), .B(n1361), .ZN(n1323) );
NOR2_X1 U1076 ( .A1(n1120), .A2(n1254), .ZN(n1100) );
XOR2_X1 U1077 ( .A(n1123), .B(n1122), .Z(n1254) );
INV_X1 U1078 ( .A(G475), .ZN(n1122) );
NAND2_X1 U1079 ( .A1(n1182), .A2(n1276), .ZN(n1123) );
XOR2_X1 U1080 ( .A(n1362), .B(n1363), .Z(n1182) );
XOR2_X1 U1081 ( .A(n1364), .B(n1365), .Z(n1363) );
NAND2_X1 U1082 ( .A1(KEYINPUT0), .A2(n1143), .ZN(n1365) );
INV_X1 U1083 ( .A(G131), .ZN(n1143) );
NAND3_X1 U1084 ( .A1(n1303), .A2(n1145), .A3(G214), .ZN(n1364) );
INV_X1 U1085 ( .A(G237), .ZN(n1303) );
XOR2_X1 U1086 ( .A(n1366), .B(n1367), .Z(n1362) );
NOR2_X1 U1087 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
XOR2_X1 U1088 ( .A(KEYINPUT48), .B(n1370), .Z(n1369) );
NOR2_X1 U1089 ( .A1(n1361), .A2(n1371), .ZN(n1370) );
AND2_X1 U1090 ( .A1(n1361), .A2(n1371), .ZN(n1368) );
XOR2_X1 U1091 ( .A(G122), .B(n1372), .Z(n1371) );
NOR2_X1 U1092 ( .A1(G113), .A2(KEYINPUT15), .ZN(n1372) );
INV_X1 U1093 ( .A(G104), .ZN(n1361) );
XNOR2_X1 U1094 ( .A(n1373), .B(n1255), .ZN(n1366) );
NAND3_X1 U1095 ( .A1(n1374), .A2(n1375), .A3(n1376), .ZN(n1373) );
OR2_X1 U1096 ( .A1(n1377), .A2(n1279), .ZN(n1376) );
NAND3_X1 U1097 ( .A1(n1279), .A2(n1377), .A3(n1134), .ZN(n1375) );
NAND2_X1 U1098 ( .A1(n1378), .A2(n1379), .ZN(n1374) );
NAND2_X1 U1099 ( .A1(n1380), .A2(n1377), .ZN(n1379) );
INV_X1 U1100 ( .A(KEYINPUT50), .ZN(n1377) );
XNOR2_X1 U1101 ( .A(n1279), .B(KEYINPUT38), .ZN(n1380) );
XOR2_X1 U1102 ( .A(G146), .B(KEYINPUT51), .Z(n1279) );
INV_X1 U1103 ( .A(n1134), .ZN(n1378) );
XNOR2_X1 U1104 ( .A(G125), .B(n1208), .ZN(n1134) );
INV_X1 U1105 ( .A(n1343), .ZN(n1208) );
XOR2_X1 U1106 ( .A(G140), .B(KEYINPUT12), .Z(n1343) );
XOR2_X1 U1107 ( .A(n1381), .B(n1178), .Z(n1120) );
INV_X1 U1108 ( .A(G478), .ZN(n1178) );
NAND2_X1 U1109 ( .A1(n1176), .A2(n1276), .ZN(n1381) );
INV_X1 U1110 ( .A(G902), .ZN(n1276) );
XNOR2_X1 U1111 ( .A(n1382), .B(n1383), .ZN(n1176) );
AND2_X1 U1112 ( .A1(n1294), .A2(G217), .ZN(n1383) );
AND2_X1 U1113 ( .A1(G234), .A2(n1145), .ZN(n1294) );
INV_X1 U1114 ( .A(G953), .ZN(n1145) );
NAND2_X1 U1115 ( .A1(n1384), .A2(KEYINPUT21), .ZN(n1382) );
XOR2_X1 U1116 ( .A(n1385), .B(n1386), .Z(n1384) );
XOR2_X1 U1117 ( .A(G116), .B(n1387), .Z(n1386) );
XNOR2_X1 U1118 ( .A(n1354), .B(G122), .ZN(n1387) );
INV_X1 U1119 ( .A(G134), .ZN(n1354) );
XOR2_X1 U1120 ( .A(n1388), .B(n1360), .Z(n1385) );
XNOR2_X1 U1121 ( .A(G128), .B(n1255), .ZN(n1360) );
INV_X1 U1122 ( .A(G143), .ZN(n1255) );
NAND2_X1 U1123 ( .A1(KEYINPUT17), .A2(n1389), .ZN(n1388) );
INV_X1 U1124 ( .A(G107), .ZN(n1389) );
endmodule


