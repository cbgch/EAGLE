//Key = 0101101001010011000110000010010000010110010100100100010001001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241;

XOR2_X1 U688 ( .A(n947), .B(n948), .Z(G9) );
NOR2_X1 U689 ( .A1(n949), .A2(n950), .ZN(n948) );
INV_X1 U690 ( .A(G107), .ZN(n950) );
XNOR2_X1 U691 ( .A(KEYINPUT53), .B(KEYINPUT24), .ZN(n949) );
NOR2_X1 U692 ( .A1(n951), .A2(n952), .ZN(G75) );
NOR4_X1 U693 ( .A1(G953), .A2(n953), .A3(n954), .A4(n955), .ZN(n952) );
NOR2_X1 U694 ( .A1(n956), .A2(n957), .ZN(n954) );
NOR2_X1 U695 ( .A1(n958), .A2(n959), .ZN(n956) );
NOR2_X1 U696 ( .A1(n960), .A2(n961), .ZN(n959) );
NOR2_X1 U697 ( .A1(n962), .A2(n963), .ZN(n960) );
AND2_X1 U698 ( .A1(n964), .A2(n965), .ZN(n963) );
NOR3_X1 U699 ( .A1(n966), .A2(n967), .A3(n968), .ZN(n962) );
NOR2_X1 U700 ( .A1(n969), .A2(n970), .ZN(n968) );
AND2_X1 U701 ( .A1(n971), .A2(n964), .ZN(n970) );
NOR3_X1 U702 ( .A1(n972), .A2(n973), .A3(n974), .ZN(n969) );
NOR3_X1 U703 ( .A1(n975), .A2(n976), .A3(n977), .ZN(n974) );
NOR2_X1 U704 ( .A1(n964), .A2(n978), .ZN(n973) );
NOR4_X1 U705 ( .A1(n979), .A2(n972), .A3(n975), .A4(n980), .ZN(n958) );
NAND3_X1 U706 ( .A1(n981), .A2(n982), .A3(n983), .ZN(n979) );
NAND2_X1 U707 ( .A1(n967), .A2(n961), .ZN(n982) );
INV_X1 U708 ( .A(n984), .ZN(n961) );
OR3_X1 U709 ( .A1(n985), .A2(n986), .A3(n967), .ZN(n981) );
NOR3_X1 U710 ( .A1(n953), .A2(G953), .A3(G952), .ZN(n951) );
AND4_X1 U711 ( .A1(n987), .A2(n988), .A3(n989), .A4(n990), .ZN(n953) );
NOR4_X1 U712 ( .A1(n991), .A2(n980), .A3(n992), .A4(n993), .ZN(n990) );
XOR2_X1 U713 ( .A(n994), .B(n995), .Z(n993) );
XNOR2_X1 U714 ( .A(G469), .B(KEYINPUT23), .ZN(n995) );
INV_X1 U715 ( .A(n964), .ZN(n980) );
XOR2_X1 U716 ( .A(n996), .B(KEYINPUT3), .Z(n991) );
NOR2_X1 U717 ( .A1(n967), .A2(n975), .ZN(n989) );
INV_X1 U718 ( .A(n997), .ZN(n967) );
NAND2_X1 U719 ( .A1(n998), .A2(n999), .ZN(n988) );
XOR2_X1 U720 ( .A(KEYINPUT41), .B(n1000), .Z(n987) );
NOR2_X1 U721 ( .A1(n998), .A2(n999), .ZN(n1000) );
XOR2_X1 U722 ( .A(n1001), .B(n1002), .Z(G72) );
NOR2_X1 U723 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
XOR2_X1 U724 ( .A(n1005), .B(n1006), .Z(n1004) );
XOR2_X1 U725 ( .A(n1007), .B(n1008), .Z(n1006) );
XOR2_X1 U726 ( .A(G131), .B(G125), .Z(n1008) );
XOR2_X1 U727 ( .A(n1009), .B(n1010), .Z(n1005) );
XOR2_X1 U728 ( .A(G137), .B(G134), .Z(n1010) );
XOR2_X1 U729 ( .A(KEYINPUT44), .B(G140), .Z(n1009) );
INV_X1 U730 ( .A(n1011), .ZN(n1003) );
NAND2_X1 U731 ( .A1(n1012), .A2(n1013), .ZN(n1001) );
NAND2_X1 U732 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
XOR2_X1 U733 ( .A(n1016), .B(KEYINPUT2), .Z(n1014) );
NAND2_X1 U734 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U735 ( .A1(KEYINPUT49), .A2(n1019), .ZN(n1012) );
NAND2_X1 U736 ( .A1(n1011), .A2(n1020), .ZN(n1019) );
NAND2_X1 U737 ( .A1(G953), .A2(n1021), .ZN(n1020) );
XOR2_X1 U738 ( .A(KEYINPUT37), .B(G227), .Z(n1021) );
NAND2_X1 U739 ( .A1(G953), .A2(n1022), .ZN(n1011) );
XOR2_X1 U740 ( .A(n1023), .B(n1024), .Z(G69) );
NOR2_X1 U741 ( .A1(n1025), .A2(n1015), .ZN(n1024) );
AND2_X1 U742 ( .A1(G224), .A2(G898), .ZN(n1025) );
NAND2_X1 U743 ( .A1(n1026), .A2(n1027), .ZN(n1023) );
NAND2_X1 U744 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
XOR2_X1 U745 ( .A(n1030), .B(KEYINPUT62), .Z(n1028) );
NAND2_X1 U746 ( .A1(n1031), .A2(n1015), .ZN(n1030) );
OR3_X1 U747 ( .A1(n1031), .A2(n1032), .A3(n1029), .ZN(n1026) );
XOR2_X1 U748 ( .A(n1033), .B(n1034), .Z(n1031) );
XOR2_X1 U749 ( .A(G119), .B(n1035), .Z(n1034) );
NOR2_X1 U750 ( .A1(n1036), .A2(n1037), .ZN(G66) );
XOR2_X1 U751 ( .A(n1038), .B(n1039), .Z(n1037) );
NOR2_X1 U752 ( .A1(KEYINPUT40), .A2(n1040), .ZN(n1039) );
XOR2_X1 U753 ( .A(n1041), .B(n1042), .Z(n1040) );
NAND2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1038) );
NOR2_X1 U755 ( .A1(n1036), .A2(n1045), .ZN(G63) );
XNOR2_X1 U756 ( .A(n1046), .B(n1047), .ZN(n1045) );
AND2_X1 U757 ( .A1(G478), .A2(n1043), .ZN(n1047) );
NOR2_X1 U758 ( .A1(n1036), .A2(n1048), .ZN(G60) );
NOR3_X1 U759 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
AND3_X1 U760 ( .A1(n1052), .A2(G475), .A3(n1043), .ZN(n1051) );
NOR2_X1 U761 ( .A1(n1053), .A2(n1052), .ZN(n1050) );
AND2_X1 U762 ( .A1(n955), .A2(G475), .ZN(n1053) );
XOR2_X1 U763 ( .A(G104), .B(n1054), .Z(G6) );
NOR3_X1 U764 ( .A1(n1036), .A2(n1055), .A3(n1056), .ZN(G57) );
NOR2_X1 U765 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR3_X1 U767 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
AND2_X1 U768 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
INV_X1 U769 ( .A(KEYINPUT29), .ZN(n1061) );
INV_X1 U770 ( .A(n1064), .ZN(n1057) );
NOR2_X1 U771 ( .A1(n1065), .A2(n1064), .ZN(n1055) );
NOR2_X1 U772 ( .A1(n1062), .A2(n1063), .ZN(n1065) );
INV_X1 U773 ( .A(KEYINPUT35), .ZN(n1063) );
NAND3_X1 U774 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1062) );
NAND2_X1 U775 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND3_X1 U776 ( .A1(n1043), .A2(G472), .A3(KEYINPUT38), .ZN(n1070) );
XNOR2_X1 U777 ( .A(KEYINPUT7), .B(n1071), .ZN(n1069) );
NAND2_X1 U778 ( .A1(KEYINPUT33), .A2(n1072), .ZN(n1067) );
NAND2_X1 U779 ( .A1(n1043), .A2(G472), .ZN(n1072) );
NAND4_X1 U780 ( .A1(n1073), .A2(G472), .A3(n1074), .A4(n1075), .ZN(n1066) );
INV_X1 U781 ( .A(KEYINPUT33), .ZN(n1075) );
AND2_X1 U782 ( .A1(n1043), .A2(KEYINPUT38), .ZN(n1074) );
XOR2_X1 U783 ( .A(KEYINPUT7), .B(n1071), .Z(n1073) );
NOR2_X1 U784 ( .A1(n1036), .A2(n1076), .ZN(G54) );
XOR2_X1 U785 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND2_X1 U786 ( .A1(n1043), .A2(G469), .ZN(n1078) );
INV_X1 U787 ( .A(n1079), .ZN(n1043) );
NAND2_X1 U788 ( .A1(n1080), .A2(KEYINPUT46), .ZN(n1077) );
XOR2_X1 U789 ( .A(n1081), .B(n1082), .Z(n1080) );
XOR2_X1 U790 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U791 ( .A(n1085), .B(n1086), .Z(n1081) );
NOR2_X1 U792 ( .A1(n1087), .A2(KEYINPUT58), .ZN(n1086) );
NOR2_X1 U793 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U794 ( .A(n1090), .B(KEYINPUT19), .Z(n1089) );
NAND2_X1 U795 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U796 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
INV_X1 U797 ( .A(n1093), .ZN(n1092) );
XNOR2_X1 U798 ( .A(n1094), .B(n1095), .ZN(n1091) );
XOR2_X1 U799 ( .A(n1096), .B(KEYINPUT17), .Z(n1094) );
INV_X1 U800 ( .A(G110), .ZN(n1085) );
NOR2_X1 U801 ( .A1(n1036), .A2(n1097), .ZN(G51) );
XOR2_X1 U802 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U803 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U804 ( .A1(G125), .A2(KEYINPUT32), .ZN(n1101) );
NOR2_X1 U805 ( .A1(n1102), .A2(n1079), .ZN(n1100) );
NAND2_X1 U806 ( .A1(G902), .A2(n955), .ZN(n1079) );
NAND3_X1 U807 ( .A1(n1103), .A2(n1104), .A3(n1017), .ZN(n955) );
AND4_X1 U808 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1017) );
NOR4_X1 U809 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
INV_X1 U810 ( .A(n1113), .ZN(n1109) );
NAND3_X1 U811 ( .A1(n1114), .A2(n971), .A3(n1115), .ZN(n1107) );
XNOR2_X1 U812 ( .A(KEYINPUT11), .B(n1018), .ZN(n1104) );
INV_X1 U813 ( .A(n1029), .ZN(n1103) );
NAND4_X1 U814 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1029) );
NOR4_X1 U815 ( .A1(n1120), .A2(n1121), .A3(n1054), .A4(n1122), .ZN(n1119) );
NOR2_X1 U816 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
AND3_X1 U817 ( .A1(n1125), .A2(n964), .A3(n986), .ZN(n1054) );
NOR2_X1 U818 ( .A1(n947), .A2(n1126), .ZN(n1118) );
AND3_X1 U819 ( .A1(n985), .A2(n964), .A3(n1125), .ZN(n947) );
NOR2_X1 U820 ( .A1(n1015), .A2(G952), .ZN(n1036) );
XOR2_X1 U821 ( .A(n1127), .B(n1105), .Z(G48) );
NAND3_X1 U822 ( .A1(n986), .A2(n971), .A3(n1128), .ZN(n1105) );
XNOR2_X1 U823 ( .A(G143), .B(n1129), .ZN(G45) );
NAND3_X1 U824 ( .A1(n1115), .A2(n1130), .A3(n1131), .ZN(n1129) );
XOR2_X1 U825 ( .A(n1132), .B(KEYINPUT20), .Z(n1131) );
XOR2_X1 U826 ( .A(KEYINPUT8), .B(n971), .Z(n1130) );
AND4_X1 U827 ( .A1(n1133), .A2(n976), .A3(n992), .A4(n1134), .ZN(n1115) );
NAND2_X1 U828 ( .A1(n1135), .A2(n1136), .ZN(G42) );
NAND2_X1 U829 ( .A1(G140), .A2(n1106), .ZN(n1136) );
XOR2_X1 U830 ( .A(KEYINPUT9), .B(n1137), .Z(n1135) );
NOR2_X1 U831 ( .A1(G140), .A2(n1106), .ZN(n1137) );
NAND3_X1 U832 ( .A1(n986), .A2(n977), .A3(n1138), .ZN(n1106) );
XOR2_X1 U833 ( .A(G137), .B(n1112), .Z(G39) );
AND4_X1 U834 ( .A1(n984), .A2(n1128), .A3(n996), .A4(n978), .ZN(n1112) );
XOR2_X1 U835 ( .A(n1018), .B(n1139), .Z(G36) );
NAND2_X1 U836 ( .A1(KEYINPUT6), .A2(G134), .ZN(n1139) );
NAND3_X1 U837 ( .A1(n976), .A2(n985), .A3(n1138), .ZN(n1018) );
XOR2_X1 U838 ( .A(G131), .B(n1111), .Z(G33) );
AND3_X1 U839 ( .A1(n976), .A2(n986), .A3(n1138), .ZN(n1111) );
AND2_X1 U840 ( .A1(n965), .A2(n1134), .ZN(n1138) );
NOR3_X1 U841 ( .A1(n1132), .A2(n975), .A3(n972), .ZN(n965) );
INV_X1 U842 ( .A(n978), .ZN(n975) );
XOR2_X1 U843 ( .A(G128), .B(n1110), .Z(G30) );
AND3_X1 U844 ( .A1(n985), .A2(n971), .A3(n1128), .ZN(n1110) );
AND4_X1 U845 ( .A1(n1114), .A2(n1140), .A3(n1141), .A4(n1134), .ZN(n1128) );
XOR2_X1 U846 ( .A(G101), .B(n1121), .Z(G3) );
AND3_X1 U847 ( .A1(n976), .A2(n1125), .A3(n984), .ZN(n1121) );
XOR2_X1 U848 ( .A(G125), .B(n1142), .Z(G27) );
NOR2_X1 U849 ( .A1(KEYINPUT59), .A2(n1113), .ZN(n1142) );
NAND4_X1 U850 ( .A1(n1134), .A2(n997), .A3(n971), .A4(n1143), .ZN(n1113) );
AND3_X1 U851 ( .A1(n986), .A2(n977), .A3(n983), .ZN(n1143) );
NAND2_X1 U852 ( .A1(n957), .A2(n1144), .ZN(n1134) );
NAND4_X1 U853 ( .A1(G902), .A2(n1145), .A3(n1146), .A4(n1022), .ZN(n1144) );
INV_X1 U854 ( .A(G900), .ZN(n1022) );
XOR2_X1 U855 ( .A(KEYINPUT12), .B(G953), .Z(n1145) );
XOR2_X1 U856 ( .A(G122), .B(n1120), .Z(G24) );
AND4_X1 U857 ( .A1(n1133), .A2(n1147), .A3(n964), .A4(n992), .ZN(n1120) );
NOR2_X1 U858 ( .A1(n1141), .A2(n1140), .ZN(n964) );
NAND2_X1 U859 ( .A1(n1148), .A2(n1149), .ZN(G21) );
OR2_X1 U860 ( .A1(n1116), .A2(G119), .ZN(n1149) );
XOR2_X1 U861 ( .A(n1150), .B(KEYINPUT22), .Z(n1148) );
NAND2_X1 U862 ( .A1(G119), .A2(n1116), .ZN(n1150) );
NAND4_X1 U863 ( .A1(n1147), .A2(n984), .A3(n1140), .A4(n1141), .ZN(n1116) );
INV_X1 U864 ( .A(n1151), .ZN(n1140) );
XNOR2_X1 U865 ( .A(G116), .B(n1117), .ZN(G18) );
NAND3_X1 U866 ( .A1(n976), .A2(n985), .A3(n1147), .ZN(n1117) );
AND2_X1 U867 ( .A1(n1152), .A2(n971), .ZN(n1147) );
XNOR2_X1 U868 ( .A(n1123), .B(KEYINPUT48), .ZN(n971) );
NOR2_X1 U869 ( .A1(n1133), .A2(n1153), .ZN(n985) );
XOR2_X1 U870 ( .A(G113), .B(n1154), .Z(G15) );
NOR2_X1 U871 ( .A1(n1155), .A2(n1123), .ZN(n1154) );
XOR2_X1 U872 ( .A(n1124), .B(KEYINPUT13), .Z(n1155) );
NAND3_X1 U873 ( .A1(n976), .A2(n986), .A3(n1152), .ZN(n1124) );
AND3_X1 U874 ( .A1(n1156), .A2(n997), .A3(n983), .ZN(n1152) );
AND2_X1 U875 ( .A1(n1133), .A2(n1153), .ZN(n986) );
NOR2_X1 U876 ( .A1(n1141), .A2(n1151), .ZN(n976) );
XOR2_X1 U877 ( .A(n1126), .B(n1157), .Z(G12) );
XOR2_X1 U878 ( .A(KEYINPUT10), .B(G110), .Z(n1157) );
AND3_X1 U879 ( .A1(n977), .A2(n1125), .A3(n984), .ZN(n1126) );
NOR2_X1 U880 ( .A1(n992), .A2(n1133), .ZN(n984) );
XOR2_X1 U881 ( .A(n999), .B(n1158), .Z(n1133) );
NOR2_X1 U882 ( .A1(n1159), .A2(n998), .ZN(n1158) );
XOR2_X1 U883 ( .A(G475), .B(KEYINPUT55), .Z(n998) );
XNOR2_X1 U884 ( .A(KEYINPUT56), .B(KEYINPUT14), .ZN(n1159) );
INV_X1 U885 ( .A(n1049), .ZN(n999) );
NOR2_X1 U886 ( .A1(n1052), .A2(G902), .ZN(n1049) );
XOR2_X1 U887 ( .A(n1160), .B(n1161), .Z(n1052) );
XOR2_X1 U888 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U889 ( .A(G113), .B(G104), .Z(n1163) );
XOR2_X1 U890 ( .A(G131), .B(G122), .Z(n1162) );
XOR2_X1 U891 ( .A(n1164), .B(n1165), .Z(n1160) );
XOR2_X1 U892 ( .A(n1166), .B(n1167), .Z(n1165) );
AND2_X1 U893 ( .A1(G214), .A2(n1168), .ZN(n1167) );
NOR2_X1 U894 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
XOR2_X1 U895 ( .A(n1171), .B(KEYINPUT4), .Z(n1170) );
NAND2_X1 U896 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U897 ( .A(KEYINPUT43), .B(G146), .Z(n1172) );
NOR2_X1 U898 ( .A1(n1127), .A2(n1173), .ZN(n1169) );
XNOR2_X1 U899 ( .A(G125), .B(n1174), .ZN(n1173) );
NAND2_X1 U900 ( .A1(n1175), .A2(KEYINPUT61), .ZN(n1174) );
XNOR2_X1 U901 ( .A(n1176), .B(KEYINPUT42), .ZN(n1175) );
NAND2_X1 U902 ( .A1(KEYINPUT26), .A2(n1177), .ZN(n1164) );
INV_X1 U903 ( .A(n1153), .ZN(n992) );
XOR2_X1 U904 ( .A(n1178), .B(G478), .Z(n1153) );
NAND2_X1 U905 ( .A1(n1046), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U906 ( .A(n1180), .B(n1181), .ZN(n1046) );
AND2_X1 U907 ( .A1(n1182), .A2(G217), .ZN(n1181) );
NAND2_X1 U908 ( .A1(KEYINPUT15), .A2(n1183), .ZN(n1180) );
XOR2_X1 U909 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U910 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U911 ( .A(G107), .B(n1188), .Z(n1187) );
NOR2_X1 U912 ( .A1(KEYINPUT39), .A2(n1177), .ZN(n1188) );
NOR2_X1 U913 ( .A1(G134), .A2(KEYINPUT21), .ZN(n1186) );
XOR2_X1 U914 ( .A(n1189), .B(n1190), .Z(n1184) );
XOR2_X1 U915 ( .A(G122), .B(G116), .Z(n1190) );
XOR2_X1 U916 ( .A(KEYINPUT51), .B(G128), .Z(n1189) );
AND3_X1 U917 ( .A1(n1114), .A2(n1156), .A3(n1191), .ZN(n1125) );
INV_X1 U918 ( .A(n1123), .ZN(n1191) );
NAND2_X1 U919 ( .A1(n972), .A2(n978), .ZN(n1123) );
NAND2_X1 U920 ( .A1(n1192), .A2(n1193), .ZN(n978) );
XNOR2_X1 U921 ( .A(G214), .B(KEYINPUT1), .ZN(n1192) );
INV_X1 U922 ( .A(n996), .ZN(n972) );
XNOR2_X1 U923 ( .A(n1194), .B(n1102), .ZN(n996) );
NAND2_X1 U924 ( .A1(G210), .A2(n1193), .ZN(n1102) );
NAND2_X1 U925 ( .A1(n1195), .A2(n1179), .ZN(n1193) );
INV_X1 U926 ( .A(G237), .ZN(n1195) );
NAND2_X1 U927 ( .A1(n1196), .A2(n1179), .ZN(n1194) );
XOR2_X1 U928 ( .A(G125), .B(n1098), .Z(n1196) );
XNOR2_X1 U929 ( .A(n1033), .B(n1197), .ZN(n1098) );
XOR2_X1 U930 ( .A(n1198), .B(n1199), .Z(n1197) );
AND2_X1 U931 ( .A1(n1015), .A2(G224), .ZN(n1198) );
XOR2_X1 U932 ( .A(n1200), .B(n1201), .Z(n1033) );
XNOR2_X1 U933 ( .A(G122), .B(n1202), .ZN(n1201) );
NAND2_X1 U934 ( .A1(KEYINPUT60), .A2(n1203), .ZN(n1202) );
INV_X1 U935 ( .A(G104), .ZN(n1203) );
NAND2_X1 U936 ( .A1(n957), .A2(n1204), .ZN(n1156) );
NAND3_X1 U937 ( .A1(n1032), .A2(n1146), .A3(G902), .ZN(n1204) );
NOR2_X1 U938 ( .A1(n1015), .A2(G898), .ZN(n1032) );
NAND3_X1 U939 ( .A1(n1146), .A2(n1015), .A3(G952), .ZN(n957) );
NAND2_X1 U940 ( .A1(G237), .A2(G234), .ZN(n1146) );
INV_X1 U941 ( .A(n1132), .ZN(n1114) );
NAND2_X1 U942 ( .A1(n966), .A2(n997), .ZN(n1132) );
NAND2_X1 U943 ( .A1(G221), .A2(n1205), .ZN(n997) );
INV_X1 U944 ( .A(n983), .ZN(n966) );
XNOR2_X1 U945 ( .A(G469), .B(n1206), .ZN(n983) );
NOR2_X1 U946 ( .A1(KEYINPUT27), .A2(n994), .ZN(n1206) );
NAND2_X1 U947 ( .A1(n1207), .A2(n1179), .ZN(n994) );
XOR2_X1 U948 ( .A(n1208), .B(n1209), .Z(n1207) );
XNOR2_X1 U949 ( .A(n1083), .B(n1210), .ZN(n1209) );
XNOR2_X1 U950 ( .A(KEYINPUT30), .B(n1211), .ZN(n1210) );
NOR2_X1 U951 ( .A1(KEYINPUT0), .A2(n1093), .ZN(n1211) );
XNOR2_X1 U952 ( .A(n1007), .B(KEYINPUT28), .ZN(n1093) );
XNOR2_X1 U953 ( .A(n1212), .B(n1213), .ZN(n1007) );
INV_X1 U954 ( .A(G128), .ZN(n1212) );
XOR2_X1 U955 ( .A(n1214), .B(n1084), .Z(n1208) );
XOR2_X1 U956 ( .A(G140), .B(n1215), .Z(n1084) );
AND2_X1 U957 ( .A1(n1015), .A2(G227), .ZN(n1215) );
XOR2_X1 U958 ( .A(n1200), .B(n1095), .Z(n1214) );
XOR2_X1 U959 ( .A(G104), .B(KEYINPUT5), .Z(n1095) );
XOR2_X1 U960 ( .A(n1096), .B(G110), .Z(n1200) );
XOR2_X1 U961 ( .A(n1216), .B(n1217), .Z(n1096) );
XOR2_X1 U962 ( .A(KEYINPUT16), .B(G107), .Z(n1217) );
INV_X1 U963 ( .A(G101), .ZN(n1216) );
AND2_X1 U964 ( .A1(n1151), .A2(n1141), .ZN(n977) );
XNOR2_X1 U965 ( .A(n1218), .B(n1044), .ZN(n1141) );
AND2_X1 U966 ( .A1(G217), .A2(n1205), .ZN(n1044) );
NAND2_X1 U967 ( .A1(n1219), .A2(n1179), .ZN(n1205) );
XOR2_X1 U968 ( .A(KEYINPUT18), .B(G234), .Z(n1219) );
NAND2_X1 U969 ( .A1(n1220), .A2(n1179), .ZN(n1218) );
XNOR2_X1 U970 ( .A(n1041), .B(n1042), .ZN(n1220) );
XNOR2_X1 U971 ( .A(n1221), .B(G137), .ZN(n1042) );
NAND2_X1 U972 ( .A1(n1182), .A2(G221), .ZN(n1221) );
AND2_X1 U973 ( .A1(G234), .A2(n1015), .ZN(n1182) );
INV_X1 U974 ( .A(G953), .ZN(n1015) );
NAND2_X1 U975 ( .A1(KEYINPUT57), .A2(n1222), .ZN(n1041) );
XOR2_X1 U976 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U977 ( .A(G110), .B(n1225), .Z(n1224) );
NOR2_X1 U978 ( .A1(KEYINPUT31), .A2(n1226), .ZN(n1225) );
XOR2_X1 U979 ( .A(n1227), .B(n1228), .Z(n1226) );
XOR2_X1 U980 ( .A(n1127), .B(n1229), .Z(n1228) );
XNOR2_X1 U981 ( .A(KEYINPUT47), .B(KEYINPUT36), .ZN(n1229) );
XNOR2_X1 U982 ( .A(G125), .B(n1176), .ZN(n1227) );
XOR2_X1 U983 ( .A(G140), .B(KEYINPUT25), .Z(n1176) );
XOR2_X1 U984 ( .A(n1230), .B(G472), .Z(n1151) );
NAND2_X1 U985 ( .A1(n1231), .A2(n1179), .ZN(n1230) );
INV_X1 U986 ( .A(G902), .ZN(n1179) );
XOR2_X1 U987 ( .A(n1064), .B(n1071), .Z(n1231) );
XOR2_X1 U988 ( .A(n1232), .B(n1199), .Z(n1071) );
XNOR2_X1 U989 ( .A(n1233), .B(n1223), .ZN(n1199) );
XOR2_X1 U990 ( .A(G119), .B(G128), .Z(n1223) );
XNOR2_X1 U991 ( .A(n1035), .B(n1234), .ZN(n1233) );
NOR2_X1 U992 ( .A1(KEYINPUT50), .A2(n1213), .ZN(n1234) );
XNOR2_X1 U993 ( .A(n1235), .B(n1177), .ZN(n1213) );
XOR2_X1 U994 ( .A(G143), .B(KEYINPUT34), .Z(n1177) );
XOR2_X1 U995 ( .A(n1127), .B(KEYINPUT45), .Z(n1235) );
INV_X1 U996 ( .A(G146), .ZN(n1127) );
XOR2_X1 U997 ( .A(G113), .B(G116), .Z(n1035) );
XNOR2_X1 U998 ( .A(n1083), .B(KEYINPUT63), .ZN(n1232) );
XNOR2_X1 U999 ( .A(n1236), .B(n1237), .ZN(n1083) );
NOR2_X1 U1000 ( .A1(KEYINPUT52), .A2(n1238), .ZN(n1237) );
INV_X1 U1001 ( .A(G134), .ZN(n1238) );
XOR2_X1 U1002 ( .A(n1239), .B(n1240), .Z(n1236) );
NOR2_X1 U1003 ( .A1(G131), .A2(KEYINPUT54), .ZN(n1240) );
INV_X1 U1004 ( .A(G137), .ZN(n1239) );
XOR2_X1 U1005 ( .A(n1241), .B(G101), .Z(n1064) );
NAND2_X1 U1006 ( .A1(n1168), .A2(G210), .ZN(n1241) );
NOR2_X1 U1007 ( .A1(G953), .A2(G237), .ZN(n1168) );
endmodule


