//Key = 0000101101010011011111111101101110101010010011001100010100010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350;

XOR2_X1 U737 ( .A(n1024), .B(n1025), .Z(G9) );
NAND3_X1 U738 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(G75) );
NAND2_X1 U739 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NAND2_X1 U740 ( .A1(G952), .A2(n1031), .ZN(n1026) );
NAND3_X1 U741 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NOR3_X1 U742 ( .A1(n1035), .A2(G953), .A3(n1036), .ZN(n1034) );
NOR2_X1 U743 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U744 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR3_X1 U745 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR3_X1 U746 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1042) );
AND3_X1 U747 ( .A1(n1047), .A2(n1048), .A3(KEYINPUT0), .ZN(n1046) );
NOR2_X1 U748 ( .A1(n1049), .A2(n1047), .ZN(n1045) );
NOR3_X1 U749 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NOR2_X1 U750 ( .A1(KEYINPUT0), .A2(n1053), .ZN(n1052) );
AND2_X1 U751 ( .A1(n1054), .A2(KEYINPUT60), .ZN(n1051) );
NOR2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U754 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR3_X1 U755 ( .A1(n1047), .A2(n1061), .A3(n1056), .ZN(n1039) );
NOR2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U757 ( .A1(n1064), .A2(n1043), .ZN(n1063) );
NOR2_X1 U758 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
AND2_X1 U759 ( .A1(n1067), .A2(KEYINPUT21), .ZN(n1066) );
NOR3_X1 U760 ( .A1(n1068), .A2(KEYINPUT60), .A3(n1069), .ZN(n1065) );
NOR2_X1 U761 ( .A1(n1070), .A2(n1041), .ZN(n1062) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U763 ( .A1(KEYINPUT21), .A2(n1073), .ZN(n1035) );
NOR4_X1 U764 ( .A1(n1074), .A2(n1047), .A3(n1075), .A4(n1056), .ZN(n1073) );
INV_X1 U765 ( .A(n1054), .ZN(n1056) );
OR2_X1 U766 ( .A1(n1038), .A2(n1043), .ZN(n1074) );
INV_X1 U767 ( .A(n1076), .ZN(n1033) );
XNOR2_X1 U768 ( .A(n1029), .B(KEYINPUT40), .ZN(n1032) );
AND4_X1 U769 ( .A1(n1077), .A2(n1060), .A3(n1078), .A4(n1079), .ZN(n1029) );
NOR4_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1079) );
XOR2_X1 U771 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U772 ( .A(G469), .B(KEYINPUT50), .ZN(n1085) );
XOR2_X1 U773 ( .A(n1086), .B(n1087), .Z(n1082) );
XOR2_X1 U774 ( .A(n1088), .B(KEYINPUT32), .Z(n1087) );
NAND2_X1 U775 ( .A1(KEYINPUT30), .A2(n1089), .ZN(n1086) );
NOR3_X1 U776 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1078) );
XNOR2_X1 U777 ( .A(n1093), .B(n1094), .ZN(n1077) );
XOR2_X1 U778 ( .A(n1095), .B(KEYINPUT31), .Z(n1094) );
XOR2_X1 U779 ( .A(n1096), .B(n1097), .Z(G72) );
XOR2_X1 U780 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U781 ( .A1(G953), .A2(n1100), .ZN(n1099) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1100) );
NAND3_X1 U783 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1098) );
XOR2_X1 U784 ( .A(n1104), .B(KEYINPUT52), .Z(n1103) );
NAND2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
OR2_X1 U786 ( .A1(n1106), .A2(n1105), .ZN(n1102) );
XOR2_X1 U787 ( .A(G125), .B(n1107), .Z(n1105) );
XOR2_X1 U788 ( .A(KEYINPUT4), .B(G140), .Z(n1107) );
XNOR2_X1 U789 ( .A(n1108), .B(n1109), .ZN(n1106) );
XNOR2_X1 U790 ( .A(G131), .B(n1110), .ZN(n1109) );
NAND2_X1 U791 ( .A1(G953), .A2(n1111), .ZN(n1101) );
NOR2_X1 U792 ( .A1(n1112), .A2(G953), .ZN(n1096) );
XOR2_X1 U793 ( .A(n1113), .B(n1114), .Z(G69) );
XOR2_X1 U794 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U795 ( .A1(G953), .A2(n1117), .ZN(n1116) );
NOR2_X1 U796 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NAND2_X1 U798 ( .A1(G953), .A2(n1122), .ZN(n1121) );
XOR2_X1 U799 ( .A(n1123), .B(n1124), .Z(n1120) );
XNOR2_X1 U800 ( .A(n1125), .B(n1126), .ZN(n1124) );
XNOR2_X1 U801 ( .A(G116), .B(n1127), .ZN(n1123) );
NAND2_X1 U802 ( .A1(n1128), .A2(KEYINPUT24), .ZN(n1127) );
XOR2_X1 U803 ( .A(n1129), .B(G110), .Z(n1128) );
NAND2_X1 U804 ( .A1(G953), .A2(n1130), .ZN(n1113) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1130) );
NOR2_X1 U806 ( .A1(n1131), .A2(n1132), .ZN(G66) );
XOR2_X1 U807 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U808 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR3_X1 U809 ( .A1(n1131), .A2(n1137), .A3(n1138), .ZN(G63) );
NOR3_X1 U810 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NOR2_X1 U811 ( .A1(KEYINPUT55), .A2(n1142), .ZN(n1141) );
NOR2_X1 U812 ( .A1(n1143), .A2(n1144), .ZN(n1137) );
NOR2_X1 U813 ( .A1(n1142), .A2(n1145), .ZN(n1143) );
INV_X1 U814 ( .A(KEYINPUT55), .ZN(n1145) );
XNOR2_X1 U815 ( .A(n1140), .B(KEYINPUT53), .ZN(n1142) );
AND2_X1 U816 ( .A1(n1135), .A2(G478), .ZN(n1140) );
NOR2_X1 U817 ( .A1(n1131), .A2(n1146), .ZN(G60) );
XOR2_X1 U818 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U819 ( .A1(KEYINPUT42), .A2(n1149), .ZN(n1148) );
NAND3_X1 U820 ( .A1(G475), .A2(n1076), .A3(n1150), .ZN(n1147) );
XOR2_X1 U821 ( .A(n1151), .B(KEYINPUT15), .Z(n1150) );
XNOR2_X1 U822 ( .A(G104), .B(n1152), .ZN(G6) );
NOR2_X1 U823 ( .A1(n1153), .A2(n1154), .ZN(G57) );
XOR2_X1 U824 ( .A(KEYINPUT16), .B(n1131), .Z(n1154) );
XOR2_X1 U825 ( .A(n1155), .B(n1156), .Z(n1153) );
NAND2_X1 U826 ( .A1(n1135), .A2(G472), .ZN(n1155) );
NOR2_X1 U827 ( .A1(n1131), .A2(n1157), .ZN(G54) );
XOR2_X1 U828 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U829 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND3_X1 U830 ( .A1(n1135), .A2(G469), .A3(KEYINPUT18), .ZN(n1160) );
INV_X1 U831 ( .A(n1162), .ZN(n1135) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1158) );
NOR2_X1 U833 ( .A1(KEYINPUT54), .A2(n1110), .ZN(n1164) );
XOR2_X1 U834 ( .A(n1165), .B(n1166), .Z(n1163) );
NOR2_X1 U835 ( .A1(KEYINPUT13), .A2(n1167), .ZN(n1166) );
XOR2_X1 U836 ( .A(n1168), .B(G140), .Z(n1167) );
NOR2_X1 U837 ( .A1(n1131), .A2(n1169), .ZN(G51) );
XOR2_X1 U838 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U839 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U840 ( .A1(KEYINPUT5), .A2(n1174), .ZN(n1173) );
NOR3_X1 U841 ( .A1(n1162), .A2(KEYINPUT43), .A3(n1175), .ZN(n1172) );
NAND2_X1 U842 ( .A1(G902), .A2(n1076), .ZN(n1162) );
NAND3_X1 U843 ( .A1(n1176), .A2(n1177), .A3(n1112), .ZN(n1076) );
AND4_X1 U844 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1112) );
NOR4_X1 U845 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
INV_X1 U846 ( .A(n1186), .ZN(n1184) );
NOR3_X1 U847 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1182) );
NAND3_X1 U848 ( .A1(n1058), .A2(n1190), .A3(n1191), .ZN(n1187) );
XOR2_X1 U849 ( .A(KEYINPUT41), .B(n1192), .Z(n1190) );
AND2_X1 U850 ( .A1(n1193), .A2(n1194), .ZN(n1180) );
NAND3_X1 U851 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1178) );
INV_X1 U852 ( .A(n1198), .ZN(n1197) );
NAND2_X1 U853 ( .A1(KEYINPUT19), .A2(n1199), .ZN(n1196) );
NAND2_X1 U854 ( .A1(n1200), .A2(n1201), .ZN(n1195) );
INV_X1 U855 ( .A(KEYINPUT19), .ZN(n1201) );
OR3_X1 U856 ( .A1(n1047), .A2(n1075), .A3(n1202), .ZN(n1200) );
XOR2_X1 U857 ( .A(KEYINPUT27), .B(n1118), .Z(n1177) );
INV_X1 U858 ( .A(n1119), .ZN(n1176) );
NAND4_X1 U859 ( .A1(n1152), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1119) );
AND3_X1 U860 ( .A1(n1206), .A2(n1207), .A3(n1025), .ZN(n1205) );
NAND3_X1 U861 ( .A1(n1054), .A2(n1208), .A3(n1071), .ZN(n1025) );
NAND2_X1 U862 ( .A1(n1209), .A2(n1210), .ZN(n1204) );
NAND2_X1 U863 ( .A1(n1198), .A2(n1211), .ZN(n1210) );
NAND3_X1 U864 ( .A1(n1212), .A2(n1213), .A3(n1054), .ZN(n1211) );
NAND3_X1 U865 ( .A1(n1054), .A2(n1208), .A3(n1072), .ZN(n1152) );
INV_X1 U866 ( .A(n1028), .ZN(n1131) );
NAND2_X1 U867 ( .A1(G953), .A2(n1030), .ZN(n1028) );
XOR2_X1 U868 ( .A(G146), .B(n1214), .Z(G48) );
NOR2_X1 U869 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U870 ( .A(KEYINPUT59), .B(KEYINPUT25), .Z(n1216) );
INV_X1 U871 ( .A(n1185), .ZN(n1215) );
NOR3_X1 U872 ( .A1(n1189), .A2(n1075), .A3(n1217), .ZN(n1185) );
XOR2_X1 U873 ( .A(n1218), .B(n1219), .Z(G45) );
NAND2_X1 U874 ( .A1(KEYINPUT20), .A2(n1220), .ZN(n1219) );
INV_X1 U875 ( .A(n1179), .ZN(n1220) );
NAND4_X1 U876 ( .A1(n1067), .A2(n1058), .A3(n1048), .A4(n1221), .ZN(n1179) );
NOR3_X1 U877 ( .A1(n1192), .A2(n1222), .A3(n1223), .ZN(n1221) );
INV_X1 U878 ( .A(n1075), .ZN(n1067) );
XOR2_X1 U879 ( .A(n1224), .B(n1194), .Z(G42) );
NAND3_X1 U880 ( .A1(n1050), .A2(n1225), .A3(n1072), .ZN(n1194) );
XOR2_X1 U881 ( .A(n1226), .B(n1193), .Z(G39) );
OR3_X1 U882 ( .A1(n1189), .A2(n1199), .A3(n1043), .ZN(n1193) );
XOR2_X1 U883 ( .A(G134), .B(n1227), .Z(G36) );
NOR2_X1 U884 ( .A1(KEYINPUT1), .A2(n1186), .ZN(n1227) );
NAND3_X1 U885 ( .A1(n1225), .A2(n1071), .A3(n1048), .ZN(n1186) );
XOR2_X1 U886 ( .A(G131), .B(n1228), .Z(G33) );
NOR2_X1 U887 ( .A1(n1199), .A2(n1198), .ZN(n1228) );
INV_X1 U888 ( .A(n1225), .ZN(n1199) );
NOR3_X1 U889 ( .A1(n1075), .A2(n1192), .A3(n1047), .ZN(n1225) );
NAND2_X1 U890 ( .A1(n1229), .A2(n1060), .ZN(n1047) );
INV_X1 U891 ( .A(n1059), .ZN(n1229) );
XNOR2_X1 U892 ( .A(n1080), .B(KEYINPUT28), .ZN(n1059) );
INV_X1 U893 ( .A(n1202), .ZN(n1192) );
XOR2_X1 U894 ( .A(G128), .B(n1230), .Z(G30) );
NOR2_X1 U895 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U896 ( .A(n1233), .B(KEYINPUT39), .Z(n1231) );
NAND4_X1 U897 ( .A1(n1234), .A2(n1071), .A3(n1191), .A4(n1202), .ZN(n1233) );
XOR2_X1 U898 ( .A(n1189), .B(KEYINPUT45), .Z(n1234) );
NAND3_X1 U899 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(G3) );
OR2_X1 U900 ( .A1(n1203), .A2(G101), .ZN(n1237) );
NAND2_X1 U901 ( .A1(KEYINPUT56), .A2(n1238), .ZN(n1236) );
NAND2_X1 U902 ( .A1(G101), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U903 ( .A(KEYINPUT62), .B(n1203), .ZN(n1239) );
NAND2_X1 U904 ( .A1(n1240), .A2(n1241), .ZN(n1235) );
INV_X1 U905 ( .A(KEYINPUT56), .ZN(n1241) );
NAND2_X1 U906 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
NAND3_X1 U907 ( .A1(KEYINPUT62), .A2(G101), .A3(n1203), .ZN(n1243) );
OR2_X1 U908 ( .A1(n1203), .A2(KEYINPUT62), .ZN(n1242) );
NAND3_X1 U909 ( .A1(n1244), .A2(n1208), .A3(n1048), .ZN(n1203) );
XOR2_X1 U910 ( .A(G125), .B(n1183), .Z(G27) );
NOR3_X1 U911 ( .A1(n1217), .A2(n1245), .A3(n1041), .ZN(n1183) );
INV_X1 U912 ( .A(n1246), .ZN(n1041) );
INV_X1 U913 ( .A(n1050), .ZN(n1245) );
NAND3_X1 U914 ( .A1(n1058), .A2(n1202), .A3(n1072), .ZN(n1217) );
NAND2_X1 U915 ( .A1(n1038), .A2(n1247), .ZN(n1202) );
NAND4_X1 U916 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1111), .ZN(n1247) );
INV_X1 U917 ( .A(G900), .ZN(n1111) );
XOR2_X1 U918 ( .A(n1129), .B(n1249), .Z(G24) );
NAND4_X1 U919 ( .A1(n1209), .A2(n1250), .A3(n1212), .A4(n1213), .ZN(n1249) );
XOR2_X1 U920 ( .A(KEYINPUT10), .B(n1054), .Z(n1250) );
NOR2_X1 U921 ( .A1(n1251), .A2(n1081), .ZN(n1054) );
INV_X1 U922 ( .A(n1252), .ZN(n1081) );
XOR2_X1 U923 ( .A(G119), .B(n1118), .Z(G21) );
NOR3_X1 U924 ( .A1(n1043), .A2(n1189), .A3(n1253), .ZN(n1118) );
NAND2_X1 U925 ( .A1(n1254), .A2(n1251), .ZN(n1189) );
XOR2_X1 U926 ( .A(n1252), .B(KEYINPUT6), .Z(n1254) );
XNOR2_X1 U927 ( .A(G116), .B(n1207), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1048), .A2(n1071), .A3(n1209), .ZN(n1207) );
INV_X1 U929 ( .A(n1253), .ZN(n1209) );
INV_X1 U930 ( .A(n1188), .ZN(n1071) );
NAND2_X1 U931 ( .A1(n1223), .A2(n1213), .ZN(n1188) );
XOR2_X1 U932 ( .A(G113), .B(n1255), .Z(G15) );
NOR3_X1 U933 ( .A1(n1253), .A2(KEYINPUT58), .A3(n1198), .ZN(n1255) );
NAND2_X1 U934 ( .A1(n1048), .A2(n1072), .ZN(n1198) );
NOR2_X1 U935 ( .A1(n1213), .A2(n1223), .ZN(n1072) );
INV_X1 U936 ( .A(n1222), .ZN(n1213) );
INV_X1 U937 ( .A(n1053), .ZN(n1048) );
NAND2_X1 U938 ( .A1(n1252), .A2(n1251), .ZN(n1053) );
NAND2_X1 U939 ( .A1(n1246), .A2(n1256), .ZN(n1253) );
NOR2_X1 U940 ( .A1(n1069), .A2(n1090), .ZN(n1246) );
INV_X1 U941 ( .A(n1068), .ZN(n1090) );
XOR2_X1 U942 ( .A(n1168), .B(n1206), .Z(G12) );
NAND3_X1 U943 ( .A1(n1244), .A2(n1208), .A3(n1050), .ZN(n1206) );
NOR2_X1 U944 ( .A1(n1251), .A2(n1252), .ZN(n1050) );
XOR2_X1 U945 ( .A(n1257), .B(n1136), .Z(n1252) );
AND2_X1 U946 ( .A1(G217), .A2(n1258), .ZN(n1136) );
NAND2_X1 U947 ( .A1(n1134), .A2(n1151), .ZN(n1257) );
XOR2_X1 U948 ( .A(n1259), .B(n1260), .Z(n1134) );
XOR2_X1 U949 ( .A(G137), .B(n1261), .Z(n1260) );
XOR2_X1 U950 ( .A(G146), .B(G140), .Z(n1261) );
XOR2_X1 U951 ( .A(n1262), .B(n1263), .Z(n1259) );
XOR2_X1 U952 ( .A(n1264), .B(n1265), .Z(n1262) );
AND2_X1 U953 ( .A1(n1266), .A2(G221), .ZN(n1265) );
NAND3_X1 U954 ( .A1(n1267), .A2(n1268), .A3(KEYINPUT63), .ZN(n1264) );
NAND2_X1 U955 ( .A1(G119), .A2(n1269), .ZN(n1268) );
XOR2_X1 U956 ( .A(KEYINPUT9), .B(n1270), .Z(n1267) );
NOR2_X1 U957 ( .A1(G119), .A2(n1269), .ZN(n1270) );
XNOR2_X1 U958 ( .A(n1089), .B(n1271), .ZN(n1251) );
NOR2_X1 U959 ( .A1(KEYINPUT3), .A2(n1088), .ZN(n1271) );
NAND2_X1 U960 ( .A1(n1156), .A2(n1151), .ZN(n1088) );
XOR2_X1 U961 ( .A(n1272), .B(n1273), .Z(n1156) );
XOR2_X1 U962 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U963 ( .A(G101), .B(KEYINPUT26), .ZN(n1275) );
NAND2_X1 U964 ( .A1(G210), .A2(n1276), .ZN(n1274) );
XOR2_X1 U965 ( .A(n1277), .B(n1278), .Z(n1272) );
INV_X1 U966 ( .A(n1279), .ZN(n1278) );
INV_X1 U967 ( .A(G472), .ZN(n1089) );
AND2_X1 U968 ( .A1(n1256), .A2(n1191), .ZN(n1208) );
XOR2_X1 U969 ( .A(n1075), .B(KEYINPUT22), .Z(n1191) );
NAND2_X1 U970 ( .A1(n1069), .A2(n1068), .ZN(n1075) );
NAND2_X1 U971 ( .A1(G221), .A2(n1258), .ZN(n1068) );
NAND2_X1 U972 ( .A1(n1280), .A2(G234), .ZN(n1258) );
XOR2_X1 U973 ( .A(n1151), .B(KEYINPUT35), .Z(n1280) );
XOR2_X1 U974 ( .A(n1281), .B(G469), .Z(n1069) );
NAND2_X1 U975 ( .A1(KEYINPUT11), .A2(n1084), .ZN(n1281) );
NAND2_X1 U976 ( .A1(n1282), .A2(n1151), .ZN(n1084) );
XOR2_X1 U977 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U978 ( .A(n1165), .B(n1285), .ZN(n1284) );
NOR2_X1 U979 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U980 ( .A(n1288), .B(KEYINPUT44), .Z(n1287) );
NAND2_X1 U981 ( .A1(G140), .A2(n1289), .ZN(n1288) );
XOR2_X1 U982 ( .A(KEYINPUT17), .B(G110), .Z(n1289) );
NOR2_X1 U983 ( .A1(G140), .A2(n1168), .ZN(n1286) );
NAND2_X1 U984 ( .A1(G227), .A2(n1290), .ZN(n1165) );
XNOR2_X1 U985 ( .A(n1161), .B(n1110), .ZN(n1283) );
NAND2_X1 U986 ( .A1(n1291), .A2(n1292), .ZN(n1110) );
NAND2_X1 U987 ( .A1(n1293), .A2(n1269), .ZN(n1292) );
XOR2_X1 U988 ( .A(KEYINPUT7), .B(n1294), .Z(n1291) );
NOR2_X1 U989 ( .A1(n1293), .A2(n1269), .ZN(n1294) );
INV_X1 U990 ( .A(G128), .ZN(n1269) );
XOR2_X1 U991 ( .A(n1218), .B(G146), .Z(n1293) );
XOR2_X1 U992 ( .A(n1295), .B(n1296), .Z(n1161) );
XNOR2_X1 U993 ( .A(G104), .B(n1297), .ZN(n1296) );
NAND2_X1 U994 ( .A1(KEYINPUT36), .A2(G101), .ZN(n1297) );
XOR2_X1 U995 ( .A(n1279), .B(n1298), .Z(n1295) );
NOR2_X1 U996 ( .A1(G107), .A2(KEYINPUT2), .ZN(n1298) );
XOR2_X1 U997 ( .A(n1299), .B(n1300), .Z(n1279) );
XOR2_X1 U998 ( .A(KEYINPUT51), .B(G131), .Z(n1300) );
NAND2_X1 U999 ( .A1(KEYINPUT34), .A2(n1108), .ZN(n1299) );
XOR2_X1 U1000 ( .A(G134), .B(n1226), .Z(n1108) );
INV_X1 U1001 ( .A(G137), .ZN(n1226) );
AND2_X1 U1002 ( .A1(n1058), .A2(n1301), .ZN(n1256) );
NAND2_X1 U1003 ( .A1(n1038), .A2(n1302), .ZN(n1301) );
NAND4_X1 U1004 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1122), .ZN(n1302) );
INV_X1 U1005 ( .A(G898), .ZN(n1122) );
NAND3_X1 U1006 ( .A1(n1248), .A2(n1290), .A3(n1303), .ZN(n1038) );
XOR2_X1 U1007 ( .A(n1030), .B(KEYINPUT49), .Z(n1303) );
INV_X1 U1008 ( .A(G952), .ZN(n1030) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1248) );
INV_X1 U1010 ( .A(n1232), .ZN(n1058) );
NAND2_X1 U1011 ( .A1(n1304), .A2(n1080), .ZN(n1232) );
XOR2_X1 U1012 ( .A(n1305), .B(n1175), .Z(n1080) );
NAND2_X1 U1013 ( .A1(G210), .A2(n1306), .ZN(n1175) );
NAND2_X1 U1014 ( .A1(n1307), .A2(n1151), .ZN(n1305) );
XNOR2_X1 U1015 ( .A(n1170), .B(n1174), .ZN(n1307) );
NAND2_X1 U1016 ( .A1(G224), .A2(n1290), .ZN(n1174) );
XOR2_X1 U1017 ( .A(n1308), .B(n1309), .Z(n1170) );
XOR2_X1 U1018 ( .A(n1129), .B(n1310), .Z(n1309) );
NAND2_X1 U1019 ( .A1(KEYINPUT48), .A2(n1125), .ZN(n1310) );
XOR2_X1 U1020 ( .A(n1311), .B(n1312), .Z(n1125) );
NOR2_X1 U1021 ( .A1(KEYINPUT33), .A2(n1024), .ZN(n1312) );
INV_X1 U1022 ( .A(G107), .ZN(n1024) );
XNOR2_X1 U1023 ( .A(G104), .B(G101), .ZN(n1311) );
XOR2_X1 U1024 ( .A(n1277), .B(n1263), .Z(n1308) );
XOR2_X1 U1025 ( .A(G125), .B(G110), .Z(n1263) );
XOR2_X1 U1026 ( .A(n1313), .B(n1314), .Z(n1277) );
XOR2_X1 U1027 ( .A(n1315), .B(n1126), .Z(n1314) );
XOR2_X1 U1028 ( .A(G113), .B(G119), .Z(n1126) );
NAND2_X1 U1029 ( .A1(n1316), .A2(n1317), .ZN(n1313) );
NAND2_X1 U1030 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
INV_X1 U1031 ( .A(G146), .ZN(n1319) );
XOR2_X1 U1032 ( .A(n1218), .B(KEYINPUT46), .Z(n1318) );
INV_X1 U1033 ( .A(G143), .ZN(n1218) );
NAND2_X1 U1034 ( .A1(n1320), .A2(G146), .ZN(n1316) );
XOR2_X1 U1035 ( .A(KEYINPUT12), .B(G143), .Z(n1320) );
XOR2_X1 U1036 ( .A(n1060), .B(KEYINPUT29), .Z(n1304) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1306), .ZN(n1060) );
NAND2_X1 U1038 ( .A1(n1321), .A2(n1151), .ZN(n1306) );
INV_X1 U1039 ( .A(G237), .ZN(n1321) );
INV_X1 U1040 ( .A(n1043), .ZN(n1244) );
NAND2_X1 U1041 ( .A1(n1222), .A2(n1223), .ZN(n1043) );
INV_X1 U1042 ( .A(n1212), .ZN(n1223) );
NAND2_X1 U1043 ( .A1(n1322), .A2(n1323), .ZN(n1212) );
NAND2_X1 U1044 ( .A1(n1093), .A2(n1095), .ZN(n1323) );
XOR2_X1 U1045 ( .A(n1324), .B(KEYINPUT47), .Z(n1322) );
OR2_X1 U1046 ( .A1(n1095), .A2(n1093), .ZN(n1324) );
NOR2_X1 U1047 ( .A1(n1149), .A2(G902), .ZN(n1093) );
XNOR2_X1 U1048 ( .A(n1325), .B(n1326), .ZN(n1149) );
XNOR2_X1 U1049 ( .A(n1327), .B(n1328), .ZN(n1326) );
NOR2_X1 U1050 ( .A1(G113), .A2(KEYINPUT8), .ZN(n1328) );
NAND3_X1 U1051 ( .A1(n1329), .A2(n1330), .A3(KEYINPUT61), .ZN(n1327) );
NAND3_X1 U1052 ( .A1(KEYINPUT23), .A2(n1331), .A3(n1332), .ZN(n1330) );
NAND2_X1 U1053 ( .A1(n1333), .A2(n1334), .ZN(n1329) );
NAND2_X1 U1054 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
OR2_X1 U1055 ( .A1(n1331), .A2(KEYINPUT37), .ZN(n1336) );
NAND2_X1 U1056 ( .A1(n1331), .A2(n1337), .ZN(n1335) );
NAND2_X1 U1057 ( .A1(KEYINPUT23), .A2(n1338), .ZN(n1337) );
INV_X1 U1058 ( .A(KEYINPUT37), .ZN(n1338) );
XOR2_X1 U1059 ( .A(n1339), .B(n1340), .Z(n1331) );
XOR2_X1 U1060 ( .A(KEYINPUT38), .B(G143), .Z(n1340) );
XOR2_X1 U1061 ( .A(n1341), .B(G131), .Z(n1339) );
NAND2_X1 U1062 ( .A1(G214), .A2(n1276), .ZN(n1341) );
NOR2_X1 U1063 ( .A1(G953), .A2(G237), .ZN(n1276) );
INV_X1 U1064 ( .A(n1332), .ZN(n1333) );
XOR2_X1 U1065 ( .A(n1342), .B(n1343), .Z(n1332) );
XOR2_X1 U1066 ( .A(G146), .B(G125), .Z(n1343) );
NAND2_X1 U1067 ( .A1(KEYINPUT14), .A2(n1224), .ZN(n1342) );
INV_X1 U1068 ( .A(G140), .ZN(n1224) );
XOR2_X1 U1069 ( .A(G104), .B(n1129), .Z(n1325) );
INV_X1 U1070 ( .A(G122), .ZN(n1129) );
INV_X1 U1071 ( .A(G475), .ZN(n1095) );
NOR2_X1 U1072 ( .A1(n1344), .A2(n1092), .ZN(n1222) );
NOR3_X1 U1073 ( .A1(G478), .A2(G902), .A3(n1144), .ZN(n1092) );
XOR2_X1 U1074 ( .A(n1091), .B(KEYINPUT57), .Z(n1344) );
AND2_X1 U1075 ( .A1(G478), .A2(n1345), .ZN(n1091) );
NAND2_X1 U1076 ( .A1(n1139), .A2(n1151), .ZN(n1345) );
INV_X1 U1077 ( .A(G902), .ZN(n1151) );
INV_X1 U1078 ( .A(n1144), .ZN(n1139) );
XOR2_X1 U1079 ( .A(n1346), .B(n1347), .Z(n1144) );
XOR2_X1 U1080 ( .A(G122), .B(n1348), .Z(n1347) );
XOR2_X1 U1081 ( .A(G143), .B(G134), .Z(n1348) );
XOR2_X1 U1082 ( .A(n1349), .B(n1315), .Z(n1346) );
XOR2_X1 U1083 ( .A(G116), .B(G128), .Z(n1315) );
XOR2_X1 U1084 ( .A(n1350), .B(G107), .Z(n1349) );
NAND2_X1 U1085 ( .A1(G217), .A2(n1266), .ZN(n1350) );
AND2_X1 U1086 ( .A1(G234), .A2(n1290), .ZN(n1266) );
INV_X1 U1087 ( .A(G953), .ZN(n1290) );
INV_X1 U1088 ( .A(G110), .ZN(n1168) );
endmodule


