//Key = 0110001011101111100100010011100101011100000011111001100101011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280;

XOR2_X1 U710 ( .A(G107), .B(n976), .Z(G9) );
NOR2_X1 U711 ( .A1(KEYINPUT18), .A2(n977), .ZN(n976) );
NOR2_X1 U712 ( .A1(n978), .A2(n979), .ZN(G75) );
NOR4_X1 U713 ( .A1(n980), .A2(n981), .A3(n982), .A4(n983), .ZN(n979) );
XOR2_X1 U714 ( .A(n984), .B(KEYINPUT50), .Z(n982) );
NAND2_X1 U715 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND3_X1 U716 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
NAND2_X1 U717 ( .A1(n990), .A2(n991), .ZN(n988) );
NAND3_X1 U718 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND2_X1 U719 ( .A1(n995), .A2(n996), .ZN(n990) );
NAND2_X1 U720 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U721 ( .A1(n994), .A2(n999), .ZN(n998) );
NAND2_X1 U722 ( .A1(n992), .A2(n1000), .ZN(n997) );
NAND2_X1 U723 ( .A1(n1001), .A2(n994), .ZN(n985) );
XOR2_X1 U724 ( .A(n1002), .B(KEYINPUT55), .Z(n1001) );
NAND4_X1 U725 ( .A1(n989), .A2(n995), .A3(n1003), .A4(n992), .ZN(n1002) );
NAND3_X1 U726 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n980) );
NAND2_X1 U727 ( .A1(n989), .A2(n1007), .ZN(n1006) );
NAND2_X1 U728 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
NAND3_X1 U729 ( .A1(n995), .A2(n1010), .A3(n994), .ZN(n1009) );
NAND2_X1 U730 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND3_X1 U731 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
XNOR2_X1 U732 ( .A(KEYINPUT41), .B(n1016), .ZN(n1013) );
NAND2_X1 U733 ( .A1(n1017), .A2(n992), .ZN(n1011) );
NAND3_X1 U734 ( .A1(n992), .A2(n1018), .A3(n987), .ZN(n1008) );
NAND2_X1 U735 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND3_X1 U736 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
XOR2_X1 U737 ( .A(KEYINPUT21), .B(n994), .Z(n1022) );
NAND3_X1 U738 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1019) );
XOR2_X1 U739 ( .A(KEYINPUT32), .B(n995), .Z(n1025) );
NOR2_X1 U740 ( .A1(KEYINPUT61), .A2(n1027), .ZN(n989) );
NOR3_X1 U741 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n978) );
INV_X1 U742 ( .A(n1004), .ZN(n1028) );
NAND4_X1 U743 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1004) );
NOR4_X1 U744 ( .A1(n1033), .A2(n1016), .A3(n1034), .A4(n1035), .ZN(n1032) );
XOR2_X1 U745 ( .A(KEYINPUT25), .B(n1036), .Z(n1035) );
XOR2_X1 U746 ( .A(KEYINPUT38), .B(n1037), .Z(n1034) );
NOR2_X1 U747 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XNOR2_X1 U748 ( .A(KEYINPUT36), .B(n1040), .ZN(n1039) );
INV_X1 U749 ( .A(n987), .ZN(n1016) );
XNOR2_X1 U750 ( .A(G469), .B(n1041), .ZN(n1033) );
NOR2_X1 U751 ( .A1(n1042), .A2(KEYINPUT53), .ZN(n1041) );
INV_X1 U752 ( .A(n1043), .ZN(n1042) );
NOR3_X1 U753 ( .A1(n1044), .A2(n1026), .A3(n1023), .ZN(n1031) );
NAND2_X1 U754 ( .A1(n1038), .A2(n1040), .ZN(n1030) );
XOR2_X1 U755 ( .A(n1045), .B(n1046), .Z(n1029) );
NAND2_X1 U756 ( .A1(KEYINPUT27), .A2(n1047), .ZN(n1046) );
XOR2_X1 U757 ( .A(n1048), .B(n1049), .Z(G72) );
XOR2_X1 U758 ( .A(n1050), .B(n1051), .Z(n1049) );
NAND2_X1 U759 ( .A1(G953), .A2(n1052), .ZN(n1051) );
NAND2_X1 U760 ( .A1(G900), .A2(G227), .ZN(n1052) );
NAND2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
NAND2_X1 U762 ( .A1(G953), .A2(n1055), .ZN(n1054) );
XNOR2_X1 U763 ( .A(n1056), .B(n1057), .ZN(n1053) );
NAND2_X1 U764 ( .A1(KEYINPUT45), .A2(n1058), .ZN(n1056) );
XNOR2_X1 U765 ( .A(n1059), .B(n1060), .ZN(n1058) );
XNOR2_X1 U766 ( .A(n1061), .B(n1062), .ZN(n1060) );
NAND2_X1 U767 ( .A1(KEYINPUT1), .A2(n1063), .ZN(n1061) );
XOR2_X1 U768 ( .A(n1064), .B(G131), .Z(n1063) );
NAND2_X1 U769 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
INV_X1 U771 ( .A(KEYINPUT0), .ZN(n1068) );
NAND3_X1 U772 ( .A1(n1069), .A2(n1070), .A3(KEYINPUT0), .ZN(n1065) );
AND2_X1 U773 ( .A1(n981), .A2(n1005), .ZN(n1048) );
NAND2_X1 U774 ( .A1(n1071), .A2(n1072), .ZN(G69) );
NAND2_X1 U775 ( .A1(n1073), .A2(n1005), .ZN(n1072) );
XNOR2_X1 U776 ( .A(n1074), .B(n983), .ZN(n1073) );
NAND2_X1 U777 ( .A1(n1075), .A2(G953), .ZN(n1071) );
NAND2_X1 U778 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U779 ( .A1(n1074), .A2(n1078), .ZN(n1077) );
INV_X1 U780 ( .A(G224), .ZN(n1078) );
NAND2_X1 U781 ( .A1(G224), .A2(n1079), .ZN(n1076) );
NAND2_X1 U782 ( .A1(G898), .A2(n1074), .ZN(n1079) );
NAND3_X1 U783 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1074) );
NAND2_X1 U784 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NOR2_X1 U785 ( .A1(n1084), .A2(n1085), .ZN(G66) );
XOR2_X1 U786 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U787 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U788 ( .A1(n1084), .A2(n1090), .ZN(G63) );
XNOR2_X1 U789 ( .A(n1091), .B(n1092), .ZN(n1090) );
XNOR2_X1 U790 ( .A(KEYINPUT13), .B(n1093), .ZN(n1092) );
NOR3_X1 U791 ( .A1(n1089), .A2(KEYINPUT7), .A3(n1094), .ZN(n1093) );
NOR2_X1 U792 ( .A1(n1084), .A2(n1095), .ZN(G60) );
XOR2_X1 U793 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U794 ( .A1(n1098), .A2(n1089), .ZN(n1096) );
XNOR2_X1 U795 ( .A(G104), .B(n1099), .ZN(G6) );
NOR2_X1 U796 ( .A1(n1084), .A2(n1100), .ZN(G57) );
XOR2_X1 U797 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U798 ( .A1(KEYINPUT3), .A2(n1103), .ZN(n1102) );
XOR2_X1 U799 ( .A(n1104), .B(n1105), .Z(n1101) );
NOR2_X1 U800 ( .A1(n1040), .A2(n1089), .ZN(n1105) );
NAND2_X1 U801 ( .A1(KEYINPUT37), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U802 ( .A(G101), .B(n1107), .ZN(n1106) );
NAND2_X1 U803 ( .A1(KEYINPUT23), .A2(n1108), .ZN(n1107) );
NOR2_X1 U804 ( .A1(n1084), .A2(n1109), .ZN(G54) );
XNOR2_X1 U805 ( .A(n1110), .B(n1111), .ZN(n1109) );
XOR2_X1 U806 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U807 ( .A1(n1114), .A2(n1089), .ZN(n1113) );
INV_X1 U808 ( .A(G469), .ZN(n1114) );
NOR2_X1 U809 ( .A1(n1084), .A2(n1115), .ZN(G51) );
XOR2_X1 U810 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U811 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U812 ( .A1(n1045), .A2(n1089), .ZN(n1119) );
NAND2_X1 U813 ( .A1(G902), .A2(n1120), .ZN(n1089) );
OR2_X1 U814 ( .A1(n981), .A2(n983), .ZN(n1120) );
NAND4_X1 U815 ( .A1(n1121), .A2(n1099), .A3(n1122), .A4(n1123), .ZN(n983) );
AND4_X1 U816 ( .A1(n977), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1123) );
NAND3_X1 U817 ( .A1(n992), .A2(n1127), .A3(n1017), .ZN(n977) );
NOR2_X1 U818 ( .A1(n1128), .A2(n1129), .ZN(n1122) );
NOR2_X1 U819 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U820 ( .A(KEYINPUT62), .B(n1132), .Z(n1131) );
NOR3_X1 U821 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1128) );
NAND3_X1 U822 ( .A1(n992), .A2(n1127), .A3(n1003), .ZN(n1099) );
NAND4_X1 U823 ( .A1(n1136), .A2(n992), .A3(n1137), .A4(n1138), .ZN(n1121) );
OR2_X1 U824 ( .A1(n1139), .A2(KEYINPUT5), .ZN(n1138) );
NAND2_X1 U825 ( .A1(KEYINPUT5), .A2(n1140), .ZN(n1137) );
NAND3_X1 U826 ( .A1(n1141), .A2(n1130), .A3(n995), .ZN(n1140) );
NAND2_X1 U827 ( .A1(n1142), .A2(n1143), .ZN(n981) );
NOR4_X1 U828 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
NOR4_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1142) );
NOR3_X1 U830 ( .A1(n1152), .A2(n1130), .A3(n1153), .ZN(n1151) );
INV_X1 U831 ( .A(n1154), .ZN(n1150) );
NAND2_X1 U832 ( .A1(KEYINPUT59), .A2(n1155), .ZN(n1116) );
NOR2_X1 U833 ( .A1(n1005), .A2(G952), .ZN(n1084) );
XOR2_X1 U834 ( .A(n1156), .B(n1149), .Z(G48) );
AND3_X1 U835 ( .A1(n1003), .A2(n1000), .A3(n1157), .ZN(n1149) );
XNOR2_X1 U836 ( .A(G146), .B(KEYINPUT10), .ZN(n1156) );
XNOR2_X1 U837 ( .A(G143), .B(n1158), .ZN(G45) );
NAND3_X1 U838 ( .A1(n1159), .A2(n1160), .A3(n1136), .ZN(n1158) );
XNOR2_X1 U839 ( .A(KEYINPUT42), .B(n1130), .ZN(n1160) );
INV_X1 U840 ( .A(n1000), .ZN(n1130) );
XOR2_X1 U841 ( .A(n1161), .B(G140), .Z(G42) );
NAND2_X1 U842 ( .A1(KEYINPUT14), .A2(n1154), .ZN(n1161) );
NAND3_X1 U843 ( .A1(n1162), .A2(n993), .A3(n994), .ZN(n1154) );
XOR2_X1 U844 ( .A(n1148), .B(n1163), .Z(G39) );
XNOR2_X1 U845 ( .A(KEYINPUT43), .B(n1070), .ZN(n1163) );
AND3_X1 U846 ( .A1(n1157), .A2(n987), .A3(n994), .ZN(n1148) );
XOR2_X1 U847 ( .A(G134), .B(n1147), .Z(G36) );
AND3_X1 U848 ( .A1(n1159), .A2(n1017), .A3(n994), .ZN(n1147) );
XNOR2_X1 U849 ( .A(G131), .B(n1164), .ZN(G33) );
NAND2_X1 U850 ( .A1(KEYINPUT6), .A2(n1146), .ZN(n1164) );
AND3_X1 U851 ( .A1(n1159), .A2(n1003), .A3(n994), .ZN(n1146) );
NOR2_X1 U852 ( .A1(n1165), .A2(n1026), .ZN(n994) );
INV_X1 U853 ( .A(n1153), .ZN(n1159) );
NAND3_X1 U854 ( .A1(n993), .A2(n1166), .A3(n999), .ZN(n1153) );
XNOR2_X1 U855 ( .A(G128), .B(n1167), .ZN(G30) );
NAND2_X1 U856 ( .A1(KEYINPUT57), .A2(n1145), .ZN(n1167) );
AND3_X1 U857 ( .A1(n1017), .A2(n1000), .A3(n1157), .ZN(n1145) );
AND4_X1 U858 ( .A1(n993), .A2(n1014), .A3(n1168), .A4(n1166), .ZN(n1157) );
XNOR2_X1 U859 ( .A(G101), .B(n1169), .ZN(G3) );
NAND3_X1 U860 ( .A1(n1132), .A2(n1000), .A3(KEYINPUT2), .ZN(n1169) );
AND4_X1 U861 ( .A1(n999), .A2(n987), .A3(n993), .A4(n1141), .ZN(n1132) );
NAND2_X1 U862 ( .A1(n1170), .A2(n1171), .ZN(G27) );
OR2_X1 U863 ( .A1(n1172), .A2(G125), .ZN(n1171) );
NAND2_X1 U864 ( .A1(G125), .A2(n1173), .ZN(n1170) );
NAND2_X1 U865 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND2_X1 U866 ( .A1(n1144), .A2(n1176), .ZN(n1175) );
INV_X1 U867 ( .A(KEYINPUT52), .ZN(n1176) );
NAND2_X1 U868 ( .A1(KEYINPUT52), .A2(n1172), .ZN(n1174) );
NAND2_X1 U869 ( .A1(KEYINPUT12), .A2(n1144), .ZN(n1172) );
AND3_X1 U870 ( .A1(n1162), .A2(n1000), .A3(n995), .ZN(n1144) );
AND4_X1 U871 ( .A1(n1015), .A2(n1003), .A3(n1014), .A4(n1166), .ZN(n1162) );
NAND2_X1 U872 ( .A1(n1177), .A2(n1178), .ZN(n1166) );
NAND2_X1 U873 ( .A1(n1179), .A2(n1055), .ZN(n1178) );
INV_X1 U874 ( .A(G900), .ZN(n1055) );
XOR2_X1 U875 ( .A(G122), .B(n1180), .Z(G24) );
AND3_X1 U876 ( .A1(n1139), .A2(n992), .A3(n1136), .ZN(n1180) );
INV_X1 U877 ( .A(n1152), .ZN(n1136) );
NAND2_X1 U878 ( .A1(n1181), .A2(n1182), .ZN(n1152) );
NOR2_X1 U879 ( .A1(n1183), .A2(n1168), .ZN(n992) );
XNOR2_X1 U880 ( .A(G119), .B(n1126), .ZN(G21) );
NAND4_X1 U881 ( .A1(n1139), .A2(n987), .A3(n1014), .A4(n1168), .ZN(n1126) );
INV_X1 U882 ( .A(n1015), .ZN(n1168) );
XOR2_X1 U883 ( .A(G116), .B(n1184), .Z(G18) );
NOR4_X1 U884 ( .A1(KEYINPUT30), .A2(n1134), .A3(n1135), .A4(n1133), .ZN(n1184) );
INV_X1 U885 ( .A(n999), .ZN(n1135) );
INV_X1 U886 ( .A(n1017), .ZN(n1134) );
NOR2_X1 U887 ( .A1(n1182), .A2(n1185), .ZN(n1017) );
XNOR2_X1 U888 ( .A(G113), .B(n1125), .ZN(G15) );
NAND3_X1 U889 ( .A1(n999), .A2(n1003), .A3(n1139), .ZN(n1125) );
INV_X1 U890 ( .A(n1133), .ZN(n1139) );
NAND3_X1 U891 ( .A1(n1000), .A2(n1141), .A3(n995), .ZN(n1133) );
NOR2_X1 U892 ( .A1(n1186), .A2(n1023), .ZN(n995) );
AND2_X1 U893 ( .A1(n1185), .A2(n1182), .ZN(n1003) );
INV_X1 U894 ( .A(n1181), .ZN(n1185) );
NOR2_X1 U895 ( .A1(n1183), .A2(n1015), .ZN(n999) );
XNOR2_X1 U896 ( .A(G110), .B(n1124), .ZN(G12) );
NAND4_X1 U897 ( .A1(n987), .A2(n1127), .A3(n1015), .A4(n1014), .ZN(n1124) );
XNOR2_X1 U898 ( .A(n1183), .B(KEYINPUT19), .ZN(n1014) );
OR2_X1 U899 ( .A1(n1036), .A2(n1044), .ZN(n1183) );
NOR2_X1 U900 ( .A1(n1187), .A2(n1088), .ZN(n1044) );
AND2_X1 U901 ( .A1(n1187), .A2(n1088), .ZN(n1036) );
NAND2_X1 U902 ( .A1(G217), .A2(n1188), .ZN(n1088) );
NOR2_X1 U903 ( .A1(n1087), .A2(G902), .ZN(n1187) );
XNOR2_X1 U904 ( .A(n1189), .B(n1190), .ZN(n1087) );
XOR2_X1 U905 ( .A(G128), .B(G125), .Z(n1190) );
XOR2_X1 U906 ( .A(n1191), .B(G119), .Z(n1189) );
XOR2_X1 U907 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U908 ( .A(n1194), .B(n1195), .Z(n1193) );
XNOR2_X1 U909 ( .A(n1070), .B(n1196), .ZN(n1195) );
NOR2_X1 U910 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
INV_X1 U911 ( .A(G221), .ZN(n1198) );
INV_X1 U912 ( .A(G137), .ZN(n1070) );
XOR2_X1 U913 ( .A(n1199), .B(KEYINPUT29), .Z(n1192) );
XNOR2_X1 U914 ( .A(KEYINPUT39), .B(KEYINPUT9), .ZN(n1199) );
XOR2_X1 U915 ( .A(n1038), .B(n1040), .Z(n1015) );
INV_X1 U916 ( .A(G472), .ZN(n1040) );
AND3_X1 U917 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1038) );
NAND2_X1 U918 ( .A1(n1203), .A2(n1204), .ZN(n1201) );
INV_X1 U919 ( .A(G101), .ZN(n1204) );
XOR2_X1 U920 ( .A(n1205), .B(n1103), .Z(n1203) );
NAND2_X1 U921 ( .A1(KEYINPUT47), .A2(n1206), .ZN(n1205) );
XOR2_X1 U922 ( .A(KEYINPUT31), .B(n1108), .Z(n1206) );
NAND2_X1 U923 ( .A1(n1207), .A2(G101), .ZN(n1200) );
XOR2_X1 U924 ( .A(n1208), .B(n1103), .Z(n1207) );
XOR2_X1 U925 ( .A(n1209), .B(n1210), .Z(n1103) );
XOR2_X1 U926 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U927 ( .A(n1213), .B(n1214), .Z(n1209) );
XNOR2_X1 U928 ( .A(KEYINPUT58), .B(KEYINPUT54), .ZN(n1213) );
NAND2_X1 U929 ( .A1(KEYINPUT47), .A2(n1108), .ZN(n1208) );
AND3_X1 U930 ( .A1(n1215), .A2(n1216), .A3(G210), .ZN(n1108) );
XNOR2_X1 U931 ( .A(KEYINPUT15), .B(n1217), .ZN(n1215) );
AND3_X1 U932 ( .A1(n993), .A2(n1141), .A3(n1000), .ZN(n1127) );
NOR2_X1 U933 ( .A1(n1024), .A2(n1026), .ZN(n1000) );
AND2_X1 U934 ( .A1(G214), .A2(n1218), .ZN(n1026) );
INV_X1 U935 ( .A(n1165), .ZN(n1024) );
XOR2_X1 U936 ( .A(n1047), .B(n1045), .Z(n1165) );
NAND2_X1 U937 ( .A1(G210), .A2(n1218), .ZN(n1045) );
NAND2_X1 U938 ( .A1(n1202), .A2(n1217), .ZN(n1218) );
NAND2_X1 U939 ( .A1(n1219), .A2(n1202), .ZN(n1047) );
XOR2_X1 U940 ( .A(n1155), .B(n1118), .Z(n1219) );
AND2_X1 U941 ( .A1(n1220), .A2(n1081), .ZN(n1118) );
NAND2_X1 U942 ( .A1(n1221), .A2(n1222), .ZN(n1081) );
XNOR2_X1 U943 ( .A(KEYINPUT51), .B(n1080), .ZN(n1220) );
OR2_X1 U944 ( .A1(n1222), .A2(n1221), .ZN(n1080) );
XNOR2_X1 U945 ( .A(G110), .B(G122), .ZN(n1221) );
XNOR2_X1 U946 ( .A(n1223), .B(n1224), .ZN(n1222) );
XNOR2_X1 U947 ( .A(n1225), .B(n1226), .ZN(n1224) );
XOR2_X1 U948 ( .A(KEYINPUT22), .B(G107), .Z(n1226) );
XOR2_X1 U949 ( .A(n1212), .B(n1227), .Z(n1223) );
XOR2_X1 U950 ( .A(G113), .B(n1228), .Z(n1212) );
XOR2_X1 U951 ( .A(G119), .B(G116), .Z(n1228) );
XOR2_X1 U952 ( .A(n1229), .B(n1230), .Z(n1155) );
XOR2_X1 U953 ( .A(G125), .B(n1214), .Z(n1230) );
NOR2_X1 U954 ( .A1(KEYINPUT17), .A2(n1062), .ZN(n1214) );
XNOR2_X1 U955 ( .A(n1231), .B(n1232), .ZN(n1229) );
NAND2_X1 U956 ( .A1(G224), .A2(n1216), .ZN(n1231) );
NAND2_X1 U957 ( .A1(n1177), .A2(n1233), .ZN(n1141) );
NAND2_X1 U958 ( .A1(n1179), .A2(n1083), .ZN(n1233) );
INV_X1 U959 ( .A(G898), .ZN(n1083) );
NOR3_X1 U960 ( .A1(n1005), .A2(n1027), .A3(n1202), .ZN(n1179) );
INV_X1 U961 ( .A(n1234), .ZN(n1027) );
NAND3_X1 U962 ( .A1(n1234), .A2(n1005), .A3(G952), .ZN(n1177) );
NAND2_X1 U963 ( .A1(G237), .A2(G234), .ZN(n1234) );
NOR2_X1 U964 ( .A1(n1021), .A2(n1023), .ZN(n993) );
AND2_X1 U965 ( .A1(G221), .A2(n1188), .ZN(n1023) );
NAND2_X1 U966 ( .A1(G234), .A2(n1202), .ZN(n1188) );
INV_X1 U967 ( .A(n1186), .ZN(n1021) );
NAND2_X1 U968 ( .A1(n1235), .A2(n1236), .ZN(n1186) );
NAND2_X1 U969 ( .A1(G469), .A2(n1043), .ZN(n1236) );
XOR2_X1 U970 ( .A(KEYINPUT8), .B(n1237), .Z(n1235) );
NOR2_X1 U971 ( .A1(G469), .A2(n1043), .ZN(n1237) );
NAND2_X1 U972 ( .A1(n1238), .A2(n1202), .ZN(n1043) );
XOR2_X1 U973 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U974 ( .A(KEYINPUT33), .B(KEYINPUT11), .Z(n1240) );
XNOR2_X1 U975 ( .A(n1241), .B(n1242), .ZN(n1239) );
INV_X1 U976 ( .A(n1110), .ZN(n1242) );
XNOR2_X1 U977 ( .A(n1243), .B(n1244), .ZN(n1110) );
XOR2_X1 U978 ( .A(n1194), .B(n1211), .Z(n1244) );
XNOR2_X1 U979 ( .A(n1232), .B(n1245), .ZN(n1211) );
XOR2_X1 U980 ( .A(G131), .B(n1246), .Z(n1245) );
NOR2_X1 U981 ( .A1(KEYINPUT34), .A2(n1067), .ZN(n1246) );
XNOR2_X1 U982 ( .A(G137), .B(n1069), .ZN(n1067) );
INV_X1 U983 ( .A(n1059), .ZN(n1232) );
XOR2_X1 U984 ( .A(n1247), .B(KEYINPUT24), .Z(n1059) );
XOR2_X1 U985 ( .A(G110), .B(n1248), .Z(n1194) );
XNOR2_X1 U986 ( .A(n1062), .B(G140), .ZN(n1248) );
XOR2_X1 U987 ( .A(n1249), .B(KEYINPUT48), .Z(n1243) );
NAND2_X1 U988 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND3_X1 U989 ( .A1(n1227), .A2(n1252), .A3(n1253), .ZN(n1251) );
NAND2_X1 U990 ( .A1(n1254), .A2(n1255), .ZN(n1250) );
NAND2_X1 U991 ( .A1(n1253), .A2(n1252), .ZN(n1255) );
NAND2_X1 U992 ( .A1(n1256), .A2(n1257), .ZN(n1252) );
XOR2_X1 U993 ( .A(KEYINPUT46), .B(G107), .Z(n1257) );
XNOR2_X1 U994 ( .A(G104), .B(KEYINPUT26), .ZN(n1256) );
XOR2_X1 U995 ( .A(n1258), .B(KEYINPUT4), .Z(n1253) );
NAND2_X1 U996 ( .A1(n1259), .A2(n1225), .ZN(n1258) );
XNOR2_X1 U997 ( .A(KEYINPUT46), .B(G107), .ZN(n1259) );
XOR2_X1 U998 ( .A(n1227), .B(KEYINPUT44), .Z(n1254) );
XNOR2_X1 U999 ( .A(G101), .B(KEYINPUT63), .ZN(n1227) );
NAND2_X1 U1000 ( .A1(KEYINPUT35), .A2(n1112), .ZN(n1241) );
NAND2_X1 U1001 ( .A1(G227), .A2(n1216), .ZN(n1112) );
NOR2_X1 U1002 ( .A1(n1181), .A2(n1182), .ZN(n987) );
XOR2_X1 U1003 ( .A(n1260), .B(n1098), .Z(n1182) );
INV_X1 U1004 ( .A(G475), .ZN(n1098) );
OR2_X1 U1005 ( .A1(n1097), .A2(G902), .ZN(n1260) );
XNOR2_X1 U1006 ( .A(n1261), .B(n1262), .ZN(n1097) );
XNOR2_X1 U1007 ( .A(n1225), .B(n1263), .ZN(n1262) );
NOR2_X1 U1008 ( .A1(KEYINPUT49), .A2(n1264), .ZN(n1263) );
XOR2_X1 U1009 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U1010 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U1011 ( .A(G143), .B(G131), .Z(n1268) );
NOR2_X1 U1012 ( .A1(KEYINPUT20), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U1013 ( .A(KEYINPUT39), .B(n1062), .ZN(n1269) );
INV_X1 U1014 ( .A(G146), .ZN(n1062) );
XOR2_X1 U1015 ( .A(n1270), .B(n1057), .Z(n1265) );
XOR2_X1 U1016 ( .A(G140), .B(G125), .Z(n1057) );
NAND3_X1 U1017 ( .A1(n1216), .A2(n1217), .A3(G214), .ZN(n1270) );
INV_X1 U1018 ( .A(G237), .ZN(n1217) );
INV_X1 U1019 ( .A(G104), .ZN(n1225) );
XNOR2_X1 U1020 ( .A(G113), .B(G122), .ZN(n1261) );
XOR2_X1 U1021 ( .A(n1271), .B(n1094), .Z(n1181) );
INV_X1 U1022 ( .A(G478), .ZN(n1094) );
NAND2_X1 U1023 ( .A1(n1091), .A2(n1202), .ZN(n1271) );
INV_X1 U1024 ( .A(G902), .ZN(n1202) );
XNOR2_X1 U1025 ( .A(n1272), .B(n1273), .ZN(n1091) );
XOR2_X1 U1026 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U1027 ( .A(G122), .B(G107), .Z(n1275) );
NOR2_X1 U1028 ( .A1(n1197), .A2(n1276), .ZN(n1274) );
INV_X1 U1029 ( .A(G217), .ZN(n1276) );
NAND2_X1 U1030 ( .A1(n1277), .A2(n1216), .ZN(n1197) );
XNOR2_X1 U1031 ( .A(n1005), .B(KEYINPUT28), .ZN(n1216) );
INV_X1 U1032 ( .A(G953), .ZN(n1005) );
XOR2_X1 U1033 ( .A(KEYINPUT56), .B(G234), .Z(n1277) );
XOR2_X1 U1034 ( .A(n1278), .B(n1069), .Z(n1272) );
XOR2_X1 U1035 ( .A(G134), .B(KEYINPUT40), .Z(n1069) );
XNOR2_X1 U1036 ( .A(n1279), .B(n1280), .ZN(n1278) );
NAND2_X1 U1037 ( .A1(KEYINPUT60), .A2(G116), .ZN(n1280) );
NAND2_X1 U1038 ( .A1(KEYINPUT16), .A2(n1247), .ZN(n1279) );
XOR2_X1 U1039 ( .A(G128), .B(G143), .Z(n1247) );
endmodule


