//Key = 0011001011101000100111100011101001100010111001010110001011010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368;

XNOR2_X1 U752 ( .A(G107), .B(n1052), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(G75) );
NOR4_X1 U754 ( .A1(G953), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1054) );
NOR2_X1 U755 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR3_X1 U757 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NOR2_X1 U758 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U761 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U762 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1069) );
NOR2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR2_X1 U766 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR3_X1 U767 ( .A1(n1078), .A2(n1083), .A3(n1072), .ZN(n1065) );
NOR2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U769 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR4_X1 U770 ( .A1(n1088), .A2(n1072), .A3(n1068), .A4(n1078), .ZN(n1060) );
NOR2_X1 U771 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR3_X1 U772 ( .A1(n1055), .A2(G953), .A3(G952), .ZN(n1053) );
AND4_X1 U773 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1055) );
NOR3_X1 U774 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
XNOR2_X1 U775 ( .A(n1081), .B(KEYINPUT1), .ZN(n1097) );
NOR2_X1 U776 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NAND3_X1 U777 ( .A1(n1100), .A2(n1101), .A3(n1076), .ZN(n1095) );
NOR3_X1 U778 ( .A1(n1068), .A2(n1102), .A3(n1103), .ZN(n1093) );
AND2_X1 U779 ( .A1(n1104), .A2(KEYINPUT51), .ZN(n1103) );
NOR3_X1 U780 ( .A1(KEYINPUT51), .A2(n1104), .A3(n1105), .ZN(n1102) );
XNOR2_X1 U781 ( .A(G472), .B(n1106), .ZN(n1092) );
NAND2_X1 U782 ( .A1(KEYINPUT10), .A2(n1107), .ZN(n1106) );
XOR2_X1 U783 ( .A(n1108), .B(n1109), .Z(n1091) );
NOR2_X1 U784 ( .A1(G475), .A2(KEYINPUT55), .ZN(n1109) );
XOR2_X1 U785 ( .A(n1110), .B(n1111), .Z(G72) );
NOR2_X1 U786 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
AND2_X1 U787 ( .A1(G227), .A2(G900), .ZN(n1112) );
NAND2_X1 U788 ( .A1(n1114), .A2(n1115), .ZN(n1110) );
NAND3_X1 U789 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
NAND2_X1 U790 ( .A1(G953), .A2(n1119), .ZN(n1117) );
NAND2_X1 U791 ( .A1(n1120), .A2(n1113), .ZN(n1116) );
XOR2_X1 U792 ( .A(KEYINPUT63), .B(n1121), .Z(n1114) );
NOR3_X1 U793 ( .A1(n1118), .A2(G953), .A3(n1122), .ZN(n1121) );
INV_X1 U794 ( .A(n1120), .ZN(n1122) );
XNOR2_X1 U795 ( .A(n1123), .B(n1124), .ZN(n1118) );
XNOR2_X1 U796 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR2_X1 U797 ( .A1(KEYINPUT39), .A2(n1127), .ZN(n1126) );
XOR2_X1 U798 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U799 ( .A(G131), .B(n1130), .Z(n1129) );
NOR2_X1 U800 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U801 ( .A(n1133), .B(KEYINPUT57), .Z(n1132) );
NAND2_X1 U802 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U803 ( .A1(n1136), .A2(n1134), .ZN(n1131) );
XNOR2_X1 U804 ( .A(G137), .B(KEYINPUT37), .ZN(n1136) );
NAND2_X1 U805 ( .A1(KEYINPUT41), .A2(n1137), .ZN(n1125) );
XNOR2_X1 U806 ( .A(n1138), .B(n1139), .ZN(n1123) );
INV_X1 U807 ( .A(G140), .ZN(n1139) );
XNOR2_X1 U808 ( .A(KEYINPUT28), .B(KEYINPUT18), .ZN(n1138) );
NAND2_X1 U809 ( .A1(n1140), .A2(n1141), .ZN(G69) );
NAND2_X1 U810 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
OR2_X1 U811 ( .A1(n1113), .A2(G224), .ZN(n1143) );
NAND3_X1 U812 ( .A1(G953), .A2(n1144), .A3(n1145), .ZN(n1140) );
XNOR2_X1 U813 ( .A(n1142), .B(KEYINPUT11), .ZN(n1145) );
XNOR2_X1 U814 ( .A(n1146), .B(n1147), .ZN(n1142) );
NOR3_X1 U815 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NOR2_X1 U816 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U817 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U818 ( .A(KEYINPUT14), .B(KEYINPUT13), .Z(n1154) );
AND2_X1 U819 ( .A1(n1151), .A2(n1153), .ZN(n1149) );
AND2_X1 U820 ( .A1(n1155), .A2(n1156), .ZN(n1151) );
NAND2_X1 U821 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U822 ( .A(KEYINPUT19), .B(n1159), .Z(n1155) );
NOR2_X1 U823 ( .A1(n1158), .A2(n1157), .ZN(n1159) );
XOR2_X1 U824 ( .A(n1160), .B(KEYINPUT7), .Z(n1157) );
NAND2_X1 U825 ( .A1(n1113), .A2(n1161), .ZN(n1146) );
NAND2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
INV_X1 U827 ( .A(n1164), .ZN(n1163) );
XOR2_X1 U828 ( .A(n1165), .B(KEYINPUT9), .Z(n1162) );
NAND2_X1 U829 ( .A1(G898), .A2(G224), .ZN(n1144) );
NOR2_X1 U830 ( .A1(n1166), .A2(n1167), .ZN(G66) );
XOR2_X1 U831 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U832 ( .A1(n1170), .A2(G217), .ZN(n1169) );
NOR2_X1 U833 ( .A1(n1171), .A2(n1172), .ZN(G63) );
XOR2_X1 U834 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U835 ( .A(n1175), .B(KEYINPUT42), .Z(n1173) );
NAND2_X1 U836 ( .A1(n1170), .A2(G478), .ZN(n1175) );
NOR2_X1 U837 ( .A1(G952), .A2(n1176), .ZN(n1171) );
XNOR2_X1 U838 ( .A(G953), .B(KEYINPUT15), .ZN(n1176) );
NOR2_X1 U839 ( .A1(n1166), .A2(n1177), .ZN(G60) );
NOR3_X1 U840 ( .A1(n1108), .A2(n1178), .A3(n1179), .ZN(n1177) );
AND3_X1 U841 ( .A1(n1180), .A2(G475), .A3(n1170), .ZN(n1179) );
NOR2_X1 U842 ( .A1(n1181), .A2(n1180), .ZN(n1178) );
AND2_X1 U843 ( .A1(n1057), .A2(G475), .ZN(n1181) );
INV_X1 U844 ( .A(n1182), .ZN(n1057) );
XNOR2_X1 U845 ( .A(G104), .B(n1183), .ZN(G6) );
NAND2_X1 U846 ( .A1(n1090), .A2(n1184), .ZN(n1183) );
NOR2_X1 U847 ( .A1(n1166), .A2(n1185), .ZN(G57) );
XOR2_X1 U848 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U849 ( .A1(KEYINPUT43), .A2(n1188), .ZN(n1187) );
XOR2_X1 U850 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U851 ( .A(n1191), .B(n1192), .Z(n1189) );
NOR2_X1 U852 ( .A1(KEYINPUT52), .A2(n1193), .ZN(n1192) );
NAND2_X1 U853 ( .A1(n1170), .A2(G472), .ZN(n1191) );
NAND2_X1 U854 ( .A1(n1194), .A2(n1195), .ZN(n1186) );
NAND2_X1 U855 ( .A1(n1196), .A2(G101), .ZN(n1195) );
XOR2_X1 U856 ( .A(KEYINPUT27), .B(n1197), .Z(n1194) );
NOR2_X1 U857 ( .A1(n1196), .A2(G101), .ZN(n1197) );
NOR2_X1 U858 ( .A1(n1166), .A2(n1198), .ZN(G54) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NOR2_X1 U860 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NOR2_X1 U861 ( .A1(n1203), .A2(n1204), .ZN(n1199) );
XOR2_X1 U862 ( .A(KEYINPUT38), .B(n1201), .Z(n1204) );
AND2_X1 U863 ( .A1(n1170), .A2(G469), .ZN(n1201) );
XNOR2_X1 U864 ( .A(n1202), .B(KEYINPUT4), .ZN(n1203) );
XOR2_X1 U865 ( .A(n1205), .B(n1206), .Z(n1202) );
NOR2_X1 U866 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR2_X1 U867 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U868 ( .A(KEYINPUT0), .B(n1211), .Z(n1210) );
AND2_X1 U869 ( .A1(n1209), .A2(n1211), .ZN(n1207) );
XOR2_X1 U870 ( .A(n1212), .B(n1213), .Z(n1209) );
XNOR2_X1 U871 ( .A(n1214), .B(KEYINPUT29), .ZN(n1213) );
NAND2_X1 U872 ( .A1(KEYINPUT22), .A2(n1215), .ZN(n1214) );
INV_X1 U873 ( .A(G110), .ZN(n1215) );
NOR2_X1 U874 ( .A1(n1166), .A2(n1216), .ZN(G51) );
XOR2_X1 U875 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U876 ( .A(n1219), .B(n1220), .Z(n1218) );
NAND2_X1 U877 ( .A1(KEYINPUT40), .A2(n1221), .ZN(n1220) );
INV_X1 U878 ( .A(n1222), .ZN(n1221) );
NAND2_X1 U879 ( .A1(n1170), .A2(n1223), .ZN(n1219) );
NOR2_X1 U880 ( .A1(n1224), .A2(n1182), .ZN(n1170) );
NOR3_X1 U881 ( .A1(n1164), .A2(n1120), .A3(n1165), .ZN(n1182) );
NAND4_X1 U882 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1052), .ZN(n1165) );
NAND2_X1 U883 ( .A1(n1089), .A2(n1184), .ZN(n1052) );
NOR2_X1 U884 ( .A1(n1228), .A2(n1072), .ZN(n1184) );
INV_X1 U885 ( .A(n1229), .ZN(n1072) );
NAND4_X1 U886 ( .A1(n1090), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1225) );
OR2_X1 U887 ( .A1(n1232), .A2(KEYINPUT17), .ZN(n1231) );
NAND2_X1 U888 ( .A1(KEYINPUT17), .A2(n1233), .ZN(n1230) );
NAND3_X1 U889 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NAND4_X1 U890 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1120) );
AND4_X1 U891 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1240) );
AND2_X1 U892 ( .A1(n1245), .A2(n1246), .ZN(n1239) );
NAND4_X1 U893 ( .A1(n1247), .A2(n1074), .A3(n1064), .A4(n1062), .ZN(n1238) );
NAND2_X1 U894 ( .A1(n1248), .A2(n1249), .ZN(n1237) );
XNOR2_X1 U895 ( .A(n1250), .B(KEYINPUT21), .ZN(n1248) );
NAND4_X1 U896 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1164) );
OR2_X1 U897 ( .A1(n1255), .A2(n1234), .ZN(n1251) );
NOR2_X1 U898 ( .A1(n1256), .A2(n1257), .ZN(n1217) );
NOR2_X1 U899 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XNOR2_X1 U900 ( .A(n1260), .B(KEYINPUT32), .ZN(n1259) );
NOR2_X1 U901 ( .A1(n1261), .A2(n1260), .ZN(n1256) );
INV_X1 U902 ( .A(n1258), .ZN(n1261) );
NOR2_X1 U903 ( .A1(n1113), .A2(G952), .ZN(n1166) );
XNOR2_X1 U904 ( .A(G146), .B(n1246), .ZN(G48) );
NAND4_X1 U905 ( .A1(n1262), .A2(n1074), .A3(n1085), .A4(n1082), .ZN(n1246) );
XNOR2_X1 U906 ( .A(G143), .B(n1263), .ZN(G45) );
NAND4_X1 U907 ( .A1(n1064), .A2(n1062), .A3(n1085), .A4(n1264), .ZN(n1263) );
NOR3_X1 U908 ( .A1(n1265), .A2(n1234), .A3(n1266), .ZN(n1264) );
XNOR2_X1 U909 ( .A(KEYINPUT36), .B(n1267), .ZN(n1265) );
XNOR2_X1 U910 ( .A(G140), .B(n1245), .ZN(G42) );
NAND4_X1 U911 ( .A1(n1249), .A2(n1262), .A3(n1268), .A4(n1085), .ZN(n1245) );
INV_X1 U912 ( .A(n1269), .ZN(n1085) );
XOR2_X1 U913 ( .A(n1244), .B(n1270), .Z(G39) );
NOR2_X1 U914 ( .A1(G137), .A2(KEYINPUT24), .ZN(n1270) );
NAND3_X1 U915 ( .A1(n1271), .A2(n1082), .A3(n1272), .ZN(n1244) );
NAND2_X1 U916 ( .A1(n1273), .A2(n1274), .ZN(G36) );
OR2_X1 U917 ( .A1(n1275), .A2(G134), .ZN(n1274) );
XOR2_X1 U918 ( .A(n1276), .B(KEYINPUT62), .Z(n1273) );
NAND2_X1 U919 ( .A1(G134), .A2(n1275), .ZN(n1276) );
NAND2_X1 U920 ( .A1(n1250), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U921 ( .A(KEYINPUT53), .B(n1078), .ZN(n1277) );
AND2_X1 U922 ( .A1(n1247), .A2(n1089), .ZN(n1250) );
NOR3_X1 U923 ( .A1(n1269), .A2(n1278), .A3(n1266), .ZN(n1247) );
INV_X1 U924 ( .A(n1080), .ZN(n1266) );
XNOR2_X1 U925 ( .A(G131), .B(n1243), .ZN(G33) );
NAND3_X1 U926 ( .A1(n1090), .A2(n1080), .A3(n1272), .ZN(n1243) );
NOR3_X1 U927 ( .A1(n1269), .A2(n1278), .A3(n1078), .ZN(n1272) );
INV_X1 U928 ( .A(n1249), .ZN(n1078) );
NOR2_X1 U929 ( .A1(n1075), .A2(n1279), .ZN(n1249) );
INV_X1 U930 ( .A(n1076), .ZN(n1279) );
INV_X1 U931 ( .A(n1267), .ZN(n1278) );
XNOR2_X1 U932 ( .A(G128), .B(n1242), .ZN(G30) );
NAND4_X1 U933 ( .A1(n1267), .A2(n1280), .A3(n1236), .A4(n1281), .ZN(n1242) );
AND3_X1 U934 ( .A1(n1089), .A2(n1082), .A3(n1074), .ZN(n1281) );
XNOR2_X1 U935 ( .A(G101), .B(n1226), .ZN(G3) );
NAND4_X1 U936 ( .A1(n1080), .A2(n1282), .A3(n1283), .A4(n1232), .ZN(n1226) );
XNOR2_X1 U937 ( .A(n1241), .B(n1284), .ZN(G27) );
NOR2_X1 U938 ( .A1(KEYINPUT23), .A2(n1137), .ZN(n1284) );
INV_X1 U939 ( .A(G125), .ZN(n1137) );
NAND4_X1 U940 ( .A1(n1262), .A2(n1285), .A3(n1268), .A4(n1074), .ZN(n1241) );
AND3_X1 U941 ( .A1(n1267), .A2(n1280), .A3(n1090), .ZN(n1262) );
NAND2_X1 U942 ( .A1(n1059), .A2(n1286), .ZN(n1267) );
NAND4_X1 U943 ( .A1(G902), .A2(G953), .A3(n1287), .A4(n1119), .ZN(n1286) );
INV_X1 U944 ( .A(G900), .ZN(n1119) );
XNOR2_X1 U945 ( .A(G122), .B(n1252), .ZN(G24) );
NAND4_X1 U946 ( .A1(n1288), .A2(n1229), .A3(n1064), .A4(n1062), .ZN(n1252) );
NOR2_X1 U947 ( .A1(n1280), .A2(n1082), .ZN(n1229) );
XNOR2_X1 U948 ( .A(G119), .B(n1253), .ZN(G21) );
NAND3_X1 U949 ( .A1(n1271), .A2(n1082), .A3(n1288), .ZN(n1253) );
XNOR2_X1 U950 ( .A(G116), .B(n1289), .ZN(G18) );
NAND2_X1 U951 ( .A1(n1290), .A2(n1074), .ZN(n1289) );
XOR2_X1 U952 ( .A(n1255), .B(KEYINPUT6), .Z(n1290) );
NAND4_X1 U953 ( .A1(n1080), .A2(n1285), .A3(n1089), .A4(n1235), .ZN(n1255) );
NOR2_X1 U954 ( .A1(n1064), .A2(n1282), .ZN(n1089) );
INV_X1 U955 ( .A(n1062), .ZN(n1282) );
NAND2_X1 U956 ( .A1(n1291), .A2(n1292), .ZN(G15) );
OR2_X1 U957 ( .A1(n1254), .A2(G113), .ZN(n1292) );
XOR2_X1 U958 ( .A(n1293), .B(KEYINPUT48), .Z(n1291) );
NAND2_X1 U959 ( .A1(G113), .A2(n1254), .ZN(n1293) );
NAND3_X1 U960 ( .A1(n1090), .A2(n1080), .A3(n1288), .ZN(n1254) );
AND3_X1 U961 ( .A1(n1074), .A2(n1235), .A3(n1285), .ZN(n1288) );
INV_X1 U962 ( .A(n1068), .ZN(n1285) );
NAND2_X1 U963 ( .A1(n1294), .A2(n1087), .ZN(n1068) );
INV_X1 U964 ( .A(n1086), .ZN(n1294) );
NOR2_X1 U965 ( .A1(n1280), .A2(n1268), .ZN(n1080) );
NOR2_X1 U966 ( .A1(n1062), .A2(n1283), .ZN(n1090) );
XNOR2_X1 U967 ( .A(G110), .B(n1227), .ZN(G12) );
NAND3_X1 U968 ( .A1(n1268), .A2(n1232), .A3(n1271), .ZN(n1227) );
NOR3_X1 U969 ( .A1(n1064), .A2(n1081), .A3(n1062), .ZN(n1271) );
NAND2_X1 U970 ( .A1(n1100), .A2(n1295), .ZN(n1062) );
OR2_X1 U971 ( .A1(n1105), .A2(n1104), .ZN(n1295) );
NAND2_X1 U972 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
INV_X1 U973 ( .A(G478), .ZN(n1105) );
NOR2_X1 U974 ( .A1(n1174), .A2(G902), .ZN(n1104) );
XNOR2_X1 U975 ( .A(n1296), .B(n1297), .ZN(n1174) );
XOR2_X1 U976 ( .A(G107), .B(n1298), .Z(n1297) );
XOR2_X1 U977 ( .A(G134), .B(G116), .Z(n1298) );
XOR2_X1 U978 ( .A(n1299), .B(n1300), .Z(n1296) );
XOR2_X1 U979 ( .A(n1301), .B(n1302), .Z(n1299) );
NAND3_X1 U980 ( .A1(G217), .A2(n1303), .A3(KEYINPUT33), .ZN(n1301) );
INV_X1 U981 ( .A(n1280), .ZN(n1081) );
NAND3_X1 U982 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1280) );
OR2_X1 U983 ( .A1(n1168), .A2(n1307), .ZN(n1306) );
NAND3_X1 U984 ( .A1(n1307), .A2(n1168), .A3(n1224), .ZN(n1305) );
NAND2_X1 U985 ( .A1(n1308), .A2(n1309), .ZN(n1168) );
NAND2_X1 U986 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U987 ( .A(KEYINPUT20), .B(n1312), .Z(n1308) );
NOR2_X1 U988 ( .A1(n1310), .A2(n1311), .ZN(n1312) );
XNOR2_X1 U989 ( .A(n1313), .B(n1314), .ZN(n1311) );
XNOR2_X1 U990 ( .A(KEYINPUT26), .B(n1315), .ZN(n1313) );
NOR2_X1 U991 ( .A1(KEYINPUT44), .A2(n1316), .ZN(n1315) );
XOR2_X1 U992 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U993 ( .A(G119), .B(G110), .ZN(n1317) );
XNOR2_X1 U994 ( .A(n1319), .B(n1135), .ZN(n1310) );
NAND2_X1 U995 ( .A1(G221), .A2(n1303), .ZN(n1319) );
NOR2_X1 U996 ( .A1(n1320), .A2(G953), .ZN(n1303) );
NAND2_X1 U997 ( .A1(G217), .A2(n1320), .ZN(n1307) );
INV_X1 U998 ( .A(G234), .ZN(n1320) );
NAND2_X1 U999 ( .A1(G902), .A2(G217), .ZN(n1304) );
INV_X1 U1000 ( .A(n1283), .ZN(n1064) );
XNOR2_X1 U1001 ( .A(n1108), .B(G475), .ZN(n1283) );
NOR2_X1 U1002 ( .A1(n1180), .A2(G902), .ZN(n1108) );
XOR2_X1 U1003 ( .A(n1321), .B(n1322), .Z(n1180) );
XOR2_X1 U1004 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1005 ( .A(G143), .B(G104), .Z(n1324) );
NOR2_X1 U1006 ( .A1(KEYINPUT58), .A2(G131), .ZN(n1323) );
XOR2_X1 U1007 ( .A(n1325), .B(n1314), .Z(n1321) );
XNOR2_X1 U1008 ( .A(n1326), .B(n1327), .ZN(n1314) );
XNOR2_X1 U1009 ( .A(G125), .B(G140), .ZN(n1326) );
XOR2_X1 U1010 ( .A(n1328), .B(n1329), .Z(n1325) );
AND3_X1 U1011 ( .A1(G214), .A2(n1113), .A3(n1330), .ZN(n1329) );
NAND2_X1 U1012 ( .A1(n1331), .A2(KEYINPUT54), .ZN(n1328) );
XNOR2_X1 U1013 ( .A(G113), .B(n1300), .ZN(n1331) );
INV_X1 U1014 ( .A(n1228), .ZN(n1232) );
NAND3_X1 U1015 ( .A1(n1236), .A2(n1235), .A3(n1074), .ZN(n1228) );
INV_X1 U1016 ( .A(n1234), .ZN(n1074) );
NAND2_X1 U1017 ( .A1(n1076), .A2(n1075), .ZN(n1234) );
NAND3_X1 U1018 ( .A1(n1332), .A2(n1333), .A3(n1101), .ZN(n1075) );
NAND2_X1 U1019 ( .A1(n1098), .A2(n1099), .ZN(n1101) );
INV_X1 U1020 ( .A(n1334), .ZN(n1098) );
OR2_X1 U1021 ( .A1(n1223), .A2(KEYINPUT3), .ZN(n1333) );
NAND3_X1 U1022 ( .A1(n1223), .A2(n1334), .A3(KEYINPUT3), .ZN(n1332) );
NAND2_X1 U1023 ( .A1(n1335), .A2(n1224), .ZN(n1334) );
XNOR2_X1 U1024 ( .A(n1260), .B(n1336), .ZN(n1335) );
XNOR2_X1 U1025 ( .A(n1337), .B(n1258), .ZN(n1336) );
NAND2_X1 U1026 ( .A1(G224), .A2(n1113), .ZN(n1258) );
NAND2_X1 U1027 ( .A1(KEYINPUT47), .A2(n1222), .ZN(n1337) );
XNOR2_X1 U1028 ( .A(n1338), .B(n1339), .ZN(n1222) );
XNOR2_X1 U1029 ( .A(n1340), .B(KEYINPUT25), .ZN(n1339) );
NAND2_X1 U1030 ( .A1(KEYINPUT8), .A2(n1160), .ZN(n1340) );
XOR2_X1 U1031 ( .A(n1341), .B(KEYINPUT50), .Z(n1160) );
XNOR2_X1 U1032 ( .A(n1158), .B(n1153), .ZN(n1338) );
XOR2_X1 U1033 ( .A(G110), .B(n1300), .Z(n1153) );
XOR2_X1 U1034 ( .A(G122), .B(KEYINPUT12), .Z(n1300) );
XOR2_X1 U1035 ( .A(n1342), .B(KEYINPUT2), .Z(n1158) );
XNOR2_X1 U1036 ( .A(G125), .B(n1193), .ZN(n1260) );
INV_X1 U1037 ( .A(n1099), .ZN(n1223) );
NAND2_X1 U1038 ( .A1(G210), .A2(n1343), .ZN(n1099) );
NAND2_X1 U1039 ( .A1(G214), .A2(n1343), .ZN(n1076) );
NAND2_X1 U1040 ( .A1(n1330), .A2(n1224), .ZN(n1343) );
NAND2_X1 U1041 ( .A1(n1059), .A2(n1344), .ZN(n1235) );
NAND3_X1 U1042 ( .A1(n1148), .A2(n1287), .A3(G902), .ZN(n1344) );
NOR2_X1 U1043 ( .A1(n1113), .A2(G898), .ZN(n1148) );
NAND3_X1 U1044 ( .A1(n1287), .A2(n1113), .A3(G952), .ZN(n1059) );
NAND2_X1 U1045 ( .A1(G237), .A2(G234), .ZN(n1287) );
XNOR2_X1 U1046 ( .A(n1269), .B(KEYINPUT46), .ZN(n1236) );
NAND2_X1 U1047 ( .A1(n1086), .A2(n1087), .ZN(n1269) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1345), .ZN(n1087) );
NAND2_X1 U1049 ( .A1(G234), .A2(n1224), .ZN(n1345) );
XNOR2_X1 U1050 ( .A(n1346), .B(G469), .ZN(n1086) );
NAND2_X1 U1051 ( .A1(n1347), .A2(n1224), .ZN(n1346) );
XOR2_X1 U1052 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1053 ( .A(n1350), .B(n1211), .Z(n1349) );
AND2_X1 U1054 ( .A1(G227), .A2(n1113), .ZN(n1211) );
NOR2_X1 U1055 ( .A1(KEYINPUT31), .A2(n1351), .ZN(n1350) );
XNOR2_X1 U1056 ( .A(G110), .B(n1212), .ZN(n1351) );
XOR2_X1 U1057 ( .A(G140), .B(KEYINPUT35), .Z(n1212) );
NAND2_X1 U1058 ( .A1(n1352), .A2(n1353), .ZN(n1348) );
NAND3_X1 U1059 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1353) );
INV_X1 U1060 ( .A(KEYINPUT30), .ZN(n1356) );
NAND2_X1 U1061 ( .A1(n1205), .A2(KEYINPUT30), .ZN(n1352) );
XOR2_X1 U1062 ( .A(n1355), .B(n1354), .Z(n1205) );
XNOR2_X1 U1063 ( .A(n1357), .B(n1342), .ZN(n1354) );
XOR2_X1 U1064 ( .A(G101), .B(n1358), .Z(n1342) );
XOR2_X1 U1065 ( .A(G107), .B(G104), .Z(n1358) );
XOR2_X1 U1066 ( .A(n1128), .B(KEYINPUT34), .Z(n1357) );
XOR2_X1 U1067 ( .A(n1193), .B(KEYINPUT59), .Z(n1128) );
INV_X1 U1068 ( .A(n1082), .ZN(n1268) );
XNOR2_X1 U1069 ( .A(n1107), .B(G472), .ZN(n1082) );
NAND2_X1 U1070 ( .A1(n1359), .A2(n1224), .ZN(n1107) );
INV_X1 U1071 ( .A(G902), .ZN(n1224) );
XOR2_X1 U1072 ( .A(n1360), .B(n1361), .Z(n1359) );
XOR2_X1 U1073 ( .A(n1362), .B(n1363), .Z(n1361) );
XNOR2_X1 U1074 ( .A(G101), .B(KEYINPUT16), .ZN(n1363) );
NAND2_X1 U1075 ( .A1(KEYINPUT45), .A2(n1196), .ZN(n1362) );
AND3_X1 U1076 ( .A1(n1330), .A2(n1113), .A3(G210), .ZN(n1196) );
INV_X1 U1077 ( .A(G953), .ZN(n1113) );
INV_X1 U1078 ( .A(G237), .ZN(n1330) );
XOR2_X1 U1079 ( .A(n1190), .B(n1193), .Z(n1360) );
XNOR2_X1 U1080 ( .A(n1327), .B(n1302), .ZN(n1193) );
XOR2_X1 U1081 ( .A(G143), .B(n1318), .Z(n1302) );
XOR2_X1 U1082 ( .A(G128), .B(KEYINPUT5), .Z(n1318) );
XOR2_X1 U1083 ( .A(G146), .B(KEYINPUT56), .Z(n1327) );
XOR2_X1 U1084 ( .A(n1355), .B(n1341), .Z(n1190) );
XOR2_X1 U1085 ( .A(G113), .B(n1364), .Z(n1341) );
XOR2_X1 U1086 ( .A(G119), .B(G116), .Z(n1364) );
XNOR2_X1 U1087 ( .A(n1365), .B(n1366), .ZN(n1355) );
XNOR2_X1 U1088 ( .A(KEYINPUT60), .B(n1135), .ZN(n1366) );
INV_X1 U1089 ( .A(G137), .ZN(n1135) );
XOR2_X1 U1090 ( .A(n1367), .B(G131), .Z(n1365) );
NAND2_X1 U1091 ( .A1(KEYINPUT49), .A2(n1368), .ZN(n1367) );
INV_X1 U1092 ( .A(n1134), .ZN(n1368) );
XOR2_X1 U1093 ( .A(G134), .B(KEYINPUT61), .Z(n1134) );
endmodule


