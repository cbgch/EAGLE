//Key = 0000010100000100110110111000000101011100111111011111101010110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318;

XNOR2_X1 U733 ( .A(G107), .B(n1002), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1003), .A2(n1004), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
XOR2_X1 U736 ( .A(n1009), .B(KEYINPUT2), .Z(n1007) );
NAND3_X1 U737 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1005) );
NAND2_X1 U738 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U739 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND4_X1 U740 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NAND2_X1 U741 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U742 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
INV_X1 U743 ( .A(n1025), .ZN(n1021) );
NAND3_X1 U744 ( .A1(n1023), .A2(n1026), .A3(n1027), .ZN(n1015) );
NAND2_X1 U745 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND3_X1 U746 ( .A1(n1018), .A2(n1030), .A3(n1017), .ZN(n1029) );
OR2_X1 U747 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U748 ( .A1(n1019), .A2(n1033), .ZN(n1028) );
NAND3_X1 U749 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
XNOR2_X1 U751 ( .A(n1017), .B(KEYINPUT47), .ZN(n1037) );
NAND3_X1 U752 ( .A1(n1039), .A2(n1040), .A3(n1017), .ZN(n1035) );
NAND2_X1 U753 ( .A1(n1018), .A2(n1041), .ZN(n1034) );
NAND2_X1 U754 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
INV_X1 U756 ( .A(n1046), .ZN(n1042) );
INV_X1 U757 ( .A(n1047), .ZN(n1013) );
NOR3_X1 U758 ( .A1(n1048), .A2(G953), .A3(G952), .ZN(n1003) );
INV_X1 U759 ( .A(n1010), .ZN(n1048) );
NAND4_X1 U760 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1010) );
NOR4_X1 U761 ( .A1(n1039), .A2(n1053), .A3(n1044), .A4(n1054), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U763 ( .A(KEYINPUT5), .B(n1057), .Z(n1056) );
INV_X1 U764 ( .A(n1058), .ZN(n1055) );
NOR2_X1 U765 ( .A1(n1059), .A2(n1060), .ZN(n1051) );
XNOR2_X1 U766 ( .A(G472), .B(n1061), .ZN(n1060) );
XOR2_X1 U767 ( .A(n1062), .B(n1063), .Z(G72) );
NAND2_X1 U768 ( .A1(G953), .A2(n1064), .ZN(n1063) );
NAND2_X1 U769 ( .A1(G900), .A2(G227), .ZN(n1064) );
NAND4_X1 U770 ( .A1(KEYINPUT24), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1062) );
NAND3_X1 U771 ( .A1(n1068), .A2(n1009), .A3(n1011), .ZN(n1067) );
NAND2_X1 U772 ( .A1(G953), .A2(n1069), .ZN(n1066) );
NAND2_X1 U773 ( .A1(G900), .A2(n1068), .ZN(n1069) );
OR2_X1 U774 ( .A1(n1009), .A2(n1068), .ZN(n1065) );
XOR2_X1 U775 ( .A(n1070), .B(n1071), .Z(n1068) );
XOR2_X1 U776 ( .A(n1072), .B(n1073), .Z(n1071) );
NAND2_X1 U777 ( .A1(KEYINPUT36), .A2(n1074), .ZN(n1073) );
XNOR2_X1 U778 ( .A(n1075), .B(G134), .ZN(n1074) );
INV_X1 U779 ( .A(G137), .ZN(n1075) );
XOR2_X1 U780 ( .A(n1076), .B(n1077), .Z(G69) );
NOR2_X1 U781 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U782 ( .A1(G953), .A2(n1080), .ZN(n1079) );
NOR2_X1 U783 ( .A1(n1006), .A2(n1081), .ZN(n1080) );
XNOR2_X1 U784 ( .A(KEYINPUT45), .B(n1008), .ZN(n1081) );
NOR2_X1 U785 ( .A1(n1082), .A2(n1011), .ZN(n1078) );
NOR2_X1 U786 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
INV_X1 U787 ( .A(G224), .ZN(n1084) );
XNOR2_X1 U788 ( .A(G898), .B(KEYINPUT14), .ZN(n1083) );
NAND2_X1 U789 ( .A1(n1085), .A2(n1086), .ZN(n1076) );
NAND2_X1 U790 ( .A1(G953), .A2(n1087), .ZN(n1086) );
XNOR2_X1 U791 ( .A(n1088), .B(n1089), .ZN(n1085) );
XOR2_X1 U792 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U793 ( .A1(n1092), .A2(KEYINPUT38), .ZN(n1090) );
NOR2_X1 U794 ( .A1(n1093), .A2(n1094), .ZN(G66) );
XOR2_X1 U795 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U796 ( .A1(n1097), .A2(n1057), .ZN(n1095) );
NOR2_X1 U797 ( .A1(n1093), .A2(n1098), .ZN(G63) );
XOR2_X1 U798 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U799 ( .A1(n1097), .A2(G478), .ZN(n1099) );
NOR2_X1 U800 ( .A1(n1093), .A2(n1101), .ZN(G60) );
XOR2_X1 U801 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND3_X1 U802 ( .A1(n1097), .A2(G475), .A3(KEYINPUT50), .ZN(n1102) );
XNOR2_X1 U803 ( .A(G104), .B(n1104), .ZN(G6) );
NOR2_X1 U804 ( .A1(n1093), .A2(n1105), .ZN(G57) );
XOR2_X1 U805 ( .A(n1106), .B(n1107), .Z(n1105) );
XNOR2_X1 U806 ( .A(G101), .B(n1108), .ZN(n1107) );
NAND2_X1 U807 ( .A1(n1109), .A2(KEYINPUT49), .ZN(n1106) );
XOR2_X1 U808 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U809 ( .A(n1112), .B(n1091), .Z(n1111) );
NAND2_X1 U810 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U811 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
INV_X1 U812 ( .A(KEYINPUT11), .ZN(n1116) );
XOR2_X1 U813 ( .A(n1117), .B(n1118), .Z(n1115) );
NAND3_X1 U814 ( .A1(n1118), .A2(n1117), .A3(KEYINPUT11), .ZN(n1113) );
XOR2_X1 U815 ( .A(n1119), .B(n1120), .Z(n1110) );
NAND2_X1 U816 ( .A1(n1097), .A2(G472), .ZN(n1119) );
NOR2_X1 U817 ( .A1(n1093), .A2(n1121), .ZN(G54) );
XOR2_X1 U818 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U819 ( .A(n1124), .B(n1125), .ZN(n1123) );
NOR2_X1 U820 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
XOR2_X1 U821 ( .A(KEYINPUT8), .B(n1128), .Z(n1127) );
NOR2_X1 U822 ( .A1(n1117), .A2(n1129), .ZN(n1128) );
AND2_X1 U823 ( .A1(n1129), .A2(n1117), .ZN(n1126) );
NAND3_X1 U824 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
NAND2_X1 U825 ( .A1(KEYINPUT3), .A2(n1133), .ZN(n1132) );
INV_X1 U826 ( .A(n1134), .ZN(n1133) );
OR3_X1 U827 ( .A1(n1135), .A2(KEYINPUT3), .A3(n1136), .ZN(n1131) );
NAND2_X1 U828 ( .A1(n1136), .A2(n1135), .ZN(n1130) );
NAND2_X1 U829 ( .A1(KEYINPUT41), .A2(n1134), .ZN(n1135) );
XNOR2_X1 U830 ( .A(n1072), .B(KEYINPUT16), .ZN(n1134) );
XOR2_X1 U831 ( .A(n1137), .B(n1138), .Z(n1122) );
NAND3_X1 U832 ( .A1(n1097), .A2(G469), .A3(KEYINPUT61), .ZN(n1137) );
NOR2_X1 U833 ( .A1(n1093), .A2(n1139), .ZN(G51) );
XOR2_X1 U834 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U835 ( .A(n1142), .B(KEYINPUT20), .Z(n1141) );
NAND2_X1 U836 ( .A1(n1097), .A2(G210), .ZN(n1142) );
AND2_X1 U837 ( .A1(G902), .A2(n1143), .ZN(n1097) );
OR3_X1 U838 ( .A1(n1008), .A2(n1009), .A3(n1006), .ZN(n1143) );
NAND4_X1 U839 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1006) );
NAND4_X1 U840 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1009) );
AND4_X1 U841 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1151) );
AND2_X1 U842 ( .A1(n1156), .A2(n1157), .ZN(n1150) );
NAND2_X1 U843 ( .A1(n1158), .A2(n1017), .ZN(n1148) );
XOR2_X1 U844 ( .A(n1159), .B(KEYINPUT62), .Z(n1158) );
NAND4_X1 U845 ( .A1(n1160), .A2(n1104), .A3(n1161), .A4(n1002), .ZN(n1008) );
NAND3_X1 U846 ( .A1(n1032), .A2(n1162), .A3(n1027), .ZN(n1002) );
NAND3_X1 U847 ( .A1(n1027), .A2(n1162), .A3(n1031), .ZN(n1104) );
NAND3_X1 U848 ( .A1(n1019), .A2(n1163), .A3(n1164), .ZN(n1160) );
NOR2_X1 U849 ( .A1(n1011), .A2(G952), .ZN(n1093) );
XOR2_X1 U850 ( .A(n1156), .B(n1165), .Z(G48) );
XNOR2_X1 U851 ( .A(G146), .B(KEYINPUT1), .ZN(n1165) );
NAND3_X1 U852 ( .A1(n1031), .A2(n1046), .A3(n1166), .ZN(n1156) );
XNOR2_X1 U853 ( .A(G143), .B(n1155), .ZN(G45) );
NAND3_X1 U854 ( .A1(n1164), .A2(n1046), .A3(n1167), .ZN(n1155) );
NOR3_X1 U855 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
XOR2_X1 U856 ( .A(G140), .B(n1171), .Z(G42) );
NOR2_X1 U857 ( .A1(n1172), .A2(n1159), .ZN(n1171) );
NAND3_X1 U858 ( .A1(n1023), .A2(n1031), .A3(n1173), .ZN(n1159) );
XNOR2_X1 U859 ( .A(G137), .B(n1154), .ZN(G39) );
NAND3_X1 U860 ( .A1(n1017), .A2(n1019), .A3(n1166), .ZN(n1154) );
XOR2_X1 U861 ( .A(n1153), .B(n1174), .Z(G36) );
XNOR2_X1 U862 ( .A(G134), .B(KEYINPUT46), .ZN(n1174) );
NAND4_X1 U863 ( .A1(n1017), .A2(n1164), .A3(n1032), .A4(n1175), .ZN(n1153) );
NAND2_X1 U864 ( .A1(n1176), .A2(n1177), .ZN(G33) );
OR2_X1 U865 ( .A1(n1149), .A2(G131), .ZN(n1177) );
XOR2_X1 U866 ( .A(n1178), .B(KEYINPUT39), .Z(n1176) );
NAND2_X1 U867 ( .A1(G131), .A2(n1149), .ZN(n1178) );
NAND4_X1 U868 ( .A1(n1017), .A2(n1164), .A3(n1031), .A4(n1175), .ZN(n1149) );
INV_X1 U869 ( .A(n1179), .ZN(n1164) );
INV_X1 U870 ( .A(n1172), .ZN(n1017) );
NAND2_X1 U871 ( .A1(n1045), .A2(n1180), .ZN(n1172) );
XNOR2_X1 U872 ( .A(n1050), .B(KEYINPUT33), .ZN(n1045) );
XNOR2_X1 U873 ( .A(G128), .B(n1152), .ZN(G30) );
NAND3_X1 U874 ( .A1(n1032), .A2(n1046), .A3(n1166), .ZN(n1152) );
AND2_X1 U875 ( .A1(n1173), .A2(n1181), .ZN(n1166) );
AND3_X1 U876 ( .A1(n1175), .A2(n1024), .A3(n1038), .ZN(n1173) );
XNOR2_X1 U877 ( .A(n1182), .B(n1183), .ZN(G3) );
NOR4_X1 U878 ( .A1(KEYINPUT6), .A2(n1184), .A3(n1059), .A4(n1179), .ZN(n1183) );
NAND2_X1 U879 ( .A1(n1025), .A2(n1038), .ZN(n1179) );
XOR2_X1 U880 ( .A(G125), .B(n1185), .Z(G27) );
NOR2_X1 U881 ( .A1(KEYINPUT53), .A2(n1157), .ZN(n1185) );
NAND4_X1 U882 ( .A1(n1018), .A2(n1046), .A3(n1031), .A4(n1186), .ZN(n1157) );
NOR3_X1 U883 ( .A1(n1187), .A2(n1027), .A3(n1169), .ZN(n1186) );
INV_X1 U884 ( .A(n1175), .ZN(n1169) );
NAND2_X1 U885 ( .A1(n1047), .A2(n1188), .ZN(n1175) );
NAND4_X1 U886 ( .A1(G953), .A2(G902), .A3(n1189), .A4(n1190), .ZN(n1188) );
INV_X1 U887 ( .A(G900), .ZN(n1190) );
XNOR2_X1 U888 ( .A(G122), .B(n1144), .ZN(G24) );
NAND3_X1 U889 ( .A1(n1191), .A2(n1027), .A3(n1192), .ZN(n1144) );
NOR3_X1 U890 ( .A1(n1187), .A2(n1170), .A3(n1168), .ZN(n1192) );
XOR2_X1 U891 ( .A(n1145), .B(n1193), .Z(G21) );
NAND2_X1 U892 ( .A1(KEYINPUT7), .A2(G119), .ZN(n1193) );
NAND4_X1 U893 ( .A1(n1191), .A2(n1019), .A3(n1181), .A4(n1024), .ZN(n1145) );
XNOR2_X1 U894 ( .A(G116), .B(n1146), .ZN(G18) );
NAND3_X1 U895 ( .A1(n1191), .A2(n1032), .A3(n1025), .ZN(n1146) );
NOR2_X1 U896 ( .A1(n1194), .A2(n1168), .ZN(n1032) );
XNOR2_X1 U897 ( .A(G113), .B(n1147), .ZN(G15) );
NAND3_X1 U898 ( .A1(n1031), .A2(n1191), .A3(n1025), .ZN(n1147) );
NOR2_X1 U899 ( .A1(n1024), .A2(n1195), .ZN(n1025) );
AND2_X1 U900 ( .A1(n1018), .A2(n1163), .ZN(n1191) );
AND2_X1 U901 ( .A1(n1196), .A2(n1040), .ZN(n1018) );
XOR2_X1 U902 ( .A(n1197), .B(KEYINPUT58), .Z(n1040) );
AND2_X1 U903 ( .A1(n1168), .A2(n1194), .ZN(n1031) );
NAND2_X1 U904 ( .A1(n1198), .A2(n1199), .ZN(G12) );
NAND2_X1 U905 ( .A1(G110), .A2(n1161), .ZN(n1199) );
XOR2_X1 U906 ( .A(KEYINPUT19), .B(n1200), .Z(n1198) );
NOR2_X1 U907 ( .A1(G110), .A2(n1161), .ZN(n1200) );
NAND3_X1 U908 ( .A1(n1162), .A2(n1024), .A3(n1019), .ZN(n1161) );
INV_X1 U909 ( .A(n1059), .ZN(n1019) );
NAND2_X1 U910 ( .A1(n1168), .A2(n1170), .ZN(n1059) );
INV_X1 U911 ( .A(n1194), .ZN(n1170) );
XNOR2_X1 U912 ( .A(n1201), .B(G475), .ZN(n1194) );
NAND2_X1 U913 ( .A1(n1103), .A2(n1202), .ZN(n1201) );
XNOR2_X1 U914 ( .A(n1203), .B(n1204), .ZN(n1103) );
XOR2_X1 U915 ( .A(n1070), .B(n1205), .Z(n1204) );
XOR2_X1 U916 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U917 ( .A1(G146), .A2(KEYINPUT60), .ZN(n1207) );
NAND2_X1 U918 ( .A1(G214), .A2(n1208), .ZN(n1206) );
XOR2_X1 U919 ( .A(n1209), .B(n1210), .Z(n1070) );
XOR2_X1 U920 ( .A(n1211), .B(n1212), .Z(n1203) );
XNOR2_X1 U921 ( .A(KEYINPUT48), .B(n1213), .ZN(n1212) );
XOR2_X1 U922 ( .A(n1214), .B(G104), .Z(n1211) );
NAND2_X1 U923 ( .A1(n1215), .A2(KEYINPUT37), .ZN(n1214) );
XNOR2_X1 U924 ( .A(G113), .B(G122), .ZN(n1215) );
XOR2_X1 U925 ( .A(n1216), .B(G478), .Z(n1168) );
NAND2_X1 U926 ( .A1(n1100), .A2(n1202), .ZN(n1216) );
XOR2_X1 U927 ( .A(n1217), .B(n1218), .Z(n1100) );
XOR2_X1 U928 ( .A(n1219), .B(n1220), .Z(n1218) );
NAND2_X1 U929 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND3_X1 U930 ( .A1(n1213), .A2(n1223), .A3(n1224), .ZN(n1222) );
XNOR2_X1 U931 ( .A(n1225), .B(n1226), .ZN(n1224) );
INV_X1 U932 ( .A(G134), .ZN(n1226) );
NAND2_X1 U933 ( .A1(KEYINPUT63), .A2(G128), .ZN(n1225) );
NAND2_X1 U934 ( .A1(n1227), .A2(n1228), .ZN(n1221) );
NAND2_X1 U935 ( .A1(n1213), .A2(n1223), .ZN(n1228) );
INV_X1 U936 ( .A(KEYINPUT32), .ZN(n1223) );
INV_X1 U937 ( .A(G143), .ZN(n1213) );
XNOR2_X1 U938 ( .A(G134), .B(n1229), .ZN(n1227) );
AND2_X1 U939 ( .A1(n1230), .A2(KEYINPUT63), .ZN(n1229) );
NAND3_X1 U940 ( .A1(n1231), .A2(n1011), .A3(n1232), .ZN(n1219) );
XNOR2_X1 U941 ( .A(G217), .B(KEYINPUT51), .ZN(n1232) );
NAND2_X1 U942 ( .A1(n1233), .A2(n1234), .ZN(n1217) );
NAND2_X1 U943 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XNOR2_X1 U944 ( .A(n1237), .B(KEYINPUT35), .ZN(n1235) );
NAND2_X1 U945 ( .A1(n1238), .A2(G107), .ZN(n1233) );
XOR2_X1 U946 ( .A(KEYINPUT52), .B(n1237), .Z(n1238) );
XNOR2_X1 U947 ( .A(G116), .B(n1239), .ZN(n1237) );
INV_X1 U948 ( .A(G122), .ZN(n1239) );
INV_X1 U949 ( .A(n1027), .ZN(n1024) );
NOR2_X1 U950 ( .A1(n1240), .A2(n1053), .ZN(n1027) );
NOR2_X1 U951 ( .A1(n1058), .A2(n1057), .ZN(n1053) );
AND2_X1 U952 ( .A1(n1241), .A2(n1058), .ZN(n1240) );
NAND2_X1 U953 ( .A1(n1242), .A2(n1096), .ZN(n1058) );
XNOR2_X1 U954 ( .A(n1243), .B(n1244), .ZN(n1096) );
XNOR2_X1 U955 ( .A(G137), .B(n1245), .ZN(n1244) );
NAND3_X1 U956 ( .A1(n1231), .A2(n1011), .A3(G221), .ZN(n1245) );
XOR2_X1 U957 ( .A(G234), .B(KEYINPUT10), .Z(n1231) );
NAND2_X1 U958 ( .A1(n1246), .A2(KEYINPUT56), .ZN(n1243) );
XOR2_X1 U959 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U960 ( .A(G146), .B(G110), .Z(n1248) );
XOR2_X1 U961 ( .A(n1249), .B(n1209), .Z(n1247) );
XOR2_X1 U962 ( .A(G125), .B(G140), .Z(n1209) );
NAND2_X1 U963 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND2_X1 U964 ( .A1(G119), .A2(n1230), .ZN(n1251) );
XOR2_X1 U965 ( .A(KEYINPUT43), .B(n1252), .Z(n1250) );
NOR2_X1 U966 ( .A1(G119), .A2(n1230), .ZN(n1252) );
XNOR2_X1 U967 ( .A(KEYINPUT22), .B(n1202), .ZN(n1242) );
XOR2_X1 U968 ( .A(KEYINPUT57), .B(n1057), .Z(n1241) );
AND2_X1 U969 ( .A1(G217), .A2(n1253), .ZN(n1057) );
AND3_X1 U970 ( .A1(n1023), .A2(n1163), .A3(n1038), .ZN(n1162) );
AND2_X1 U971 ( .A1(n1196), .A2(n1197), .ZN(n1038) );
XNOR2_X1 U972 ( .A(n1049), .B(KEYINPUT34), .ZN(n1197) );
XNOR2_X1 U973 ( .A(G469), .B(n1254), .ZN(n1049) );
NOR2_X1 U974 ( .A1(G902), .A2(n1255), .ZN(n1254) );
XOR2_X1 U975 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U976 ( .A(n1258), .B(n1138), .Z(n1257) );
XOR2_X1 U977 ( .A(G140), .B(G110), .Z(n1138) );
NOR2_X1 U978 ( .A1(KEYINPUT15), .A2(n1125), .ZN(n1258) );
NAND2_X1 U979 ( .A1(G227), .A2(n1011), .ZN(n1125) );
XOR2_X1 U980 ( .A(n1117), .B(n1259), .Z(n1256) );
NOR2_X1 U981 ( .A1(KEYINPUT27), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U982 ( .A(n1136), .B(n1261), .ZN(n1260) );
NAND2_X1 U983 ( .A1(KEYINPUT17), .A2(n1072), .ZN(n1261) );
NAND3_X1 U984 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1072) );
NAND2_X1 U985 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
INV_X1 U986 ( .A(KEYINPUT23), .ZN(n1266) );
NAND3_X1 U987 ( .A1(KEYINPUT23), .A2(n1267), .A3(n1268), .ZN(n1263) );
OR2_X1 U988 ( .A1(n1268), .A2(n1267), .ZN(n1262) );
NOR2_X1 U989 ( .A1(KEYINPUT30), .A2(n1265), .ZN(n1267) );
XOR2_X1 U990 ( .A(n1269), .B(KEYINPUT44), .Z(n1268) );
AND3_X1 U991 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1136) );
NAND2_X1 U992 ( .A1(n1273), .A2(n1182), .ZN(n1271) );
XNOR2_X1 U993 ( .A(G107), .B(n1274), .ZN(n1273) );
NOR2_X1 U994 ( .A1(KEYINPUT29), .A2(n1275), .ZN(n1274) );
NAND3_X1 U995 ( .A1(n1276), .A2(n1277), .A3(G101), .ZN(n1270) );
XNOR2_X1 U996 ( .A(KEYINPUT29), .B(G107), .ZN(n1276) );
XNOR2_X1 U997 ( .A(n1039), .B(KEYINPUT4), .ZN(n1196) );
AND2_X1 U998 ( .A1(G221), .A2(n1253), .ZN(n1039) );
NAND2_X1 U999 ( .A1(G234), .A2(n1202), .ZN(n1253) );
INV_X1 U1000 ( .A(n1184), .ZN(n1163) );
NAND2_X1 U1001 ( .A1(n1046), .A2(n1278), .ZN(n1184) );
NAND2_X1 U1002 ( .A1(n1279), .A2(n1047), .ZN(n1278) );
NAND3_X1 U1003 ( .A1(n1189), .A2(n1011), .A3(G952), .ZN(n1047) );
NAND4_X1 U1004 ( .A1(G953), .A2(G902), .A3(n1189), .A4(n1087), .ZN(n1279) );
INV_X1 U1005 ( .A(G898), .ZN(n1087) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1189) );
NOR2_X1 U1007 ( .A1(n1050), .A2(n1044), .ZN(n1046) );
INV_X1 U1008 ( .A(n1180), .ZN(n1044) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1280), .ZN(n1180) );
OR2_X1 U1010 ( .A1(G237), .A2(G902), .ZN(n1280) );
AND3_X1 U1011 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1050) );
NAND2_X1 U1012 ( .A1(G210), .A2(G902), .ZN(n1283) );
NAND3_X1 U1013 ( .A1(n1284), .A2(n1202), .A3(n1285), .ZN(n1282) );
OR2_X1 U1014 ( .A1(n1284), .A2(n1285), .ZN(n1281) );
NAND2_X1 U1015 ( .A1(G237), .A2(G210), .ZN(n1285) );
XOR2_X1 U1016 ( .A(n1140), .B(n1286), .Z(n1284) );
XOR2_X1 U1017 ( .A(KEYINPUT31), .B(KEYINPUT21), .Z(n1286) );
XOR2_X1 U1018 ( .A(n1287), .B(n1288), .Z(n1140) );
XOR2_X1 U1019 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U1020 ( .A(G125), .B(KEYINPUT13), .ZN(n1290) );
NAND2_X1 U1021 ( .A1(n1291), .A2(n1011), .ZN(n1289) );
INV_X1 U1022 ( .A(G953), .ZN(n1011) );
XNOR2_X1 U1023 ( .A(G224), .B(KEYINPUT40), .ZN(n1291) );
XNOR2_X1 U1024 ( .A(n1292), .B(n1293), .ZN(n1287) );
INV_X1 U1025 ( .A(n1088), .ZN(n1293) );
XNOR2_X1 U1026 ( .A(n1294), .B(n1295), .ZN(n1088) );
NOR2_X1 U1027 ( .A1(KEYINPUT25), .A2(G122), .ZN(n1295) );
XNOR2_X1 U1028 ( .A(G110), .B(G116), .ZN(n1294) );
XNOR2_X1 U1029 ( .A(n1092), .B(n1296), .ZN(n1292) );
AND3_X1 U1030 ( .A1(n1297), .A2(n1298), .A3(n1272), .ZN(n1092) );
NAND3_X1 U1031 ( .A1(G107), .A2(n1275), .A3(G101), .ZN(n1272) );
NAND2_X1 U1032 ( .A1(n1299), .A2(n1236), .ZN(n1298) );
INV_X1 U1033 ( .A(G107), .ZN(n1236) );
XNOR2_X1 U1034 ( .A(n1182), .B(n1275), .ZN(n1299) );
NAND3_X1 U1035 ( .A1(n1277), .A2(n1182), .A3(G107), .ZN(n1297) );
INV_X1 U1036 ( .A(n1275), .ZN(n1277) );
XOR2_X1 U1037 ( .A(G104), .B(KEYINPUT59), .Z(n1275) );
INV_X1 U1038 ( .A(n1187), .ZN(n1023) );
XOR2_X1 U1039 ( .A(n1181), .B(KEYINPUT9), .Z(n1187) );
INV_X1 U1040 ( .A(n1195), .ZN(n1181) );
NAND2_X1 U1041 ( .A1(n1300), .A2(n1301), .ZN(n1195) );
NAND2_X1 U1042 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n1303) );
XOR2_X1 U1044 ( .A(n1061), .B(G472), .Z(n1302) );
NAND3_X1 U1045 ( .A1(G472), .A2(n1061), .A3(KEYINPUT55), .ZN(n1300) );
NAND2_X1 U1046 ( .A1(n1304), .A2(n1202), .ZN(n1061) );
INV_X1 U1047 ( .A(G902), .ZN(n1202) );
XOR2_X1 U1048 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1049 ( .A(n1117), .B(n1296), .ZN(n1306) );
XOR2_X1 U1050 ( .A(n1091), .B(n1118), .Z(n1296) );
XNOR2_X1 U1051 ( .A(n1269), .B(n1265), .ZN(n1118) );
XNOR2_X1 U1052 ( .A(n1230), .B(KEYINPUT18), .ZN(n1265) );
INV_X1 U1053 ( .A(G128), .ZN(n1230) );
XNOR2_X1 U1054 ( .A(G143), .B(G146), .ZN(n1269) );
XOR2_X1 U1055 ( .A(G113), .B(G119), .Z(n1091) );
NAND2_X1 U1056 ( .A1(n1307), .A2(n1308), .ZN(n1117) );
NAND2_X1 U1057 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND2_X1 U1058 ( .A1(KEYINPUT54), .A2(n1311), .ZN(n1310) );
OR2_X1 U1059 ( .A1(n1210), .A2(KEYINPUT28), .ZN(n1311) );
INV_X1 U1060 ( .A(n1312), .ZN(n1309) );
NAND2_X1 U1061 ( .A1(n1210), .A2(n1313), .ZN(n1307) );
NAND2_X1 U1062 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND2_X1 U1063 ( .A1(KEYINPUT54), .A2(n1312), .ZN(n1315) );
XOR2_X1 U1064 ( .A(G137), .B(n1316), .Z(n1312) );
NOR2_X1 U1065 ( .A1(G134), .A2(KEYINPUT12), .ZN(n1316) );
INV_X1 U1066 ( .A(KEYINPUT28), .ZN(n1314) );
XNOR2_X1 U1067 ( .A(G131), .B(KEYINPUT42), .ZN(n1210) );
XOR2_X1 U1068 ( .A(n1317), .B(n1318), .Z(n1305) );
XNOR2_X1 U1069 ( .A(n1182), .B(n1120), .ZN(n1318) );
NOR2_X1 U1070 ( .A1(KEYINPUT26), .A2(G116), .ZN(n1120) );
INV_X1 U1071 ( .A(G101), .ZN(n1182) );
NOR2_X1 U1072 ( .A1(KEYINPUT0), .A2(n1108), .ZN(n1317) );
NAND2_X1 U1073 ( .A1(G210), .A2(n1208), .ZN(n1108) );
NOR2_X1 U1074 ( .A1(G953), .A2(G237), .ZN(n1208) );
endmodule


