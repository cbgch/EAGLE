//Key = 1011001001100100111010000011111001100111100001100100111011001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335;

XNOR2_X1 U737 ( .A(G107), .B(n1020), .ZN(G9) );
NOR2_X1 U738 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR2_X1 U739 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND4_X1 U740 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
NAND3_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND2_X1 U742 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND3_X1 U743 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NAND2_X1 U745 ( .A1(n1039), .A2(n1040), .ZN(n1032) );
NAND2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1043), .ZN(n1042) );
NAND2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U749 ( .A1(n1034), .A2(n1046), .ZN(n1041) );
NAND2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1027) );
XNOR2_X1 U753 ( .A(n1053), .B(KEYINPUT27), .ZN(n1051) );
XNOR2_X1 U754 ( .A(n1054), .B(KEYINPUT39), .ZN(n1025) );
NAND4_X1 U755 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1023) );
NAND3_X1 U756 ( .A1(n1059), .A2(n1060), .A3(n1053), .ZN(n1055) );
AND4_X1 U757 ( .A1(n1029), .A2(n1036), .A3(n1039), .A4(n1034), .ZN(n1053) );
INV_X1 U758 ( .A(n1061), .ZN(n1029) );
NOR3_X1 U759 ( .A1(n1062), .A2(G953), .A3(G952), .ZN(n1021) );
INV_X1 U760 ( .A(n1057), .ZN(n1062) );
NAND4_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1057) );
NOR4_X1 U762 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
XOR2_X1 U763 ( .A(KEYINPUT18), .B(n1071), .Z(n1070) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U765 ( .A(KEYINPUT12), .B(n1074), .Z(n1073) );
NOR2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XNOR2_X1 U767 ( .A(KEYINPUT3), .B(n1077), .ZN(n1076) );
NOR3_X1 U768 ( .A1(n1060), .A2(n1078), .A3(n1079), .ZN(n1065) );
XOR2_X1 U769 ( .A(n1080), .B(n1081), .Z(G72) );
NOR2_X1 U770 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U771 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U772 ( .A(n1086), .B(n1087), .ZN(n1085) );
XNOR2_X1 U773 ( .A(n1088), .B(n1089), .ZN(n1084) );
NOR2_X1 U774 ( .A1(G900), .A2(n1058), .ZN(n1082) );
NAND3_X1 U775 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1080) );
OR2_X1 U776 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND3_X1 U777 ( .A1(n1094), .A2(n1093), .A3(G953), .ZN(n1091) );
NAND2_X1 U778 ( .A1(G900), .A2(G227), .ZN(n1094) );
NAND2_X1 U779 ( .A1(n1095), .A2(n1058), .ZN(n1090) );
NAND4_X1 U780 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1093), .ZN(n1095) );
INV_X1 U781 ( .A(KEYINPUT32), .ZN(n1093) );
XOR2_X1 U782 ( .A(n1099), .B(n1100), .Z(G69) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
AND2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR3_X1 U785 ( .A1(n1103), .A2(n1105), .A3(n1104), .ZN(n1101) );
XNOR2_X1 U786 ( .A(n1106), .B(n1107), .ZN(n1104) );
XOR2_X1 U787 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U788 ( .A(n1110), .B(KEYINPUT53), .Z(n1106) );
NOR2_X1 U789 ( .A1(G898), .A2(n1058), .ZN(n1105) );
AND2_X1 U790 ( .A1(n1111), .A2(n1058), .ZN(n1103) );
NAND2_X1 U791 ( .A1(n1026), .A2(n1112), .ZN(n1111) );
XNOR2_X1 U792 ( .A(KEYINPUT33), .B(n1056), .ZN(n1112) );
NAND3_X1 U793 ( .A1(G953), .A2(n1113), .A3(KEYINPUT20), .ZN(n1099) );
NAND2_X1 U794 ( .A1(G898), .A2(G224), .ZN(n1113) );
NOR2_X1 U795 ( .A1(n1114), .A2(n1115), .ZN(G66) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U797 ( .A(KEYINPUT28), .B(n1118), .Z(n1117) );
NOR2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR3_X1 U799 ( .A1(n1114), .A2(n1121), .A3(n1122), .ZN(G63) );
NOR3_X1 U800 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
NOR2_X1 U801 ( .A1(KEYINPUT52), .A2(n1126), .ZN(n1125) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1128), .ZN(n1121) );
INV_X1 U803 ( .A(n1123), .ZN(n1128) );
NOR2_X1 U804 ( .A1(n1126), .A2(n1129), .ZN(n1127) );
INV_X1 U805 ( .A(KEYINPUT52), .ZN(n1129) );
XNOR2_X1 U806 ( .A(n1124), .B(KEYINPUT34), .ZN(n1126) );
AND2_X1 U807 ( .A1(n1130), .A2(G478), .ZN(n1124) );
NOR2_X1 U808 ( .A1(n1114), .A2(n1131), .ZN(G60) );
XNOR2_X1 U809 ( .A(n1132), .B(n1133), .ZN(n1131) );
AND2_X1 U810 ( .A1(G475), .A2(n1130), .ZN(n1133) );
XNOR2_X1 U811 ( .A(G104), .B(n1134), .ZN(G6) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(G57) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U814 ( .A(n1139), .B(n1140), .ZN(n1138) );
NOR2_X1 U815 ( .A1(KEYINPUT58), .A2(n1141), .ZN(n1140) );
NAND3_X1 U816 ( .A1(KEYINPUT17), .A2(n1130), .A3(n1142), .ZN(n1139) );
XNOR2_X1 U817 ( .A(G472), .B(KEYINPUT37), .ZN(n1142) );
XNOR2_X1 U818 ( .A(n1114), .B(KEYINPUT6), .ZN(n1135) );
NOR3_X1 U819 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(G54) );
AND2_X1 U820 ( .A1(KEYINPUT49), .A2(n1114), .ZN(n1145) );
NOR3_X1 U821 ( .A1(KEYINPUT49), .A2(G953), .A3(G952), .ZN(n1144) );
XOR2_X1 U822 ( .A(n1146), .B(n1147), .Z(n1143) );
AND2_X1 U823 ( .A1(G469), .A2(n1130), .ZN(n1147) );
INV_X1 U824 ( .A(n1120), .ZN(n1130) );
NOR2_X1 U825 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
XOR2_X1 U826 ( .A(n1150), .B(KEYINPUT40), .Z(n1149) );
NAND4_X1 U827 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
NAND3_X1 U828 ( .A1(n1155), .A2(n1089), .A3(n1156), .ZN(n1154) );
OR2_X1 U829 ( .A1(n1156), .A2(n1155), .ZN(n1153) );
INV_X1 U830 ( .A(KEYINPUT62), .ZN(n1156) );
INV_X1 U831 ( .A(n1157), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1158), .A2(n1151), .ZN(n1148) );
NOR2_X1 U833 ( .A1(n1157), .A2(n1159), .ZN(n1158) );
NOR2_X1 U834 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XNOR2_X1 U835 ( .A(n1155), .B(KEYINPUT62), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1089), .ZN(n1157) );
XNOR2_X1 U837 ( .A(n1162), .B(n1163), .ZN(n1155) );
NAND2_X1 U838 ( .A1(KEYINPUT38), .A2(n1164), .ZN(n1162) );
NOR2_X1 U839 ( .A1(n1114), .A2(n1165), .ZN(G51) );
XOR2_X1 U840 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(n1166) );
NOR2_X1 U842 ( .A1(n1170), .A2(n1120), .ZN(n1169) );
NAND2_X1 U843 ( .A1(G902), .A2(n1171), .ZN(n1120) );
NAND3_X1 U844 ( .A1(n1054), .A2(n1056), .A3(n1026), .ZN(n1171) );
AND4_X1 U845 ( .A1(n1134), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1026) );
AND3_X1 U846 ( .A1(n1175), .A2(n1020), .A3(n1176), .ZN(n1174) );
NAND3_X1 U847 ( .A1(n1177), .A2(n1039), .A3(n1178), .ZN(n1020) );
NAND2_X1 U848 ( .A1(n1052), .A2(n1179), .ZN(n1173) );
NAND2_X1 U849 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND4_X1 U850 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1180) );
XNOR2_X1 U851 ( .A(n1036), .B(KEYINPUT26), .ZN(n1182) );
NAND3_X1 U852 ( .A1(n1178), .A2(n1039), .A3(n1183), .ZN(n1134) );
AND3_X1 U853 ( .A1(n1186), .A2(n1098), .A3(n1096), .ZN(n1054) );
AND3_X1 U854 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1096) );
NAND2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1098) );
XOR2_X1 U856 ( .A(KEYINPUT22), .B(n1097), .Z(n1186) );
AND4_X1 U857 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1097) );
NAND3_X1 U858 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1192) );
OR2_X1 U859 ( .A1(n1190), .A2(KEYINPUT35), .ZN(n1197) );
NAND2_X1 U860 ( .A1(KEYINPUT35), .A2(n1199), .ZN(n1196) );
NAND2_X1 U861 ( .A1(n1200), .A2(n1047), .ZN(n1199) );
NAND2_X1 U862 ( .A1(n1201), .A2(KEYINPUT13), .ZN(n1168) );
XOR2_X1 U863 ( .A(n1141), .B(KEYINPUT31), .Z(n1201) );
NOR2_X1 U864 ( .A1(n1058), .A2(G952), .ZN(n1114) );
XNOR2_X1 U865 ( .A(G146), .B(n1193), .ZN(G48) );
NAND2_X1 U866 ( .A1(n1202), .A2(n1183), .ZN(n1193) );
NAND2_X1 U867 ( .A1(n1203), .A2(n1204), .ZN(G45) );
NAND2_X1 U868 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U869 ( .A(KEYINPUT42), .B(G143), .Z(n1206) );
XOR2_X1 U870 ( .A(n1194), .B(KEYINPUT24), .Z(n1205) );
XOR2_X1 U871 ( .A(KEYINPUT63), .B(n1207), .Z(n1203) );
NOR2_X1 U872 ( .A1(G143), .A2(n1194), .ZN(n1207) );
NAND3_X1 U873 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1194) );
NOR3_X1 U874 ( .A1(n1037), .A2(n1047), .A3(n1063), .ZN(n1210) );
XNOR2_X1 U875 ( .A(G140), .B(n1195), .ZN(G42) );
NAND3_X1 U876 ( .A1(n1183), .A2(n1211), .A3(n1190), .ZN(n1195) );
XOR2_X1 U877 ( .A(n1212), .B(n1213), .Z(G39) );
NOR2_X1 U878 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U879 ( .A1(KEYINPUT44), .A2(n1216), .ZN(n1212) );
XNOR2_X1 U880 ( .A(G134), .B(n1217), .ZN(G36) );
NAND4_X1 U881 ( .A1(n1031), .A2(n1191), .A3(n1218), .A4(n1219), .ZN(n1217) );
XNOR2_X1 U882 ( .A(KEYINPUT57), .B(n1220), .ZN(n1219) );
XNOR2_X1 U883 ( .A(G131), .B(n1189), .ZN(G33) );
NAND3_X1 U884 ( .A1(n1183), .A2(n1184), .A3(n1190), .ZN(n1189) );
INV_X1 U885 ( .A(n1215), .ZN(n1190) );
NAND2_X1 U886 ( .A1(n1200), .A2(n1218), .ZN(n1215) );
AND2_X1 U887 ( .A1(n1031), .A2(n1220), .ZN(n1200) );
AND2_X1 U888 ( .A1(n1059), .A2(n1221), .ZN(n1031) );
XNOR2_X1 U889 ( .A(G128), .B(n1187), .ZN(G30) );
NAND2_X1 U890 ( .A1(n1202), .A2(n1177), .ZN(n1187) );
AND4_X1 U891 ( .A1(n1209), .A2(n1218), .A3(n1067), .A4(n1222), .ZN(n1202) );
XNOR2_X1 U892 ( .A(G101), .B(n1056), .ZN(G3) );
NAND3_X1 U893 ( .A1(n1178), .A2(n1034), .A3(n1184), .ZN(n1056) );
XNOR2_X1 U894 ( .A(G125), .B(n1188), .ZN(G27) );
NAND4_X1 U895 ( .A1(n1209), .A2(n1183), .A3(n1036), .A4(n1211), .ZN(n1188) );
AND2_X1 U896 ( .A1(n1052), .A2(n1220), .ZN(n1209) );
NAND2_X1 U897 ( .A1(n1061), .A2(n1223), .ZN(n1220) );
NAND4_X1 U898 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1225), .ZN(n1223) );
INV_X1 U899 ( .A(G900), .ZN(n1225) );
XOR2_X1 U900 ( .A(G122), .B(n1226), .Z(G24) );
NOR2_X1 U901 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XOR2_X1 U902 ( .A(n1181), .B(KEYINPUT47), .Z(n1227) );
NAND3_X1 U903 ( .A1(n1208), .A2(n1036), .A3(n1229), .ZN(n1181) );
NOR3_X1 U904 ( .A1(n1230), .A2(n1231), .A3(n1063), .ZN(n1229) );
INV_X1 U905 ( .A(n1039), .ZN(n1230) );
NOR2_X1 U906 ( .A1(n1222), .A2(n1067), .ZN(n1039) );
INV_X1 U907 ( .A(n1232), .ZN(n1036) );
XNOR2_X1 U908 ( .A(G119), .B(n1172), .ZN(G21) );
NAND2_X1 U909 ( .A1(n1198), .A2(n1233), .ZN(n1172) );
INV_X1 U910 ( .A(n1214), .ZN(n1198) );
NAND3_X1 U911 ( .A1(n1067), .A2(n1222), .A3(n1034), .ZN(n1214) );
INV_X1 U912 ( .A(n1234), .ZN(n1222) );
XOR2_X1 U913 ( .A(n1175), .B(n1235), .Z(G18) );
NAND2_X1 U914 ( .A1(KEYINPUT60), .A2(G116), .ZN(n1235) );
NAND2_X1 U915 ( .A1(n1191), .A2(n1233), .ZN(n1175) );
NOR2_X1 U916 ( .A1(n1037), .A2(n1044), .ZN(n1191) );
INV_X1 U917 ( .A(n1184), .ZN(n1037) );
XOR2_X1 U918 ( .A(n1236), .B(n1237), .Z(G15) );
NOR2_X1 U919 ( .A1(KEYINPUT7), .A2(n1238), .ZN(n1237) );
AND3_X1 U920 ( .A1(n1183), .A2(n1184), .A3(n1233), .ZN(n1236) );
NOR3_X1 U921 ( .A1(n1228), .A2(n1231), .A3(n1232), .ZN(n1233) );
NAND2_X1 U922 ( .A1(n1050), .A2(n1064), .ZN(n1232) );
XNOR2_X1 U923 ( .A(n1069), .B(KEYINPUT4), .ZN(n1050) );
NOR2_X1 U924 ( .A1(n1067), .A2(n1234), .ZN(n1184) );
INV_X1 U925 ( .A(n1045), .ZN(n1183) );
NAND2_X1 U926 ( .A1(n1208), .A2(n1063), .ZN(n1045) );
XNOR2_X1 U927 ( .A(G110), .B(n1176), .ZN(G12) );
NAND3_X1 U928 ( .A1(n1178), .A2(n1034), .A3(n1211), .ZN(n1176) );
INV_X1 U929 ( .A(n1038), .ZN(n1211) );
NAND2_X1 U930 ( .A1(n1234), .A2(n1067), .ZN(n1038) );
XOR2_X1 U931 ( .A(n1239), .B(n1119), .Z(n1067) );
NAND2_X1 U932 ( .A1(G217), .A2(n1240), .ZN(n1119) );
NAND2_X1 U933 ( .A1(n1116), .A2(n1241), .ZN(n1239) );
XNOR2_X1 U934 ( .A(n1242), .B(n1243), .ZN(n1116) );
XOR2_X1 U935 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND2_X1 U936 ( .A1(n1246), .A2(G221), .ZN(n1245) );
NAND2_X1 U937 ( .A1(KEYINPUT0), .A2(n1247), .ZN(n1244) );
XNOR2_X1 U938 ( .A(n1248), .B(n1249), .ZN(n1247) );
XOR2_X1 U939 ( .A(G128), .B(G119), .Z(n1249) );
XOR2_X1 U940 ( .A(n1250), .B(n1251), .Z(n1242) );
NAND2_X1 U941 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
NAND2_X1 U942 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XNOR2_X1 U943 ( .A(n1256), .B(n1087), .ZN(n1255) );
XNOR2_X1 U944 ( .A(G146), .B(KEYINPUT14), .ZN(n1254) );
XOR2_X1 U945 ( .A(n1257), .B(KEYINPUT61), .Z(n1252) );
NAND2_X1 U946 ( .A1(n1258), .A2(G146), .ZN(n1257) );
XOR2_X1 U947 ( .A(n1256), .B(n1087), .Z(n1258) );
NAND2_X1 U948 ( .A1(KEYINPUT2), .A2(n1086), .ZN(n1256) );
NOR2_X1 U949 ( .A1(n1259), .A2(n1072), .ZN(n1234) );
NOR2_X1 U950 ( .A1(n1260), .A2(G472), .ZN(n1072) );
NOR2_X1 U951 ( .A1(n1077), .A2(n1075), .ZN(n1259) );
INV_X1 U952 ( .A(n1260), .ZN(n1075) );
NAND2_X1 U953 ( .A1(n1261), .A2(n1241), .ZN(n1260) );
XOR2_X1 U954 ( .A(n1137), .B(n1262), .Z(n1261) );
XOR2_X1 U955 ( .A(KEYINPUT30), .B(n1263), .Z(n1262) );
NOR2_X1 U956 ( .A1(KEYINPUT43), .A2(n1141), .ZN(n1263) );
XOR2_X1 U957 ( .A(n1264), .B(n1265), .Z(n1137) );
XOR2_X1 U958 ( .A(G101), .B(n1266), .Z(n1265) );
NOR3_X1 U959 ( .A1(n1170), .A2(G953), .A3(G237), .ZN(n1266) );
INV_X1 U960 ( .A(G210), .ZN(n1170) );
XNOR2_X1 U961 ( .A(n1267), .B(n1268), .ZN(n1264) );
XNOR2_X1 U962 ( .A(n1269), .B(n1089), .ZN(n1268) );
NOR2_X1 U963 ( .A1(KEYINPUT51), .A2(n1238), .ZN(n1269) );
INV_X1 U964 ( .A(G472), .ZN(n1077) );
NAND2_X1 U965 ( .A1(n1270), .A2(n1271), .ZN(n1034) );
OR2_X1 U966 ( .A1(n1044), .A2(KEYINPUT16), .ZN(n1271) );
INV_X1 U967 ( .A(n1177), .ZN(n1044) );
NOR2_X1 U968 ( .A1(n1063), .A2(n1208), .ZN(n1177) );
INV_X1 U969 ( .A(n1272), .ZN(n1208) );
NAND3_X1 U970 ( .A1(n1272), .A2(n1063), .A3(KEYINPUT16), .ZN(n1270) );
XNOR2_X1 U971 ( .A(n1273), .B(n1274), .ZN(n1063) );
XOR2_X1 U972 ( .A(KEYINPUT46), .B(G478), .Z(n1274) );
NAND2_X1 U973 ( .A1(n1123), .A2(n1241), .ZN(n1273) );
XNOR2_X1 U974 ( .A(n1275), .B(n1276), .ZN(n1123) );
XOR2_X1 U975 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U976 ( .A(G122), .B(G116), .Z(n1278) );
XOR2_X1 U977 ( .A(KEYINPUT21), .B(G134), .Z(n1277) );
XOR2_X1 U978 ( .A(n1279), .B(n1280), .Z(n1275) );
XOR2_X1 U979 ( .A(n1281), .B(G107), .Z(n1279) );
NAND2_X1 U980 ( .A1(G217), .A2(n1246), .ZN(n1281) );
AND2_X1 U981 ( .A1(G234), .A2(n1058), .ZN(n1246) );
XOR2_X1 U982 ( .A(n1068), .B(KEYINPUT56), .Z(n1272) );
XNOR2_X1 U983 ( .A(n1282), .B(G475), .ZN(n1068) );
NAND2_X1 U984 ( .A1(n1241), .A2(n1132), .ZN(n1282) );
NAND2_X1 U985 ( .A1(n1283), .A2(n1284), .ZN(n1132) );
NAND2_X1 U986 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XOR2_X1 U987 ( .A(n1287), .B(KEYINPUT8), .Z(n1283) );
OR2_X1 U988 ( .A1(n1286), .A2(n1285), .ZN(n1287) );
XNOR2_X1 U989 ( .A(n1288), .B(n1289), .ZN(n1285) );
XNOR2_X1 U990 ( .A(G131), .B(n1290), .ZN(n1289) );
NAND2_X1 U991 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND2_X1 U992 ( .A1(n1293), .A2(n1086), .ZN(n1292) );
XNOR2_X1 U993 ( .A(n1294), .B(KEYINPUT59), .ZN(n1293) );
NAND2_X1 U994 ( .A1(n1295), .A2(G140), .ZN(n1291) );
XNOR2_X1 U995 ( .A(KEYINPUT19), .B(n1296), .ZN(n1295) );
INV_X1 U996 ( .A(n1294), .ZN(n1296) );
XOR2_X1 U997 ( .A(n1087), .B(n1297), .Z(n1294) );
NOR4_X1 U998 ( .A1(KEYINPUT25), .A2(G237), .A3(n1298), .A4(n1299), .ZN(n1297) );
XNOR2_X1 U999 ( .A(KEYINPUT15), .B(n1058), .ZN(n1299) );
INV_X1 U1000 ( .A(G214), .ZN(n1298) );
XNOR2_X1 U1001 ( .A(G143), .B(G146), .ZN(n1288) );
XNOR2_X1 U1002 ( .A(G104), .B(n1300), .ZN(n1286) );
XNOR2_X1 U1003 ( .A(G122), .B(n1238), .ZN(n1300) );
INV_X1 U1004 ( .A(G113), .ZN(n1238) );
NOR3_X1 U1005 ( .A1(n1228), .A2(n1231), .A3(n1047), .ZN(n1178) );
INV_X1 U1006 ( .A(n1218), .ZN(n1047) );
NOR2_X1 U1007 ( .A1(n1301), .A2(n1049), .ZN(n1218) );
INV_X1 U1008 ( .A(n1064), .ZN(n1049) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1240), .ZN(n1064) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1241), .ZN(n1240) );
INV_X1 U1011 ( .A(n1069), .ZN(n1301) );
XNOR2_X1 U1012 ( .A(n1302), .B(G469), .ZN(n1069) );
NAND2_X1 U1013 ( .A1(n1303), .A2(n1241), .ZN(n1302) );
XOR2_X1 U1014 ( .A(n1304), .B(n1151), .Z(n1303) );
XNOR2_X1 U1015 ( .A(n1305), .B(n1306), .ZN(n1151) );
XNOR2_X1 U1016 ( .A(n1086), .B(G110), .ZN(n1306) );
INV_X1 U1017 ( .A(G140), .ZN(n1086) );
NAND2_X1 U1018 ( .A1(G227), .A2(n1058), .ZN(n1305) );
NAND2_X1 U1019 ( .A1(n1307), .A2(KEYINPUT29), .ZN(n1304) );
XOR2_X1 U1020 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1021 ( .A(n1164), .B(n1163), .ZN(n1309) );
XNOR2_X1 U1022 ( .A(n1310), .B(n1311), .ZN(n1163) );
NOR2_X1 U1023 ( .A1(KEYINPUT23), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1024 ( .A(G101), .B(KEYINPUT10), .ZN(n1310) );
XNOR2_X1 U1025 ( .A(n1088), .B(KEYINPUT36), .ZN(n1164) );
NAND2_X1 U1026 ( .A1(n1313), .A2(n1314), .ZN(n1088) );
NAND2_X1 U1027 ( .A1(n1280), .A2(n1315), .ZN(n1314) );
INV_X1 U1028 ( .A(G146), .ZN(n1315) );
NAND2_X1 U1029 ( .A1(n1316), .A2(G146), .ZN(n1313) );
XOR2_X1 U1030 ( .A(KEYINPUT9), .B(n1280), .Z(n1316) );
XNOR2_X1 U1031 ( .A(n1317), .B(n1089), .ZN(n1308) );
INV_X1 U1032 ( .A(n1161), .ZN(n1089) );
XNOR2_X1 U1033 ( .A(n1318), .B(n1251), .ZN(n1161) );
XNOR2_X1 U1034 ( .A(n1216), .B(KEYINPUT55), .ZN(n1251) );
INV_X1 U1035 ( .A(G137), .ZN(n1216) );
XNOR2_X1 U1036 ( .A(G131), .B(G134), .ZN(n1318) );
XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(KEYINPUT1), .ZN(n1317) );
INV_X1 U1038 ( .A(n1185), .ZN(n1231) );
NAND2_X1 U1039 ( .A1(n1061), .A2(n1319), .ZN(n1185) );
NAND4_X1 U1040 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1320), .ZN(n1319) );
INV_X1 U1041 ( .A(G898), .ZN(n1320) );
NAND3_X1 U1042 ( .A1(n1224), .A2(n1058), .A3(G952), .ZN(n1061) );
NAND2_X1 U1043 ( .A1(G237), .A2(G234), .ZN(n1224) );
INV_X1 U1044 ( .A(n1052), .ZN(n1228) );
NOR2_X1 U1045 ( .A1(n1060), .A2(n1059), .ZN(n1052) );
NOR2_X1 U1046 ( .A1(n1321), .A2(n1079), .ZN(n1059) );
NOR2_X1 U1047 ( .A1(n1322), .A2(n1323), .ZN(n1079) );
AND2_X1 U1048 ( .A1(G210), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1049 ( .A(n1078), .B(KEYINPUT50), .Z(n1321) );
AND3_X1 U1050 ( .A1(n1322), .A2(n1324), .A3(G210), .ZN(n1078) );
NAND2_X1 U1051 ( .A1(n1325), .A2(n1241), .ZN(n1322) );
INV_X1 U1052 ( .A(G902), .ZN(n1241) );
XOR2_X1 U1053 ( .A(n1167), .B(n1141), .Z(n1325) );
XOR2_X1 U1054 ( .A(n1326), .B(n1280), .Z(n1141) );
XOR2_X1 U1055 ( .A(G128), .B(G143), .Z(n1280) );
XNOR2_X1 U1056 ( .A(G146), .B(KEYINPUT5), .ZN(n1326) );
XNOR2_X1 U1057 ( .A(n1327), .B(n1328), .ZN(n1167) );
XOR2_X1 U1058 ( .A(n1087), .B(n1109), .Z(n1328) );
XNOR2_X1 U1059 ( .A(n1329), .B(G122), .ZN(n1109) );
NAND2_X1 U1060 ( .A1(KEYINPUT45), .A2(n1248), .ZN(n1329) );
INV_X1 U1061 ( .A(G110), .ZN(n1248) );
XOR2_X1 U1062 ( .A(G125), .B(KEYINPUT11), .Z(n1087) );
XOR2_X1 U1063 ( .A(n1330), .B(n1331), .Z(n1327) );
AND2_X1 U1064 ( .A1(n1058), .A2(G224), .ZN(n1331) );
INV_X1 U1065 ( .A(G953), .ZN(n1058) );
NAND2_X1 U1066 ( .A1(n1332), .A2(n1333), .ZN(n1330) );
OR2_X1 U1067 ( .A1(n1108), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1068 ( .A(n1335), .B(KEYINPUT41), .Z(n1332) );
NAND2_X1 U1069 ( .A1(n1334), .A2(n1108), .ZN(n1335) );
XOR2_X1 U1070 ( .A(G113), .B(n1267), .Z(n1108) );
XOR2_X1 U1071 ( .A(G116), .B(G119), .Z(n1267) );
XNOR2_X1 U1072 ( .A(n1110), .B(KEYINPUT48), .ZN(n1334) );
XOR2_X1 U1073 ( .A(G101), .B(n1312), .Z(n1110) );
XNOR2_X1 U1074 ( .A(G104), .B(G107), .ZN(n1312) );
INV_X1 U1075 ( .A(n1221), .ZN(n1060) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1324), .ZN(n1221) );
OR2_X1 U1077 ( .A1(G902), .A2(G237), .ZN(n1324) );
endmodule


