//Key = 1111111100110000111000011110001000010110100001001100110110010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424, n1425, n1426, n1427, n1428;

XOR2_X1 U786 ( .A(n1094), .B(n1095), .Z(G9) );
XOR2_X1 U787 ( .A(KEYINPUT17), .B(G107), .Z(n1095) );
NAND4_X1 U788 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1094) );
AND2_X1 U789 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
XOR2_X1 U790 ( .A(n1102), .B(KEYINPUT18), .Z(n1096) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(G75) );
NOR4_X1 U792 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1104) );
NOR2_X1 U793 ( .A1(n1102), .A2(n1109), .ZN(n1107) );
INV_X1 U794 ( .A(n1110), .ZN(n1102) );
NAND4_X1 U795 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1105) );
NAND3_X1 U796 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1112) );
XNOR2_X1 U797 ( .A(KEYINPUT46), .B(n1109), .ZN(n1116) );
NAND4_X1 U798 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1101), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1111) );
NAND2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U801 ( .A1(KEYINPUT44), .A2(n1125), .ZN(n1124) );
NAND4_X1 U802 ( .A1(n1118), .A2(n1119), .A3(n1097), .A4(n1101), .ZN(n1125) );
NAND2_X1 U803 ( .A1(n1118), .A2(n1126), .ZN(n1123) );
NAND2_X1 U804 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND3_X1 U805 ( .A1(n1101), .A2(n1129), .A3(n1120), .ZN(n1128) );
OR2_X1 U806 ( .A1(n1130), .A2(n1099), .ZN(n1129) );
NAND2_X1 U807 ( .A1(n1119), .A2(n1131), .ZN(n1127) );
NAND2_X1 U808 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U809 ( .A1(n1101), .A2(n1134), .ZN(n1133) );
NAND2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
OR2_X1 U811 ( .A1(n1137), .A2(KEYINPUT44), .ZN(n1136) );
NAND2_X1 U812 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
NAND2_X1 U813 ( .A1(n1120), .A2(n1140), .ZN(n1132) );
OR2_X1 U814 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U815 ( .A(n1143), .ZN(n1118) );
NOR3_X1 U816 ( .A1(n1144), .A2(G953), .A3(G952), .ZN(n1103) );
INV_X1 U817 ( .A(n1113), .ZN(n1144) );
NAND4_X1 U818 ( .A1(n1145), .A2(n1121), .A3(n1146), .A4(n1147), .ZN(n1113) );
NOR4_X1 U819 ( .A1(n1138), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1147) );
XOR2_X1 U820 ( .A(n1151), .B(KEYINPUT4), .Z(n1149) );
NOR2_X1 U821 ( .A1(G478), .A2(n1152), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1153), .A2(n1154), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1155), .B(n1156), .Z(n1145) );
NAND2_X1 U824 ( .A1(KEYINPUT16), .A2(G475), .ZN(n1155) );
XOR2_X1 U825 ( .A(n1157), .B(n1158), .Z(G72) );
XOR2_X1 U826 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U827 ( .A1(n1161), .A2(n1114), .ZN(n1160) );
AND2_X1 U828 ( .A1(G227), .A2(G900), .ZN(n1161) );
NAND2_X1 U829 ( .A1(n1162), .A2(n1163), .ZN(n1159) );
NAND2_X1 U830 ( .A1(G953), .A2(n1164), .ZN(n1163) );
XOR2_X1 U831 ( .A(n1165), .B(n1166), .Z(n1162) );
XOR2_X1 U832 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U833 ( .A(n1169), .B(KEYINPUT15), .ZN(n1165) );
NAND2_X1 U834 ( .A1(KEYINPUT49), .A2(n1170), .ZN(n1169) );
XNOR2_X1 U835 ( .A(n1171), .B(n1172), .ZN(n1170) );
NAND2_X1 U836 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
OR2_X1 U837 ( .A1(n1175), .A2(G137), .ZN(n1174) );
XOR2_X1 U838 ( .A(n1176), .B(KEYINPUT54), .Z(n1173) );
NAND2_X1 U839 ( .A1(G137), .A2(n1175), .ZN(n1176) );
NAND2_X1 U840 ( .A1(n1114), .A2(n1108), .ZN(n1157) );
XOR2_X1 U841 ( .A(n1177), .B(n1178), .Z(G69) );
NAND2_X1 U842 ( .A1(G953), .A2(n1179), .ZN(n1178) );
NAND2_X1 U843 ( .A1(n1180), .A2(G898), .ZN(n1179) );
XNOR2_X1 U844 ( .A(G224), .B(KEYINPUT23), .ZN(n1180) );
NAND2_X1 U845 ( .A1(KEYINPUT0), .A2(n1181), .ZN(n1177) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1181) );
AND2_X1 U847 ( .A1(n1106), .A2(n1114), .ZN(n1183) );
NOR3_X1 U848 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1182) );
INV_X1 U849 ( .A(n1187), .ZN(n1185) );
XOR2_X1 U850 ( .A(n1188), .B(KEYINPUT53), .Z(n1184) );
NOR2_X1 U851 ( .A1(n1189), .A2(n1190), .ZN(G66) );
NOR2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U853 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U854 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U855 ( .A1(KEYINPUT56), .A2(n1197), .ZN(n1193) );
NOR2_X1 U856 ( .A1(KEYINPUT56), .A2(n1197), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1189), .A2(n1198), .ZN(G63) );
XNOR2_X1 U858 ( .A(n1199), .B(n1200), .ZN(n1198) );
NOR2_X1 U859 ( .A1(n1201), .A2(n1196), .ZN(n1200) );
INV_X1 U860 ( .A(G478), .ZN(n1201) );
NOR2_X1 U861 ( .A1(n1189), .A2(n1202), .ZN(G60) );
XOR2_X1 U862 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U863 ( .A1(n1205), .A2(n1196), .ZN(n1204) );
INV_X1 U864 ( .A(G475), .ZN(n1205) );
NAND2_X1 U865 ( .A1(n1206), .A2(n1207), .ZN(G6) );
NAND2_X1 U866 ( .A1(G104), .A2(n1208), .ZN(n1207) );
XOR2_X1 U867 ( .A(n1209), .B(KEYINPUT33), .Z(n1206) );
OR2_X1 U868 ( .A1(n1208), .A2(G104), .ZN(n1209) );
NOR2_X1 U869 ( .A1(n1189), .A2(n1210), .ZN(G57) );
XOR2_X1 U870 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U871 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U872 ( .A(n1215), .B(n1216), .Z(n1211) );
NOR2_X1 U873 ( .A1(n1217), .A2(n1196), .ZN(n1216) );
INV_X1 U874 ( .A(G472), .ZN(n1217) );
NAND2_X1 U875 ( .A1(KEYINPUT62), .A2(n1218), .ZN(n1215) );
NOR3_X1 U876 ( .A1(n1189), .A2(n1219), .A3(n1220), .ZN(G54) );
NOR2_X1 U877 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XOR2_X1 U878 ( .A(n1223), .B(n1224), .Z(n1222) );
NAND2_X1 U879 ( .A1(KEYINPUT5), .A2(n1225), .ZN(n1223) );
NOR2_X1 U880 ( .A1(n1226), .A2(n1227), .ZN(n1219) );
XOR2_X1 U881 ( .A(n1228), .B(n1224), .Z(n1227) );
XNOR2_X1 U882 ( .A(n1229), .B(n1230), .ZN(n1224) );
NOR2_X1 U883 ( .A1(n1231), .A2(n1196), .ZN(n1230) );
INV_X1 U884 ( .A(G469), .ZN(n1231) );
NAND2_X1 U885 ( .A1(n1232), .A2(n1233), .ZN(n1229) );
NAND3_X1 U886 ( .A1(n1234), .A2(KEYINPUT11), .A3(n1235), .ZN(n1233) );
XOR2_X1 U887 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND2_X1 U888 ( .A1(n1168), .A2(n1238), .ZN(n1236) );
INV_X1 U889 ( .A(n1239), .ZN(n1168) );
NAND2_X1 U890 ( .A1(n1240), .A2(n1241), .ZN(n1232) );
NAND2_X1 U891 ( .A1(KEYINPUT11), .A2(n1234), .ZN(n1241) );
XOR2_X1 U892 ( .A(n1242), .B(n1237), .Z(n1240) );
NAND2_X1 U893 ( .A1(n1239), .A2(n1238), .ZN(n1242) );
INV_X1 U894 ( .A(KEYINPUT22), .ZN(n1238) );
NAND2_X1 U895 ( .A1(KEYINPUT5), .A2(n1243), .ZN(n1228) );
INV_X1 U896 ( .A(n1225), .ZN(n1243) );
INV_X1 U897 ( .A(n1221), .ZN(n1226) );
NOR2_X1 U898 ( .A1(n1189), .A2(n1244), .ZN(G51) );
XOR2_X1 U899 ( .A(n1245), .B(n1246), .Z(n1244) );
NOR2_X1 U900 ( .A1(n1247), .A2(n1196), .ZN(n1246) );
NAND2_X1 U901 ( .A1(G902), .A2(n1248), .ZN(n1196) );
OR2_X1 U902 ( .A1(n1106), .A2(n1108), .ZN(n1248) );
NAND2_X1 U903 ( .A1(n1249), .A2(n1250), .ZN(n1108) );
NOR4_X1 U904 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1250) );
INV_X1 U905 ( .A(n1255), .ZN(n1253) );
AND4_X1 U906 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1249) );
OR2_X1 U907 ( .A1(n1137), .A2(n1260), .ZN(n1259) );
NAND2_X1 U908 ( .A1(n1261), .A2(n1262), .ZN(n1106) );
NOR4_X1 U909 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1262) );
NOR4_X1 U910 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1261) );
AND3_X1 U911 ( .A1(n1271), .A2(n1101), .A3(n1099), .ZN(n1270) );
INV_X1 U912 ( .A(n1208), .ZN(n1269) );
NAND3_X1 U913 ( .A1(n1271), .A2(n1101), .A3(n1130), .ZN(n1208) );
INV_X1 U914 ( .A(n1272), .ZN(n1268) );
NAND2_X1 U915 ( .A1(n1273), .A2(KEYINPUT35), .ZN(n1245) );
XOR2_X1 U916 ( .A(n1274), .B(n1275), .Z(n1273) );
NOR2_X1 U917 ( .A1(KEYINPUT47), .A2(n1276), .ZN(n1275) );
XOR2_X1 U918 ( .A(n1277), .B(n1278), .Z(n1276) );
AND2_X1 U919 ( .A1(G953), .A2(n1279), .ZN(n1189) );
XOR2_X1 U920 ( .A(KEYINPUT1), .B(G952), .Z(n1279) );
XOR2_X1 U921 ( .A(n1257), .B(n1280), .Z(G48) );
NAND2_X1 U922 ( .A1(KEYINPUT38), .A2(G146), .ZN(n1280) );
NAND3_X1 U923 ( .A1(n1130), .A2(n1110), .A3(n1281), .ZN(n1257) );
NAND3_X1 U924 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(G45) );
NAND2_X1 U925 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U926 ( .A1(KEYINPUT34), .A2(n1287), .ZN(n1283) );
NAND2_X1 U927 ( .A1(n1288), .A2(G143), .ZN(n1287) );
XNOR2_X1 U928 ( .A(KEYINPUT39), .B(n1285), .ZN(n1288) );
NAND2_X1 U929 ( .A1(n1289), .A2(n1290), .ZN(n1282) );
INV_X1 U930 ( .A(KEYINPUT34), .ZN(n1290) );
NAND2_X1 U931 ( .A1(n1291), .A2(n1292), .ZN(n1289) );
OR3_X1 U932 ( .A1(n1286), .A2(n1285), .A3(KEYINPUT39), .ZN(n1292) );
NAND2_X1 U933 ( .A1(KEYINPUT39), .A2(n1285), .ZN(n1291) );
NOR2_X1 U934 ( .A1(n1260), .A2(n1293), .ZN(n1285) );
XOR2_X1 U935 ( .A(KEYINPUT31), .B(n1137), .Z(n1293) );
NAND3_X1 U936 ( .A1(n1141), .A2(n1110), .A3(n1294), .ZN(n1260) );
NOR3_X1 U937 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
XOR2_X1 U938 ( .A(n1298), .B(n1256), .Z(G42) );
NAND3_X1 U939 ( .A1(n1130), .A2(n1142), .A3(n1299), .ZN(n1256) );
XOR2_X1 U940 ( .A(G137), .B(n1254), .Z(G39) );
AND3_X1 U941 ( .A1(n1119), .A2(n1121), .A3(n1281), .ZN(n1254) );
XOR2_X1 U942 ( .A(n1175), .B(n1255), .Z(G36) );
NAND3_X1 U943 ( .A1(n1141), .A2(n1099), .A3(n1299), .ZN(n1255) );
XOR2_X1 U944 ( .A(G131), .B(n1252), .Z(G33) );
AND3_X1 U945 ( .A1(n1130), .A2(n1141), .A3(n1299), .ZN(n1252) );
AND3_X1 U946 ( .A1(n1097), .A2(n1300), .A3(n1121), .ZN(n1299) );
NOR2_X1 U947 ( .A1(n1301), .A2(n1117), .ZN(n1121) );
INV_X1 U948 ( .A(n1115), .ZN(n1301) );
NAND2_X1 U949 ( .A1(n1302), .A2(n1303), .ZN(G30) );
NAND2_X1 U950 ( .A1(G128), .A2(n1258), .ZN(n1303) );
XOR2_X1 U951 ( .A(KEYINPUT25), .B(n1304), .Z(n1302) );
NOR2_X1 U952 ( .A1(G128), .A2(n1258), .ZN(n1304) );
NAND3_X1 U953 ( .A1(n1099), .A2(n1110), .A3(n1281), .ZN(n1258) );
NOR4_X1 U954 ( .A1(n1137), .A2(n1305), .A3(n1306), .A4(n1297), .ZN(n1281) );
INV_X1 U955 ( .A(n1300), .ZN(n1297) );
INV_X1 U956 ( .A(n1097), .ZN(n1137) );
XOR2_X1 U957 ( .A(G101), .B(n1265), .Z(G3) );
AND3_X1 U958 ( .A1(n1119), .A2(n1141), .A3(n1271), .ZN(n1265) );
XOR2_X1 U959 ( .A(n1307), .B(n1308), .Z(G27) );
NAND2_X1 U960 ( .A1(KEYINPUT63), .A2(n1251), .ZN(n1308) );
AND4_X1 U961 ( .A1(n1110), .A2(n1300), .A3(n1120), .A4(n1309), .ZN(n1251) );
AND2_X1 U962 ( .A1(n1142), .A2(n1130), .ZN(n1309) );
NAND2_X1 U963 ( .A1(n1143), .A2(n1310), .ZN(n1300) );
NAND4_X1 U964 ( .A1(G902), .A2(G953), .A3(n1311), .A4(n1164), .ZN(n1310) );
INV_X1 U965 ( .A(G900), .ZN(n1164) );
XOR2_X1 U966 ( .A(n1312), .B(n1272), .Z(G24) );
NAND4_X1 U967 ( .A1(n1313), .A2(n1101), .A3(n1314), .A4(n1315), .ZN(n1272) );
AND2_X1 U968 ( .A1(n1306), .A2(n1316), .ZN(n1101) );
XOR2_X1 U969 ( .A(KEYINPUT61), .B(n1153), .Z(n1316) );
XOR2_X1 U970 ( .A(n1264), .B(n1317), .Z(G21) );
NOR2_X1 U971 ( .A1(KEYINPUT21), .A2(n1318), .ZN(n1317) );
AND4_X1 U972 ( .A1(n1119), .A2(n1313), .A3(n1153), .A4(n1154), .ZN(n1264) );
XOR2_X1 U973 ( .A(n1263), .B(n1319), .Z(G18) );
NOR2_X1 U974 ( .A1(KEYINPUT50), .A2(n1320), .ZN(n1319) );
AND3_X1 U975 ( .A1(n1313), .A2(n1099), .A3(n1141), .ZN(n1263) );
NOR2_X1 U976 ( .A1(n1314), .A2(n1296), .ZN(n1099) );
INV_X1 U977 ( .A(n1315), .ZN(n1296) );
XOR2_X1 U978 ( .A(G113), .B(n1267), .Z(G15) );
AND3_X1 U979 ( .A1(n1141), .A2(n1313), .A3(n1130), .ZN(n1267) );
NOR2_X1 U980 ( .A1(n1315), .A2(n1295), .ZN(n1130) );
INV_X1 U981 ( .A(n1314), .ZN(n1295) );
AND3_X1 U982 ( .A1(n1110), .A2(n1100), .A3(n1120), .ZN(n1313) );
AND2_X1 U983 ( .A1(n1139), .A2(n1321), .ZN(n1120) );
NOR2_X1 U984 ( .A1(n1153), .A2(n1306), .ZN(n1141) );
INV_X1 U985 ( .A(n1305), .ZN(n1153) );
XOR2_X1 U986 ( .A(n1322), .B(n1266), .Z(G12) );
AND3_X1 U987 ( .A1(n1271), .A2(n1119), .A3(n1142), .ZN(n1266) );
NOR2_X1 U988 ( .A1(n1154), .A2(n1305), .ZN(n1142) );
XNOR2_X1 U989 ( .A(n1323), .B(n1195), .ZN(n1305) );
NAND2_X1 U990 ( .A1(G217), .A2(n1324), .ZN(n1195) );
NAND2_X1 U991 ( .A1(G234), .A2(n1325), .ZN(n1324) );
OR2_X1 U992 ( .A1(n1197), .A2(G902), .ZN(n1323) );
XNOR2_X1 U993 ( .A(n1326), .B(n1327), .ZN(n1197) );
XNOR2_X1 U994 ( .A(G137), .B(n1328), .ZN(n1327) );
NAND2_X1 U995 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
OR2_X1 U996 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U997 ( .A(n1333), .B(KEYINPUT51), .Z(n1329) );
NAND2_X1 U998 ( .A1(n1332), .A2(n1331), .ZN(n1333) );
XNOR2_X1 U999 ( .A(n1334), .B(G110), .ZN(n1331) );
NAND2_X1 U1000 ( .A1(KEYINPUT2), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1001 ( .A(G119), .B(n1336), .Z(n1335) );
NOR2_X1 U1002 ( .A1(G128), .A2(KEYINPUT42), .ZN(n1336) );
XOR2_X1 U1003 ( .A(G146), .B(n1337), .Z(n1332) );
NOR2_X1 U1004 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NOR2_X1 U1005 ( .A1(KEYINPUT36), .A2(n1167), .ZN(n1339) );
NOR2_X1 U1006 ( .A1(KEYINPUT48), .A2(n1340), .ZN(n1338) );
INV_X1 U1007 ( .A(n1167), .ZN(n1340) );
XNOR2_X1 U1008 ( .A(n1307), .B(G140), .ZN(n1167) );
NAND3_X1 U1009 ( .A1(G234), .A2(n1114), .A3(G221), .ZN(n1326) );
INV_X1 U1010 ( .A(n1306), .ZN(n1154) );
XOR2_X1 U1011 ( .A(n1341), .B(G472), .Z(n1306) );
NAND2_X1 U1012 ( .A1(n1342), .A2(n1325), .ZN(n1341) );
XOR2_X1 U1013 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1014 ( .A(n1345), .B(KEYINPUT28), .ZN(n1344) );
NAND2_X1 U1015 ( .A1(KEYINPUT7), .A2(n1213), .ZN(n1345) );
XOR2_X1 U1016 ( .A(n1346), .B(n1347), .Z(n1213) );
XOR2_X1 U1017 ( .A(G119), .B(n1348), .Z(n1347) );
NOR2_X1 U1018 ( .A1(G116), .A2(KEYINPUT43), .ZN(n1348) );
INV_X1 U1019 ( .A(n1349), .ZN(n1346) );
XOR2_X1 U1020 ( .A(n1218), .B(n1214), .Z(n1343) );
XNOR2_X1 U1021 ( .A(n1350), .B(n1237), .ZN(n1214) );
XOR2_X1 U1022 ( .A(n1351), .B(G101), .Z(n1218) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1352), .ZN(n1351) );
NOR2_X1 U1024 ( .A1(n1315), .A2(n1314), .ZN(n1119) );
XOR2_X1 U1025 ( .A(n1156), .B(G475), .Z(n1314) );
NOR2_X1 U1026 ( .A1(n1203), .A2(G902), .ZN(n1156) );
XOR2_X1 U1027 ( .A(n1353), .B(n1354), .Z(n1203) );
XOR2_X1 U1028 ( .A(n1355), .B(n1356), .Z(n1354) );
NAND2_X1 U1029 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
OR2_X1 U1030 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
XOR2_X1 U1031 ( .A(n1361), .B(KEYINPUT60), .Z(n1357) );
NAND2_X1 U1032 ( .A1(n1360), .A2(n1359), .ZN(n1361) );
XNOR2_X1 U1033 ( .A(n1362), .B(n1363), .ZN(n1359) );
NOR2_X1 U1034 ( .A1(KEYINPUT41), .A2(n1307), .ZN(n1363) );
INV_X1 U1035 ( .A(G125), .ZN(n1307) );
XOR2_X1 U1036 ( .A(n1298), .B(G146), .Z(n1362) );
XNOR2_X1 U1037 ( .A(n1364), .B(n1365), .ZN(n1360) );
XOR2_X1 U1038 ( .A(G143), .B(G131), .Z(n1365) );
NAND2_X1 U1039 ( .A1(G214), .A2(n1352), .ZN(n1364) );
NOR2_X1 U1040 ( .A1(G953), .A2(G237), .ZN(n1352) );
NAND2_X1 U1041 ( .A1(n1366), .A2(KEYINPUT59), .ZN(n1355) );
XOR2_X1 U1042 ( .A(n1349), .B(KEYINPUT24), .Z(n1366) );
XOR2_X1 U1043 ( .A(n1312), .B(n1367), .Z(n1353) );
NOR2_X1 U1044 ( .A1(G104), .A2(KEYINPUT13), .ZN(n1367) );
NAND2_X1 U1045 ( .A1(n1368), .A2(n1151), .ZN(n1315) );
NAND2_X1 U1046 ( .A1(G478), .A2(n1152), .ZN(n1151) );
OR2_X1 U1047 ( .A1(n1152), .A2(G478), .ZN(n1368) );
NAND2_X1 U1048 ( .A1(n1199), .A2(n1325), .ZN(n1152) );
XNOR2_X1 U1049 ( .A(n1369), .B(n1370), .ZN(n1199) );
NOR2_X1 U1050 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
NOR2_X1 U1051 ( .A1(n1175), .A2(n1373), .ZN(n1372) );
XOR2_X1 U1052 ( .A(n1374), .B(KEYINPUT30), .Z(n1373) );
NOR2_X1 U1053 ( .A1(G134), .A2(n1375), .ZN(n1371) );
XOR2_X1 U1054 ( .A(n1374), .B(KEYINPUT19), .Z(n1375) );
XNOR2_X1 U1055 ( .A(G128), .B(n1376), .ZN(n1374) );
XOR2_X1 U1056 ( .A(KEYINPUT52), .B(G143), .Z(n1376) );
XOR2_X1 U1057 ( .A(n1377), .B(n1378), .Z(n1369) );
NOR2_X1 U1058 ( .A1(KEYINPUT9), .A2(n1379), .ZN(n1378) );
XOR2_X1 U1059 ( .A(n1380), .B(n1381), .Z(n1379) );
NAND2_X1 U1060 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
NAND2_X1 U1061 ( .A1(G122), .A2(n1320), .ZN(n1383) );
INV_X1 U1062 ( .A(G116), .ZN(n1320) );
XOR2_X1 U1063 ( .A(n1384), .B(KEYINPUT32), .Z(n1382) );
NAND2_X1 U1064 ( .A1(G116), .A2(n1312), .ZN(n1384) );
INV_X1 U1065 ( .A(G122), .ZN(n1312) );
INV_X1 U1066 ( .A(G107), .ZN(n1380) );
NAND3_X1 U1067 ( .A1(G234), .A2(n1114), .A3(G217), .ZN(n1377) );
AND3_X1 U1068 ( .A1(n1110), .A2(n1100), .A3(n1097), .ZN(n1271) );
NOR2_X1 U1069 ( .A1(n1139), .A2(n1138), .ZN(n1097) );
INV_X1 U1070 ( .A(n1321), .ZN(n1138) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1385), .ZN(n1321) );
XOR2_X1 U1072 ( .A(KEYINPUT37), .B(n1386), .Z(n1385) );
AND2_X1 U1073 ( .A1(n1325), .A2(G234), .ZN(n1386) );
XOR2_X1 U1074 ( .A(n1150), .B(KEYINPUT45), .Z(n1139) );
XNOR2_X1 U1075 ( .A(n1387), .B(G469), .ZN(n1150) );
NAND2_X1 U1076 ( .A1(n1388), .A2(n1325), .ZN(n1387) );
XOR2_X1 U1077 ( .A(n1389), .B(n1390), .Z(n1388) );
XNOR2_X1 U1078 ( .A(n1234), .B(n1391), .ZN(n1390) );
NOR2_X1 U1079 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
AND3_X1 U1080 ( .A1(KEYINPUT29), .A2(n1394), .A3(G140), .ZN(n1393) );
NOR2_X1 U1081 ( .A1(KEYINPUT29), .A2(n1225), .ZN(n1392) );
XNOR2_X1 U1082 ( .A(n1298), .B(G110), .ZN(n1225) );
INV_X1 U1083 ( .A(G140), .ZN(n1298) );
XOR2_X1 U1084 ( .A(n1395), .B(n1396), .Z(n1389) );
XOR2_X1 U1085 ( .A(n1221), .B(n1397), .Z(n1396) );
NOR2_X1 U1086 ( .A1(KEYINPUT12), .A2(n1239), .ZN(n1397) );
XOR2_X1 U1087 ( .A(n1286), .B(n1398), .Z(n1239) );
NAND2_X1 U1088 ( .A1(G227), .A2(n1114), .ZN(n1221) );
NAND2_X1 U1089 ( .A1(KEYINPUT3), .A2(n1237), .ZN(n1395) );
AND2_X1 U1090 ( .A1(n1399), .A2(n1400), .ZN(n1237) );
NAND2_X1 U1091 ( .A1(n1172), .A2(n1401), .ZN(n1400) );
XOR2_X1 U1092 ( .A(n1402), .B(KEYINPUT8), .Z(n1399) );
OR2_X1 U1093 ( .A1(n1401), .A2(n1172), .ZN(n1402) );
XOR2_X1 U1094 ( .A(G131), .B(KEYINPUT58), .Z(n1172) );
NAND3_X1 U1095 ( .A1(n1403), .A2(n1404), .A3(n1405), .ZN(n1401) );
NAND2_X1 U1096 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
NAND2_X1 U1097 ( .A1(n1408), .A2(KEYINPUT55), .ZN(n1407) );
XOR2_X1 U1098 ( .A(n1175), .B(KEYINPUT57), .Z(n1408) );
NAND3_X1 U1099 ( .A1(KEYINPUT55), .A2(n1409), .A3(n1175), .ZN(n1404) );
INV_X1 U1100 ( .A(n1406), .ZN(n1409) );
XNOR2_X1 U1101 ( .A(G137), .B(KEYINPUT27), .ZN(n1406) );
OR2_X1 U1102 ( .A1(n1175), .A2(KEYINPUT55), .ZN(n1403) );
INV_X1 U1103 ( .A(G134), .ZN(n1175) );
NAND2_X1 U1104 ( .A1(n1143), .A2(n1410), .ZN(n1100) );
NAND3_X1 U1105 ( .A1(n1186), .A2(n1311), .A3(G902), .ZN(n1410) );
NOR2_X1 U1106 ( .A1(n1114), .A2(G898), .ZN(n1186) );
NAND3_X1 U1107 ( .A1(n1311), .A2(n1114), .A3(G952), .ZN(n1143) );
NAND2_X1 U1108 ( .A1(G237), .A2(G234), .ZN(n1311) );
NOR2_X1 U1109 ( .A1(n1115), .A2(n1117), .ZN(n1110) );
AND2_X1 U1110 ( .A1(G214), .A2(n1411), .ZN(n1117) );
XNOR2_X1 U1111 ( .A(n1412), .B(n1247), .ZN(n1115) );
NAND2_X1 U1112 ( .A1(G210), .A2(n1411), .ZN(n1247) );
NAND2_X1 U1113 ( .A1(n1325), .A2(n1413), .ZN(n1411) );
INV_X1 U1114 ( .A(G237), .ZN(n1413) );
NAND2_X1 U1115 ( .A1(n1414), .A2(n1325), .ZN(n1412) );
INV_X1 U1116 ( .A(G902), .ZN(n1325) );
XOR2_X1 U1117 ( .A(n1415), .B(n1416), .Z(n1414) );
XOR2_X1 U1118 ( .A(n1277), .B(n1274), .Z(n1416) );
NAND2_X1 U1119 ( .A1(n1187), .A2(n1188), .ZN(n1274) );
NAND3_X1 U1120 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n1188) );
XOR2_X1 U1121 ( .A(n1394), .B(n1420), .Z(n1419) );
NAND2_X1 U1122 ( .A1(n1421), .A2(n1422), .ZN(n1187) );
NAND2_X1 U1123 ( .A1(n1417), .A2(n1418), .ZN(n1422) );
NAND2_X1 U1124 ( .A1(n1423), .A2(n1424), .ZN(n1418) );
XNOR2_X1 U1125 ( .A(KEYINPUT20), .B(n1425), .ZN(n1424) );
XOR2_X1 U1126 ( .A(G119), .B(G116), .Z(n1423) );
NAND2_X1 U1127 ( .A1(n1426), .A2(n1425), .ZN(n1417) );
XNOR2_X1 U1128 ( .A(n1234), .B(n1349), .ZN(n1425) );
XNOR2_X1 U1129 ( .A(G113), .B(KEYINPUT26), .ZN(n1349) );
XNOR2_X1 U1130 ( .A(G101), .B(n1427), .ZN(n1234) );
XOR2_X1 U1131 ( .A(G107), .B(G104), .Z(n1427) );
XOR2_X1 U1132 ( .A(n1318), .B(G116), .Z(n1426) );
INV_X1 U1133 ( .A(G119), .ZN(n1318) );
XOR2_X1 U1134 ( .A(G110), .B(n1420), .Z(n1421) );
NOR2_X1 U1135 ( .A1(KEYINPUT14), .A2(G122), .ZN(n1420) );
NAND2_X1 U1136 ( .A1(G224), .A2(n1114), .ZN(n1277) );
INV_X1 U1137 ( .A(G953), .ZN(n1114) );
NAND2_X1 U1138 ( .A1(KEYINPUT10), .A2(n1278), .ZN(n1415) );
XOR2_X1 U1139 ( .A(n1350), .B(G125), .Z(n1278) );
XOR2_X1 U1140 ( .A(n1428), .B(n1398), .Z(n1350) );
XOR2_X1 U1141 ( .A(G128), .B(G146), .Z(n1398) );
NAND2_X1 U1142 ( .A1(KEYINPUT6), .A2(n1286), .ZN(n1428) );
INV_X1 U1143 ( .A(G143), .ZN(n1286) );
NAND2_X1 U1144 ( .A1(KEYINPUT40), .A2(n1394), .ZN(n1322) );
INV_X1 U1145 ( .A(G110), .ZN(n1394) );
endmodule


