//Key = 1100001011011110011011100000110010011000001101101111000001111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286;

XNOR2_X1 U699 ( .A(G107), .B(n979), .ZN(G9) );
NAND4_X1 U700 ( .A1(KEYINPUT11), .A2(n980), .A3(n981), .A4(n982), .ZN(n979) );
NOR2_X1 U701 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR3_X1 U702 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
NOR2_X1 U703 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR2_X1 U704 ( .A1(n990), .A2(n991), .ZN(n988) );
XOR2_X1 U705 ( .A(KEYINPUT33), .B(n992), .Z(n991) );
NOR3_X1 U706 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NOR3_X1 U707 ( .A1(n994), .A2(n996), .A3(n997), .ZN(n990) );
NAND3_X1 U708 ( .A1(n982), .A2(n998), .A3(n999), .ZN(n994) );
NAND3_X1 U709 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n985) );
NAND3_X1 U710 ( .A1(n1003), .A2(n1004), .A3(n999), .ZN(n1002) );
INV_X1 U711 ( .A(n1005), .ZN(n999) );
NAND2_X1 U712 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NAND3_X1 U713 ( .A1(n982), .A2(n1008), .A3(n1009), .ZN(n1007) );
NAND2_X1 U714 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NAND2_X1 U715 ( .A1(n998), .A2(n1012), .ZN(n1006) );
NAND2_X1 U716 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U717 ( .A1(n1009), .A2(n1015), .ZN(n1014) );
NAND2_X1 U718 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U719 ( .A1(n982), .A2(n1018), .ZN(n1013) );
NAND2_X1 U720 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U721 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
AND3_X1 U722 ( .A1(n1000), .A2(n1001), .A3(n1023), .ZN(n983) );
NAND4_X1 U723 ( .A1(n1024), .A2(n1003), .A3(n1025), .A4(n1026), .ZN(n1000) );
NOR4_X1 U724 ( .A1(n1021), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1026) );
XNOR2_X1 U725 ( .A(n1030), .B(KEYINPUT63), .ZN(n1028) );
XNOR2_X1 U726 ( .A(n1031), .B(n1032), .ZN(n1027) );
NOR2_X1 U727 ( .A1(n1033), .A2(KEYINPUT15), .ZN(n1032) );
XNOR2_X1 U728 ( .A(n1034), .B(KEYINPUT25), .ZN(n1025) );
XNOR2_X1 U729 ( .A(n1035), .B(n1036), .ZN(n1024) );
XOR2_X1 U730 ( .A(n1037), .B(n1038), .Z(G72) );
XOR2_X1 U731 ( .A(n1039), .B(n1040), .Z(n1038) );
NOR2_X1 U732 ( .A1(n1041), .A2(n1001), .ZN(n1040) );
AND2_X1 U733 ( .A1(G227), .A2(G900), .ZN(n1041) );
NAND2_X1 U734 ( .A1(n1042), .A2(n1043), .ZN(n1039) );
NAND2_X1 U735 ( .A1(G953), .A2(n1044), .ZN(n1043) );
XOR2_X1 U736 ( .A(n1045), .B(n1046), .Z(n1042) );
XNOR2_X1 U737 ( .A(n1047), .B(n1048), .ZN(n1046) );
XNOR2_X1 U738 ( .A(n1049), .B(n1050), .ZN(n1045) );
NAND2_X1 U739 ( .A1(n1051), .A2(KEYINPUT57), .ZN(n1049) );
XNOR2_X1 U740 ( .A(G140), .B(KEYINPUT43), .ZN(n1051) );
NAND2_X1 U741 ( .A1(n1001), .A2(n1052), .ZN(n1037) );
NAND2_X1 U742 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
XOR2_X1 U743 ( .A(n1055), .B(n1056), .Z(G69) );
NAND2_X1 U744 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U745 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U746 ( .A(n1061), .ZN(n1060) );
NAND3_X1 U747 ( .A1(n1062), .A2(n1063), .A3(n1061), .ZN(n1057) );
XNOR2_X1 U748 ( .A(n1064), .B(n1065), .ZN(n1061) );
XOR2_X1 U749 ( .A(KEYINPUT48), .B(KEYINPUT35), .Z(n1065) );
XNOR2_X1 U750 ( .A(n1059), .B(KEYINPUT4), .ZN(n1062) );
NOR2_X1 U751 ( .A1(n1066), .A2(G953), .ZN(n1059) );
NAND2_X1 U752 ( .A1(n1063), .A2(n1067), .ZN(n1055) );
NAND2_X1 U753 ( .A1(G953), .A2(n1068), .ZN(n1067) );
INV_X1 U754 ( .A(n1069), .ZN(n1063) );
NOR2_X1 U755 ( .A1(n1070), .A2(n1071), .ZN(G66) );
NOR3_X1 U756 ( .A1(n1072), .A2(n1036), .A3(n1073), .ZN(n1071) );
NOR2_X1 U757 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U758 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
XOR2_X1 U759 ( .A(n1078), .B(KEYINPUT45), .Z(n1072) );
NAND3_X1 U760 ( .A1(n1035), .A2(n1075), .A3(n1079), .ZN(n1078) );
NOR2_X1 U761 ( .A1(n1070), .A2(n1080), .ZN(G63) );
XOR2_X1 U762 ( .A(n1081), .B(n1082), .Z(n1080) );
XOR2_X1 U763 ( .A(n1083), .B(KEYINPUT52), .Z(n1081) );
NAND2_X1 U764 ( .A1(n1079), .A2(G478), .ZN(n1083) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1084), .ZN(G60) );
XNOR2_X1 U766 ( .A(n1085), .B(n1086), .ZN(n1084) );
NAND2_X1 U767 ( .A1(KEYINPUT36), .A2(n1087), .ZN(n1085) );
NAND2_X1 U768 ( .A1(n1079), .A2(G475), .ZN(n1087) );
XNOR2_X1 U769 ( .A(G104), .B(n1088), .ZN(G6) );
NOR2_X1 U770 ( .A1(n1089), .A2(n1090), .ZN(G57) );
XOR2_X1 U771 ( .A(KEYINPUT30), .B(n1070), .Z(n1090) );
NOR2_X1 U772 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
XOR2_X1 U773 ( .A(KEYINPUT53), .B(n1093), .Z(n1092) );
NOR2_X1 U774 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
AND2_X1 U775 ( .A1(n1095), .A2(n1094), .ZN(n1091) );
AND2_X1 U776 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND2_X1 U777 ( .A1(G101), .A2(n1098), .ZN(n1097) );
XNOR2_X1 U778 ( .A(KEYINPUT39), .B(n1099), .ZN(n1098) );
XOR2_X1 U779 ( .A(KEYINPUT21), .B(n1100), .Z(n1096) );
NOR2_X1 U780 ( .A1(n1101), .A2(G101), .ZN(n1100) );
XNOR2_X1 U781 ( .A(n1102), .B(n1103), .ZN(n1095) );
NOR2_X1 U782 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
AND2_X1 U783 ( .A1(KEYINPUT49), .A2(n1106), .ZN(n1105) );
NOR3_X1 U784 ( .A1(KEYINPUT49), .A2(n1107), .A3(n1048), .ZN(n1104) );
XOR2_X1 U785 ( .A(n1108), .B(n1109), .Z(n1102) );
NOR2_X1 U786 ( .A1(KEYINPUT40), .A2(n1110), .ZN(n1109) );
NAND2_X1 U787 ( .A1(n1079), .A2(G472), .ZN(n1108) );
NOR2_X1 U788 ( .A1(n1070), .A2(n1111), .ZN(G54) );
XOR2_X1 U789 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U790 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U791 ( .A(G110), .B(G140), .ZN(n1115) );
XOR2_X1 U792 ( .A(n1116), .B(n1117), .Z(n1112) );
XOR2_X1 U793 ( .A(n1118), .B(n1119), .Z(n1116) );
NOR2_X1 U794 ( .A1(KEYINPUT23), .A2(n1120), .ZN(n1119) );
NAND2_X1 U795 ( .A1(n1079), .A2(G469), .ZN(n1118) );
NOR2_X1 U796 ( .A1(n1070), .A2(n1121), .ZN(G51) );
XOR2_X1 U797 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U798 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U799 ( .A1(KEYINPUT51), .A2(n1107), .ZN(n1124) );
XNOR2_X1 U800 ( .A(n1126), .B(n1050), .ZN(n1122) );
NAND2_X1 U801 ( .A1(n1079), .A2(n1031), .ZN(n1126) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1076), .ZN(n1079) );
INV_X1 U803 ( .A(n987), .ZN(n1076) );
NAND3_X1 U804 ( .A1(n1066), .A2(n1128), .A3(n1053), .ZN(n987) );
AND4_X1 U805 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1053) );
AND4_X1 U806 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1132) );
OR2_X1 U807 ( .A1(n1137), .A2(n1016), .ZN(n1129) );
XNOR2_X1 U808 ( .A(KEYINPUT59), .B(n1054), .ZN(n1128) );
AND4_X1 U809 ( .A1(n1088), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1066) );
AND4_X1 U810 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
NOR2_X1 U812 ( .A1(n1147), .A2(n1019), .ZN(n1146) );
XOR2_X1 U813 ( .A(n1148), .B(KEYINPUT31), .Z(n1147) );
NOR3_X1 U814 ( .A1(n1149), .A2(n1150), .A3(n1010), .ZN(n1145) );
NAND3_X1 U815 ( .A1(n980), .A2(n982), .A3(n1151), .ZN(n1088) );
AND2_X1 U816 ( .A1(n1152), .A2(n1023), .ZN(n1070) );
INV_X1 U817 ( .A(G952), .ZN(n1023) );
XNOR2_X1 U818 ( .A(G953), .B(KEYINPUT50), .ZN(n1152) );
XNOR2_X1 U819 ( .A(n1153), .B(n1130), .ZN(G48) );
NAND2_X1 U820 ( .A1(n1154), .A2(n1155), .ZN(n1130) );
NAND2_X1 U821 ( .A1(KEYINPUT13), .A2(n1156), .ZN(n1153) );
XOR2_X1 U822 ( .A(G143), .B(n1157), .Z(G45) );
NOR2_X1 U823 ( .A1(n1137), .A2(n1158), .ZN(n1157) );
XNOR2_X1 U824 ( .A(KEYINPUT32), .B(n1016), .ZN(n1158) );
NAND4_X1 U825 ( .A1(n1159), .A2(n1160), .A3(n1030), .A4(n1034), .ZN(n1137) );
XOR2_X1 U826 ( .A(n1161), .B(G140), .Z(G42) );
NAND2_X1 U827 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
OR2_X1 U828 ( .A1(n1131), .A2(KEYINPUT19), .ZN(n1163) );
NAND3_X1 U829 ( .A1(n1154), .A2(n1164), .A3(n1009), .ZN(n1131) );
NAND4_X1 U830 ( .A1(n1164), .A2(n989), .A3(n1154), .A4(KEYINPUT19), .ZN(n1162) );
XNOR2_X1 U831 ( .A(G137), .B(n1136), .ZN(G39) );
NAND4_X1 U832 ( .A1(n1165), .A2(n1029), .A3(n998), .A4(n1166), .ZN(n1136) );
NOR2_X1 U833 ( .A1(n1167), .A2(n989), .ZN(n1166) );
XOR2_X1 U834 ( .A(n1168), .B(G134), .Z(G36) );
NAND2_X1 U835 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
OR2_X1 U836 ( .A1(n1054), .A2(KEYINPUT27), .ZN(n1170) );
OR2_X1 U837 ( .A1(n1171), .A2(n989), .ZN(n1054) );
NAND3_X1 U838 ( .A1(n1009), .A2(n1171), .A3(KEYINPUT27), .ZN(n1169) );
NAND3_X1 U839 ( .A1(n1159), .A2(n981), .A3(n1172), .ZN(n1171) );
XNOR2_X1 U840 ( .A(G131), .B(n1135), .ZN(G33) );
NAND3_X1 U841 ( .A1(n1009), .A2(n1154), .A3(n1172), .ZN(n1135) );
NOR2_X1 U842 ( .A1(n1167), .A2(n1011), .ZN(n1154) );
INV_X1 U843 ( .A(n1159), .ZN(n1167) );
INV_X1 U844 ( .A(n989), .ZN(n1009) );
NAND2_X1 U845 ( .A1(n1022), .A2(n1173), .ZN(n989) );
XOR2_X1 U846 ( .A(n1174), .B(G128), .Z(G30) );
NAND2_X1 U847 ( .A1(KEYINPUT61), .A2(n1134), .ZN(n1174) );
NAND3_X1 U848 ( .A1(n1155), .A2(n981), .A3(n1159), .ZN(n1134) );
NOR3_X1 U849 ( .A1(n1175), .A2(n996), .A3(n997), .ZN(n1159) );
INV_X1 U850 ( .A(n995), .ZN(n997) );
XNOR2_X1 U851 ( .A(G101), .B(n1138), .ZN(G3) );
NAND3_X1 U852 ( .A1(n980), .A2(n998), .A3(n1172), .ZN(n1138) );
XNOR2_X1 U853 ( .A(G125), .B(n1133), .ZN(G27) );
NAND4_X1 U854 ( .A1(n1151), .A2(n1164), .A3(n1176), .A4(n1003), .ZN(n1133) );
NOR2_X1 U855 ( .A1(n1175), .A2(n1019), .ZN(n1176) );
AND2_X1 U856 ( .A1(n1005), .A2(n1177), .ZN(n1175) );
NAND4_X1 U857 ( .A1(G902), .A2(G953), .A3(n1178), .A4(n1044), .ZN(n1177) );
INV_X1 U858 ( .A(G900), .ZN(n1044) );
XNOR2_X1 U859 ( .A(n1179), .B(n1180), .ZN(G24) );
NOR2_X1 U860 ( .A1(n1019), .A2(n1148), .ZN(n1180) );
NAND4_X1 U861 ( .A1(n1181), .A2(n982), .A3(n1030), .A4(n1034), .ZN(n1148) );
INV_X1 U862 ( .A(n1150), .ZN(n982) );
NAND2_X1 U863 ( .A1(n1182), .A2(n1183), .ZN(n1150) );
XNOR2_X1 U864 ( .A(G119), .B(n1144), .ZN(G21) );
NAND3_X1 U865 ( .A1(n1155), .A2(n998), .A3(n1181), .ZN(n1144) );
AND3_X1 U866 ( .A1(n1165), .A2(n1029), .A3(n1160), .ZN(n1155) );
XNOR2_X1 U867 ( .A(G116), .B(n1143), .ZN(G18) );
NAND4_X1 U868 ( .A1(n1181), .A2(n1172), .A3(n981), .A4(n1160), .ZN(n1143) );
AND2_X1 U869 ( .A1(n1003), .A2(n1184), .ZN(n1181) );
XNOR2_X1 U870 ( .A(G113), .B(n1142), .ZN(G15) );
NAND4_X1 U871 ( .A1(n1172), .A2(n1151), .A3(n1003), .A4(n1185), .ZN(n1142) );
NOR2_X1 U872 ( .A1(n995), .A2(n996), .ZN(n1003) );
INV_X1 U873 ( .A(n993), .ZN(n996) );
INV_X1 U874 ( .A(n1011), .ZN(n1151) );
NAND2_X1 U875 ( .A1(n1186), .A2(n1187), .ZN(n1011) );
XNOR2_X1 U876 ( .A(KEYINPUT46), .B(n1188), .ZN(n1187) );
XNOR2_X1 U877 ( .A(n1030), .B(KEYINPUT14), .ZN(n1186) );
INV_X1 U878 ( .A(n1016), .ZN(n1172) );
NAND2_X1 U879 ( .A1(n1029), .A2(n1183), .ZN(n1016) );
XNOR2_X1 U880 ( .A(n1189), .B(n1141), .ZN(G12) );
NAND3_X1 U881 ( .A1(n980), .A2(n998), .A3(n1164), .ZN(n1141) );
INV_X1 U882 ( .A(n1017), .ZN(n1164) );
NAND2_X1 U883 ( .A1(n1182), .A2(n1165), .ZN(n1017) );
XNOR2_X1 U884 ( .A(n1183), .B(KEYINPUT5), .ZN(n1165) );
NAND3_X1 U885 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1183) );
NAND2_X1 U886 ( .A1(n1036), .A2(n1193), .ZN(n1192) );
OR3_X1 U887 ( .A1(n1193), .A2(n1036), .A3(KEYINPUT55), .ZN(n1191) );
NOR2_X1 U888 ( .A1(n1075), .A2(G902), .ZN(n1036) );
XNOR2_X1 U889 ( .A(n1194), .B(n1195), .ZN(n1075) );
XOR2_X1 U890 ( .A(G137), .B(n1196), .Z(n1195) );
NOR2_X1 U891 ( .A1(KEYINPUT47), .A2(n1197), .ZN(n1196) );
XOR2_X1 U892 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U893 ( .A(n1200), .B(n1201), .ZN(n1199) );
XNOR2_X1 U894 ( .A(G128), .B(G119), .ZN(n1198) );
NAND2_X1 U895 ( .A1(n1202), .A2(G221), .ZN(n1194) );
NAND2_X1 U896 ( .A1(KEYINPUT6), .A2(n1077), .ZN(n1193) );
NAND2_X1 U897 ( .A1(KEYINPUT55), .A2(n1035), .ZN(n1190) );
INV_X1 U898 ( .A(n1077), .ZN(n1035) );
NAND2_X1 U899 ( .A1(G217), .A2(n1203), .ZN(n1077) );
INV_X1 U900 ( .A(n1029), .ZN(n1182) );
XNOR2_X1 U901 ( .A(n1204), .B(G472), .ZN(n1029) );
NAND3_X1 U902 ( .A1(n1205), .A2(n1206), .A3(n1127), .ZN(n1204) );
NAND2_X1 U903 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
INV_X1 U904 ( .A(KEYINPUT44), .ZN(n1208) );
XOR2_X1 U905 ( .A(n1209), .B(n1210), .Z(n1207) );
NAND3_X1 U906 ( .A1(n1210), .A2(n1209), .A3(KEYINPUT44), .ZN(n1205) );
XNOR2_X1 U907 ( .A(n1101), .B(G101), .ZN(n1209) );
INV_X1 U908 ( .A(n1099), .ZN(n1101) );
NAND3_X1 U909 ( .A1(n1211), .A2(n1001), .A3(G210), .ZN(n1099) );
XNOR2_X1 U910 ( .A(n1110), .B(n1106), .ZN(n1210) );
XNOR2_X1 U911 ( .A(n1120), .B(n1107), .ZN(n1106) );
XNOR2_X1 U912 ( .A(n1212), .B(n1213), .ZN(n1110) );
XOR2_X1 U913 ( .A(G119), .B(G113), .Z(n1213) );
NAND2_X1 U914 ( .A1(KEYINPUT29), .A2(n1214), .ZN(n1212) );
XNOR2_X1 U915 ( .A(KEYINPUT28), .B(n1215), .ZN(n1214) );
NAND2_X1 U916 ( .A1(n1216), .A2(n1217), .ZN(n998) );
OR2_X1 U917 ( .A1(n1010), .A2(KEYINPUT46), .ZN(n1217) );
INV_X1 U918 ( .A(n981), .ZN(n1010) );
NOR2_X1 U919 ( .A1(n1030), .A2(n1188), .ZN(n981) );
NAND3_X1 U920 ( .A1(n1218), .A2(n1188), .A3(KEYINPUT46), .ZN(n1216) );
INV_X1 U921 ( .A(n1034), .ZN(n1188) );
XNOR2_X1 U922 ( .A(n1219), .B(G478), .ZN(n1034) );
NAND2_X1 U923 ( .A1(n1220), .A2(n1127), .ZN(n1219) );
XNOR2_X1 U924 ( .A(n1082), .B(KEYINPUT60), .ZN(n1220) );
XNOR2_X1 U925 ( .A(n1221), .B(n1222), .ZN(n1082) );
XOR2_X1 U926 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U927 ( .A(G107), .B(n1225), .Z(n1224) );
NOR2_X1 U928 ( .A1(KEYINPUT41), .A2(n1226), .ZN(n1225) );
AND2_X1 U929 ( .A1(n1202), .A2(G217), .ZN(n1223) );
AND2_X1 U930 ( .A1(G234), .A2(n1001), .ZN(n1202) );
XNOR2_X1 U931 ( .A(G116), .B(n1227), .ZN(n1221) );
XNOR2_X1 U932 ( .A(G134), .B(n1179), .ZN(n1227) );
INV_X1 U933 ( .A(n1030), .ZN(n1218) );
XNOR2_X1 U934 ( .A(n1228), .B(G475), .ZN(n1030) );
NAND2_X1 U935 ( .A1(n1127), .A2(n1086), .ZN(n1228) );
NAND3_X1 U936 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1086) );
NAND2_X1 U937 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND2_X1 U938 ( .A1(n1234), .A2(n1235), .ZN(n1232) );
XOR2_X1 U939 ( .A(KEYINPUT3), .B(n1236), .Z(n1234) );
NAND3_X1 U940 ( .A1(n1237), .A2(n1236), .A3(n1235), .ZN(n1230) );
INV_X1 U941 ( .A(n1233), .ZN(n1237) );
NAND2_X1 U942 ( .A1(n1238), .A2(n1239), .ZN(n1233) );
NAND2_X1 U943 ( .A1(n1240), .A2(G104), .ZN(n1239) );
XOR2_X1 U944 ( .A(KEYINPUT0), .B(n1241), .Z(n1238) );
NOR2_X1 U945 ( .A1(G104), .A2(n1240), .ZN(n1241) );
XNOR2_X1 U946 ( .A(G122), .B(n1242), .ZN(n1240) );
NOR2_X1 U947 ( .A1(G113), .A2(KEYINPUT54), .ZN(n1242) );
OR2_X1 U948 ( .A1(n1235), .A2(n1236), .ZN(n1229) );
XNOR2_X1 U949 ( .A(n1243), .B(n1244), .ZN(n1236) );
XNOR2_X1 U950 ( .A(n1245), .B(n1246), .ZN(n1244) );
AND3_X1 U951 ( .A1(G214), .A2(n1001), .A3(n1211), .ZN(n1246) );
INV_X1 U952 ( .A(G131), .ZN(n1245) );
XOR2_X1 U953 ( .A(n1200), .B(n1247), .Z(n1243) );
XNOR2_X1 U954 ( .A(G125), .B(n1248), .ZN(n1200) );
XNOR2_X1 U955 ( .A(n1156), .B(G140), .ZN(n1248) );
INV_X1 U956 ( .A(KEYINPUT24), .ZN(n1235) );
INV_X1 U957 ( .A(n1149), .ZN(n980) );
NAND3_X1 U958 ( .A1(n995), .A2(n993), .A3(n1185), .ZN(n1149) );
AND2_X1 U959 ( .A1(n1249), .A2(n1184), .ZN(n1185) );
NAND2_X1 U960 ( .A1(n1005), .A2(n1250), .ZN(n1184) );
NAND3_X1 U961 ( .A1(n1069), .A2(n1178), .A3(G902), .ZN(n1250) );
NOR2_X1 U962 ( .A1(G898), .A2(n1001), .ZN(n1069) );
NAND3_X1 U963 ( .A1(n1178), .A2(n1001), .A3(G952), .ZN(n1005) );
NAND2_X1 U964 ( .A1(G237), .A2(G234), .ZN(n1178) );
XNOR2_X1 U965 ( .A(KEYINPUT56), .B(n1019), .ZN(n1249) );
INV_X1 U966 ( .A(n1160), .ZN(n1019) );
NOR2_X1 U967 ( .A1(n1022), .A2(n1021), .ZN(n1160) );
INV_X1 U968 ( .A(n1173), .ZN(n1021) );
NAND2_X1 U969 ( .A1(G214), .A2(n1251), .ZN(n1173) );
XOR2_X1 U970 ( .A(n1252), .B(n1033), .Z(n1022) );
AND2_X1 U971 ( .A1(n1253), .A2(n1127), .ZN(n1033) );
XOR2_X1 U972 ( .A(n1125), .B(n1254), .Z(n1253) );
NOR2_X1 U973 ( .A1(KEYINPUT34), .A2(n1255), .ZN(n1254) );
XNOR2_X1 U974 ( .A(n1107), .B(n1050), .ZN(n1255) );
INV_X1 U975 ( .A(G125), .ZN(n1050) );
XNOR2_X1 U976 ( .A(G146), .B(n1256), .ZN(n1107) );
XOR2_X1 U977 ( .A(n1064), .B(n1257), .Z(n1125) );
NOR2_X1 U978 ( .A1(G953), .A2(n1068), .ZN(n1257) );
INV_X1 U979 ( .A(G224), .ZN(n1068) );
XOR2_X1 U980 ( .A(n1258), .B(n1259), .Z(n1064) );
XOR2_X1 U981 ( .A(n1260), .B(n1261), .Z(n1259) );
XNOR2_X1 U982 ( .A(n1215), .B(G113), .ZN(n1261) );
INV_X1 U983 ( .A(G116), .ZN(n1215) );
XNOR2_X1 U984 ( .A(KEYINPUT22), .B(n1179), .ZN(n1260) );
INV_X1 U985 ( .A(G122), .ZN(n1179) );
XOR2_X1 U986 ( .A(n1262), .B(n1263), .Z(n1258) );
XOR2_X1 U987 ( .A(n1264), .B(n1265), .Z(n1263) );
NOR2_X1 U988 ( .A1(G119), .A2(KEYINPUT10), .ZN(n1264) );
XNOR2_X1 U989 ( .A(G110), .B(n1266), .ZN(n1262) );
NOR2_X1 U990 ( .A1(G101), .A2(KEYINPUT38), .ZN(n1266) );
NAND2_X1 U991 ( .A1(KEYINPUT9), .A2(n1031), .ZN(n1252) );
AND2_X1 U992 ( .A1(G210), .A2(n1251), .ZN(n1031) );
NAND2_X1 U993 ( .A1(n1211), .A2(n1127), .ZN(n1251) );
INV_X1 U994 ( .A(G237), .ZN(n1211) );
NAND2_X1 U995 ( .A1(G221), .A2(n1203), .ZN(n993) );
NAND2_X1 U996 ( .A1(G234), .A2(n1127), .ZN(n1203) );
XNOR2_X1 U997 ( .A(n1267), .B(G469), .ZN(n995) );
NAND3_X1 U998 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1267) );
XNOR2_X1 U999 ( .A(KEYINPUT20), .B(n1127), .ZN(n1270) );
INV_X1 U1000 ( .A(G902), .ZN(n1127) );
NAND2_X1 U1001 ( .A1(n1271), .A2(n1048), .ZN(n1269) );
INV_X1 U1002 ( .A(n1120), .ZN(n1048) );
XNOR2_X1 U1003 ( .A(n1272), .B(KEYINPUT58), .ZN(n1271) );
NAND2_X1 U1004 ( .A1(n1273), .A2(n1120), .ZN(n1268) );
XNOR2_X1 U1005 ( .A(n1274), .B(n1275), .ZN(n1120) );
XOR2_X1 U1006 ( .A(KEYINPUT2), .B(G137), .Z(n1275) );
XNOR2_X1 U1007 ( .A(G131), .B(G134), .ZN(n1274) );
XNOR2_X1 U1008 ( .A(KEYINPUT12), .B(n1276), .ZN(n1273) );
INV_X1 U1009 ( .A(n1272), .ZN(n1276) );
XNOR2_X1 U1010 ( .A(n1277), .B(n1278), .ZN(n1272) );
XOR2_X1 U1011 ( .A(KEYINPUT7), .B(n1279), .Z(n1278) );
NOR2_X1 U1012 ( .A1(KEYINPUT37), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U1013 ( .A(G140), .B(n1281), .ZN(n1280) );
NAND2_X1 U1014 ( .A1(KEYINPUT17), .A2(n1201), .ZN(n1281) );
INV_X1 U1015 ( .A(G110), .ZN(n1201) );
XOR2_X1 U1016 ( .A(n1117), .B(n1114), .Z(n1277) );
NAND2_X1 U1017 ( .A1(n1282), .A2(n1001), .ZN(n1114) );
INV_X1 U1018 ( .A(G953), .ZN(n1001) );
XNOR2_X1 U1019 ( .A(G227), .B(KEYINPUT8), .ZN(n1282) );
XNOR2_X1 U1020 ( .A(n1283), .B(n1284), .ZN(n1117) );
XOR2_X1 U1021 ( .A(KEYINPUT16), .B(G101), .Z(n1284) );
XOR2_X1 U1022 ( .A(n1047), .B(n1265), .Z(n1283) );
XOR2_X1 U1023 ( .A(G107), .B(G104), .Z(n1265) );
XNOR2_X1 U1024 ( .A(n1256), .B(n1285), .ZN(n1047) );
NOR2_X1 U1025 ( .A1(KEYINPUT62), .A2(n1286), .ZN(n1285) );
XNOR2_X1 U1026 ( .A(KEYINPUT26), .B(n1156), .ZN(n1286) );
INV_X1 U1027 ( .A(G146), .ZN(n1156) );
XOR2_X1 U1028 ( .A(n1226), .B(KEYINPUT1), .Z(n1256) );
XOR2_X1 U1029 ( .A(G128), .B(n1247), .Z(n1226) );
XOR2_X1 U1030 ( .A(G143), .B(KEYINPUT42), .Z(n1247) );
XNOR2_X1 U1031 ( .A(G110), .B(KEYINPUT18), .ZN(n1189) );
endmodule


