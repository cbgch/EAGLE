//Key = 1101011111000010011100100000110110101110101110101011000110011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423;

NAND2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(G9) );
NAND2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U776 ( .A(KEYINPUT28), .B(n1080), .Z(n1076) );
NOR2_X1 U777 ( .A1(n1078), .A2(n1079), .ZN(n1080) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(G75) );
NOR4_X1 U779 ( .A1(G953), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1082) );
NOR2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR3_X1 U782 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
NOR3_X1 U783 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1091) );
NOR3_X1 U784 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
NOR2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(n1093) );
NOR2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR3_X1 U787 ( .A1(n1100), .A2(n1103), .A3(n1098), .ZN(n1088) );
NOR3_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
NOR2_X1 U789 ( .A1(n1107), .A2(n1092), .ZN(n1106) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1090), .ZN(n1104) );
NOR3_X1 U793 ( .A1(n1083), .A2(G953), .A3(G952), .ZN(n1081) );
AND4_X1 U794 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1083) );
NOR3_X1 U795 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
XOR2_X1 U796 ( .A(KEYINPUT45), .B(n1120), .Z(n1119) );
NOR2_X1 U797 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1118) );
XOR2_X1 U799 ( .A(KEYINPUT38), .B(n1125), .Z(n1124) );
NOR2_X1 U800 ( .A1(G475), .A2(KEYINPUT49), .ZN(n1123) );
NAND3_X1 U801 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1117) );
XOR2_X1 U802 ( .A(KEYINPUT43), .B(n1129), .Z(n1127) );
NOR3_X1 U803 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1115) );
AND2_X1 U804 ( .A1(n1122), .A2(n1121), .ZN(n1130) );
NAND2_X1 U805 ( .A1(G469), .A2(n1133), .ZN(n1114) );
XNOR2_X1 U806 ( .A(KEYINPUT42), .B(n1134), .ZN(n1113) );
XOR2_X1 U807 ( .A(n1135), .B(n1136), .Z(G72) );
NOR2_X1 U808 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U809 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NAND2_X1 U810 ( .A1(n1141), .A2(n1142), .ZN(n1135) );
NAND2_X1 U811 ( .A1(n1143), .A2(n1138), .ZN(n1142) );
XOR2_X1 U812 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND3_X1 U813 ( .A1(G900), .A2(n1145), .A3(G953), .ZN(n1141) );
XNOR2_X1 U814 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U815 ( .A(n1148), .B(n1149), .Z(n1146) );
XOR2_X1 U816 ( .A(n1150), .B(n1151), .Z(G69) );
XOR2_X1 U817 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U818 ( .A1(n1154), .A2(n1138), .ZN(n1153) );
XOR2_X1 U819 ( .A(n1155), .B(KEYINPUT46), .Z(n1154) );
NAND2_X1 U820 ( .A1(G898), .A2(G224), .ZN(n1155) );
NAND2_X1 U821 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
INV_X1 U822 ( .A(n1158), .ZN(n1157) );
NAND2_X1 U823 ( .A1(n1138), .A2(n1159), .ZN(n1150) );
NOR2_X1 U824 ( .A1(n1160), .A2(n1161), .ZN(G66) );
XOR2_X1 U825 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U826 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NOR2_X1 U827 ( .A1(n1160), .A2(n1166), .ZN(G63) );
XOR2_X1 U828 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND2_X1 U829 ( .A1(n1164), .A2(G478), .ZN(n1167) );
NOR2_X1 U830 ( .A1(n1160), .A2(n1169), .ZN(G60) );
NOR2_X1 U831 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U832 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U833 ( .A1(n1174), .A2(n1175), .ZN(n1170) );
XOR2_X1 U834 ( .A(KEYINPUT6), .B(n1173), .Z(n1175) );
AND2_X1 U835 ( .A1(n1164), .A2(G475), .ZN(n1173) );
XNOR2_X1 U836 ( .A(n1172), .B(KEYINPUT10), .ZN(n1174) );
XNOR2_X1 U837 ( .A(G104), .B(n1176), .ZN(G6) );
NOR2_X1 U838 ( .A1(n1160), .A2(n1177), .ZN(G57) );
XOR2_X1 U839 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U840 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U841 ( .A1(n1164), .A2(G472), .ZN(n1181) );
NAND3_X1 U842 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1180) );
NAND3_X1 U843 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NOR2_X1 U844 ( .A1(n1160), .A2(n1188), .ZN(G54) );
XOR2_X1 U845 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U846 ( .A(n1191), .B(n1192), .Z(n1190) );
NAND2_X1 U847 ( .A1(n1164), .A2(G469), .ZN(n1192) );
NAND2_X1 U848 ( .A1(n1193), .A2(n1194), .ZN(n1191) );
NAND2_X1 U849 ( .A1(G140), .A2(n1195), .ZN(n1194) );
XOR2_X1 U850 ( .A(KEYINPUT22), .B(n1196), .Z(n1193) );
NOR2_X1 U851 ( .A1(G140), .A2(n1195), .ZN(n1196) );
XNOR2_X1 U852 ( .A(n1197), .B(n1198), .ZN(n1189) );
NOR2_X1 U853 ( .A1(KEYINPUT2), .A2(n1149), .ZN(n1198) );
NOR2_X1 U854 ( .A1(n1160), .A2(n1199), .ZN(G51) );
XOR2_X1 U855 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND3_X1 U856 ( .A1(n1164), .A2(G210), .A3(KEYINPUT34), .ZN(n1201) );
AND2_X1 U857 ( .A1(G902), .A2(n1085), .ZN(n1164) );
OR2_X1 U858 ( .A1(n1144), .A2(n1159), .ZN(n1085) );
NAND4_X1 U859 ( .A1(n1176), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1159) );
NOR4_X1 U860 ( .A1(n1078), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1204) );
AND2_X1 U861 ( .A1(n1101), .A2(n1208), .ZN(n1078) );
NAND2_X1 U862 ( .A1(n1109), .A2(n1209), .ZN(n1203) );
NAND2_X1 U863 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XNOR2_X1 U864 ( .A(KEYINPUT50), .B(n1212), .ZN(n1210) );
NAND2_X1 U865 ( .A1(n1102), .A2(n1208), .ZN(n1176) );
NOR3_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1092), .ZN(n1208) );
NAND4_X1 U867 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1144) );
AND3_X1 U868 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1218) );
OR2_X1 U869 ( .A1(n1222), .A2(KEYINPUT25), .ZN(n1217) );
NAND2_X1 U870 ( .A1(n1223), .A2(n1224), .ZN(n1216) );
NAND2_X1 U871 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND2_X1 U872 ( .A1(n1105), .A2(n1101), .ZN(n1226) );
NAND2_X1 U873 ( .A1(n1102), .A2(n1227), .ZN(n1225) );
NAND3_X1 U874 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1227) );
NAND2_X1 U875 ( .A1(n1231), .A2(n1109), .ZN(n1230) );
OR3_X1 U876 ( .A1(n1090), .A2(n1232), .A3(KEYINPUT40), .ZN(n1229) );
NAND2_X1 U877 ( .A1(KEYINPUT40), .A2(n1105), .ZN(n1228) );
NOR2_X1 U878 ( .A1(n1233), .A2(n1090), .ZN(n1105) );
INV_X1 U879 ( .A(n1234), .ZN(n1090) );
NAND2_X1 U880 ( .A1(n1109), .A2(n1235), .ZN(n1215) );
NAND2_X1 U881 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND4_X1 U882 ( .A1(KEYINPUT25), .A2(n1223), .A3(n1101), .A4(n1238), .ZN(n1237) );
XNOR2_X1 U883 ( .A(KEYINPUT14), .B(n1239), .ZN(n1236) );
NAND3_X1 U884 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1200) );
NAND2_X1 U885 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NAND3_X1 U886 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1241) );
NAND2_X1 U887 ( .A1(n1248), .A2(n1249), .ZN(n1240) );
XNOR2_X1 U888 ( .A(n1246), .B(n1244), .ZN(n1248) );
INV_X1 U889 ( .A(n1245), .ZN(n1244) );
NOR2_X1 U890 ( .A1(KEYINPUT39), .A2(n1156), .ZN(n1245) );
NOR2_X1 U891 ( .A1(n1138), .A2(G952), .ZN(n1160) );
XOR2_X1 U892 ( .A(n1250), .B(n1251), .Z(G48) );
NAND2_X1 U893 ( .A1(n1252), .A2(KEYINPUT37), .ZN(n1251) );
XNOR2_X1 U894 ( .A(G146), .B(KEYINPUT19), .ZN(n1252) );
NAND4_X1 U895 ( .A1(n1253), .A2(n1102), .A3(n1254), .A4(n1231), .ZN(n1250) );
NOR2_X1 U896 ( .A1(n1255), .A2(n1214), .ZN(n1254) );
XNOR2_X1 U897 ( .A(n1256), .B(KEYINPUT15), .ZN(n1253) );
XOR2_X1 U898 ( .A(n1219), .B(n1257), .Z(G45) );
XNOR2_X1 U899 ( .A(G143), .B(KEYINPUT53), .ZN(n1257) );
NAND3_X1 U900 ( .A1(n1232), .A2(n1223), .A3(n1258), .ZN(n1219) );
NOR3_X1 U901 ( .A1(n1255), .A2(n1128), .A3(n1259), .ZN(n1258) );
XOR2_X1 U902 ( .A(n1221), .B(n1260), .Z(G42) );
XNOR2_X1 U903 ( .A(G140), .B(KEYINPUT41), .ZN(n1260) );
OR2_X1 U904 ( .A1(n1261), .A2(n1112), .ZN(n1221) );
INV_X1 U905 ( .A(n1262), .ZN(n1112) );
XNOR2_X1 U906 ( .A(G137), .B(n1220), .ZN(G39) );
NAND4_X1 U907 ( .A1(n1231), .A2(n1094), .A3(n1234), .A4(n1263), .ZN(n1220) );
XNOR2_X1 U908 ( .A(G134), .B(n1264), .ZN(G36) );
NAND4_X1 U909 ( .A1(n1265), .A2(n1232), .A3(n1223), .A4(n1101), .ZN(n1264) );
XNOR2_X1 U910 ( .A(n1234), .B(KEYINPUT17), .ZN(n1265) );
XOR2_X1 U911 ( .A(G131), .B(n1266), .Z(G33) );
NOR2_X1 U912 ( .A1(n1261), .A2(n1233), .ZN(n1266) );
NAND3_X1 U913 ( .A1(n1223), .A2(n1234), .A3(n1102), .ZN(n1261) );
NOR2_X1 U914 ( .A1(n1110), .A2(n1132), .ZN(n1234) );
XNOR2_X1 U915 ( .A(G128), .B(n1222), .ZN(G30) );
NAND4_X1 U916 ( .A1(n1223), .A2(n1231), .A3(n1101), .A4(n1109), .ZN(n1222) );
INV_X1 U917 ( .A(n1238), .ZN(n1231) );
NOR2_X1 U918 ( .A1(n1214), .A2(n1256), .ZN(n1223) );
INV_X1 U919 ( .A(n1263), .ZN(n1256) );
XNOR2_X1 U920 ( .A(G101), .B(n1202), .ZN(G3) );
NAND3_X1 U921 ( .A1(n1094), .A2(n1267), .A3(n1232), .ZN(n1202) );
INV_X1 U922 ( .A(n1233), .ZN(n1232) );
INV_X1 U923 ( .A(n1213), .ZN(n1267) );
XOR2_X1 U924 ( .A(G125), .B(n1268), .Z(G27) );
NOR2_X1 U925 ( .A1(n1239), .A2(n1269), .ZN(n1268) );
XNOR2_X1 U926 ( .A(KEYINPUT63), .B(n1255), .ZN(n1269) );
NAND4_X1 U927 ( .A1(n1270), .A2(n1102), .A3(n1262), .A4(n1263), .ZN(n1239) );
NAND2_X1 U928 ( .A1(n1087), .A2(n1271), .ZN(n1263) );
NAND4_X1 U929 ( .A1(G902), .A2(G953), .A3(n1272), .A4(n1140), .ZN(n1271) );
INV_X1 U930 ( .A(G900), .ZN(n1140) );
XNOR2_X1 U931 ( .A(n1273), .B(n1274), .ZN(G24) );
NOR2_X1 U932 ( .A1(n1255), .A2(n1212), .ZN(n1274) );
NAND3_X1 U933 ( .A1(n1270), .A2(n1275), .A3(n1276), .ZN(n1212) );
NOR3_X1 U934 ( .A1(n1259), .A2(n1277), .A3(n1128), .ZN(n1276) );
INV_X1 U935 ( .A(n1278), .ZN(n1277) );
INV_X1 U936 ( .A(n1100), .ZN(n1270) );
XNOR2_X1 U937 ( .A(n1279), .B(n1207), .ZN(G21) );
NOR4_X1 U938 ( .A1(n1100), .A2(n1238), .A3(n1098), .A4(n1213), .ZN(n1207) );
NAND2_X1 U939 ( .A1(n1280), .A2(n1281), .ZN(n1238) );
XNOR2_X1 U940 ( .A(KEYINPUT13), .B(n1134), .ZN(n1280) );
NAND2_X1 U941 ( .A1(n1282), .A2(n1283), .ZN(G18) );
NAND2_X1 U942 ( .A1(G116), .A2(n1284), .ZN(n1283) );
NAND2_X1 U943 ( .A1(n1206), .A2(n1285), .ZN(n1284) );
NAND2_X1 U944 ( .A1(KEYINPUT23), .A2(KEYINPUT1), .ZN(n1285) );
NAND3_X1 U945 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1282) );
INV_X1 U946 ( .A(KEYINPUT23), .ZN(n1288) );
NAND2_X1 U947 ( .A1(n1206), .A2(n1289), .ZN(n1287) );
INV_X1 U948 ( .A(KEYINPUT1), .ZN(n1289) );
NAND2_X1 U949 ( .A1(KEYINPUT1), .A2(n1290), .ZN(n1286) );
NAND2_X1 U950 ( .A1(n1206), .A2(n1291), .ZN(n1290) );
AND2_X1 U951 ( .A1(n1292), .A2(n1101), .ZN(n1206) );
NOR2_X1 U952 ( .A1(n1293), .A2(n1128), .ZN(n1101) );
XNOR2_X1 U953 ( .A(n1294), .B(n1205), .ZN(G15) );
AND2_X1 U954 ( .A1(n1292), .A2(n1102), .ZN(n1205) );
AND2_X1 U955 ( .A1(n1128), .A2(n1293), .ZN(n1102) );
NOR3_X1 U956 ( .A1(n1233), .A2(n1213), .A3(n1100), .ZN(n1292) );
NAND2_X1 U957 ( .A1(n1295), .A2(n1296), .ZN(n1100) );
NAND2_X1 U958 ( .A1(n1109), .A2(n1278), .ZN(n1213) );
NAND2_X1 U959 ( .A1(n1297), .A2(n1298), .ZN(n1233) );
XNOR2_X1 U960 ( .A(KEYINPUT51), .B(n1126), .ZN(n1297) );
INV_X1 U961 ( .A(n1281), .ZN(n1126) );
XNOR2_X1 U962 ( .A(n1195), .B(n1299), .ZN(G12) );
NOR2_X1 U963 ( .A1(n1300), .A2(n1255), .ZN(n1299) );
INV_X1 U964 ( .A(n1109), .ZN(n1255) );
NOR2_X1 U965 ( .A1(n1301), .A2(n1132), .ZN(n1109) );
INV_X1 U966 ( .A(n1111), .ZN(n1132) );
NAND2_X1 U967 ( .A1(G214), .A2(n1302), .ZN(n1111) );
INV_X1 U968 ( .A(n1110), .ZN(n1301) );
XNOR2_X1 U969 ( .A(n1121), .B(n1122), .ZN(n1110) );
NAND2_X1 U970 ( .A1(G210), .A2(n1302), .ZN(n1122) );
NAND2_X1 U971 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
INV_X1 U972 ( .A(G237), .ZN(n1303) );
AND2_X1 U973 ( .A1(n1305), .A2(n1304), .ZN(n1121) );
XOR2_X1 U974 ( .A(n1156), .B(n1306), .Z(n1305) );
NOR2_X1 U975 ( .A1(n1243), .A2(n1307), .ZN(n1306) );
XOR2_X1 U976 ( .A(n1308), .B(KEYINPUT59), .Z(n1307) );
NAND2_X1 U977 ( .A1(n1246), .A2(n1309), .ZN(n1308) );
XOR2_X1 U978 ( .A(KEYINPUT3), .B(n1247), .Z(n1309) );
INV_X1 U979 ( .A(n1249), .ZN(n1247) );
NOR2_X1 U980 ( .A1(n1249), .A2(n1246), .ZN(n1243) );
XOR2_X1 U981 ( .A(n1310), .B(n1311), .Z(n1246) );
XOR2_X1 U982 ( .A(KEYINPUT61), .B(G125), .Z(n1311) );
NAND2_X1 U983 ( .A1(n1312), .A2(n1138), .ZN(n1249) );
XOR2_X1 U984 ( .A(KEYINPUT21), .B(G224), .Z(n1312) );
XOR2_X1 U985 ( .A(n1313), .B(n1314), .Z(n1156) );
XOR2_X1 U986 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U987 ( .A(n1195), .B(n1317), .ZN(n1316) );
NOR2_X1 U988 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XOR2_X1 U989 ( .A(KEYINPUT5), .B(KEYINPUT31), .Z(n1319) );
NOR2_X1 U990 ( .A1(n1320), .A2(n1321), .ZN(n1315) );
XOR2_X1 U991 ( .A(n1322), .B(n1323), .Z(n1313) );
NOR2_X1 U992 ( .A1(KEYINPUT27), .A2(n1324), .ZN(n1323) );
XOR2_X1 U993 ( .A(n1211), .B(KEYINPUT30), .Z(n1300) );
NAND3_X1 U994 ( .A1(n1262), .A2(n1278), .A3(n1094), .ZN(n1211) );
NOR2_X1 U995 ( .A1(n1098), .A2(n1214), .ZN(n1094) );
NAND2_X1 U996 ( .A1(n1296), .A2(n1096), .ZN(n1214) );
INV_X1 U997 ( .A(n1295), .ZN(n1096) );
NOR2_X1 U998 ( .A1(n1325), .A2(n1129), .ZN(n1295) );
NOR2_X1 U999 ( .A1(n1133), .A2(G469), .ZN(n1129) );
AND2_X1 U1000 ( .A1(n1326), .A2(n1133), .ZN(n1325) );
NAND2_X1 U1001 ( .A1(n1327), .A2(n1328), .ZN(n1133) );
XNOR2_X1 U1002 ( .A(n1329), .B(n1330), .ZN(n1328) );
XNOR2_X1 U1003 ( .A(n1331), .B(n1149), .ZN(n1330) );
XNOR2_X1 U1004 ( .A(n1332), .B(n1333), .ZN(n1149) );
NOR2_X1 U1005 ( .A1(G143), .A2(KEYINPUT24), .ZN(n1333) );
NAND2_X1 U1006 ( .A1(KEYINPUT48), .A2(n1334), .ZN(n1331) );
XNOR2_X1 U1007 ( .A(G140), .B(n1195), .ZN(n1334) );
INV_X1 U1008 ( .A(n1197), .ZN(n1329) );
XNOR2_X1 U1009 ( .A(n1335), .B(n1336), .ZN(n1197) );
XNOR2_X1 U1010 ( .A(n1318), .B(n1185), .ZN(n1336) );
XOR2_X1 U1011 ( .A(n1337), .B(n1338), .Z(n1335) );
NOR2_X1 U1012 ( .A1(G953), .A2(n1139), .ZN(n1338) );
INV_X1 U1013 ( .A(G227), .ZN(n1139) );
XOR2_X1 U1014 ( .A(n1339), .B(KEYINPUT8), .Z(n1337) );
NAND3_X1 U1015 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1339) );
NAND2_X1 U1016 ( .A1(n1324), .A2(n1343), .ZN(n1342) );
INV_X1 U1017 ( .A(KEYINPUT56), .ZN(n1343) );
NAND3_X1 U1018 ( .A1(KEYINPUT56), .A2(n1344), .A3(n1079), .ZN(n1341) );
OR2_X1 U1019 ( .A1(n1079), .A2(n1344), .ZN(n1340) );
NOR2_X1 U1020 ( .A1(KEYINPUT54), .A2(n1324), .ZN(n1344) );
XOR2_X1 U1021 ( .A(G104), .B(KEYINPUT4), .Z(n1324) );
INV_X1 U1022 ( .A(G107), .ZN(n1079) );
XNOR2_X1 U1023 ( .A(KEYINPUT18), .B(n1304), .ZN(n1327) );
XNOR2_X1 U1024 ( .A(G469), .B(KEYINPUT32), .ZN(n1326) );
XNOR2_X1 U1025 ( .A(n1131), .B(KEYINPUT20), .ZN(n1296) );
INV_X1 U1026 ( .A(n1097), .ZN(n1131) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1345), .ZN(n1097) );
NAND2_X1 U1028 ( .A1(n1128), .A2(n1259), .ZN(n1098) );
INV_X1 U1029 ( .A(n1293), .ZN(n1259) );
XOR2_X1 U1030 ( .A(n1125), .B(G475), .Z(n1293) );
NOR2_X1 U1031 ( .A1(n1172), .A2(G902), .ZN(n1125) );
AND2_X1 U1032 ( .A1(n1346), .A2(n1347), .ZN(n1172) );
NAND2_X1 U1033 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1034 ( .A(KEYINPUT35), .B(n1350), .Z(n1348) );
XOR2_X1 U1035 ( .A(n1351), .B(KEYINPUT62), .Z(n1346) );
OR2_X1 U1036 ( .A1(n1349), .A2(n1350), .ZN(n1351) );
XOR2_X1 U1037 ( .A(G104), .B(n1352), .Z(n1350) );
XNOR2_X1 U1038 ( .A(n1273), .B(G113), .ZN(n1352) );
INV_X1 U1039 ( .A(G122), .ZN(n1273) );
XNOR2_X1 U1040 ( .A(n1353), .B(n1354), .ZN(n1349) );
XNOR2_X1 U1041 ( .A(n1355), .B(G131), .ZN(n1354) );
XOR2_X1 U1042 ( .A(n1356), .B(n1357), .Z(n1353) );
AND2_X1 U1043 ( .A1(n1358), .A2(G214), .ZN(n1357) );
NAND3_X1 U1044 ( .A1(n1359), .A2(n1360), .A3(KEYINPUT44), .ZN(n1356) );
NAND2_X1 U1045 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
NAND2_X1 U1046 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1047 ( .A1(G146), .A2(n1365), .ZN(n1364) );
INV_X1 U1048 ( .A(n1147), .ZN(n1361) );
NAND2_X1 U1049 ( .A1(n1366), .A2(n1367), .ZN(n1359) );
NAND2_X1 U1050 ( .A1(n1365), .A2(n1368), .ZN(n1366) );
NAND2_X1 U1051 ( .A1(n1147), .A2(n1363), .ZN(n1368) );
INV_X1 U1052 ( .A(KEYINPUT16), .ZN(n1363) );
XOR2_X1 U1053 ( .A(G125), .B(G140), .Z(n1147) );
INV_X1 U1054 ( .A(KEYINPUT52), .ZN(n1365) );
XOR2_X1 U1055 ( .A(n1369), .B(G478), .Z(n1128) );
NAND2_X1 U1056 ( .A1(n1168), .A2(n1304), .ZN(n1369) );
XNOR2_X1 U1057 ( .A(n1370), .B(n1371), .ZN(n1168) );
XOR2_X1 U1058 ( .A(n1372), .B(n1322), .Z(n1371) );
XNOR2_X1 U1059 ( .A(G122), .B(G107), .ZN(n1322) );
NAND2_X1 U1060 ( .A1(KEYINPUT55), .A2(n1373), .ZN(n1372) );
XOR2_X1 U1061 ( .A(G128), .B(n1374), .Z(n1373) );
XNOR2_X1 U1062 ( .A(n1355), .B(G134), .ZN(n1374) );
XNOR2_X1 U1063 ( .A(n1375), .B(n1291), .ZN(n1370) );
NAND3_X1 U1064 ( .A1(G217), .A2(n1138), .A3(G234), .ZN(n1375) );
NAND2_X1 U1065 ( .A1(n1087), .A2(n1376), .ZN(n1278) );
NAND3_X1 U1066 ( .A1(n1158), .A2(n1272), .A3(G902), .ZN(n1376) );
NOR2_X1 U1067 ( .A1(n1138), .A2(G898), .ZN(n1158) );
NAND3_X1 U1068 ( .A1(n1272), .A2(n1138), .A3(G952), .ZN(n1087) );
NAND2_X1 U1069 ( .A1(G237), .A2(G234), .ZN(n1272) );
NAND2_X1 U1070 ( .A1(n1377), .A2(n1378), .ZN(n1262) );
OR2_X1 U1071 ( .A1(n1092), .A2(KEYINPUT29), .ZN(n1378) );
INV_X1 U1072 ( .A(n1275), .ZN(n1092) );
NOR2_X1 U1073 ( .A1(n1281), .A2(n1298), .ZN(n1275) );
NAND3_X1 U1074 ( .A1(n1281), .A2(n1134), .A3(KEYINPUT29), .ZN(n1377) );
INV_X1 U1075 ( .A(n1298), .ZN(n1134) );
XNOR2_X1 U1076 ( .A(n1379), .B(G472), .ZN(n1298) );
NAND2_X1 U1077 ( .A1(n1380), .A2(n1304), .ZN(n1379) );
XOR2_X1 U1078 ( .A(n1381), .B(n1178), .Z(n1380) );
XOR2_X1 U1079 ( .A(n1382), .B(n1318), .Z(n1178) );
XOR2_X1 U1080 ( .A(G101), .B(KEYINPUT26), .Z(n1318) );
NAND2_X1 U1081 ( .A1(G210), .A2(n1358), .ZN(n1382) );
NOR2_X1 U1082 ( .A1(G953), .A2(G237), .ZN(n1358) );
NAND4_X1 U1083 ( .A1(n1383), .A2(n1183), .A3(n1384), .A4(n1385), .ZN(n1381) );
NAND3_X1 U1084 ( .A1(KEYINPUT33), .A2(n1386), .A3(n1387), .ZN(n1385) );
NAND3_X1 U1085 ( .A1(n1388), .A2(n1186), .A3(n1187), .ZN(n1384) );
OR2_X1 U1086 ( .A1(n1185), .A2(KEYINPUT33), .ZN(n1388) );
NAND3_X1 U1087 ( .A1(n1185), .A2(n1387), .A3(n1386), .ZN(n1183) );
INV_X1 U1088 ( .A(n1389), .ZN(n1185) );
OR2_X1 U1089 ( .A1(n1182), .A2(KEYINPUT33), .ZN(n1383) );
NAND2_X1 U1090 ( .A1(n1390), .A2(n1389), .ZN(n1182) );
XNOR2_X1 U1091 ( .A(n1148), .B(KEYINPUT58), .ZN(n1389) );
XNOR2_X1 U1092 ( .A(G131), .B(n1391), .ZN(n1148) );
XOR2_X1 U1093 ( .A(G137), .B(G134), .Z(n1391) );
XNOR2_X1 U1094 ( .A(n1386), .B(n1187), .ZN(n1390) );
INV_X1 U1095 ( .A(n1387), .ZN(n1187) );
XNOR2_X1 U1096 ( .A(n1310), .B(KEYINPUT36), .ZN(n1387) );
XOR2_X1 U1097 ( .A(n1392), .B(G128), .Z(n1310) );
NAND3_X1 U1098 ( .A1(n1393), .A2(n1394), .A3(n1395), .ZN(n1392) );
OR2_X1 U1099 ( .A1(n1367), .A2(KEYINPUT7), .ZN(n1395) );
NAND3_X1 U1100 ( .A1(KEYINPUT7), .A2(n1367), .A3(G143), .ZN(n1394) );
INV_X1 U1101 ( .A(G146), .ZN(n1367) );
NAND2_X1 U1102 ( .A1(n1396), .A2(n1355), .ZN(n1393) );
INV_X1 U1103 ( .A(G143), .ZN(n1355) );
NAND2_X1 U1104 ( .A1(n1397), .A2(KEYINPUT7), .ZN(n1396) );
XNOR2_X1 U1105 ( .A(G146), .B(KEYINPUT12), .ZN(n1397) );
INV_X1 U1106 ( .A(n1186), .ZN(n1386) );
NAND3_X1 U1107 ( .A1(n1398), .A2(n1399), .A3(n1400), .ZN(n1186) );
INV_X1 U1108 ( .A(n1320), .ZN(n1400) );
NOR3_X1 U1109 ( .A1(n1291), .A2(G119), .A3(n1294), .ZN(n1320) );
NAND2_X1 U1110 ( .A1(n1321), .A2(n1401), .ZN(n1399) );
INV_X1 U1111 ( .A(KEYINPUT57), .ZN(n1401) );
NAND2_X1 U1112 ( .A1(n1402), .A2(n1403), .ZN(n1321) );
NAND2_X1 U1113 ( .A1(n1404), .A2(n1294), .ZN(n1403) );
XNOR2_X1 U1114 ( .A(G116), .B(G119), .ZN(n1404) );
NAND3_X1 U1115 ( .A1(n1405), .A2(n1402), .A3(KEYINPUT57), .ZN(n1398) );
NAND3_X1 U1116 ( .A1(G113), .A2(n1291), .A3(G119), .ZN(n1402) );
NAND2_X1 U1117 ( .A1(n1406), .A2(n1294), .ZN(n1405) );
INV_X1 U1118 ( .A(G113), .ZN(n1294) );
NAND2_X1 U1119 ( .A1(G119), .A2(n1291), .ZN(n1406) );
INV_X1 U1120 ( .A(G116), .ZN(n1291) );
XNOR2_X1 U1121 ( .A(n1407), .B(n1165), .ZN(n1281) );
AND2_X1 U1122 ( .A1(G217), .A2(n1345), .ZN(n1165) );
NAND2_X1 U1123 ( .A1(G234), .A2(n1304), .ZN(n1345) );
NAND2_X1 U1124 ( .A1(n1163), .A2(n1304), .ZN(n1407) );
INV_X1 U1125 ( .A(G902), .ZN(n1304) );
XOR2_X1 U1126 ( .A(n1408), .B(n1409), .Z(n1163) );
XOR2_X1 U1127 ( .A(n1410), .B(n1332), .Z(n1409) );
XNOR2_X1 U1128 ( .A(G128), .B(G146), .ZN(n1332) );
NAND2_X1 U1129 ( .A1(KEYINPUT9), .A2(n1279), .ZN(n1410) );
INV_X1 U1130 ( .A(G119), .ZN(n1279) );
XOR2_X1 U1131 ( .A(n1411), .B(n1412), .Z(n1408) );
NOR3_X1 U1132 ( .A1(n1413), .A2(n1414), .A3(n1415), .ZN(n1412) );
AND2_X1 U1133 ( .A1(n1416), .A2(G137), .ZN(n1415) );
NOR3_X1 U1134 ( .A1(G137), .A2(KEYINPUT47), .A3(n1416), .ZN(n1414) );
NAND2_X1 U1135 ( .A1(KEYINPUT0), .A2(n1417), .ZN(n1416) );
NOR2_X1 U1136 ( .A1(n1417), .A2(n1418), .ZN(n1413) );
INV_X1 U1137 ( .A(KEYINPUT47), .ZN(n1418) );
AND3_X1 U1138 ( .A1(G234), .A2(n1138), .A3(G221), .ZN(n1417) );
INV_X1 U1139 ( .A(G953), .ZN(n1138) );
XNOR2_X1 U1140 ( .A(n1419), .B(n1195), .ZN(n1411) );
NAND2_X1 U1141 ( .A1(n1420), .A2(n1421), .ZN(n1419) );
OR2_X1 U1142 ( .A1(n1422), .A2(G125), .ZN(n1421) );
XOR2_X1 U1143 ( .A(n1423), .B(KEYINPUT11), .Z(n1420) );
NAND2_X1 U1144 ( .A1(G125), .A2(n1422), .ZN(n1423) );
XOR2_X1 U1145 ( .A(G140), .B(KEYINPUT60), .Z(n1422) );
INV_X1 U1146 ( .A(G110), .ZN(n1195) );
endmodule


