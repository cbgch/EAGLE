//Key = 1110011100110101100100111100001111011111001011001000100110000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362;

XNOR2_X1 U742 ( .A(G107), .B(n1033), .ZN(G9) );
NOR2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR4_X1 U744 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
XOR2_X1 U745 ( .A(n1040), .B(KEYINPUT7), .Z(n1039) );
NAND3_X1 U746 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1038) );
XNOR2_X1 U748 ( .A(n1046), .B(KEYINPUT60), .ZN(n1044) );
NAND4_X1 U749 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1036) );
NAND3_X1 U750 ( .A1(n1041), .A2(n1051), .A3(n1052), .ZN(n1048) );
NAND2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND3_X1 U752 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U753 ( .A1(n1058), .A2(n1059), .ZN(n1053) );
NAND2_X1 U754 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U755 ( .A1(n1055), .A2(n1062), .ZN(n1061) );
NAND2_X1 U756 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U757 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U758 ( .A1(n1057), .A2(n1067), .ZN(n1060) );
NAND2_X1 U759 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U760 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND3_X1 U761 ( .A1(n1072), .A2(n1073), .A3(n1046), .ZN(n1047) );
AND2_X1 U762 ( .A1(n1043), .A2(n1058), .ZN(n1046) );
AND3_X1 U763 ( .A1(n1057), .A2(n1055), .A3(n1052), .ZN(n1043) );
INV_X1 U764 ( .A(n1074), .ZN(n1052) );
NOR3_X1 U765 ( .A1(n1075), .A2(G953), .A3(G952), .ZN(n1034) );
INV_X1 U766 ( .A(n1049), .ZN(n1075) );
NAND4_X1 U767 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1049) );
NOR4_X1 U768 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1079) );
XOR2_X1 U769 ( .A(n1084), .B(n1085), .Z(n1083) );
XOR2_X1 U770 ( .A(KEYINPUT5), .B(n1086), .Z(n1082) );
NOR4_X1 U771 ( .A1(n1072), .A2(n1065), .A3(n1087), .A4(n1088), .ZN(n1086) );
XOR2_X1 U772 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR3_X1 U773 ( .A1(n1091), .A2(KEYINPUT12), .A3(n1092), .ZN(n1081) );
AND2_X1 U774 ( .A1(n1091), .A2(KEYINPUT12), .ZN(n1080) );
XOR2_X1 U775 ( .A(n1093), .B(G478), .Z(n1078) );
NAND2_X1 U776 ( .A1(KEYINPUT52), .A2(n1094), .ZN(n1093) );
XOR2_X1 U777 ( .A(n1095), .B(n1096), .Z(G72) );
NOR2_X1 U778 ( .A1(n1097), .A2(n1050), .ZN(n1096) );
AND2_X1 U779 ( .A1(G227), .A2(G900), .ZN(n1097) );
NAND2_X1 U780 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
NAND2_X1 U781 ( .A1(n1100), .A2(n1050), .ZN(n1099) );
XOR2_X1 U782 ( .A(n1101), .B(n1102), .Z(n1100) );
OR3_X1 U783 ( .A1(n1103), .A2(n1102), .A3(n1050), .ZN(n1098) );
XNOR2_X1 U784 ( .A(n1104), .B(n1105), .ZN(n1102) );
XOR2_X1 U785 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U786 ( .A(KEYINPUT58), .B(G140), .Z(n1107) );
NOR2_X1 U787 ( .A1(G125), .A2(KEYINPUT53), .ZN(n1106) );
XOR2_X1 U788 ( .A(n1108), .B(n1109), .Z(n1104) );
XOR2_X1 U789 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(G69) );
NAND2_X1 U791 ( .A1(n1114), .A2(n1050), .ZN(n1113) );
XOR2_X1 U792 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U793 ( .A1(n1117), .A2(G953), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U795 ( .A1(n1115), .A2(n1120), .ZN(n1119) );
NAND2_X1 U796 ( .A1(G224), .A2(n1121), .ZN(n1118) );
NAND2_X1 U797 ( .A1(G898), .A2(n1115), .ZN(n1121) );
NAND2_X1 U798 ( .A1(n1122), .A2(n1123), .ZN(n1115) );
NAND2_X1 U799 ( .A1(G953), .A2(n1124), .ZN(n1123) );
XOR2_X1 U800 ( .A(n1125), .B(n1126), .Z(n1122) );
XNOR2_X1 U801 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U802 ( .A1(KEYINPUT4), .A2(n1129), .ZN(n1128) );
XOR2_X1 U803 ( .A(G101), .B(n1130), .Z(n1129) );
NAND2_X1 U804 ( .A1(KEYINPUT55), .A2(n1131), .ZN(n1127) );
NOR2_X1 U805 ( .A1(n1132), .A2(n1133), .ZN(G66) );
NOR2_X1 U806 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U807 ( .A(n1136), .B(KEYINPUT37), .Z(n1135) );
NAND2_X1 U808 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U809 ( .A1(n1139), .A2(n1037), .ZN(n1138) );
NOR3_X1 U810 ( .A1(n1140), .A2(n1141), .A3(n1137), .ZN(n1134) );
NOR2_X1 U811 ( .A1(n1132), .A2(n1142), .ZN(G63) );
XOR2_X1 U812 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U813 ( .A(KEYINPUT42), .B(n1145), .Z(n1144) );
NOR2_X1 U814 ( .A1(n1146), .A2(n1140), .ZN(n1145) );
INV_X1 U815 ( .A(G478), .ZN(n1146) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1147), .ZN(G60) );
NOR2_X1 U817 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U818 ( .A(n1150), .B(KEYINPUT35), .Z(n1149) );
NAND2_X1 U819 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U820 ( .A1(n1151), .A2(n1152), .ZN(n1148) );
NOR2_X1 U821 ( .A1(n1140), .A2(n1153), .ZN(n1151) );
XOR2_X1 U822 ( .A(G104), .B(n1154), .Z(G6) );
NOR2_X1 U823 ( .A1(KEYINPUT28), .A2(n1155), .ZN(n1154) );
NOR2_X1 U824 ( .A1(n1132), .A2(n1156), .ZN(G57) );
XOR2_X1 U825 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U826 ( .A1(n1084), .A2(n1140), .ZN(n1157) );
NOR2_X1 U827 ( .A1(n1132), .A2(n1159), .ZN(G54) );
XOR2_X1 U828 ( .A(n1160), .B(n1161), .Z(n1159) );
NOR2_X1 U829 ( .A1(n1162), .A2(n1140), .ZN(n1161) );
INV_X1 U830 ( .A(G469), .ZN(n1162) );
NAND2_X1 U831 ( .A1(n1163), .A2(KEYINPUT25), .ZN(n1160) );
XNOR2_X1 U832 ( .A(n1164), .B(n1165), .ZN(n1163) );
XOR2_X1 U833 ( .A(n1166), .B(n1167), .Z(n1164) );
NOR2_X1 U834 ( .A1(n1132), .A2(n1168), .ZN(G51) );
XOR2_X1 U835 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U836 ( .A1(n1090), .A2(n1140), .ZN(n1170) );
NAND2_X1 U837 ( .A1(G902), .A2(n1037), .ZN(n1140) );
NAND2_X1 U838 ( .A1(n1116), .A2(n1101), .ZN(n1037) );
AND4_X1 U839 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1101) );
NOR4_X1 U840 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
INV_X1 U841 ( .A(n1179), .ZN(n1178) );
NOR3_X1 U842 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1176) );
NOR2_X1 U843 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
INV_X1 U844 ( .A(KEYINPUT54), .ZN(n1184) );
NOR3_X1 U845 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1183) );
NOR2_X1 U846 ( .A1(KEYINPUT54), .A2(n1188), .ZN(n1181) );
NOR3_X1 U847 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1173) );
NOR2_X1 U848 ( .A1(n1045), .A2(n1192), .ZN(n1191) );
NOR3_X1 U849 ( .A1(n1193), .A2(KEYINPUT23), .A3(n1194), .ZN(n1190) );
AND2_X1 U850 ( .A1(n1195), .A2(KEYINPUT23), .ZN(n1189) );
AND4_X1 U851 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1116) );
NOR4_X1 U852 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NOR2_X1 U853 ( .A1(n1045), .A2(n1204), .ZN(n1203) );
INV_X1 U854 ( .A(n1155), .ZN(n1202) );
NAND3_X1 U855 ( .A1(n1205), .A2(n1055), .A3(n1042), .ZN(n1155) );
AND2_X1 U856 ( .A1(n1206), .A2(n1033), .ZN(n1198) );
NAND3_X1 U857 ( .A1(n1055), .A2(n1056), .A3(n1205), .ZN(n1033) );
NAND2_X1 U858 ( .A1(n1207), .A2(KEYINPUT36), .ZN(n1169) );
XOR2_X1 U859 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U860 ( .A(KEYINPUT41), .B(n1210), .Z(n1209) );
NOR2_X1 U861 ( .A1(n1050), .A2(G952), .ZN(n1132) );
XNOR2_X1 U862 ( .A(G146), .B(n1171), .ZN(G48) );
NAND3_X1 U863 ( .A1(n1211), .A2(n1042), .A3(n1212), .ZN(n1171) );
XOR2_X1 U864 ( .A(n1213), .B(n1214), .Z(G45) );
NAND3_X1 U865 ( .A1(n1193), .A2(n1215), .A3(KEYINPUT39), .ZN(n1214) );
XNOR2_X1 U866 ( .A(KEYINPUT27), .B(n1192), .ZN(n1215) );
NAND3_X1 U867 ( .A1(n1216), .A2(n1217), .A3(n1212), .ZN(n1192) );
XOR2_X1 U868 ( .A(n1172), .B(n1218), .Z(G42) );
XOR2_X1 U869 ( .A(n1219), .B(KEYINPUT59), .Z(n1218) );
NAND2_X1 U870 ( .A1(n1220), .A2(n1188), .ZN(n1172) );
XOR2_X1 U871 ( .A(n1221), .B(n1222), .Z(G39) );
NOR2_X1 U872 ( .A1(KEYINPUT34), .A2(n1223), .ZN(n1222) );
INV_X1 U873 ( .A(G137), .ZN(n1223) );
NAND2_X1 U874 ( .A1(n1224), .A2(n1225), .ZN(n1221) );
NAND4_X1 U875 ( .A1(n1226), .A2(n1188), .A3(n1227), .A4(n1228), .ZN(n1225) );
INV_X1 U876 ( .A(KEYINPUT2), .ZN(n1228) );
NOR2_X1 U877 ( .A1(n1058), .A2(n1229), .ZN(n1227) );
NAND2_X1 U878 ( .A1(n1175), .A2(KEYINPUT2), .ZN(n1224) );
AND4_X1 U879 ( .A1(n1226), .A2(n1188), .A3(n1058), .A4(n1071), .ZN(n1175) );
XNOR2_X1 U880 ( .A(G134), .B(n1230), .ZN(G36) );
NAND2_X1 U881 ( .A1(n1188), .A2(n1231), .ZN(n1230) );
XOR2_X1 U882 ( .A(n1232), .B(n1179), .Z(G33) );
NAND3_X1 U883 ( .A1(n1042), .A2(n1217), .A3(n1188), .ZN(n1179) );
AND2_X1 U884 ( .A1(n1041), .A2(n1212), .ZN(n1188) );
INV_X1 U885 ( .A(n1185), .ZN(n1041) );
NAND2_X1 U886 ( .A1(n1073), .A2(n1233), .ZN(n1185) );
XNOR2_X1 U887 ( .A(n1177), .B(n1234), .ZN(G30) );
NOR2_X1 U888 ( .A1(G128), .A2(KEYINPUT51), .ZN(n1234) );
AND3_X1 U889 ( .A1(n1211), .A2(n1056), .A3(n1212), .ZN(n1177) );
NOR2_X1 U890 ( .A1(n1063), .A2(n1187), .ZN(n1212) );
INV_X1 U891 ( .A(n1235), .ZN(n1187) );
INV_X1 U892 ( .A(n1186), .ZN(n1063) );
XOR2_X1 U893 ( .A(n1206), .B(n1236), .Z(G3) );
XOR2_X1 U894 ( .A(KEYINPUT11), .B(G101), .Z(n1236) );
NAND3_X1 U895 ( .A1(n1058), .A2(n1205), .A3(n1217), .ZN(n1206) );
NAND3_X1 U896 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(G27) );
NAND2_X1 U897 ( .A1(KEYINPUT3), .A2(n1240), .ZN(n1239) );
OR3_X1 U898 ( .A1(n1240), .A2(KEYINPUT3), .A3(G125), .ZN(n1238) );
INV_X1 U899 ( .A(n1195), .ZN(n1240) );
NAND2_X1 U900 ( .A1(G125), .A2(n1241), .ZN(n1237) );
NAND2_X1 U901 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
INV_X1 U902 ( .A(KEYINPUT3), .ZN(n1243) );
XOR2_X1 U903 ( .A(KEYINPUT50), .B(n1195), .Z(n1242) );
NOR2_X1 U904 ( .A1(n1194), .A2(n1045), .ZN(n1195) );
NAND3_X1 U905 ( .A1(n1057), .A2(n1235), .A3(n1220), .ZN(n1194) );
AND3_X1 U906 ( .A1(n1070), .A2(n1071), .A3(n1042), .ZN(n1220) );
NAND2_X1 U907 ( .A1(n1074), .A2(n1244), .ZN(n1235) );
NAND4_X1 U908 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1103), .ZN(n1244) );
INV_X1 U909 ( .A(G900), .ZN(n1103) );
NAND2_X1 U910 ( .A1(n1246), .A2(n1247), .ZN(G24) );
NAND2_X1 U911 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
INV_X1 U912 ( .A(G122), .ZN(n1249) );
NAND2_X1 U913 ( .A1(G122), .A2(n1250), .ZN(n1246) );
NAND2_X1 U914 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U915 ( .A1(n1201), .A2(n1253), .ZN(n1252) );
INV_X1 U916 ( .A(n1254), .ZN(n1201) );
OR2_X1 U917 ( .A1(n1253), .A2(n1248), .ZN(n1251) );
NOR2_X1 U918 ( .A1(KEYINPUT20), .A2(n1254), .ZN(n1248) );
NAND4_X1 U919 ( .A1(n1216), .A2(n1255), .A3(n1055), .A4(n1193), .ZN(n1254) );
AND2_X1 U920 ( .A1(n1229), .A2(n1070), .ZN(n1055) );
AND2_X1 U921 ( .A1(n1256), .A2(n1257), .ZN(n1216) );
XOR2_X1 U922 ( .A(KEYINPUT40), .B(n1258), .Z(n1256) );
INV_X1 U923 ( .A(KEYINPUT30), .ZN(n1253) );
XOR2_X1 U924 ( .A(n1200), .B(n1259), .Z(G21) );
NOR2_X1 U925 ( .A1(KEYINPUT47), .A2(n1260), .ZN(n1259) );
AND3_X1 U926 ( .A1(n1255), .A2(n1058), .A3(n1211), .ZN(n1200) );
AND3_X1 U927 ( .A1(n1193), .A2(n1071), .A3(n1226), .ZN(n1211) );
XOR2_X1 U928 ( .A(G116), .B(n1261), .Z(G18) );
NOR3_X1 U929 ( .A1(n1262), .A2(KEYINPUT63), .A3(n1045), .ZN(n1261) );
INV_X1 U930 ( .A(n1193), .ZN(n1045) );
XNOR2_X1 U931 ( .A(KEYINPUT56), .B(n1204), .ZN(n1262) );
NAND2_X1 U932 ( .A1(n1231), .A2(n1255), .ZN(n1204) );
INV_X1 U933 ( .A(n1180), .ZN(n1231) );
NAND2_X1 U934 ( .A1(n1217), .A2(n1056), .ZN(n1180) );
AND2_X1 U935 ( .A1(n1076), .A2(n1257), .ZN(n1056) );
XNOR2_X1 U936 ( .A(G113), .B(n1196), .ZN(G15) );
NAND4_X1 U937 ( .A1(n1042), .A2(n1217), .A3(n1255), .A4(n1193), .ZN(n1196) );
AND2_X1 U938 ( .A1(n1057), .A2(n1263), .ZN(n1255) );
AND2_X1 U939 ( .A1(n1066), .A2(n1264), .ZN(n1057) );
INV_X1 U940 ( .A(n1068), .ZN(n1217) );
NAND2_X1 U941 ( .A1(n1226), .A2(n1229), .ZN(n1068) );
INV_X1 U942 ( .A(n1071), .ZN(n1229) );
XOR2_X1 U943 ( .A(n1265), .B(KEYINPUT17), .Z(n1226) );
NOR2_X1 U944 ( .A1(n1257), .A2(n1076), .ZN(n1042) );
INV_X1 U945 ( .A(n1258), .ZN(n1076) );
XNOR2_X1 U946 ( .A(G110), .B(n1197), .ZN(G12) );
NAND4_X1 U947 ( .A1(n1058), .A2(n1205), .A3(n1070), .A4(n1071), .ZN(n1197) );
NAND2_X1 U948 ( .A1(n1266), .A2(n1267), .ZN(n1071) );
NAND2_X1 U949 ( .A1(n1268), .A2(n1141), .ZN(n1267) );
NAND2_X1 U950 ( .A1(n1269), .A2(n1091), .ZN(n1268) );
NAND2_X1 U951 ( .A1(n1139), .A2(n1269), .ZN(n1266) );
INV_X1 U952 ( .A(KEYINPUT14), .ZN(n1269) );
INV_X1 U953 ( .A(n1077), .ZN(n1139) );
NAND2_X1 U954 ( .A1(n1092), .A2(n1091), .ZN(n1077) );
NAND2_X1 U955 ( .A1(n1137), .A2(n1270), .ZN(n1091) );
XNOR2_X1 U956 ( .A(n1271), .B(n1272), .ZN(n1137) );
XOR2_X1 U957 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U958 ( .A(n1275), .B(n1276), .ZN(n1274) );
NAND2_X1 U959 ( .A1(KEYINPUT45), .A2(n1277), .ZN(n1276) );
NAND2_X1 U960 ( .A1(KEYINPUT61), .A2(n1278), .ZN(n1275) );
XOR2_X1 U961 ( .A(G125), .B(n1279), .Z(n1278) );
XOR2_X1 U962 ( .A(G146), .B(G140), .Z(n1279) );
NAND2_X1 U963 ( .A1(n1280), .A2(G221), .ZN(n1273) );
XOR2_X1 U964 ( .A(n1281), .B(n1282), .Z(n1271) );
XOR2_X1 U965 ( .A(KEYINPUT0), .B(G137), .Z(n1282) );
XOR2_X1 U966 ( .A(n1260), .B(G110), .Z(n1281) );
INV_X1 U967 ( .A(G119), .ZN(n1260) );
INV_X1 U968 ( .A(n1141), .ZN(n1092) );
NAND2_X1 U969 ( .A1(G217), .A2(n1283), .ZN(n1141) );
XNOR2_X1 U970 ( .A(n1265), .B(KEYINPUT18), .ZN(n1070) );
NAND2_X1 U971 ( .A1(n1284), .A2(n1285), .ZN(n1265) );
NAND2_X1 U972 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U973 ( .A1(G472), .A2(n1288), .ZN(n1287) );
NAND2_X1 U974 ( .A1(KEYINPUT49), .A2(KEYINPUT32), .ZN(n1288) );
NAND3_X1 U975 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1284) );
INV_X1 U976 ( .A(KEYINPUT49), .ZN(n1291) );
OR2_X1 U977 ( .A1(n1084), .A2(KEYINPUT32), .ZN(n1290) );
INV_X1 U978 ( .A(G472), .ZN(n1084) );
NAND2_X1 U979 ( .A1(KEYINPUT32), .A2(n1292), .ZN(n1289) );
NAND2_X1 U980 ( .A1(G472), .A2(n1085), .ZN(n1292) );
INV_X1 U981 ( .A(n1286), .ZN(n1085) );
NOR2_X1 U982 ( .A1(n1158), .A2(G902), .ZN(n1286) );
XNOR2_X1 U983 ( .A(n1293), .B(n1294), .ZN(n1158) );
XOR2_X1 U984 ( .A(KEYINPUT6), .B(n1295), .Z(n1294) );
AND2_X1 U985 ( .A1(G210), .A2(n1296), .ZN(n1295) );
XOR2_X1 U986 ( .A(n1297), .B(n1167), .Z(n1293) );
AND3_X1 U987 ( .A1(n1186), .A2(n1263), .A3(n1193), .ZN(n1205) );
NOR2_X1 U988 ( .A1(n1073), .A2(n1072), .ZN(n1193) );
INV_X1 U989 ( .A(n1233), .ZN(n1072) );
NAND2_X1 U990 ( .A1(G214), .A2(n1298), .ZN(n1233) );
XNOR2_X1 U991 ( .A(n1089), .B(n1299), .ZN(n1073) );
NOR2_X1 U992 ( .A1(n1300), .A2(KEYINPUT46), .ZN(n1299) );
INV_X1 U993 ( .A(n1090), .ZN(n1300) );
NAND2_X1 U994 ( .A1(G210), .A2(n1298), .ZN(n1090) );
NAND2_X1 U995 ( .A1(n1301), .A2(n1270), .ZN(n1298) );
INV_X1 U996 ( .A(G237), .ZN(n1301) );
NAND2_X1 U997 ( .A1(n1302), .A2(n1270), .ZN(n1089) );
XOR2_X1 U998 ( .A(n1303), .B(n1304), .Z(n1302) );
INV_X1 U999 ( .A(n1208), .ZN(n1304) );
XOR2_X1 U1000 ( .A(n1305), .B(n1306), .Z(n1208) );
XOR2_X1 U1001 ( .A(n1131), .B(n1130), .Z(n1306) );
XNOR2_X1 U1002 ( .A(n1307), .B(n1308), .ZN(n1130) );
NOR2_X1 U1003 ( .A1(KEYINPUT21), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1004 ( .A(G107), .B(KEYINPUT10), .ZN(n1307) );
XOR2_X1 U1005 ( .A(G122), .B(n1310), .Z(n1131) );
NOR2_X1 U1006 ( .A1(G110), .A2(KEYINPUT29), .ZN(n1310) );
XOR2_X1 U1007 ( .A(n1297), .B(G125), .Z(n1305) );
XOR2_X1 U1008 ( .A(n1311), .B(n1312), .Z(n1297) );
XOR2_X1 U1009 ( .A(G128), .B(G101), .Z(n1312) );
XOR2_X1 U1010 ( .A(n1313), .B(n1125), .Z(n1311) );
XOR2_X1 U1011 ( .A(G113), .B(n1314), .Z(n1125) );
XOR2_X1 U1012 ( .A(G119), .B(G116), .Z(n1314) );
NAND2_X1 U1013 ( .A1(n1315), .A2(n1316), .ZN(n1313) );
OR2_X1 U1014 ( .A1(n1317), .A2(G146), .ZN(n1316) );
XOR2_X1 U1015 ( .A(n1318), .B(KEYINPUT8), .Z(n1315) );
NAND2_X1 U1016 ( .A1(G146), .A2(n1317), .ZN(n1318) );
XNOR2_X1 U1017 ( .A(n1213), .B(KEYINPUT1), .ZN(n1317) );
INV_X1 U1018 ( .A(G143), .ZN(n1213) );
NAND2_X1 U1019 ( .A1(KEYINPUT38), .A2(n1210), .ZN(n1303) );
NOR2_X1 U1020 ( .A1(n1120), .A2(G953), .ZN(n1210) );
INV_X1 U1021 ( .A(G224), .ZN(n1120) );
NAND2_X1 U1022 ( .A1(n1074), .A2(n1319), .ZN(n1263) );
NAND4_X1 U1023 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1124), .ZN(n1319) );
INV_X1 U1024 ( .A(G898), .ZN(n1124) );
NAND3_X1 U1025 ( .A1(n1245), .A2(n1050), .A3(G952), .ZN(n1074) );
NAND2_X1 U1026 ( .A1(G237), .A2(n1320), .ZN(n1245) );
NOR2_X1 U1027 ( .A1(n1066), .A2(n1065), .ZN(n1186) );
INV_X1 U1028 ( .A(n1264), .ZN(n1065) );
NAND2_X1 U1029 ( .A1(G221), .A2(n1283), .ZN(n1264) );
NAND2_X1 U1030 ( .A1(n1320), .A2(n1270), .ZN(n1283) );
XOR2_X1 U1031 ( .A(G234), .B(KEYINPUT26), .Z(n1320) );
XOR2_X1 U1032 ( .A(n1087), .B(KEYINPUT22), .Z(n1066) );
XNOR2_X1 U1033 ( .A(n1321), .B(G469), .ZN(n1087) );
NAND2_X1 U1034 ( .A1(n1322), .A2(n1270), .ZN(n1321) );
XOR2_X1 U1035 ( .A(n1323), .B(n1324), .Z(n1322) );
XNOR2_X1 U1036 ( .A(n1325), .B(KEYINPUT43), .ZN(n1324) );
NAND2_X1 U1037 ( .A1(KEYINPUT15), .A2(n1165), .ZN(n1325) );
XOR2_X1 U1038 ( .A(G110), .B(n1219), .Z(n1165) );
NAND2_X1 U1039 ( .A1(n1326), .A2(n1327), .ZN(n1323) );
NAND2_X1 U1040 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1041 ( .A(KEYINPUT9), .B(n1330), .Z(n1328) );
NAND2_X1 U1042 ( .A1(n1331), .A2(n1167), .ZN(n1326) );
INV_X1 U1043 ( .A(n1329), .ZN(n1167) );
XOR2_X1 U1044 ( .A(n1332), .B(n1111), .Z(n1329) );
XOR2_X1 U1045 ( .A(G134), .B(G137), .Z(n1111) );
NAND2_X1 U1046 ( .A1(KEYINPUT13), .A2(n1232), .ZN(n1332) );
INV_X1 U1047 ( .A(G131), .ZN(n1232) );
XOR2_X1 U1048 ( .A(KEYINPUT24), .B(n1330), .Z(n1331) );
INV_X1 U1049 ( .A(n1166), .ZN(n1330) );
XOR2_X1 U1050 ( .A(n1333), .B(n1334), .Z(n1166) );
XOR2_X1 U1051 ( .A(G101), .B(n1335), .Z(n1334) );
XOR2_X1 U1052 ( .A(KEYINPUT16), .B(G104), .Z(n1335) );
XOR2_X1 U1053 ( .A(n1336), .B(n1337), .Z(n1333) );
INV_X1 U1054 ( .A(n1108), .ZN(n1337) );
XOR2_X1 U1055 ( .A(n1338), .B(G146), .Z(n1108) );
NAND2_X1 U1056 ( .A1(KEYINPUT19), .A2(n1277), .ZN(n1338) );
XOR2_X1 U1057 ( .A(n1339), .B(n1340), .Z(n1336) );
NAND2_X1 U1058 ( .A1(G227), .A2(n1050), .ZN(n1339) );
NOR2_X1 U1059 ( .A1(n1257), .A2(n1258), .ZN(n1058) );
XOR2_X1 U1060 ( .A(n1341), .B(n1153), .Z(n1258) );
INV_X1 U1061 ( .A(G475), .ZN(n1153) );
OR2_X1 U1062 ( .A1(n1152), .A2(G902), .ZN(n1341) );
XNOR2_X1 U1063 ( .A(n1342), .B(n1343), .ZN(n1152) );
XOR2_X1 U1064 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1065 ( .A1(KEYINPUT31), .A2(n1219), .ZN(n1345) );
INV_X1 U1066 ( .A(G140), .ZN(n1219) );
NAND2_X1 U1067 ( .A1(n1346), .A2(KEYINPUT33), .ZN(n1344) );
XOR2_X1 U1068 ( .A(n1347), .B(n1110), .Z(n1346) );
XOR2_X1 U1069 ( .A(G131), .B(G143), .Z(n1110) );
NAND2_X1 U1070 ( .A1(n1296), .A2(G214), .ZN(n1347) );
NOR2_X1 U1071 ( .A1(G953), .A2(G237), .ZN(n1296) );
XOR2_X1 U1072 ( .A(n1348), .B(n1349), .Z(n1342) );
XOR2_X1 U1073 ( .A(G146), .B(G125), .Z(n1349) );
NAND3_X1 U1074 ( .A1(n1350), .A2(n1351), .A3(KEYINPUT44), .ZN(n1348) );
NAND2_X1 U1075 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
INV_X1 U1076 ( .A(KEYINPUT57), .ZN(n1353) );
XOR2_X1 U1077 ( .A(n1309), .B(n1354), .Z(n1352) );
NAND2_X1 U1078 ( .A1(KEYINPUT48), .A2(n1355), .ZN(n1354) );
NAND3_X1 U1079 ( .A1(n1355), .A2(n1356), .A3(KEYINPUT57), .ZN(n1350) );
XOR2_X1 U1080 ( .A(KEYINPUT48), .B(n1309), .Z(n1356) );
INV_X1 U1081 ( .A(G104), .ZN(n1309) );
XOR2_X1 U1082 ( .A(G113), .B(G122), .Z(n1355) );
XOR2_X1 U1083 ( .A(n1094), .B(G478), .Z(n1257) );
AND2_X1 U1084 ( .A1(n1143), .A2(n1270), .ZN(n1094) );
INV_X1 U1085 ( .A(G902), .ZN(n1270) );
XOR2_X1 U1086 ( .A(n1357), .B(n1358), .Z(n1143) );
XNOR2_X1 U1087 ( .A(n1359), .B(n1340), .ZN(n1358) );
XOR2_X1 U1088 ( .A(G107), .B(G143), .Z(n1340) );
NAND2_X1 U1089 ( .A1(n1280), .A2(G217), .ZN(n1359) );
AND2_X1 U1090 ( .A1(G234), .A2(n1050), .ZN(n1280) );
INV_X1 U1091 ( .A(G953), .ZN(n1050) );
XOR2_X1 U1092 ( .A(n1360), .B(n1361), .Z(n1357) );
NOR2_X1 U1093 ( .A1(KEYINPUT62), .A2(n1362), .ZN(n1361) );
XOR2_X1 U1094 ( .A(G122), .B(G116), .Z(n1362) );
XOR2_X1 U1095 ( .A(G134), .B(n1277), .Z(n1360) );
INV_X1 U1096 ( .A(G128), .ZN(n1277) );
endmodule


