//Key = 1001011011001100010000011101000000011011011101000110011111100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312;

XNOR2_X1 U725 ( .A(G107), .B(n997), .ZN(G9) );
NOR2_X1 U726 ( .A1(n998), .A2(n999), .ZN(G75) );
NOR4_X1 U727 ( .A1(n1000), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n999) );
NOR3_X1 U728 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1002) );
NOR2_X1 U729 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR2_X1 U730 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NOR2_X1 U731 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U732 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
XOR2_X1 U733 ( .A(n1015), .B(KEYINPUT32), .Z(n1013) );
NAND2_X1 U734 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
AND3_X1 U735 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1011) );
AND4_X1 U736 ( .A1(n1021), .A2(n1018), .A3(n1022), .A4(n1023), .ZN(n1007) );
XOR2_X1 U737 ( .A(KEYINPUT36), .B(n1024), .Z(n1001) );
NOR2_X1 U738 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR2_X1 U739 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
INV_X1 U740 ( .A(n1029), .ZN(n1028) );
NOR2_X1 U741 ( .A1(n1030), .A2(n1031), .ZN(n1027) );
AND2_X1 U742 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
AND2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(n1030) );
NOR4_X1 U744 ( .A1(n1036), .A2(n1006), .A3(n1010), .A4(n1004), .ZN(n1025) );
NOR2_X1 U745 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U746 ( .A1(n1039), .A2(n1014), .ZN(n1038) );
NOR2_X1 U747 ( .A1(n1040), .A2(n1041), .ZN(n1037) );
NAND3_X1 U748 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1000) );
NAND3_X1 U749 ( .A1(n1034), .A2(n1045), .A3(n1029), .ZN(n1044) );
NOR3_X1 U750 ( .A1(n1040), .A2(n1014), .A3(n1004), .ZN(n1029) );
NOR3_X1 U751 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n998) );
INV_X1 U752 ( .A(n1042), .ZN(n1046) );
NAND4_X1 U753 ( .A1(n1020), .A2(n1018), .A3(n1047), .A4(n1048), .ZN(n1042) );
NOR4_X1 U754 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
XNOR2_X1 U755 ( .A(KEYINPUT20), .B(n1053), .ZN(n1052) );
XNOR2_X1 U756 ( .A(n1054), .B(n1055), .ZN(n1051) );
XNOR2_X1 U757 ( .A(KEYINPUT4), .B(n1056), .ZN(n1050) );
XOR2_X1 U758 ( .A(n1057), .B(n1058), .Z(n1049) );
NAND2_X1 U759 ( .A1(KEYINPUT49), .A2(n1059), .ZN(n1058) );
NOR2_X1 U760 ( .A1(n1022), .A2(n1060), .ZN(n1047) );
NOR2_X1 U761 ( .A1(KEYINPUT49), .A2(n1059), .ZN(n1060) );
XNOR2_X1 U762 ( .A(n1061), .B(KEYINPUT45), .ZN(n1059) );
XOR2_X1 U763 ( .A(n1062), .B(n1063), .Z(G72) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1043), .ZN(n1063) );
AND2_X1 U765 ( .A1(G227), .A2(G900), .ZN(n1064) );
NAND3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1062) );
NAND3_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
INV_X1 U768 ( .A(n1071), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1072), .A2(n1043), .ZN(n1069) );
NAND2_X1 U770 ( .A1(G953), .A2(n1073), .ZN(n1068) );
NAND3_X1 U771 ( .A1(KEYINPUT24), .A2(n1071), .A3(n1074), .ZN(n1066) );
NAND2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1071) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XNOR2_X1 U774 ( .A(n1079), .B(n1080), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1075) );
XNOR2_X1 U776 ( .A(n1083), .B(n1084), .ZN(n1082) );
OR2_X1 U777 ( .A1(n1074), .A2(KEYINPUT24), .ZN(n1065) );
AND2_X1 U778 ( .A1(n1043), .A2(n1072), .ZN(n1074) );
NAND2_X1 U779 ( .A1(n1085), .A2(n1086), .ZN(n1072) );
XNOR2_X1 U780 ( .A(KEYINPUT13), .B(n1087), .ZN(n1086) );
XOR2_X1 U781 ( .A(n1088), .B(n1089), .Z(G69) );
XOR2_X1 U782 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U784 ( .A(KEYINPUT54), .B(n1043), .ZN(n1093) );
AND2_X1 U785 ( .A1(G224), .A2(G898), .ZN(n1092) );
NAND2_X1 U786 ( .A1(n1043), .A2(n1094), .ZN(n1090) );
NAND2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XNOR2_X1 U788 ( .A(KEYINPUT17), .B(n1097), .ZN(n1096) );
NAND2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1088) );
INV_X1 U790 ( .A(n1100), .ZN(n1099) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(n1098) );
XNOR2_X1 U792 ( .A(n1103), .B(G110), .ZN(n1102) );
NOR2_X1 U793 ( .A1(KEYINPUT60), .A2(n1104), .ZN(n1101) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(G66) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U796 ( .A1(KEYINPUT59), .A2(n1109), .ZN(n1108) );
NOR2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NOR2_X1 U798 ( .A1(n1105), .A2(n1112), .ZN(G63) );
NOR3_X1 U799 ( .A1(n1055), .A2(n1113), .A3(n1114), .ZN(n1112) );
NOR4_X1 U800 ( .A1(n1115), .A2(n1111), .A3(KEYINPUT46), .A4(n1054), .ZN(n1114) );
NOR2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
NOR3_X1 U802 ( .A1(n1054), .A2(KEYINPUT46), .A3(n1118), .ZN(n1116) );
INV_X1 U803 ( .A(G478), .ZN(n1054) );
NOR2_X1 U804 ( .A1(n1105), .A2(n1119), .ZN(G60) );
XNOR2_X1 U805 ( .A(n1120), .B(n1121), .ZN(n1119) );
AND2_X1 U806 ( .A1(G475), .A2(n1122), .ZN(n1121) );
XNOR2_X1 U807 ( .A(n1123), .B(n1124), .ZN(G6) );
NAND2_X1 U808 ( .A1(KEYINPUT38), .A2(n1125), .ZN(n1123) );
NOR3_X1 U809 ( .A1(n1105), .A2(n1126), .A3(n1127), .ZN(G57) );
NOR2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1129) );
AND2_X1 U812 ( .A1(n1132), .A2(KEYINPUT50), .ZN(n1131) );
INV_X1 U813 ( .A(n1133), .ZN(n1128) );
NOR2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(n1126) );
XOR2_X1 U815 ( .A(n1130), .B(n1135), .Z(n1134) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1132), .ZN(n1135) );
XOR2_X1 U817 ( .A(n1080), .B(n1137), .Z(n1132) );
NOR2_X1 U818 ( .A1(KEYINPUT22), .A2(n1138), .ZN(n1137) );
INV_X1 U819 ( .A(KEYINPUT50), .ZN(n1136) );
XOR2_X1 U820 ( .A(n1139), .B(n1140), .Z(n1130) );
XOR2_X1 U821 ( .A(n1141), .B(n1142), .Z(n1140) );
AND2_X1 U822 ( .A1(G472), .A2(n1122), .ZN(n1142) );
NOR2_X1 U823 ( .A1(KEYINPUT21), .A2(n1143), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1144), .B(KEYINPUT14), .Z(n1143) );
XNOR2_X1 U825 ( .A(G101), .B(KEYINPUT26), .ZN(n1139) );
NOR2_X1 U826 ( .A1(n1105), .A2(n1145), .ZN(G54) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U828 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U829 ( .A1(KEYINPUT5), .A2(n1150), .ZN(n1148) );
NAND2_X1 U830 ( .A1(n1122), .A2(G469), .ZN(n1150) );
XNOR2_X1 U831 ( .A(n1151), .B(KEYINPUT15), .ZN(n1146) );
NAND2_X1 U832 ( .A1(KEYINPUT35), .A2(G140), .ZN(n1151) );
NOR2_X1 U833 ( .A1(n1105), .A2(n1152), .ZN(G51) );
XOR2_X1 U834 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1111), .ZN(n1154) );
INV_X1 U836 ( .A(n1122), .ZN(n1111) );
NOR2_X1 U837 ( .A1(n1156), .A2(n1118), .ZN(n1122) );
INV_X1 U838 ( .A(n1003), .ZN(n1118) );
NAND4_X1 U839 ( .A1(n1095), .A2(n1085), .A3(n1087), .A4(n1097), .ZN(n1003) );
AND4_X1 U840 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1085) );
NOR3_X1 U841 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
NAND2_X1 U842 ( .A1(n1045), .A2(n1164), .ZN(n1159) );
NAND2_X1 U843 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U844 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XNOR2_X1 U845 ( .A(n1169), .B(KEYINPUT58), .ZN(n1167) );
NAND2_X1 U846 ( .A1(n1170), .A2(n1018), .ZN(n1165) );
NAND3_X1 U847 ( .A1(n1035), .A2(n1018), .A3(n1170), .ZN(n1157) );
AND4_X1 U848 ( .A1(n1124), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1095) );
AND4_X1 U849 ( .A1(n997), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1173) );
NAND3_X1 U850 ( .A1(n1045), .A2(n1021), .A3(n1177), .ZN(n997) );
NAND4_X1 U851 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1045), .ZN(n1172) );
XNOR2_X1 U852 ( .A(n1169), .B(KEYINPUT9), .ZN(n1178) );
NAND3_X1 U853 ( .A1(n1177), .A2(n1021), .A3(n1035), .ZN(n1124) );
NOR2_X1 U854 ( .A1(n1181), .A2(n1182), .ZN(n1153) );
XOR2_X1 U855 ( .A(KEYINPUT40), .B(n1183), .Z(n1182) );
AND2_X1 U856 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U857 ( .A1(n1185), .A2(n1184), .ZN(n1181) );
XOR2_X1 U858 ( .A(n1186), .B(n1187), .Z(n1184) );
INV_X1 U859 ( .A(G110), .ZN(n1187) );
XNOR2_X1 U860 ( .A(n1188), .B(n1189), .ZN(n1185) );
XNOR2_X1 U861 ( .A(KEYINPUT52), .B(n1190), .ZN(n1189) );
XOR2_X1 U862 ( .A(n1191), .B(n1192), .Z(n1188) );
NAND2_X1 U863 ( .A1(KEYINPUT8), .A2(n1079), .ZN(n1191) );
NOR2_X1 U864 ( .A1(n1043), .A2(G952), .ZN(n1105) );
XNOR2_X1 U865 ( .A(G146), .B(n1158), .ZN(G48) );
NAND3_X1 U866 ( .A1(n1035), .A2(n1169), .A3(n1168), .ZN(n1158) );
INV_X1 U867 ( .A(n1193), .ZN(n1168) );
XNOR2_X1 U868 ( .A(n1194), .B(n1161), .ZN(G45) );
AND2_X1 U869 ( .A1(n1170), .A2(n1195), .ZN(n1161) );
XNOR2_X1 U870 ( .A(G140), .B(n1087), .ZN(G42) );
NAND3_X1 U871 ( .A1(n1018), .A2(n1032), .A3(n1196), .ZN(n1087) );
XOR2_X1 U872 ( .A(G137), .B(n1163), .Z(G39) );
NOR3_X1 U873 ( .A1(n1006), .A2(n1040), .A3(n1193), .ZN(n1163) );
INV_X1 U874 ( .A(n1033), .ZN(n1006) );
XOR2_X1 U875 ( .A(n1197), .B(G134), .Z(G36) );
NAND2_X1 U876 ( .A1(KEYINPUT23), .A2(n1198), .ZN(n1197) );
NAND3_X1 U877 ( .A1(n1170), .A2(n1045), .A3(n1199), .ZN(n1198) );
XNOR2_X1 U878 ( .A(n1018), .B(KEYINPUT3), .ZN(n1199) );
XNOR2_X1 U879 ( .A(G131), .B(n1200), .ZN(G33) );
NAND3_X1 U880 ( .A1(n1170), .A2(n1035), .A3(n1201), .ZN(n1200) );
XNOR2_X1 U881 ( .A(n1018), .B(KEYINPUT57), .ZN(n1201) );
INV_X1 U882 ( .A(n1040), .ZN(n1018) );
NAND2_X1 U883 ( .A1(n1017), .A2(n1202), .ZN(n1040) );
AND3_X1 U884 ( .A1(n1032), .A2(n1203), .A3(n1179), .ZN(n1170) );
XNOR2_X1 U885 ( .A(n1084), .B(n1204), .ZN(G30) );
NOR3_X1 U886 ( .A1(n1193), .A2(n1205), .A3(n1206), .ZN(n1204) );
XNOR2_X1 U887 ( .A(n1169), .B(KEYINPUT18), .ZN(n1205) );
NAND4_X1 U888 ( .A1(n1032), .A2(n1207), .A3(n1019), .A4(n1203), .ZN(n1193) );
XOR2_X1 U889 ( .A(n1097), .B(n1208), .Z(G3) );
NOR2_X1 U890 ( .A1(G101), .A2(KEYINPUT1), .ZN(n1208) );
NAND3_X1 U891 ( .A1(n1033), .A2(n1177), .A3(n1179), .ZN(n1097) );
XNOR2_X1 U892 ( .A(n1190), .B(n1162), .ZN(G27) );
AND3_X1 U893 ( .A1(n1034), .A2(n1169), .A3(n1196), .ZN(n1162) );
AND4_X1 U894 ( .A1(n1020), .A2(n1035), .A3(n1019), .A4(n1203), .ZN(n1196) );
NAND2_X1 U895 ( .A1(n1004), .A2(n1209), .ZN(n1203) );
NAND4_X1 U896 ( .A1(G902), .A2(G953), .A3(n1210), .A4(n1073), .ZN(n1209) );
INV_X1 U897 ( .A(G900), .ZN(n1073) );
XNOR2_X1 U898 ( .A(G122), .B(n1171), .ZN(G24) );
NAND3_X1 U899 ( .A1(n1180), .A2(n1021), .A3(n1195), .ZN(n1171) );
NOR3_X1 U900 ( .A1(n1039), .A2(n1053), .A3(n1211), .ZN(n1195) );
INV_X1 U901 ( .A(n1169), .ZN(n1039) );
INV_X1 U902 ( .A(n1014), .ZN(n1021) );
NAND2_X1 U903 ( .A1(n1056), .A2(n1020), .ZN(n1014) );
NAND3_X1 U904 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(G21) );
NAND2_X1 U905 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U906 ( .A1(n1217), .A2(KEYINPUT25), .ZN(n1216) );
XOR2_X1 U907 ( .A(n1176), .B(KEYINPUT11), .Z(n1217) );
INV_X1 U908 ( .A(n1218), .ZN(n1215) );
NAND3_X1 U909 ( .A1(KEYINPUT25), .A2(n1218), .A3(n1176), .ZN(n1213) );
XOR2_X1 U910 ( .A(G119), .B(KEYINPUT31), .Z(n1218) );
OR2_X1 U911 ( .A1(n1176), .A2(KEYINPUT25), .ZN(n1212) );
NAND4_X1 U912 ( .A1(n1180), .A2(n1033), .A3(n1219), .A4(n1169), .ZN(n1176) );
NOR2_X1 U913 ( .A1(n1056), .A2(n1220), .ZN(n1219) );
INV_X1 U914 ( .A(n1019), .ZN(n1056) );
XNOR2_X1 U915 ( .A(G116), .B(n1221), .ZN(G18) );
NAND4_X1 U916 ( .A1(n1222), .A2(n1223), .A3(n1169), .A4(n1224), .ZN(n1221) );
NOR2_X1 U917 ( .A1(n1206), .A2(n1041), .ZN(n1224) );
INV_X1 U918 ( .A(n1179), .ZN(n1041) );
INV_X1 U919 ( .A(n1045), .ZN(n1206) );
NOR2_X1 U920 ( .A1(n1225), .A2(n1211), .ZN(n1045) );
XNOR2_X1 U921 ( .A(KEYINPUT19), .B(n1010), .ZN(n1222) );
XOR2_X1 U922 ( .A(G113), .B(n1226), .Z(G15) );
NOR2_X1 U923 ( .A1(KEYINPUT33), .A2(n1175), .ZN(n1226) );
NAND4_X1 U924 ( .A1(n1035), .A2(n1179), .A3(n1227), .A4(n1180), .ZN(n1175) );
AND2_X1 U925 ( .A1(n1034), .A2(n1223), .ZN(n1180) );
INV_X1 U926 ( .A(n1010), .ZN(n1034) );
NAND2_X1 U927 ( .A1(n1023), .A2(n1228), .ZN(n1010) );
NOR2_X1 U928 ( .A1(n1019), .A2(n1220), .ZN(n1179) );
INV_X1 U929 ( .A(n1207), .ZN(n1220) );
XNOR2_X1 U930 ( .A(n1020), .B(KEYINPUT63), .ZN(n1207) );
NOR2_X1 U931 ( .A1(n1229), .A2(n1053), .ZN(n1035) );
INV_X1 U932 ( .A(n1225), .ZN(n1053) );
XNOR2_X1 U933 ( .A(G110), .B(n1174), .ZN(G12) );
NAND4_X1 U934 ( .A1(n1033), .A2(n1177), .A3(n1020), .A4(n1019), .ZN(n1174) );
XOR2_X1 U935 ( .A(n1230), .B(n1110), .Z(n1019) );
NAND2_X1 U936 ( .A1(G217), .A2(n1231), .ZN(n1110) );
NAND2_X1 U937 ( .A1(n1156), .A2(n1109), .ZN(n1230) );
NAND2_X1 U938 ( .A1(n1232), .A2(n1233), .ZN(n1109) );
NAND2_X1 U939 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U940 ( .A(KEYINPUT41), .B(n1236), .Z(n1232) );
NOR2_X1 U941 ( .A1(n1234), .A2(n1235), .ZN(n1236) );
XOR2_X1 U942 ( .A(n1237), .B(n1238), .Z(n1235) );
XNOR2_X1 U943 ( .A(G119), .B(n1239), .ZN(n1238) );
NAND2_X1 U944 ( .A1(KEYINPUT39), .A2(n1240), .ZN(n1237) );
XOR2_X1 U945 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U946 ( .A(n1243), .B(G140), .Z(n1242) );
NAND2_X1 U947 ( .A1(KEYINPUT55), .A2(n1190), .ZN(n1243) );
XNOR2_X1 U948 ( .A(G146), .B(KEYINPUT42), .ZN(n1241) );
XOR2_X1 U949 ( .A(n1244), .B(n1245), .Z(n1234) );
AND3_X1 U950 ( .A1(n1246), .A2(G234), .A3(G221), .ZN(n1245) );
XNOR2_X1 U951 ( .A(G137), .B(KEYINPUT7), .ZN(n1244) );
XOR2_X1 U952 ( .A(n1247), .B(G472), .Z(n1020) );
NAND2_X1 U953 ( .A1(n1248), .A2(n1156), .ZN(n1247) );
XOR2_X1 U954 ( .A(n1249), .B(n1250), .Z(n1248) );
XNOR2_X1 U955 ( .A(n1144), .B(n1251), .ZN(n1250) );
XOR2_X1 U956 ( .A(KEYINPUT61), .B(G101), .Z(n1251) );
NAND3_X1 U957 ( .A1(n1246), .A2(n1252), .A3(G210), .ZN(n1144) );
XNOR2_X1 U958 ( .A(n1133), .B(n1253), .ZN(n1249) );
XNOR2_X1 U959 ( .A(n1254), .B(n1079), .ZN(n1253) );
INV_X1 U960 ( .A(n1138), .ZN(n1079) );
XOR2_X1 U961 ( .A(G128), .B(n1255), .Z(n1138) );
NOR2_X1 U962 ( .A1(KEYINPUT28), .A2(n1256), .ZN(n1254) );
INV_X1 U963 ( .A(n1080), .ZN(n1256) );
XOR2_X1 U964 ( .A(n1257), .B(n1258), .Z(n1133) );
NOR2_X1 U965 ( .A1(KEYINPUT51), .A2(n1259), .ZN(n1258) );
XNOR2_X1 U966 ( .A(G119), .B(n1260), .ZN(n1259) );
NOR2_X1 U967 ( .A1(G116), .A2(KEYINPUT44), .ZN(n1260) );
AND3_X1 U968 ( .A1(n1227), .A2(n1223), .A3(n1032), .ZN(n1177) );
NOR2_X1 U969 ( .A1(n1023), .A2(n1022), .ZN(n1032) );
INV_X1 U970 ( .A(n1228), .ZN(n1022) );
NAND2_X1 U971 ( .A1(G221), .A2(n1231), .ZN(n1228) );
NAND2_X1 U972 ( .A1(G234), .A2(n1156), .ZN(n1231) );
XNOR2_X1 U973 ( .A(n1057), .B(n1261), .ZN(n1023) );
INV_X1 U974 ( .A(n1061), .ZN(n1261) );
XOR2_X1 U975 ( .A(G469), .B(KEYINPUT62), .Z(n1061) );
NAND2_X1 U976 ( .A1(n1262), .A2(n1156), .ZN(n1057) );
XOR2_X1 U977 ( .A(n1149), .B(n1263), .Z(n1262) );
XOR2_X1 U978 ( .A(KEYINPUT43), .B(G140), .Z(n1263) );
XOR2_X1 U979 ( .A(n1264), .B(n1265), .Z(n1149) );
XOR2_X1 U980 ( .A(n1266), .B(n1239), .Z(n1265) );
AND2_X1 U981 ( .A1(n1246), .A2(G227), .ZN(n1266) );
XOR2_X1 U982 ( .A(n1083), .B(n1267), .Z(n1264) );
XNOR2_X1 U983 ( .A(n1255), .B(n1080), .ZN(n1083) );
XNOR2_X1 U984 ( .A(n1268), .B(n1269), .ZN(n1080) );
XNOR2_X1 U985 ( .A(G131), .B(G137), .ZN(n1268) );
NAND2_X1 U986 ( .A1(n1004), .A2(n1270), .ZN(n1223) );
NAND3_X1 U987 ( .A1(n1100), .A2(n1210), .A3(G902), .ZN(n1270) );
NOR2_X1 U988 ( .A1(n1043), .A2(G898), .ZN(n1100) );
NAND3_X1 U989 ( .A1(n1210), .A2(n1043), .A3(G952), .ZN(n1004) );
INV_X1 U990 ( .A(G953), .ZN(n1043) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1210) );
XNOR2_X1 U992 ( .A(n1169), .B(KEYINPUT12), .ZN(n1227) );
NOR2_X1 U993 ( .A1(n1017), .A2(n1016), .ZN(n1169) );
INV_X1 U994 ( .A(n1202), .ZN(n1016) );
NAND2_X1 U995 ( .A1(G214), .A2(n1271), .ZN(n1202) );
XNOR2_X1 U996 ( .A(n1272), .B(n1155), .ZN(n1017) );
NAND2_X1 U997 ( .A1(G210), .A2(n1271), .ZN(n1155) );
NAND2_X1 U998 ( .A1(n1252), .A2(n1156), .ZN(n1271) );
NAND2_X1 U999 ( .A1(n1273), .A2(n1156), .ZN(n1272) );
XOR2_X1 U1000 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U1001 ( .A(n1186), .B(n1276), .Z(n1275) );
XNOR2_X1 U1002 ( .A(n1239), .B(n1255), .ZN(n1276) );
XNOR2_X1 U1003 ( .A(G110), .B(n1084), .ZN(n1239) );
XNOR2_X1 U1004 ( .A(n1104), .B(G122), .ZN(n1186) );
XNOR2_X1 U1005 ( .A(n1277), .B(n1278), .ZN(n1104) );
XNOR2_X1 U1006 ( .A(n1279), .B(G116), .ZN(n1278) );
INV_X1 U1007 ( .A(G119), .ZN(n1279) );
XNOR2_X1 U1008 ( .A(n1267), .B(n1257), .ZN(n1277) );
XOR2_X1 U1009 ( .A(G113), .B(KEYINPUT10), .Z(n1257) );
XOR2_X1 U1010 ( .A(G101), .B(n1280), .Z(n1267) );
XNOR2_X1 U1011 ( .A(G107), .B(n1125), .ZN(n1280) );
XOR2_X1 U1012 ( .A(n1281), .B(n1282), .Z(n1274) );
XOR2_X1 U1013 ( .A(n1283), .B(n1192), .Z(n1282) );
AND2_X1 U1014 ( .A1(n1246), .A2(n1284), .ZN(n1192) );
XOR2_X1 U1015 ( .A(KEYINPUT37), .B(G224), .Z(n1284) );
NAND2_X1 U1016 ( .A1(KEYINPUT27), .A2(n1190), .ZN(n1283) );
INV_X1 U1017 ( .A(G125), .ZN(n1190) );
XNOR2_X1 U1018 ( .A(KEYINPUT47), .B(KEYINPUT0), .ZN(n1281) );
NOR2_X1 U1019 ( .A1(n1225), .A2(n1229), .ZN(n1033) );
INV_X1 U1020 ( .A(n1211), .ZN(n1229) );
XOR2_X1 U1021 ( .A(n1055), .B(n1285), .Z(n1211) );
NOR2_X1 U1022 ( .A1(G478), .A2(KEYINPUT16), .ZN(n1285) );
NOR2_X1 U1023 ( .A1(n1117), .A2(G902), .ZN(n1055) );
INV_X1 U1024 ( .A(n1115), .ZN(n1117) );
XNOR2_X1 U1025 ( .A(n1286), .B(n1287), .ZN(n1115) );
XNOR2_X1 U1026 ( .A(n1269), .B(n1288), .ZN(n1287) );
XOR2_X1 U1027 ( .A(n1289), .B(n1290), .Z(n1288) );
NOR3_X1 U1028 ( .A1(KEYINPUT29), .A2(n1291), .A3(n1292), .ZN(n1290) );
NOR2_X1 U1029 ( .A1(n1194), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U1030 ( .A(G128), .B(KEYINPUT2), .ZN(n1293) );
NOR2_X1 U1031 ( .A1(G143), .A2(n1294), .ZN(n1291) );
XNOR2_X1 U1032 ( .A(KEYINPUT30), .B(n1084), .ZN(n1294) );
INV_X1 U1033 ( .A(G128), .ZN(n1084) );
NAND3_X1 U1034 ( .A1(n1246), .A2(G234), .A3(G217), .ZN(n1289) );
XOR2_X1 U1035 ( .A(G134), .B(KEYINPUT48), .Z(n1269) );
XNOR2_X1 U1036 ( .A(G107), .B(n1295), .ZN(n1286) );
XNOR2_X1 U1037 ( .A(n1103), .B(G116), .ZN(n1295) );
XNOR2_X1 U1038 ( .A(n1296), .B(G475), .ZN(n1225) );
NAND2_X1 U1039 ( .A1(n1120), .A2(n1156), .ZN(n1296) );
INV_X1 U1040 ( .A(G902), .ZN(n1156) );
XNOR2_X1 U1041 ( .A(n1297), .B(n1298), .ZN(n1120) );
XNOR2_X1 U1042 ( .A(n1255), .B(n1078), .ZN(n1298) );
INV_X1 U1043 ( .A(n1081), .ZN(n1078) );
XOR2_X1 U1044 ( .A(G125), .B(G140), .Z(n1081) );
XNOR2_X1 U1045 ( .A(G146), .B(n1194), .ZN(n1255) );
INV_X1 U1046 ( .A(G143), .ZN(n1194) );
XOR2_X1 U1047 ( .A(n1299), .B(n1300), .Z(n1297) );
XNOR2_X1 U1048 ( .A(G131), .B(n1301), .ZN(n1300) );
NAND3_X1 U1049 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1301) );
NAND2_X1 U1050 ( .A1(n1305), .A2(n1125), .ZN(n1304) );
INV_X1 U1051 ( .A(G104), .ZN(n1125) );
NAND2_X1 U1052 ( .A1(n1306), .A2(n1307), .ZN(n1303) );
INV_X1 U1053 ( .A(KEYINPUT53), .ZN(n1307) );
NAND2_X1 U1054 ( .A1(n1308), .A2(G104), .ZN(n1306) );
XNOR2_X1 U1055 ( .A(KEYINPUT56), .B(n1309), .ZN(n1308) );
NAND2_X1 U1056 ( .A1(KEYINPUT53), .A2(n1310), .ZN(n1302) );
NAND2_X1 U1057 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
OR2_X1 U1058 ( .A1(n1309), .A2(KEYINPUT56), .ZN(n1312) );
NAND3_X1 U1059 ( .A1(G104), .A2(n1309), .A3(KEYINPUT56), .ZN(n1311) );
INV_X1 U1060 ( .A(n1305), .ZN(n1309) );
XOR2_X1 U1061 ( .A(G113), .B(n1103), .Z(n1305) );
INV_X1 U1062 ( .A(G122), .ZN(n1103) );
NAND4_X1 U1063 ( .A1(KEYINPUT6), .A2(G214), .A3(n1246), .A4(n1252), .ZN(n1299) );
INV_X1 U1064 ( .A(G237), .ZN(n1252) );
XNOR2_X1 U1065 ( .A(G953), .B(KEYINPUT34), .ZN(n1246) );
endmodule


