//Key = 1111111011011100011101101011010010101011000110110111001000011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;

XOR2_X1 U690 ( .A(G107), .B(n950), .Z(G9) );
NOR2_X1 U691 ( .A1(n951), .A2(n952), .ZN(G75) );
NOR4_X1 U692 ( .A1(n953), .A2(n954), .A3(n955), .A4(n956), .ZN(n952) );
NOR3_X1 U693 ( .A1(n957), .A2(n958), .A3(n959), .ZN(n956) );
NOR2_X1 U694 ( .A1(n960), .A2(n961), .ZN(n958) );
NOR2_X1 U695 ( .A1(n962), .A2(n963), .ZN(n961) );
NOR2_X1 U696 ( .A1(n964), .A2(n965), .ZN(n962) );
NOR2_X1 U697 ( .A1(n966), .A2(n967), .ZN(n965) );
NOR2_X1 U698 ( .A1(n968), .A2(n969), .ZN(n966) );
NOR2_X1 U699 ( .A1(n970), .A2(n971), .ZN(n968) );
NOR2_X1 U700 ( .A1(n972), .A2(n973), .ZN(n964) );
NOR2_X1 U701 ( .A1(n974), .A2(n975), .ZN(n972) );
NOR2_X1 U702 ( .A1(n976), .A2(n977), .ZN(n974) );
NOR3_X1 U703 ( .A1(n973), .A2(n978), .A3(n967), .ZN(n960) );
NOR2_X1 U704 ( .A1(n979), .A2(n980), .ZN(n978) );
NOR2_X1 U705 ( .A1(n981), .A2(n973), .ZN(n954) );
NOR2_X1 U706 ( .A1(n982), .A2(n983), .ZN(n981) );
XOR2_X1 U707 ( .A(n984), .B(KEYINPUT3), .Z(n983) );
NAND4_X1 U708 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n984) );
NOR2_X1 U709 ( .A1(n957), .A2(n989), .ZN(n988) );
XOR2_X1 U710 ( .A(KEYINPUT59), .B(n990), .Z(n989) );
NOR4_X1 U711 ( .A1(n967), .A2(n963), .A3(n991), .A4(n957), .ZN(n982) );
NAND2_X1 U712 ( .A1(n992), .A2(n993), .ZN(n953) );
NOR3_X1 U713 ( .A1(n994), .A2(G952), .A3(n955), .ZN(n951) );
AND4_X1 U714 ( .A1(n995), .A2(n996), .A3(n997), .A4(n998), .ZN(n955) );
NOR4_X1 U715 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(n998) );
XOR2_X1 U716 ( .A(KEYINPUT40), .B(n1003), .Z(n1002) );
NAND2_X1 U717 ( .A1(n1004), .A2(n1005), .ZN(n1000) );
XOR2_X1 U718 ( .A(n1006), .B(n1007), .Z(n1005) );
XOR2_X1 U719 ( .A(n1008), .B(KEYINPUT13), .Z(n1007) );
XNOR2_X1 U720 ( .A(n1009), .B(n1010), .ZN(n1004) );
NAND2_X1 U721 ( .A1(KEYINPUT36), .A2(n1011), .ZN(n1010) );
XOR2_X1 U722 ( .A(n1012), .B(n1013), .Z(n999) );
XOR2_X1 U723 ( .A(n1014), .B(KEYINPUT44), .Z(n1012) );
NOR3_X1 U724 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n997) );
NAND2_X1 U725 ( .A1(n1018), .A2(n1019), .ZN(n995) );
XOR2_X1 U726 ( .A(KEYINPUT45), .B(n1020), .Z(n1018) );
INV_X1 U727 ( .A(n992), .ZN(n994) );
XOR2_X1 U728 ( .A(n1021), .B(n1022), .Z(G72) );
NOR2_X1 U729 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
AND2_X1 U730 ( .A1(G227), .A2(G900), .ZN(n1023) );
NAND2_X1 U731 ( .A1(n1025), .A2(n1026), .ZN(n1021) );
NAND2_X1 U732 ( .A1(n1027), .A2(n1024), .ZN(n1026) );
XOR2_X1 U733 ( .A(n1028), .B(n1029), .Z(n1027) );
NOR2_X1 U734 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
OR3_X1 U735 ( .A1(n1032), .A2(n1029), .A3(n1024), .ZN(n1025) );
XNOR2_X1 U736 ( .A(n1033), .B(n1034), .ZN(n1029) );
XOR2_X1 U737 ( .A(G131), .B(n1035), .Z(n1034) );
XOR2_X1 U738 ( .A(KEYINPUT22), .B(G137), .Z(n1035) );
XOR2_X1 U739 ( .A(n1036), .B(n1037), .Z(n1033) );
XOR2_X1 U740 ( .A(n1038), .B(n1039), .Z(n1036) );
NAND2_X1 U741 ( .A1(KEYINPUT47), .A2(n1040), .ZN(n1038) );
XOR2_X1 U742 ( .A(n1041), .B(n1042), .Z(G69) );
NOR2_X1 U743 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U744 ( .A1(n1024), .A2(n1045), .ZN(n1044) );
XOR2_X1 U745 ( .A(n1046), .B(KEYINPUT27), .Z(n1045) );
NAND2_X1 U746 ( .A1(G898), .A2(G224), .ZN(n1046) );
NOR2_X1 U747 ( .A1(G953), .A2(n1047), .ZN(n1043) );
NAND3_X1 U748 ( .A1(n1048), .A2(n1049), .A3(KEYINPUT49), .ZN(n1041) );
NAND2_X1 U749 ( .A1(G953), .A2(n1050), .ZN(n1049) );
XNOR2_X1 U750 ( .A(n1051), .B(n1052), .ZN(n1048) );
NOR2_X1 U751 ( .A1(KEYINPUT15), .A2(n1053), .ZN(n1051) );
NOR2_X1 U752 ( .A1(n1054), .A2(n1055), .ZN(G66) );
NOR3_X1 U753 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NOR3_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
AND2_X1 U755 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND3_X1 U756 ( .A1(n1062), .A2(n1063), .A3(KEYINPUT54), .ZN(n1059) );
INV_X1 U757 ( .A(n1006), .ZN(n1062) );
NOR2_X1 U758 ( .A1(n1054), .A2(n1064), .ZN(G63) );
XNOR2_X1 U759 ( .A(n1065), .B(n1066), .ZN(n1064) );
NAND3_X1 U760 ( .A1(n1067), .A2(G478), .A3(KEYINPUT60), .ZN(n1065) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1068), .ZN(G60) );
XOR2_X1 U762 ( .A(n1069), .B(n1070), .Z(n1068) );
NAND2_X1 U763 ( .A1(n1067), .A2(G475), .ZN(n1069) );
XNOR2_X1 U764 ( .A(G104), .B(n1071), .ZN(G6) );
NOR2_X1 U765 ( .A1(n1054), .A2(n1072), .ZN(G57) );
NOR3_X1 U766 ( .A1(n1009), .A2(n1073), .A3(n1074), .ZN(n1072) );
AND3_X1 U767 ( .A1(n1075), .A2(G472), .A3(n1067), .ZN(n1074) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1075), .ZN(n1073) );
NOR2_X1 U769 ( .A1(n993), .A2(n1011), .ZN(n1076) );
INV_X1 U770 ( .A(G472), .ZN(n1011) );
NOR2_X1 U771 ( .A1(n1054), .A2(n1077), .ZN(G54) );
XOR2_X1 U772 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U773 ( .A(n1080), .B(n1081), .Z(n1078) );
NOR3_X1 U774 ( .A1(n1082), .A2(n993), .A3(n1083), .ZN(n1081) );
XOR2_X1 U775 ( .A(KEYINPUT61), .B(G902), .Z(n1082) );
NAND2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1080) );
OR2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U778 ( .A(n1088), .B(KEYINPUT62), .Z(n1084) );
NAND2_X1 U779 ( .A1(n1086), .A2(n1087), .ZN(n1088) );
XNOR2_X1 U780 ( .A(n1089), .B(n1090), .ZN(n1086) );
XNOR2_X1 U781 ( .A(KEYINPUT63), .B(n1091), .ZN(n1089) );
NOR2_X1 U782 ( .A1(n1054), .A2(n1092), .ZN(G51) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U784 ( .A1(KEYINPUT48), .A2(n1095), .ZN(n1094) );
XNOR2_X1 U785 ( .A(n1096), .B(n1097), .ZN(n1095) );
XOR2_X1 U786 ( .A(KEYINPUT38), .B(n1098), .Z(n1097) );
NAND2_X1 U787 ( .A1(n1067), .A2(n1013), .ZN(n1093) );
INV_X1 U788 ( .A(n1099), .ZN(n1013) );
NOR2_X1 U789 ( .A1(n1061), .A2(n993), .ZN(n1067) );
INV_X1 U790 ( .A(n1063), .ZN(n993) );
NAND3_X1 U791 ( .A1(n1047), .A2(n1100), .A3(n1101), .ZN(n1063) );
XNOR2_X1 U792 ( .A(n1030), .B(KEYINPUT14), .ZN(n1101) );
INV_X1 U793 ( .A(n1031), .ZN(n1100) );
NAND4_X1 U794 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1031) );
NOR4_X1 U795 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1105) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1104) );
XOR2_X1 U797 ( .A(n973), .B(KEYINPUT26), .Z(n1110) );
INV_X1 U798 ( .A(n1112), .ZN(n973) );
NAND2_X1 U799 ( .A1(n969), .A2(n1113), .ZN(n1102) );
XOR2_X1 U800 ( .A(KEYINPUT20), .B(n1114), .Z(n1113) );
AND4_X1 U801 ( .A1(n1071), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1047) );
NOR4_X1 U802 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n950), .ZN(n1117) );
AND3_X1 U803 ( .A1(n1121), .A2(n1122), .A3(n979), .ZN(n950) );
NAND2_X1 U804 ( .A1(n990), .A2(n1123), .ZN(n1116) );
NAND2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND3_X1 U806 ( .A1(n1126), .A2(n986), .A3(n1127), .ZN(n1125) );
NAND2_X1 U807 ( .A1(n1128), .A2(n1122), .ZN(n1124) );
NAND3_X1 U808 ( .A1(n1121), .A2(n1122), .A3(n980), .ZN(n1071) );
INV_X1 U809 ( .A(n1129), .ZN(n1122) );
NOR2_X1 U810 ( .A1(n1024), .A2(G952), .ZN(n1054) );
XNOR2_X1 U811 ( .A(G146), .B(n1130), .ZN(G48) );
NAND2_X1 U812 ( .A1(n1114), .A2(n969), .ZN(n1130) );
AND2_X1 U813 ( .A1(n1131), .A2(n980), .ZN(n1114) );
XOR2_X1 U814 ( .A(n1132), .B(n1103), .Z(G45) );
NAND4_X1 U815 ( .A1(n969), .A2(n975), .A3(n1128), .A4(n1133), .ZN(n1103) );
AND3_X1 U816 ( .A1(n1001), .A2(n1134), .A3(n1135), .ZN(n1133) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(G42) );
NAND2_X1 U818 ( .A1(n1111), .A2(n1112), .ZN(n1137) );
AND2_X1 U819 ( .A1(n1138), .A2(n975), .ZN(n1111) );
NAND2_X1 U820 ( .A1(KEYINPUT21), .A2(G140), .ZN(n1136) );
XOR2_X1 U821 ( .A(G137), .B(n1108), .Z(G39) );
AND3_X1 U822 ( .A1(n1112), .A2(n990), .A3(n1131), .ZN(n1108) );
XOR2_X1 U823 ( .A(G134), .B(n1107), .Z(G36) );
AND2_X1 U824 ( .A1(n1139), .A2(n979), .ZN(n1107) );
XOR2_X1 U825 ( .A(G131), .B(n1106), .Z(G33) );
AND2_X1 U826 ( .A1(n1139), .A2(n980), .ZN(n1106) );
AND4_X1 U827 ( .A1(n1112), .A2(n1128), .A3(n975), .A4(n1135), .ZN(n1139) );
NOR2_X1 U828 ( .A1(n970), .A2(n1015), .ZN(n1112) );
INV_X1 U829 ( .A(n971), .ZN(n1015) );
XOR2_X1 U830 ( .A(G128), .B(n1030), .Z(G30) );
AND3_X1 U831 ( .A1(n979), .A2(n969), .A3(n1131), .ZN(n1030) );
AND4_X1 U832 ( .A1(n975), .A2(n1126), .A3(n986), .A4(n1135), .ZN(n1131) );
XOR2_X1 U833 ( .A(G101), .B(n1140), .Z(G3) );
NOR3_X1 U834 ( .A1(n963), .A2(n1141), .A3(n1129), .ZN(n1140) );
XOR2_X1 U835 ( .A(n991), .B(KEYINPUT30), .Z(n1141) );
NAND2_X1 U836 ( .A1(n1142), .A2(n1143), .ZN(G27) );
NAND2_X1 U837 ( .A1(G125), .A2(n1144), .ZN(n1143) );
XOR2_X1 U838 ( .A(n1145), .B(KEYINPUT35), .Z(n1142) );
NAND2_X1 U839 ( .A1(n1109), .A2(n1146), .ZN(n1145) );
INV_X1 U840 ( .A(n1144), .ZN(n1109) );
NAND3_X1 U841 ( .A1(n969), .A2(n985), .A3(n1138), .ZN(n1144) );
AND4_X1 U842 ( .A1(n987), .A2(n980), .A3(n986), .A4(n1135), .ZN(n1138) );
NAND2_X1 U843 ( .A1(n957), .A2(n1147), .ZN(n1135) );
NAND4_X1 U844 ( .A1(G953), .A2(G902), .A3(n1148), .A4(n1032), .ZN(n1147) );
INV_X1 U845 ( .A(G900), .ZN(n1032) );
INV_X1 U846 ( .A(n1149), .ZN(n986) );
XOR2_X1 U847 ( .A(n1150), .B(n1115), .Z(G24) );
NAND4_X1 U848 ( .A1(n1127), .A2(n1121), .A3(n1001), .A4(n1134), .ZN(n1115) );
INV_X1 U849 ( .A(n959), .ZN(n1121) );
NAND2_X1 U850 ( .A1(n1149), .A2(n987), .ZN(n959) );
XNOR2_X1 U851 ( .A(G119), .B(n1151), .ZN(G21) );
NAND4_X1 U852 ( .A1(n990), .A2(n985), .A3(n1152), .A4(n1153), .ZN(n1151) );
NOR3_X1 U853 ( .A1(n987), .A2(n1154), .A3(n1149), .ZN(n1153) );
INV_X1 U854 ( .A(n1126), .ZN(n987) );
XOR2_X1 U855 ( .A(n1155), .B(KEYINPUT6), .Z(n1152) );
XOR2_X1 U856 ( .A(G116), .B(n1120), .Z(G18) );
AND3_X1 U857 ( .A1(n1128), .A2(n979), .A3(n1127), .ZN(n1120) );
AND2_X1 U858 ( .A1(n1156), .A2(n1134), .ZN(n979) );
XOR2_X1 U859 ( .A(n1157), .B(n1119), .Z(G15) );
AND3_X1 U860 ( .A1(n1128), .A2(n980), .A3(n1127), .ZN(n1119) );
NOR3_X1 U861 ( .A1(n967), .A2(n1154), .A3(n1155), .ZN(n1127) );
INV_X1 U862 ( .A(n1158), .ZN(n1154) );
INV_X1 U863 ( .A(n985), .ZN(n967) );
NAND2_X1 U864 ( .A1(n1159), .A2(n1160), .ZN(n985) );
OR3_X1 U865 ( .A1(n977), .A2(n1003), .A3(KEYINPUT33), .ZN(n1160) );
INV_X1 U866 ( .A(n1161), .ZN(n977) );
NAND2_X1 U867 ( .A1(KEYINPUT33), .A2(n975), .ZN(n1159) );
NOR2_X1 U868 ( .A1(n1134), .A2(n1156), .ZN(n980) );
INV_X1 U869 ( .A(n991), .ZN(n1128) );
NAND2_X1 U870 ( .A1(n1149), .A2(n1126), .ZN(n991) );
XNOR2_X1 U871 ( .A(G113), .B(KEYINPUT5), .ZN(n1157) );
XNOR2_X1 U872 ( .A(G110), .B(n1162), .ZN(G12) );
NOR2_X1 U873 ( .A1(n1118), .A2(KEYINPUT56), .ZN(n1162) );
NOR4_X1 U874 ( .A1(n963), .A2(n1129), .A3(n1126), .A4(n1149), .ZN(n1118) );
XOR2_X1 U875 ( .A(n1163), .B(n1164), .Z(n1149) );
XOR2_X1 U876 ( .A(KEYINPUT17), .B(n1056), .Z(n1164) );
INV_X1 U877 ( .A(n1008), .ZN(n1056) );
NAND2_X1 U878 ( .A1(n1060), .A2(n1061), .ZN(n1008) );
XOR2_X1 U879 ( .A(n1165), .B(n1166), .Z(n1060) );
XOR2_X1 U880 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U881 ( .A(G128), .B(G119), .Z(n1168) );
XOR2_X1 U882 ( .A(KEYINPUT9), .B(G146), .Z(n1167) );
XOR2_X1 U883 ( .A(n1169), .B(n1037), .Z(n1165) );
XOR2_X1 U884 ( .A(n1170), .B(G110), .Z(n1169) );
NAND2_X1 U885 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND4_X1 U886 ( .A1(G221), .A2(G137), .A3(G234), .A4(n1024), .ZN(n1172) );
NAND2_X1 U887 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NAND3_X1 U888 ( .A1(G234), .A2(n1024), .A3(G221), .ZN(n1174) );
XOR2_X1 U889 ( .A(KEYINPUT4), .B(G137), .Z(n1173) );
NAND2_X1 U890 ( .A1(KEYINPUT11), .A2(n1006), .ZN(n1163) );
NAND2_X1 U891 ( .A1(G217), .A2(n1175), .ZN(n1006) );
XOR2_X1 U892 ( .A(n1009), .B(G472), .Z(n1126) );
NOR2_X1 U893 ( .A1(n1075), .A2(G902), .ZN(n1009) );
XNOR2_X1 U894 ( .A(n1176), .B(n1177), .ZN(n1075) );
XOR2_X1 U895 ( .A(n1178), .B(n1090), .Z(n1177) );
XOR2_X1 U896 ( .A(G101), .B(n1039), .Z(n1090) );
XOR2_X1 U897 ( .A(n1179), .B(n1180), .Z(n1176) );
INV_X1 U898 ( .A(n1181), .ZN(n1180) );
NAND2_X1 U899 ( .A1(G210), .A2(n1182), .ZN(n1179) );
NAND3_X1 U900 ( .A1(n975), .A2(n1158), .A3(n969), .ZN(n1129) );
INV_X1 U901 ( .A(n1155), .ZN(n969) );
NAND2_X1 U902 ( .A1(n970), .A2(n971), .ZN(n1155) );
NAND2_X1 U903 ( .A1(G214), .A2(n1183), .ZN(n971) );
XNOR2_X1 U904 ( .A(n1184), .B(n1014), .ZN(n970) );
NAND2_X1 U905 ( .A1(n1185), .A2(n1061), .ZN(n1014) );
XOR2_X1 U906 ( .A(n1186), .B(n1098), .Z(n1185) );
XOR2_X1 U907 ( .A(n1187), .B(n1053), .Z(n1098) );
XOR2_X1 U908 ( .A(n1188), .B(n1178), .Z(n1053) );
XNOR2_X1 U909 ( .A(n1189), .B(n1190), .ZN(n1178) );
XOR2_X1 U910 ( .A(KEYINPUT18), .B(G119), .Z(n1190) );
XNOR2_X1 U911 ( .A(G113), .B(G116), .ZN(n1189) );
XOR2_X1 U912 ( .A(n1191), .B(G101), .Z(n1188) );
NAND2_X1 U913 ( .A1(KEYINPUT29), .A2(n1192), .ZN(n1191) );
NAND2_X1 U914 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U915 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XNOR2_X1 U916 ( .A(n1197), .B(KEYINPUT53), .ZN(n1195) );
XOR2_X1 U917 ( .A(n1198), .B(KEYINPUT52), .Z(n1193) );
NAND2_X1 U918 ( .A1(n1199), .A2(n1197), .ZN(n1198) );
XOR2_X1 U919 ( .A(G104), .B(KEYINPUT8), .Z(n1197) );
XOR2_X1 U920 ( .A(n1196), .B(KEYINPUT32), .Z(n1199) );
INV_X1 U921 ( .A(G107), .ZN(n1196) );
NAND2_X1 U922 ( .A1(KEYINPUT12), .A2(n1052), .ZN(n1187) );
XOR2_X1 U923 ( .A(G110), .B(n1150), .Z(n1052) );
INV_X1 U924 ( .A(G122), .ZN(n1150) );
NOR2_X1 U925 ( .A1(KEYINPUT16), .A2(n1096), .ZN(n1186) );
XOR2_X1 U926 ( .A(n1200), .B(n1039), .Z(n1096) );
XOR2_X1 U927 ( .A(n1146), .B(n1201), .Z(n1200) );
AND2_X1 U928 ( .A1(n1024), .A2(G224), .ZN(n1201) );
INV_X1 U929 ( .A(G125), .ZN(n1146) );
NAND2_X1 U930 ( .A1(n1202), .A2(KEYINPUT1), .ZN(n1184) );
XOR2_X1 U931 ( .A(n1099), .B(KEYINPUT55), .Z(n1202) );
NAND2_X1 U932 ( .A1(G210), .A2(n1183), .ZN(n1099) );
NAND2_X1 U933 ( .A1(n1203), .A2(n1061), .ZN(n1183) );
INV_X1 U934 ( .A(G237), .ZN(n1203) );
NAND2_X1 U935 ( .A1(n957), .A2(n1204), .ZN(n1158) );
NAND4_X1 U936 ( .A1(G953), .A2(G902), .A3(n1148), .A4(n1050), .ZN(n1204) );
INV_X1 U937 ( .A(G898), .ZN(n1050) );
NAND3_X1 U938 ( .A1(n992), .A2(n1148), .A3(G952), .ZN(n957) );
NAND2_X1 U939 ( .A1(G237), .A2(G234), .ZN(n1148) );
XOR2_X1 U940 ( .A(n1024), .B(KEYINPUT10), .Z(n992) );
NOR2_X1 U941 ( .A1(n1003), .A2(n1161), .ZN(n975) );
NOR2_X1 U942 ( .A1(n1205), .A2(n1017), .ZN(n1161) );
NOR2_X1 U943 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
AND2_X1 U944 ( .A1(n1020), .A2(n1019), .ZN(n1205) );
NAND3_X1 U945 ( .A1(n1206), .A2(n1207), .A3(n1061), .ZN(n1019) );
NAND2_X1 U946 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
INV_X1 U947 ( .A(KEYINPUT37), .ZN(n1209) );
XOR2_X1 U948 ( .A(n1210), .B(n1211), .Z(n1208) );
NAND3_X1 U949 ( .A1(n1211), .A2(n1210), .A3(KEYINPUT37), .ZN(n1206) );
XNOR2_X1 U950 ( .A(n1079), .B(KEYINPUT2), .ZN(n1210) );
XNOR2_X1 U951 ( .A(n1212), .B(n1213), .ZN(n1079) );
XOR2_X1 U952 ( .A(G140), .B(G110), .Z(n1213) );
NAND2_X1 U953 ( .A1(G227), .A2(n1024), .ZN(n1212) );
XOR2_X1 U954 ( .A(n1214), .B(n1215), .Z(n1211) );
XOR2_X1 U955 ( .A(G101), .B(n1216), .Z(n1215) );
NOR2_X1 U956 ( .A1(KEYINPUT57), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U957 ( .A(n1039), .B(KEYINPUT63), .ZN(n1217) );
XOR2_X1 U958 ( .A(G146), .B(n1218), .Z(n1039) );
XNOR2_X1 U959 ( .A(n1091), .B(n1087), .ZN(n1214) );
XNOR2_X1 U960 ( .A(n1181), .B(KEYINPUT31), .ZN(n1087) );
XOR2_X1 U961 ( .A(n1219), .B(n1220), .Z(n1181) );
NOR2_X1 U962 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XOR2_X1 U963 ( .A(n1223), .B(KEYINPUT19), .Z(n1222) );
NAND2_X1 U964 ( .A1(G137), .A2(n1040), .ZN(n1223) );
NOR2_X1 U965 ( .A1(G137), .A2(n1040), .ZN(n1221) );
XOR2_X1 U966 ( .A(G134), .B(KEYINPUT34), .Z(n1040) );
NAND2_X1 U967 ( .A1(KEYINPUT43), .A2(n1224), .ZN(n1219) );
INV_X1 U968 ( .A(G131), .ZN(n1224) );
XOR2_X1 U969 ( .A(G104), .B(G107), .Z(n1091) );
XNOR2_X1 U970 ( .A(n1083), .B(KEYINPUT28), .ZN(n1020) );
INV_X1 U971 ( .A(G469), .ZN(n1083) );
INV_X1 U972 ( .A(n976), .ZN(n1003) );
NAND2_X1 U973 ( .A1(G221), .A2(n1175), .ZN(n976) );
NAND2_X1 U974 ( .A1(G234), .A2(n1061), .ZN(n1175) );
INV_X1 U975 ( .A(n990), .ZN(n963) );
NOR2_X1 U976 ( .A1(n1134), .A2(n1001), .ZN(n990) );
INV_X1 U977 ( .A(n1156), .ZN(n1001) );
XOR2_X1 U978 ( .A(n1225), .B(G475), .Z(n1156) );
NAND2_X1 U979 ( .A1(n1070), .A2(n1061), .ZN(n1225) );
INV_X1 U980 ( .A(G902), .ZN(n1061) );
XNOR2_X1 U981 ( .A(n1226), .B(n1227), .ZN(n1070) );
XOR2_X1 U982 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U983 ( .A(G122), .B(G113), .Z(n1229) );
NOR2_X1 U984 ( .A1(n1230), .A2(n1231), .ZN(n1228) );
XOR2_X1 U985 ( .A(KEYINPUT25), .B(n1232), .Z(n1231) );
NOR2_X1 U986 ( .A1(G131), .A2(n1233), .ZN(n1232) );
AND2_X1 U987 ( .A1(n1233), .A2(G131), .ZN(n1230) );
NAND3_X1 U988 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NAND2_X1 U989 ( .A1(n1132), .A2(n1237), .ZN(n1236) );
OR3_X1 U990 ( .A1(n1237), .A2(n1132), .A3(n1238), .ZN(n1235) );
INV_X1 U991 ( .A(KEYINPUT39), .ZN(n1237) );
NAND2_X1 U992 ( .A1(n1239), .A2(n1238), .ZN(n1234) );
NAND2_X1 U993 ( .A1(G214), .A2(n1182), .ZN(n1238) );
AND2_X1 U994 ( .A1(n1240), .A2(n1024), .ZN(n1182) );
XOR2_X1 U995 ( .A(KEYINPUT0), .B(G237), .Z(n1240) );
NAND2_X1 U996 ( .A1(n1241), .A2(KEYINPUT39), .ZN(n1239) );
XOR2_X1 U997 ( .A(n1132), .B(KEYINPUT24), .Z(n1241) );
INV_X1 U998 ( .A(G143), .ZN(n1132) );
XOR2_X1 U999 ( .A(n1242), .B(n1243), .Z(n1226) );
XNOR2_X1 U1000 ( .A(n1244), .B(n1245), .ZN(n1243) );
NOR2_X1 U1001 ( .A1(G104), .A2(KEYINPUT41), .ZN(n1245) );
NAND2_X1 U1002 ( .A1(KEYINPUT46), .A2(G146), .ZN(n1244) );
INV_X1 U1003 ( .A(n1037), .ZN(n1242) );
XOR2_X1 U1004 ( .A(G140), .B(G125), .Z(n1037) );
NAND2_X1 U1005 ( .A1(n1246), .A2(n996), .ZN(n1134) );
NAND2_X1 U1006 ( .A1(G478), .A2(n1247), .ZN(n996) );
OR2_X1 U1007 ( .A1(n1066), .A2(G902), .ZN(n1247) );
XNOR2_X1 U1008 ( .A(n1016), .B(KEYINPUT42), .ZN(n1246) );
NOR3_X1 U1009 ( .A1(G478), .A2(G902), .A3(n1066), .ZN(n1016) );
XOR2_X1 U1010 ( .A(n1248), .B(n1249), .Z(n1066) );
AND3_X1 U1011 ( .A1(G234), .A2(n1024), .A3(G217), .ZN(n1249) );
INV_X1 U1012 ( .A(G953), .ZN(n1024) );
NAND3_X1 U1013 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1248) );
NAND2_X1 U1014 ( .A1(KEYINPUT23), .A2(n1253), .ZN(n1252) );
NAND3_X1 U1015 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1251) );
INV_X1 U1016 ( .A(KEYINPUT23), .ZN(n1255) );
OR2_X1 U1017 ( .A1(n1256), .A2(n1254), .ZN(n1250) );
NOR2_X1 U1018 ( .A1(KEYINPUT58), .A2(n1253), .ZN(n1254) );
XOR2_X1 U1019 ( .A(G134), .B(n1218), .Z(n1253) );
XOR2_X1 U1020 ( .A(G128), .B(G143), .Z(n1218) );
NAND3_X1 U1021 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
NAND2_X1 U1022 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
OR3_X1 U1023 ( .A1(n1261), .A2(n1260), .A3(n1262), .ZN(n1258) );
INV_X1 U1024 ( .A(KEYINPUT50), .ZN(n1261) );
NAND2_X1 U1025 ( .A1(n1262), .A2(n1263), .ZN(n1257) );
NAND2_X1 U1026 ( .A1(KEYINPUT50), .A2(n1264), .ZN(n1263) );
XNOR2_X1 U1027 ( .A(KEYINPUT7), .B(n1260), .ZN(n1264) );
XNOR2_X1 U1028 ( .A(G107), .B(KEYINPUT51), .ZN(n1260) );
XOR2_X1 U1029 ( .A(G116), .B(G122), .Z(n1262) );
endmodule


