//Key = 1111111101010011101100111010000101011010111010100011001000110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371;

NAND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(G9) );
NAND2_X1 U758 ( .A1(G107), .A2(n1050), .ZN(n1049) );
XOR2_X1 U759 ( .A(KEYINPUT54), .B(n1051), .Z(n1048) );
NOR2_X1 U760 ( .A1(G107), .A2(n1050), .ZN(n1051) );
NOR2_X1 U761 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
NOR4_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1056) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NAND4_X1 U765 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XNOR2_X1 U767 ( .A(n1070), .B(KEYINPUT19), .ZN(n1068) );
NAND2_X1 U768 ( .A1(KEYINPUT7), .A2(n1071), .ZN(n1066) );
NAND2_X1 U769 ( .A1(n1070), .A2(n1072), .ZN(n1065) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1058) );
NOR2_X1 U772 ( .A1(KEYINPUT7), .A2(n1077), .ZN(n1075) );
INV_X1 U773 ( .A(n1071), .ZN(n1077) );
NAND3_X1 U774 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1054) );
NAND4_X1 U775 ( .A1(n1070), .A2(n1074), .A3(n1081), .A4(n1076), .ZN(n1080) );
NAND4_X1 U776 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
NAND2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U779 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
INV_X1 U780 ( .A(KEYINPUT56), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NAND3_X1 U782 ( .A1(KEYINPUT56), .A2(n1090), .A3(n1060), .ZN(n1084) );
OR3_X1 U783 ( .A1(n1094), .A2(n1061), .A3(n1095), .ZN(n1082) );
NOR3_X1 U784 ( .A1(n1096), .A2(G953), .A3(G952), .ZN(n1052) );
INV_X1 U785 ( .A(n1078), .ZN(n1096) );
NAND4_X1 U786 ( .A1(n1097), .A2(n1086), .A3(n1098), .A4(n1099), .ZN(n1078) );
NOR4_X1 U787 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
XOR2_X1 U788 ( .A(n1104), .B(n1105), .Z(n1098) );
XOR2_X1 U789 ( .A(n1106), .B(n1107), .Z(G72) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U792 ( .A(n1112), .B(n1113), .Z(n1111) );
XNOR2_X1 U793 ( .A(n1114), .B(n1115), .ZN(n1113) );
XNOR2_X1 U794 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U795 ( .A1(KEYINPUT46), .A2(G134), .ZN(n1116) );
XNOR2_X1 U796 ( .A(n1118), .B(n1119), .ZN(n1112) );
NOR2_X1 U797 ( .A1(G900), .A2(n1079), .ZN(n1110) );
NAND2_X1 U798 ( .A1(n1120), .A2(n1055), .ZN(n1108) );
XNOR2_X1 U799 ( .A(G953), .B(KEYINPUT47), .ZN(n1120) );
NAND2_X1 U800 ( .A1(G953), .A2(n1121), .ZN(n1106) );
NAND2_X1 U801 ( .A1(G900), .A2(G227), .ZN(n1121) );
XOR2_X1 U802 ( .A(n1122), .B(n1123), .Z(G69) );
NAND2_X1 U803 ( .A1(G953), .A2(n1124), .ZN(n1123) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1124) );
NAND2_X1 U805 ( .A1(KEYINPUT5), .A2(n1125), .ZN(n1122) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U807 ( .A1(n1079), .A2(n1057), .ZN(n1127) );
NAND3_X1 U808 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1126) );
XOR2_X1 U809 ( .A(KEYINPUT63), .B(n1131), .Z(n1130) );
NOR2_X1 U810 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
OR3_X1 U812 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1129) );
AND2_X1 U813 ( .A1(KEYINPUT3), .A2(n1137), .ZN(n1135) );
NOR3_X1 U814 ( .A1(n1138), .A2(KEYINPUT3), .A3(n1139), .ZN(n1134) );
NAND2_X1 U815 ( .A1(G953), .A2(n1140), .ZN(n1128) );
NOR3_X1 U816 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(G66) );
AND2_X1 U817 ( .A1(KEYINPUT14), .A2(n1144), .ZN(n1143) );
NOR3_X1 U818 ( .A1(KEYINPUT14), .A2(G953), .A3(G952), .ZN(n1142) );
XOR2_X1 U819 ( .A(n1145), .B(n1146), .Z(n1141) );
NAND2_X1 U820 ( .A1(n1147), .A2(n1105), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1148), .ZN(G63) );
NOR2_X1 U822 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U823 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U824 ( .A1(n1153), .A2(n1154), .ZN(n1149) );
XOR2_X1 U825 ( .A(KEYINPUT38), .B(n1151), .Z(n1154) );
AND2_X1 U826 ( .A1(n1147), .A2(G478), .ZN(n1151) );
XNOR2_X1 U827 ( .A(n1152), .B(KEYINPUT34), .ZN(n1153) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(G60) );
XOR2_X1 U829 ( .A(KEYINPUT39), .B(n1144), .Z(n1156) );
XNOR2_X1 U830 ( .A(n1157), .B(n1158), .ZN(n1155) );
NAND2_X1 U831 ( .A1(n1147), .A2(G475), .ZN(n1157) );
XNOR2_X1 U832 ( .A(G104), .B(n1159), .ZN(G6) );
NOR3_X1 U833 ( .A1(n1160), .A2(n1144), .A3(n1161), .ZN(G57) );
NOR3_X1 U834 ( .A1(n1162), .A2(KEYINPUT17), .A3(n1163), .ZN(n1161) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1162) );
NAND2_X1 U836 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
INV_X1 U837 ( .A(KEYINPUT27), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1168), .A2(n1169), .ZN(n1160) );
XNOR2_X1 U839 ( .A(n1164), .B(n1170), .ZN(n1169) );
NOR2_X1 U840 ( .A1(KEYINPUT27), .A2(n1167), .ZN(n1170) );
NAND2_X1 U841 ( .A1(n1147), .A2(G472), .ZN(n1167) );
NAND3_X1 U842 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1164) );
OR2_X1 U843 ( .A1(n1174), .A2(KEYINPUT40), .ZN(n1173) );
NAND4_X1 U844 ( .A1(n1174), .A2(n1175), .A3(KEYINPUT40), .A4(n1176), .ZN(n1172) );
INV_X1 U845 ( .A(G101), .ZN(n1176) );
NAND2_X1 U846 ( .A1(G101), .A2(n1177), .ZN(n1171) );
NAND2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(n1177) );
INV_X1 U848 ( .A(KEYINPUT55), .ZN(n1175) );
NOR2_X1 U849 ( .A1(KEYINPUT17), .A2(n1163), .ZN(n1168) );
XNOR2_X1 U850 ( .A(n1178), .B(n1179), .ZN(n1163) );
NOR2_X1 U851 ( .A1(n1144), .A2(n1180), .ZN(G54) );
NOR2_X1 U852 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U853 ( .A(n1183), .B(KEYINPUT11), .Z(n1182) );
NAND2_X1 U854 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U855 ( .A1(n1184), .A2(n1185), .ZN(n1181) );
XNOR2_X1 U856 ( .A(n1186), .B(KEYINPUT62), .ZN(n1185) );
AND2_X1 U857 ( .A1(n1147), .A2(G469), .ZN(n1184) );
NOR2_X1 U858 ( .A1(n1144), .A2(n1187), .ZN(G51) );
XOR2_X1 U859 ( .A(n1188), .B(n1189), .Z(n1187) );
XNOR2_X1 U860 ( .A(n1190), .B(n1191), .ZN(n1189) );
XNOR2_X1 U861 ( .A(n1192), .B(n1193), .ZN(n1188) );
NAND2_X1 U862 ( .A1(n1147), .A2(G210), .ZN(n1192) );
AND2_X1 U863 ( .A1(G902), .A2(n1194), .ZN(n1147) );
NAND2_X1 U864 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XNOR2_X1 U865 ( .A(KEYINPUT57), .B(n1057), .ZN(n1196) );
NAND4_X1 U866 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1057) );
AND4_X1 U867 ( .A1(n1201), .A2(n1202), .A3(n1159), .A4(n1050), .ZN(n1200) );
NAND3_X1 U868 ( .A1(n1069), .A2(n1070), .A3(n1203), .ZN(n1050) );
NAND3_X1 U869 ( .A1(n1070), .A2(n1072), .A3(n1203), .ZN(n1159) );
NAND2_X1 U870 ( .A1(n1204), .A2(n1205), .ZN(n1199) );
NAND2_X1 U871 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND3_X1 U872 ( .A1(n1070), .A2(n1208), .A3(n1209), .ZN(n1207) );
NAND3_X1 U873 ( .A1(n1073), .A2(n1072), .A3(n1210), .ZN(n1206) );
XNOR2_X1 U874 ( .A(KEYINPUT33), .B(n1208), .ZN(n1210) );
INV_X1 U875 ( .A(n1055), .ZN(n1195) );
NAND4_X1 U876 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1055) );
NOR4_X1 U877 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NOR3_X1 U878 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1213) );
NOR2_X1 U879 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NAND4_X1 U880 ( .A1(n1073), .A2(n1209), .A3(n1224), .A4(n1225), .ZN(n1223) );
INV_X1 U881 ( .A(KEYINPUT45), .ZN(n1222) );
NOR2_X1 U882 ( .A1(KEYINPUT45), .A2(n1226), .ZN(n1220) );
AND2_X1 U883 ( .A1(n1227), .A2(n1228), .ZN(n1219) );
NOR2_X1 U884 ( .A1(n1079), .A2(G952), .ZN(n1144) );
XOR2_X1 U885 ( .A(G146), .B(n1218), .Z(G48) );
AND2_X1 U886 ( .A1(n1229), .A2(n1072), .ZN(n1218) );
XNOR2_X1 U887 ( .A(G143), .B(n1226), .ZN(G45) );
NAND4_X1 U888 ( .A1(n1073), .A2(n1230), .A3(n1209), .A4(n1224), .ZN(n1226) );
XNOR2_X1 U889 ( .A(G140), .B(n1231), .ZN(G42) );
NAND3_X1 U890 ( .A1(n1228), .A2(n1227), .A3(KEYINPUT16), .ZN(n1231) );
NAND2_X1 U891 ( .A1(n1232), .A2(n1233), .ZN(G39) );
NAND2_X1 U892 ( .A1(n1234), .A2(n1117), .ZN(n1233) );
XOR2_X1 U893 ( .A(n1211), .B(KEYINPUT50), .Z(n1234) );
NAND2_X1 U894 ( .A1(n1235), .A2(G137), .ZN(n1232) );
XNOR2_X1 U895 ( .A(KEYINPUT35), .B(n1211), .ZN(n1235) );
NAND3_X1 U896 ( .A1(n1102), .A2(n1228), .A3(n1236), .ZN(n1211) );
XOR2_X1 U897 ( .A(G134), .B(n1217), .Z(G36) );
AND3_X1 U898 ( .A1(n1228), .A2(n1069), .A3(n1073), .ZN(n1217) );
XNOR2_X1 U899 ( .A(G131), .B(n1212), .ZN(G33) );
NAND3_X1 U900 ( .A1(n1228), .A2(n1072), .A3(n1073), .ZN(n1212) );
AND3_X1 U901 ( .A1(n1086), .A2(n1090), .A3(n1230), .ZN(n1228) );
INV_X1 U902 ( .A(n1060), .ZN(n1086) );
NAND2_X1 U903 ( .A1(n1237), .A2(n1095), .ZN(n1060) );
INV_X1 U904 ( .A(n1094), .ZN(n1237) );
XOR2_X1 U905 ( .A(G128), .B(n1216), .Z(G30) );
AND2_X1 U906 ( .A1(n1229), .A2(n1069), .ZN(n1216) );
AND4_X1 U907 ( .A1(n1238), .A2(n1230), .A3(n1102), .A4(n1224), .ZN(n1229) );
XNOR2_X1 U908 ( .A(G101), .B(n1239), .ZN(G3) );
NOR2_X1 U909 ( .A1(n1240), .A2(KEYINPUT29), .ZN(n1239) );
INV_X1 U910 ( .A(n1202), .ZN(n1240) );
NAND3_X1 U911 ( .A1(n1203), .A2(n1074), .A3(n1073), .ZN(n1202) );
XOR2_X1 U912 ( .A(n1215), .B(n1241), .Z(G27) );
NOR2_X1 U913 ( .A1(KEYINPUT43), .A2(n1193), .ZN(n1241) );
AND3_X1 U914 ( .A1(n1230), .A2(n1227), .A3(n1204), .ZN(n1215) );
NOR3_X1 U915 ( .A1(n1242), .A2(n1102), .A3(n1243), .ZN(n1227) );
INV_X1 U916 ( .A(n1225), .ZN(n1230) );
NAND3_X1 U917 ( .A1(n1244), .A2(n1245), .A3(n1076), .ZN(n1225) );
NAND2_X1 U918 ( .A1(G953), .A2(n1246), .ZN(n1245) );
OR2_X1 U919 ( .A1(n1247), .A2(G900), .ZN(n1246) );
NAND2_X1 U920 ( .A1(n1248), .A2(n1079), .ZN(n1244) );
NAND2_X1 U921 ( .A1(n1249), .A2(n1250), .ZN(G24) );
NAND2_X1 U922 ( .A1(G122), .A2(n1251), .ZN(n1250) );
XOR2_X1 U923 ( .A(KEYINPUT42), .B(n1252), .Z(n1249) );
NOR2_X1 U924 ( .A1(G122), .A2(n1251), .ZN(n1252) );
NAND4_X1 U925 ( .A1(n1204), .A2(n1209), .A3(n1253), .A4(n1070), .ZN(n1251) );
AND2_X1 U926 ( .A1(n1254), .A2(n1243), .ZN(n1070) );
XOR2_X1 U927 ( .A(n1102), .B(KEYINPUT59), .Z(n1254) );
XOR2_X1 U928 ( .A(n1208), .B(KEYINPUT32), .Z(n1253) );
XNOR2_X1 U929 ( .A(G119), .B(n1197), .ZN(G21) );
NAND4_X1 U930 ( .A1(n1236), .A2(n1204), .A3(n1102), .A4(n1208), .ZN(n1197) );
INV_X1 U931 ( .A(n1255), .ZN(n1236) );
XNOR2_X1 U932 ( .A(G116), .B(n1198), .ZN(G18) );
NAND2_X1 U933 ( .A1(n1256), .A2(n1069), .ZN(n1198) );
INV_X1 U934 ( .A(n1257), .ZN(n1256) );
XNOR2_X1 U935 ( .A(n1258), .B(n1259), .ZN(G15) );
NOR2_X1 U936 ( .A1(n1242), .A2(n1257), .ZN(n1259) );
NAND3_X1 U937 ( .A1(n1204), .A2(n1208), .A3(n1073), .ZN(n1257) );
AND2_X1 U938 ( .A1(n1260), .A2(n1102), .ZN(n1073) );
XNOR2_X1 U939 ( .A(n1243), .B(KEYINPUT51), .ZN(n1260) );
INV_X1 U940 ( .A(n1083), .ZN(n1204) );
NAND3_X1 U941 ( .A1(n1094), .A2(n1095), .A3(n1097), .ZN(n1083) );
INV_X1 U942 ( .A(n1061), .ZN(n1097) );
NAND2_X1 U943 ( .A1(n1093), .A2(n1261), .ZN(n1061) );
INV_X1 U944 ( .A(n1072), .ZN(n1242) );
NAND2_X1 U945 ( .A1(n1262), .A2(n1263), .ZN(n1072) );
NAND2_X1 U946 ( .A1(n1209), .A2(n1264), .ZN(n1263) );
NOR2_X1 U947 ( .A1(n1265), .A2(n1266), .ZN(n1209) );
NAND3_X1 U948 ( .A1(n1265), .A2(n1267), .A3(KEYINPUT0), .ZN(n1262) );
NAND2_X1 U949 ( .A1(n1268), .A2(n1269), .ZN(G12) );
NAND2_X1 U950 ( .A1(G110), .A2(n1201), .ZN(n1269) );
XOR2_X1 U951 ( .A(n1270), .B(KEYINPUT25), .Z(n1268) );
OR2_X1 U952 ( .A1(n1201), .A2(G110), .ZN(n1270) );
NAND2_X1 U953 ( .A1(n1071), .A2(n1203), .ZN(n1201) );
AND2_X1 U954 ( .A1(n1224), .A2(n1208), .ZN(n1203) );
NAND2_X1 U955 ( .A1(n1271), .A2(n1272), .ZN(n1208) );
OR3_X1 U956 ( .A1(n1248), .A2(n1062), .A3(G953), .ZN(n1272) );
INV_X1 U957 ( .A(n1076), .ZN(n1062) );
XOR2_X1 U958 ( .A(G952), .B(KEYINPUT44), .Z(n1248) );
NAND4_X1 U959 ( .A1(n1273), .A2(n1140), .A3(G902), .A4(G953), .ZN(n1271) );
INV_X1 U960 ( .A(G898), .ZN(n1140) );
XNOR2_X1 U961 ( .A(KEYINPUT1), .B(n1076), .ZN(n1273) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1076) );
AND3_X1 U963 ( .A1(n1094), .A2(n1095), .A3(n1090), .ZN(n1224) );
NOR2_X1 U964 ( .A1(n1093), .A2(n1092), .ZN(n1090) );
INV_X1 U965 ( .A(n1261), .ZN(n1092) );
NAND2_X1 U966 ( .A1(n1274), .A2(n1275), .ZN(n1261) );
XOR2_X1 U967 ( .A(KEYINPUT8), .B(G221), .Z(n1274) );
XOR2_X1 U968 ( .A(n1276), .B(G469), .Z(n1093) );
NAND2_X1 U969 ( .A1(n1186), .A2(n1247), .ZN(n1276) );
XNOR2_X1 U970 ( .A(n1277), .B(KEYINPUT18), .ZN(n1186) );
XOR2_X1 U971 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U972 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U973 ( .A(n1282), .B(G104), .ZN(n1281) );
XNOR2_X1 U974 ( .A(n1283), .B(G110), .ZN(n1280) );
INV_X1 U975 ( .A(G140), .ZN(n1283) );
XOR2_X1 U976 ( .A(n1284), .B(n1285), .Z(n1278) );
XOR2_X1 U977 ( .A(n1286), .B(n1287), .Z(n1285) );
NOR2_X1 U978 ( .A1(G101), .A2(KEYINPUT53), .ZN(n1287) );
AND2_X1 U979 ( .A1(n1079), .A2(G227), .ZN(n1286) );
XNOR2_X1 U980 ( .A(n1178), .B(n1118), .ZN(n1284) );
NAND2_X1 U981 ( .A1(G214), .A2(n1288), .ZN(n1095) );
XNOR2_X1 U982 ( .A(n1289), .B(n1290), .ZN(n1094) );
AND2_X1 U983 ( .A1(n1288), .A2(G210), .ZN(n1290) );
NAND2_X1 U984 ( .A1(n1291), .A2(n1247), .ZN(n1288) );
XNOR2_X1 U985 ( .A(KEYINPUT24), .B(n1292), .ZN(n1291) );
NAND2_X1 U986 ( .A1(n1293), .A2(n1247), .ZN(n1289) );
XOR2_X1 U987 ( .A(n1190), .B(n1294), .Z(n1293) );
XNOR2_X1 U988 ( .A(n1193), .B(n1295), .ZN(n1294) );
NOR2_X1 U989 ( .A1(KEYINPUT13), .A2(n1191), .ZN(n1295) );
INV_X1 U990 ( .A(G125), .ZN(n1193) );
XNOR2_X1 U991 ( .A(n1296), .B(n1133), .ZN(n1190) );
INV_X1 U992 ( .A(n1136), .ZN(n1133) );
XOR2_X1 U993 ( .A(G110), .B(n1297), .Z(n1136) );
XOR2_X1 U994 ( .A(n1137), .B(n1298), .Z(n1296) );
AND2_X1 U995 ( .A1(n1079), .A2(G224), .ZN(n1298) );
XOR2_X1 U996 ( .A(n1139), .B(n1138), .Z(n1137) );
XNOR2_X1 U997 ( .A(n1299), .B(n1300), .ZN(n1138) );
NOR2_X1 U998 ( .A1(G104), .A2(n1301), .ZN(n1300) );
XNOR2_X1 U999 ( .A(KEYINPUT22), .B(KEYINPUT20), .ZN(n1301) );
XNOR2_X1 U1000 ( .A(G107), .B(G101), .ZN(n1299) );
NAND3_X1 U1001 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1139) );
NAND2_X1 U1002 ( .A1(KEYINPUT48), .A2(n1305), .ZN(n1304) );
OR3_X1 U1003 ( .A1(n1305), .A2(KEYINPUT48), .A3(n1306), .ZN(n1303) );
NAND2_X1 U1004 ( .A1(n1306), .A2(n1307), .ZN(n1302) );
NAND2_X1 U1005 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
INV_X1 U1006 ( .A(KEYINPUT48), .ZN(n1309) );
XNOR2_X1 U1007 ( .A(n1305), .B(KEYINPUT52), .ZN(n1308) );
AND2_X1 U1008 ( .A1(n1310), .A2(n1311), .ZN(n1305) );
NOR2_X1 U1009 ( .A1(n1255), .A2(n1102), .ZN(n1071) );
XOR2_X1 U1010 ( .A(n1312), .B(n1313), .Z(n1102) );
XOR2_X1 U1011 ( .A(KEYINPUT36), .B(G472), .Z(n1313) );
NAND2_X1 U1012 ( .A1(n1314), .A2(n1247), .ZN(n1312) );
XOR2_X1 U1013 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1014 ( .A(n1317), .B(n1174), .Z(n1316) );
AND3_X1 U1015 ( .A1(n1292), .A2(n1079), .A3(G210), .ZN(n1174) );
NAND2_X1 U1016 ( .A1(n1318), .A2(KEYINPUT9), .ZN(n1317) );
XOR2_X1 U1017 ( .A(n1319), .B(n1179), .Z(n1318) );
XNOR2_X1 U1018 ( .A(n1191), .B(n1320), .ZN(n1179) );
XNOR2_X1 U1019 ( .A(n1321), .B(n1306), .ZN(n1320) );
XOR2_X1 U1020 ( .A(G113), .B(KEYINPUT2), .Z(n1306) );
NAND2_X1 U1021 ( .A1(n1322), .A2(n1310), .ZN(n1321) );
NAND2_X1 U1022 ( .A1(G116), .A2(n1323), .ZN(n1310) );
INV_X1 U1023 ( .A(G119), .ZN(n1323) );
XOR2_X1 U1024 ( .A(n1311), .B(KEYINPUT60), .Z(n1322) );
NAND2_X1 U1025 ( .A1(G119), .A2(n1324), .ZN(n1311) );
INV_X1 U1026 ( .A(G116), .ZN(n1324) );
XNOR2_X1 U1027 ( .A(n1118), .B(KEYINPUT4), .ZN(n1191) );
XOR2_X1 U1028 ( .A(G143), .B(n1325), .Z(n1118) );
NAND2_X1 U1029 ( .A1(KEYINPUT26), .A2(n1326), .ZN(n1319) );
XNOR2_X1 U1030 ( .A(KEYINPUT28), .B(n1327), .ZN(n1326) );
INV_X1 U1031 ( .A(n1178), .ZN(n1327) );
XNOR2_X1 U1032 ( .A(n1328), .B(n1119), .ZN(n1178) );
XOR2_X1 U1033 ( .A(G131), .B(KEYINPUT58), .Z(n1119) );
NAND2_X1 U1034 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1035 ( .A1(G134), .A2(n1117), .ZN(n1330) );
XOR2_X1 U1036 ( .A(KEYINPUT23), .B(n1331), .Z(n1329) );
NOR2_X1 U1037 ( .A1(G134), .A2(n1117), .ZN(n1331) );
XNOR2_X1 U1038 ( .A(G101), .B(KEYINPUT21), .ZN(n1315) );
NAND2_X1 U1039 ( .A1(n1238), .A2(n1074), .ZN(n1255) );
NAND2_X1 U1040 ( .A1(n1332), .A2(n1333), .ZN(n1074) );
NAND2_X1 U1041 ( .A1(n1069), .A2(n1264), .ZN(n1333) );
INV_X1 U1042 ( .A(KEYINPUT0), .ZN(n1264) );
NOR2_X1 U1043 ( .A1(n1267), .A2(n1265), .ZN(n1069) );
INV_X1 U1044 ( .A(n1266), .ZN(n1267) );
NAND3_X1 U1045 ( .A1(n1266), .A2(n1265), .A3(KEYINPUT0), .ZN(n1332) );
INV_X1 U1046 ( .A(n1103), .ZN(n1265) );
XNOR2_X1 U1047 ( .A(n1334), .B(G478), .ZN(n1103) );
NAND2_X1 U1048 ( .A1(n1335), .A2(n1247), .ZN(n1334) );
INV_X1 U1049 ( .A(n1152), .ZN(n1335) );
XNOR2_X1 U1050 ( .A(n1336), .B(n1337), .ZN(n1152) );
XNOR2_X1 U1051 ( .A(n1282), .B(n1338), .ZN(n1337) );
XNOR2_X1 U1052 ( .A(n1339), .B(G128), .ZN(n1338) );
INV_X1 U1053 ( .A(G107), .ZN(n1282) );
XOR2_X1 U1054 ( .A(n1340), .B(n1341), .Z(n1336) );
XNOR2_X1 U1055 ( .A(n1342), .B(n1343), .ZN(n1341) );
NOR2_X1 U1056 ( .A1(G134), .A2(KEYINPUT10), .ZN(n1343) );
NAND2_X1 U1057 ( .A1(n1344), .A2(KEYINPUT41), .ZN(n1342) );
XNOR2_X1 U1058 ( .A(G116), .B(n1297), .ZN(n1344) );
NAND2_X1 U1059 ( .A1(G217), .A2(n1345), .ZN(n1340) );
NOR2_X1 U1060 ( .A1(n1346), .A2(n1101), .ZN(n1266) );
NOR3_X1 U1061 ( .A1(G475), .A2(G902), .A3(n1158), .ZN(n1101) );
XOR2_X1 U1062 ( .A(n1100), .B(KEYINPUT30), .Z(n1346) );
AND2_X1 U1063 ( .A1(G475), .A2(n1347), .ZN(n1100) );
OR2_X1 U1064 ( .A1(n1158), .A2(G902), .ZN(n1347) );
XOR2_X1 U1065 ( .A(n1348), .B(n1349), .Z(n1158) );
XOR2_X1 U1066 ( .A(n1114), .B(n1350), .Z(n1349) );
XOR2_X1 U1067 ( .A(n1351), .B(n1352), .Z(n1350) );
NAND2_X1 U1068 ( .A1(n1353), .A2(KEYINPUT15), .ZN(n1352) );
XOR2_X1 U1069 ( .A(n1354), .B(n1355), .Z(n1353) );
AND3_X1 U1070 ( .A1(G214), .A2(n1079), .A3(n1292), .ZN(n1355) );
INV_X1 U1071 ( .A(G237), .ZN(n1292) );
NAND2_X1 U1072 ( .A1(KEYINPUT31), .A2(n1339), .ZN(n1354) );
INV_X1 U1073 ( .A(G143), .ZN(n1339) );
NAND2_X1 U1074 ( .A1(n1356), .A2(n1357), .ZN(n1351) );
NAND2_X1 U1075 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
NAND2_X1 U1076 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
NAND2_X1 U1077 ( .A1(n1258), .A2(n1362), .ZN(n1361) );
INV_X1 U1078 ( .A(G113), .ZN(n1258) );
INV_X1 U1079 ( .A(KEYINPUT12), .ZN(n1360) );
NAND2_X1 U1080 ( .A1(G113), .A2(n1363), .ZN(n1356) );
NAND2_X1 U1081 ( .A1(n1362), .A2(n1364), .ZN(n1363) );
OR2_X1 U1082 ( .A1(n1358), .A2(KEYINPUT12), .ZN(n1364) );
XOR2_X1 U1083 ( .A(n1297), .B(KEYINPUT37), .Z(n1358) );
XOR2_X1 U1084 ( .A(G122), .B(KEYINPUT6), .Z(n1297) );
INV_X1 U1085 ( .A(KEYINPUT49), .ZN(n1362) );
XNOR2_X1 U1086 ( .A(G104), .B(n1365), .ZN(n1348) );
XOR2_X1 U1087 ( .A(G146), .B(G131), .Z(n1365) );
INV_X1 U1088 ( .A(n1243), .ZN(n1238) );
XNOR2_X1 U1089 ( .A(n1104), .B(n1366), .ZN(n1243) );
NOR2_X1 U1090 ( .A1(n1105), .A2(KEYINPUT61), .ZN(n1366) );
AND2_X1 U1091 ( .A1(G217), .A2(n1275), .ZN(n1105) );
NAND2_X1 U1092 ( .A1(G234), .A2(n1247), .ZN(n1275) );
NAND2_X1 U1093 ( .A1(n1146), .A2(n1247), .ZN(n1104) );
INV_X1 U1094 ( .A(G902), .ZN(n1247) );
XNOR2_X1 U1095 ( .A(n1367), .B(n1368), .ZN(n1146) );
XOR2_X1 U1096 ( .A(G110), .B(n1369), .Z(n1368) );
XNOR2_X1 U1097 ( .A(n1117), .B(G119), .ZN(n1369) );
INV_X1 U1098 ( .A(G137), .ZN(n1117) );
XOR2_X1 U1099 ( .A(n1370), .B(n1325), .Z(n1367) );
XOR2_X1 U1100 ( .A(G128), .B(G146), .Z(n1325) );
XOR2_X1 U1101 ( .A(n1371), .B(n1114), .Z(n1370) );
XOR2_X1 U1102 ( .A(G140), .B(G125), .Z(n1114) );
NAND2_X1 U1103 ( .A1(n1345), .A2(G221), .ZN(n1371) );
AND2_X1 U1104 ( .A1(G234), .A2(n1079), .ZN(n1345) );
INV_X1 U1105 ( .A(G953), .ZN(n1079) );
endmodule


