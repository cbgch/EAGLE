//Key = 1000011111110100000000000101110000010110111110000011101111111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335;

XOR2_X1 U724 ( .A(n1019), .B(n1020), .Z(G9) );
NAND4_X1 U725 ( .A1(KEYINPUT11), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1020) );
XOR2_X1 U726 ( .A(KEYINPUT49), .B(n1024), .Z(n1023) );
NOR2_X1 U727 ( .A1(n1025), .A2(n1026), .ZN(G75) );
AND4_X1 U728 ( .A1(n1027), .A2(n1028), .A3(KEYINPUT58), .A4(n1029), .ZN(n1026) );
NOR4_X1 U729 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
NOR2_X1 U730 ( .A1(KEYINPUT43), .A2(n1034), .ZN(n1033) );
NOR4_X1 U731 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
NOR2_X1 U732 ( .A1(n1039), .A2(n1038), .ZN(n1032) );
NAND4_X1 U733 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1038) );
INV_X1 U734 ( .A(n1044), .ZN(n1040) );
NOR2_X1 U735 ( .A1(n1045), .A2(n1046), .ZN(n1039) );
NOR2_X1 U736 ( .A1(n1047), .A2(n1035), .ZN(n1046) );
NOR2_X1 U737 ( .A1(n1048), .A2(n1024), .ZN(n1047) );
AND3_X1 U738 ( .A1(KEYINPUT43), .A2(n1049), .A3(n1050), .ZN(n1048) );
NOR2_X1 U739 ( .A1(n1051), .A2(n1052), .ZN(n1045) );
NOR2_X1 U740 ( .A1(n1053), .A2(n1021), .ZN(n1051) );
NOR4_X1 U741 ( .A1(n1054), .A2(n1035), .A3(n1052), .A4(n1044), .ZN(n1031) );
NOR2_X1 U742 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
AND2_X1 U743 ( .A1(n1057), .A2(n1041), .ZN(n1056) );
NOR2_X1 U744 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
NOR2_X1 U745 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
AND2_X1 U746 ( .A1(n1062), .A2(n1041), .ZN(n1061) );
NOR2_X1 U747 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NOR2_X1 U748 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U749 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U750 ( .A1(n1069), .A2(G952), .A3(n1030), .ZN(n1025) );
AND4_X1 U751 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1030) );
NOR4_X1 U752 ( .A1(n1049), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1073) );
XNOR2_X1 U753 ( .A(n1077), .B(n1078), .ZN(n1076) );
XOR2_X1 U754 ( .A(n1079), .B(KEYINPUT13), .Z(n1077) );
XNOR2_X1 U755 ( .A(n1080), .B(n1081), .ZN(n1075) );
NAND2_X1 U756 ( .A1(KEYINPUT63), .A2(n1082), .ZN(n1080) );
NOR2_X1 U757 ( .A1(n1036), .A2(n1083), .ZN(n1072) );
INV_X1 U758 ( .A(n1050), .ZN(n1036) );
XOR2_X1 U759 ( .A(n1084), .B(KEYINPUT28), .Z(n1071) );
NAND2_X1 U760 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U761 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U762 ( .A(n1089), .B(KEYINPUT1), .Z(n1085) );
OR2_X1 U763 ( .A1(n1088), .A2(n1087), .ZN(n1089) );
XNOR2_X1 U764 ( .A(n1090), .B(KEYINPUT59), .ZN(n1088) );
XOR2_X1 U765 ( .A(n1042), .B(KEYINPUT48), .Z(n1070) );
INV_X1 U766 ( .A(n1027), .ZN(n1069) );
XOR2_X1 U767 ( .A(n1091), .B(n1092), .Z(G72) );
NOR2_X1 U768 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U769 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND2_X1 U770 ( .A1(n1097), .A2(n1098), .ZN(n1091) );
NAND2_X1 U771 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U772 ( .A(n1101), .B(n1102), .ZN(n1099) );
OR3_X1 U773 ( .A1(n1096), .A2(n1101), .A3(n1100), .ZN(n1097) );
NAND2_X1 U774 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NAND2_X1 U775 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U776 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
INV_X1 U777 ( .A(n1109), .ZN(n1105) );
NAND3_X1 U778 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1103) );
NAND2_X1 U779 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
XOR2_X1 U780 ( .A(KEYINPUT8), .B(n1112), .Z(n1111) );
XOR2_X1 U781 ( .A(n1113), .B(KEYINPUT37), .Z(n1110) );
XNOR2_X1 U782 ( .A(KEYINPUT51), .B(n1114), .ZN(n1107) );
NAND2_X1 U783 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U784 ( .A(KEYINPUT37), .B(n1117), .Z(n1116) );
INV_X1 U785 ( .A(n1113), .ZN(n1117) );
XOR2_X1 U786 ( .A(KEYINPUT8), .B(n1118), .Z(n1115) );
XOR2_X1 U787 ( .A(n1119), .B(n1120), .Z(G69) );
NOR2_X1 U788 ( .A1(n1121), .A2(n1094), .ZN(n1120) );
XOR2_X1 U789 ( .A(n1100), .B(KEYINPUT23), .Z(n1094) );
NOR2_X1 U790 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U791 ( .A1(n1124), .A2(n1125), .ZN(n1119) );
NAND3_X1 U792 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1125) );
NAND2_X1 U793 ( .A1(G953), .A2(n1123), .ZN(n1127) );
NAND2_X1 U794 ( .A1(n1129), .A2(n1100), .ZN(n1126) );
XOR2_X1 U795 ( .A(n1130), .B(KEYINPUT12), .Z(n1124) );
NAND3_X1 U796 ( .A1(n1129), .A2(n1100), .A3(n1131), .ZN(n1130) );
NOR2_X1 U797 ( .A1(n1132), .A2(n1133), .ZN(G66) );
NOR3_X1 U798 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR3_X1 U799 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
NOR2_X1 U800 ( .A1(n1140), .A2(n1141), .ZN(n1135) );
INV_X1 U801 ( .A(n1137), .ZN(n1141) );
NOR2_X1 U802 ( .A1(n1028), .A2(n1138), .ZN(n1140) );
XOR2_X1 U803 ( .A(G217), .B(KEYINPUT27), .Z(n1138) );
NOR2_X1 U804 ( .A1(n1132), .A2(n1142), .ZN(G63) );
XNOR2_X1 U805 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U806 ( .A1(n1145), .A2(n1139), .ZN(n1144) );
INV_X1 U807 ( .A(G478), .ZN(n1145) );
NOR2_X1 U808 ( .A1(n1132), .A2(n1146), .ZN(G60) );
NOR3_X1 U809 ( .A1(n1147), .A2(n1087), .A3(n1148), .ZN(n1146) );
NOR2_X1 U810 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U811 ( .A1(n1028), .A2(n1090), .ZN(n1149) );
XOR2_X1 U812 ( .A(KEYINPUT16), .B(n1151), .Z(n1147) );
NOR3_X1 U813 ( .A1(n1139), .A2(n1152), .A3(n1090), .ZN(n1151) );
INV_X1 U814 ( .A(G475), .ZN(n1090) );
XNOR2_X1 U815 ( .A(G104), .B(n1153), .ZN(G6) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1154), .ZN(G57) );
XOR2_X1 U817 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U818 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U819 ( .A(n1159), .B(n1160), .Z(n1155) );
NOR3_X1 U820 ( .A1(n1139), .A2(KEYINPUT14), .A3(n1161), .ZN(n1160) );
INV_X1 U821 ( .A(G472), .ZN(n1161) );
XNOR2_X1 U822 ( .A(KEYINPUT46), .B(n1162), .ZN(n1159) );
NOR2_X1 U823 ( .A1(KEYINPUT53), .A2(n1163), .ZN(n1162) );
NOR2_X1 U824 ( .A1(n1132), .A2(n1164), .ZN(G54) );
XOR2_X1 U825 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U826 ( .A(n1167), .B(n1112), .Z(n1166) );
NOR2_X1 U827 ( .A1(n1168), .A2(n1139), .ZN(n1167) );
INV_X1 U828 ( .A(G469), .ZN(n1168) );
XOR2_X1 U829 ( .A(n1169), .B(n1170), .Z(n1165) );
XOR2_X1 U830 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U831 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U832 ( .A(KEYINPUT33), .B(n1175), .Z(n1174) );
NOR2_X1 U833 ( .A1(n1113), .A2(n1176), .ZN(n1175) );
AND2_X1 U834 ( .A1(n1113), .A2(n1176), .ZN(n1173) );
NOR3_X1 U835 ( .A1(KEYINPUT3), .A2(n1177), .A3(n1178), .ZN(n1169) );
NOR3_X1 U836 ( .A1(KEYINPUT40), .A2(G110), .A3(n1179), .ZN(n1178) );
NOR2_X1 U837 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
INV_X1 U838 ( .A(KEYINPUT40), .ZN(n1181) );
NOR2_X1 U839 ( .A1(n1132), .A2(n1182), .ZN(G51) );
XOR2_X1 U840 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U841 ( .A1(n1081), .A2(n1139), .ZN(n1184) );
OR2_X1 U842 ( .A1(n1185), .A2(n1028), .ZN(n1139) );
NOR2_X1 U843 ( .A1(n1129), .A2(n1102), .ZN(n1028) );
NAND4_X1 U844 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1102) );
AND4_X1 U845 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
AND2_X1 U846 ( .A1(n1194), .A2(n1195), .ZN(n1188) );
NAND3_X1 U847 ( .A1(n1196), .A2(n1197), .A3(n1041), .ZN(n1186) );
NAND4_X1 U848 ( .A1(n1153), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1129) );
AND4_X1 U849 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NAND2_X1 U850 ( .A1(n1022), .A2(n1205), .ZN(n1199) );
NAND2_X1 U851 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND3_X1 U852 ( .A1(n1083), .A2(n1208), .A3(n1209), .ZN(n1207) );
NAND2_X1 U853 ( .A1(n1021), .A2(n1024), .ZN(n1206) );
NAND3_X1 U854 ( .A1(n1022), .A2(n1024), .A3(n1053), .ZN(n1153) );
NAND4_X1 U855 ( .A1(KEYINPUT5), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1183) );
NAND3_X1 U856 ( .A1(KEYINPUT25), .A2(n1213), .A3(n1131), .ZN(n1212) );
OR2_X1 U857 ( .A1(n1131), .A2(n1213), .ZN(n1211) );
NOR2_X1 U858 ( .A1(KEYINPUT32), .A2(n1214), .ZN(n1213) );
INV_X1 U859 ( .A(n1128), .ZN(n1131) );
NAND2_X1 U860 ( .A1(n1214), .A2(n1215), .ZN(n1210) );
INV_X1 U861 ( .A(KEYINPUT25), .ZN(n1215) );
XNOR2_X1 U862 ( .A(n1216), .B(n1217), .ZN(n1214) );
XOR2_X1 U863 ( .A(KEYINPUT61), .B(n1218), .Z(n1217) );
NAND2_X1 U864 ( .A1(n1219), .A2(n1220), .ZN(n1216) );
OR2_X1 U865 ( .A1(n1221), .A2(G125), .ZN(n1220) );
XOR2_X1 U866 ( .A(n1222), .B(KEYINPUT26), .Z(n1219) );
NAND2_X1 U867 ( .A1(G125), .A2(n1221), .ZN(n1222) );
NOR2_X1 U868 ( .A1(n1100), .A2(G952), .ZN(n1132) );
XNOR2_X1 U869 ( .A(G146), .B(n1190), .ZN(G48) );
NAND3_X1 U870 ( .A1(n1053), .A2(n1066), .A3(n1196), .ZN(n1190) );
XOR2_X1 U871 ( .A(n1223), .B(n1187), .Z(G45) );
NAND4_X1 U872 ( .A1(n1224), .A2(n1066), .A3(n1083), .A4(n1208), .ZN(n1187) );
XOR2_X1 U873 ( .A(n1179), .B(n1195), .Z(G42) );
NAND3_X1 U874 ( .A1(n1225), .A2(n1226), .A3(n1041), .ZN(n1195) );
XOR2_X1 U875 ( .A(n1227), .B(n1228), .Z(G39) );
NAND2_X1 U876 ( .A1(n1229), .A2(G137), .ZN(n1228) );
XNOR2_X1 U877 ( .A(KEYINPUT30), .B(KEYINPUT24), .ZN(n1229) );
NAND2_X1 U878 ( .A1(n1041), .A2(n1230), .ZN(n1227) );
XOR2_X1 U879 ( .A(KEYINPUT34), .B(n1231), .Z(n1230) );
NOR2_X1 U880 ( .A1(n1035), .A2(n1232), .ZN(n1231) );
INV_X1 U881 ( .A(n1197), .ZN(n1035) );
XNOR2_X1 U882 ( .A(G134), .B(n1194), .ZN(G36) );
NAND3_X1 U883 ( .A1(n1224), .A2(n1021), .A3(n1041), .ZN(n1194) );
XOR2_X1 U884 ( .A(n1193), .B(n1233), .Z(G33) );
XNOR2_X1 U885 ( .A(G131), .B(KEYINPUT17), .ZN(n1233) );
NAND3_X1 U886 ( .A1(n1224), .A2(n1053), .A3(n1041), .ZN(n1193) );
NOR2_X1 U887 ( .A1(n1067), .A2(n1074), .ZN(n1041) );
INV_X1 U888 ( .A(n1068), .ZN(n1074) );
AND2_X1 U889 ( .A1(n1226), .A2(n1057), .ZN(n1224) );
NAND2_X1 U890 ( .A1(n1234), .A2(n1235), .ZN(G30) );
NAND2_X1 U891 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
XOR2_X1 U892 ( .A(n1238), .B(KEYINPUT19), .Z(n1234) );
OR2_X1 U893 ( .A1(n1237), .A2(n1236), .ZN(n1238) );
INV_X1 U894 ( .A(n1192), .ZN(n1236) );
NAND3_X1 U895 ( .A1(n1021), .A2(n1066), .A3(n1196), .ZN(n1192) );
INV_X1 U896 ( .A(n1232), .ZN(n1196) );
NAND3_X1 U897 ( .A1(n1062), .A2(n1059), .A3(n1226), .ZN(n1232) );
AND2_X1 U898 ( .A1(n1024), .A2(n1239), .ZN(n1226) );
XNOR2_X1 U899 ( .A(n1240), .B(KEYINPUT60), .ZN(n1237) );
XOR2_X1 U900 ( .A(n1241), .B(n1198), .Z(G3) );
NAND4_X1 U901 ( .A1(n1057), .A2(n1024), .A3(n1242), .A4(n1197), .ZN(n1198) );
XOR2_X1 U902 ( .A(n1191), .B(n1243), .Z(G27) );
XNOR2_X1 U903 ( .A(G125), .B(KEYINPUT36), .ZN(n1243) );
NAND4_X1 U904 ( .A1(n1225), .A2(n1209), .A3(n1066), .A4(n1239), .ZN(n1191) );
NAND2_X1 U905 ( .A1(n1044), .A2(n1244), .ZN(n1239) );
NAND4_X1 U906 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1096), .ZN(n1244) );
INV_X1 U907 ( .A(G900), .ZN(n1096) );
AND3_X1 U908 ( .A1(n1042), .A2(n1062), .A3(n1053), .ZN(n1225) );
XNOR2_X1 U909 ( .A(G122), .B(n1246), .ZN(G24) );
NAND3_X1 U910 ( .A1(n1209), .A2(n1022), .A3(n1247), .ZN(n1246) );
NOR3_X1 U911 ( .A1(n1248), .A2(KEYINPUT21), .A3(n1249), .ZN(n1247) );
AND3_X1 U912 ( .A1(n1042), .A2(n1043), .A3(n1242), .ZN(n1022) );
INV_X1 U913 ( .A(n1064), .ZN(n1043) );
XNOR2_X1 U914 ( .A(n1204), .B(n1250), .ZN(G21) );
NOR2_X1 U915 ( .A1(KEYINPUT22), .A2(n1251), .ZN(n1250) );
XOR2_X1 U916 ( .A(KEYINPUT54), .B(G119), .Z(n1251) );
NAND3_X1 U917 ( .A1(n1252), .A2(n1059), .A3(n1209), .ZN(n1204) );
INV_X1 U918 ( .A(n1042), .ZN(n1059) );
XNOR2_X1 U919 ( .A(G116), .B(n1203), .ZN(G18) );
NAND2_X1 U920 ( .A1(n1253), .A2(n1021), .ZN(n1203) );
XOR2_X1 U921 ( .A(n1202), .B(n1254), .Z(G15) );
XOR2_X1 U922 ( .A(KEYINPUT7), .B(G113), .Z(n1254) );
NAND2_X1 U923 ( .A1(n1053), .A2(n1253), .ZN(n1202) );
AND3_X1 U924 ( .A1(n1209), .A2(n1242), .A3(n1057), .ZN(n1253) );
NOR2_X1 U925 ( .A1(n1064), .A2(n1042), .ZN(n1057) );
INV_X1 U926 ( .A(n1052), .ZN(n1209) );
NAND2_X1 U927 ( .A1(n1255), .A2(n1037), .ZN(n1052) );
XOR2_X1 U928 ( .A(n1050), .B(KEYINPUT2), .Z(n1255) );
AND2_X1 U929 ( .A1(n1256), .A2(n1208), .ZN(n1053) );
XOR2_X1 U930 ( .A(KEYINPUT56), .B(n1083), .Z(n1256) );
INV_X1 U931 ( .A(n1248), .ZN(n1083) );
XNOR2_X1 U932 ( .A(G110), .B(n1201), .ZN(G12) );
NAND3_X1 U933 ( .A1(n1042), .A2(n1024), .A3(n1252), .ZN(n1201) );
AND3_X1 U934 ( .A1(n1197), .A2(n1062), .A3(n1242), .ZN(n1252) );
AND2_X1 U935 ( .A1(n1066), .A2(n1257), .ZN(n1242) );
NAND2_X1 U936 ( .A1(n1044), .A2(n1258), .ZN(n1257) );
NAND4_X1 U937 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1123), .ZN(n1258) );
INV_X1 U938 ( .A(G898), .ZN(n1123) );
NAND3_X1 U939 ( .A1(n1027), .A2(n1245), .A3(G952), .ZN(n1044) );
NAND2_X1 U940 ( .A1(G237), .A2(G234), .ZN(n1245) );
XOR2_X1 U941 ( .A(n1100), .B(KEYINPUT39), .Z(n1027) );
AND2_X1 U942 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U943 ( .A1(G214), .A2(n1259), .ZN(n1068) );
XOR2_X1 U944 ( .A(n1082), .B(n1081), .Z(n1067) );
NAND2_X1 U945 ( .A1(G210), .A2(n1259), .ZN(n1081) );
NAND2_X1 U946 ( .A1(n1260), .A2(n1185), .ZN(n1259) );
INV_X1 U947 ( .A(G237), .ZN(n1260) );
NAND2_X1 U948 ( .A1(n1261), .A2(n1185), .ZN(n1082) );
XOR2_X1 U949 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U950 ( .A(n1128), .B(n1221), .Z(n1263) );
XOR2_X1 U951 ( .A(n1264), .B(n1265), .Z(n1128) );
XOR2_X1 U952 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U953 ( .A(n1019), .B(G110), .Z(n1267) );
NAND2_X1 U954 ( .A1(KEYINPUT57), .A2(G122), .ZN(n1266) );
XOR2_X1 U955 ( .A(n1268), .B(n1269), .Z(n1264) );
XNOR2_X1 U956 ( .A(n1218), .B(n1270), .ZN(n1262) );
XOR2_X1 U957 ( .A(KEYINPUT55), .B(G125), .Z(n1270) );
NOR2_X1 U958 ( .A1(n1122), .A2(G953), .ZN(n1218) );
INV_X1 U959 ( .A(G224), .ZN(n1122) );
XNOR2_X1 U960 ( .A(n1064), .B(KEYINPUT42), .ZN(n1062) );
XOR2_X1 U961 ( .A(n1271), .B(n1134), .Z(n1064) );
INV_X1 U962 ( .A(n1079), .ZN(n1134) );
NAND2_X1 U963 ( .A1(n1137), .A2(n1185), .ZN(n1079) );
XOR2_X1 U964 ( .A(n1272), .B(n1273), .Z(n1137) );
XOR2_X1 U965 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U966 ( .A(G137), .B(G128), .Z(n1275) );
XOR2_X1 U967 ( .A(KEYINPUT0), .B(G146), .Z(n1274) );
XOR2_X1 U968 ( .A(n1276), .B(n1277), .Z(n1272) );
XOR2_X1 U969 ( .A(G125), .B(G119), .Z(n1277) );
XOR2_X1 U970 ( .A(n1278), .B(n1180), .Z(n1276) );
NAND2_X1 U971 ( .A1(G221), .A2(n1279), .ZN(n1278) );
NAND2_X1 U972 ( .A1(KEYINPUT52), .A2(n1078), .ZN(n1271) );
NAND2_X1 U973 ( .A1(G217), .A2(n1280), .ZN(n1078) );
NAND2_X1 U974 ( .A1(n1281), .A2(n1282), .ZN(n1197) );
NAND2_X1 U975 ( .A1(n1021), .A2(n1283), .ZN(n1282) );
INV_X1 U976 ( .A(KEYINPUT56), .ZN(n1283) );
NOR2_X1 U977 ( .A1(n1208), .A2(n1248), .ZN(n1021) );
NAND3_X1 U978 ( .A1(n1249), .A2(n1248), .A3(KEYINPUT56), .ZN(n1281) );
XOR2_X1 U979 ( .A(n1284), .B(G478), .Z(n1248) );
NAND2_X1 U980 ( .A1(n1143), .A2(n1185), .ZN(n1284) );
XNOR2_X1 U981 ( .A(n1285), .B(n1286), .ZN(n1143) );
XOR2_X1 U982 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U983 ( .A(n1289), .B(n1290), .Z(n1288) );
NAND2_X1 U984 ( .A1(KEYINPUT35), .A2(n1019), .ZN(n1289) );
XOR2_X1 U985 ( .A(n1291), .B(n1292), .Z(n1285) );
XOR2_X1 U986 ( .A(KEYINPUT20), .B(G128), .Z(n1292) );
XOR2_X1 U987 ( .A(n1293), .B(G116), .Z(n1291) );
NAND2_X1 U988 ( .A1(G217), .A2(n1279), .ZN(n1293) );
AND2_X1 U989 ( .A1(G234), .A2(n1100), .ZN(n1279) );
INV_X1 U990 ( .A(G953), .ZN(n1100) );
INV_X1 U991 ( .A(n1208), .ZN(n1249) );
XOR2_X1 U992 ( .A(n1087), .B(G475), .Z(n1208) );
NOR2_X1 U993 ( .A1(n1150), .A2(G902), .ZN(n1087) );
INV_X1 U994 ( .A(n1152), .ZN(n1150) );
XOR2_X1 U995 ( .A(n1294), .B(n1295), .Z(n1152) );
XOR2_X1 U996 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U997 ( .A(G131), .B(G113), .Z(n1297) );
XOR2_X1 U998 ( .A(KEYINPUT10), .B(G146), .Z(n1296) );
XOR2_X1 U999 ( .A(n1298), .B(n1299), .Z(n1294) );
XOR2_X1 U1000 ( .A(n1300), .B(n1287), .Z(n1299) );
XOR2_X1 U1001 ( .A(G122), .B(n1223), .Z(n1287) );
NAND3_X1 U1002 ( .A1(G214), .A2(n1301), .A3(KEYINPUT9), .ZN(n1300) );
XNOR2_X1 U1003 ( .A(G104), .B(n1302), .ZN(n1298) );
NOR2_X1 U1004 ( .A1(KEYINPUT31), .A2(n1109), .ZN(n1302) );
XOR2_X1 U1005 ( .A(n1179), .B(G125), .Z(n1109) );
INV_X1 U1006 ( .A(G140), .ZN(n1179) );
NOR2_X1 U1007 ( .A1(n1050), .A2(n1049), .ZN(n1024) );
INV_X1 U1008 ( .A(n1037), .ZN(n1049) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1280), .ZN(n1037) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1185), .ZN(n1280) );
XOR2_X1 U1011 ( .A(n1303), .B(G469), .Z(n1050) );
NAND4_X1 U1012 ( .A1(n1304), .A2(n1305), .A3(n1306), .A4(n1307), .ZN(n1303) );
OR4_X1 U1013 ( .A1(n1308), .A2(KEYINPUT4), .A3(n1118), .A4(n1309), .ZN(n1307) );
NAND2_X1 U1014 ( .A1(n1309), .A2(n1310), .ZN(n1306) );
NAND3_X1 U1015 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1310) );
NAND2_X1 U1016 ( .A1(KEYINPUT47), .A2(n1308), .ZN(n1313) );
OR3_X1 U1017 ( .A1(n1308), .A2(KEYINPUT47), .A3(n1112), .ZN(n1312) );
NAND2_X1 U1018 ( .A1(n1112), .A2(n1314), .ZN(n1311) );
OR2_X1 U1019 ( .A1(n1308), .A2(KEYINPUT4), .ZN(n1314) );
NAND3_X1 U1020 ( .A1(n1118), .A2(n1315), .A3(n1316), .ZN(n1305) );
XOR2_X1 U1021 ( .A(KEYINPUT47), .B(n1308), .Z(n1316) );
XOR2_X1 U1022 ( .A(n1317), .B(n1176), .Z(n1308) );
NAND2_X1 U1023 ( .A1(n1318), .A2(n1319), .ZN(n1176) );
NAND2_X1 U1024 ( .A1(n1320), .A2(n1019), .ZN(n1319) );
INV_X1 U1025 ( .A(G107), .ZN(n1019) );
XOR2_X1 U1026 ( .A(KEYINPUT41), .B(n1269), .Z(n1320) );
NAND2_X1 U1027 ( .A1(n1269), .A2(G107), .ZN(n1318) );
XOR2_X1 U1028 ( .A(G101), .B(G104), .Z(n1269) );
XOR2_X1 U1029 ( .A(n1113), .B(KEYINPUT38), .Z(n1317) );
NAND2_X1 U1030 ( .A1(n1321), .A2(n1322), .ZN(n1113) );
NAND2_X1 U1031 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1032 ( .A(KEYINPUT62), .B(n1325), .Z(n1321) );
NOR2_X1 U1033 ( .A1(n1324), .A2(n1323), .ZN(n1325) );
XOR2_X1 U1034 ( .A(G143), .B(n1326), .Z(n1323) );
NOR2_X1 U1035 ( .A1(G146), .A2(KEYINPUT15), .ZN(n1326) );
XNOR2_X1 U1036 ( .A(KEYINPUT4), .B(n1309), .ZN(n1315) );
XNOR2_X1 U1037 ( .A(n1171), .B(n1180), .ZN(n1309) );
XOR2_X1 U1038 ( .A(G110), .B(G140), .Z(n1180) );
NOR2_X1 U1039 ( .A1(n1095), .A2(G953), .ZN(n1171) );
INV_X1 U1040 ( .A(G227), .ZN(n1095) );
XOR2_X1 U1041 ( .A(n1185), .B(KEYINPUT45), .Z(n1304) );
XOR2_X1 U1042 ( .A(n1327), .B(G472), .Z(n1042) );
NAND2_X1 U1043 ( .A1(n1328), .A2(n1185), .ZN(n1327) );
INV_X1 U1044 ( .A(G902), .ZN(n1185) );
XOR2_X1 U1045 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1046 ( .A(n1158), .B(n1163), .Z(n1330) );
XNOR2_X1 U1047 ( .A(n1268), .B(KEYINPUT29), .ZN(n1163) );
XNOR2_X1 U1048 ( .A(G113), .B(n1331), .ZN(n1268) );
XOR2_X1 U1049 ( .A(G119), .B(G116), .Z(n1331) );
XOR2_X1 U1050 ( .A(n1221), .B(n1112), .Z(n1158) );
INV_X1 U1051 ( .A(n1118), .ZN(n1112) );
XOR2_X1 U1052 ( .A(n1332), .B(n1290), .Z(n1118) );
XOR2_X1 U1053 ( .A(G134), .B(KEYINPUT6), .Z(n1290) );
XNOR2_X1 U1054 ( .A(G131), .B(G137), .ZN(n1332) );
XOR2_X1 U1055 ( .A(n1324), .B(n1333), .Z(n1221) );
NOR2_X1 U1056 ( .A1(KEYINPUT18), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1057 ( .A(n1223), .B(G146), .Z(n1334) );
INV_X1 U1058 ( .A(G143), .ZN(n1223) );
XNOR2_X1 U1059 ( .A(n1240), .B(KEYINPUT44), .ZN(n1324) );
INV_X1 U1060 ( .A(G128), .ZN(n1240) );
XOR2_X1 U1061 ( .A(KEYINPUT50), .B(n1157), .Z(n1329) );
XOR2_X1 U1062 ( .A(n1335), .B(n1241), .Z(n1157) );
INV_X1 U1063 ( .A(G101), .ZN(n1241) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1301), .ZN(n1335) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1301) );
endmodule


