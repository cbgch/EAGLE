//Key = 0111000011100101001111010101110101001001001101001011011000010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425;

XOR2_X1 U778 ( .A(n1083), .B(n1084), .Z(G9) );
NAND2_X1 U779 ( .A1(KEYINPUT33), .A2(G107), .ZN(n1084) );
NOR2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(G75) );
NOR3_X1 U781 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NAND3_X1 U782 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1087) );
NAND2_X1 U783 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND4_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
OR2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1103), .A2(n1104), .ZN(n1095) );
NAND2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND3_X1 U789 ( .A1(n1099), .A2(n1107), .A3(n1097), .ZN(n1106) );
NAND2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U792 ( .A1(n1098), .A2(n1112), .ZN(n1105) );
NAND2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1097), .A2(n1115), .ZN(n1114) );
OR2_X1 U795 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U796 ( .A1(n1099), .A2(n1118), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U798 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
INV_X1 U799 ( .A(n1123), .ZN(n1093) );
AND3_X1 U800 ( .A1(n1092), .A2(n1124), .A3(n1091), .ZN(n1085) );
NAND2_X1 U801 ( .A1(n1125), .A2(n1126), .ZN(n1091) );
NOR4_X1 U802 ( .A1(n1127), .A2(n1128), .A3(n1110), .A4(n1121), .ZN(n1126) );
XOR2_X1 U803 ( .A(n1129), .B(KEYINPUT40), .Z(n1128) );
NAND3_X1 U804 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
OR3_X1 U805 ( .A1(n1133), .A2(n1134), .A3(KEYINPUT60), .ZN(n1131) );
NAND2_X1 U806 ( .A1(KEYINPUT60), .A2(n1133), .ZN(n1130) );
NAND3_X1 U807 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1127) );
NOR4_X1 U808 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1125) );
XNOR2_X1 U809 ( .A(n1142), .B(n1143), .ZN(n1140) );
NOR2_X1 U810 ( .A1(G475), .A2(KEYINPUT44), .ZN(n1143) );
NAND4_X1 U811 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1138) );
OR3_X1 U812 ( .A1(n1148), .A2(n1149), .A3(KEYINPUT26), .ZN(n1147) );
NAND2_X1 U813 ( .A1(KEYINPUT26), .A2(n1148), .ZN(n1146) );
NAND2_X1 U814 ( .A1(n1150), .A2(n1151), .ZN(n1145) );
INV_X1 U815 ( .A(KEYINPUT52), .ZN(n1151) );
NAND2_X1 U816 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
NAND3_X1 U817 ( .A1(n1153), .A2(n1152), .A3(KEYINPUT52), .ZN(n1144) );
OR3_X1 U818 ( .A1(n1154), .A2(KEYINPUT35), .A3(n1155), .ZN(n1152) );
NAND2_X1 U819 ( .A1(KEYINPUT35), .A2(n1154), .ZN(n1153) );
INV_X1 U820 ( .A(G952), .ZN(n1124) );
XOR2_X1 U821 ( .A(n1156), .B(n1157), .Z(G72) );
XOR2_X1 U822 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U823 ( .A1(G953), .A2(n1160), .ZN(n1159) );
NAND2_X1 U824 ( .A1(G900), .A2(G227), .ZN(n1160) );
NAND2_X1 U825 ( .A1(n1161), .A2(n1162), .ZN(n1158) );
NAND2_X1 U826 ( .A1(G953), .A2(n1163), .ZN(n1162) );
XNOR2_X1 U827 ( .A(n1164), .B(n1165), .ZN(n1161) );
NAND2_X1 U828 ( .A1(n1166), .A2(KEYINPUT45), .ZN(n1164) );
XOR2_X1 U829 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U830 ( .A(G134), .B(G131), .Z(n1168) );
XOR2_X1 U831 ( .A(n1169), .B(n1170), .Z(n1167) );
NOR2_X1 U832 ( .A1(n1171), .A2(n1172), .ZN(n1156) );
NOR2_X1 U833 ( .A1(KEYINPUT37), .A2(n1173), .ZN(n1172) );
INV_X1 U834 ( .A(n1174), .ZN(n1173) );
NOR2_X1 U835 ( .A1(KEYINPUT29), .A2(n1174), .ZN(n1171) );
NAND2_X1 U836 ( .A1(n1175), .A2(n1089), .ZN(n1174) );
NAND2_X1 U837 ( .A1(n1176), .A2(n1177), .ZN(G69) );
NAND2_X1 U838 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U839 ( .A1(G953), .A2(n1180), .ZN(n1179) );
NAND3_X1 U840 ( .A1(n1181), .A2(n1182), .A3(G953), .ZN(n1176) );
NAND2_X1 U841 ( .A1(G898), .A2(G224), .ZN(n1182) );
XOR2_X1 U842 ( .A(KEYINPUT43), .B(n1178), .Z(n1181) );
XNOR2_X1 U843 ( .A(n1183), .B(n1184), .ZN(n1178) );
NOR3_X1 U844 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NOR2_X1 U845 ( .A1(KEYINPUT22), .A2(n1188), .ZN(n1187) );
NOR2_X1 U846 ( .A1(n1189), .A2(n1190), .ZN(n1186) );
INV_X1 U847 ( .A(KEYINPUT22), .ZN(n1190) );
NOR2_X1 U848 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NAND2_X1 U849 ( .A1(n1175), .A2(n1088), .ZN(n1183) );
NOR2_X1 U850 ( .A1(n1193), .A2(n1194), .ZN(G66) );
XOR2_X1 U851 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U852 ( .A1(n1133), .A2(n1197), .ZN(n1195) );
NOR2_X1 U853 ( .A1(n1193), .A2(n1198), .ZN(G63) );
XOR2_X1 U854 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U855 ( .A1(n1148), .A2(n1197), .ZN(n1199) );
NOR2_X1 U856 ( .A1(n1193), .A2(n1201), .ZN(G60) );
NOR3_X1 U857 ( .A1(n1142), .A2(n1202), .A3(n1203), .ZN(n1201) );
NOR3_X1 U858 ( .A1(n1204), .A2(n1205), .A3(n1197), .ZN(n1203) );
INV_X1 U859 ( .A(n1206), .ZN(n1204) );
NOR2_X1 U860 ( .A1(n1207), .A2(n1206), .ZN(n1202) );
NOR2_X1 U861 ( .A1(n1208), .A2(n1205), .ZN(n1207) );
INV_X1 U862 ( .A(G475), .ZN(n1205) );
NOR2_X1 U863 ( .A1(n1088), .A2(n1089), .ZN(n1208) );
XNOR2_X1 U864 ( .A(G104), .B(n1209), .ZN(G6) );
NAND4_X1 U865 ( .A1(n1210), .A2(n1101), .A3(n1211), .A4(n1212), .ZN(n1209) );
NOR2_X1 U866 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
XOR2_X1 U867 ( .A(n1119), .B(KEYINPUT7), .Z(n1214) );
XOR2_X1 U868 ( .A(n1215), .B(KEYINPUT21), .Z(n1210) );
NOR3_X1 U869 ( .A1(n1193), .A2(n1216), .A3(n1217), .ZN(G57) );
NOR3_X1 U870 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
AND2_X1 U871 ( .A1(KEYINPUT9), .A2(n1221), .ZN(n1220) );
NOR2_X1 U872 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
AND2_X1 U873 ( .A1(n1224), .A2(KEYINPUT9), .ZN(n1222) );
INV_X1 U874 ( .A(n1225), .ZN(n1218) );
NOR2_X1 U875 ( .A1(n1226), .A2(n1225), .ZN(n1216) );
XOR2_X1 U876 ( .A(n1227), .B(n1228), .Z(n1225) );
NOR2_X1 U877 ( .A1(n1221), .A2(n1229), .ZN(n1226) );
NOR2_X1 U878 ( .A1(n1224), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U879 ( .A(KEYINPUT9), .B(n1223), .ZN(n1230) );
AND2_X1 U880 ( .A1(n1224), .A2(n1223), .ZN(n1221) );
XNOR2_X1 U881 ( .A(n1231), .B(n1232), .ZN(n1223) );
NOR2_X1 U882 ( .A1(n1233), .A2(n1197), .ZN(n1232) );
INV_X1 U883 ( .A(G472), .ZN(n1233) );
NAND2_X1 U884 ( .A1(n1234), .A2(n1235), .ZN(n1231) );
NAND2_X1 U885 ( .A1(n1236), .A2(G101), .ZN(n1235) );
XOR2_X1 U886 ( .A(KEYINPUT1), .B(n1237), .Z(n1234) );
NOR2_X1 U887 ( .A1(n1236), .A2(G101), .ZN(n1237) );
INV_X1 U888 ( .A(n1238), .ZN(n1236) );
XNOR2_X1 U889 ( .A(n1239), .B(n1240), .ZN(n1224) );
NAND2_X1 U890 ( .A1(KEYINPUT15), .A2(n1241), .ZN(n1239) );
NOR3_X1 U891 ( .A1(n1193), .A2(n1242), .A3(n1243), .ZN(G54) );
NOR4_X1 U892 ( .A1(n1244), .A2(n1197), .A3(KEYINPUT4), .A4(n1155), .ZN(n1243) );
INV_X1 U893 ( .A(n1245), .ZN(n1244) );
NOR2_X1 U894 ( .A1(n1245), .A2(n1246), .ZN(n1242) );
NOR3_X1 U895 ( .A1(n1197), .A2(n1247), .A3(n1155), .ZN(n1246) );
AND2_X1 U896 ( .A1(n1248), .A2(KEYINPUT4), .ZN(n1247) );
NOR2_X1 U897 ( .A1(KEYINPUT32), .A2(n1248), .ZN(n1245) );
XNOR2_X1 U898 ( .A(n1249), .B(n1250), .ZN(n1248) );
NOR2_X1 U899 ( .A1(n1193), .A2(n1251), .ZN(G51) );
XOR2_X1 U900 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U901 ( .A(n1254), .B(n1255), .Z(n1253) );
NOR3_X1 U902 ( .A1(n1197), .A2(KEYINPUT55), .A3(n1256), .ZN(n1255) );
NAND2_X1 U903 ( .A1(G902), .A2(n1257), .ZN(n1197) );
OR2_X1 U904 ( .A1(n1089), .A2(n1088), .ZN(n1257) );
NAND4_X1 U905 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1088) );
AND4_X1 U906 ( .A1(n1262), .A2(n1263), .A3(n1083), .A4(n1264), .ZN(n1261) );
NAND3_X1 U907 ( .A1(n1102), .A2(n1099), .A3(n1265), .ZN(n1083) );
NOR3_X1 U908 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1260) );
NOR2_X1 U909 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
INV_X1 U910 ( .A(KEYINPUT8), .ZN(n1269) );
NOR2_X1 U911 ( .A1(KEYINPUT8), .A2(n1271), .ZN(n1267) );
NAND4_X1 U912 ( .A1(n1213), .A2(n1103), .A3(n1272), .A4(n1098), .ZN(n1271) );
NOR2_X1 U913 ( .A1(n1119), .A2(n1273), .ZN(n1266) );
NAND3_X1 U914 ( .A1(n1265), .A2(n1099), .A3(n1101), .ZN(n1258) );
NAND4_X1 U915 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1089) );
AND4_X1 U916 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1277) );
NOR3_X1 U917 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n1276) );
NOR4_X1 U918 ( .A1(n1285), .A2(n1286), .A3(n1101), .A4(n1287), .ZN(n1284) );
INV_X1 U919 ( .A(n1288), .ZN(n1286) );
AND2_X1 U920 ( .A1(n1285), .A2(n1289), .ZN(n1283) );
INV_X1 U921 ( .A(KEYINPUT49), .ZN(n1285) );
AND2_X1 U922 ( .A1(n1290), .A2(KEYINPUT2), .ZN(n1282) );
NAND3_X1 U923 ( .A1(n1291), .A2(n1292), .A3(n1097), .ZN(n1274) );
NAND2_X1 U924 ( .A1(n1293), .A2(n1294), .ZN(n1291) );
NAND3_X1 U925 ( .A1(n1108), .A2(n1101), .A3(n1295), .ZN(n1294) );
NOR3_X1 U926 ( .A1(n1139), .A2(KEYINPUT2), .A3(n1296), .ZN(n1295) );
NOR2_X1 U927 ( .A1(n1297), .A2(n1298), .ZN(n1254) );
XOR2_X1 U928 ( .A(n1299), .B(KEYINPUT59), .Z(n1298) );
NAND2_X1 U929 ( .A1(G125), .A2(n1241), .ZN(n1299) );
NOR2_X1 U930 ( .A1(G125), .A2(n1241), .ZN(n1297) );
NOR2_X1 U931 ( .A1(n1175), .A2(G952), .ZN(n1193) );
XOR2_X1 U932 ( .A(n1300), .B(n1289), .Z(G48) );
AND3_X1 U933 ( .A1(n1272), .A2(n1101), .A3(n1288), .ZN(n1289) );
NOR2_X1 U934 ( .A1(KEYINPUT41), .A2(n1301), .ZN(n1300) );
XNOR2_X1 U935 ( .A(G146), .B(KEYINPUT34), .ZN(n1301) );
XOR2_X1 U936 ( .A(n1302), .B(n1275), .Z(G45) );
NAND3_X1 U937 ( .A1(n1116), .A2(n1288), .A3(n1303), .ZN(n1275) );
NOR3_X1 U938 ( .A1(n1304), .A2(n1305), .A3(n1119), .ZN(n1303) );
INV_X1 U939 ( .A(n1306), .ZN(n1119) );
XOR2_X1 U940 ( .A(G140), .B(n1290), .Z(G42) );
AND2_X1 U941 ( .A1(n1307), .A2(n1117), .ZN(n1290) );
XOR2_X1 U942 ( .A(G137), .B(n1308), .Z(G39) );
NOR4_X1 U943 ( .A1(KEYINPUT62), .A2(n1309), .A3(n1293), .A4(n1310), .ZN(n1308) );
XOR2_X1 U944 ( .A(KEYINPUT23), .B(n1097), .Z(n1310) );
NAND3_X1 U945 ( .A1(n1288), .A2(n1139), .A3(n1103), .ZN(n1293) );
XOR2_X1 U946 ( .A(n1281), .B(n1311), .Z(G36) );
XOR2_X1 U947 ( .A(KEYINPUT53), .B(G134), .Z(n1311) );
NAND4_X1 U948 ( .A1(n1116), .A2(n1097), .A3(n1288), .A4(n1102), .ZN(n1281) );
XOR2_X1 U949 ( .A(n1312), .B(n1280), .Z(G33) );
NAND2_X1 U950 ( .A1(n1116), .A2(n1307), .ZN(n1280) );
AND3_X1 U951 ( .A1(n1288), .A2(n1101), .A3(n1097), .ZN(n1307) );
AND2_X1 U952 ( .A1(n1122), .A2(n1313), .ZN(n1097) );
NOR2_X1 U953 ( .A1(n1108), .A2(n1296), .ZN(n1288) );
INV_X1 U954 ( .A(n1314), .ZN(n1296) );
XNOR2_X1 U955 ( .A(n1212), .B(KEYINPUT16), .ZN(n1108) );
XOR2_X1 U956 ( .A(n1279), .B(n1315), .Z(G30) );
XOR2_X1 U957 ( .A(n1316), .B(KEYINPUT56), .Z(n1315) );
NAND4_X1 U958 ( .A1(n1272), .A2(n1102), .A3(n1212), .A4(n1314), .ZN(n1279) );
XNOR2_X1 U959 ( .A(G101), .B(n1259), .ZN(G3) );
NAND3_X1 U960 ( .A1(n1116), .A2(n1265), .A3(n1103), .ZN(n1259) );
XOR2_X1 U961 ( .A(n1317), .B(n1278), .Z(G27) );
NAND4_X1 U962 ( .A1(n1306), .A2(n1314), .A3(n1117), .A4(n1318), .ZN(n1278) );
AND2_X1 U963 ( .A1(n1101), .A2(n1098), .ZN(n1318) );
NAND2_X1 U964 ( .A1(n1123), .A2(n1319), .ZN(n1314) );
NAND4_X1 U965 ( .A1(G902), .A2(G953), .A3(n1320), .A4(n1163), .ZN(n1319) );
INV_X1 U966 ( .A(G900), .ZN(n1163) );
XOR2_X1 U967 ( .A(n1321), .B(n1322), .Z(G24) );
NAND2_X1 U968 ( .A1(n1323), .A2(n1306), .ZN(n1322) );
XOR2_X1 U969 ( .A(n1273), .B(KEYINPUT36), .Z(n1323) );
NAND3_X1 U970 ( .A1(n1324), .A2(n1098), .A3(n1325), .ZN(n1273) );
NOR3_X1 U971 ( .A1(n1215), .A2(n1213), .A3(n1305), .ZN(n1325) );
INV_X1 U972 ( .A(n1326), .ZN(n1213) );
INV_X1 U973 ( .A(n1099), .ZN(n1215) );
NOR2_X1 U974 ( .A1(n1292), .A2(n1139), .ZN(n1099) );
INV_X1 U975 ( .A(n1304), .ZN(n1324) );
XNOR2_X1 U976 ( .A(G119), .B(n1270), .ZN(G21) );
NAND4_X1 U977 ( .A1(n1103), .A2(n1272), .A3(n1098), .A4(n1326), .ZN(n1270) );
INV_X1 U978 ( .A(n1287), .ZN(n1272) );
NAND3_X1 U979 ( .A1(n1139), .A2(n1292), .A3(n1306), .ZN(n1287) );
XOR2_X1 U980 ( .A(n1327), .B(n1263), .Z(G18) );
NAND2_X1 U981 ( .A1(n1328), .A2(n1102), .ZN(n1263) );
NOR2_X1 U982 ( .A1(n1329), .A2(n1305), .ZN(n1102) );
XOR2_X1 U983 ( .A(n1330), .B(KEYINPUT48), .Z(n1305) );
XOR2_X1 U984 ( .A(n1262), .B(n1331), .Z(G15) );
XOR2_X1 U985 ( .A(KEYINPUT42), .B(G113), .Z(n1331) );
NAND2_X1 U986 ( .A1(n1328), .A2(n1101), .ZN(n1262) );
NOR2_X1 U987 ( .A1(n1304), .A2(n1330), .ZN(n1101) );
XOR2_X1 U988 ( .A(n1329), .B(KEYINPUT28), .Z(n1304) );
AND4_X1 U989 ( .A1(n1116), .A2(n1098), .A3(n1306), .A4(n1326), .ZN(n1328) );
NOR2_X1 U990 ( .A1(n1332), .A2(n1110), .ZN(n1098) );
AND2_X1 U991 ( .A1(n1309), .A2(n1139), .ZN(n1116) );
XOR2_X1 U992 ( .A(n1333), .B(n1264), .Z(G12) );
NAND3_X1 U993 ( .A1(n1117), .A2(n1265), .A3(n1103), .ZN(n1264) );
NOR2_X1 U994 ( .A1(n1329), .A2(n1330), .ZN(n1103) );
NAND2_X1 U995 ( .A1(n1334), .A2(n1136), .ZN(n1330) );
NAND2_X1 U996 ( .A1(n1149), .A2(n1148), .ZN(n1136) );
OR2_X1 U997 ( .A1(n1148), .A2(n1149), .ZN(n1334) );
NOR2_X1 U998 ( .A1(n1200), .A2(G902), .ZN(n1149) );
XNOR2_X1 U999 ( .A(n1335), .B(n1336), .ZN(n1200) );
NOR2_X1 U1000 ( .A1(KEYINPUT30), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1001 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1002 ( .A(G128), .B(n1340), .Z(n1339) );
XOR2_X1 U1003 ( .A(G143), .B(G134), .Z(n1340) );
XOR2_X1 U1004 ( .A(n1341), .B(G107), .Z(n1338) );
NAND2_X1 U1005 ( .A1(n1342), .A2(KEYINPUT25), .ZN(n1341) );
XOR2_X1 U1006 ( .A(n1327), .B(G122), .Z(n1342) );
NAND3_X1 U1007 ( .A1(G234), .A2(n1175), .A3(n1343), .ZN(n1335) );
XNOR2_X1 U1008 ( .A(G217), .B(KEYINPUT20), .ZN(n1343) );
INV_X1 U1009 ( .A(G478), .ZN(n1148) );
XOR2_X1 U1010 ( .A(n1142), .B(G475), .Z(n1329) );
NOR2_X1 U1011 ( .A1(n1206), .A2(G902), .ZN(n1142) );
XOR2_X1 U1012 ( .A(n1344), .B(n1345), .Z(n1206) );
XOR2_X1 U1013 ( .A(G104), .B(n1346), .Z(n1345) );
XOR2_X1 U1014 ( .A(G122), .B(G113), .Z(n1346) );
XNOR2_X1 U1015 ( .A(n1347), .B(n1348), .ZN(n1344) );
XOR2_X1 U1016 ( .A(n1349), .B(n1350), .Z(n1347) );
NOR2_X1 U1017 ( .A1(n1351), .A2(KEYINPUT17), .ZN(n1350) );
NOR2_X1 U1018 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1019 ( .A(n1354), .B(KEYINPUT63), .Z(n1353) );
NAND2_X1 U1020 ( .A1(G125), .A2(n1355), .ZN(n1354) );
NOR2_X1 U1021 ( .A1(G125), .A2(n1355), .ZN(n1352) );
NAND2_X1 U1022 ( .A1(n1356), .A2(n1357), .ZN(n1349) );
NAND2_X1 U1023 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1024 ( .A(KEYINPUT19), .B(n1360), .Z(n1356) );
NOR2_X1 U1025 ( .A1(n1359), .A2(n1361), .ZN(n1360) );
XNOR2_X1 U1026 ( .A(KEYINPUT18), .B(n1358), .ZN(n1361) );
XNOR2_X1 U1027 ( .A(G131), .B(KEYINPUT11), .ZN(n1358) );
XOR2_X1 U1028 ( .A(n1302), .B(n1362), .Z(n1359) );
NAND3_X1 U1029 ( .A1(n1363), .A2(n1175), .A3(n1364), .ZN(n1362) );
XOR2_X1 U1030 ( .A(KEYINPUT5), .B(G214), .Z(n1364) );
AND3_X1 U1031 ( .A1(n1306), .A2(n1326), .A3(n1212), .ZN(n1265) );
NOR2_X1 U1032 ( .A1(n1111), .A2(n1110), .ZN(n1212) );
AND2_X1 U1033 ( .A1(G221), .A2(n1365), .ZN(n1110) );
INV_X1 U1034 ( .A(n1332), .ZN(n1111) );
NAND2_X1 U1035 ( .A1(n1137), .A2(n1366), .ZN(n1332) );
NAND2_X1 U1036 ( .A1(G469), .A2(n1367), .ZN(n1366) );
NAND2_X1 U1037 ( .A1(n1154), .A2(n1155), .ZN(n1137) );
INV_X1 U1038 ( .A(G469), .ZN(n1155) );
INV_X1 U1039 ( .A(n1367), .ZN(n1154) );
NAND2_X1 U1040 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
XOR2_X1 U1041 ( .A(n1370), .B(n1371), .Z(n1368) );
INV_X1 U1042 ( .A(n1249), .ZN(n1371) );
XOR2_X1 U1043 ( .A(n1372), .B(n1373), .Z(n1249) );
XOR2_X1 U1044 ( .A(n1374), .B(n1375), .Z(n1373) );
XOR2_X1 U1045 ( .A(n1376), .B(n1377), .Z(n1375) );
AND2_X1 U1046 ( .A1(n1175), .A2(G227), .ZN(n1377) );
NOR2_X1 U1047 ( .A1(KEYINPUT6), .A2(n1378), .ZN(n1376) );
INV_X1 U1048 ( .A(G107), .ZN(n1378) );
XOR2_X1 U1049 ( .A(n1379), .B(n1380), .Z(n1372) );
XOR2_X1 U1050 ( .A(G128), .B(G104), .Z(n1380) );
XOR2_X1 U1051 ( .A(n1240), .B(G101), .Z(n1379) );
NAND2_X1 U1052 ( .A1(KEYINPUT10), .A2(n1250), .ZN(n1370) );
XOR2_X1 U1053 ( .A(G110), .B(G140), .Z(n1250) );
NAND2_X1 U1054 ( .A1(n1123), .A2(n1381), .ZN(n1326) );
NAND3_X1 U1055 ( .A1(n1185), .A2(n1320), .A3(G902), .ZN(n1381) );
NOR2_X1 U1056 ( .A1(n1175), .A2(G898), .ZN(n1185) );
NAND3_X1 U1057 ( .A1(n1092), .A2(n1320), .A3(G952), .ZN(n1123) );
NAND2_X1 U1058 ( .A1(G237), .A2(G234), .ZN(n1320) );
XNOR2_X1 U1059 ( .A(G953), .B(KEYINPUT24), .ZN(n1092) );
NOR2_X1 U1060 ( .A1(n1122), .A2(n1121), .ZN(n1306) );
INV_X1 U1061 ( .A(n1313), .ZN(n1121) );
NAND2_X1 U1062 ( .A1(G214), .A2(n1382), .ZN(n1313) );
NAND2_X1 U1063 ( .A1(n1363), .A2(n1369), .ZN(n1382) );
NOR2_X1 U1064 ( .A1(n1383), .A2(n1141), .ZN(n1122) );
NAND2_X1 U1065 ( .A1(n1384), .A2(n1385), .ZN(n1141) );
NAND2_X1 U1066 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
NAND2_X1 U1067 ( .A1(G210), .A2(G902), .ZN(n1384) );
XNOR2_X1 U1068 ( .A(n1135), .B(KEYINPUT46), .ZN(n1383) );
OR3_X1 U1069 ( .A1(n1386), .A2(G902), .A3(n1387), .ZN(n1135) );
XNOR2_X1 U1070 ( .A(n1388), .B(n1252), .ZN(n1387) );
XNOR2_X1 U1071 ( .A(n1188), .B(n1389), .ZN(n1252) );
NOR2_X1 U1072 ( .A1(G953), .A2(n1180), .ZN(n1389) );
INV_X1 U1073 ( .A(G224), .ZN(n1180) );
XOR2_X1 U1074 ( .A(n1192), .B(n1191), .Z(n1188) );
AND2_X1 U1075 ( .A1(n1390), .A2(n1391), .ZN(n1191) );
NAND2_X1 U1076 ( .A1(G122), .A2(n1333), .ZN(n1391) );
XOR2_X1 U1077 ( .A(n1392), .B(KEYINPUT14), .Z(n1390) );
NAND2_X1 U1078 ( .A1(n1393), .A2(n1321), .ZN(n1392) );
INV_X1 U1079 ( .A(G122), .ZN(n1321) );
XOR2_X1 U1080 ( .A(KEYINPUT61), .B(G110), .Z(n1393) );
XOR2_X1 U1081 ( .A(n1394), .B(n1395), .Z(n1192) );
XOR2_X1 U1082 ( .A(G116), .B(G107), .Z(n1395) );
XOR2_X1 U1083 ( .A(n1396), .B(n1397), .Z(n1394) );
NOR2_X1 U1084 ( .A1(G104), .A2(KEYINPUT47), .ZN(n1397) );
XOR2_X1 U1085 ( .A(n1398), .B(G125), .Z(n1388) );
NAND2_X1 U1086 ( .A1(KEYINPUT54), .A2(n1241), .ZN(n1398) );
NOR2_X1 U1087 ( .A1(n1256), .A2(n1363), .ZN(n1386) );
INV_X1 U1088 ( .A(G210), .ZN(n1256) );
NOR2_X1 U1089 ( .A1(n1139), .A2(n1309), .ZN(n1117) );
INV_X1 U1090 ( .A(n1292), .ZN(n1309) );
NAND3_X1 U1091 ( .A1(n1399), .A2(n1400), .A3(n1132), .ZN(n1292) );
NAND2_X1 U1092 ( .A1(n1134), .A2(n1133), .ZN(n1132) );
OR3_X1 U1093 ( .A1(n1133), .A2(n1134), .A3(KEYINPUT58), .ZN(n1400) );
NOR2_X1 U1094 ( .A1(n1196), .A2(G902), .ZN(n1134) );
XNOR2_X1 U1095 ( .A(n1401), .B(n1402), .ZN(n1196) );
XNOR2_X1 U1096 ( .A(n1403), .B(n1170), .ZN(n1402) );
XOR2_X1 U1097 ( .A(G137), .B(G128), .Z(n1170) );
NAND4_X1 U1098 ( .A1(KEYINPUT31), .A2(G221), .A3(G234), .A4(n1175), .ZN(n1403) );
XOR2_X1 U1099 ( .A(n1404), .B(n1405), .Z(n1401) );
XOR2_X1 U1100 ( .A(G119), .B(G110), .Z(n1405) );
NAND3_X1 U1101 ( .A1(n1406), .A2(n1407), .A3(n1408), .ZN(n1404) );
NAND2_X1 U1102 ( .A1(n1348), .A2(n1409), .ZN(n1408) );
OR3_X1 U1103 ( .A1(n1409), .A2(n1348), .A3(KEYINPUT12), .ZN(n1407) );
NAND2_X1 U1104 ( .A1(KEYINPUT27), .A2(n1410), .ZN(n1409) );
INV_X1 U1105 ( .A(n1165), .ZN(n1410) );
NAND2_X1 U1106 ( .A1(KEYINPUT12), .A2(n1165), .ZN(n1406) );
XNOR2_X1 U1107 ( .A(n1355), .B(n1317), .ZN(n1165) );
INV_X1 U1108 ( .A(G125), .ZN(n1317) );
INV_X1 U1109 ( .A(G140), .ZN(n1355) );
NAND2_X1 U1110 ( .A1(KEYINPUT58), .A2(n1133), .ZN(n1399) );
NAND2_X1 U1111 ( .A1(G217), .A2(n1365), .ZN(n1133) );
NAND2_X1 U1112 ( .A1(G234), .A2(n1369), .ZN(n1365) );
XNOR2_X1 U1113 ( .A(n1411), .B(G472), .ZN(n1139) );
NAND2_X1 U1114 ( .A1(n1412), .A2(n1369), .ZN(n1411) );
INV_X1 U1115 ( .A(G902), .ZN(n1369) );
XOR2_X1 U1116 ( .A(n1413), .B(n1414), .Z(n1412) );
XOR2_X1 U1117 ( .A(n1227), .B(n1415), .Z(n1414) );
XNOR2_X1 U1118 ( .A(KEYINPUT38), .B(n1416), .ZN(n1415) );
NOR2_X1 U1119 ( .A1(KEYINPUT57), .A2(n1240), .ZN(n1416) );
NAND3_X1 U1120 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n1240) );
NAND2_X1 U1121 ( .A1(n1420), .A2(n1312), .ZN(n1419) );
INV_X1 U1122 ( .A(G131), .ZN(n1312) );
NAND2_X1 U1123 ( .A1(n1421), .A2(KEYINPUT39), .ZN(n1420) );
XNOR2_X1 U1124 ( .A(n1422), .B(KEYINPUT3), .ZN(n1421) );
NAND3_X1 U1125 ( .A1(KEYINPUT39), .A2(G131), .A3(n1422), .ZN(n1418) );
OR2_X1 U1126 ( .A1(n1422), .A2(KEYINPUT39), .ZN(n1417) );
XOR2_X1 U1127 ( .A(G137), .B(G134), .Z(n1422) );
NAND2_X1 U1128 ( .A1(KEYINPUT51), .A2(n1327), .ZN(n1227) );
INV_X1 U1129 ( .A(G116), .ZN(n1327) );
XNOR2_X1 U1130 ( .A(n1423), .B(n1241), .ZN(n1413) );
XNOR2_X1 U1131 ( .A(n1424), .B(n1169), .ZN(n1241) );
INV_X1 U1132 ( .A(n1374), .ZN(n1169) );
XOR2_X1 U1133 ( .A(n1302), .B(n1348), .Z(n1374) );
XNOR2_X1 U1134 ( .A(G146), .B(KEYINPUT50), .ZN(n1348) );
INV_X1 U1135 ( .A(G143), .ZN(n1302) );
NAND2_X1 U1136 ( .A1(KEYINPUT13), .A2(n1316), .ZN(n1424) );
INV_X1 U1137 ( .A(G128), .ZN(n1316) );
XOR2_X1 U1138 ( .A(n1396), .B(n1425), .Z(n1423) );
NOR2_X1 U1139 ( .A1(KEYINPUT0), .A2(n1238), .ZN(n1425) );
NAND3_X1 U1140 ( .A1(n1363), .A2(n1175), .A3(G210), .ZN(n1238) );
INV_X1 U1141 ( .A(G953), .ZN(n1175) );
INV_X1 U1142 ( .A(G237), .ZN(n1363) );
XNOR2_X1 U1143 ( .A(G101), .B(n1228), .ZN(n1396) );
XOR2_X1 U1144 ( .A(G113), .B(G119), .Z(n1228) );
INV_X1 U1145 ( .A(G110), .ZN(n1333) );
endmodule


