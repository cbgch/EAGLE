//Key = 1110100110110100010100000100011111110011001011000111110111101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;

XOR2_X1 U761 ( .A(G107), .B(n1055), .Z(G9) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(G75) );
NOR4_X1 U763 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR4_X1 U765 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1062) );
NAND4_X1 U766 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1064) );
NAND3_X1 U767 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1058) );
NAND2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND4_X1 U770 ( .A1(n1069), .A2(n1079), .A3(n1071), .A4(n1080), .ZN(n1078) );
NAND2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U775 ( .A1(n1070), .A2(n1089), .ZN(n1081) );
NAND2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND3_X1 U777 ( .A1(n1068), .A2(n1063), .A3(n1092), .ZN(n1091) );
INV_X1 U778 ( .A(KEYINPUT28), .ZN(n1063) );
INV_X1 U779 ( .A(n1093), .ZN(n1090) );
NAND3_X1 U780 ( .A1(n1070), .A2(n1094), .A3(n1083), .ZN(n1077) );
NAND2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND3_X1 U782 ( .A1(n1069), .A2(n1097), .A3(n1079), .ZN(n1096) );
NAND3_X1 U783 ( .A1(n1098), .A2(n1099), .A3(n1071), .ZN(n1095) );
NAND2_X1 U784 ( .A1(n1100), .A2(n1066), .ZN(n1099) );
NAND3_X1 U785 ( .A1(n1101), .A2(n1102), .A3(n1069), .ZN(n1098) );
INV_X1 U786 ( .A(n1065), .ZN(n1075) );
AND3_X1 U787 ( .A1(n1072), .A2(n1073), .A3(n1103), .ZN(n1056) );
NAND4_X1 U788 ( .A1(n1104), .A2(n1070), .A3(n1105), .A4(n1106), .ZN(n1072) );
NOR4_X1 U789 ( .A1(n1097), .A2(n1092), .A3(n1107), .A4(n1108), .ZN(n1106) );
XNOR2_X1 U790 ( .A(n1100), .B(KEYINPUT13), .ZN(n1108) );
XOR2_X1 U791 ( .A(n1109), .B(n1110), .Z(n1107) );
XOR2_X1 U792 ( .A(KEYINPUT44), .B(KEYINPUT15), .Z(n1110) );
XNOR2_X1 U793 ( .A(G478), .B(n1111), .ZN(n1109) );
XNOR2_X1 U794 ( .A(n1112), .B(n1113), .ZN(n1105) );
XOR2_X1 U795 ( .A(n1114), .B(n1115), .Z(G72) );
AND2_X1 U796 ( .A1(n1059), .A2(n1073), .ZN(n1115) );
NAND2_X1 U797 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NAND2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U799 ( .A1(G953), .A2(n1120), .ZN(n1119) );
INV_X1 U800 ( .A(n1121), .ZN(n1118) );
NAND3_X1 U801 ( .A1(G953), .A2(n1122), .A3(n1121), .ZN(n1116) );
NAND3_X1 U802 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1121) );
NAND2_X1 U803 ( .A1(G953), .A2(n1126), .ZN(n1125) );
NAND2_X1 U804 ( .A1(n1127), .A2(n1128), .ZN(n1124) );
NAND2_X1 U805 ( .A1(KEYINPUT32), .A2(n1129), .ZN(n1128) );
XOR2_X1 U806 ( .A(n1130), .B(n1131), .Z(n1127) );
NOR2_X1 U807 ( .A1(G140), .A2(KEYINPUT20), .ZN(n1131) );
NAND3_X1 U808 ( .A1(n1132), .A2(n1129), .A3(KEYINPUT32), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1130), .B(n1133), .Z(n1132) );
NOR2_X1 U810 ( .A1(KEYINPUT20), .A2(n1134), .ZN(n1133) );
NAND2_X1 U811 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
NAND2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U813 ( .A(KEYINPUT24), .B(n1139), .ZN(n1137) );
NAND2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(n1135) );
XOR2_X1 U815 ( .A(n1139), .B(KEYINPUT59), .Z(n1140) );
NAND2_X1 U816 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
NAND2_X1 U817 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U818 ( .A(KEYINPUT49), .B(n1146), .Z(n1144) );
NAND2_X1 U819 ( .A1(n1146), .A2(G137), .ZN(n1142) );
NAND2_X1 U820 ( .A1(G900), .A2(G227), .ZN(n1122) );
XOR2_X1 U821 ( .A(n1147), .B(n1148), .Z(G69) );
NAND2_X1 U822 ( .A1(G953), .A2(n1149), .ZN(n1148) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1149) );
NAND3_X1 U824 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1147) );
XOR2_X1 U825 ( .A(KEYINPUT43), .B(KEYINPUT17), .Z(n1152) );
NAND2_X1 U826 ( .A1(KEYINPUT34), .A2(n1153), .ZN(n1151) );
NAND2_X1 U827 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U828 ( .A1(G953), .A2(n1156), .ZN(n1155) );
XNOR2_X1 U829 ( .A(n1061), .B(n1157), .ZN(n1154) );
NAND4_X1 U830 ( .A1(n1061), .A2(n1073), .A3(n1157), .A4(n1158), .ZN(n1150) );
INV_X1 U831 ( .A(KEYINPUT34), .ZN(n1158) );
XOR2_X1 U832 ( .A(n1159), .B(n1160), .Z(n1157) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U834 ( .A1(KEYINPUT38), .A2(n1163), .ZN(n1162) );
XNOR2_X1 U835 ( .A(KEYINPUT46), .B(n1164), .ZN(n1163) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(G66) );
XNOR2_X1 U837 ( .A(n1167), .B(n1168), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U839 ( .A1(n1165), .A2(n1171), .ZN(G63) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U841 ( .A(n1174), .B(KEYINPUT19), .Z(n1173) );
NAND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U843 ( .A1(n1175), .A2(n1176), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1170), .A2(n1177), .ZN(n1175) );
NOR3_X1 U845 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(G60) );
NOR3_X1 U846 ( .A1(n1181), .A2(n1073), .A3(n1103), .ZN(n1180) );
INV_X1 U847 ( .A(G952), .ZN(n1103) );
AND2_X1 U848 ( .A1(n1181), .A2(n1165), .ZN(n1179) );
INV_X1 U849 ( .A(KEYINPUT41), .ZN(n1181) );
XOR2_X1 U850 ( .A(n1182), .B(n1183), .Z(n1178) );
AND2_X1 U851 ( .A1(G475), .A2(n1184), .ZN(n1182) );
XOR2_X1 U852 ( .A(G104), .B(n1185), .Z(G6) );
NOR3_X1 U853 ( .A1(n1101), .A2(n1186), .A3(n1187), .ZN(n1185) );
NOR2_X1 U854 ( .A1(n1165), .A2(n1188), .ZN(G57) );
XOR2_X1 U855 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U856 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U857 ( .A(KEYINPUT36), .B(n1193), .Z(n1192) );
AND2_X1 U858 ( .A1(G472), .A2(n1184), .ZN(n1193) );
NOR2_X1 U859 ( .A1(n1194), .A2(n1195), .ZN(n1191) );
XOR2_X1 U860 ( .A(KEYINPUT26), .B(n1196), .Z(n1195) );
NOR2_X1 U861 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U862 ( .A1(n1199), .A2(n1200), .ZN(n1194) );
XNOR2_X1 U863 ( .A(n1201), .B(n1202), .ZN(n1189) );
NOR2_X1 U864 ( .A1(n1165), .A2(n1203), .ZN(G54) );
XOR2_X1 U865 ( .A(n1204), .B(n1205), .Z(n1203) );
XNOR2_X1 U866 ( .A(n1199), .B(n1206), .ZN(n1205) );
XNOR2_X1 U867 ( .A(n1207), .B(n1208), .ZN(n1206) );
NOR2_X1 U868 ( .A1(KEYINPUT37), .A2(n1209), .ZN(n1208) );
XOR2_X1 U869 ( .A(n1210), .B(n1211), .Z(n1209) );
XNOR2_X1 U870 ( .A(n1134), .B(G110), .ZN(n1211) );
INV_X1 U871 ( .A(G140), .ZN(n1134) );
NAND2_X1 U872 ( .A1(KEYINPUT31), .A2(n1212), .ZN(n1207) );
NAND2_X1 U873 ( .A1(n1184), .A2(G469), .ZN(n1212) );
INV_X1 U874 ( .A(n1170), .ZN(n1184) );
XNOR2_X1 U875 ( .A(n1213), .B(n1138), .ZN(n1204) );
NOR2_X1 U876 ( .A1(n1165), .A2(n1214), .ZN(G51) );
XOR2_X1 U877 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U878 ( .A(n1217), .B(n1218), .ZN(n1216) );
NOR3_X1 U879 ( .A1(n1170), .A2(KEYINPUT62), .A3(n1113), .ZN(n1218) );
NAND2_X1 U880 ( .A1(G902), .A2(n1219), .ZN(n1170) );
OR2_X1 U881 ( .A1(n1059), .A2(n1061), .ZN(n1219) );
NAND2_X1 U882 ( .A1(n1220), .A2(n1221), .ZN(n1061) );
NOR4_X1 U883 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
NOR4_X1 U884 ( .A1(n1226), .A2(n1055), .A3(n1227), .A4(n1228), .ZN(n1220) );
NOR3_X1 U885 ( .A1(n1101), .A2(n1229), .A3(n1187), .ZN(n1227) );
XNOR2_X1 U886 ( .A(n1070), .B(KEYINPUT16), .ZN(n1229) );
NOR3_X1 U887 ( .A1(n1102), .A2(n1186), .A3(n1187), .ZN(n1055) );
INV_X1 U888 ( .A(n1070), .ZN(n1186) );
INV_X1 U889 ( .A(n1230), .ZN(n1102) );
NAND4_X1 U890 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1059) );
AND4_X1 U891 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1234) );
NOR2_X1 U892 ( .A1(n1239), .A2(n1240), .ZN(n1233) );
NAND2_X1 U893 ( .A1(KEYINPUT25), .A2(n1197), .ZN(n1217) );
NOR2_X1 U894 ( .A1(n1073), .A2(G952), .ZN(n1165) );
XNOR2_X1 U895 ( .A(G146), .B(n1238), .ZN(G48) );
NAND2_X1 U896 ( .A1(n1241), .A2(n1242), .ZN(n1238) );
XNOR2_X1 U897 ( .A(G143), .B(n1237), .ZN(G45) );
NAND4_X1 U898 ( .A1(n1243), .A2(n1093), .A3(n1244), .A4(n1245), .ZN(n1237) );
XNOR2_X1 U899 ( .A(G140), .B(n1236), .ZN(G42) );
NAND4_X1 U900 ( .A1(n1246), .A2(n1083), .A3(n1087), .A4(n1242), .ZN(n1236) );
XNOR2_X1 U901 ( .A(G137), .B(n1235), .ZN(G39) );
NAND4_X1 U902 ( .A1(n1079), .A2(n1246), .A3(n1083), .A4(n1247), .ZN(n1235) );
XNOR2_X1 U903 ( .A(n1248), .B(n1240), .ZN(G36) );
AND3_X1 U904 ( .A1(n1243), .A2(n1230), .A3(n1083), .ZN(n1240) );
XOR2_X1 U905 ( .A(G131), .B(n1239), .Z(G33) );
AND3_X1 U906 ( .A1(n1243), .A2(n1242), .A3(n1083), .ZN(n1239) );
NOR2_X1 U907 ( .A1(n1249), .A2(n1092), .ZN(n1083) );
AND4_X1 U908 ( .A1(n1250), .A2(n1071), .A3(n1100), .A4(n1251), .ZN(n1243) );
XNOR2_X1 U909 ( .A(G128), .B(n1231), .ZN(G30) );
NAND2_X1 U910 ( .A1(n1241), .A2(n1230), .ZN(n1231) );
AND3_X1 U911 ( .A1(n1093), .A2(n1247), .A3(n1246), .ZN(n1241) );
AND4_X1 U912 ( .A1(n1071), .A2(n1100), .A3(n1088), .A4(n1251), .ZN(n1246) );
XNOR2_X1 U913 ( .A(n1252), .B(n1226), .ZN(G3) );
NOR3_X1 U914 ( .A1(n1085), .A2(n1187), .A3(n1066), .ZN(n1226) );
INV_X1 U915 ( .A(n1250), .ZN(n1085) );
XNOR2_X1 U916 ( .A(G125), .B(n1232), .ZN(G27) );
NAND4_X1 U917 ( .A1(n1088), .A2(n1251), .A3(n1253), .A4(n1254), .ZN(n1232) );
NOR3_X1 U918 ( .A1(n1101), .A2(n1247), .A3(n1100), .ZN(n1254) );
INV_X1 U919 ( .A(n1242), .ZN(n1101) );
NAND2_X1 U920 ( .A1(n1255), .A2(n1065), .ZN(n1251) );
NAND4_X1 U921 ( .A1(G953), .A2(G902), .A3(n1256), .A4(n1126), .ZN(n1255) );
INV_X1 U922 ( .A(G900), .ZN(n1126) );
XNOR2_X1 U923 ( .A(G122), .B(n1257), .ZN(G24) );
NAND2_X1 U924 ( .A1(KEYINPUT33), .A2(n1228), .ZN(n1257) );
AND4_X1 U925 ( .A1(n1258), .A2(n1070), .A3(n1244), .A4(n1245), .ZN(n1228) );
NOR2_X1 U926 ( .A1(n1088), .A2(n1247), .ZN(n1070) );
XOR2_X1 U927 ( .A(n1225), .B(n1259), .Z(G21) );
NOR2_X1 U928 ( .A1(KEYINPUT47), .A2(n1260), .ZN(n1259) );
AND4_X1 U929 ( .A1(n1258), .A2(n1079), .A3(n1247), .A4(n1088), .ZN(n1225) );
XNOR2_X1 U930 ( .A(n1261), .B(n1224), .ZN(G18) );
AND3_X1 U931 ( .A1(n1250), .A2(n1230), .A3(n1258), .ZN(n1224) );
NOR2_X1 U932 ( .A1(n1245), .A2(n1262), .ZN(n1230) );
INV_X1 U933 ( .A(n1244), .ZN(n1262) );
XOR2_X1 U934 ( .A(n1263), .B(n1223), .Z(G15) );
AND3_X1 U935 ( .A1(n1242), .A2(n1250), .A3(n1258), .ZN(n1223) );
AND3_X1 U936 ( .A1(n1253), .A2(n1264), .A3(n1069), .ZN(n1258) );
INV_X1 U937 ( .A(n1100), .ZN(n1069) );
NOR2_X1 U938 ( .A1(n1088), .A2(n1087), .ZN(n1250) );
INV_X1 U939 ( .A(n1247), .ZN(n1087) );
NOR2_X1 U940 ( .A1(n1244), .A2(n1104), .ZN(n1242) );
INV_X1 U941 ( .A(n1245), .ZN(n1104) );
XNOR2_X1 U942 ( .A(G113), .B(KEYINPUT4), .ZN(n1263) );
XNOR2_X1 U943 ( .A(G110), .B(n1265), .ZN(G12) );
NOR2_X1 U944 ( .A1(n1222), .A2(KEYINPUT48), .ZN(n1265) );
NOR4_X1 U945 ( .A1(n1066), .A2(n1187), .A3(n1247), .A4(n1266), .ZN(n1222) );
INV_X1 U946 ( .A(n1088), .ZN(n1266) );
XOR2_X1 U947 ( .A(n1267), .B(n1169), .Z(n1088) );
NAND2_X1 U948 ( .A1(G217), .A2(n1268), .ZN(n1169) );
NAND2_X1 U949 ( .A1(n1167), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U950 ( .A(n1270), .B(n1271), .ZN(n1167) );
AND3_X1 U951 ( .A1(G221), .A2(n1073), .A3(G234), .ZN(n1271) );
XNOR2_X1 U952 ( .A(n1272), .B(n1145), .ZN(n1270) );
INV_X1 U953 ( .A(G137), .ZN(n1145) );
NAND2_X1 U954 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U955 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XOR2_X1 U956 ( .A(KEYINPUT56), .B(n1277), .Z(n1276) );
XOR2_X1 U957 ( .A(n1278), .B(n1279), .Z(n1275) );
NAND2_X1 U958 ( .A1(n1280), .A2(n1281), .ZN(n1273) );
XNOR2_X1 U959 ( .A(n1278), .B(n1279), .ZN(n1281) );
XNOR2_X1 U960 ( .A(n1282), .B(G128), .ZN(n1279) );
NAND2_X1 U961 ( .A1(KEYINPUT30), .A2(n1260), .ZN(n1278) );
XOR2_X1 U962 ( .A(KEYINPUT27), .B(n1277), .Z(n1280) );
XNOR2_X1 U963 ( .A(n1283), .B(KEYINPUT57), .ZN(n1277) );
XNOR2_X1 U964 ( .A(n1284), .B(G472), .ZN(n1247) );
NAND2_X1 U965 ( .A1(n1285), .A2(n1269), .ZN(n1284) );
XNOR2_X1 U966 ( .A(n1286), .B(n1202), .ZN(n1285) );
XOR2_X1 U967 ( .A(n1287), .B(n1252), .Z(n1202) );
INV_X1 U968 ( .A(G101), .ZN(n1252) );
NAND2_X1 U969 ( .A1(n1288), .A2(G210), .ZN(n1287) );
NAND2_X1 U970 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
NAND2_X1 U971 ( .A1(n1291), .A2(n1201), .ZN(n1290) );
XOR2_X1 U972 ( .A(KEYINPUT29), .B(n1292), .Z(n1289) );
NOR2_X1 U973 ( .A1(n1291), .A2(n1201), .ZN(n1292) );
XOR2_X1 U974 ( .A(n1293), .B(n1294), .Z(n1201) );
INV_X1 U975 ( .A(n1295), .ZN(n1294) );
XNOR2_X1 U976 ( .A(n1296), .B(n1260), .ZN(n1293) );
NAND2_X1 U977 ( .A1(KEYINPUT11), .A2(n1261), .ZN(n1296) );
XNOR2_X1 U978 ( .A(n1297), .B(n1197), .ZN(n1291) );
NAND2_X1 U979 ( .A1(KEYINPUT60), .A2(n1198), .ZN(n1297) );
NAND3_X1 U980 ( .A1(n1100), .A2(n1264), .A3(n1253), .ZN(n1187) );
AND2_X1 U981 ( .A1(n1093), .A2(n1071), .ZN(n1253) );
XOR2_X1 U982 ( .A(n1097), .B(KEYINPUT53), .Z(n1071) );
AND2_X1 U983 ( .A1(G221), .A2(n1268), .ZN(n1097) );
NAND2_X1 U984 ( .A1(G234), .A2(n1269), .ZN(n1268) );
NOR2_X1 U985 ( .A1(n1068), .A2(n1092), .ZN(n1093) );
INV_X1 U986 ( .A(n1067), .ZN(n1092) );
NAND2_X1 U987 ( .A1(G214), .A2(n1298), .ZN(n1067) );
INV_X1 U988 ( .A(n1249), .ZN(n1068) );
XNOR2_X1 U989 ( .A(n1299), .B(n1300), .ZN(n1249) );
XNOR2_X1 U990 ( .A(KEYINPUT1), .B(n1113), .ZN(n1300) );
NAND2_X1 U991 ( .A1(G210), .A2(n1298), .ZN(n1113) );
NAND2_X1 U992 ( .A1(n1301), .A2(n1269), .ZN(n1298) );
INV_X1 U993 ( .A(G237), .ZN(n1301) );
NAND2_X1 U994 ( .A1(KEYINPUT8), .A2(n1112), .ZN(n1299) );
NAND2_X1 U995 ( .A1(n1302), .A2(n1269), .ZN(n1112) );
XNOR2_X1 U996 ( .A(n1197), .B(n1303), .ZN(n1302) );
XOR2_X1 U997 ( .A(n1215), .B(KEYINPUT5), .Z(n1303) );
XOR2_X1 U998 ( .A(n1304), .B(n1305), .Z(n1215) );
XOR2_X1 U999 ( .A(n1161), .B(n1306), .Z(n1305) );
NAND2_X1 U1000 ( .A1(G224), .A2(n1073), .ZN(n1306) );
NAND2_X1 U1001 ( .A1(n1307), .A2(n1308), .ZN(n1161) );
NAND2_X1 U1002 ( .A1(G122), .A2(n1282), .ZN(n1308) );
XOR2_X1 U1003 ( .A(KEYINPUT51), .B(n1309), .Z(n1307) );
NOR2_X1 U1004 ( .A1(G122), .A2(n1282), .ZN(n1309) );
INV_X1 U1005 ( .A(G110), .ZN(n1282) );
XNOR2_X1 U1006 ( .A(n1310), .B(n1129), .ZN(n1304) );
INV_X1 U1007 ( .A(G125), .ZN(n1129) );
NAND3_X1 U1008 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1310) );
NAND2_X1 U1009 ( .A1(KEYINPUT63), .A2(n1164), .ZN(n1313) );
NAND3_X1 U1010 ( .A1(n1314), .A2(n1315), .A3(n1159), .ZN(n1312) );
INV_X1 U1011 ( .A(KEYINPUT63), .ZN(n1315) );
OR2_X1 U1012 ( .A1(n1159), .A2(n1314), .ZN(n1311) );
NOR2_X1 U1013 ( .A1(KEYINPUT6), .A2(n1164), .ZN(n1314) );
XOR2_X1 U1014 ( .A(n1213), .B(KEYINPUT9), .Z(n1164) );
XOR2_X1 U1015 ( .A(n1295), .B(n1316), .Z(n1159) );
NOR2_X1 U1016 ( .A1(KEYINPUT12), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1017 ( .A(n1261), .B(n1318), .ZN(n1317) );
NOR2_X1 U1018 ( .A1(KEYINPUT23), .A2(n1319), .ZN(n1318) );
XNOR2_X1 U1019 ( .A(KEYINPUT18), .B(n1260), .ZN(n1319) );
INV_X1 U1020 ( .A(G119), .ZN(n1260) );
INV_X1 U1021 ( .A(G116), .ZN(n1261) );
INV_X1 U1022 ( .A(n1200), .ZN(n1197) );
NAND2_X1 U1023 ( .A1(n1320), .A2(n1321), .ZN(n1200) );
NAND2_X1 U1024 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
INV_X1 U1025 ( .A(n1324), .ZN(n1323) );
NAND2_X1 U1026 ( .A1(n1325), .A2(n1326), .ZN(n1322) );
NAND2_X1 U1027 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1028 ( .A1(n1329), .A2(G146), .ZN(n1325) );
NAND2_X1 U1029 ( .A1(n1324), .A2(n1330), .ZN(n1320) );
NAND2_X1 U1030 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND2_X1 U1031 ( .A1(G146), .A2(n1327), .ZN(n1332) );
NAND2_X1 U1032 ( .A1(n1329), .A2(n1328), .ZN(n1331) );
XNOR2_X1 U1033 ( .A(n1333), .B(G128), .ZN(n1329) );
XNOR2_X1 U1034 ( .A(KEYINPUT61), .B(KEYINPUT52), .ZN(n1333) );
NOR2_X1 U1035 ( .A1(KEYINPUT40), .A2(n1334), .ZN(n1324) );
NAND2_X1 U1036 ( .A1(n1065), .A2(n1335), .ZN(n1264) );
NAND4_X1 U1037 ( .A1(n1336), .A2(G953), .A3(G902), .A4(n1156), .ZN(n1335) );
INV_X1 U1038 ( .A(G898), .ZN(n1156) );
XOR2_X1 U1039 ( .A(n1256), .B(KEYINPUT54), .Z(n1336) );
NAND3_X1 U1040 ( .A1(n1256), .A2(n1073), .A3(G952), .ZN(n1065) );
NAND2_X1 U1041 ( .A1(G237), .A2(G234), .ZN(n1256) );
XNOR2_X1 U1042 ( .A(n1337), .B(G469), .ZN(n1100) );
NAND2_X1 U1043 ( .A1(n1338), .A2(n1269), .ZN(n1337) );
INV_X1 U1044 ( .A(G902), .ZN(n1269) );
XOR2_X1 U1045 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1046 ( .A(n1341), .B(n1342), .Z(n1340) );
NAND2_X1 U1047 ( .A1(KEYINPUT42), .A2(G140), .ZN(n1342) );
NAND2_X1 U1048 ( .A1(n1343), .A2(n1344), .ZN(n1341) );
NAND2_X1 U1049 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1050 ( .A1(KEYINPUT2), .A2(n1347), .ZN(n1346) );
NAND2_X1 U1051 ( .A1(n1199), .A2(n1348), .ZN(n1347) );
INV_X1 U1052 ( .A(n1198), .ZN(n1199) );
NAND2_X1 U1053 ( .A1(n1198), .A2(n1349), .ZN(n1343) );
NAND2_X1 U1054 ( .A1(n1348), .A2(n1350), .ZN(n1349) );
NAND2_X1 U1055 ( .A1(n1351), .A2(KEYINPUT2), .ZN(n1350) );
INV_X1 U1056 ( .A(n1345), .ZN(n1351) );
XNOR2_X1 U1057 ( .A(n1213), .B(n1352), .ZN(n1345) );
NOR2_X1 U1058 ( .A1(KEYINPUT22), .A2(n1138), .ZN(n1352) );
INV_X1 U1059 ( .A(n1141), .ZN(n1138) );
XOR2_X1 U1060 ( .A(n1353), .B(n1327), .Z(n1141) );
NAND3_X1 U1061 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1353) );
OR2_X1 U1062 ( .A1(G146), .A2(KEYINPUT7), .ZN(n1356) );
NAND3_X1 U1063 ( .A1(KEYINPUT7), .A2(n1357), .A3(n1358), .ZN(n1355) );
OR2_X1 U1064 ( .A1(n1358), .A2(n1357), .ZN(n1354) );
AND2_X1 U1065 ( .A1(KEYINPUT10), .A2(G146), .ZN(n1357) );
XOR2_X1 U1066 ( .A(G143), .B(KEYINPUT3), .Z(n1358) );
XNOR2_X1 U1067 ( .A(G101), .B(n1359), .ZN(n1213) );
XOR2_X1 U1068 ( .A(G107), .B(G104), .Z(n1359) );
INV_X1 U1069 ( .A(KEYINPUT21), .ZN(n1348) );
XOR2_X1 U1070 ( .A(G137), .B(n1146), .Z(n1198) );
XOR2_X1 U1071 ( .A(G131), .B(G134), .Z(n1146) );
XNOR2_X1 U1072 ( .A(G110), .B(n1360), .ZN(n1339) );
NOR2_X1 U1073 ( .A1(KEYINPUT14), .A2(n1361), .ZN(n1360) );
XOR2_X1 U1074 ( .A(KEYINPUT35), .B(n1210), .Z(n1361) );
NOR2_X1 U1075 ( .A1(n1120), .A2(G953), .ZN(n1210) );
INV_X1 U1076 ( .A(G227), .ZN(n1120) );
INV_X1 U1077 ( .A(n1079), .ZN(n1066) );
NOR2_X1 U1078 ( .A1(n1244), .A2(n1245), .ZN(n1079) );
XNOR2_X1 U1079 ( .A(n1362), .B(G475), .ZN(n1245) );
OR2_X1 U1080 ( .A1(n1183), .A2(G902), .ZN(n1362) );
XNOR2_X1 U1081 ( .A(n1363), .B(n1364), .ZN(n1183) );
XOR2_X1 U1082 ( .A(n1283), .B(n1365), .Z(n1364) );
XOR2_X1 U1083 ( .A(n1366), .B(n1367), .Z(n1365) );
NOR2_X1 U1084 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
XOR2_X1 U1085 ( .A(n1370), .B(KEYINPUT39), .Z(n1369) );
NAND2_X1 U1086 ( .A1(n1371), .A2(G104), .ZN(n1370) );
NOR2_X1 U1087 ( .A1(G104), .A2(n1371), .ZN(n1368) );
XNOR2_X1 U1088 ( .A(G122), .B(n1295), .ZN(n1371) );
XOR2_X1 U1089 ( .A(G113), .B(KEYINPUT45), .Z(n1295) );
NAND2_X1 U1090 ( .A1(n1288), .A2(G214), .ZN(n1366) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1288) );
XNOR2_X1 U1092 ( .A(G125), .B(n1372), .ZN(n1283) );
XNOR2_X1 U1093 ( .A(n1328), .B(G140), .ZN(n1372) );
INV_X1 U1094 ( .A(G146), .ZN(n1328) );
XNOR2_X1 U1095 ( .A(G131), .B(n1373), .ZN(n1363) );
XNOR2_X1 U1096 ( .A(KEYINPUT58), .B(n1334), .ZN(n1373) );
INV_X1 U1097 ( .A(G143), .ZN(n1334) );
XOR2_X1 U1098 ( .A(n1374), .B(n1177), .Z(n1244) );
INV_X1 U1099 ( .A(G478), .ZN(n1177) );
NAND2_X1 U1100 ( .A1(KEYINPUT50), .A2(n1111), .ZN(n1374) );
NOR2_X1 U1101 ( .A1(n1176), .A2(G902), .ZN(n1111) );
XOR2_X1 U1102 ( .A(n1375), .B(n1376), .Z(n1176) );
XOR2_X1 U1103 ( .A(n1377), .B(n1378), .Z(n1376) );
XOR2_X1 U1104 ( .A(n1379), .B(n1380), .Z(n1378) );
AND3_X1 U1105 ( .A1(G217), .A2(n1073), .A3(G234), .ZN(n1380) );
INV_X1 U1106 ( .A(G953), .ZN(n1073) );
NAND2_X1 U1107 ( .A1(KEYINPUT55), .A2(n1248), .ZN(n1379) );
INV_X1 U1108 ( .A(G134), .ZN(n1248) );
XNOR2_X1 U1109 ( .A(G107), .B(G116), .ZN(n1377) );
XOR2_X1 U1110 ( .A(n1381), .B(n1382), .Z(n1375) );
XNOR2_X1 U1111 ( .A(n1327), .B(G122), .ZN(n1382) );
INV_X1 U1112 ( .A(G128), .ZN(n1327) );
XNOR2_X1 U1113 ( .A(G143), .B(KEYINPUT0), .ZN(n1381) );
endmodule


