//Key = 0110110000101100011100000010101001100011110110111101011111001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306;

NAND2_X1 U726 ( .A1(n996), .A2(n997), .ZN(G9) );
NAND3_X1 U727 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
XOR2_X1 U728 ( .A(n1001), .B(KEYINPUT16), .Z(n996) );
NAND2_X1 U729 ( .A1(G107), .A2(n1002), .ZN(n1001) );
NAND2_X1 U730 ( .A1(n1000), .A2(n998), .ZN(n1002) );
XNOR2_X1 U731 ( .A(n1003), .B(KEYINPUT22), .ZN(n998) );
NOR2_X1 U732 ( .A1(n1004), .A2(n1005), .ZN(G75) );
XOR2_X1 U733 ( .A(KEYINPUT37), .B(n1006), .Z(n1005) );
NOR4_X1 U734 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
NOR3_X1 U735 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1010) );
NOR2_X1 U736 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
XOR2_X1 U737 ( .A(n1016), .B(KEYINPUT60), .Z(n1015) );
NOR2_X1 U738 ( .A1(n1017), .A2(n1018), .ZN(n1012) );
NOR3_X1 U739 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NOR2_X1 U740 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U741 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U742 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1022) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR3_X1 U746 ( .A1(n1034), .A2(n1035), .A3(n1019), .ZN(n1009) );
NAND3_X1 U747 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1034) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1016), .ZN(n1008) );
OR4_X1 U749 ( .A1(n1019), .A2(n1025), .A3(n1021), .A4(n1029), .ZN(n1016) );
INV_X1 U750 ( .A(n1036), .ZN(n1029) );
INV_X1 U751 ( .A(n1040), .ZN(n1021) );
NAND3_X1 U752 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1007) );
INV_X1 U753 ( .A(n1044), .ZN(n1042) );
NOR2_X1 U754 ( .A1(G952), .A2(n1044), .ZN(n1004) );
NAND2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND4_X1 U756 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
NOR3_X1 U757 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
XNOR2_X1 U758 ( .A(n1054), .B(n1055), .ZN(n1052) );
NAND2_X1 U759 ( .A1(KEYINPUT5), .A2(n1056), .ZN(n1054) );
NAND3_X1 U760 ( .A1(n1033), .A2(n1057), .A3(n1014), .ZN(n1051) );
NOR3_X1 U761 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1049) );
AND3_X1 U762 ( .A1(KEYINPUT43), .A2(n1061), .A3(G478), .ZN(n1060) );
NOR2_X1 U763 ( .A1(KEYINPUT43), .A2(G478), .ZN(n1059) );
XNOR2_X1 U764 ( .A(G475), .B(n1062), .ZN(n1058) );
XOR2_X1 U765 ( .A(n1063), .B(n1064), .Z(n1048) );
XNOR2_X1 U766 ( .A(KEYINPUT27), .B(n1065), .ZN(n1064) );
XNOR2_X1 U767 ( .A(n1032), .B(KEYINPUT52), .ZN(n1047) );
XOR2_X1 U768 ( .A(n1066), .B(n1067), .Z(G72) );
XOR2_X1 U769 ( .A(n1068), .B(n1069), .Z(n1067) );
NAND2_X1 U770 ( .A1(G953), .A2(n1070), .ZN(n1069) );
NAND2_X1 U771 ( .A1(G900), .A2(G227), .ZN(n1070) );
NAND2_X1 U772 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
NAND2_X1 U773 ( .A1(G953), .A2(n1073), .ZN(n1072) );
XOR2_X1 U774 ( .A(n1074), .B(n1075), .Z(n1071) );
XOR2_X1 U775 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U776 ( .A(n1078), .B(KEYINPUT26), .Z(n1077) );
XOR2_X1 U777 ( .A(n1079), .B(n1080), .Z(n1074) );
NOR2_X1 U778 ( .A1(n1041), .A2(G953), .ZN(n1066) );
XOR2_X1 U779 ( .A(n1081), .B(n1082), .Z(G69) );
NOR2_X1 U780 ( .A1(n1083), .A2(n1045), .ZN(n1082) );
AND2_X1 U781 ( .A1(G224), .A2(G898), .ZN(n1083) );
NOR2_X1 U782 ( .A1(KEYINPUT11), .A2(n1084), .ZN(n1081) );
XOR2_X1 U783 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U784 ( .A1(n1043), .A2(G953), .ZN(n1086) );
NAND3_X1 U785 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
NAND2_X1 U786 ( .A1(G953), .A2(n1090), .ZN(n1087) );
NOR2_X1 U787 ( .A1(n1091), .A2(n1092), .ZN(G66) );
XNOR2_X1 U788 ( .A(n1093), .B(n1094), .ZN(n1092) );
NOR2_X1 U789 ( .A1(n1056), .A2(n1095), .ZN(n1094) );
NOR2_X1 U790 ( .A1(n1091), .A2(n1096), .ZN(G63) );
XNOR2_X1 U791 ( .A(n1097), .B(n1098), .ZN(n1096) );
AND2_X1 U792 ( .A1(G478), .A2(n1099), .ZN(n1098) );
NOR2_X1 U793 ( .A1(n1091), .A2(n1100), .ZN(G60) );
XNOR2_X1 U794 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR2_X1 U795 ( .A1(n1103), .A2(n1095), .ZN(n1102) );
XNOR2_X1 U796 ( .A(G104), .B(n1104), .ZN(G6) );
NOR2_X1 U797 ( .A1(n1105), .A2(KEYINPUT14), .ZN(n1104) );
NOR2_X1 U798 ( .A1(n1091), .A2(n1106), .ZN(G57) );
NOR2_X1 U799 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XOR2_X1 U800 ( .A(KEYINPUT24), .B(n1109), .Z(n1108) );
NOR2_X1 U801 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U802 ( .A(n1112), .B(KEYINPUT46), .Z(n1111) );
INV_X1 U803 ( .A(n1113), .ZN(n1110) );
NOR2_X1 U804 ( .A1(n1113), .A2(n1114), .ZN(n1107) );
XNOR2_X1 U805 ( .A(KEYINPUT46), .B(n1112), .ZN(n1114) );
XNOR2_X1 U806 ( .A(n1115), .B(n1116), .ZN(n1113) );
XOR2_X1 U807 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U808 ( .A(n1119), .B(n1120), .Z(n1115) );
NAND3_X1 U809 ( .A1(n1099), .A2(G472), .A3(KEYINPUT44), .ZN(n1119) );
NOR2_X1 U810 ( .A1(n1091), .A2(n1121), .ZN(G54) );
XOR2_X1 U811 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U813 ( .A(n1126), .B(n1127), .Z(n1122) );
AND2_X1 U814 ( .A1(G469), .A2(n1099), .ZN(n1127) );
INV_X1 U815 ( .A(n1095), .ZN(n1099) );
XOR2_X1 U816 ( .A(n1128), .B(n1129), .Z(n1126) );
NOR2_X1 U817 ( .A1(KEYINPUT50), .A2(n1120), .ZN(n1129) );
NAND2_X1 U818 ( .A1(KEYINPUT61), .A2(n1130), .ZN(n1128) );
XOR2_X1 U819 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U820 ( .A(G110), .B(n1133), .ZN(n1132) );
NAND2_X1 U821 ( .A1(KEYINPUT49), .A2(G140), .ZN(n1131) );
NOR2_X1 U822 ( .A1(n1091), .A2(n1134), .ZN(G51) );
XOR2_X1 U823 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U824 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U825 ( .A1(n1065), .A2(n1095), .ZN(n1137) );
NAND2_X1 U826 ( .A1(G902), .A2(n1139), .ZN(n1095) );
NAND2_X1 U827 ( .A1(n1043), .A2(n1140), .ZN(n1139) );
XOR2_X1 U828 ( .A(KEYINPUT29), .B(n1041), .Z(n1140) );
AND4_X1 U829 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1041) );
NOR4_X1 U830 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1144) );
NOR2_X1 U831 ( .A1(n1149), .A2(n1150), .ZN(n1143) );
NAND3_X1 U832 ( .A1(n1151), .A2(n1038), .A3(n1152), .ZN(n1141) );
XNOR2_X1 U833 ( .A(n1153), .B(KEYINPUT10), .ZN(n1152) );
AND4_X1 U834 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1043) );
NOR4_X1 U835 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1105), .ZN(n1157) );
AND3_X1 U836 ( .A1(n1031), .A2(n1161), .A3(n1162), .ZN(n1105) );
NAND2_X1 U837 ( .A1(n1000), .A2(n1031), .ZN(n1156) );
AND2_X1 U838 ( .A1(n1161), .A2(n1163), .ZN(n1000) );
NAND4_X1 U839 ( .A1(n1027), .A2(n1038), .A3(n1164), .A4(n1037), .ZN(n1154) );
OR2_X1 U840 ( .A1(n1162), .A2(n1163), .ZN(n1037) );
XOR2_X1 U841 ( .A(KEYINPUT58), .B(KEYINPUT15), .Z(n1135) );
NOR2_X1 U842 ( .A1(n1165), .A2(G952), .ZN(n1091) );
XNOR2_X1 U843 ( .A(n1045), .B(KEYINPUT1), .ZN(n1165) );
XNOR2_X1 U844 ( .A(n1150), .B(n1166), .ZN(G48) );
NAND2_X1 U845 ( .A1(KEYINPUT54), .A2(G146), .ZN(n1166) );
AND3_X1 U846 ( .A1(n1162), .A2(n1153), .A3(n1167), .ZN(n1150) );
XOR2_X1 U847 ( .A(n1168), .B(G143), .Z(G45) );
NAND2_X1 U848 ( .A1(KEYINPUT55), .A2(n1142), .ZN(n1168) );
NAND4_X1 U849 ( .A1(n1169), .A2(n1031), .A3(n1170), .A4(n1153), .ZN(n1142) );
AND2_X1 U850 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U851 ( .A(n1149), .B(n1173), .Z(G42) );
NOR2_X1 U852 ( .A1(KEYINPUT32), .A2(n1174), .ZN(n1173) );
XNOR2_X1 U853 ( .A(KEYINPUT38), .B(n1175), .ZN(n1174) );
AND2_X1 U854 ( .A1(n1151), .A2(n1176), .ZN(n1149) );
XOR2_X1 U855 ( .A(G137), .B(n1148), .Z(G39) );
AND3_X1 U856 ( .A1(n1167), .A2(n1040), .A3(n1177), .ZN(n1148) );
XOR2_X1 U857 ( .A(G134), .B(n1147), .Z(G36) );
AND3_X1 U858 ( .A1(n1169), .A2(n1163), .A3(n1176), .ZN(n1147) );
XOR2_X1 U859 ( .A(G131), .B(n1146), .Z(G33) );
AND3_X1 U860 ( .A1(n1169), .A2(n1162), .A3(n1176), .ZN(n1146) );
NOR2_X1 U861 ( .A1(n1035), .A2(n1003), .ZN(n1176) );
INV_X1 U862 ( .A(n1177), .ZN(n1035) );
NOR2_X1 U863 ( .A1(n1011), .A2(n1017), .ZN(n1177) );
INV_X1 U864 ( .A(n1014), .ZN(n1017) );
AND2_X1 U865 ( .A1(n1027), .A2(n1178), .ZN(n1169) );
XOR2_X1 U866 ( .A(n1179), .B(n1145), .Z(G30) );
AND3_X1 U867 ( .A1(n1163), .A2(n1153), .A3(n1167), .ZN(n1145) );
AND4_X1 U868 ( .A1(n1031), .A2(n1053), .A3(n1180), .A4(n1178), .ZN(n1167) );
XNOR2_X1 U869 ( .A(G128), .B(KEYINPUT18), .ZN(n1179) );
XNOR2_X1 U870 ( .A(n1181), .B(n1160), .ZN(G3) );
AND2_X1 U871 ( .A1(n1027), .A2(n1182), .ZN(n1160) );
XOR2_X1 U872 ( .A(n1183), .B(n1184), .Z(G27) );
NAND3_X1 U873 ( .A1(n1038), .A2(n1153), .A3(n1151), .ZN(n1184) );
AND3_X1 U874 ( .A1(n1026), .A2(n1178), .A3(n1162), .ZN(n1151) );
NAND2_X1 U875 ( .A1(n1019), .A2(n1185), .ZN(n1178) );
NAND4_X1 U876 ( .A1(G953), .A2(G902), .A3(n1186), .A4(n1073), .ZN(n1185) );
INV_X1 U877 ( .A(G900), .ZN(n1073) );
NAND2_X1 U878 ( .A1(n1187), .A2(KEYINPUT57), .ZN(n1183) );
XNOR2_X1 U879 ( .A(G125), .B(KEYINPUT47), .ZN(n1187) );
XNOR2_X1 U880 ( .A(G122), .B(n1188), .ZN(G24) );
NOR2_X1 U881 ( .A1(n1159), .A2(KEYINPUT8), .ZN(n1188) );
AND4_X1 U882 ( .A1(n1038), .A2(n1161), .A3(n1172), .A4(n1171), .ZN(n1159) );
XNOR2_X1 U883 ( .A(n1189), .B(KEYINPUT48), .ZN(n1172) );
AND2_X1 U884 ( .A1(n1164), .A2(n1036), .ZN(n1161) );
NOR2_X1 U885 ( .A1(n1180), .A2(n1053), .ZN(n1036) );
NAND2_X1 U886 ( .A1(n1190), .A2(n1191), .ZN(G21) );
NAND2_X1 U887 ( .A1(G119), .A2(n1155), .ZN(n1191) );
XOR2_X1 U888 ( .A(n1192), .B(KEYINPUT0), .Z(n1190) );
OR2_X1 U889 ( .A1(n1155), .A2(G119), .ZN(n1192) );
NAND4_X1 U890 ( .A1(n1038), .A2(n1040), .A3(n1193), .A4(n1164), .ZN(n1155) );
NOR2_X1 U891 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U892 ( .A(G116), .B(n1196), .ZN(G18) );
NAND4_X1 U893 ( .A1(n1027), .A2(n1163), .A3(n1164), .A4(n1197), .ZN(n1196) );
XNOR2_X1 U894 ( .A(KEYINPUT42), .B(n1025), .ZN(n1197) );
AND2_X1 U895 ( .A1(n1198), .A2(n1171), .ZN(n1163) );
XNOR2_X1 U896 ( .A(G113), .B(n1199), .ZN(G15) );
NAND4_X1 U897 ( .A1(n1200), .A2(n1162), .A3(n1038), .A4(n1164), .ZN(n1199) );
INV_X1 U898 ( .A(n1025), .ZN(n1038) );
NAND2_X1 U899 ( .A1(n1201), .A2(n1033), .ZN(n1025) );
INV_X1 U900 ( .A(n1032), .ZN(n1201) );
NOR2_X1 U901 ( .A1(n1198), .A2(n1171), .ZN(n1162) );
INV_X1 U902 ( .A(n1189), .ZN(n1198) );
XNOR2_X1 U903 ( .A(n1027), .B(KEYINPUT40), .ZN(n1200) );
NOR2_X1 U904 ( .A1(n1180), .A2(n1195), .ZN(n1027) );
INV_X1 U905 ( .A(n1053), .ZN(n1195) );
INV_X1 U906 ( .A(n1194), .ZN(n1180) );
XNOR2_X1 U907 ( .A(G110), .B(n1202), .ZN(G12) );
NAND2_X1 U908 ( .A1(KEYINPUT12), .A2(n1158), .ZN(n1202) );
AND2_X1 U909 ( .A1(n1182), .A2(n1026), .ZN(n1158) );
NOR2_X1 U910 ( .A1(n1053), .A2(n1194), .ZN(n1026) );
XNOR2_X1 U911 ( .A(n1055), .B(n1056), .ZN(n1194) );
NAND2_X1 U912 ( .A1(G217), .A2(n1203), .ZN(n1056) );
NAND2_X1 U913 ( .A1(n1093), .A2(n1204), .ZN(n1055) );
XNOR2_X1 U914 ( .A(n1205), .B(n1206), .ZN(n1093) );
XNOR2_X1 U915 ( .A(n1207), .B(n1208), .ZN(n1206) );
XNOR2_X1 U916 ( .A(n1209), .B(n1210), .ZN(n1208) );
NOR2_X1 U917 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
INV_X1 U918 ( .A(G221), .ZN(n1212) );
XOR2_X1 U919 ( .A(n1213), .B(n1214), .Z(n1205) );
XOR2_X1 U920 ( .A(G137), .B(G110), .Z(n1214) );
NAND2_X1 U921 ( .A1(n1215), .A2(KEYINPUT56), .ZN(n1213) );
XNOR2_X1 U922 ( .A(n1216), .B(n1217), .ZN(n1215) );
XNOR2_X1 U923 ( .A(G119), .B(KEYINPUT28), .ZN(n1216) );
XNOR2_X1 U924 ( .A(n1218), .B(G472), .ZN(n1053) );
NAND2_X1 U925 ( .A1(n1219), .A2(n1204), .ZN(n1218) );
XOR2_X1 U926 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U927 ( .A(n1112), .B(n1118), .Z(n1221) );
XOR2_X1 U928 ( .A(n1222), .B(n1223), .Z(n1118) );
XNOR2_X1 U929 ( .A(KEYINPUT4), .B(n1224), .ZN(n1223) );
INV_X1 U930 ( .A(G113), .ZN(n1224) );
NAND2_X1 U931 ( .A1(KEYINPUT41), .A2(n1225), .ZN(n1222) );
XNOR2_X1 U932 ( .A(n1226), .B(G116), .ZN(n1225) );
XNOR2_X1 U933 ( .A(n1227), .B(n1181), .ZN(n1112) );
INV_X1 U934 ( .A(G101), .ZN(n1181) );
NAND2_X1 U935 ( .A1(n1228), .A2(G210), .ZN(n1227) );
XOR2_X1 U936 ( .A(n1229), .B(n1117), .Z(n1220) );
XOR2_X1 U937 ( .A(n1230), .B(KEYINPUT33), .Z(n1117) );
NAND2_X1 U938 ( .A1(KEYINPUT62), .A2(n1120), .ZN(n1229) );
AND3_X1 U939 ( .A1(n1031), .A2(n1164), .A3(n1040), .ZN(n1182) );
NOR2_X1 U940 ( .A1(n1171), .A2(n1189), .ZN(n1040) );
XNOR2_X1 U941 ( .A(n1231), .B(n1062), .ZN(n1189) );
NAND2_X1 U942 ( .A1(n1101), .A2(n1204), .ZN(n1062) );
XNOR2_X1 U943 ( .A(n1232), .B(n1233), .ZN(n1101) );
XOR2_X1 U944 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND2_X1 U945 ( .A1(n1228), .A2(G214), .ZN(n1235) );
NOR2_X1 U946 ( .A1(G953), .A2(G237), .ZN(n1228) );
NAND2_X1 U947 ( .A1(n1236), .A2(n1237), .ZN(n1234) );
NAND2_X1 U948 ( .A1(n1238), .A2(G104), .ZN(n1237) );
XOR2_X1 U949 ( .A(KEYINPUT51), .B(n1239), .Z(n1236) );
NOR2_X1 U950 ( .A1(G104), .A2(n1238), .ZN(n1239) );
XNOR2_X1 U951 ( .A(G122), .B(n1240), .ZN(n1238) );
NOR2_X1 U952 ( .A1(G113), .A2(KEYINPUT9), .ZN(n1240) );
XOR2_X1 U953 ( .A(n1079), .B(n1207), .Z(n1232) );
XOR2_X1 U954 ( .A(n1080), .B(KEYINPUT25), .Z(n1207) );
XNOR2_X1 U955 ( .A(G125), .B(n1175), .ZN(n1080) );
XOR2_X1 U956 ( .A(n1241), .B(G131), .Z(n1079) );
NAND2_X1 U957 ( .A1(KEYINPUT2), .A2(n1103), .ZN(n1231) );
INV_X1 U958 ( .A(G475), .ZN(n1103) );
NAND2_X1 U959 ( .A1(n1057), .A2(n1242), .ZN(n1171) );
NAND2_X1 U960 ( .A1(G478), .A2(n1061), .ZN(n1242) );
OR2_X1 U961 ( .A1(n1061), .A2(G478), .ZN(n1057) );
NAND2_X1 U962 ( .A1(n1097), .A2(n1204), .ZN(n1061) );
XNOR2_X1 U963 ( .A(n1243), .B(n1244), .ZN(n1097) );
XNOR2_X1 U964 ( .A(n1245), .B(n1246), .ZN(n1244) );
NAND3_X1 U965 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1245) );
NAND2_X1 U966 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND2_X1 U967 ( .A1(n1252), .A2(KEYINPUT17), .ZN(n1251) );
XNOR2_X1 U968 ( .A(G107), .B(KEYINPUT63), .ZN(n1252) );
NAND3_X1 U969 ( .A1(KEYINPUT17), .A2(n1253), .A3(n999), .ZN(n1248) );
INV_X1 U970 ( .A(n1250), .ZN(n1253) );
XOR2_X1 U971 ( .A(G116), .B(n1254), .Z(n1250) );
NOR2_X1 U972 ( .A1(KEYINPUT36), .A2(n1255), .ZN(n1254) );
INV_X1 U973 ( .A(G122), .ZN(n1255) );
OR2_X1 U974 ( .A1(n999), .A2(KEYINPUT17), .ZN(n1247) );
INV_X1 U975 ( .A(G107), .ZN(n999) );
XOR2_X1 U976 ( .A(n1256), .B(n1257), .Z(n1243) );
NOR2_X1 U977 ( .A1(n1211), .A2(n1258), .ZN(n1257) );
INV_X1 U978 ( .A(G217), .ZN(n1258) );
NAND2_X1 U979 ( .A1(n1259), .A2(n1045), .ZN(n1211) );
XNOR2_X1 U980 ( .A(G234), .B(KEYINPUT34), .ZN(n1259) );
XNOR2_X1 U981 ( .A(G134), .B(G143), .ZN(n1256) );
AND2_X1 U982 ( .A1(n1153), .A2(n1260), .ZN(n1164) );
NAND2_X1 U983 ( .A1(n1019), .A2(n1261), .ZN(n1260) );
NAND4_X1 U984 ( .A1(G953), .A2(G902), .A3(n1186), .A4(n1090), .ZN(n1261) );
INV_X1 U985 ( .A(G898), .ZN(n1090) );
NAND3_X1 U986 ( .A1(n1186), .A2(n1045), .A3(G952), .ZN(n1019) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1186) );
INV_X1 U988 ( .A(n1039), .ZN(n1153) );
NAND2_X1 U989 ( .A1(n1011), .A2(n1014), .ZN(n1039) );
NAND2_X1 U990 ( .A1(G214), .A2(n1262), .ZN(n1014) );
XNOR2_X1 U991 ( .A(n1263), .B(n1065), .ZN(n1011) );
NAND2_X1 U992 ( .A1(G210), .A2(n1262), .ZN(n1065) );
NAND2_X1 U993 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
INV_X1 U994 ( .A(G237), .ZN(n1264) );
NAND2_X1 U995 ( .A1(KEYINPUT13), .A2(n1063), .ZN(n1263) );
NAND2_X1 U996 ( .A1(n1266), .A2(n1204), .ZN(n1063) );
XNOR2_X1 U997 ( .A(n1138), .B(KEYINPUT6), .ZN(n1266) );
XNOR2_X1 U998 ( .A(n1267), .B(n1268), .ZN(n1138) );
XOR2_X1 U999 ( .A(n1269), .B(n1270), .Z(n1268) );
NAND3_X1 U1000 ( .A1(n1271), .A2(n1272), .A3(n1088), .ZN(n1270) );
NAND2_X1 U1001 ( .A1(n1273), .A2(n1274), .ZN(n1088) );
NAND2_X1 U1002 ( .A1(KEYINPUT45), .A2(n1275), .ZN(n1272) );
NAND3_X1 U1003 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1275) );
INV_X1 U1004 ( .A(n1273), .ZN(n1278) );
NOR2_X1 U1005 ( .A1(n1279), .A2(n1280), .ZN(n1273) );
NAND3_X1 U1006 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1277) );
NAND2_X1 U1007 ( .A1(n1274), .A2(n1282), .ZN(n1276) );
OR2_X1 U1008 ( .A1(n1089), .A2(KEYINPUT45), .ZN(n1271) );
AND2_X1 U1009 ( .A1(n1283), .A2(n1284), .ZN(n1089) );
NAND2_X1 U1010 ( .A1(n1285), .A2(n1280), .ZN(n1284) );
INV_X1 U1011 ( .A(n1282), .ZN(n1280) );
XNOR2_X1 U1012 ( .A(n1279), .B(n1274), .ZN(n1285) );
INV_X1 U1013 ( .A(n1281), .ZN(n1274) );
NAND3_X1 U1014 ( .A1(n1281), .A2(n1279), .A3(n1282), .ZN(n1283) );
XOR2_X1 U1015 ( .A(G122), .B(G110), .Z(n1282) );
XOR2_X1 U1016 ( .A(n1286), .B(n1287), .Z(n1279) );
NOR2_X1 U1017 ( .A1(KEYINPUT31), .A2(n1226), .ZN(n1287) );
INV_X1 U1018 ( .A(G119), .ZN(n1226) );
XNOR2_X1 U1019 ( .A(G113), .B(G116), .ZN(n1286) );
XOR2_X1 U1020 ( .A(n1288), .B(n1289), .Z(n1281) );
XNOR2_X1 U1021 ( .A(G101), .B(KEYINPUT39), .ZN(n1288) );
NAND2_X1 U1022 ( .A1(G224), .A2(n1045), .ZN(n1269) );
XOR2_X1 U1023 ( .A(n1230), .B(G125), .Z(n1267) );
NAND2_X1 U1024 ( .A1(n1290), .A2(n1291), .ZN(n1230) );
OR2_X1 U1025 ( .A1(n1292), .A2(n1217), .ZN(n1291) );
XOR2_X1 U1026 ( .A(n1293), .B(KEYINPUT3), .Z(n1290) );
NAND2_X1 U1027 ( .A1(n1217), .A2(n1292), .ZN(n1293) );
XOR2_X1 U1028 ( .A(G143), .B(n1294), .Z(n1292) );
NOR2_X1 U1029 ( .A1(KEYINPUT21), .A2(n1209), .ZN(n1294) );
INV_X1 U1030 ( .A(n1003), .ZN(n1031) );
NAND2_X1 U1031 ( .A1(n1032), .A2(n1033), .ZN(n1003) );
NAND2_X1 U1032 ( .A1(G221), .A2(n1203), .ZN(n1033) );
NAND2_X1 U1033 ( .A1(G234), .A2(n1265), .ZN(n1203) );
XNOR2_X1 U1034 ( .A(n1295), .B(G469), .ZN(n1032) );
NAND2_X1 U1035 ( .A1(n1296), .A2(n1204), .ZN(n1295) );
XNOR2_X1 U1036 ( .A(n1265), .B(KEYINPUT53), .ZN(n1204) );
INV_X1 U1037 ( .A(G902), .ZN(n1265) );
XOR2_X1 U1038 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U1039 ( .A(n1120), .B(n1125), .ZN(n1298) );
XNOR2_X1 U1040 ( .A(G101), .B(n1299), .ZN(n1125) );
NOR2_X1 U1041 ( .A1(KEYINPUT20), .A2(n1289), .ZN(n1299) );
XNOR2_X1 U1042 ( .A(G104), .B(G107), .ZN(n1289) );
XNOR2_X1 U1043 ( .A(n1076), .B(G131), .ZN(n1120) );
XNOR2_X1 U1044 ( .A(G134), .B(n1300), .ZN(n1076) );
XOR2_X1 U1045 ( .A(KEYINPUT23), .B(G137), .Z(n1300) );
XOR2_X1 U1046 ( .A(n1301), .B(n1302), .Z(n1297) );
NOR2_X1 U1047 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XOR2_X1 U1048 ( .A(KEYINPUT7), .B(n1305), .Z(n1304) );
NOR2_X1 U1049 ( .A1(G110), .A2(n1175), .ZN(n1305) );
AND2_X1 U1050 ( .A1(n1175), .A2(G110), .ZN(n1303) );
INV_X1 U1051 ( .A(G140), .ZN(n1175) );
XOR2_X1 U1052 ( .A(n1306), .B(n1133), .Z(n1301) );
AND2_X1 U1053 ( .A1(G227), .A2(n1045), .ZN(n1133) );
INV_X1 U1054 ( .A(G953), .ZN(n1045) );
NAND2_X1 U1055 ( .A1(KEYINPUT30), .A2(n1124), .ZN(n1306) );
XNOR2_X1 U1056 ( .A(n1241), .B(n1078), .ZN(n1124) );
NAND2_X1 U1057 ( .A1(KEYINPUT19), .A2(n1217), .ZN(n1078) );
INV_X1 U1058 ( .A(n1246), .ZN(n1217) );
XOR2_X1 U1059 ( .A(G128), .B(KEYINPUT59), .Z(n1246) );
XNOR2_X1 U1060 ( .A(G143), .B(n1209), .ZN(n1241) );
XOR2_X1 U1061 ( .A(G146), .B(KEYINPUT35), .Z(n1209) );
endmodule


