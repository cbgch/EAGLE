//Key = 1001100011101111101011100100001010100100100011010010001111111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377;

XOR2_X1 U762 ( .A(n1048), .B(n1049), .Z(G9) );
NOR2_X1 U763 ( .A1(KEYINPUT48), .A2(n1050), .ZN(n1049) );
NOR2_X1 U764 ( .A1(n1051), .A2(n1052), .ZN(G75) );
NOR4_X1 U765 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NOR2_X1 U766 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U767 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
XOR2_X1 U768 ( .A(n1061), .B(KEYINPUT62), .Z(n1060) );
NAND4_X1 U769 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
NOR3_X1 U770 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1059) );
INV_X1 U771 ( .A(n1069), .ZN(n1068) );
NOR2_X1 U772 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
NOR2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1070) );
NOR2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND3_X1 U776 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1053) );
NAND3_X1 U777 ( .A1(n1065), .A2(n1081), .A3(n1062), .ZN(n1080) );
INV_X1 U778 ( .A(n1066), .ZN(n1062) );
NAND2_X1 U779 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND3_X1 U780 ( .A1(n1084), .A2(n1085), .A3(n1063), .ZN(n1083) );
NAND2_X1 U781 ( .A1(n1069), .A2(n1086), .ZN(n1082) );
NAND2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U783 ( .A1(n1089), .A2(n1090), .A3(n1084), .ZN(n1088) );
NAND2_X1 U784 ( .A1(n1063), .A2(n1091), .ZN(n1087) );
NAND2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XOR2_X1 U787 ( .A(n1096), .B(KEYINPUT50), .Z(n1094) );
NOR3_X1 U788 ( .A1(n1097), .A2(G953), .A3(n1098), .ZN(n1051) );
INV_X1 U789 ( .A(n1078), .ZN(n1098) );
NAND4_X1 U790 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1078) );
NOR3_X1 U791 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NOR3_X1 U792 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
NOR2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U794 ( .A1(G475), .A2(n1111), .ZN(n1109) );
NOR2_X1 U795 ( .A1(KEYINPUT13), .A2(G475), .ZN(n1107) );
INV_X1 U796 ( .A(KEYINPUT18), .ZN(n1106) );
NOR2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1104) );
NOR2_X1 U798 ( .A1(n1114), .A2(G475), .ZN(n1113) );
NOR2_X1 U799 ( .A1(KEYINPUT18), .A2(n1110), .ZN(n1114) );
INV_X1 U800 ( .A(KEYINPUT13), .ZN(n1110) );
NAND3_X1 U801 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1103) );
NOR3_X1 U802 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1101) );
XOR2_X1 U803 ( .A(n1121), .B(KEYINPUT58), .Z(n1120) );
NOR2_X1 U804 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
XNOR2_X1 U805 ( .A(n1124), .B(n1125), .ZN(n1099) );
XNOR2_X1 U806 ( .A(G952), .B(KEYINPUT32), .ZN(n1097) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(G72) );
NOR2_X1 U808 ( .A1(n1128), .A2(n1079), .ZN(n1127) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1126) );
NAND2_X1 U811 ( .A1(n1133), .A2(n1079), .ZN(n1132) );
XOR2_X1 U812 ( .A(n1134), .B(n1135), .Z(n1133) );
OR3_X1 U813 ( .A1(n1130), .A2(n1135), .A3(n1079), .ZN(n1131) );
XOR2_X1 U814 ( .A(n1136), .B(n1137), .Z(n1135) );
INV_X1 U815 ( .A(n1138), .ZN(n1137) );
XOR2_X1 U816 ( .A(n1139), .B(G140), .Z(n1136) );
NAND2_X1 U817 ( .A1(KEYINPUT57), .A2(n1140), .ZN(n1139) );
XOR2_X1 U818 ( .A(n1141), .B(n1142), .Z(G69) );
AND2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND3_X1 U820 ( .A1(n1145), .A2(n1146), .A3(n1143), .ZN(n1141) );
INV_X1 U821 ( .A(n1147), .ZN(n1143) );
NAND2_X1 U822 ( .A1(G953), .A2(n1148), .ZN(n1146) );
NAND2_X1 U823 ( .A1(n1149), .A2(n1079), .ZN(n1145) );
NAND2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XNOR2_X1 U825 ( .A(KEYINPUT22), .B(n1152), .ZN(n1151) );
NOR2_X1 U826 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U828 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
NOR3_X1 U829 ( .A1(n1153), .A2(n1159), .A3(n1160), .ZN(G63) );
NOR4_X1 U830 ( .A1(n1161), .A2(n1162), .A3(KEYINPUT23), .A4(n1163), .ZN(n1160) );
INV_X1 U831 ( .A(n1164), .ZN(n1161) );
NOR2_X1 U832 ( .A1(n1164), .A2(n1165), .ZN(n1159) );
NOR3_X1 U833 ( .A1(n1162), .A2(n1166), .A3(n1163), .ZN(n1165) );
AND2_X1 U834 ( .A1(n1167), .A2(KEYINPUT23), .ZN(n1166) );
NOR2_X1 U835 ( .A1(KEYINPUT11), .A2(n1167), .ZN(n1164) );
NOR2_X1 U836 ( .A1(n1168), .A2(n1169), .ZN(G60) );
XOR2_X1 U837 ( .A(KEYINPUT42), .B(n1153), .Z(n1169) );
NOR3_X1 U838 ( .A1(n1170), .A2(n1112), .A3(n1171), .ZN(n1168) );
NOR2_X1 U839 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
AND2_X1 U840 ( .A1(n1054), .A2(G475), .ZN(n1172) );
XOR2_X1 U841 ( .A(n1174), .B(KEYINPUT47), .Z(n1170) );
NAND3_X1 U842 ( .A1(n1157), .A2(G475), .A3(n1173), .ZN(n1174) );
XNOR2_X1 U843 ( .A(G104), .B(n1175), .ZN(G6) );
NOR2_X1 U844 ( .A1(n1153), .A2(n1176), .ZN(G57) );
XOR2_X1 U845 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U846 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U847 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U849 ( .A(KEYINPUT12), .B(n1185), .Z(n1181) );
NOR2_X1 U850 ( .A1(n1184), .A2(n1183), .ZN(n1185) );
XNOR2_X1 U851 ( .A(G113), .B(n1186), .ZN(n1183) );
XNOR2_X1 U852 ( .A(n1187), .B(n1188), .ZN(n1184) );
NAND2_X1 U853 ( .A1(KEYINPUT59), .A2(n1189), .ZN(n1187) );
NAND2_X1 U854 ( .A1(n1157), .A2(G472), .ZN(n1179) );
XNOR2_X1 U855 ( .A(n1190), .B(n1191), .ZN(n1177) );
INV_X1 U856 ( .A(G101), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1153), .A2(n1192), .ZN(G54) );
XOR2_X1 U858 ( .A(n1193), .B(n1194), .Z(n1192) );
XNOR2_X1 U859 ( .A(n1195), .B(n1196), .ZN(n1194) );
XOR2_X1 U860 ( .A(KEYINPUT14), .B(G140), .Z(n1196) );
XNOR2_X1 U861 ( .A(n1138), .B(n1197), .ZN(n1193) );
XOR2_X1 U862 ( .A(n1198), .B(n1199), .Z(n1197) );
NAND2_X1 U863 ( .A1(n1157), .A2(G469), .ZN(n1198) );
INV_X1 U864 ( .A(n1162), .ZN(n1157) );
XNOR2_X1 U865 ( .A(n1200), .B(n1201), .ZN(n1138) );
NOR2_X1 U866 ( .A1(n1153), .A2(n1202), .ZN(G51) );
XOR2_X1 U867 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U868 ( .A(n1205), .B(n1144), .Z(n1204) );
NAND2_X1 U869 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U870 ( .A1(n1188), .A2(G125), .ZN(n1207) );
XOR2_X1 U871 ( .A(n1208), .B(KEYINPUT33), .Z(n1206) );
OR2_X1 U872 ( .A1(n1188), .A2(G125), .ZN(n1208) );
XOR2_X1 U873 ( .A(n1209), .B(n1210), .Z(n1203) );
XOR2_X1 U874 ( .A(KEYINPUT20), .B(n1211), .Z(n1210) );
OR2_X1 U875 ( .A1(n1162), .A2(n1125), .ZN(n1209) );
NAND2_X1 U876 ( .A1(G902), .A2(n1054), .ZN(n1162) );
NAND3_X1 U877 ( .A1(n1150), .A2(n1152), .A3(n1134), .ZN(n1054) );
AND4_X1 U878 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1134) );
AND3_X1 U879 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
OR2_X1 U880 ( .A1(n1219), .A2(n1058), .ZN(n1214) );
NAND3_X1 U881 ( .A1(n1220), .A2(n1221), .A3(n1064), .ZN(n1213) );
NAND2_X1 U882 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
NAND3_X1 U883 ( .A1(n1076), .A2(n1224), .A3(n1084), .ZN(n1223) );
NAND3_X1 U884 ( .A1(n1077), .A2(n1225), .A3(n1063), .ZN(n1222) );
NAND2_X1 U885 ( .A1(n1226), .A2(n1227), .ZN(n1212) );
NAND2_X1 U886 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U887 ( .A1(n1084), .A2(n1069), .ZN(n1229) );
NAND2_X1 U888 ( .A1(n1085), .A2(n1225), .ZN(n1228) );
AND4_X1 U889 ( .A1(n1230), .A2(n1231), .A3(n1175), .A4(n1232), .ZN(n1150) );
NOR4_X1 U890 ( .A1(n1048), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1232) );
AND3_X1 U891 ( .A1(n1065), .A2(n1236), .A3(n1085), .ZN(n1048) );
NAND3_X1 U892 ( .A1(n1065), .A2(n1236), .A3(n1064), .ZN(n1175) );
AND2_X1 U893 ( .A1(n1237), .A2(n1056), .ZN(n1153) );
INV_X1 U894 ( .A(G952), .ZN(n1056) );
XNOR2_X1 U895 ( .A(KEYINPUT1), .B(n1079), .ZN(n1237) );
XNOR2_X1 U896 ( .A(G146), .B(n1216), .ZN(G48) );
NAND3_X1 U897 ( .A1(n1064), .A2(n1225), .A3(n1226), .ZN(n1216) );
INV_X1 U898 ( .A(n1238), .ZN(n1226) );
XOR2_X1 U899 ( .A(n1239), .B(G143), .Z(G45) );
NAND2_X1 U900 ( .A1(KEYINPUT0), .A2(n1217), .ZN(n1239) );
NAND4_X1 U901 ( .A1(n1240), .A2(n1076), .A3(n1241), .A4(n1225), .ZN(n1217) );
NOR2_X1 U902 ( .A1(n1100), .A2(n1242), .ZN(n1241) );
XNOR2_X1 U903 ( .A(G140), .B(n1218), .ZN(G42) );
NAND4_X1 U904 ( .A1(n1084), .A2(n1077), .A3(n1240), .A4(n1064), .ZN(n1218) );
XNOR2_X1 U905 ( .A(G137), .B(n1243), .ZN(G39) );
NAND4_X1 U906 ( .A1(n1244), .A2(n1245), .A3(n1084), .A4(n1221), .ZN(n1243) );
XNOR2_X1 U907 ( .A(n1224), .B(KEYINPUT34), .ZN(n1244) );
XNOR2_X1 U908 ( .A(G134), .B(n1246), .ZN(G36) );
NAND2_X1 U909 ( .A1(n1247), .A2(n1084), .ZN(n1246) );
XOR2_X1 U910 ( .A(n1219), .B(KEYINPUT37), .Z(n1247) );
NAND3_X1 U911 ( .A1(n1076), .A2(n1085), .A3(n1240), .ZN(n1219) );
XNOR2_X1 U912 ( .A(n1248), .B(n1249), .ZN(G33) );
NOR2_X1 U913 ( .A1(n1250), .A2(n1058), .ZN(n1249) );
INV_X1 U914 ( .A(n1084), .ZN(n1058) );
NOR2_X1 U915 ( .A1(n1096), .A2(n1095), .ZN(n1084) );
INV_X1 U916 ( .A(n1115), .ZN(n1095) );
XOR2_X1 U917 ( .A(n1251), .B(KEYINPUT35), .Z(n1250) );
NAND3_X1 U918 ( .A1(n1240), .A2(n1064), .A3(n1252), .ZN(n1251) );
XNOR2_X1 U919 ( .A(n1076), .B(KEYINPUT9), .ZN(n1252) );
XOR2_X1 U920 ( .A(G128), .B(n1253), .Z(G30) );
NOR4_X1 U921 ( .A1(KEYINPUT5), .A2(n1092), .A3(n1254), .A4(n1238), .ZN(n1253) );
NAND3_X1 U922 ( .A1(n1255), .A2(n1256), .A3(n1240), .ZN(n1238) );
NOR2_X1 U923 ( .A1(n1072), .A2(n1257), .ZN(n1240) );
XNOR2_X1 U924 ( .A(G101), .B(n1258), .ZN(G3) );
NAND2_X1 U925 ( .A1(KEYINPUT55), .A2(n1259), .ZN(n1258) );
INV_X1 U926 ( .A(n1152), .ZN(n1259) );
NAND3_X1 U927 ( .A1(n1236), .A2(n1069), .A3(n1076), .ZN(n1152) );
XNOR2_X1 U928 ( .A(G125), .B(n1260), .ZN(G27) );
NAND4_X1 U929 ( .A1(n1063), .A2(n1064), .A3(n1261), .A4(n1262), .ZN(n1260) );
NOR3_X1 U930 ( .A1(n1092), .A2(KEYINPUT41), .A3(n1257), .ZN(n1262) );
INV_X1 U931 ( .A(n1221), .ZN(n1257) );
NAND2_X1 U932 ( .A1(n1066), .A2(n1263), .ZN(n1221) );
NAND4_X1 U933 ( .A1(G902), .A2(G953), .A3(n1264), .A4(n1130), .ZN(n1263) );
INV_X1 U934 ( .A(G900), .ZN(n1130) );
XNOR2_X1 U935 ( .A(n1077), .B(KEYINPUT15), .ZN(n1261) );
XNOR2_X1 U936 ( .A(G122), .B(n1230), .ZN(G24) );
NAND4_X1 U937 ( .A1(n1265), .A2(n1065), .A3(n1266), .A4(n1267), .ZN(n1230) );
INV_X1 U938 ( .A(n1073), .ZN(n1065) );
NAND2_X1 U939 ( .A1(n1268), .A2(n1269), .ZN(n1073) );
XNOR2_X1 U940 ( .A(G119), .B(n1231), .ZN(G21) );
NAND2_X1 U941 ( .A1(n1245), .A2(n1265), .ZN(n1231) );
AND3_X1 U942 ( .A1(n1069), .A2(n1256), .A3(n1255), .ZN(n1245) );
XNOR2_X1 U943 ( .A(n1270), .B(n1235), .ZN(G18) );
AND3_X1 U944 ( .A1(n1076), .A2(n1085), .A3(n1265), .ZN(n1235) );
INV_X1 U945 ( .A(n1254), .ZN(n1085) );
NAND2_X1 U946 ( .A1(n1271), .A2(n1267), .ZN(n1254) );
XNOR2_X1 U947 ( .A(n1272), .B(n1266), .ZN(n1271) );
INV_X1 U948 ( .A(n1242), .ZN(n1266) );
XOR2_X1 U949 ( .A(G113), .B(n1234), .Z(G15) );
AND3_X1 U950 ( .A1(n1076), .A2(n1064), .A3(n1265), .ZN(n1234) );
AND2_X1 U951 ( .A1(n1063), .A2(n1273), .ZN(n1265) );
INV_X1 U952 ( .A(n1075), .ZN(n1063) );
NAND2_X1 U953 ( .A1(n1089), .A2(n1274), .ZN(n1075) );
XNOR2_X1 U954 ( .A(KEYINPUT10), .B(n1117), .ZN(n1274) );
INV_X1 U955 ( .A(n1118), .ZN(n1089) );
AND2_X1 U956 ( .A1(n1269), .A2(n1256), .ZN(n1076) );
XNOR2_X1 U957 ( .A(n1255), .B(KEYINPUT49), .ZN(n1269) );
XNOR2_X1 U958 ( .A(n1195), .B(n1233), .ZN(G12) );
AND3_X1 U959 ( .A1(n1236), .A2(n1069), .A3(n1077), .ZN(n1233) );
AND2_X1 U960 ( .A1(n1268), .A2(n1255), .ZN(n1077) );
XOR2_X1 U961 ( .A(n1121), .B(n1275), .Z(n1255) );
XOR2_X1 U962 ( .A(KEYINPUT24), .B(KEYINPUT16), .Z(n1275) );
XOR2_X1 U963 ( .A(n1276), .B(n1158), .Z(n1121) );
AND2_X1 U964 ( .A1(G217), .A2(n1277), .ZN(n1158) );
NAND2_X1 U965 ( .A1(n1156), .A2(n1278), .ZN(n1276) );
XOR2_X1 U966 ( .A(n1279), .B(n1280), .Z(n1156) );
XNOR2_X1 U967 ( .A(n1281), .B(n1282), .ZN(n1279) );
NOR2_X1 U968 ( .A1(KEYINPUT28), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U969 ( .A(n1284), .B(n1285), .ZN(n1283) );
NAND2_X1 U970 ( .A1(G221), .A2(n1286), .ZN(n1284) );
INV_X1 U971 ( .A(n1287), .ZN(n1286) );
NOR2_X1 U972 ( .A1(KEYINPUT36), .A2(n1288), .ZN(n1281) );
XOR2_X1 U973 ( .A(G128), .B(n1289), .Z(n1288) );
INV_X1 U974 ( .A(n1256), .ZN(n1268) );
NAND3_X1 U975 ( .A1(n1290), .A2(n1291), .A3(n1116), .ZN(n1256) );
NAND2_X1 U976 ( .A1(n1122), .A2(n1123), .ZN(n1116) );
NAND2_X1 U977 ( .A1(KEYINPUT63), .A2(n1123), .ZN(n1291) );
OR3_X1 U978 ( .A1(n1122), .A2(KEYINPUT63), .A3(n1123), .ZN(n1290) );
INV_X1 U979 ( .A(G472), .ZN(n1123) );
AND2_X1 U980 ( .A1(n1292), .A2(n1278), .ZN(n1122) );
XOR2_X1 U981 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U982 ( .A(n1295), .B(n1296), .Z(n1294) );
NAND2_X1 U983 ( .A1(n1297), .A2(KEYINPUT45), .ZN(n1295) );
XOR2_X1 U984 ( .A(n1298), .B(n1299), .Z(n1297) );
XNOR2_X1 U985 ( .A(n1201), .B(n1300), .ZN(n1299) );
XOR2_X1 U986 ( .A(G128), .B(n1301), .Z(n1201) );
XOR2_X1 U987 ( .A(KEYINPUT6), .B(KEYINPUT14), .Z(n1298) );
XOR2_X1 U988 ( .A(n1190), .B(n1186), .Z(n1293) );
NOR2_X1 U989 ( .A1(KEYINPUT2), .A2(n1302), .ZN(n1186) );
XNOR2_X1 U990 ( .A(G119), .B(G116), .ZN(n1302) );
NAND3_X1 U991 ( .A1(n1303), .A2(n1079), .A3(G210), .ZN(n1190) );
NAND2_X1 U992 ( .A1(n1304), .A2(n1305), .ZN(n1069) );
NAND2_X1 U993 ( .A1(n1064), .A2(n1272), .ZN(n1305) );
INV_X1 U994 ( .A(KEYINPUT3), .ZN(n1272) );
NOR2_X1 U995 ( .A1(n1267), .A2(n1242), .ZN(n1064) );
NAND3_X1 U996 ( .A1(n1242), .A2(n1100), .A3(KEYINPUT3), .ZN(n1304) );
INV_X1 U997 ( .A(n1267), .ZN(n1100) );
XOR2_X1 U998 ( .A(n1306), .B(n1163), .Z(n1267) );
INV_X1 U999 ( .A(G478), .ZN(n1163) );
NAND2_X1 U1000 ( .A1(n1307), .A2(n1278), .ZN(n1306) );
XNOR2_X1 U1001 ( .A(KEYINPUT19), .B(n1167), .ZN(n1307) );
XOR2_X1 U1002 ( .A(n1308), .B(n1309), .Z(n1167) );
XNOR2_X1 U1003 ( .A(n1310), .B(n1311), .ZN(n1309) );
NAND2_X1 U1004 ( .A1(KEYINPUT30), .A2(n1312), .ZN(n1310) );
INV_X1 U1005 ( .A(G134), .ZN(n1312) );
XOR2_X1 U1006 ( .A(n1313), .B(n1314), .Z(n1308) );
NOR3_X1 U1007 ( .A1(n1315), .A2(KEYINPUT46), .A3(n1287), .ZN(n1314) );
NAND2_X1 U1008 ( .A1(G234), .A2(n1079), .ZN(n1287) );
INV_X1 U1009 ( .A(G217), .ZN(n1315) );
XOR2_X1 U1010 ( .A(n1316), .B(G128), .Z(n1313) );
NAND2_X1 U1011 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND3_X1 U1012 ( .A1(n1270), .A2(n1319), .A3(n1320), .ZN(n1318) );
XNOR2_X1 U1013 ( .A(n1321), .B(n1050), .ZN(n1320) );
NAND2_X1 U1014 ( .A1(G122), .A2(n1322), .ZN(n1321) );
INV_X1 U1015 ( .A(KEYINPUT61), .ZN(n1322) );
NAND2_X1 U1016 ( .A1(n1323), .A2(n1324), .ZN(n1317) );
NAND2_X1 U1017 ( .A1(n1270), .A2(n1319), .ZN(n1324) );
INV_X1 U1018 ( .A(KEYINPUT26), .ZN(n1319) );
XNOR2_X1 U1019 ( .A(G107), .B(n1325), .ZN(n1323) );
NOR2_X1 U1020 ( .A1(G122), .A2(KEYINPUT61), .ZN(n1325) );
XOR2_X1 U1021 ( .A(n1111), .B(G475), .Z(n1242) );
INV_X1 U1022 ( .A(n1112), .ZN(n1111) );
NOR2_X1 U1023 ( .A1(n1173), .A2(G902), .ZN(n1112) );
XOR2_X1 U1024 ( .A(n1326), .B(n1327), .Z(n1173) );
XOR2_X1 U1025 ( .A(n1328), .B(n1280), .Z(n1327) );
XNOR2_X1 U1026 ( .A(n1140), .B(n1329), .ZN(n1280) );
XOR2_X1 U1027 ( .A(G146), .B(G140), .Z(n1329) );
NOR2_X1 U1028 ( .A1(KEYINPUT38), .A2(n1330), .ZN(n1328) );
NOR2_X1 U1029 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1030 ( .A(n1333), .B(KEYINPUT44), .Z(n1332) );
NAND2_X1 U1031 ( .A1(n1334), .A2(n1248), .ZN(n1333) );
NOR2_X1 U1032 ( .A1(n1334), .A2(n1248), .ZN(n1331) );
INV_X1 U1033 ( .A(G131), .ZN(n1248) );
XNOR2_X1 U1034 ( .A(n1335), .B(n1336), .ZN(n1334) );
NAND3_X1 U1035 ( .A1(n1303), .A2(n1079), .A3(n1337), .ZN(n1335) );
XOR2_X1 U1036 ( .A(KEYINPUT29), .B(G214), .Z(n1337) );
XNOR2_X1 U1037 ( .A(G104), .B(n1338), .ZN(n1326) );
XOR2_X1 U1038 ( .A(G122), .B(G113), .Z(n1338) );
AND2_X1 U1039 ( .A1(n1273), .A2(n1224), .ZN(n1236) );
INV_X1 U1040 ( .A(n1072), .ZN(n1224) );
NAND2_X1 U1041 ( .A1(n1339), .A2(n1118), .ZN(n1072) );
XNOR2_X1 U1042 ( .A(n1340), .B(G469), .ZN(n1118) );
NAND2_X1 U1043 ( .A1(n1341), .A2(n1278), .ZN(n1340) );
XOR2_X1 U1044 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1045 ( .A(n1344), .B(n1345), .Z(n1343) );
XOR2_X1 U1046 ( .A(G128), .B(n1346), .Z(n1345) );
NOR2_X1 U1047 ( .A1(KEYINPUT27), .A2(n1189), .ZN(n1346) );
XOR2_X1 U1048 ( .A(KEYINPUT14), .B(n1301), .Z(n1189) );
XNOR2_X1 U1049 ( .A(n1347), .B(n1285), .ZN(n1301) );
XOR2_X1 U1050 ( .A(G137), .B(KEYINPUT60), .Z(n1285) );
XNOR2_X1 U1051 ( .A(G134), .B(G131), .ZN(n1347) );
XOR2_X1 U1052 ( .A(KEYINPUT54), .B(G140), .Z(n1344) );
XOR2_X1 U1053 ( .A(n1199), .B(n1348), .Z(n1342) );
XOR2_X1 U1054 ( .A(n1349), .B(n1200), .Z(n1348) );
XNOR2_X1 U1055 ( .A(KEYINPUT8), .B(n1350), .ZN(n1200) );
NOR2_X1 U1056 ( .A1(KEYINPUT52), .A2(n1351), .ZN(n1350) );
XNOR2_X1 U1057 ( .A(G146), .B(n1311), .ZN(n1351) );
NAND2_X1 U1058 ( .A1(KEYINPUT25), .A2(n1195), .ZN(n1349) );
XOR2_X1 U1059 ( .A(n1352), .B(n1353), .Z(n1199) );
XOR2_X1 U1060 ( .A(n1354), .B(n1355), .Z(n1353) );
NOR2_X1 U1061 ( .A1(G953), .A2(n1129), .ZN(n1355) );
INV_X1 U1062 ( .A(G227), .ZN(n1129) );
NOR2_X1 U1063 ( .A1(KEYINPUT31), .A2(n1050), .ZN(n1354) );
INV_X1 U1064 ( .A(G107), .ZN(n1050) );
XNOR2_X1 U1065 ( .A(G101), .B(G104), .ZN(n1352) );
XNOR2_X1 U1066 ( .A(n1090), .B(KEYINPUT17), .ZN(n1339) );
INV_X1 U1067 ( .A(n1117), .ZN(n1090) );
NAND2_X1 U1068 ( .A1(G221), .A2(n1277), .ZN(n1117) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1278), .ZN(n1277) );
AND2_X1 U1070 ( .A1(n1225), .A2(n1356), .ZN(n1273) );
NAND2_X1 U1071 ( .A1(n1066), .A2(n1357), .ZN(n1356) );
NAND3_X1 U1072 ( .A1(n1147), .A2(n1264), .A3(G902), .ZN(n1357) );
NOR2_X1 U1073 ( .A1(G898), .A2(n1079), .ZN(n1147) );
NAND3_X1 U1074 ( .A1(n1264), .A2(n1079), .A3(G952), .ZN(n1066) );
INV_X1 U1075 ( .A(G953), .ZN(n1079) );
NAND2_X1 U1076 ( .A1(G237), .A2(G234), .ZN(n1264) );
INV_X1 U1077 ( .A(n1092), .ZN(n1225) );
NAND2_X1 U1078 ( .A1(n1096), .A2(n1115), .ZN(n1092) );
NAND2_X1 U1079 ( .A1(G214), .A2(n1358), .ZN(n1115) );
NAND2_X1 U1080 ( .A1(n1359), .A2(n1360), .ZN(n1096) );
OR2_X1 U1081 ( .A1(n1125), .A2(n1361), .ZN(n1360) );
XOR2_X1 U1082 ( .A(n1362), .B(KEYINPUT53), .Z(n1359) );
NAND2_X1 U1083 ( .A1(n1361), .A2(n1125), .ZN(n1362) );
NAND2_X1 U1084 ( .A1(G210), .A2(n1358), .ZN(n1125) );
NAND2_X1 U1085 ( .A1(n1303), .A2(n1278), .ZN(n1358) );
INV_X1 U1086 ( .A(G237), .ZN(n1303) );
XNOR2_X1 U1087 ( .A(n1124), .B(KEYINPUT51), .ZN(n1361) );
NAND2_X1 U1088 ( .A1(n1363), .A2(n1278), .ZN(n1124) );
INV_X1 U1089 ( .A(G902), .ZN(n1278) );
XNOR2_X1 U1090 ( .A(n1211), .B(n1364), .ZN(n1363) );
XNOR2_X1 U1091 ( .A(n1365), .B(n1366), .ZN(n1364) );
NOR2_X1 U1092 ( .A1(KEYINPUT43), .A2(n1144), .ZN(n1366) );
XNOR2_X1 U1093 ( .A(n1367), .B(n1368), .ZN(n1144) );
XNOR2_X1 U1094 ( .A(n1270), .B(n1369), .ZN(n1368) );
XOR2_X1 U1095 ( .A(KEYINPUT21), .B(G122), .Z(n1369) );
INV_X1 U1096 ( .A(G116), .ZN(n1270) );
XOR2_X1 U1097 ( .A(n1296), .B(n1370), .Z(n1367) );
XOR2_X1 U1098 ( .A(n1371), .B(n1289), .Z(n1370) );
XOR2_X1 U1099 ( .A(G119), .B(G110), .Z(n1289) );
NOR2_X1 U1100 ( .A1(KEYINPUT39), .A2(n1372), .ZN(n1371) );
XOR2_X1 U1101 ( .A(G104), .B(n1373), .Z(n1372) );
NOR2_X1 U1102 ( .A1(G107), .A2(KEYINPUT7), .ZN(n1373) );
XNOR2_X1 U1103 ( .A(G101), .B(G113), .ZN(n1296) );
NAND2_X1 U1104 ( .A1(n1374), .A2(KEYINPUT40), .ZN(n1365) );
XNOR2_X1 U1105 ( .A(n1140), .B(n1188), .ZN(n1374) );
XNOR2_X1 U1106 ( .A(n1300), .B(G128), .ZN(n1188) );
NAND2_X1 U1107 ( .A1(n1375), .A2(n1376), .ZN(n1300) );
NAND2_X1 U1108 ( .A1(n1377), .A2(n1336), .ZN(n1376) );
INV_X1 U1109 ( .A(n1311), .ZN(n1336) );
XOR2_X1 U1110 ( .A(KEYINPUT56), .B(G146), .Z(n1377) );
NAND2_X1 U1111 ( .A1(G146), .A2(n1311), .ZN(n1375) );
XOR2_X1 U1112 ( .A(G143), .B(KEYINPUT4), .Z(n1311) );
INV_X1 U1113 ( .A(G125), .ZN(n1140) );
NOR2_X1 U1114 ( .A1(n1148), .A2(G953), .ZN(n1211) );
INV_X1 U1115 ( .A(G224), .ZN(n1148) );
INV_X1 U1116 ( .A(G110), .ZN(n1195) );
endmodule


