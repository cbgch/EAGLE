//Key = 1101011100110100011010100111110001101011001111010011100100011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
n1503;

XOR2_X1 U809 ( .A(G107), .B(n1133), .Z(G9) );
NOR2_X1 U810 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(G75) );
NOR4_X1 U812 ( .A1(n1138), .A2(n1139), .A3(G953), .A4(n1140), .ZN(n1137) );
NOR2_X1 U813 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NOR2_X1 U814 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NOR2_X1 U815 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR2_X1 U816 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
NOR2_X1 U817 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U818 ( .A1(n1151), .A2(n1152), .ZN(n1147) );
NOR2_X1 U819 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
NOR3_X1 U821 ( .A1(n1149), .A2(n1152), .A3(n1135), .ZN(n1143) );
NAND3_X1 U822 ( .A1(G952), .A2(n1157), .A3(n1158), .ZN(n1138) );
NAND2_X1 U823 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND4_X1 U824 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
NAND2_X1 U825 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U826 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
OR3_X1 U827 ( .A1(n1152), .A2(KEYINPUT24), .A3(n1169), .ZN(n1168) );
NAND3_X1 U828 ( .A1(n1170), .A2(n1171), .A3(KEYINPUT42), .ZN(n1167) );
NAND4_X1 U829 ( .A1(n1172), .A2(n1170), .A3(n1173), .A4(n1174), .ZN(n1163) );
NAND2_X1 U830 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U831 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U832 ( .A1(n1179), .A2(n1180), .ZN(n1162) );
INV_X1 U833 ( .A(KEYINPUT42), .ZN(n1180) );
NAND3_X1 U834 ( .A1(n1181), .A2(n1170), .A3(n1172), .ZN(n1179) );
NAND2_X1 U835 ( .A1(KEYINPUT24), .A2(n1182), .ZN(n1161) );
NAND3_X1 U836 ( .A1(n1183), .A2(n1173), .A3(n1165), .ZN(n1182) );
INV_X1 U837 ( .A(n1142), .ZN(n1165) );
NAND2_X1 U838 ( .A1(n1172), .A2(n1184), .ZN(n1142) );
INV_X1 U839 ( .A(n1185), .ZN(n1172) );
NOR3_X1 U840 ( .A1(n1186), .A2(G953), .A3(n1140), .ZN(n1136) );
AND4_X1 U841 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1140) );
NOR4_X1 U842 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1177), .ZN(n1190) );
NAND2_X1 U843 ( .A1(n1194), .A2(n1195), .ZN(n1191) );
NOR3_X1 U844 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1189) );
XOR2_X1 U845 ( .A(n1199), .B(n1200), .Z(n1198) );
NAND2_X1 U846 ( .A1(KEYINPUT6), .A2(n1201), .ZN(n1199) );
XOR2_X1 U847 ( .A(KEYINPUT29), .B(G478), .Z(n1201) );
XOR2_X1 U848 ( .A(n1202), .B(KEYINPUT63), .Z(n1197) );
NAND3_X1 U849 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
OR2_X1 U850 ( .A1(n1206), .A2(KEYINPUT7), .ZN(n1204) );
NAND3_X1 U851 ( .A1(n1207), .A2(n1206), .A3(KEYINPUT7), .ZN(n1203) );
XOR2_X1 U852 ( .A(n1208), .B(KEYINPUT62), .Z(n1187) );
XOR2_X1 U853 ( .A(KEYINPUT16), .B(G952), .Z(n1186) );
XOR2_X1 U854 ( .A(n1209), .B(n1210), .Z(G72) );
XOR2_X1 U855 ( .A(n1211), .B(n1212), .Z(n1210) );
NOR2_X1 U856 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NOR2_X1 U857 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
NAND2_X1 U858 ( .A1(n1217), .A2(n1218), .ZN(n1211) );
NAND2_X1 U859 ( .A1(G953), .A2(n1216), .ZN(n1218) );
XOR2_X1 U860 ( .A(n1219), .B(n1220), .Z(n1217) );
XOR2_X1 U861 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U862 ( .A(n1223), .B(n1224), .Z(n1219) );
XOR2_X1 U863 ( .A(n1225), .B(KEYINPUT0), .Z(n1223) );
NAND2_X1 U864 ( .A1(n1214), .A2(n1226), .ZN(n1209) );
NAND2_X1 U865 ( .A1(n1227), .A2(n1228), .ZN(G69) );
NAND2_X1 U866 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND2_X1 U867 ( .A1(G953), .A2(n1231), .ZN(n1230) );
INV_X1 U868 ( .A(n1232), .ZN(n1229) );
NAND3_X1 U869 ( .A1(G953), .A2(n1233), .A3(n1232), .ZN(n1227) );
XOR2_X1 U870 ( .A(n1234), .B(n1235), .Z(n1232) );
NOR4_X1 U871 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NOR3_X1 U872 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
NOR2_X1 U873 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NOR2_X1 U874 ( .A1(n1245), .A2(n1246), .ZN(n1241) );
NOR2_X1 U875 ( .A1(G898), .A2(n1214), .ZN(n1238) );
NOR3_X1 U876 ( .A1(n1244), .A2(n1247), .A3(n1243), .ZN(n1237) );
INV_X1 U877 ( .A(KEYINPUT5), .ZN(n1243) );
NOR3_X1 U878 ( .A1(n1246), .A2(n1245), .A3(n1248), .ZN(n1236) );
AND2_X1 U879 ( .A1(KEYINPUT5), .A2(n1249), .ZN(n1245) );
NAND2_X1 U880 ( .A1(n1250), .A2(n1214), .ZN(n1234) );
XOR2_X1 U881 ( .A(n1251), .B(KEYINPUT41), .Z(n1250) );
NAND2_X1 U882 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U883 ( .A1(G898), .A2(G224), .ZN(n1233) );
NOR2_X1 U884 ( .A1(n1254), .A2(n1255), .ZN(G66) );
XOR2_X1 U885 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U886 ( .A1(KEYINPUT21), .A2(n1258), .ZN(n1257) );
NAND2_X1 U887 ( .A1(n1259), .A2(n1207), .ZN(n1256) );
NOR2_X1 U888 ( .A1(n1254), .A2(n1260), .ZN(G63) );
NOR3_X1 U889 ( .A1(n1200), .A2(n1261), .A3(n1262), .ZN(n1260) );
AND3_X1 U890 ( .A1(n1263), .A2(G478), .A3(n1259), .ZN(n1262) );
NOR2_X1 U891 ( .A1(n1264), .A2(n1263), .ZN(n1261) );
NOR2_X1 U892 ( .A1(n1158), .A2(n1265), .ZN(n1264) );
NOR2_X1 U893 ( .A1(n1254), .A2(n1266), .ZN(G60) );
XOR2_X1 U894 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U895 ( .A(n1269), .B(KEYINPUT53), .Z(n1267) );
NAND2_X1 U896 ( .A1(n1259), .A2(G475), .ZN(n1269) );
XOR2_X1 U897 ( .A(G104), .B(n1270), .Z(G6) );
NOR2_X1 U898 ( .A1(n1134), .A2(n1169), .ZN(n1270) );
NOR2_X1 U899 ( .A1(n1254), .A2(n1271), .ZN(G57) );
XOR2_X1 U900 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U901 ( .A(n1274), .B(n1240), .Z(n1273) );
NAND2_X1 U902 ( .A1(KEYINPUT52), .A2(n1275), .ZN(n1274) );
NAND2_X1 U903 ( .A1(n1259), .A2(G472), .ZN(n1275) );
XOR2_X1 U904 ( .A(n1276), .B(n1277), .Z(n1272) );
NOR2_X1 U905 ( .A1(KEYINPUT9), .A2(n1278), .ZN(n1277) );
XOR2_X1 U906 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U907 ( .A(KEYINPUT60), .B(n1281), .Z(n1280) );
NAND2_X1 U908 ( .A1(n1282), .A2(n1283), .ZN(n1276) );
INV_X1 U909 ( .A(n1284), .ZN(n1283) );
XOR2_X1 U910 ( .A(KEYINPUT33), .B(n1285), .Z(n1282) );
NOR2_X1 U911 ( .A1(n1254), .A2(n1286), .ZN(G54) );
XOR2_X1 U912 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U913 ( .A(n1289), .B(n1290), .Z(n1288) );
NAND3_X1 U914 ( .A1(G227), .A2(n1214), .A3(KEYINPUT34), .ZN(n1289) );
XOR2_X1 U915 ( .A(n1291), .B(n1292), .Z(n1287) );
NOR2_X1 U916 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U917 ( .A(n1295), .B(KEYINPUT50), .Z(n1294) );
NAND2_X1 U918 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NOR2_X1 U919 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
XOR2_X1 U920 ( .A(n1298), .B(n1222), .Z(n1297) );
NAND3_X1 U921 ( .A1(n1259), .A2(G469), .A3(KEYINPUT17), .ZN(n1291) );
NOR2_X1 U922 ( .A1(n1254), .A2(n1299), .ZN(G51) );
XOR2_X1 U923 ( .A(n1300), .B(n1301), .Z(n1299) );
NAND2_X1 U924 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U925 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
XOR2_X1 U926 ( .A(KEYINPUT20), .B(n1306), .Z(n1302) );
NOR2_X1 U927 ( .A1(n1304), .A2(n1305), .ZN(n1306) );
NAND2_X1 U928 ( .A1(n1307), .A2(n1308), .ZN(n1305) );
NAND2_X1 U929 ( .A1(G125), .A2(n1309), .ZN(n1308) );
NAND2_X1 U930 ( .A1(n1310), .A2(n1311), .ZN(n1307) );
XOR2_X1 U931 ( .A(n1309), .B(KEYINPUT51), .Z(n1310) );
XOR2_X1 U932 ( .A(n1312), .B(n1281), .Z(n1309) );
XNOR2_X1 U933 ( .A(n1313), .B(KEYINPUT31), .ZN(n1312) );
NAND2_X1 U934 ( .A1(n1259), .A2(G210), .ZN(n1300) );
NOR2_X1 U935 ( .A1(n1314), .A2(n1158), .ZN(n1259) );
AND3_X1 U936 ( .A1(n1315), .A2(n1252), .A3(n1316), .ZN(n1158) );
XNOR2_X1 U937 ( .A(n1253), .B(KEYINPUT59), .ZN(n1316) );
AND3_X1 U938 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(n1253) );
NAND2_X1 U939 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U940 ( .A1(n1322), .A2(n1169), .ZN(n1321) );
XOR2_X1 U941 ( .A(KEYINPUT38), .B(n1323), .Z(n1322) );
INV_X1 U942 ( .A(n1134), .ZN(n1320) );
NAND4_X1 U943 ( .A1(n1324), .A2(n1173), .A3(n1325), .A4(n1326), .ZN(n1134) );
NAND3_X1 U944 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1317) );
XOR2_X1 U945 ( .A(n1326), .B(KEYINPUT30), .Z(n1329) );
AND3_X1 U946 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1252) );
NAND2_X1 U947 ( .A1(n1325), .A2(n1333), .ZN(n1332) );
XOR2_X1 U948 ( .A(KEYINPUT14), .B(n1334), .Z(n1333) );
NAND2_X1 U949 ( .A1(n1335), .A2(n1336), .ZN(n1330) );
NAND2_X1 U950 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND3_X1 U951 ( .A1(n1196), .A2(n1339), .A3(n1340), .ZN(n1338) );
XOR2_X1 U952 ( .A(KEYINPUT49), .B(n1170), .Z(n1340) );
NAND2_X1 U953 ( .A1(n1171), .A2(n1323), .ZN(n1337) );
INV_X1 U954 ( .A(n1226), .ZN(n1315) );
NAND4_X1 U955 ( .A1(n1341), .A2(n1342), .A3(n1343), .A4(n1344), .ZN(n1226) );
NOR4_X1 U956 ( .A1(n1345), .A2(n1346), .A3(n1347), .A4(n1348), .ZN(n1344) );
INV_X1 U957 ( .A(n1349), .ZN(n1346) );
NOR2_X1 U958 ( .A1(n1350), .A2(n1351), .ZN(n1343) );
INV_X1 U959 ( .A(n1352), .ZN(n1350) );
NAND3_X1 U960 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1342) );
INV_X1 U961 ( .A(n1356), .ZN(n1355) );
OR2_X1 U962 ( .A1(n1357), .A2(KEYINPUT32), .ZN(n1354) );
NAND2_X1 U963 ( .A1(KEYINPUT32), .A2(n1358), .ZN(n1353) );
OR3_X1 U964 ( .A1(n1149), .A2(n1175), .A3(n1359), .ZN(n1358) );
INV_X1 U965 ( .A(n1159), .ZN(n1149) );
NOR2_X1 U966 ( .A1(n1214), .A2(G952), .ZN(n1254) );
XOR2_X1 U967 ( .A(G146), .B(n1351), .Z(G48) );
AND2_X1 U968 ( .A1(n1360), .A2(n1183), .ZN(n1351) );
XOR2_X1 U969 ( .A(n1361), .B(n1362), .Z(G45) );
NAND2_X1 U970 ( .A1(KEYINPUT45), .A2(n1363), .ZN(n1362) );
INV_X1 U971 ( .A(n1341), .ZN(n1363) );
NAND3_X1 U972 ( .A1(n1171), .A2(n1364), .A3(n1365), .ZN(n1341) );
NOR3_X1 U973 ( .A1(n1175), .A2(n1366), .A3(n1367), .ZN(n1365) );
INV_X1 U974 ( .A(n1324), .ZN(n1175) );
XOR2_X1 U975 ( .A(n1368), .B(n1345), .Z(G42) );
NOR3_X1 U976 ( .A1(n1150), .A2(n1169), .A3(n1369), .ZN(n1345) );
NAND2_X1 U977 ( .A1(KEYINPUT27), .A2(n1370), .ZN(n1368) );
XOR2_X1 U978 ( .A(G137), .B(n1371), .Z(G39) );
NOR2_X1 U979 ( .A1(n1369), .A2(n1356), .ZN(n1371) );
NAND2_X1 U980 ( .A1(n1372), .A2(n1373), .ZN(G36) );
NAND2_X1 U981 ( .A1(G134), .A2(n1352), .ZN(n1373) );
XOR2_X1 U982 ( .A(n1374), .B(KEYINPUT35), .Z(n1372) );
OR2_X1 U983 ( .A1(n1352), .A2(G134), .ZN(n1374) );
NAND3_X1 U984 ( .A1(n1357), .A2(n1323), .A3(n1171), .ZN(n1352) );
NAND2_X1 U985 ( .A1(n1375), .A2(n1376), .ZN(G33) );
NAND2_X1 U986 ( .A1(n1348), .A2(n1225), .ZN(n1376) );
INV_X1 U987 ( .A(n1377), .ZN(n1348) );
XOR2_X1 U988 ( .A(n1378), .B(KEYINPUT40), .Z(n1375) );
NAND2_X1 U989 ( .A1(G131), .A2(n1377), .ZN(n1378) );
NAND3_X1 U990 ( .A1(n1357), .A2(n1183), .A3(n1171), .ZN(n1377) );
INV_X1 U991 ( .A(n1369), .ZN(n1357) );
NAND3_X1 U992 ( .A1(n1324), .A2(n1359), .A3(n1159), .ZN(n1369) );
NOR2_X1 U993 ( .A1(n1155), .A2(n1192), .ZN(n1159) );
XNOR2_X1 U994 ( .A(n1188), .B(KEYINPUT8), .ZN(n1155) );
XOR2_X1 U995 ( .A(G128), .B(n1347), .Z(G30) );
AND2_X1 U996 ( .A1(n1360), .A2(n1323), .ZN(n1347) );
AND4_X1 U997 ( .A1(n1364), .A2(n1324), .A3(n1196), .A4(n1339), .ZN(n1360) );
XOR2_X1 U998 ( .A(n1379), .B(n1318), .Z(G3) );
NAND3_X1 U999 ( .A1(n1171), .A2(n1326), .A3(n1327), .ZN(n1318) );
INV_X1 U1000 ( .A(n1380), .ZN(n1327) );
XOR2_X1 U1001 ( .A(G125), .B(n1381), .Z(G27) );
NOR2_X1 U1002 ( .A1(KEYINPUT2), .A2(n1349), .ZN(n1381) );
NAND4_X1 U1003 ( .A1(n1184), .A2(n1364), .A3(n1328), .A4(n1183), .ZN(n1349) );
INV_X1 U1004 ( .A(n1150), .ZN(n1328) );
AND2_X1 U1005 ( .A1(n1154), .A2(n1359), .ZN(n1364) );
NAND2_X1 U1006 ( .A1(n1185), .A2(n1382), .ZN(n1359) );
NAND4_X1 U1007 ( .A1(G953), .A2(G902), .A3(n1383), .A4(n1216), .ZN(n1382) );
INV_X1 U1008 ( .A(G900), .ZN(n1216) );
XNOR2_X1 U1009 ( .A(G122), .B(n1331), .ZN(G24) );
NAND4_X1 U1010 ( .A1(n1335), .A2(n1173), .A3(n1384), .A4(n1385), .ZN(n1331) );
INV_X1 U1011 ( .A(n1152), .ZN(n1173) );
NAND2_X1 U1012 ( .A1(n1386), .A2(n1387), .ZN(n1152) );
XNOR2_X1 U1013 ( .A(KEYINPUT46), .B(n1339), .ZN(n1387) );
INV_X1 U1014 ( .A(n1388), .ZN(n1335) );
XOR2_X1 U1015 ( .A(G119), .B(n1389), .Z(G21) );
NOR2_X1 U1016 ( .A1(n1356), .A2(n1388), .ZN(n1389) );
NAND3_X1 U1017 ( .A1(n1154), .A2(n1326), .A3(n1184), .ZN(n1388) );
NAND3_X1 U1018 ( .A1(n1196), .A2(n1339), .A3(n1170), .ZN(n1356) );
INV_X1 U1019 ( .A(n1386), .ZN(n1196) );
XNOR2_X1 U1020 ( .A(G116), .B(n1390), .ZN(G18) );
NAND4_X1 U1021 ( .A1(n1181), .A2(n1323), .A3(n1154), .A4(n1391), .ZN(n1390) );
XOR2_X1 U1022 ( .A(KEYINPUT39), .B(n1392), .Z(n1391) );
INV_X1 U1023 ( .A(n1135), .ZN(n1323) );
NAND2_X1 U1024 ( .A1(n1366), .A2(n1384), .ZN(n1135) );
INV_X1 U1025 ( .A(n1367), .ZN(n1384) );
XOR2_X1 U1026 ( .A(n1393), .B(n1394), .Z(G15) );
XNOR2_X1 U1027 ( .A(G113), .B(KEYINPUT12), .ZN(n1394) );
NAND2_X1 U1028 ( .A1(n1334), .A2(n1325), .ZN(n1393) );
AND3_X1 U1029 ( .A1(n1183), .A2(n1326), .A3(n1181), .ZN(n1334) );
AND2_X1 U1030 ( .A1(n1171), .A2(n1184), .ZN(n1181) );
NOR2_X1 U1031 ( .A1(n1395), .A2(n1177), .ZN(n1184) );
NOR2_X1 U1032 ( .A1(n1339), .A2(n1386), .ZN(n1171) );
INV_X1 U1033 ( .A(n1169), .ZN(n1183) );
NAND2_X1 U1034 ( .A1(n1367), .A2(n1385), .ZN(n1169) );
XOR2_X1 U1035 ( .A(G110), .B(n1396), .Z(G12) );
NOR3_X1 U1036 ( .A1(n1380), .A2(n1392), .A3(n1150), .ZN(n1396) );
NAND2_X1 U1037 ( .A1(n1386), .A2(n1339), .ZN(n1150) );
NAND2_X1 U1038 ( .A1(n1205), .A2(n1397), .ZN(n1339) );
NAND2_X1 U1039 ( .A1(n1207), .A2(n1206), .ZN(n1397) );
INV_X1 U1040 ( .A(n1398), .ZN(n1206) );
INV_X1 U1041 ( .A(n1399), .ZN(n1207) );
NAND2_X1 U1042 ( .A1(n1398), .A2(n1399), .ZN(n1205) );
NAND2_X1 U1043 ( .A1(G217), .A2(n1400), .ZN(n1399) );
NOR2_X1 U1044 ( .A1(n1258), .A2(G902), .ZN(n1398) );
XNOR2_X1 U1045 ( .A(n1401), .B(n1402), .ZN(n1258) );
XOR2_X1 U1046 ( .A(G146), .B(n1403), .Z(n1402) );
NOR2_X1 U1047 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
XOR2_X1 U1048 ( .A(n1406), .B(KEYINPUT10), .Z(n1405) );
NAND3_X1 U1049 ( .A1(n1407), .A2(n1408), .A3(G221), .ZN(n1406) );
NOR2_X1 U1050 ( .A1(n1409), .A2(n1408), .ZN(n1404) );
XOR2_X1 U1051 ( .A(G137), .B(KEYINPUT54), .Z(n1408) );
AND2_X1 U1052 ( .A1(n1407), .A2(G221), .ZN(n1409) );
XOR2_X1 U1053 ( .A(n1410), .B(n1411), .Z(n1401) );
NAND2_X1 U1054 ( .A1(n1412), .A2(n1413), .ZN(n1410) );
NAND2_X1 U1055 ( .A1(n1414), .A2(n1415), .ZN(n1413) );
XOR2_X1 U1056 ( .A(KEYINPUT13), .B(n1416), .Z(n1415) );
XOR2_X1 U1057 ( .A(KEYINPUT55), .B(G110), .Z(n1414) );
XOR2_X1 U1058 ( .A(n1417), .B(KEYINPUT57), .Z(n1412) );
NAND2_X1 U1059 ( .A1(n1418), .A2(n1416), .ZN(n1417) );
XOR2_X1 U1060 ( .A(G119), .B(G128), .Z(n1416) );
XOR2_X1 U1061 ( .A(KEYINPUT55), .B(n1419), .Z(n1418) );
XOR2_X1 U1062 ( .A(n1420), .B(G472), .Z(n1386) );
NAND2_X1 U1063 ( .A1(n1421), .A2(n1314), .ZN(n1420) );
XOR2_X1 U1064 ( .A(n1422), .B(n1423), .Z(n1421) );
XOR2_X1 U1065 ( .A(n1424), .B(n1248), .Z(n1423) );
INV_X1 U1066 ( .A(n1240), .ZN(n1248) );
NOR3_X1 U1067 ( .A1(n1285), .A2(KEYINPUT37), .A3(n1284), .ZN(n1424) );
NOR2_X1 U1068 ( .A1(n1425), .A2(n1379), .ZN(n1284) );
AND2_X1 U1069 ( .A1(n1425), .A2(n1379), .ZN(n1285) );
NAND3_X1 U1070 ( .A1(n1426), .A2(n1214), .A3(G210), .ZN(n1425) );
XOR2_X1 U1071 ( .A(n1427), .B(KEYINPUT44), .Z(n1422) );
NAND3_X1 U1072 ( .A1(n1428), .A2(n1429), .A3(n1430), .ZN(n1427) );
OR2_X1 U1073 ( .A1(n1296), .A2(KEYINPUT22), .ZN(n1430) );
NAND3_X1 U1074 ( .A1(KEYINPUT22), .A2(n1296), .A3(n1281), .ZN(n1429) );
NAND2_X1 U1075 ( .A1(n1431), .A2(n1432), .ZN(n1428) );
NAND2_X1 U1076 ( .A1(KEYINPUT22), .A2(n1433), .ZN(n1432) );
XOR2_X1 U1077 ( .A(n1279), .B(KEYINPUT36), .Z(n1433) );
INV_X1 U1078 ( .A(n1326), .ZN(n1392) );
NAND2_X1 U1079 ( .A1(n1434), .A2(n1185), .ZN(n1326) );
NAND3_X1 U1080 ( .A1(n1383), .A2(n1214), .A3(G952), .ZN(n1185) );
NAND4_X1 U1081 ( .A1(G953), .A2(G902), .A3(n1383), .A4(n1435), .ZN(n1434) );
INV_X1 U1082 ( .A(G898), .ZN(n1435) );
NAND2_X1 U1083 ( .A1(G234), .A2(G237), .ZN(n1383) );
NAND3_X1 U1084 ( .A1(n1325), .A2(n1324), .A3(n1170), .ZN(n1380) );
INV_X1 U1085 ( .A(n1146), .ZN(n1170) );
NAND2_X1 U1086 ( .A1(n1367), .A2(n1366), .ZN(n1146) );
INV_X1 U1087 ( .A(n1385), .ZN(n1366) );
NAND2_X1 U1088 ( .A1(n1436), .A2(n1195), .ZN(n1385) );
NAND2_X1 U1089 ( .A1(G475), .A2(n1437), .ZN(n1195) );
XOR2_X1 U1090 ( .A(KEYINPUT47), .B(n1193), .Z(n1436) );
NOR2_X1 U1091 ( .A1(n1437), .A2(G475), .ZN(n1193) );
NAND2_X1 U1092 ( .A1(n1268), .A2(n1314), .ZN(n1437) );
XNOR2_X1 U1093 ( .A(n1438), .B(n1439), .ZN(n1268) );
XOR2_X1 U1094 ( .A(n1440), .B(n1441), .Z(n1439) );
XOR2_X1 U1095 ( .A(G122), .B(G113), .Z(n1441) );
XOR2_X1 U1096 ( .A(KEYINPUT43), .B(G131), .Z(n1440) );
XOR2_X1 U1097 ( .A(n1442), .B(n1443), .Z(n1438) );
XOR2_X1 U1098 ( .A(n1444), .B(n1445), .Z(n1443) );
NAND3_X1 U1099 ( .A1(G214), .A2(n1214), .A3(n1446), .ZN(n1445) );
XOR2_X1 U1100 ( .A(n1426), .B(KEYINPUT48), .Z(n1446) );
XOR2_X1 U1101 ( .A(n1447), .B(n1411), .Z(n1442) );
XOR2_X1 U1102 ( .A(n1224), .B(KEYINPUT25), .Z(n1411) );
XOR2_X1 U1103 ( .A(n1370), .B(n1311), .Z(n1224) );
INV_X1 U1104 ( .A(G125), .ZN(n1311) );
XOR2_X1 U1105 ( .A(n1448), .B(n1449), .Z(n1367) );
XOR2_X1 U1106 ( .A(KEYINPUT11), .B(n1200), .Z(n1449) );
NOR2_X1 U1107 ( .A1(n1263), .A2(G902), .ZN(n1200) );
XOR2_X1 U1108 ( .A(n1450), .B(n1451), .Z(n1263) );
XOR2_X1 U1109 ( .A(G128), .B(n1452), .Z(n1451) );
XOR2_X1 U1110 ( .A(G143), .B(G134), .Z(n1452) );
XOR2_X1 U1111 ( .A(n1453), .B(n1454), .Z(n1450) );
AND2_X1 U1112 ( .A1(n1407), .A2(G217), .ZN(n1454) );
AND2_X1 U1113 ( .A1(G234), .A2(n1214), .ZN(n1407) );
INV_X1 U1114 ( .A(G953), .ZN(n1214) );
NAND3_X1 U1115 ( .A1(n1455), .A2(n1456), .A3(n1457), .ZN(n1453) );
NAND2_X1 U1116 ( .A1(G107), .A2(n1458), .ZN(n1457) );
NAND2_X1 U1117 ( .A1(KEYINPUT58), .A2(n1459), .ZN(n1456) );
NAND2_X1 U1118 ( .A1(n1460), .A2(n1461), .ZN(n1459) );
XOR2_X1 U1119 ( .A(KEYINPUT18), .B(n1458), .Z(n1460) );
NAND2_X1 U1120 ( .A1(n1462), .A2(n1463), .ZN(n1455) );
INV_X1 U1121 ( .A(KEYINPUT58), .ZN(n1463) );
NAND2_X1 U1122 ( .A1(n1464), .A2(n1465), .ZN(n1462) );
NAND2_X1 U1123 ( .A1(n1458), .A2(n1466), .ZN(n1465) );
OR3_X1 U1124 ( .A1(n1458), .A2(G107), .A3(n1466), .ZN(n1464) );
INV_X1 U1125 ( .A(KEYINPUT18), .ZN(n1466) );
XOR2_X1 U1126 ( .A(G116), .B(G122), .Z(n1458) );
NAND2_X1 U1127 ( .A1(KEYINPUT3), .A2(n1265), .ZN(n1448) );
INV_X1 U1128 ( .A(G478), .ZN(n1265) );
NOR2_X1 U1129 ( .A1(n1177), .A2(n1178), .ZN(n1324) );
INV_X1 U1130 ( .A(n1395), .ZN(n1178) );
NAND2_X1 U1131 ( .A1(n1208), .A2(n1194), .ZN(n1395) );
NAND2_X1 U1132 ( .A1(G469), .A2(n1467), .ZN(n1194) );
OR2_X1 U1133 ( .A1(n1467), .A2(G469), .ZN(n1208) );
NAND2_X1 U1134 ( .A1(n1468), .A2(n1314), .ZN(n1467) );
XOR2_X1 U1135 ( .A(n1469), .B(n1470), .Z(n1468) );
XOR2_X1 U1136 ( .A(n1471), .B(n1296), .Z(n1470) );
INV_X1 U1137 ( .A(n1279), .ZN(n1296) );
XOR2_X1 U1138 ( .A(n1225), .B(n1472), .Z(n1279) );
NOR2_X1 U1139 ( .A1(n1473), .A2(n1474), .ZN(n1472) );
AND3_X1 U1140 ( .A1(KEYINPUT15), .A2(n1475), .A3(G134), .ZN(n1474) );
INV_X1 U1141 ( .A(G137), .ZN(n1475) );
NOR2_X1 U1142 ( .A1(KEYINPUT15), .A2(n1221), .ZN(n1473) );
XOR2_X1 U1143 ( .A(G134), .B(G137), .Z(n1221) );
INV_X1 U1144 ( .A(G131), .ZN(n1225) );
NOR2_X1 U1145 ( .A1(KEYINPUT23), .A2(n1222), .ZN(n1471) );
XOR2_X1 U1146 ( .A(n1476), .B(n1477), .Z(n1222) );
INV_X1 U1147 ( .A(n1447), .ZN(n1477) );
XOR2_X1 U1148 ( .A(n1361), .B(G146), .Z(n1447) );
XNOR2_X1 U1149 ( .A(G128), .B(KEYINPUT61), .ZN(n1476) );
XOR2_X1 U1150 ( .A(n1298), .B(n1478), .Z(n1469) );
NOR2_X1 U1151 ( .A1(n1479), .A2(n1480), .ZN(n1478) );
NOR2_X1 U1152 ( .A1(n1481), .A2(n1290), .ZN(n1480) );
INV_X1 U1153 ( .A(n1482), .ZN(n1290) );
NOR2_X1 U1154 ( .A1(G953), .A2(n1215), .ZN(n1481) );
NOR3_X1 U1155 ( .A1(n1483), .A2(G953), .A3(n1215), .ZN(n1479) );
INV_X1 U1156 ( .A(G227), .ZN(n1215) );
XOR2_X1 U1157 ( .A(KEYINPUT56), .B(n1482), .Z(n1483) );
XNOR2_X1 U1158 ( .A(n1370), .B(G110), .ZN(n1482) );
INV_X1 U1159 ( .A(G140), .ZN(n1370) );
NAND3_X1 U1160 ( .A1(n1484), .A2(n1485), .A3(n1486), .ZN(n1298) );
OR2_X1 U1161 ( .A1(n1487), .A2(KEYINPUT26), .ZN(n1486) );
NAND3_X1 U1162 ( .A1(KEYINPUT26), .A2(n1487), .A3(G101), .ZN(n1485) );
NAND2_X1 U1163 ( .A1(n1488), .A2(n1379), .ZN(n1484) );
INV_X1 U1164 ( .A(G101), .ZN(n1379) );
NAND2_X1 U1165 ( .A1(n1489), .A2(KEYINPUT26), .ZN(n1488) );
XNOR2_X1 U1166 ( .A(n1487), .B(KEYINPUT1), .ZN(n1489) );
XNOR2_X1 U1167 ( .A(n1461), .B(n1490), .ZN(n1487) );
NOR2_X1 U1168 ( .A1(KEYINPUT4), .A2(n1444), .ZN(n1490) );
INV_X1 U1169 ( .A(G104), .ZN(n1444) );
INV_X1 U1170 ( .A(G107), .ZN(n1461) );
AND2_X1 U1171 ( .A1(G221), .A2(n1400), .ZN(n1177) );
NAND2_X1 U1172 ( .A1(G234), .A2(n1314), .ZN(n1400) );
XNOR2_X1 U1173 ( .A(n1154), .B(KEYINPUT28), .ZN(n1325) );
NOR2_X1 U1174 ( .A1(n1192), .A2(n1188), .ZN(n1154) );
AND3_X1 U1175 ( .A1(n1491), .A2(n1492), .A3(n1493), .ZN(n1188) );
NAND3_X1 U1176 ( .A1(G210), .A2(G237), .A3(n1494), .ZN(n1493) );
NAND3_X1 U1177 ( .A1(n1495), .A2(n1496), .A3(n1314), .ZN(n1492) );
NAND2_X1 U1178 ( .A1(G210), .A2(G237), .ZN(n1496) );
INV_X1 U1179 ( .A(n1494), .ZN(n1495) );
XOR2_X1 U1180 ( .A(n1497), .B(n1498), .Z(n1494) );
XOR2_X1 U1181 ( .A(G125), .B(n1313), .Z(n1498) );
NOR2_X1 U1182 ( .A1(n1231), .A2(G953), .ZN(n1313) );
INV_X1 U1183 ( .A(G224), .ZN(n1231) );
XOR2_X1 U1184 ( .A(n1304), .B(n1281), .Z(n1497) );
INV_X1 U1185 ( .A(n1431), .ZN(n1281) );
XOR2_X1 U1186 ( .A(n1499), .B(n1500), .Z(n1431) );
NOR2_X1 U1187 ( .A1(KEYINPUT19), .A2(n1361), .ZN(n1500) );
INV_X1 U1188 ( .A(G143), .ZN(n1361) );
XNOR2_X1 U1189 ( .A(G128), .B(G146), .ZN(n1499) );
XOR2_X1 U1190 ( .A(n1247), .B(n1244), .Z(n1304) );
INV_X1 U1191 ( .A(n1246), .ZN(n1244) );
XOR2_X1 U1192 ( .A(n1419), .B(G122), .Z(n1246) );
INV_X1 U1193 ( .A(G110), .ZN(n1419) );
XOR2_X1 U1194 ( .A(n1240), .B(n1249), .Z(n1247) );
XOR2_X1 U1195 ( .A(G101), .B(n1501), .Z(n1249) );
XOR2_X1 U1196 ( .A(G107), .B(G104), .Z(n1501) );
XNOR2_X1 U1197 ( .A(G113), .B(n1502), .ZN(n1240) );
XOR2_X1 U1198 ( .A(G119), .B(G116), .Z(n1502) );
NAND2_X1 U1199 ( .A1(G210), .A2(G902), .ZN(n1491) );
INV_X1 U1200 ( .A(n1156), .ZN(n1192) );
NAND2_X1 U1201 ( .A1(G214), .A2(n1503), .ZN(n1156) );
NAND2_X1 U1202 ( .A1(n1426), .A2(n1314), .ZN(n1503) );
INV_X1 U1203 ( .A(G902), .ZN(n1314) );
INV_X1 U1204 ( .A(G237), .ZN(n1426) );
endmodule


