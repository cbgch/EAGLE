//Key = 1011101100111110100101011101101000100010111111000011111010000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;

XNOR2_X1 U733 ( .A(G107), .B(n1006), .ZN(G9) );
NAND3_X1 U734 ( .A1(n1007), .A2(n1008), .A3(KEYINPUT52), .ZN(n1006) );
NOR2_X1 U735 ( .A1(n1009), .A2(n1010), .ZN(G75) );
XOR2_X1 U736 ( .A(KEYINPUT32), .B(n1011), .Z(n1010) );
NOR3_X1 U737 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
NOR2_X1 U738 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U739 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U740 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U741 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U742 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U743 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U744 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U745 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U746 ( .A1(n1031), .A2(n1032), .ZN(n1025) );
NOR2_X1 U747 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U749 ( .A1(n1028), .A2(n1037), .A3(n1032), .ZN(n1021) );
NOR2_X1 U750 ( .A1(n1007), .A2(n1038), .ZN(n1037) );
NOR4_X1 U751 ( .A1(n1039), .A2(n1032), .A3(n1028), .A4(n1024), .ZN(n1017) );
INV_X1 U752 ( .A(n1040), .ZN(n1024) );
NOR2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
XNOR2_X1 U754 ( .A(n1043), .B(KEYINPUT21), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1041) );
NOR2_X1 U756 ( .A1(G952), .A2(n1014), .ZN(n1009) );
NAND2_X1 U757 ( .A1(n1046), .A2(n1047), .ZN(n1014) );
NAND4_X1 U758 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
NOR4_X1 U759 ( .A1(n1028), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1051) );
XNOR2_X1 U760 ( .A(KEYINPUT26), .B(n1055), .ZN(n1054) );
XOR2_X1 U761 ( .A(n1056), .B(n1057), .Z(n1053) );
NAND2_X1 U762 ( .A1(KEYINPUT40), .A2(n1058), .ZN(n1057) );
XOR2_X1 U763 ( .A(n1059), .B(n1060), .Z(n1052) );
XOR2_X1 U764 ( .A(KEYINPUT30), .B(G472), .Z(n1060) );
NOR2_X1 U765 ( .A1(n1061), .A2(KEYINPUT15), .ZN(n1059) );
NOR3_X1 U766 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1050) );
NOR2_X1 U767 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
XOR2_X1 U768 ( .A(KEYINPUT61), .B(G478), .Z(n1066) );
XOR2_X1 U769 ( .A(n1067), .B(n1068), .Z(G72) );
XOR2_X1 U770 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR3_X1 U771 ( .A1(n1071), .A2(KEYINPUT5), .A3(G953), .ZN(n1070) );
AND2_X1 U772 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
XOR2_X1 U774 ( .A(n1076), .B(n1077), .Z(n1075) );
NOR2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U776 ( .A(n1080), .B(KEYINPUT6), .Z(n1079) );
NAND2_X1 U777 ( .A1(G125), .A2(n1081), .ZN(n1080) );
NOR2_X1 U778 ( .A1(G125), .A2(n1081), .ZN(n1078) );
NOR2_X1 U779 ( .A1(KEYINPUT22), .A2(n1082), .ZN(n1076) );
XOR2_X1 U780 ( .A(n1083), .B(n1084), .Z(n1082) );
XNOR2_X1 U781 ( .A(n1085), .B(n1086), .ZN(n1084) );
NOR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U783 ( .A(KEYINPUT46), .B(n1089), .Z(n1088) );
NOR2_X1 U784 ( .A1(G134), .A2(n1090), .ZN(n1089) );
XNOR2_X1 U785 ( .A(G131), .B(KEYINPUT19), .ZN(n1083) );
NOR2_X1 U786 ( .A1(n1091), .A2(n1092), .ZN(n1074) );
XNOR2_X1 U787 ( .A(G900), .B(KEYINPUT24), .ZN(n1091) );
NOR2_X1 U788 ( .A1(n1093), .A2(n1046), .ZN(n1067) );
AND2_X1 U789 ( .A1(G227), .A2(G900), .ZN(n1093) );
XOR2_X1 U790 ( .A(n1094), .B(n1095), .Z(G69) );
NOR2_X1 U791 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U792 ( .A1(n1098), .A2(n1046), .ZN(n1097) );
NOR2_X1 U793 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U794 ( .A(KEYINPUT7), .B(n1101), .ZN(n1100) );
NOR2_X1 U795 ( .A1(G953), .A2(n1102), .ZN(n1096) );
NAND3_X1 U796 ( .A1(n1103), .A2(n1104), .A3(KEYINPUT50), .ZN(n1094) );
NAND2_X1 U797 ( .A1(n1105), .A2(n1101), .ZN(n1104) );
XNOR2_X1 U798 ( .A(n1106), .B(n1107), .ZN(n1103) );
NAND2_X1 U799 ( .A1(KEYINPUT10), .A2(n1108), .ZN(n1106) );
NOR2_X1 U800 ( .A1(n1109), .A2(n1110), .ZN(G66) );
NOR3_X1 U801 ( .A1(n1058), .A2(n1111), .A3(n1112), .ZN(n1110) );
NOR3_X1 U802 ( .A1(n1113), .A2(n1056), .A3(n1114), .ZN(n1112) );
INV_X1 U803 ( .A(n1115), .ZN(n1113) );
NOR2_X1 U804 ( .A1(n1116), .A2(n1115), .ZN(n1111) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1056), .ZN(n1116) );
NOR2_X1 U806 ( .A1(n1109), .A2(n1118), .ZN(G63) );
NOR2_X1 U807 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U808 ( .A(n1121), .B(KEYINPUT53), .Z(n1120) );
NAND2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U810 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
AND2_X1 U811 ( .A1(n1124), .A2(G478), .ZN(n1122) );
NOR3_X1 U812 ( .A1(n1109), .A2(n1125), .A3(n1126), .ZN(G60) );
NOR2_X1 U813 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U814 ( .A(KEYINPUT9), .B(n1129), .ZN(n1128) );
NOR2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1125) );
XOR2_X1 U816 ( .A(n1129), .B(KEYINPUT37), .Z(n1131) );
NAND2_X1 U817 ( .A1(n1124), .A2(G475), .ZN(n1129) );
XOR2_X1 U818 ( .A(G104), .B(n1132), .Z(G6) );
NOR2_X1 U819 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U820 ( .A1(n1109), .A2(n1135), .ZN(G57) );
XOR2_X1 U821 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U822 ( .A(n1138), .B(n1139), .Z(n1137) );
XNOR2_X1 U823 ( .A(G101), .B(KEYINPUT18), .ZN(n1139) );
XNOR2_X1 U824 ( .A(n1140), .B(n1141), .ZN(n1136) );
AND2_X1 U825 ( .A1(G472), .A2(n1124), .ZN(n1141) );
NOR2_X1 U826 ( .A1(n1109), .A2(n1142), .ZN(G54) );
XOR2_X1 U827 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U828 ( .A(n1145), .B(n1146), .ZN(n1144) );
NAND2_X1 U829 ( .A1(KEYINPUT38), .A2(n1147), .ZN(n1145) );
INV_X1 U830 ( .A(n1148), .ZN(n1147) );
XOR2_X1 U831 ( .A(n1149), .B(n1150), .Z(n1143) );
NOR2_X1 U832 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U833 ( .A(n1153), .B(KEYINPUT12), .Z(n1152) );
NAND2_X1 U834 ( .A1(G110), .A2(n1081), .ZN(n1153) );
NAND3_X1 U835 ( .A1(n1154), .A2(n1012), .A3(G469), .ZN(n1149) );
XNOR2_X1 U836 ( .A(KEYINPUT8), .B(n1155), .ZN(n1154) );
NOR2_X1 U837 ( .A1(n1109), .A2(n1156), .ZN(G51) );
XOR2_X1 U838 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U839 ( .A1(KEYINPUT36), .A2(n1159), .ZN(n1158) );
NOR2_X1 U840 ( .A1(n1160), .A2(n1114), .ZN(n1157) );
INV_X1 U841 ( .A(n1124), .ZN(n1114) );
NOR2_X1 U842 ( .A1(n1155), .A2(n1117), .ZN(n1124) );
INV_X1 U843 ( .A(n1012), .ZN(n1117) );
NAND3_X1 U844 ( .A1(n1102), .A2(n1161), .A3(n1073), .ZN(n1012) );
AND4_X1 U845 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1073) );
AND3_X1 U846 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
NAND3_X1 U847 ( .A1(n1169), .A2(n1170), .A3(n1043), .ZN(n1164) );
NAND2_X1 U848 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
NAND4_X1 U849 ( .A1(n1029), .A2(n1034), .A3(n1173), .A4(n1174), .ZN(n1172) );
NAND3_X1 U850 ( .A1(n1038), .A2(n1175), .A3(n1030), .ZN(n1171) );
XNOR2_X1 U851 ( .A(KEYINPUT16), .B(n1072), .ZN(n1161) );
AND2_X1 U852 ( .A1(n1176), .A2(n1177), .ZN(n1102) );
AND4_X1 U853 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR4_X1 U854 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1176) );
AND2_X1 U855 ( .A1(n1008), .A2(n1007), .ZN(n1185) );
INV_X1 U856 ( .A(n1133), .ZN(n1008) );
NAND2_X1 U857 ( .A1(n1186), .A2(n1187), .ZN(n1133) );
NOR4_X1 U858 ( .A1(n1188), .A2(n1189), .A3(n1032), .A4(n1134), .ZN(n1184) );
INV_X1 U859 ( .A(n1187), .ZN(n1032) );
NOR2_X1 U860 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
INV_X1 U861 ( .A(KEYINPUT29), .ZN(n1191) );
NOR3_X1 U862 ( .A1(n1192), .A2(n1193), .A3(n1043), .ZN(n1190) );
NOR2_X1 U863 ( .A1(KEYINPUT29), .A2(n1186), .ZN(n1188) );
INV_X1 U864 ( .A(n1194), .ZN(n1182) );
NOR2_X1 U865 ( .A1(n1046), .A2(G952), .ZN(n1109) );
XOR2_X1 U866 ( .A(n1162), .B(n1195), .Z(G48) );
NAND2_X1 U867 ( .A1(KEYINPUT28), .A2(n1196), .ZN(n1195) );
XOR2_X1 U868 ( .A(KEYINPUT57), .B(G146), .Z(n1196) );
NAND3_X1 U869 ( .A1(n1197), .A2(n1043), .A3(n1038), .ZN(n1162) );
XNOR2_X1 U870 ( .A(G143), .B(n1198), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1029), .A2(n1043), .A3(n1199), .A4(n1200), .ZN(n1198) );
NOR4_X1 U872 ( .A1(KEYINPUT33), .A2(n1201), .A3(n1202), .A4(n1048), .ZN(n1200) );
XNOR2_X1 U873 ( .A(n1034), .B(KEYINPUT23), .ZN(n1199) );
XNOR2_X1 U874 ( .A(G140), .B(n1072), .ZN(G42) );
NAND3_X1 U875 ( .A1(n1038), .A2(n1203), .A3(n1030), .ZN(n1072) );
XNOR2_X1 U876 ( .A(G137), .B(n1167), .ZN(G39) );
NAND3_X1 U877 ( .A1(n1204), .A2(n1197), .A3(n1040), .ZN(n1167) );
XNOR2_X1 U878 ( .A(n1205), .B(n1206), .ZN(G36) );
NAND2_X1 U879 ( .A1(KEYINPUT63), .A2(n1168), .ZN(n1205) );
NAND3_X1 U880 ( .A1(n1203), .A2(n1007), .A3(n1029), .ZN(n1168) );
NAND2_X1 U881 ( .A1(n1207), .A2(n1208), .ZN(G33) );
NAND2_X1 U882 ( .A1(G131), .A2(n1163), .ZN(n1208) );
XOR2_X1 U883 ( .A(n1209), .B(KEYINPUT39), .Z(n1207) );
OR2_X1 U884 ( .A1(n1163), .A2(G131), .ZN(n1209) );
NAND3_X1 U885 ( .A1(n1029), .A2(n1203), .A3(n1038), .ZN(n1163) );
NOR3_X1 U886 ( .A1(n1192), .A2(n1202), .A3(n1020), .ZN(n1203) );
INV_X1 U887 ( .A(n1204), .ZN(n1020) );
NOR2_X1 U888 ( .A1(n1044), .A2(n1064), .ZN(n1204) );
INV_X1 U889 ( .A(n1045), .ZN(n1064) );
XNOR2_X1 U890 ( .A(n1210), .B(KEYINPUT2), .ZN(n1044) );
INV_X1 U891 ( .A(n1170), .ZN(n1202) );
NAND2_X1 U892 ( .A1(n1211), .A2(n1212), .ZN(G30) );
NAND2_X1 U893 ( .A1(G128), .A2(n1166), .ZN(n1212) );
XOR2_X1 U894 ( .A(KEYINPUT27), .B(n1213), .Z(n1211) );
NOR2_X1 U895 ( .A1(G128), .A2(n1166), .ZN(n1213) );
NAND3_X1 U896 ( .A1(n1007), .A2(n1043), .A3(n1197), .ZN(n1166) );
AND4_X1 U897 ( .A1(n1034), .A2(n1170), .A3(n1214), .A4(n1215), .ZN(n1197) );
OR2_X1 U898 ( .A1(n1029), .A2(KEYINPUT11), .ZN(n1215) );
NAND2_X1 U899 ( .A1(KEYINPUT11), .A2(n1216), .ZN(n1214) );
NAND2_X1 U900 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
INV_X1 U901 ( .A(n1192), .ZN(n1034) );
INV_X1 U902 ( .A(n1219), .ZN(n1043) );
XNOR2_X1 U903 ( .A(G101), .B(n1179), .ZN(G3) );
NAND3_X1 U904 ( .A1(n1040), .A2(n1186), .A3(n1029), .ZN(n1179) );
XOR2_X1 U905 ( .A(G125), .B(n1220), .Z(G27) );
NOR2_X1 U906 ( .A1(n1221), .A2(n1219), .ZN(n1220) );
XOR2_X1 U907 ( .A(n1222), .B(KEYINPUT31), .Z(n1221) );
NAND4_X1 U908 ( .A1(n1030), .A2(n1175), .A3(n1223), .A4(n1170), .ZN(n1222) );
NAND2_X1 U909 ( .A1(n1016), .A2(n1224), .ZN(n1170) );
NAND2_X1 U910 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U911 ( .A(KEYINPUT24), .B(G900), .Z(n1226) );
XNOR2_X1 U912 ( .A(KEYINPUT48), .B(n1134), .ZN(n1223) );
INV_X1 U913 ( .A(n1038), .ZN(n1134) );
INV_X1 U914 ( .A(n1028), .ZN(n1175) );
XNOR2_X1 U915 ( .A(G122), .B(n1178), .ZN(G24) );
NAND4_X1 U916 ( .A1(n1227), .A2(n1187), .A3(n1173), .A4(n1174), .ZN(n1178) );
NOR2_X1 U917 ( .A1(n1218), .A2(n1217), .ZN(n1187) );
XOR2_X1 U918 ( .A(G119), .B(n1183), .Z(G21) );
AND4_X1 U919 ( .A1(n1227), .A2(n1040), .A3(n1228), .A4(n1218), .ZN(n1183) );
XNOR2_X1 U920 ( .A(KEYINPUT11), .B(n1217), .ZN(n1228) );
INV_X1 U921 ( .A(n1229), .ZN(n1217) );
NAND2_X1 U922 ( .A1(n1230), .A2(n1231), .ZN(G18) );
NAND2_X1 U923 ( .A1(G116), .A2(n1194), .ZN(n1231) );
XOR2_X1 U924 ( .A(n1232), .B(KEYINPUT1), .Z(n1230) );
OR2_X1 U925 ( .A1(n1194), .A2(G116), .ZN(n1232) );
NAND3_X1 U926 ( .A1(n1029), .A2(n1007), .A3(n1227), .ZN(n1194) );
NOR2_X1 U927 ( .A1(n1173), .A2(n1201), .ZN(n1007) );
XNOR2_X1 U928 ( .A(G113), .B(n1181), .ZN(G15) );
NAND3_X1 U929 ( .A1(n1038), .A2(n1029), .A3(n1227), .ZN(n1181) );
NOR3_X1 U930 ( .A1(n1219), .A2(n1193), .A3(n1028), .ZN(n1227) );
NAND2_X1 U931 ( .A1(n1233), .A2(n1036), .ZN(n1028) );
INV_X1 U932 ( .A(n1035), .ZN(n1233) );
AND2_X1 U933 ( .A1(n1229), .A2(n1218), .ZN(n1029) );
NOR2_X1 U934 ( .A1(n1174), .A2(n1048), .ZN(n1038) );
INV_X1 U935 ( .A(n1173), .ZN(n1048) );
XNOR2_X1 U936 ( .A(G110), .B(n1180), .ZN(G12) );
NAND3_X1 U937 ( .A1(n1040), .A2(n1186), .A3(n1030), .ZN(n1180) );
NOR2_X1 U938 ( .A1(n1229), .A2(n1218), .ZN(n1030) );
XNOR2_X1 U939 ( .A(n1234), .B(n1235), .ZN(n1218) );
NOR2_X1 U940 ( .A1(KEYINPUT58), .A2(G472), .ZN(n1235) );
XNOR2_X1 U941 ( .A(n1061), .B(KEYINPUT51), .ZN(n1234) );
AND2_X1 U942 ( .A1(n1236), .A2(n1155), .ZN(n1061) );
NAND2_X1 U943 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND2_X1 U944 ( .A1(n1239), .A2(n1140), .ZN(n1238) );
XOR2_X1 U945 ( .A(KEYINPUT41), .B(n1240), .Z(n1237) );
NOR2_X1 U946 ( .A1(n1239), .A2(n1140), .ZN(n1240) );
XOR2_X1 U947 ( .A(n1241), .B(n1242), .Z(n1140) );
XOR2_X1 U948 ( .A(n1243), .B(n1244), .Z(n1242) );
NAND2_X1 U949 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
OR2_X1 U950 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
XOR2_X1 U951 ( .A(n1249), .B(KEYINPUT59), .Z(n1245) );
NAND2_X1 U952 ( .A1(n1247), .A2(n1248), .ZN(n1249) );
XOR2_X1 U953 ( .A(G113), .B(KEYINPUT49), .Z(n1247) );
XNOR2_X1 U954 ( .A(G101), .B(n1250), .ZN(n1239) );
NOR2_X1 U955 ( .A1(KEYINPUT20), .A2(n1138), .ZN(n1250) );
NAND2_X1 U956 ( .A1(G210), .A2(n1251), .ZN(n1138) );
XNOR2_X1 U957 ( .A(n1056), .B(n1252), .ZN(n1229) );
NOR2_X1 U958 ( .A1(n1058), .A2(KEYINPUT17), .ZN(n1252) );
NOR2_X1 U959 ( .A1(n1115), .A2(G902), .ZN(n1058) );
XNOR2_X1 U960 ( .A(n1253), .B(n1254), .ZN(n1115) );
XOR2_X1 U961 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U962 ( .A(n1257), .B(G119), .ZN(n1256) );
XNOR2_X1 U963 ( .A(G146), .B(n1090), .ZN(n1255) );
XNOR2_X1 U964 ( .A(n1258), .B(n1259), .ZN(n1253) );
XOR2_X1 U965 ( .A(n1260), .B(n1261), .Z(n1258) );
NOR2_X1 U966 ( .A1(KEYINPUT35), .A2(G110), .ZN(n1261) );
NAND2_X1 U967 ( .A1(G221), .A2(n1262), .ZN(n1260) );
NAND2_X1 U968 ( .A1(G217), .A2(n1263), .ZN(n1056) );
NOR3_X1 U969 ( .A1(n1219), .A2(n1193), .A3(n1192), .ZN(n1186) );
NAND2_X1 U970 ( .A1(n1035), .A2(n1036), .ZN(n1192) );
NAND2_X1 U971 ( .A1(G221), .A2(n1263), .ZN(n1036) );
NAND2_X1 U972 ( .A1(G234), .A2(n1155), .ZN(n1263) );
XNOR2_X1 U973 ( .A(n1264), .B(G469), .ZN(n1035) );
NAND4_X1 U974 ( .A1(n1265), .A2(n1155), .A3(n1266), .A4(n1267), .ZN(n1264) );
OR3_X1 U975 ( .A1(n1268), .A2(n1269), .A3(n1081), .ZN(n1267) );
NAND2_X1 U976 ( .A1(n1270), .A2(n1081), .ZN(n1266) );
XNOR2_X1 U977 ( .A(G110), .B(n1269), .ZN(n1270) );
NAND2_X1 U978 ( .A1(n1151), .A2(n1269), .ZN(n1265) );
XOR2_X1 U979 ( .A(n1271), .B(n1272), .Z(n1269) );
INV_X1 U980 ( .A(n1146), .ZN(n1272) );
XNOR2_X1 U981 ( .A(n1243), .B(n1273), .ZN(n1146) );
AND2_X1 U982 ( .A1(n1046), .A2(G227), .ZN(n1273) );
NAND3_X1 U983 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1243) );
NAND2_X1 U984 ( .A1(n1087), .A2(G131), .ZN(n1276) );
NOR2_X1 U985 ( .A1(n1206), .A2(G137), .ZN(n1087) );
NAND3_X1 U986 ( .A1(n1277), .A2(n1206), .A3(n1090), .ZN(n1275) );
INV_X1 U987 ( .A(G137), .ZN(n1090) );
INV_X1 U988 ( .A(G131), .ZN(n1277) );
NAND2_X1 U989 ( .A1(n1278), .A2(G137), .ZN(n1274) );
XNOR2_X1 U990 ( .A(n1206), .B(G131), .ZN(n1278) );
NAND2_X1 U991 ( .A1(KEYINPUT42), .A2(n1148), .ZN(n1271) );
XOR2_X1 U992 ( .A(n1279), .B(n1280), .Z(n1148) );
INV_X1 U993 ( .A(n1085), .ZN(n1280) );
XOR2_X1 U994 ( .A(n1241), .B(KEYINPUT47), .Z(n1085) );
XNOR2_X1 U995 ( .A(n1281), .B(n1282), .ZN(n1279) );
INV_X1 U996 ( .A(G101), .ZN(n1282) );
NAND2_X1 U997 ( .A1(n1283), .A2(KEYINPUT43), .ZN(n1281) );
XOR2_X1 U998 ( .A(n1284), .B(G107), .Z(n1283) );
NAND2_X1 U999 ( .A1(KEYINPUT54), .A2(n1285), .ZN(n1284) );
NOR2_X1 U1000 ( .A1(n1081), .A2(G110), .ZN(n1151) );
AND2_X1 U1001 ( .A1(n1286), .A2(n1287), .ZN(n1193) );
NAND2_X1 U1002 ( .A1(n1225), .A2(n1101), .ZN(n1287) );
INV_X1 U1003 ( .A(G898), .ZN(n1101) );
AND3_X1 U1004 ( .A1(n1105), .A2(n1288), .A3(G902), .ZN(n1225) );
INV_X1 U1005 ( .A(n1092), .ZN(n1105) );
XOR2_X1 U1006 ( .A(G953), .B(KEYINPUT44), .Z(n1092) );
XNOR2_X1 U1007 ( .A(KEYINPUT34), .B(n1016), .ZN(n1286) );
NAND3_X1 U1008 ( .A1(n1288), .A2(n1046), .A3(G952), .ZN(n1016) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1288) );
NAND2_X1 U1010 ( .A1(n1210), .A2(n1045), .ZN(n1219) );
NAND2_X1 U1011 ( .A1(G214), .A2(n1289), .ZN(n1045) );
NAND2_X1 U1012 ( .A1(n1055), .A2(n1049), .ZN(n1210) );
NAND2_X1 U1013 ( .A1(n1290), .A2(n1291), .ZN(n1049) );
OR2_X1 U1014 ( .A1(n1291), .A2(n1290), .ZN(n1055) );
INV_X1 U1015 ( .A(n1160), .ZN(n1290) );
NAND2_X1 U1016 ( .A1(G210), .A2(n1289), .ZN(n1160) );
NAND2_X1 U1017 ( .A1(n1292), .A2(n1155), .ZN(n1289) );
INV_X1 U1018 ( .A(G237), .ZN(n1292) );
NAND2_X1 U1019 ( .A1(n1159), .A2(n1155), .ZN(n1291) );
XNOR2_X1 U1020 ( .A(n1293), .B(n1294), .ZN(n1159) );
XOR2_X1 U1021 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1022 ( .A(G125), .B(n1297), .ZN(n1296) );
NOR2_X1 U1023 ( .A1(G953), .A2(n1099), .ZN(n1297) );
INV_X1 U1024 ( .A(G224), .ZN(n1099) );
NAND2_X1 U1025 ( .A1(KEYINPUT14), .A2(n1107), .ZN(n1295) );
XNOR2_X1 U1026 ( .A(G122), .B(n1268), .ZN(n1107) );
INV_X1 U1027 ( .A(G110), .ZN(n1268) );
XNOR2_X1 U1028 ( .A(n1108), .B(n1298), .ZN(n1293) );
INV_X1 U1029 ( .A(n1241), .ZN(n1298) );
XOR2_X1 U1030 ( .A(G128), .B(n1299), .Z(n1241) );
XOR2_X1 U1031 ( .A(n1300), .B(n1301), .Z(n1108) );
XNOR2_X1 U1032 ( .A(n1302), .B(n1285), .ZN(n1301) );
NAND2_X1 U1033 ( .A1(n1303), .A2(KEYINPUT3), .ZN(n1302) );
XNOR2_X1 U1034 ( .A(G101), .B(KEYINPUT60), .ZN(n1303) );
XOR2_X1 U1035 ( .A(n1304), .B(G107), .Z(n1300) );
NAND2_X1 U1036 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U1037 ( .A1(G113), .A2(n1248), .ZN(n1306) );
XOR2_X1 U1038 ( .A(KEYINPUT45), .B(n1307), .Z(n1305) );
NOR2_X1 U1039 ( .A1(G113), .A2(n1248), .ZN(n1307) );
XOR2_X1 U1040 ( .A(G119), .B(G116), .Z(n1248) );
NOR2_X1 U1041 ( .A1(n1174), .A2(n1173), .ZN(n1040) );
XNOR2_X1 U1042 ( .A(n1308), .B(G475), .ZN(n1173) );
NAND2_X1 U1043 ( .A1(n1127), .A2(n1155), .ZN(n1308) );
INV_X1 U1044 ( .A(G902), .ZN(n1155) );
INV_X1 U1045 ( .A(n1130), .ZN(n1127) );
XNOR2_X1 U1046 ( .A(n1309), .B(n1310), .ZN(n1130) );
XNOR2_X1 U1047 ( .A(n1311), .B(n1299), .ZN(n1310) );
XOR2_X1 U1048 ( .A(G143), .B(G146), .Z(n1299) );
NAND2_X1 U1049 ( .A1(KEYINPUT13), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1050 ( .A(n1313), .B(n1314), .ZN(n1312) );
XOR2_X1 U1051 ( .A(G122), .B(G113), .Z(n1314) );
INV_X1 U1052 ( .A(n1285), .ZN(n1313) );
XOR2_X1 U1053 ( .A(G104), .B(KEYINPUT25), .Z(n1285) );
NAND2_X1 U1054 ( .A1(n1315), .A2(n1316), .ZN(n1309) );
NAND2_X1 U1055 ( .A1(n1317), .A2(n1259), .ZN(n1316) );
XOR2_X1 U1056 ( .A(KEYINPUT4), .B(n1318), .Z(n1317) );
NAND2_X1 U1057 ( .A1(n1319), .A2(n1320), .ZN(n1315) );
INV_X1 U1058 ( .A(n1259), .ZN(n1320) );
XOR2_X1 U1059 ( .A(G125), .B(n1081), .Z(n1259) );
INV_X1 U1060 ( .A(G140), .ZN(n1081) );
XOR2_X1 U1061 ( .A(KEYINPUT55), .B(n1318), .Z(n1319) );
XNOR2_X1 U1062 ( .A(n1321), .B(G131), .ZN(n1318) );
NAND2_X1 U1063 ( .A1(G214), .A2(n1251), .ZN(n1321) );
NOR2_X1 U1064 ( .A1(G953), .A2(G237), .ZN(n1251) );
INV_X1 U1065 ( .A(n1201), .ZN(n1174) );
NOR2_X1 U1066 ( .A1(n1322), .A2(n1063), .ZN(n1201) );
NOR2_X1 U1067 ( .A1(n1323), .A2(G478), .ZN(n1063) );
AND2_X1 U1068 ( .A1(n1324), .A2(n1323), .ZN(n1322) );
INV_X1 U1069 ( .A(n1065), .ZN(n1323) );
NOR2_X1 U1070 ( .A1(n1123), .A2(G902), .ZN(n1065) );
XOR2_X1 U1071 ( .A(n1325), .B(n1326), .Z(n1123) );
XOR2_X1 U1072 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1073 ( .A(G116), .B(G107), .Z(n1328) );
XNOR2_X1 U1074 ( .A(n1329), .B(G122), .ZN(n1327) );
INV_X1 U1075 ( .A(G143), .ZN(n1329) );
XOR2_X1 U1076 ( .A(n1330), .B(n1331), .Z(n1325) );
AND2_X1 U1077 ( .A1(n1262), .A2(G217), .ZN(n1331) );
AND2_X1 U1078 ( .A1(G234), .A2(n1046), .ZN(n1262) );
INV_X1 U1079 ( .A(G953), .ZN(n1046) );
XNOR2_X1 U1080 ( .A(n1332), .B(n1333), .ZN(n1330) );
NAND2_X1 U1081 ( .A1(KEYINPUT0), .A2(n1206), .ZN(n1333) );
INV_X1 U1082 ( .A(G134), .ZN(n1206) );
NAND2_X1 U1083 ( .A1(KEYINPUT56), .A2(n1257), .ZN(n1332) );
INV_X1 U1084 ( .A(G128), .ZN(n1257) );
XOR2_X1 U1085 ( .A(KEYINPUT62), .B(G478), .Z(n1324) );
endmodule


