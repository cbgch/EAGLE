//Key = 0010010001011010110101101001011100101100100010110111001111100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;

XOR2_X1 U739 ( .A(n1010), .B(G107), .Z(G9) );
NAND2_X1 U740 ( .A1(KEYINPUT34), .A2(n1011), .ZN(n1010) );
NOR2_X1 U741 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
INV_X1 U743 ( .A(G952), .ZN(n1017) );
XOR2_X1 U744 ( .A(n1018), .B(KEYINPUT28), .Z(n1016) );
NAND2_X1 U745 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND3_X1 U746 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NAND2_X1 U747 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NAND3_X1 U748 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NAND2_X1 U749 ( .A1(n1029), .A2(n1030), .ZN(n1024) );
NAND2_X1 U750 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND3_X1 U751 ( .A1(n1033), .A2(n1027), .A3(n1034), .ZN(n1032) );
NAND2_X1 U752 ( .A1(n1026), .A2(n1035), .ZN(n1031) );
XOR2_X1 U753 ( .A(KEYINPUT45), .B(n1036), .Z(n1035) );
NOR2_X1 U754 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U755 ( .A1(n1039), .A2(n1040), .ZN(n1019) );
NAND4_X1 U756 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1014) );
NAND3_X1 U757 ( .A1(n1021), .A2(n1045), .A3(n1023), .ZN(n1042) );
NAND2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND3_X1 U759 ( .A1(n1048), .A2(n1049), .A3(n1026), .ZN(n1047) );
XOR2_X1 U760 ( .A(KEYINPUT26), .B(n1027), .Z(n1049) );
NAND2_X1 U761 ( .A1(n1029), .A2(n1050), .ZN(n1046) );
NAND2_X1 U762 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U763 ( .A1(n1026), .A2(n1053), .ZN(n1052) );
NAND2_X1 U764 ( .A1(n1027), .A2(n1054), .ZN(n1051) );
NAND2_X1 U765 ( .A1(n1039), .A2(n1055), .ZN(n1041) );
AND4_X1 U766 ( .A1(n1023), .A2(n1026), .A3(n1027), .A4(n1029), .ZN(n1039) );
INV_X1 U767 ( .A(n1056), .ZN(n1023) );
NOR3_X1 U768 ( .A1(n1057), .A2(G953), .A3(n1058), .ZN(n1012) );
INV_X1 U769 ( .A(n1043), .ZN(n1058) );
NAND4_X1 U770 ( .A1(n1059), .A2(n1029), .A3(n1060), .A4(n1061), .ZN(n1043) );
NOR4_X1 U771 ( .A1(n1034), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1061) );
XOR2_X1 U772 ( .A(n1065), .B(n1066), .Z(n1063) );
NOR2_X1 U773 ( .A1(G475), .A2(KEYINPUT33), .ZN(n1066) );
XNOR2_X1 U774 ( .A(n1067), .B(n1068), .ZN(n1060) );
NAND2_X1 U775 ( .A1(KEYINPUT19), .A2(G478), .ZN(n1067) );
XOR2_X1 U776 ( .A(KEYINPUT42), .B(G952), .Z(n1057) );
NAND2_X1 U777 ( .A1(n1069), .A2(n1070), .ZN(G72) );
NAND2_X1 U778 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U779 ( .A(n1073), .B(KEYINPUT2), .Z(n1071) );
XOR2_X1 U780 ( .A(KEYINPUT29), .B(n1074), .Z(n1069) );
NOR2_X1 U781 ( .A1(n1072), .A2(n1075), .ZN(n1074) );
XOR2_X1 U782 ( .A(KEYINPUT7), .B(n1076), .Z(n1075) );
INV_X1 U783 ( .A(n1073), .ZN(n1076) );
XOR2_X1 U784 ( .A(n1077), .B(n1078), .Z(n1073) );
NOR2_X1 U785 ( .A1(KEYINPUT38), .A2(n1079), .ZN(n1078) );
NOR3_X1 U786 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U787 ( .A1(G900), .A2(n1044), .ZN(n1082) );
NOR2_X1 U788 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
XOR2_X1 U789 ( .A(KEYINPUT23), .B(n1085), .Z(n1080) );
AND2_X1 U790 ( .A1(n1084), .A2(n1083), .ZN(n1085) );
XNOR2_X1 U791 ( .A(n1086), .B(n1087), .ZN(n1084) );
XNOR2_X1 U792 ( .A(n1088), .B(n1089), .ZN(n1086) );
NOR2_X1 U793 ( .A1(KEYINPUT53), .A2(n1090), .ZN(n1089) );
NAND2_X1 U794 ( .A1(n1044), .A2(n1091), .ZN(n1077) );
AND2_X1 U795 ( .A1(G953), .A2(n1092), .ZN(n1072) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1092) );
XOR2_X1 U797 ( .A(n1093), .B(n1094), .Z(G69) );
XOR2_X1 U798 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR3_X1 U799 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NOR2_X1 U800 ( .A1(G898), .A2(n1044), .ZN(n1099) );
NOR2_X1 U801 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
XOR2_X1 U802 ( .A(n1102), .B(KEYINPUT24), .Z(n1097) );
NAND2_X1 U803 ( .A1(n1101), .A2(n1100), .ZN(n1102) );
XOR2_X1 U804 ( .A(n1103), .B(n1104), .Z(n1101) );
NOR2_X1 U805 ( .A1(KEYINPUT6), .A2(n1105), .ZN(n1104) );
NOR3_X1 U806 ( .A1(n1106), .A2(KEYINPUT25), .A3(n1107), .ZN(n1095) );
NOR2_X1 U807 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U808 ( .A(KEYINPUT36), .B(n1110), .ZN(n1109) );
XOR2_X1 U809 ( .A(n1044), .B(KEYINPUT17), .Z(n1106) );
NOR2_X1 U810 ( .A1(n1111), .A2(n1044), .ZN(n1093) );
AND2_X1 U811 ( .A1(G224), .A2(G898), .ZN(n1111) );
NOR2_X1 U812 ( .A1(n1112), .A2(n1113), .ZN(G66) );
XOR2_X1 U813 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U814 ( .A1(KEYINPUT10), .A2(n1116), .ZN(n1115) );
NAND3_X1 U815 ( .A1(G902), .A2(n1117), .A3(G217), .ZN(n1114) );
XOR2_X1 U816 ( .A(KEYINPUT31), .B(n1118), .Z(n1117) );
NOR2_X1 U817 ( .A1(n1112), .A2(n1119), .ZN(G63) );
XOR2_X1 U818 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U819 ( .A1(n1122), .A2(G478), .ZN(n1120) );
NOR2_X1 U820 ( .A1(n1112), .A2(n1123), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
AND3_X1 U822 ( .A1(n1127), .A2(G475), .A3(n1122), .ZN(n1126) );
NOR2_X1 U823 ( .A1(n1128), .A2(n1127), .ZN(n1125) );
AND2_X1 U824 ( .A1(n1015), .A2(G475), .ZN(n1128) );
INV_X1 U825 ( .A(n1118), .ZN(n1015) );
XNOR2_X1 U826 ( .A(G104), .B(n1129), .ZN(G6) );
NOR2_X1 U827 ( .A1(n1130), .A2(n1131), .ZN(G57) );
XOR2_X1 U828 ( .A(KEYINPUT62), .B(n1112), .Z(n1131) );
XOR2_X1 U829 ( .A(n1132), .B(n1133), .Z(n1130) );
XOR2_X1 U830 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U831 ( .A(n1136), .B(n1105), .ZN(n1135) );
NAND2_X1 U832 ( .A1(n1122), .A2(G472), .ZN(n1136) );
XOR2_X1 U833 ( .A(n1137), .B(n1138), .Z(n1132) );
NOR2_X1 U834 ( .A1(KEYINPUT35), .A2(n1139), .ZN(n1138) );
XOR2_X1 U835 ( .A(n1140), .B(n1141), .Z(n1137) );
NOR2_X1 U836 ( .A1(G101), .A2(KEYINPUT0), .ZN(n1141) );
NOR2_X1 U837 ( .A1(n1112), .A2(n1142), .ZN(G54) );
XOR2_X1 U838 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U839 ( .A1(KEYINPUT18), .A2(n1145), .ZN(n1144) );
XOR2_X1 U840 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U841 ( .A(n1148), .B(n1149), .ZN(n1147) );
XOR2_X1 U842 ( .A(n1150), .B(n1151), .Z(n1146) );
XOR2_X1 U843 ( .A(KEYINPUT8), .B(n1152), .Z(n1151) );
NAND2_X1 U844 ( .A1(KEYINPUT9), .A2(n1153), .ZN(n1150) );
NAND2_X1 U845 ( .A1(n1122), .A2(G469), .ZN(n1143) );
NOR2_X1 U846 ( .A1(n1112), .A2(n1154), .ZN(G51) );
XOR2_X1 U847 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U848 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U849 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U850 ( .A1(n1122), .A2(n1161), .ZN(n1159) );
NOR2_X1 U851 ( .A1(n1162), .A2(n1118), .ZN(n1122) );
NOR3_X1 U852 ( .A1(n1091), .A2(n1110), .A3(n1108), .ZN(n1118) );
NAND4_X1 U853 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1108) );
NAND2_X1 U854 ( .A1(n1054), .A2(n1167), .ZN(n1164) );
NAND2_X1 U855 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND4_X1 U856 ( .A1(n1055), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1169) );
INV_X1 U857 ( .A(KEYINPUT27), .ZN(n1172) );
XNOR2_X1 U858 ( .A(KEYINPUT44), .B(n1173), .ZN(n1168) );
NAND2_X1 U859 ( .A1(KEYINPUT27), .A2(n1174), .ZN(n1163) );
NAND4_X1 U860 ( .A1(n1129), .A2(n1175), .A3(n1176), .A4(n1011), .ZN(n1110) );
NAND3_X1 U861 ( .A1(n1040), .A2(n1029), .A3(n1177), .ZN(n1011) );
NAND3_X1 U862 ( .A1(n1177), .A2(n1029), .A3(n1055), .ZN(n1129) );
NAND2_X1 U863 ( .A1(n1178), .A2(n1179), .ZN(n1091) );
AND4_X1 U864 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
NOR4_X1 U865 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1178) );
NOR3_X1 U866 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
NOR4_X1 U867 ( .A1(n1191), .A2(n1192), .A3(n1171), .A4(n1193), .ZN(n1186) );
NOR2_X1 U868 ( .A1(KEYINPUT57), .A2(n1194), .ZN(n1192) );
NOR3_X1 U869 ( .A1(n1195), .A2(n1196), .A3(n1053), .ZN(n1194) );
AND2_X1 U870 ( .A1(n1188), .A2(KEYINPUT57), .ZN(n1191) );
XOR2_X1 U871 ( .A(n1197), .B(n1198), .Z(n1155) );
XOR2_X1 U872 ( .A(KEYINPUT37), .B(G125), .Z(n1198) );
NOR2_X1 U873 ( .A1(KEYINPUT13), .A2(n1199), .ZN(n1197) );
NOR2_X1 U874 ( .A1(n1044), .A2(G952), .ZN(n1112) );
XOR2_X1 U875 ( .A(n1200), .B(n1201), .Z(G48) );
NOR3_X1 U876 ( .A1(n1202), .A2(n1189), .A3(n1188), .ZN(n1201) );
XOR2_X1 U877 ( .A(KEYINPUT58), .B(n1203), .Z(n1202) );
NAND2_X1 U878 ( .A1(KEYINPUT63), .A2(n1204), .ZN(n1200) );
XOR2_X1 U879 ( .A(G143), .B(n1185), .Z(G45) );
AND2_X1 U880 ( .A1(n1205), .A2(n1206), .ZN(n1185) );
XOR2_X1 U881 ( .A(n1153), .B(n1181), .Z(G42) );
NAND3_X1 U882 ( .A1(n1028), .A2(n1026), .A3(n1207), .ZN(n1181) );
XNOR2_X1 U883 ( .A(G137), .B(n1180), .ZN(G39) );
NAND3_X1 U884 ( .A1(n1053), .A2(n1026), .A3(n1208), .ZN(n1180) );
NOR3_X1 U885 ( .A1(n1209), .A2(n1196), .A3(n1190), .ZN(n1208) );
XOR2_X1 U886 ( .A(G134), .B(n1184), .Z(G36) );
AND3_X1 U887 ( .A1(n1026), .A2(n1040), .A3(n1205), .ZN(n1184) );
AND3_X1 U888 ( .A1(n1048), .A2(n1210), .A3(n1053), .ZN(n1205) );
NAND2_X1 U889 ( .A1(n1211), .A2(n1212), .ZN(G33) );
NAND2_X1 U890 ( .A1(G131), .A2(n1213), .ZN(n1212) );
XOR2_X1 U891 ( .A(KEYINPUT16), .B(n1214), .Z(n1211) );
NOR2_X1 U892 ( .A1(G131), .A2(n1213), .ZN(n1214) );
NAND3_X1 U893 ( .A1(n1026), .A2(n1048), .A3(n1207), .ZN(n1213) );
INV_X1 U894 ( .A(n1188), .ZN(n1207) );
NAND3_X1 U895 ( .A1(n1055), .A2(n1210), .A3(n1053), .ZN(n1188) );
XNOR2_X1 U896 ( .A(n1215), .B(KEYINPUT14), .ZN(n1053) );
INV_X1 U897 ( .A(n1193), .ZN(n1026) );
NAND2_X1 U898 ( .A1(n1033), .A2(n1216), .ZN(n1193) );
XOR2_X1 U899 ( .A(KEYINPUT12), .B(n1034), .Z(n1216) );
INV_X1 U900 ( .A(n1217), .ZN(n1034) );
XOR2_X1 U901 ( .A(n1218), .B(n1183), .Z(G30) );
NAND3_X1 U902 ( .A1(n1203), .A2(n1040), .A3(n1219), .ZN(n1183) );
AND3_X1 U903 ( .A1(n1054), .A2(n1210), .A3(n1215), .ZN(n1219) );
XNOR2_X1 U904 ( .A(n1220), .B(n1175), .ZN(G3) );
NAND3_X1 U905 ( .A1(n1048), .A2(n1177), .A3(n1021), .ZN(n1175) );
NAND2_X1 U906 ( .A1(KEYINPUT54), .A2(n1221), .ZN(n1220) );
XOR2_X1 U907 ( .A(n1222), .B(n1182), .Z(G27) );
NAND4_X1 U908 ( .A1(n1028), .A2(n1055), .A3(n1223), .A4(n1027), .ZN(n1182) );
NOR2_X1 U909 ( .A1(n1196), .A2(n1189), .ZN(n1223) );
INV_X1 U910 ( .A(n1210), .ZN(n1196) );
NAND2_X1 U911 ( .A1(n1056), .A2(n1224), .ZN(n1210) );
NAND4_X1 U912 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1226), .ZN(n1224) );
INV_X1 U913 ( .A(G900), .ZN(n1226) );
XNOR2_X1 U914 ( .A(G122), .B(n1165), .ZN(G24) );
NAND3_X1 U915 ( .A1(n1170), .A2(n1029), .A3(n1206), .ZN(n1165) );
AND3_X1 U916 ( .A1(n1054), .A2(n1227), .A3(n1228), .ZN(n1206) );
AND2_X1 U917 ( .A1(n1229), .A2(n1230), .ZN(n1029) );
XOR2_X1 U918 ( .A(G119), .B(n1231), .Z(G21) );
NOR2_X1 U919 ( .A1(n1189), .A2(n1173), .ZN(n1231) );
NAND3_X1 U920 ( .A1(n1203), .A2(n1170), .A3(n1021), .ZN(n1173) );
INV_X1 U921 ( .A(n1190), .ZN(n1203) );
NAND2_X1 U922 ( .A1(n1232), .A2(n1233), .ZN(n1190) );
XOR2_X1 U923 ( .A(n1234), .B(n1166), .Z(G18) );
NAND2_X1 U924 ( .A1(n1235), .A2(n1040), .ZN(n1166) );
AND2_X1 U925 ( .A1(n1236), .A2(n1237), .ZN(n1040) );
XOR2_X1 U926 ( .A(KEYINPUT4), .B(n1227), .Z(n1236) );
INV_X1 U927 ( .A(n1238), .ZN(n1227) );
XOR2_X1 U928 ( .A(G113), .B(n1174), .Z(G15) );
AND2_X1 U929 ( .A1(n1055), .A2(n1235), .ZN(n1174) );
AND3_X1 U930 ( .A1(n1170), .A2(n1054), .A3(n1048), .ZN(n1235) );
INV_X1 U931 ( .A(n1171), .ZN(n1048) );
NAND2_X1 U932 ( .A1(n1232), .A2(n1229), .ZN(n1171) );
INV_X1 U933 ( .A(n1233), .ZN(n1229) );
XOR2_X1 U934 ( .A(n1230), .B(KEYINPUT56), .Z(n1232) );
AND2_X1 U935 ( .A1(n1027), .A2(n1239), .ZN(n1170) );
NOR2_X1 U936 ( .A1(n1037), .A2(n1062), .ZN(n1027) );
XNOR2_X1 U937 ( .A(n1059), .B(KEYINPUT43), .ZN(n1037) );
INV_X1 U938 ( .A(n1195), .ZN(n1055) );
NAND2_X1 U939 ( .A1(n1238), .A2(n1228), .ZN(n1195) );
XNOR2_X1 U940 ( .A(G110), .B(n1176), .ZN(G12) );
NAND3_X1 U941 ( .A1(n1021), .A2(n1177), .A3(n1028), .ZN(n1176) );
AND2_X1 U942 ( .A1(n1230), .A2(n1233), .ZN(n1028) );
NAND3_X1 U943 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1233) );
NAND2_X1 U944 ( .A1(n1243), .A2(n1116), .ZN(n1242) );
OR3_X1 U945 ( .A1(n1116), .A2(n1243), .A3(G902), .ZN(n1241) );
NOR2_X1 U946 ( .A1(n1244), .A2(G234), .ZN(n1243) );
INV_X1 U947 ( .A(G217), .ZN(n1244) );
XNOR2_X1 U948 ( .A(n1245), .B(n1246), .ZN(n1116) );
XOR2_X1 U949 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U950 ( .A(G137), .B(G110), .Z(n1248) );
XOR2_X1 U951 ( .A(KEYINPUT22), .B(G146), .Z(n1247) );
XNOR2_X1 U952 ( .A(n1249), .B(n1083), .ZN(n1245) );
XOR2_X1 U953 ( .A(n1250), .B(n1251), .Z(n1249) );
AND3_X1 U954 ( .A1(G221), .A2(n1044), .A3(G234), .ZN(n1251) );
NAND2_X1 U955 ( .A1(KEYINPUT21), .A2(n1252), .ZN(n1250) );
XOR2_X1 U956 ( .A(G128), .B(n1253), .Z(n1252) );
NOR2_X1 U957 ( .A1(KEYINPUT48), .A2(n1254), .ZN(n1253) );
INV_X1 U958 ( .A(G119), .ZN(n1254) );
NAND2_X1 U959 ( .A1(G217), .A2(G902), .ZN(n1240) );
XOR2_X1 U960 ( .A(n1255), .B(G472), .Z(n1230) );
NAND2_X1 U961 ( .A1(n1256), .A2(n1162), .ZN(n1255) );
XOR2_X1 U962 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U963 ( .A(n1134), .B(n1139), .Z(n1258) );
INV_X1 U964 ( .A(n1259), .ZN(n1134) );
XOR2_X1 U965 ( .A(n1260), .B(n1261), .Z(n1257) );
XNOR2_X1 U966 ( .A(KEYINPUT51), .B(n1262), .ZN(n1261) );
NOR2_X1 U967 ( .A1(KEYINPUT15), .A2(n1263), .ZN(n1262) );
XOR2_X1 U968 ( .A(n1221), .B(n1140), .Z(n1263) );
NAND3_X1 U969 ( .A1(n1264), .A2(n1044), .A3(G210), .ZN(n1140) );
NAND2_X1 U970 ( .A1(KEYINPUT5), .A2(n1105), .ZN(n1260) );
AND3_X1 U971 ( .A1(n1215), .A2(n1239), .A3(n1054), .ZN(n1177) );
INV_X1 U972 ( .A(n1189), .ZN(n1054) );
NAND2_X1 U973 ( .A1(n1265), .A2(n1217), .ZN(n1189) );
NAND2_X1 U974 ( .A1(G214), .A2(n1266), .ZN(n1217) );
XOR2_X1 U975 ( .A(KEYINPUT41), .B(n1064), .Z(n1265) );
INV_X1 U976 ( .A(n1033), .ZN(n1064) );
XOR2_X1 U977 ( .A(n1267), .B(n1161), .Z(n1033) );
AND2_X1 U978 ( .A1(G210), .A2(n1266), .ZN(n1161) );
NAND2_X1 U979 ( .A1(n1268), .A2(n1162), .ZN(n1266) );
NAND2_X1 U980 ( .A1(n1269), .A2(n1162), .ZN(n1267) );
XOR2_X1 U981 ( .A(n1270), .B(n1157), .Z(n1269) );
XOR2_X1 U982 ( .A(n1271), .B(n1100), .Z(n1157) );
XNOR2_X1 U983 ( .A(G110), .B(G122), .ZN(n1100) );
XOR2_X1 U984 ( .A(n1105), .B(n1103), .Z(n1271) );
XOR2_X1 U985 ( .A(G113), .B(n1272), .Z(n1105) );
XOR2_X1 U986 ( .A(G119), .B(G116), .Z(n1272) );
NAND2_X1 U987 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
NAND2_X1 U988 ( .A1(n1275), .A2(n1199), .ZN(n1274) );
XOR2_X1 U989 ( .A(n1276), .B(KEYINPUT59), .Z(n1273) );
NAND2_X1 U990 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
INV_X1 U991 ( .A(n1199), .ZN(n1278) );
NAND2_X1 U992 ( .A1(G224), .A2(n1044), .ZN(n1199) );
XNOR2_X1 U993 ( .A(n1275), .B(KEYINPUT20), .ZN(n1277) );
XNOR2_X1 U994 ( .A(n1222), .B(n1279), .ZN(n1275) );
NOR2_X1 U995 ( .A1(KEYINPUT1), .A2(n1160), .ZN(n1279) );
INV_X1 U996 ( .A(n1139), .ZN(n1160) );
XOR2_X1 U997 ( .A(n1218), .B(n1280), .Z(n1139) );
INV_X1 U998 ( .A(G128), .ZN(n1218) );
INV_X1 U999 ( .A(G125), .ZN(n1222) );
NAND2_X1 U1000 ( .A1(n1056), .A2(n1281), .ZN(n1239) );
NAND4_X1 U1001 ( .A1(G953), .A2(G902), .A3(n1225), .A4(n1282), .ZN(n1281) );
INV_X1 U1002 ( .A(G898), .ZN(n1282) );
NAND3_X1 U1003 ( .A1(n1225), .A2(n1044), .A3(G952), .ZN(n1056) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1225) );
NOR2_X1 U1005 ( .A1(n1059), .A2(n1062), .ZN(n1215) );
INV_X1 U1006 ( .A(n1038), .ZN(n1062) );
NAND2_X1 U1007 ( .A1(G221), .A2(n1283), .ZN(n1038) );
NAND2_X1 U1008 ( .A1(G234), .A2(n1162), .ZN(n1283) );
XOR2_X1 U1009 ( .A(n1284), .B(G469), .Z(n1059) );
NAND2_X1 U1010 ( .A1(n1285), .A2(n1162), .ZN(n1284) );
XOR2_X1 U1011 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U1012 ( .A(n1153), .B(n1288), .Z(n1287) );
NAND2_X1 U1013 ( .A1(KEYINPUT40), .A2(n1152), .ZN(n1288) );
AND2_X1 U1014 ( .A1(G227), .A2(n1044), .ZN(n1152) );
XOR2_X1 U1015 ( .A(n1289), .B(n1148), .Z(n1286) );
XNOR2_X1 U1016 ( .A(n1259), .B(G110), .ZN(n1148) );
XOR2_X1 U1017 ( .A(n1090), .B(n1088), .Z(n1259) );
XOR2_X1 U1018 ( .A(G137), .B(G134), .Z(n1088) );
INV_X1 U1019 ( .A(G131), .ZN(n1090) );
NAND2_X1 U1020 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
OR3_X1 U1021 ( .A1(n1087), .A2(n1292), .A3(KEYINPUT49), .ZN(n1291) );
NAND2_X1 U1022 ( .A1(n1149), .A2(KEYINPUT49), .ZN(n1290) );
XOR2_X1 U1023 ( .A(n1292), .B(n1087), .Z(n1149) );
XNOR2_X1 U1024 ( .A(n1293), .B(G128), .ZN(n1087) );
NAND3_X1 U1025 ( .A1(n1294), .A2(n1295), .A3(KEYINPUT30), .ZN(n1293) );
NAND2_X1 U1026 ( .A1(KEYINPUT55), .A2(n1280), .ZN(n1295) );
OR3_X1 U1027 ( .A1(n1204), .A2(G143), .A3(KEYINPUT55), .ZN(n1294) );
INV_X1 U1028 ( .A(n1103), .ZN(n1292) );
XOR2_X1 U1029 ( .A(n1296), .B(n1297), .Z(n1103) );
XOR2_X1 U1030 ( .A(G104), .B(n1221), .Z(n1296) );
INV_X1 U1031 ( .A(G101), .ZN(n1221) );
INV_X1 U1032 ( .A(n1209), .ZN(n1021) );
NAND2_X1 U1033 ( .A1(n1238), .A2(n1237), .ZN(n1209) );
XNOR2_X1 U1034 ( .A(n1228), .B(KEYINPUT32), .ZN(n1237) );
XOR2_X1 U1035 ( .A(n1298), .B(G475), .Z(n1228) );
NAND2_X1 U1036 ( .A1(KEYINPUT11), .A2(n1065), .ZN(n1298) );
INV_X1 U1037 ( .A(n1124), .ZN(n1065) );
NOR2_X1 U1038 ( .A1(n1127), .A2(G902), .ZN(n1124) );
XOR2_X1 U1039 ( .A(n1299), .B(n1300), .Z(n1127) );
XNOR2_X1 U1040 ( .A(n1280), .B(n1301), .ZN(n1300) );
XOR2_X1 U1041 ( .A(n1302), .B(n1303), .Z(n1301) );
NOR2_X1 U1042 ( .A1(KEYINPUT39), .A2(n1083), .ZN(n1303) );
XOR2_X1 U1043 ( .A(G125), .B(n1153), .Z(n1083) );
INV_X1 U1044 ( .A(G140), .ZN(n1153) );
AND3_X1 U1045 ( .A1(n1304), .A2(n1264), .A3(G214), .ZN(n1302) );
XNOR2_X1 U1046 ( .A(n1268), .B(KEYINPUT46), .ZN(n1264) );
INV_X1 U1047 ( .A(G237), .ZN(n1268) );
XOR2_X1 U1048 ( .A(KEYINPUT3), .B(n1044), .Z(n1304) );
XOR2_X1 U1049 ( .A(G143), .B(n1204), .Z(n1280) );
INV_X1 U1050 ( .A(G146), .ZN(n1204) );
XOR2_X1 U1051 ( .A(n1305), .B(n1306), .Z(n1299) );
XOR2_X1 U1052 ( .A(G131), .B(G122), .Z(n1306) );
XNOR2_X1 U1053 ( .A(G104), .B(G113), .ZN(n1305) );
XOR2_X1 U1054 ( .A(n1068), .B(G478), .Z(n1238) );
NAND2_X1 U1055 ( .A1(n1121), .A2(n1162), .ZN(n1068) );
INV_X1 U1056 ( .A(G902), .ZN(n1162) );
XOR2_X1 U1057 ( .A(n1307), .B(n1308), .Z(n1121) );
XOR2_X1 U1058 ( .A(n1309), .B(n1310), .Z(n1308) );
NAND2_X1 U1059 ( .A1(KEYINPUT47), .A2(n1311), .ZN(n1310) );
XOR2_X1 U1060 ( .A(G122), .B(n1312), .Z(n1311) );
NOR2_X1 U1061 ( .A1(KEYINPUT60), .A2(n1234), .ZN(n1312) );
INV_X1 U1062 ( .A(G116), .ZN(n1234) );
NAND2_X1 U1063 ( .A1(KEYINPUT61), .A2(n1313), .ZN(n1309) );
NAND3_X1 U1064 ( .A1(G234), .A2(n1044), .A3(G217), .ZN(n1313) );
INV_X1 U1065 ( .A(G953), .ZN(n1044) );
XNOR2_X1 U1066 ( .A(n1297), .B(n1314), .ZN(n1307) );
NOR2_X1 U1067 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U1068 ( .A(n1317), .B(KEYINPUT50), .Z(n1316) );
NAND2_X1 U1069 ( .A1(G134), .A2(n1318), .ZN(n1317) );
NOR2_X1 U1070 ( .A1(G134), .A2(n1318), .ZN(n1315) );
XOR2_X1 U1071 ( .A(G143), .B(G128), .Z(n1318) );
XOR2_X1 U1072 ( .A(G107), .B(KEYINPUT52), .Z(n1297) );
endmodule


