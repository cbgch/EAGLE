//Key = 0011001111110101101001010111001010111110100011000000010101000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
n1439;

NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(G9) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U790 ( .A(KEYINPUT32), .B(n1103), .Z(n1099) );
NOR2_X1 U791 ( .A1(n1101), .A2(n1102), .ZN(n1103) );
NOR2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(G75) );
NOR3_X1 U793 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
NAND3_X1 U794 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1106) );
NAND2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U796 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND3_X1 U797 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
NAND2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NAND3_X1 U799 ( .A1(n1121), .A2(n1122), .A3(KEYINPUT61), .ZN(n1119) );
NAND3_X1 U800 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1116) );
NAND2_X1 U801 ( .A1(n1121), .A2(n1126), .ZN(n1124) );
NAND2_X1 U802 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U803 ( .A1(n1122), .A2(n1129), .ZN(n1128) );
INV_X1 U804 ( .A(KEYINPUT61), .ZN(n1129) );
NAND2_X1 U805 ( .A1(n1130), .A2(n1131), .ZN(n1123) );
XNOR2_X1 U806 ( .A(n1132), .B(n1133), .ZN(n1130) );
NAND3_X1 U807 ( .A1(n1131), .A2(n1134), .A3(n1121), .ZN(n1114) );
NAND2_X1 U808 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U809 ( .A1(n1125), .A2(n1137), .ZN(n1136) );
NAND2_X1 U810 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U811 ( .A1(n1118), .A2(n1140), .ZN(n1135) );
NAND2_X1 U812 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
INV_X1 U814 ( .A(n1145), .ZN(n1112) );
NOR3_X1 U815 ( .A1(n1146), .A2(G953), .A3(G952), .ZN(n1104) );
INV_X1 U816 ( .A(n1109), .ZN(n1146) );
NAND4_X1 U817 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1109) );
NOR4_X1 U818 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
XNOR2_X1 U819 ( .A(n1155), .B(n1156), .ZN(n1152) );
NAND2_X1 U820 ( .A1(n1157), .A2(KEYINPUT10), .ZN(n1155) );
XOR2_X1 U821 ( .A(n1158), .B(KEYINPUT24), .Z(n1157) );
AND2_X1 U822 ( .A1(n1159), .A2(G469), .ZN(n1151) );
NOR3_X1 U823 ( .A1(n1143), .A2(n1160), .A3(n1161), .ZN(n1149) );
INV_X1 U824 ( .A(n1162), .ZN(n1143) );
NAND2_X1 U825 ( .A1(G475), .A2(n1163), .ZN(n1147) );
XOR2_X1 U826 ( .A(n1164), .B(n1165), .Z(G72) );
NOR2_X1 U827 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U828 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U829 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U830 ( .A(KEYINPUT5), .B(n1172), .ZN(n1171) );
XOR2_X1 U831 ( .A(n1173), .B(n1174), .Z(n1168) );
NAND2_X1 U832 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
NAND2_X1 U833 ( .A1(G140), .A2(n1177), .ZN(n1176) );
XOR2_X1 U834 ( .A(KEYINPUT35), .B(n1178), .Z(n1175) );
NOR2_X1 U835 ( .A1(G140), .A2(n1177), .ZN(n1178) );
NAND2_X1 U836 ( .A1(n1179), .A2(n1180), .ZN(n1164) );
NAND2_X1 U837 ( .A1(n1108), .A2(n1110), .ZN(n1180) );
NAND3_X1 U838 ( .A1(KEYINPUT8), .A2(n1181), .A3(G953), .ZN(n1179) );
NAND2_X1 U839 ( .A1(G900), .A2(G227), .ZN(n1181) );
NAND2_X1 U840 ( .A1(n1182), .A2(n1183), .ZN(G69) );
NAND2_X1 U841 ( .A1(n1184), .A2(n1110), .ZN(n1183) );
XNOR2_X1 U842 ( .A(n1107), .B(n1185), .ZN(n1184) );
NAND2_X1 U843 ( .A1(n1186), .A2(G953), .ZN(n1182) );
NAND2_X1 U844 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U845 ( .A1(n1185), .A2(n1189), .ZN(n1188) );
INV_X1 U846 ( .A(G224), .ZN(n1189) );
NAND2_X1 U847 ( .A1(G224), .A2(n1190), .ZN(n1187) );
NAND2_X1 U848 ( .A1(G898), .A2(n1185), .ZN(n1190) );
NAND2_X1 U849 ( .A1(n1191), .A2(n1192), .ZN(n1185) );
NAND2_X1 U850 ( .A1(G953), .A2(n1193), .ZN(n1192) );
XOR2_X1 U851 ( .A(n1194), .B(n1195), .Z(n1191) );
XNOR2_X1 U852 ( .A(n1196), .B(n1197), .ZN(n1195) );
NOR2_X1 U853 ( .A1(n1198), .A2(n1199), .ZN(G66) );
XOR2_X1 U854 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U855 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U856 ( .A(G217), .B(KEYINPUT59), .ZN(n1202) );
NOR2_X1 U857 ( .A1(n1198), .A2(n1204), .ZN(G63) );
XOR2_X1 U858 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U859 ( .A1(n1207), .A2(n1203), .ZN(n1206) );
INV_X1 U860 ( .A(G478), .ZN(n1207) );
NOR3_X1 U861 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(G60) );
AND2_X1 U862 ( .A1(KEYINPUT26), .A2(n1198), .ZN(n1210) );
NOR3_X1 U863 ( .A1(KEYINPUT26), .A2(n1211), .A3(n1110), .ZN(n1209) );
XOR2_X1 U864 ( .A(n1212), .B(n1213), .Z(n1208) );
NAND3_X1 U865 ( .A1(G475), .A2(n1214), .A3(n1215), .ZN(n1212) );
XNOR2_X1 U866 ( .A(G902), .B(KEYINPUT7), .ZN(n1215) );
XNOR2_X1 U867 ( .A(n1216), .B(n1217), .ZN(G6) );
NOR2_X1 U868 ( .A1(n1141), .A2(n1218), .ZN(n1217) );
NOR2_X1 U869 ( .A1(n1198), .A2(n1219), .ZN(G57) );
XOR2_X1 U870 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U871 ( .A(n1222), .B(n1223), .Z(n1221) );
NAND2_X1 U872 ( .A1(KEYINPUT44), .A2(n1224), .ZN(n1222) );
XOR2_X1 U873 ( .A(n1225), .B(n1226), .Z(n1220) );
XNOR2_X1 U874 ( .A(G101), .B(n1227), .ZN(n1226) );
NAND3_X1 U875 ( .A1(G472), .A2(G902), .A3(n1228), .ZN(n1225) );
XOR2_X1 U876 ( .A(n1214), .B(KEYINPUT12), .Z(n1228) );
NOR2_X1 U877 ( .A1(n1198), .A2(n1229), .ZN(G54) );
XOR2_X1 U878 ( .A(n1230), .B(n1231), .Z(n1229) );
XNOR2_X1 U879 ( .A(n1232), .B(n1224), .ZN(n1231) );
NOR2_X1 U880 ( .A1(n1233), .A2(n1203), .ZN(n1232) );
INV_X1 U881 ( .A(G469), .ZN(n1233) );
NAND2_X1 U882 ( .A1(n1234), .A2(n1235), .ZN(n1230) );
NAND2_X1 U883 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
INV_X1 U884 ( .A(KEYINPUT17), .ZN(n1237) );
XOR2_X1 U885 ( .A(n1238), .B(n1239), .Z(n1236) );
NAND2_X1 U886 ( .A1(n1240), .A2(KEYINPUT17), .ZN(n1234) );
XOR2_X1 U887 ( .A(n1238), .B(n1241), .Z(n1240) );
NOR2_X1 U888 ( .A1(KEYINPUT46), .A2(n1242), .ZN(n1238) );
NOR3_X1 U889 ( .A1(n1243), .A2(n1198), .A3(n1244), .ZN(G51) );
NOR3_X1 U890 ( .A1(n1245), .A2(n1158), .A3(n1203), .ZN(n1244) );
AND2_X1 U891 ( .A1(n1211), .A2(G953), .ZN(n1198) );
XNOR2_X1 U892 ( .A(G952), .B(KEYINPUT28), .ZN(n1211) );
NOR2_X1 U893 ( .A1(n1246), .A2(n1247), .ZN(n1243) );
XNOR2_X1 U894 ( .A(n1245), .B(KEYINPUT51), .ZN(n1247) );
XNOR2_X1 U895 ( .A(n1248), .B(n1249), .ZN(n1245) );
XNOR2_X1 U896 ( .A(n1250), .B(n1251), .ZN(n1249) );
NOR2_X1 U897 ( .A1(KEYINPUT1), .A2(n1252), .ZN(n1251) );
NOR2_X1 U898 ( .A1(n1158), .A2(n1203), .ZN(n1246) );
NAND2_X1 U899 ( .A1(G902), .A2(n1214), .ZN(n1203) );
NAND2_X1 U900 ( .A1(n1253), .A2(n1254), .ZN(n1214) );
INV_X1 U901 ( .A(n1107), .ZN(n1254) );
NAND4_X1 U902 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1107) );
NOR4_X1 U903 ( .A1(n1259), .A2(n1260), .A3(n1101), .A4(n1261), .ZN(n1258) );
AND3_X1 U904 ( .A1(n1118), .A2(n1122), .A3(n1262), .ZN(n1101) );
NOR2_X1 U905 ( .A1(n1263), .A2(n1264), .ZN(n1257) );
NOR2_X1 U906 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NOR2_X1 U907 ( .A1(n1141), .A2(n1267), .ZN(n1263) );
XNOR2_X1 U908 ( .A(KEYINPUT27), .B(n1218), .ZN(n1267) );
NAND4_X1 U909 ( .A1(n1268), .A2(n1269), .A3(n1148), .A4(n1270), .ZN(n1218) );
NOR2_X1 U910 ( .A1(n1153), .A2(n1127), .ZN(n1270) );
INV_X1 U911 ( .A(n1118), .ZN(n1153) );
XOR2_X1 U912 ( .A(n1108), .B(KEYINPUT45), .Z(n1253) );
NAND4_X1 U913 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1108) );
AND4_X1 U914 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1274) );
NOR3_X1 U915 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1273) );
AND4_X1 U916 ( .A1(KEYINPUT31), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1281) );
AND2_X1 U917 ( .A1(n1122), .A2(n1120), .ZN(n1282) );
NOR2_X1 U918 ( .A1(KEYINPUT31), .A2(n1285), .ZN(n1280) );
INV_X1 U919 ( .A(n1286), .ZN(n1279) );
XNOR2_X1 U920 ( .A(G146), .B(n1278), .ZN(G48) );
NAND3_X1 U921 ( .A1(n1287), .A2(n1283), .A3(n1288), .ZN(n1278) );
XNOR2_X1 U922 ( .A(G143), .B(n1286), .ZN(G45) );
NAND3_X1 U923 ( .A1(n1284), .A2(n1283), .A3(n1289), .ZN(n1286) );
NOR3_X1 U924 ( .A1(n1141), .A2(n1290), .A3(n1291), .ZN(n1289) );
XNOR2_X1 U925 ( .A(G140), .B(n1277), .ZN(G42) );
NAND3_X1 U926 ( .A1(n1292), .A2(n1287), .A3(n1293), .ZN(n1277) );
XNOR2_X1 U927 ( .A(G137), .B(n1276), .ZN(G39) );
OR2_X1 U928 ( .A1(n1265), .A2(n1294), .ZN(n1276) );
NAND3_X1 U929 ( .A1(n1295), .A2(n1296), .A3(n1131), .ZN(n1265) );
XNOR2_X1 U930 ( .A(n1297), .B(n1285), .ZN(G36) );
NAND3_X1 U931 ( .A1(n1292), .A2(n1122), .A3(n1284), .ZN(n1285) );
NAND2_X1 U932 ( .A1(KEYINPUT15), .A2(n1172), .ZN(n1297) );
XNOR2_X1 U933 ( .A(G131), .B(n1275), .ZN(G33) );
NAND3_X1 U934 ( .A1(n1292), .A2(n1287), .A3(n1284), .ZN(n1275) );
INV_X1 U935 ( .A(n1294), .ZN(n1292) );
NAND2_X1 U936 ( .A1(n1283), .A2(n1125), .ZN(n1294) );
INV_X1 U937 ( .A(n1120), .ZN(n1125) );
NAND2_X1 U938 ( .A1(n1144), .A2(n1162), .ZN(n1120) );
XNOR2_X1 U939 ( .A(G128), .B(n1271), .ZN(G30) );
NAND3_X1 U940 ( .A1(n1283), .A2(n1122), .A3(n1288), .ZN(n1271) );
NOR3_X1 U941 ( .A1(n1133), .A2(n1132), .A3(n1298), .ZN(n1283) );
XNOR2_X1 U942 ( .A(G101), .B(n1255), .ZN(G3) );
NAND3_X1 U943 ( .A1(n1284), .A2(n1262), .A3(n1131), .ZN(n1255) );
XNOR2_X1 U944 ( .A(G125), .B(n1272), .ZN(G27) );
NAND4_X1 U945 ( .A1(n1121), .A2(n1293), .A3(n1299), .A4(n1287), .ZN(n1272) );
INV_X1 U946 ( .A(n1127), .ZN(n1287) );
NOR2_X1 U947 ( .A1(n1298), .A2(n1141), .ZN(n1299) );
AND2_X1 U948 ( .A1(n1145), .A2(n1300), .ZN(n1298) );
NAND3_X1 U949 ( .A1(G902), .A2(n1301), .A3(n1166), .ZN(n1300) );
NOR2_X1 U950 ( .A1(n1110), .A2(G900), .ZN(n1166) );
XNOR2_X1 U951 ( .A(G122), .B(n1256), .ZN(G24) );
NAND4_X1 U952 ( .A1(n1302), .A2(n1118), .A3(n1154), .A4(n1303), .ZN(n1256) );
NOR2_X1 U953 ( .A1(n1296), .A2(n1295), .ZN(n1118) );
XOR2_X1 U954 ( .A(n1304), .B(n1305), .Z(G21) );
XNOR2_X1 U955 ( .A(G119), .B(KEYINPUT0), .ZN(n1305) );
NAND4_X1 U956 ( .A1(n1121), .A2(n1288), .A3(n1131), .A4(n1306), .ZN(n1304) );
XNOR2_X1 U957 ( .A(KEYINPUT16), .B(n1268), .ZN(n1306) );
AND3_X1 U958 ( .A1(n1307), .A2(n1296), .A3(n1295), .ZN(n1288) );
INV_X1 U959 ( .A(n1308), .ZN(n1295) );
NAND2_X1 U960 ( .A1(n1309), .A2(n1310), .ZN(G18) );
NAND2_X1 U961 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND2_X1 U962 ( .A1(n1313), .A2(G116), .ZN(n1309) );
NAND2_X1 U963 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND2_X1 U964 ( .A1(n1261), .A2(n1316), .ZN(n1315) );
INV_X1 U965 ( .A(n1317), .ZN(n1261) );
OR2_X1 U966 ( .A1(n1316), .A2(n1311), .ZN(n1314) );
NOR2_X1 U967 ( .A1(KEYINPUT56), .A2(n1317), .ZN(n1311) );
NAND3_X1 U968 ( .A1(n1284), .A2(n1122), .A3(n1302), .ZN(n1317) );
INV_X1 U969 ( .A(n1266), .ZN(n1302) );
AND2_X1 U970 ( .A1(n1318), .A2(n1154), .ZN(n1122) );
XNOR2_X1 U971 ( .A(n1290), .B(KEYINPUT53), .ZN(n1318) );
INV_X1 U972 ( .A(KEYINPUT21), .ZN(n1316) );
XOR2_X1 U973 ( .A(G113), .B(n1260), .Z(G15) );
NOR3_X1 U974 ( .A1(n1138), .A2(n1127), .A3(n1266), .ZN(n1260) );
NAND3_X1 U975 ( .A1(n1307), .A2(n1268), .A3(n1121), .ZN(n1266) );
NOR2_X1 U976 ( .A1(n1269), .A2(n1133), .ZN(n1121) );
INV_X1 U977 ( .A(n1148), .ZN(n1133) );
NAND2_X1 U978 ( .A1(n1319), .A2(n1303), .ZN(n1127) );
INV_X1 U979 ( .A(n1284), .ZN(n1138) );
NOR2_X1 U980 ( .A1(n1308), .A2(n1296), .ZN(n1284) );
XOR2_X1 U981 ( .A(G110), .B(n1259), .Z(G12) );
AND3_X1 U982 ( .A1(n1131), .A2(n1262), .A3(n1293), .ZN(n1259) );
INV_X1 U983 ( .A(n1139), .ZN(n1293) );
NAND2_X1 U984 ( .A1(n1308), .A2(n1296), .ZN(n1139) );
NAND3_X1 U985 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1296) );
NAND2_X1 U986 ( .A1(n1323), .A2(n1200), .ZN(n1322) );
OR3_X1 U987 ( .A1(n1200), .A2(n1323), .A3(G902), .ZN(n1321) );
NOR2_X1 U988 ( .A1(n1324), .A2(G234), .ZN(n1323) );
INV_X1 U989 ( .A(G217), .ZN(n1324) );
XOR2_X1 U990 ( .A(n1325), .B(n1326), .Z(n1200) );
XNOR2_X1 U991 ( .A(n1327), .B(n1328), .ZN(n1326) );
XOR2_X1 U992 ( .A(G137), .B(G128), .Z(n1328) );
XNOR2_X1 U993 ( .A(n1329), .B(n1330), .ZN(n1325) );
XOR2_X1 U994 ( .A(n1331), .B(n1332), .Z(n1330) );
NAND2_X1 U995 ( .A1(n1333), .A2(G221), .ZN(n1332) );
NAND2_X1 U996 ( .A1(n1334), .A2(KEYINPUT34), .ZN(n1331) );
XNOR2_X1 U997 ( .A(n1335), .B(KEYINPUT58), .ZN(n1334) );
NAND2_X1 U998 ( .A1(G217), .A2(G902), .ZN(n1320) );
XNOR2_X1 U999 ( .A(n1336), .B(n1337), .ZN(n1308) );
XOR2_X1 U1000 ( .A(KEYINPUT9), .B(G472), .Z(n1337) );
NAND2_X1 U1001 ( .A1(n1338), .A2(n1339), .ZN(n1336) );
XOR2_X1 U1002 ( .A(n1340), .B(n1341), .Z(n1338) );
XNOR2_X1 U1003 ( .A(n1224), .B(n1223), .ZN(n1341) );
XOR2_X1 U1004 ( .A(n1342), .B(n1252), .Z(n1223) );
XNOR2_X1 U1005 ( .A(n1343), .B(n1344), .ZN(n1342) );
NOR2_X1 U1006 ( .A1(KEYINPUT39), .A2(n1327), .ZN(n1344) );
INV_X1 U1007 ( .A(n1345), .ZN(n1224) );
XOR2_X1 U1008 ( .A(n1227), .B(n1346), .Z(n1340) );
NOR2_X1 U1009 ( .A1(KEYINPUT22), .A2(G101), .ZN(n1346) );
NAND3_X1 U1010 ( .A1(n1347), .A2(n1110), .A3(G210), .ZN(n1227) );
AND4_X1 U1011 ( .A1(n1307), .A2(n1148), .A3(n1268), .A4(n1269), .ZN(n1262) );
INV_X1 U1012 ( .A(n1132), .ZN(n1269) );
NOR2_X1 U1013 ( .A1(n1348), .A2(n1160), .ZN(n1132) );
NOR2_X1 U1014 ( .A1(n1159), .A2(G469), .ZN(n1160) );
AND2_X1 U1015 ( .A1(n1349), .A2(n1159), .ZN(n1348) );
NAND2_X1 U1016 ( .A1(n1350), .A2(n1339), .ZN(n1159) );
XOR2_X1 U1017 ( .A(n1351), .B(n1239), .Z(n1350) );
XOR2_X1 U1018 ( .A(n1241), .B(n1352), .Z(n1239) );
AND2_X1 U1019 ( .A1(n1110), .A2(G227), .ZN(n1352) );
XOR2_X1 U1020 ( .A(G140), .B(n1329), .Z(n1241) );
XNOR2_X1 U1021 ( .A(n1345), .B(n1353), .ZN(n1351) );
NOR2_X1 U1022 ( .A1(KEYINPUT41), .A2(n1242), .ZN(n1353) );
XOR2_X1 U1023 ( .A(n1354), .B(n1355), .Z(n1242) );
NOR2_X1 U1024 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1025 ( .A(n1358), .B(KEYINPUT11), .Z(n1357) );
NAND2_X1 U1026 ( .A1(n1359), .A2(n1102), .ZN(n1358) );
XNOR2_X1 U1027 ( .A(KEYINPUT42), .B(n1360), .ZN(n1359) );
XNOR2_X1 U1028 ( .A(G101), .B(n1170), .ZN(n1354) );
AND2_X1 U1029 ( .A1(n1361), .A2(n1362), .ZN(n1170) );
NAND2_X1 U1030 ( .A1(G128), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1031 ( .A(n1364), .B(KEYINPUT14), .Z(n1361) );
OR2_X1 U1032 ( .A1(n1363), .A2(G128), .ZN(n1364) );
NAND3_X1 U1033 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1363) );
NAND2_X1 U1034 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
NAND2_X1 U1035 ( .A1(n1370), .A2(n1371), .ZN(n1368) );
INV_X1 U1036 ( .A(KEYINPUT50), .ZN(n1371) );
XNOR2_X1 U1037 ( .A(G146), .B(KEYINPUT43), .ZN(n1370) );
OR3_X1 U1038 ( .A1(n1369), .A2(G146), .A3(KEYINPUT50), .ZN(n1366) );
NAND2_X1 U1039 ( .A1(G146), .A2(KEYINPUT50), .ZN(n1365) );
XNOR2_X1 U1040 ( .A(n1372), .B(n1174), .ZN(n1345) );
XOR2_X1 U1041 ( .A(G137), .B(G131), .Z(n1174) );
NAND2_X1 U1042 ( .A1(KEYINPUT3), .A2(n1172), .ZN(n1372) );
XNOR2_X1 U1043 ( .A(G469), .B(KEYINPUT6), .ZN(n1349) );
NAND2_X1 U1044 ( .A1(n1145), .A2(n1373), .ZN(n1268) );
NAND4_X1 U1045 ( .A1(G953), .A2(G902), .A3(n1301), .A4(n1193), .ZN(n1373) );
INV_X1 U1046 ( .A(G898), .ZN(n1193) );
NAND3_X1 U1047 ( .A1(n1301), .A2(n1110), .A3(G952), .ZN(n1145) );
NAND2_X1 U1048 ( .A1(G237), .A2(G234), .ZN(n1301) );
NAND2_X1 U1049 ( .A1(G221), .A2(n1374), .ZN(n1148) );
NAND2_X1 U1050 ( .A1(G234), .A2(n1339), .ZN(n1374) );
INV_X1 U1051 ( .A(n1141), .ZN(n1307) );
NAND2_X1 U1052 ( .A1(n1375), .A2(n1162), .ZN(n1141) );
NAND2_X1 U1053 ( .A1(G214), .A2(n1376), .ZN(n1162) );
XNOR2_X1 U1054 ( .A(n1144), .B(KEYINPUT29), .ZN(n1375) );
XOR2_X1 U1055 ( .A(n1377), .B(n1158), .Z(n1144) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1376), .ZN(n1158) );
NAND2_X1 U1057 ( .A1(n1347), .A2(n1339), .ZN(n1376) );
XOR2_X1 U1058 ( .A(n1156), .B(KEYINPUT36), .Z(n1377) );
NAND2_X1 U1059 ( .A1(n1378), .A2(n1339), .ZN(n1156) );
XOR2_X1 U1060 ( .A(n1248), .B(n1379), .Z(n1378) );
XNOR2_X1 U1061 ( .A(n1380), .B(n1252), .ZN(n1379) );
XNOR2_X1 U1062 ( .A(G128), .B(n1381), .ZN(n1252) );
NOR2_X1 U1063 ( .A1(KEYINPUT52), .A2(n1382), .ZN(n1381) );
XOR2_X1 U1064 ( .A(G146), .B(n1383), .Z(n1382) );
NOR2_X1 U1065 ( .A1(KEYINPUT47), .A2(n1369), .ZN(n1383) );
NOR2_X1 U1066 ( .A1(KEYINPUT60), .A2(n1250), .ZN(n1380) );
NAND2_X1 U1067 ( .A1(G224), .A2(n1110), .ZN(n1250) );
XNOR2_X1 U1068 ( .A(n1384), .B(n1177), .ZN(n1248) );
INV_X1 U1069 ( .A(G125), .ZN(n1177) );
NAND2_X1 U1070 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
NAND2_X1 U1071 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
NAND2_X1 U1072 ( .A1(KEYINPUT2), .A2(n1389), .ZN(n1388) );
OR2_X1 U1073 ( .A1(n1197), .A2(KEYINPUT20), .ZN(n1389) );
INV_X1 U1074 ( .A(n1390), .ZN(n1387) );
NAND2_X1 U1075 ( .A1(n1197), .A2(n1391), .ZN(n1385) );
NAND2_X1 U1076 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NAND2_X1 U1077 ( .A1(KEYINPUT2), .A2(n1390), .ZN(n1393) );
XNOR2_X1 U1078 ( .A(n1394), .B(n1194), .ZN(n1390) );
XNOR2_X1 U1079 ( .A(n1327), .B(n1343), .ZN(n1194) );
XNOR2_X1 U1080 ( .A(G113), .B(n1312), .ZN(n1343) );
INV_X1 U1081 ( .A(G116), .ZN(n1312) );
INV_X1 U1082 ( .A(G119), .ZN(n1327) );
NAND2_X1 U1083 ( .A1(KEYINPUT37), .A2(n1196), .ZN(n1394) );
AND3_X1 U1084 ( .A1(n1395), .A2(n1396), .A3(n1397), .ZN(n1196) );
NAND2_X1 U1085 ( .A1(n1356), .A2(n1398), .ZN(n1397) );
AND2_X1 U1086 ( .A1(G107), .A2(n1360), .ZN(n1356) );
OR3_X1 U1087 ( .A1(n1398), .A2(n1360), .A3(n1102), .ZN(n1396) );
NAND2_X1 U1088 ( .A1(n1399), .A2(n1102), .ZN(n1395) );
XOR2_X1 U1089 ( .A(n1398), .B(n1360), .Z(n1399) );
XNOR2_X1 U1090 ( .A(G104), .B(KEYINPUT48), .ZN(n1360) );
NAND2_X1 U1091 ( .A1(KEYINPUT55), .A2(n1400), .ZN(n1398) );
INV_X1 U1092 ( .A(G101), .ZN(n1400) );
INV_X1 U1093 ( .A(KEYINPUT20), .ZN(n1392) );
XNOR2_X1 U1094 ( .A(G122), .B(n1329), .ZN(n1197) );
XOR2_X1 U1095 ( .A(G110), .B(KEYINPUT63), .Z(n1329) );
AND2_X1 U1096 ( .A1(n1290), .A2(n1319), .ZN(n1131) );
XNOR2_X1 U1097 ( .A(KEYINPUT57), .B(n1291), .ZN(n1319) );
INV_X1 U1098 ( .A(n1154), .ZN(n1291) );
XOR2_X1 U1099 ( .A(G478), .B(n1401), .Z(n1154) );
NOR2_X1 U1100 ( .A1(G902), .A2(n1205), .ZN(n1401) );
XOR2_X1 U1101 ( .A(n1402), .B(n1403), .Z(n1205) );
NOR2_X1 U1102 ( .A1(KEYINPUT54), .A2(n1404), .ZN(n1403) );
XOR2_X1 U1103 ( .A(n1405), .B(n1406), .Z(n1404) );
XNOR2_X1 U1104 ( .A(n1102), .B(n1407), .ZN(n1406) );
NOR2_X1 U1105 ( .A1(KEYINPUT33), .A2(n1408), .ZN(n1407) );
NOR2_X1 U1106 ( .A1(n1409), .A2(n1410), .ZN(n1408) );
XOR2_X1 U1107 ( .A(n1411), .B(KEYINPUT38), .Z(n1410) );
NAND2_X1 U1108 ( .A1(G116), .A2(n1412), .ZN(n1411) );
NOR2_X1 U1109 ( .A1(G116), .A2(n1412), .ZN(n1409) );
INV_X1 U1110 ( .A(G107), .ZN(n1102) );
NAND2_X1 U1111 ( .A1(n1413), .A2(n1414), .ZN(n1405) );
OR2_X1 U1112 ( .A1(n1172), .A2(n1415), .ZN(n1414) );
XOR2_X1 U1113 ( .A(n1416), .B(KEYINPUT19), .Z(n1413) );
NAND2_X1 U1114 ( .A1(n1172), .A2(n1415), .ZN(n1416) );
NAND3_X1 U1115 ( .A1(n1417), .A2(n1418), .A3(n1419), .ZN(n1415) );
NAND2_X1 U1116 ( .A1(n1420), .A2(n1369), .ZN(n1419) );
NAND3_X1 U1117 ( .A1(n1421), .A2(G143), .A3(KEYINPUT13), .ZN(n1418) );
INV_X1 U1118 ( .A(n1420), .ZN(n1421) );
NAND2_X1 U1119 ( .A1(KEYINPUT40), .A2(G128), .ZN(n1420) );
OR2_X1 U1120 ( .A1(G128), .A2(KEYINPUT13), .ZN(n1417) );
INV_X1 U1121 ( .A(G134), .ZN(n1172) );
NAND2_X1 U1122 ( .A1(n1333), .A2(G217), .ZN(n1402) );
AND2_X1 U1123 ( .A1(n1422), .A2(n1110), .ZN(n1333) );
XNOR2_X1 U1124 ( .A(G234), .B(KEYINPUT25), .ZN(n1422) );
INV_X1 U1125 ( .A(n1303), .ZN(n1290) );
NAND3_X1 U1126 ( .A1(n1423), .A2(n1424), .A3(n1425), .ZN(n1303) );
INV_X1 U1127 ( .A(n1161), .ZN(n1425) );
NOR2_X1 U1128 ( .A1(n1163), .A2(G475), .ZN(n1161) );
NAND3_X1 U1129 ( .A1(KEYINPUT30), .A2(G475), .A3(n1163), .ZN(n1424) );
OR2_X1 U1130 ( .A1(n1163), .A2(KEYINPUT30), .ZN(n1423) );
NAND2_X1 U1131 ( .A1(n1213), .A2(n1339), .ZN(n1163) );
INV_X1 U1132 ( .A(G902), .ZN(n1339) );
XOR2_X1 U1133 ( .A(n1426), .B(n1427), .Z(n1213) );
XNOR2_X1 U1134 ( .A(n1216), .B(n1428), .ZN(n1427) );
XNOR2_X1 U1135 ( .A(n1412), .B(G113), .ZN(n1428) );
INV_X1 U1136 ( .A(G122), .ZN(n1412) );
INV_X1 U1137 ( .A(G104), .ZN(n1216) );
XOR2_X1 U1138 ( .A(n1429), .B(n1335), .Z(n1426) );
XOR2_X1 U1139 ( .A(G125), .B(n1430), .Z(n1335) );
XOR2_X1 U1140 ( .A(G146), .B(G140), .Z(n1430) );
NAND2_X1 U1141 ( .A1(n1431), .A2(n1432), .ZN(n1429) );
NAND2_X1 U1142 ( .A1(n1433), .A2(n1434), .ZN(n1432) );
XOR2_X1 U1143 ( .A(KEYINPUT62), .B(n1435), .Z(n1434) );
XOR2_X1 U1144 ( .A(KEYINPUT4), .B(G131), .Z(n1433) );
XOR2_X1 U1145 ( .A(KEYINPUT23), .B(n1436), .Z(n1431) );
NOR2_X1 U1146 ( .A1(n1435), .A2(n1437), .ZN(n1436) );
XOR2_X1 U1147 ( .A(KEYINPUT49), .B(G131), .Z(n1437) );
XNOR2_X1 U1148 ( .A(n1438), .B(n1439), .ZN(n1435) );
AND3_X1 U1149 ( .A1(G214), .A2(n1110), .A3(n1347), .ZN(n1439) );
INV_X1 U1150 ( .A(G237), .ZN(n1347) );
INV_X1 U1151 ( .A(G953), .ZN(n1110) );
NAND2_X1 U1152 ( .A1(KEYINPUT18), .A2(n1369), .ZN(n1438) );
INV_X1 U1153 ( .A(G143), .ZN(n1369) );
endmodule


