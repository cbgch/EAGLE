//Key = 0001111000011011000000101011111111101001110001111110011000001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;

XNOR2_X1 U748 ( .A(G107), .B(n1031), .ZN(G9) );
NAND2_X1 U749 ( .A1(KEYINPUT22), .A2(n1032), .ZN(n1031) );
NAND3_X1 U750 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(G75) );
NAND2_X1 U751 ( .A1(G952), .A2(n1036), .ZN(n1035) );
NAND3_X1 U752 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NAND2_X1 U753 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND2_X1 U754 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U755 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U758 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U759 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U760 ( .A1(n1055), .A2(n1056), .ZN(n1047) );
NAND2_X1 U761 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
OR2_X1 U762 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U763 ( .A1(n1055), .A2(n1061), .A3(n1049), .ZN(n1042) );
NAND2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U765 ( .A1(n1044), .A2(n1064), .ZN(n1063) );
OR2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1046), .A2(n1067), .ZN(n1062) );
NAND3_X1 U768 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NAND3_X1 U769 ( .A1(n1071), .A2(KEYINPUT31), .A3(n1072), .ZN(n1069) );
OR2_X1 U770 ( .A1(n1072), .A2(KEYINPUT31), .ZN(n1068) );
XNOR2_X1 U771 ( .A(KEYINPUT3), .B(n1073), .ZN(n1040) );
NAND4_X1 U772 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1033) );
XOR2_X1 U773 ( .A(KEYINPUT1), .B(n1078), .Z(n1077) );
NOR3_X1 U774 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
XNOR2_X1 U775 ( .A(KEYINPUT0), .B(n1054), .ZN(n1081) );
INV_X1 U776 ( .A(n1046), .ZN(n1080) );
XOR2_X1 U777 ( .A(KEYINPUT7), .B(n1082), .Z(n1079) );
NOR2_X1 U778 ( .A1(n1083), .A2(n1071), .ZN(n1076) );
XNOR2_X1 U779 ( .A(n1084), .B(n1085), .ZN(n1075) );
XNOR2_X1 U780 ( .A(n1086), .B(G469), .ZN(n1074) );
XOR2_X1 U781 ( .A(n1087), .B(n1088), .Z(G72) );
NOR2_X1 U782 ( .A1(n1089), .A2(n1034), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR3_X1 U784 ( .A1(KEYINPUT43), .A2(n1092), .A3(n1093), .ZN(n1087) );
NOR2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
INV_X1 U786 ( .A(n1096), .ZN(n1095) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
NOR2_X1 U788 ( .A1(G900), .A2(n1034), .ZN(n1097) );
NOR2_X1 U789 ( .A1(n1098), .A2(n1096), .ZN(n1092) );
XOR2_X1 U790 ( .A(n1099), .B(n1100), .Z(n1096) );
XNOR2_X1 U791 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U793 ( .A(n1105), .B(KEYINPUT33), .Z(n1104) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U795 ( .A1(n1107), .A2(n1106), .ZN(n1103) );
XOR2_X1 U796 ( .A(n1108), .B(G131), .Z(n1106) );
NAND3_X1 U797 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1108) );
OR2_X1 U798 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U799 ( .A1(n1113), .A2(n1112), .A3(KEYINPUT53), .ZN(n1110) );
NOR2_X1 U800 ( .A1(KEYINPUT42), .A2(n1114), .ZN(n1113) );
OR2_X1 U801 ( .A1(n1115), .A2(KEYINPUT53), .ZN(n1109) );
NOR2_X1 U802 ( .A1(G953), .A2(n1039), .ZN(n1098) );
XOR2_X1 U803 ( .A(n1116), .B(n1117), .Z(G69) );
NOR2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U805 ( .A(KEYINPUT17), .B(n1120), .ZN(n1119) );
INV_X1 U806 ( .A(n1121), .ZN(n1120) );
NOR2_X1 U807 ( .A1(G898), .A2(n1034), .ZN(n1118) );
XNOR2_X1 U808 ( .A(n1122), .B(n1123), .ZN(n1116) );
NOR3_X1 U809 ( .A1(n1034), .A2(KEYINPUT2), .A3(n1124), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U811 ( .A1(KEYINPUT52), .A2(n1127), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1128), .A2(G953), .ZN(n1127) );
NOR3_X1 U813 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
XOR2_X1 U814 ( .A(KEYINPUT58), .B(n1132), .Z(n1129) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U816 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1133), .A2(n1139), .ZN(G63) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U820 ( .A1(n1142), .A2(n1138), .ZN(n1140) );
NOR2_X1 U821 ( .A1(n1133), .A2(n1143), .ZN(G60) );
XOR2_X1 U822 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U823 ( .A1(n1146), .A2(KEYINPUT9), .ZN(n1144) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1138), .ZN(n1146) );
XOR2_X1 U825 ( .A(G104), .B(n1130), .Z(G6) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1149), .ZN(G57) );
XNOR2_X1 U827 ( .A(n1133), .B(KEYINPUT27), .ZN(n1149) );
XNOR2_X1 U828 ( .A(n1150), .B(n1151), .ZN(n1148) );
NOR2_X1 U829 ( .A1(KEYINPUT10), .A2(n1152), .ZN(n1151) );
XOR2_X1 U830 ( .A(n1153), .B(n1154), .Z(n1152) );
XNOR2_X1 U831 ( .A(n1155), .B(n1156), .ZN(n1154) );
XOR2_X1 U832 ( .A(n1157), .B(n1158), .Z(n1153) );
NOR2_X1 U833 ( .A1(KEYINPUT23), .A2(n1159), .ZN(n1158) );
NOR2_X1 U834 ( .A1(n1160), .A2(n1138), .ZN(n1157) );
NOR2_X1 U835 ( .A1(n1133), .A2(n1161), .ZN(G54) );
XOR2_X1 U836 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U837 ( .A(n1164), .B(n1165), .ZN(n1163) );
XNOR2_X1 U838 ( .A(n1155), .B(n1166), .ZN(n1165) );
NOR2_X1 U839 ( .A1(KEYINPUT25), .A2(n1167), .ZN(n1166) );
XOR2_X1 U840 ( .A(n1168), .B(n1169), .Z(n1162) );
NOR2_X1 U841 ( .A1(n1170), .A2(n1138), .ZN(n1169) );
XOR2_X1 U842 ( .A(n1171), .B(KEYINPUT21), .Z(n1168) );
NAND2_X1 U843 ( .A1(KEYINPUT39), .A2(n1172), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1133), .A2(n1173), .ZN(G51) );
XNOR2_X1 U845 ( .A(n1121), .B(n1174), .ZN(n1173) );
XOR2_X1 U846 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR3_X1 U847 ( .A1(n1138), .A2(KEYINPUT59), .A3(n1085), .ZN(n1176) );
NAND2_X1 U848 ( .A1(G902), .A2(n1177), .ZN(n1138) );
NAND2_X1 U849 ( .A1(n1178), .A2(n1037), .ZN(n1177) );
NOR3_X1 U850 ( .A1(n1179), .A2(n1132), .A3(n1131), .ZN(n1037) );
NAND4_X1 U851 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1131) );
NOR3_X1 U852 ( .A1(n1184), .A2(n1032), .A3(n1185), .ZN(n1183) );
AND3_X1 U853 ( .A1(n1066), .A2(n1055), .A3(n1186), .ZN(n1032) );
NAND2_X1 U854 ( .A1(n1187), .A2(n1188), .ZN(n1182) );
XOR2_X1 U855 ( .A(n1189), .B(KEYINPUT24), .Z(n1187) );
NAND4_X1 U856 ( .A1(n1046), .A2(n1190), .A3(n1191), .A4(n1044), .ZN(n1180) );
XOR2_X1 U857 ( .A(KEYINPUT56), .B(n1192), .Z(n1191) );
INV_X1 U858 ( .A(n1193), .ZN(n1190) );
XNOR2_X1 U859 ( .A(KEYINPUT36), .B(n1130), .ZN(n1179) );
AND3_X1 U860 ( .A1(n1186), .A2(n1055), .A3(n1065), .ZN(n1130) );
XNOR2_X1 U861 ( .A(n1039), .B(KEYINPUT49), .ZN(n1178) );
AND4_X1 U862 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1039) );
AND4_X1 U863 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
NAND2_X1 U864 ( .A1(n1049), .A2(n1202), .ZN(n1196) );
NAND2_X1 U865 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NAND4_X1 U866 ( .A1(n1065), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1204) );
OR2_X1 U867 ( .A1(n1208), .A2(KEYINPUT38), .ZN(n1207) );
NAND2_X1 U868 ( .A1(KEYINPUT38), .A2(n1209), .ZN(n1206) );
NAND2_X1 U869 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1175) );
INV_X1 U871 ( .A(n1214), .ZN(n1213) );
NOR2_X1 U872 ( .A1(n1034), .A2(G952), .ZN(n1133) );
XOR2_X1 U873 ( .A(G146), .B(n1215), .Z(G48) );
NOR2_X1 U874 ( .A1(KEYINPUT35), .A2(n1194), .ZN(n1215) );
NAND2_X1 U875 ( .A1(n1216), .A2(n1065), .ZN(n1194) );
XNOR2_X1 U876 ( .A(G143), .B(n1198), .ZN(G45) );
NAND4_X1 U877 ( .A1(n1217), .A2(n1218), .A3(n1188), .A4(n1219), .ZN(n1198) );
AND2_X1 U878 ( .A1(n1208), .A2(n1205), .ZN(n1219) );
XNOR2_X1 U879 ( .A(G140), .B(n1220), .ZN(G42) );
NAND2_X1 U880 ( .A1(n1049), .A2(n1221), .ZN(n1220) );
XNOR2_X1 U881 ( .A(KEYINPUT55), .B(n1203), .ZN(n1221) );
NAND2_X1 U882 ( .A1(n1222), .A2(n1208), .ZN(n1203) );
XNOR2_X1 U883 ( .A(G137), .B(n1195), .ZN(G39) );
NAND4_X1 U884 ( .A1(n1049), .A2(n1192), .A3(n1208), .A4(n1046), .ZN(n1195) );
XNOR2_X1 U885 ( .A(G134), .B(n1201), .ZN(G36) );
NAND2_X1 U886 ( .A1(n1223), .A2(n1066), .ZN(n1201) );
XNOR2_X1 U887 ( .A(G131), .B(n1224), .ZN(G33) );
NAND2_X1 U888 ( .A1(n1223), .A2(n1065), .ZN(n1224) );
AND3_X1 U889 ( .A1(n1205), .A2(n1208), .A3(n1049), .ZN(n1223) );
NOR2_X1 U890 ( .A1(n1059), .A2(n1083), .ZN(n1049) );
INV_X1 U891 ( .A(n1060), .ZN(n1083) );
XNOR2_X1 U892 ( .A(G128), .B(n1200), .ZN(G30) );
NAND2_X1 U893 ( .A1(n1216), .A2(n1066), .ZN(n1200) );
AND3_X1 U894 ( .A1(n1208), .A2(n1188), .A3(n1192), .ZN(n1216) );
NOR2_X1 U895 ( .A1(n1070), .A2(n1210), .ZN(n1208) );
INV_X1 U896 ( .A(n1225), .ZN(n1210) );
XNOR2_X1 U897 ( .A(G101), .B(n1181), .ZN(G3) );
NAND3_X1 U898 ( .A1(n1046), .A2(n1186), .A3(n1205), .ZN(n1181) );
XNOR2_X1 U899 ( .A(G125), .B(n1199), .ZN(G27) );
NAND4_X1 U900 ( .A1(n1222), .A2(n1188), .A3(n1044), .A4(n1225), .ZN(n1199) );
NAND2_X1 U901 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND2_X1 U902 ( .A1(n1228), .A2(n1091), .ZN(n1226) );
INV_X1 U903 ( .A(G900), .ZN(n1091) );
AND3_X1 U904 ( .A1(n1054), .A2(n1053), .A3(n1065), .ZN(n1222) );
XNOR2_X1 U905 ( .A(n1229), .B(n1230), .ZN(G24) );
NOR2_X1 U906 ( .A1(n1057), .A2(n1189), .ZN(n1230) );
NAND3_X1 U907 ( .A1(n1055), .A2(n1044), .A3(n1231), .ZN(n1189) );
NOR3_X1 U908 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
NOR2_X1 U909 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
AND2_X1 U910 ( .A1(n1126), .A2(n1228), .ZN(n1236) );
INV_X1 U911 ( .A(n1227), .ZN(n1235) );
AND2_X1 U912 ( .A1(n1054), .A2(n1237), .ZN(n1055) );
XNOR2_X1 U913 ( .A(G119), .B(n1238), .ZN(G21) );
NAND4_X1 U914 ( .A1(KEYINPUT34), .A2(n1192), .A3(n1239), .A4(n1046), .ZN(n1238) );
NOR2_X1 U915 ( .A1(n1240), .A2(n1193), .ZN(n1239) );
NOR2_X1 U916 ( .A1(n1237), .A2(n1054), .ZN(n1192) );
XOR2_X1 U917 ( .A(G116), .B(n1184), .Z(G18) );
AND2_X1 U918 ( .A1(n1241), .A2(n1066), .ZN(n1184) );
NOR2_X1 U919 ( .A1(n1217), .A2(n1234), .ZN(n1066) );
INV_X1 U920 ( .A(n1218), .ZN(n1234) );
XOR2_X1 U921 ( .A(G113), .B(n1132), .Z(G15) );
AND2_X1 U922 ( .A1(n1241), .A2(n1065), .ZN(n1132) );
NOR2_X1 U923 ( .A1(n1218), .A2(n1232), .ZN(n1065) );
INV_X1 U924 ( .A(n1217), .ZN(n1232) );
NOR3_X1 U925 ( .A1(n1193), .A2(n1240), .A3(n1051), .ZN(n1241) );
INV_X1 U926 ( .A(n1205), .ZN(n1051) );
NOR2_X1 U927 ( .A1(n1054), .A2(n1053), .ZN(n1205) );
INV_X1 U928 ( .A(n1044), .ZN(n1240) );
NAND2_X1 U929 ( .A1(n1242), .A2(n1243), .ZN(n1044) );
OR2_X1 U930 ( .A1(n1070), .A2(KEYINPUT31), .ZN(n1243) );
NAND3_X1 U931 ( .A1(n1244), .A2(n1072), .A3(KEYINPUT31), .ZN(n1242) );
XOR2_X1 U932 ( .A(G110), .B(n1185), .Z(G12) );
AND4_X1 U933 ( .A1(n1053), .A2(n1046), .A3(n1054), .A4(n1186), .ZN(n1185) );
NOR2_X1 U934 ( .A1(n1193), .A2(n1070), .ZN(n1186) );
INV_X1 U935 ( .A(n1211), .ZN(n1070) );
NOR2_X1 U936 ( .A1(n1072), .A2(n1071), .ZN(n1211) );
INV_X1 U937 ( .A(n1244), .ZN(n1071) );
NAND2_X1 U938 ( .A1(G221), .A2(n1245), .ZN(n1244) );
XOR2_X1 U939 ( .A(KEYINPUT32), .B(n1246), .Z(n1245) );
NOR2_X1 U940 ( .A1(G902), .A2(n1247), .ZN(n1246) );
NAND2_X1 U941 ( .A1(n1248), .A2(n1249), .ZN(n1072) );
NAND2_X1 U942 ( .A1(n1086), .A2(n1250), .ZN(n1249) );
NAND2_X1 U943 ( .A1(KEYINPUT14), .A2(n1251), .ZN(n1250) );
NAND2_X1 U944 ( .A1(KEYINPUT11), .A2(G469), .ZN(n1251) );
INV_X1 U945 ( .A(n1252), .ZN(n1086) );
NAND2_X1 U946 ( .A1(n1253), .A2(n1170), .ZN(n1248) );
INV_X1 U947 ( .A(G469), .ZN(n1170) );
NAND2_X1 U948 ( .A1(KEYINPUT11), .A2(n1254), .ZN(n1253) );
NAND2_X1 U949 ( .A1(KEYINPUT14), .A2(n1252), .ZN(n1254) );
NAND3_X1 U950 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1252) );
NAND2_X1 U951 ( .A1(n1258), .A2(n1259), .ZN(n1256) );
INV_X1 U952 ( .A(KEYINPUT8), .ZN(n1259) );
XOR2_X1 U953 ( .A(n1167), .B(n1260), .Z(n1258) );
NAND3_X1 U954 ( .A1(n1260), .A2(n1167), .A3(KEYINPUT8), .ZN(n1255) );
XNOR2_X1 U955 ( .A(n1261), .B(n1262), .ZN(n1167) );
XOR2_X1 U956 ( .A(KEYINPUT26), .B(n1263), .Z(n1262) );
NOR2_X1 U957 ( .A1(G953), .A2(n1090), .ZN(n1263) );
INV_X1 U958 ( .A(G227), .ZN(n1090) );
XNOR2_X1 U959 ( .A(n1264), .B(n1265), .ZN(n1260) );
XNOR2_X1 U960 ( .A(n1172), .B(n1107), .ZN(n1265) );
INV_X1 U961 ( .A(n1164), .ZN(n1107) );
XOR2_X1 U962 ( .A(G143), .B(n1266), .Z(n1164) );
XNOR2_X1 U963 ( .A(n1267), .B(n1268), .ZN(n1172) );
XNOR2_X1 U964 ( .A(n1155), .B(KEYINPUT16), .ZN(n1264) );
NAND2_X1 U965 ( .A1(n1188), .A2(n1269), .ZN(n1193) );
NAND2_X1 U966 ( .A1(n1227), .A2(n1270), .ZN(n1269) );
NAND2_X1 U967 ( .A1(n1228), .A2(n1126), .ZN(n1270) );
INV_X1 U968 ( .A(G898), .ZN(n1126) );
AND3_X1 U969 ( .A1(G902), .A2(n1073), .A3(G953), .ZN(n1228) );
NAND3_X1 U970 ( .A1(n1073), .A2(n1034), .A3(G952), .ZN(n1227) );
NAND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n1073) );
INV_X1 U972 ( .A(n1057), .ZN(n1188) );
NAND2_X1 U973 ( .A1(n1059), .A2(n1271), .ZN(n1057) );
XNOR2_X1 U974 ( .A(KEYINPUT60), .B(n1060), .ZN(n1271) );
NAND2_X1 U975 ( .A1(G214), .A2(n1272), .ZN(n1060) );
NAND2_X1 U976 ( .A1(n1273), .A2(n1274), .ZN(n1059) );
NAND2_X1 U977 ( .A1(n1275), .A2(n1085), .ZN(n1274) );
INV_X1 U978 ( .A(n1084), .ZN(n1275) );
NAND2_X1 U979 ( .A1(n1276), .A2(n1084), .ZN(n1273) );
NAND2_X1 U980 ( .A1(n1277), .A2(n1257), .ZN(n1084) );
XNOR2_X1 U981 ( .A(n1121), .B(n1278), .ZN(n1277) );
NOR3_X1 U982 ( .A1(n1279), .A2(KEYINPUT51), .A3(n1214), .ZN(n1278) );
NOR3_X1 U983 ( .A1(n1280), .A2(G953), .A3(n1125), .ZN(n1214) );
INV_X1 U984 ( .A(G224), .ZN(n1125) );
XOR2_X1 U985 ( .A(n1212), .B(KEYINPUT47), .Z(n1279) );
NAND2_X1 U986 ( .A1(n1280), .A2(n1281), .ZN(n1212) );
NAND2_X1 U987 ( .A1(G224), .A2(n1034), .ZN(n1281) );
XOR2_X1 U988 ( .A(n1156), .B(G125), .Z(n1280) );
XNOR2_X1 U989 ( .A(n1282), .B(n1283), .ZN(n1121) );
XOR2_X1 U990 ( .A(n1284), .B(n1285), .Z(n1283) );
XOR2_X1 U991 ( .A(G113), .B(G110), .Z(n1285) );
NOR2_X1 U992 ( .A1(KEYINPUT61), .A2(n1229), .ZN(n1284) );
XOR2_X1 U993 ( .A(n1286), .B(n1287), .Z(n1282) );
XNOR2_X1 U994 ( .A(n1288), .B(n1289), .ZN(n1287) );
NAND2_X1 U995 ( .A1(n1290), .A2(n1291), .ZN(n1286) );
OR2_X1 U996 ( .A1(n1267), .A2(n1268), .ZN(n1291) );
NAND2_X1 U997 ( .A1(n1292), .A2(n1268), .ZN(n1290) );
XNOR2_X1 U998 ( .A(KEYINPUT45), .B(n1267), .ZN(n1292) );
XNOR2_X1 U999 ( .A(G101), .B(G104), .ZN(n1267) );
XOR2_X1 U1000 ( .A(n1085), .B(KEYINPUT46), .Z(n1276) );
NAND2_X1 U1001 ( .A1(G210), .A2(n1272), .ZN(n1085) );
NAND2_X1 U1002 ( .A1(n1293), .A2(n1257), .ZN(n1272) );
XNOR2_X1 U1003 ( .A(n1294), .B(n1160), .ZN(n1054) );
INV_X1 U1004 ( .A(G472), .ZN(n1160) );
NAND2_X1 U1005 ( .A1(n1295), .A2(n1257), .ZN(n1294) );
XOR2_X1 U1006 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U1007 ( .A(n1298), .B(n1299), .ZN(n1297) );
INV_X1 U1008 ( .A(n1150), .ZN(n1299) );
XOR2_X1 U1009 ( .A(G101), .B(n1300), .Z(n1150) );
NOR3_X1 U1010 ( .A1(n1301), .A2(G237), .A3(n1302), .ZN(n1300) );
INV_X1 U1011 ( .A(G210), .ZN(n1302) );
XNOR2_X1 U1012 ( .A(KEYINPUT57), .B(n1034), .ZN(n1301) );
NOR2_X1 U1013 ( .A1(KEYINPUT13), .A2(n1155), .ZN(n1298) );
XOR2_X1 U1014 ( .A(n1303), .B(n1114), .Z(n1155) );
XNOR2_X1 U1015 ( .A(n1304), .B(n1112), .ZN(n1303) );
INV_X1 U1016 ( .A(G137), .ZN(n1112) );
NAND2_X1 U1017 ( .A1(KEYINPUT63), .A2(G131), .ZN(n1304) );
XOR2_X1 U1018 ( .A(n1156), .B(n1159), .Z(n1296) );
XNOR2_X1 U1019 ( .A(n1305), .B(G113), .ZN(n1159) );
NAND3_X1 U1020 ( .A1(n1306), .A2(n1307), .A3(KEYINPUT5), .ZN(n1305) );
NAND2_X1 U1021 ( .A1(n1308), .A2(n1288), .ZN(n1307) );
XOR2_X1 U1022 ( .A(n1309), .B(KEYINPUT4), .Z(n1308) );
NAND2_X1 U1023 ( .A1(n1310), .A2(n1311), .ZN(n1306) );
XOR2_X1 U1024 ( .A(n1309), .B(KEYINPUT62), .Z(n1311) );
XNOR2_X1 U1025 ( .A(n1289), .B(KEYINPUT40), .ZN(n1309) );
XOR2_X1 U1026 ( .A(G116), .B(KEYINPUT41), .Z(n1289) );
XOR2_X1 U1027 ( .A(n1312), .B(n1266), .Z(n1156) );
NAND2_X1 U1028 ( .A1(KEYINPUT6), .A2(n1313), .ZN(n1312) );
NOR2_X1 U1029 ( .A1(n1218), .A2(n1217), .ZN(n1046) );
XOR2_X1 U1030 ( .A(n1314), .B(n1147), .Z(n1217) );
INV_X1 U1031 ( .A(G475), .ZN(n1147) );
NAND2_X1 U1032 ( .A1(n1145), .A2(n1257), .ZN(n1314) );
XNOR2_X1 U1033 ( .A(n1315), .B(n1316), .ZN(n1145) );
XNOR2_X1 U1034 ( .A(n1317), .B(n1318), .ZN(n1316) );
NOR2_X1 U1035 ( .A1(G122), .A2(KEYINPUT44), .ZN(n1318) );
NAND2_X1 U1036 ( .A1(KEYINPUT48), .A2(n1319), .ZN(n1317) );
XOR2_X1 U1037 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1038 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1039 ( .A(n1324), .B(n1325), .ZN(n1323) );
NOR2_X1 U1040 ( .A1(KEYINPUT19), .A2(n1326), .ZN(n1325) );
XNOR2_X1 U1041 ( .A(G146), .B(KEYINPUT20), .ZN(n1326) );
NAND2_X1 U1042 ( .A1(KEYINPUT54), .A2(n1099), .ZN(n1324) );
NAND3_X1 U1043 ( .A1(n1293), .A2(n1034), .A3(G214), .ZN(n1322) );
INV_X1 U1044 ( .A(G953), .ZN(n1034) );
INV_X1 U1045 ( .A(G237), .ZN(n1293) );
XNOR2_X1 U1046 ( .A(G125), .B(n1327), .ZN(n1320) );
XNOR2_X1 U1047 ( .A(n1313), .B(G131), .ZN(n1327) );
INV_X1 U1048 ( .A(G143), .ZN(n1313) );
XNOR2_X1 U1049 ( .A(G104), .B(n1328), .ZN(n1315) );
XOR2_X1 U1050 ( .A(KEYINPUT18), .B(G113), .Z(n1328) );
XOR2_X1 U1051 ( .A(n1329), .B(n1142), .Z(n1218) );
INV_X1 U1052 ( .A(G478), .ZN(n1142) );
OR2_X1 U1053 ( .A1(n1141), .A2(G902), .ZN(n1329) );
XNOR2_X1 U1054 ( .A(n1330), .B(n1331), .ZN(n1141) );
XOR2_X1 U1055 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1056 ( .A(n1334), .B(n1229), .ZN(n1333) );
INV_X1 U1057 ( .A(G122), .ZN(n1229) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1335), .ZN(n1334) );
XNOR2_X1 U1059 ( .A(G128), .B(G143), .ZN(n1332) );
XNOR2_X1 U1060 ( .A(n1268), .B(n1336), .ZN(n1330) );
XNOR2_X1 U1061 ( .A(n1337), .B(n1114), .ZN(n1336) );
INV_X1 U1062 ( .A(n1115), .ZN(n1114) );
XOR2_X1 U1063 ( .A(G134), .B(KEYINPUT29), .Z(n1115) );
NOR2_X1 U1064 ( .A1(G116), .A2(KEYINPUT37), .ZN(n1337) );
XOR2_X1 U1065 ( .A(G107), .B(KEYINPUT50), .Z(n1268) );
INV_X1 U1066 ( .A(n1237), .ZN(n1053) );
XOR2_X1 U1067 ( .A(n1082), .B(KEYINPUT28), .Z(n1237) );
XOR2_X1 U1068 ( .A(n1338), .B(n1137), .Z(n1082) );
NAND2_X1 U1069 ( .A1(G217), .A2(n1339), .ZN(n1137) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1257), .ZN(n1339) );
INV_X1 U1071 ( .A(G902), .ZN(n1257) );
OR2_X1 U1072 ( .A1(n1136), .A2(G902), .ZN(n1338) );
XNOR2_X1 U1073 ( .A(n1340), .B(n1341), .ZN(n1136) );
XOR2_X1 U1074 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1075 ( .A(n1344), .B(n1101), .ZN(n1343) );
INV_X1 U1076 ( .A(G125), .ZN(n1101) );
NAND2_X1 U1077 ( .A1(n1335), .A2(G221), .ZN(n1344) );
NOR2_X1 U1078 ( .A1(n1247), .A2(G953), .ZN(n1335) );
INV_X1 U1079 ( .A(G234), .ZN(n1247) );
XNOR2_X1 U1080 ( .A(KEYINPUT20), .B(G137), .ZN(n1342) );
XOR2_X1 U1081 ( .A(n1345), .B(n1261), .Z(n1340) );
XNOR2_X1 U1082 ( .A(G110), .B(n1346), .ZN(n1261) );
INV_X1 U1083 ( .A(n1099), .ZN(n1346) );
XOR2_X1 U1084 ( .A(G140), .B(KEYINPUT30), .Z(n1099) );
XOR2_X1 U1085 ( .A(n1347), .B(n1266), .Z(n1345) );
XNOR2_X1 U1086 ( .A(n1348), .B(G146), .ZN(n1266) );
INV_X1 U1087 ( .A(G128), .ZN(n1348) );
NAND2_X1 U1088 ( .A1(KEYINPUT12), .A2(n1288), .ZN(n1347) );
INV_X1 U1089 ( .A(n1310), .ZN(n1288) );
XOR2_X1 U1090 ( .A(G119), .B(KEYINPUT15), .Z(n1310) );
endmodule


