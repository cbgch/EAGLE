//Key = 0010010011010110000001000001011000011110011111011011011111111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322;

XNOR2_X1 U734 ( .A(G107), .B(n1009), .ZN(G9) );
NOR2_X1 U735 ( .A1(n1010), .A2(n1011), .ZN(G75) );
NOR4_X1 U736 ( .A1(G953), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1011) );
NOR2_X1 U737 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U738 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR3_X1 U739 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NOR2_X1 U740 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U741 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U742 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(n1022) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR3_X1 U747 ( .A1(n1031), .A2(n1036), .A3(n1025), .ZN(n1017) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1019), .ZN(n1038) );
INV_X1 U750 ( .A(n1040), .ZN(n1019) );
NOR2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U753 ( .A1(n1045), .A2(n1021), .ZN(n1037) );
INV_X1 U754 ( .A(n1046), .ZN(n1021) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
INV_X1 U756 ( .A(n1049), .ZN(n1031) );
NOR3_X1 U757 ( .A1(n1012), .A2(G953), .A3(G952), .ZN(n1010) );
AND4_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1012) );
NOR4_X1 U759 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
XOR2_X1 U760 ( .A(n1058), .B(n1059), .Z(n1057) );
NOR2_X1 U761 ( .A1(n1060), .A2(KEYINPUT40), .ZN(n1059) );
NOR4_X1 U762 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1052) );
AND2_X1 U763 ( .A1(G469), .A2(n1065), .ZN(n1064) );
NOR2_X1 U764 ( .A1(G469), .A2(n1066), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U766 ( .A1(KEYINPUT39), .A2(n1065), .ZN(n1068) );
AND2_X1 U767 ( .A1(KEYINPUT47), .A2(n1069), .ZN(n1065) );
AND2_X1 U768 ( .A1(n1069), .A2(KEYINPUT39), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1062) );
INV_X1 U770 ( .A(KEYINPUT25), .ZN(n1071) );
NOR2_X1 U771 ( .A1(KEYINPUT25), .A2(n1072), .ZN(n1061) );
XNOR2_X1 U772 ( .A(n1073), .B(n1074), .ZN(n1051) );
NAND2_X1 U773 ( .A1(KEYINPUT43), .A2(n1075), .ZN(n1074) );
XOR2_X1 U774 ( .A(n1076), .B(n1077), .Z(G72) );
XOR2_X1 U775 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U776 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U777 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U778 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U779 ( .A1(KEYINPUT11), .A2(n1086), .ZN(n1084) );
NOR2_X1 U780 ( .A1(G900), .A2(n1087), .ZN(n1080) );
NOR3_X1 U781 ( .A1(KEYINPUT31), .A2(n1088), .A3(n1089), .ZN(n1078) );
NOR2_X1 U782 ( .A1(KEYINPUT44), .A2(n1090), .ZN(n1089) );
NOR3_X1 U783 ( .A1(n1091), .A2(n1092), .A3(n1087), .ZN(n1090) );
NOR2_X1 U784 ( .A1(n1093), .A2(n1094), .ZN(n1088) );
INV_X1 U785 ( .A(KEYINPUT44), .ZN(n1094) );
NOR2_X1 U786 ( .A1(n1095), .A2(n1087), .ZN(n1093) );
NOR2_X1 U787 ( .A1(n1092), .A2(n1091), .ZN(n1095) );
NOR2_X1 U788 ( .A1(n1096), .A2(G953), .ZN(n1076) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U790 ( .A(KEYINPUT3), .B(n1099), .Z(n1098) );
NAND2_X1 U791 ( .A1(n1100), .A2(n1101), .ZN(G69) );
NAND2_X1 U792 ( .A1(n1102), .A2(n1087), .ZN(n1101) );
XNOR2_X1 U793 ( .A(n1103), .B(n1104), .ZN(n1102) );
NAND2_X1 U794 ( .A1(n1105), .A2(G953), .ZN(n1100) );
NAND2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U796 ( .A1(n1104), .A2(n1108), .ZN(n1107) );
NAND2_X1 U797 ( .A1(G224), .A2(n1109), .ZN(n1106) );
NAND2_X1 U798 ( .A1(G898), .A2(n1104), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1110), .A2(n1111), .ZN(n1104) );
NAND2_X1 U800 ( .A1(G953), .A2(n1112), .ZN(n1111) );
XOR2_X1 U801 ( .A(n1113), .B(n1114), .Z(n1110) );
XNOR2_X1 U802 ( .A(n1115), .B(KEYINPUT24), .ZN(n1114) );
NAND2_X1 U803 ( .A1(KEYINPUT35), .A2(n1116), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1117), .A2(n1118), .ZN(G66) );
XOR2_X1 U805 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U806 ( .A1(n1121), .A2(n1073), .ZN(n1119) );
INV_X1 U807 ( .A(n1122), .ZN(n1073) );
NOR2_X1 U808 ( .A1(n1117), .A2(n1123), .ZN(G63) );
NOR3_X1 U809 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U811 ( .A1(KEYINPUT1), .A2(n1129), .ZN(n1127) );
XOR2_X1 U812 ( .A(KEYINPUT63), .B(n1130), .Z(n1129) );
NOR3_X1 U813 ( .A1(n1131), .A2(KEYINPUT1), .A3(n1130), .ZN(n1125) );
AND2_X1 U814 ( .A1(n1130), .A2(KEYINPUT1), .ZN(n1124) );
AND2_X1 U815 ( .A1(n1121), .A2(G478), .ZN(n1130) );
NOR2_X1 U816 ( .A1(n1117), .A2(n1132), .ZN(G60) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND3_X1 U818 ( .A1(n1121), .A2(G475), .A3(KEYINPUT41), .ZN(n1133) );
XNOR2_X1 U819 ( .A(G104), .B(n1135), .ZN(G6) );
NOR2_X1 U820 ( .A1(n1117), .A2(n1136), .ZN(G57) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U822 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U823 ( .A1(KEYINPUT27), .A2(n1141), .ZN(n1140) );
NAND2_X1 U824 ( .A1(n1121), .A2(G472), .ZN(n1139) );
XOR2_X1 U825 ( .A(G101), .B(n1142), .Z(n1137) );
NOR2_X1 U826 ( .A1(KEYINPUT26), .A2(n1143), .ZN(n1142) );
XOR2_X1 U827 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U828 ( .A1(KEYINPUT0), .A2(n1146), .ZN(n1144) );
NOR2_X1 U829 ( .A1(n1117), .A2(n1147), .ZN(G54) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U831 ( .A(n1150), .B(n1151), .ZN(n1149) );
NAND2_X1 U832 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
OR2_X1 U833 ( .A1(KEYINPUT57), .A2(n1154), .ZN(n1153) );
NAND2_X1 U834 ( .A1(KEYINPUT38), .A2(n1154), .ZN(n1152) );
NAND2_X1 U835 ( .A1(n1121), .A2(G469), .ZN(n1154) );
NOR2_X1 U836 ( .A1(n1117), .A2(n1155), .ZN(G51) );
XOR2_X1 U837 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U838 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U839 ( .A1(n1160), .A2(KEYINPUT13), .ZN(n1159) );
XOR2_X1 U840 ( .A(n1161), .B(KEYINPUT56), .Z(n1160) );
NAND2_X1 U841 ( .A1(n1162), .A2(n1121), .ZN(n1158) );
AND2_X1 U842 ( .A1(n1163), .A2(n1014), .ZN(n1121) );
OR3_X1 U843 ( .A1(n1097), .A2(n1099), .A3(n1103), .ZN(n1014) );
NAND4_X1 U844 ( .A1(n1135), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1103) );
NOR4_X1 U845 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
INV_X1 U846 ( .A(n1009), .ZN(n1170) );
NAND3_X1 U847 ( .A1(n1047), .A2(n1171), .A3(n1042), .ZN(n1009) );
NAND2_X1 U848 ( .A1(n1027), .A2(n1172), .ZN(n1165) );
NAND2_X1 U849 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XNOR2_X1 U850 ( .A(KEYINPUT55), .B(n1175), .ZN(n1174) );
XOR2_X1 U851 ( .A(n1176), .B(KEYINPUT4), .Z(n1173) );
NAND3_X1 U852 ( .A1(n1042), .A2(n1171), .A3(n1048), .ZN(n1135) );
NAND4_X1 U853 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1097) );
AND4_X1 U854 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
XNOR2_X1 U855 ( .A(G902), .B(KEYINPUT58), .ZN(n1163) );
XNOR2_X1 U856 ( .A(n1060), .B(KEYINPUT51), .ZN(n1162) );
INV_X1 U857 ( .A(n1185), .ZN(n1060) );
NOR2_X1 U858 ( .A1(n1087), .A2(G952), .ZN(n1117) );
XNOR2_X1 U859 ( .A(n1181), .B(n1186), .ZN(G48) );
XNOR2_X1 U860 ( .A(KEYINPUT7), .B(n1187), .ZN(n1186) );
NAND3_X1 U861 ( .A1(n1048), .A2(n1027), .A3(n1188), .ZN(n1181) );
NAND2_X1 U862 ( .A1(n1189), .A2(n1190), .ZN(G45) );
NAND2_X1 U863 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U864 ( .A(KEYINPUT30), .B(n1193), .Z(n1189) );
NOR2_X1 U865 ( .A1(n1191), .A2(n1192), .ZN(n1193) );
INV_X1 U866 ( .A(n1179), .ZN(n1191) );
NAND4_X1 U867 ( .A1(n1056), .A2(n1194), .A3(n1027), .A4(n1195), .ZN(n1179) );
XNOR2_X1 U868 ( .A(G140), .B(n1177), .ZN(G42) );
NAND3_X1 U869 ( .A1(n1196), .A2(n1042), .A3(n1049), .ZN(n1177) );
XNOR2_X1 U870 ( .A(G137), .B(n1178), .ZN(G39) );
NAND3_X1 U871 ( .A1(n1188), .A2(n1040), .A3(n1049), .ZN(n1178) );
XNOR2_X1 U872 ( .A(G134), .B(n1184), .ZN(G36) );
NAND3_X1 U873 ( .A1(n1194), .A2(n1047), .A3(n1049), .ZN(n1184) );
XNOR2_X1 U874 ( .A(G131), .B(n1183), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1194), .A2(n1048), .A3(n1049), .ZN(n1183) );
NOR2_X1 U876 ( .A1(n1028), .A2(n1055), .ZN(n1049) );
AND3_X1 U877 ( .A1(n1042), .A2(n1197), .A3(n1033), .ZN(n1194) );
XNOR2_X1 U878 ( .A(n1198), .B(n1199), .ZN(G30) );
NOR2_X1 U879 ( .A1(KEYINPUT19), .A2(n1182), .ZN(n1199) );
NAND3_X1 U880 ( .A1(n1047), .A2(n1027), .A3(n1188), .ZN(n1182) );
AND4_X1 U881 ( .A1(n1200), .A2(n1042), .A3(n1201), .A4(n1197), .ZN(n1188) );
XOR2_X1 U882 ( .A(G101), .B(n1202), .Z(G3) );
NOR2_X1 U883 ( .A1(n1203), .A2(n1176), .ZN(n1202) );
NAND4_X1 U884 ( .A1(n1033), .A2(n1040), .A3(n1042), .A4(n1204), .ZN(n1176) );
XOR2_X1 U885 ( .A(n1205), .B(n1099), .Z(G27) );
AND3_X1 U886 ( .A1(n1196), .A2(n1027), .A3(n1046), .ZN(n1099) );
AND4_X1 U887 ( .A1(n1048), .A2(n1072), .A3(n1201), .A4(n1197), .ZN(n1196) );
NAND2_X1 U888 ( .A1(n1206), .A2(n1207), .ZN(n1197) );
NAND2_X1 U889 ( .A1(n1208), .A2(n1091), .ZN(n1207) );
INV_X1 U890 ( .A(G900), .ZN(n1091) );
XNOR2_X1 U891 ( .A(G125), .B(KEYINPUT54), .ZN(n1205) );
XNOR2_X1 U892 ( .A(n1164), .B(n1209), .ZN(G24) );
NOR2_X1 U893 ( .A1(KEYINPUT12), .A2(n1210), .ZN(n1209) );
NAND4_X1 U894 ( .A1(n1056), .A2(n1046), .A3(n1171), .A4(n1195), .ZN(n1164) );
NOR3_X1 U895 ( .A1(n1025), .A2(n1211), .A3(n1203), .ZN(n1171) );
NAND2_X1 U896 ( .A1(n1072), .A2(n1034), .ZN(n1025) );
XOR2_X1 U897 ( .A(G119), .B(n1212), .Z(G21) );
NOR2_X1 U898 ( .A1(n1203), .A2(n1175), .ZN(n1212) );
NAND4_X1 U899 ( .A1(n1200), .A2(n1040), .A3(n1213), .A4(n1046), .ZN(n1175) );
NOR2_X1 U900 ( .A1(n1211), .A2(n1034), .ZN(n1213) );
INV_X1 U901 ( .A(n1027), .ZN(n1203) );
XNOR2_X1 U902 ( .A(n1214), .B(n1169), .ZN(G18) );
AND2_X1 U903 ( .A1(n1215), .A2(n1047), .ZN(n1169) );
NOR2_X1 U904 ( .A1(n1216), .A2(n1056), .ZN(n1047) );
XOR2_X1 U905 ( .A(n1168), .B(n1217), .Z(G15) );
XNOR2_X1 U906 ( .A(KEYINPUT22), .B(n1218), .ZN(n1217) );
AND2_X1 U907 ( .A1(n1215), .A2(n1048), .ZN(n1168) );
AND2_X1 U908 ( .A1(n1056), .A2(n1216), .ZN(n1048) );
INV_X1 U909 ( .A(n1195), .ZN(n1216) );
AND4_X1 U910 ( .A1(n1033), .A2(n1046), .A3(n1027), .A4(n1204), .ZN(n1215) );
NOR2_X1 U911 ( .A1(n1043), .A2(n1054), .ZN(n1046) );
INV_X1 U912 ( .A(n1044), .ZN(n1054) );
AND2_X1 U913 ( .A1(n1200), .A2(n1034), .ZN(n1033) );
XNOR2_X1 U914 ( .A(n1072), .B(KEYINPUT49), .ZN(n1200) );
NAND2_X1 U915 ( .A1(n1219), .A2(n1220), .ZN(G12) );
NAND2_X1 U916 ( .A1(n1167), .A2(n1221), .ZN(n1220) );
XOR2_X1 U917 ( .A(KEYINPUT9), .B(n1222), .Z(n1219) );
NOR2_X1 U918 ( .A1(n1167), .A2(n1221), .ZN(n1222) );
AND4_X1 U919 ( .A1(n1042), .A2(n1027), .A3(n1040), .A4(n1223), .ZN(n1167) );
NOR3_X1 U920 ( .A1(n1035), .A2(n1211), .A3(n1034), .ZN(n1223) );
INV_X1 U921 ( .A(n1201), .ZN(n1034) );
XOR2_X1 U922 ( .A(n1075), .B(n1122), .Z(n1201) );
NAND2_X1 U923 ( .A1(G217), .A2(n1224), .ZN(n1122) );
NAND2_X1 U924 ( .A1(n1120), .A2(n1225), .ZN(n1075) );
XNOR2_X1 U925 ( .A(KEYINPUT42), .B(n1226), .ZN(n1225) );
XOR2_X1 U926 ( .A(n1227), .B(n1228), .Z(n1120) );
XOR2_X1 U927 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U928 ( .A(G137), .B(n1198), .ZN(n1230) );
XNOR2_X1 U929 ( .A(KEYINPUT62), .B(n1187), .ZN(n1229) );
XOR2_X1 U930 ( .A(n1231), .B(n1232), .Z(n1227) );
XOR2_X1 U931 ( .A(n1233), .B(n1085), .Z(n1232) );
NAND2_X1 U932 ( .A1(KEYINPUT36), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U933 ( .A(KEYINPUT21), .B(n1221), .ZN(n1234) );
INV_X1 U934 ( .A(G110), .ZN(n1221) );
XOR2_X1 U935 ( .A(n1235), .B(G119), .Z(n1231) );
NAND3_X1 U936 ( .A1(G221), .A2(n1087), .A3(n1236), .ZN(n1235) );
XNOR2_X1 U937 ( .A(G234), .B(KEYINPUT37), .ZN(n1236) );
INV_X1 U938 ( .A(n1204), .ZN(n1211) );
NAND2_X1 U939 ( .A1(n1206), .A2(n1237), .ZN(n1204) );
NAND2_X1 U940 ( .A1(n1208), .A2(n1112), .ZN(n1237) );
INV_X1 U941 ( .A(G898), .ZN(n1112) );
NOR3_X1 U942 ( .A1(n1226), .A2(n1015), .A3(n1087), .ZN(n1208) );
INV_X1 U943 ( .A(n1238), .ZN(n1015) );
NAND3_X1 U944 ( .A1(n1238), .A2(n1087), .A3(G952), .ZN(n1206) );
NAND2_X1 U945 ( .A1(n1239), .A2(G234), .ZN(n1238) );
XNOR2_X1 U946 ( .A(G237), .B(KEYINPUT14), .ZN(n1239) );
INV_X1 U947 ( .A(n1072), .ZN(n1035) );
NOR2_X1 U948 ( .A1(n1070), .A2(n1240), .ZN(n1072) );
AND2_X1 U949 ( .A1(G472), .A2(n1241), .ZN(n1240) );
NAND2_X1 U950 ( .A1(n1242), .A2(n1226), .ZN(n1241) );
XOR2_X1 U951 ( .A(n1243), .B(n1244), .Z(n1242) );
NOR3_X1 U952 ( .A1(G472), .A2(G902), .A3(n1245), .ZN(n1070) );
XNOR2_X1 U953 ( .A(n1243), .B(n1244), .ZN(n1245) );
XNOR2_X1 U954 ( .A(n1246), .B(G101), .ZN(n1244) );
NAND2_X1 U955 ( .A1(KEYINPUT5), .A2(n1141), .ZN(n1246) );
AND3_X1 U956 ( .A1(n1247), .A2(n1087), .A3(G210), .ZN(n1141) );
NOR2_X1 U957 ( .A1(KEYINPUT17), .A2(n1248), .ZN(n1243) );
XOR2_X1 U958 ( .A(n1145), .B(n1146), .Z(n1248) );
XNOR2_X1 U959 ( .A(n1249), .B(n1250), .ZN(n1145) );
XNOR2_X1 U960 ( .A(G119), .B(n1251), .ZN(n1250) );
NAND2_X1 U961 ( .A1(KEYINPUT50), .A2(n1214), .ZN(n1251) );
INV_X1 U962 ( .A(G116), .ZN(n1214) );
XOR2_X1 U963 ( .A(n1252), .B(n1082), .Z(n1249) );
NAND2_X1 U964 ( .A1(KEYINPUT48), .A2(n1218), .ZN(n1252) );
NOR2_X1 U965 ( .A1(n1195), .A2(n1056), .ZN(n1040) );
XOR2_X1 U966 ( .A(n1253), .B(n1254), .Z(n1056) );
XOR2_X1 U967 ( .A(KEYINPUT53), .B(G475), .Z(n1254) );
NAND2_X1 U968 ( .A1(n1134), .A2(n1226), .ZN(n1253) );
XNOR2_X1 U969 ( .A(n1255), .B(n1256), .ZN(n1134) );
NOR2_X1 U970 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U971 ( .A(n1259), .B(KEYINPUT60), .Z(n1258) );
NAND3_X1 U972 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1259) );
OR2_X1 U973 ( .A1(n1187), .A2(n1085), .ZN(n1261) );
NOR2_X1 U974 ( .A1(n1263), .A2(n1262), .ZN(n1257) );
XNOR2_X1 U975 ( .A(G131), .B(n1264), .ZN(n1262) );
NAND2_X1 U976 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND4_X1 U977 ( .A1(G214), .A2(G143), .A3(n1247), .A4(n1087), .ZN(n1266) );
XOR2_X1 U978 ( .A(n1267), .B(KEYINPUT16), .Z(n1265) );
NAND2_X1 U979 ( .A1(n1192), .A2(n1268), .ZN(n1267) );
NAND3_X1 U980 ( .A1(n1247), .A2(n1087), .A3(G214), .ZN(n1268) );
NOR2_X1 U981 ( .A1(n1269), .A2(n1270), .ZN(n1263) );
INV_X1 U982 ( .A(n1260), .ZN(n1270) );
XNOR2_X1 U983 ( .A(n1271), .B(KEYINPUT29), .ZN(n1260) );
NAND2_X1 U984 ( .A1(n1085), .A2(n1187), .ZN(n1271) );
NOR2_X1 U985 ( .A1(n1085), .A2(n1187), .ZN(n1269) );
XNOR2_X1 U986 ( .A(G125), .B(G140), .ZN(n1085) );
NAND2_X1 U987 ( .A1(n1272), .A2(n1273), .ZN(n1255) );
NAND2_X1 U988 ( .A1(G104), .A2(n1274), .ZN(n1273) );
XOR2_X1 U989 ( .A(n1275), .B(KEYINPUT34), .Z(n1272) );
OR2_X1 U990 ( .A1(n1274), .A2(G104), .ZN(n1275) );
XOR2_X1 U991 ( .A(G113), .B(n1276), .Z(n1274) );
XNOR2_X1 U992 ( .A(KEYINPUT52), .B(n1210), .ZN(n1276) );
XNOR2_X1 U993 ( .A(n1050), .B(KEYINPUT18), .ZN(n1195) );
XOR2_X1 U994 ( .A(n1277), .B(G478), .Z(n1050) );
NAND2_X1 U995 ( .A1(n1128), .A2(n1226), .ZN(n1277) );
INV_X1 U996 ( .A(n1131), .ZN(n1128) );
XNOR2_X1 U997 ( .A(n1278), .B(n1279), .ZN(n1131) );
AND4_X1 U998 ( .A1(n1280), .A2(n1087), .A3(G234), .A4(G217), .ZN(n1279) );
INV_X1 U999 ( .A(G953), .ZN(n1087) );
INV_X1 U1000 ( .A(KEYINPUT20), .ZN(n1280) );
NAND2_X1 U1001 ( .A1(n1281), .A2(n1282), .ZN(n1278) );
NAND2_X1 U1002 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U1003 ( .A(n1285), .B(KEYINPUT23), .Z(n1281) );
OR2_X1 U1004 ( .A1(n1284), .A2(n1283), .ZN(n1285) );
XOR2_X1 U1005 ( .A(n1286), .B(n1287), .Z(n1283) );
NOR2_X1 U1006 ( .A1(G122), .A2(KEYINPUT33), .ZN(n1287) );
XNOR2_X1 U1007 ( .A(G107), .B(G116), .ZN(n1286) );
XNOR2_X1 U1008 ( .A(n1288), .B(n1289), .ZN(n1284) );
NOR2_X1 U1009 ( .A1(KEYINPUT10), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U1010 ( .A(KEYINPUT46), .B(n1192), .ZN(n1290) );
INV_X1 U1011 ( .A(G143), .ZN(n1192) );
XNOR2_X1 U1012 ( .A(G134), .B(G128), .ZN(n1288) );
NOR2_X1 U1013 ( .A1(n1291), .A2(n1055), .ZN(n1027) );
INV_X1 U1014 ( .A(n1029), .ZN(n1055) );
NAND2_X1 U1015 ( .A1(G214), .A2(n1292), .ZN(n1029) );
INV_X1 U1016 ( .A(n1028), .ZN(n1291) );
XOR2_X1 U1017 ( .A(n1058), .B(n1185), .Z(n1028) );
NAND2_X1 U1018 ( .A1(G210), .A2(n1292), .ZN(n1185) );
NAND2_X1 U1019 ( .A1(n1247), .A2(n1226), .ZN(n1292) );
INV_X1 U1020 ( .A(G237), .ZN(n1247) );
NAND2_X1 U1021 ( .A1(n1293), .A2(n1226), .ZN(n1058) );
XNOR2_X1 U1022 ( .A(n1156), .B(n1294), .ZN(n1293) );
XOR2_X1 U1023 ( .A(n1161), .B(KEYINPUT61), .Z(n1294) );
XNOR2_X1 U1024 ( .A(n1295), .B(n1146), .ZN(n1161) );
XNOR2_X1 U1025 ( .A(n1296), .B(n1297), .ZN(n1146) );
XNOR2_X1 U1026 ( .A(n1298), .B(KEYINPUT2), .ZN(n1297) );
NAND2_X1 U1027 ( .A1(KEYINPUT59), .A2(n1198), .ZN(n1298) );
XNOR2_X1 U1028 ( .A(G125), .B(n1299), .ZN(n1295) );
NOR2_X1 U1029 ( .A1(G953), .A2(n1108), .ZN(n1299) );
INV_X1 U1030 ( .A(G224), .ZN(n1108) );
XOR2_X1 U1031 ( .A(n1113), .B(n1300), .Z(n1156) );
NOR2_X1 U1032 ( .A1(KEYINPUT32), .A2(n1301), .ZN(n1300) );
INV_X1 U1033 ( .A(n1116), .ZN(n1301) );
XNOR2_X1 U1034 ( .A(n1302), .B(n1303), .ZN(n1116) );
XNOR2_X1 U1035 ( .A(G119), .B(n1218), .ZN(n1303) );
INV_X1 U1036 ( .A(G113), .ZN(n1218) );
XOR2_X1 U1037 ( .A(n1304), .B(n1305), .Z(n1302) );
NOR2_X1 U1038 ( .A1(G116), .A2(KEYINPUT15), .ZN(n1305) );
XNOR2_X1 U1039 ( .A(G110), .B(n1210), .ZN(n1113) );
INV_X1 U1040 ( .A(G122), .ZN(n1210) );
AND2_X1 U1041 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1224), .ZN(n1044) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1226), .ZN(n1224) );
XNOR2_X1 U1044 ( .A(n1069), .B(G469), .ZN(n1043) );
NAND2_X1 U1045 ( .A1(n1306), .A2(n1226), .ZN(n1069) );
INV_X1 U1046 ( .A(G902), .ZN(n1226) );
XNOR2_X1 U1047 ( .A(n1307), .B(n1308), .ZN(n1306) );
INV_X1 U1048 ( .A(n1150), .ZN(n1308) );
XNOR2_X1 U1049 ( .A(n1309), .B(n1310), .ZN(n1150) );
XOR2_X1 U1050 ( .A(n1086), .B(n1311), .Z(n1310) );
NOR2_X1 U1051 ( .A1(G953), .A2(n1092), .ZN(n1311) );
INV_X1 U1052 ( .A(G227), .ZN(n1092) );
AND2_X1 U1053 ( .A1(n1312), .A2(n1313), .ZN(n1086) );
NAND2_X1 U1054 ( .A1(n1314), .A2(n1296), .ZN(n1313) );
XNOR2_X1 U1055 ( .A(KEYINPUT8), .B(G128), .ZN(n1314) );
XOR2_X1 U1056 ( .A(n1315), .B(KEYINPUT6), .Z(n1312) );
NAND2_X1 U1057 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XNOR2_X1 U1058 ( .A(KEYINPUT8), .B(n1198), .ZN(n1317) );
INV_X1 U1059 ( .A(G128), .ZN(n1198) );
XNOR2_X1 U1060 ( .A(n1296), .B(KEYINPUT28), .ZN(n1316) );
XNOR2_X1 U1061 ( .A(G143), .B(n1187), .ZN(n1296) );
INV_X1 U1062 ( .A(G146), .ZN(n1187) );
XOR2_X1 U1063 ( .A(n1304), .B(n1082), .Z(n1309) );
XNOR2_X1 U1064 ( .A(n1318), .B(n1319), .ZN(n1082) );
XNOR2_X1 U1065 ( .A(G137), .B(n1320), .ZN(n1319) );
INV_X1 U1066 ( .A(G134), .ZN(n1320) );
INV_X1 U1067 ( .A(G131), .ZN(n1318) );
XNOR2_X1 U1068 ( .A(G101), .B(n1321), .ZN(n1304) );
XNOR2_X1 U1069 ( .A(n1322), .B(G104), .ZN(n1321) );
INV_X1 U1070 ( .A(G107), .ZN(n1322) );
NAND2_X1 U1071 ( .A1(KEYINPUT45), .A2(n1151), .ZN(n1307) );
XNOR2_X1 U1072 ( .A(G140), .B(G110), .ZN(n1151) );
endmodule


