//Key = 0100101111011111100100001001111000101101100001001000110110110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376;

XNOR2_X1 U754 ( .A(G107), .B(n1046), .ZN(G9) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1049), .A2(n1050), .A3(G953), .A4(n1051), .ZN(n1048) );
NOR2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR3_X1 U759 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NOR2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U761 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR3_X1 U762 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
AND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1061) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1057) );
NOR3_X1 U768 ( .A1(n1071), .A2(n1076), .A3(n1063), .ZN(n1075) );
NOR2_X1 U769 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR4_X1 U770 ( .A1(n1079), .A2(n1063), .A3(n1059), .A4(n1071), .ZN(n1054) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR3_X1 U772 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1047) );
AND4_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1051) );
NOR4_X1 U774 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1085) );
XNOR2_X1 U775 ( .A(G472), .B(n1090), .ZN(n1089) );
XOR2_X1 U776 ( .A(n1091), .B(n1092), .Z(n1087) );
NOR2_X1 U777 ( .A1(KEYINPUT22), .A2(n1093), .ZN(n1092) );
XOR2_X1 U778 ( .A(KEYINPUT21), .B(G469), .Z(n1093) );
XOR2_X1 U779 ( .A(n1094), .B(KEYINPUT19), .Z(n1086) );
NOR3_X1 U780 ( .A1(n1095), .A2(n1096), .A3(n1067), .ZN(n1084) );
NAND2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1083) );
XOR2_X1 U782 ( .A(n1099), .B(KEYINPUT52), .Z(n1097) );
XOR2_X1 U783 ( .A(n1100), .B(n1101), .Z(n1082) );
XOR2_X1 U784 ( .A(KEYINPUT7), .B(n1102), .Z(n1101) );
NOR2_X1 U785 ( .A1(KEYINPUT44), .A2(n1103), .ZN(n1100) );
NAND2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(G72) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U789 ( .A1(G953), .A2(n1110), .ZN(n1109) );
INV_X1 U790 ( .A(n1111), .ZN(n1108) );
INV_X1 U791 ( .A(n1112), .ZN(n1106) );
NAND2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1104) );
NAND2_X1 U793 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1114) );
XOR2_X1 U795 ( .A(n1115), .B(n1116), .Z(n1112) );
NOR2_X1 U796 ( .A1(n1111), .A2(n1117), .ZN(n1116) );
XOR2_X1 U797 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U798 ( .A(G131), .B(n1120), .Z(n1119) );
XOR2_X1 U799 ( .A(G137), .B(G134), .Z(n1120) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(n1118) );
NAND2_X1 U801 ( .A1(KEYINPUT40), .A2(n1123), .ZN(n1121) );
NAND2_X1 U802 ( .A1(KEYINPUT12), .A2(n1124), .ZN(n1115) );
NAND2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U804 ( .A(n1127), .B(n1128), .Z(G69) );
XOR2_X1 U805 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR3_X1 U806 ( .A1(n1131), .A2(KEYINPUT5), .A3(G953), .ZN(n1130) );
NAND2_X1 U807 ( .A1(n1132), .A2(n1133), .ZN(n1129) );
INV_X1 U808 ( .A(n1134), .ZN(n1133) );
NAND2_X1 U809 ( .A1(G953), .A2(n1135), .ZN(n1127) );
NAND2_X1 U810 ( .A1(G898), .A2(G224), .ZN(n1135) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(G66) );
NOR3_X1 U812 ( .A1(n1102), .A2(n1138), .A3(n1139), .ZN(n1137) );
AND3_X1 U813 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
NOR2_X1 U814 ( .A1(n1143), .A2(n1140), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1144), .A2(n1103), .ZN(n1143) );
NOR2_X1 U816 ( .A1(n1125), .A2(n1145), .ZN(n1144) );
NOR2_X1 U817 ( .A1(n1136), .A2(n1146), .ZN(G63) );
XNOR2_X1 U818 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U819 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XNOR2_X1 U820 ( .A(G478), .B(KEYINPUT25), .ZN(n1149) );
NOR2_X1 U821 ( .A1(n1136), .A2(n1151), .ZN(G60) );
XOR2_X1 U822 ( .A(n1152), .B(n1153), .Z(n1151) );
AND2_X1 U823 ( .A1(G475), .A2(n1142), .ZN(n1153) );
NAND2_X1 U824 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
INV_X1 U825 ( .A(n1156), .ZN(n1155) );
XNOR2_X1 U826 ( .A(KEYINPUT41), .B(KEYINPUT23), .ZN(n1154) );
XOR2_X1 U827 ( .A(n1157), .B(n1158), .Z(G6) );
NOR2_X1 U828 ( .A1(n1159), .A2(n1160), .ZN(G57) );
XOR2_X1 U829 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U830 ( .A(n1163), .B(n1164), .ZN(n1161) );
NAND3_X1 U831 ( .A1(n1142), .A2(G472), .A3(KEYINPUT34), .ZN(n1163) );
NOR2_X1 U832 ( .A1(n1165), .A2(n1126), .ZN(n1159) );
XNOR2_X1 U833 ( .A(G952), .B(KEYINPUT28), .ZN(n1165) );
NOR2_X1 U834 ( .A1(n1136), .A2(n1166), .ZN(G54) );
XOR2_X1 U835 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U836 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U837 ( .A(n1171), .B(KEYINPUT62), .ZN(n1170) );
NAND2_X1 U838 ( .A1(n1172), .A2(n1173), .ZN(n1169) );
OR2_X1 U839 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U840 ( .A(n1176), .B(KEYINPUT46), .Z(n1172) );
NAND2_X1 U841 ( .A1(n1175), .A2(n1174), .ZN(n1176) );
XNOR2_X1 U842 ( .A(n1177), .B(n1178), .ZN(n1174) );
XOR2_X1 U843 ( .A(n1179), .B(G101), .Z(n1177) );
NAND2_X1 U844 ( .A1(KEYINPUT16), .A2(n1180), .ZN(n1179) );
XNOR2_X1 U845 ( .A(n1181), .B(n1182), .ZN(n1167) );
AND2_X1 U846 ( .A1(G469), .A2(n1142), .ZN(n1182) );
INV_X1 U847 ( .A(n1150), .ZN(n1142) );
NOR2_X1 U848 ( .A1(n1136), .A2(n1183), .ZN(G51) );
XOR2_X1 U849 ( .A(n1184), .B(n1185), .Z(n1183) );
XNOR2_X1 U850 ( .A(n1186), .B(n1187), .ZN(n1184) );
NOR2_X1 U851 ( .A1(n1098), .A2(n1150), .ZN(n1187) );
NAND2_X1 U852 ( .A1(G902), .A2(n1049), .ZN(n1150) );
NAND2_X1 U853 ( .A1(n1131), .A2(n1188), .ZN(n1049) );
INV_X1 U854 ( .A(n1125), .ZN(n1188) );
NAND4_X1 U855 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1125) );
AND4_X1 U856 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
AND2_X1 U857 ( .A1(n1197), .A2(n1198), .ZN(n1191) );
NAND2_X1 U858 ( .A1(n1199), .A2(n1081), .ZN(n1189) );
INV_X1 U859 ( .A(n1145), .ZN(n1131) );
NAND2_X1 U860 ( .A1(n1200), .A2(n1201), .ZN(n1145) );
AND4_X1 U861 ( .A1(n1046), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1201) );
NAND3_X1 U862 ( .A1(n1080), .A2(n1068), .A3(n1205), .ZN(n1046) );
AND4_X1 U863 ( .A1(n1206), .A2(n1207), .A3(n1158), .A4(n1208), .ZN(n1200) );
NAND2_X1 U864 ( .A1(n1065), .A2(n1209), .ZN(n1208) );
INV_X1 U865 ( .A(n1210), .ZN(n1209) );
NAND3_X1 U866 ( .A1(n1205), .A2(n1068), .A3(n1081), .ZN(n1158) );
NOR2_X1 U867 ( .A1(n1126), .A2(G952), .ZN(n1136) );
XOR2_X1 U868 ( .A(n1211), .B(n1212), .Z(G48) );
NAND3_X1 U869 ( .A1(n1199), .A2(n1081), .A3(KEYINPUT24), .ZN(n1212) );
XNOR2_X1 U870 ( .A(G143), .B(n1190), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1065), .A2(n1213), .A3(n1214), .A4(n1088), .ZN(n1190) );
NAND3_X1 U872 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(G42) );
NAND2_X1 U873 ( .A1(G140), .A2(n1198), .ZN(n1217) );
NAND2_X1 U874 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
INV_X1 U875 ( .A(KEYINPUT15), .ZN(n1219) );
NAND2_X1 U876 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
INV_X1 U877 ( .A(n1198), .ZN(n1221) );
XNOR2_X1 U878 ( .A(KEYINPUT49), .B(G140), .ZN(n1220) );
NAND2_X1 U879 ( .A1(KEYINPUT15), .A2(n1222), .ZN(n1215) );
NAND2_X1 U880 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
OR3_X1 U881 ( .A1(n1198), .A2(G140), .A3(KEYINPUT49), .ZN(n1224) );
NAND4_X1 U882 ( .A1(n1225), .A2(n1226), .A3(n1081), .A4(n1073), .ZN(n1198) );
NAND2_X1 U883 ( .A1(KEYINPUT49), .A2(G140), .ZN(n1223) );
XOR2_X1 U884 ( .A(n1227), .B(n1197), .Z(G39) );
NAND4_X1 U885 ( .A1(n1225), .A2(n1226), .A3(n1228), .A4(n1229), .ZN(n1197) );
XNOR2_X1 U886 ( .A(G134), .B(n1196), .ZN(G36) );
NAND3_X1 U887 ( .A1(n1225), .A2(n1080), .A3(n1213), .ZN(n1196) );
XOR2_X1 U888 ( .A(G131), .B(n1230), .Z(G33) );
NOR2_X1 U889 ( .A1(KEYINPUT50), .A2(n1195), .ZN(n1230) );
NAND3_X1 U890 ( .A1(n1225), .A2(n1081), .A3(n1213), .ZN(n1195) );
AND4_X1 U891 ( .A1(n1072), .A2(n1228), .A3(n1231), .A4(n1232), .ZN(n1213) );
INV_X1 U892 ( .A(n1071), .ZN(n1225) );
NAND2_X1 U893 ( .A1(n1066), .A2(n1233), .ZN(n1071) );
XNOR2_X1 U894 ( .A(G128), .B(n1194), .ZN(G30) );
NAND2_X1 U895 ( .A1(n1199), .A2(n1080), .ZN(n1194) );
AND3_X1 U896 ( .A1(n1065), .A2(n1228), .A3(n1226), .ZN(n1199) );
AND3_X1 U897 ( .A1(n1234), .A2(n1232), .A3(n1231), .ZN(n1226) );
XOR2_X1 U898 ( .A(n1235), .B(n1207), .Z(G3) );
NAND4_X1 U899 ( .A1(n1228), .A2(n1229), .A3(n1072), .A4(n1205), .ZN(n1207) );
XOR2_X1 U900 ( .A(n1123), .B(n1193), .Z(G27) );
NAND4_X1 U901 ( .A1(n1081), .A2(n1074), .A3(n1065), .A4(n1236), .ZN(n1193) );
AND3_X1 U902 ( .A1(n1073), .A2(n1232), .A3(n1234), .ZN(n1236) );
NAND2_X1 U903 ( .A1(n1053), .A2(n1237), .ZN(n1232) );
NAND3_X1 U904 ( .A1(G902), .A2(n1238), .A3(n1111), .ZN(n1237) );
NOR2_X1 U905 ( .A1(n1126), .A2(G900), .ZN(n1111) );
NAND2_X1 U906 ( .A1(n1239), .A2(n1240), .ZN(G24) );
OR2_X1 U907 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U908 ( .A(n1243), .B(KEYINPUT63), .Z(n1239) );
NAND2_X1 U909 ( .A1(n1242), .A2(n1241), .ZN(n1243) );
NOR2_X1 U910 ( .A1(n1210), .A2(n1244), .ZN(n1242) );
XOR2_X1 U911 ( .A(KEYINPUT6), .B(n1065), .Z(n1244) );
NAND3_X1 U912 ( .A1(n1074), .A2(n1068), .A3(n1245), .ZN(n1210) );
NOR3_X1 U913 ( .A1(n1094), .A2(n1246), .A3(n1247), .ZN(n1245) );
INV_X1 U914 ( .A(n1063), .ZN(n1068) );
NAND2_X1 U915 ( .A1(n1072), .A2(n1073), .ZN(n1063) );
INV_X1 U916 ( .A(n1059), .ZN(n1074) );
XOR2_X1 U917 ( .A(n1248), .B(n1206), .Z(G21) );
NAND4_X1 U918 ( .A1(n1065), .A2(n1249), .A3(n1229), .A4(n1234), .ZN(n1206) );
XOR2_X1 U919 ( .A(n1250), .B(n1204), .Z(G18) );
NAND4_X1 U920 ( .A1(n1065), .A2(n1249), .A3(n1072), .A4(n1080), .ZN(n1204) );
NOR2_X1 U921 ( .A1(n1214), .A2(n1247), .ZN(n1080) );
INV_X1 U922 ( .A(n1094), .ZN(n1214) );
XNOR2_X1 U923 ( .A(n1251), .B(KEYINPUT58), .ZN(n1065) );
XNOR2_X1 U924 ( .A(G113), .B(n1203), .ZN(G15) );
NAND4_X1 U925 ( .A1(n1081), .A2(n1249), .A3(n1072), .A4(n1251), .ZN(n1203) );
NOR3_X1 U926 ( .A1(n1073), .A2(n1246), .A3(n1059), .ZN(n1249) );
NAND2_X1 U927 ( .A1(n1077), .A2(n1078), .ZN(n1059) );
INV_X1 U928 ( .A(n1252), .ZN(n1246) );
NOR2_X1 U929 ( .A1(n1088), .A2(n1094), .ZN(n1081) );
INV_X1 U930 ( .A(n1247), .ZN(n1088) );
NAND3_X1 U931 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(G12) );
NAND2_X1 U932 ( .A1(G110), .A2(n1202), .ZN(n1255) );
NAND2_X1 U933 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
INV_X1 U934 ( .A(KEYINPUT30), .ZN(n1257) );
NAND2_X1 U935 ( .A1(n1258), .A2(n1259), .ZN(n1256) );
XNOR2_X1 U936 ( .A(KEYINPUT18), .B(n1202), .ZN(n1258) );
NAND2_X1 U937 ( .A1(KEYINPUT30), .A2(n1260), .ZN(n1253) );
NAND2_X1 U938 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NAND2_X1 U939 ( .A1(KEYINPUT18), .A2(n1202), .ZN(n1262) );
OR3_X1 U940 ( .A1(G110), .A2(KEYINPUT18), .A3(n1202), .ZN(n1261) );
NAND4_X1 U941 ( .A1(n1229), .A2(n1205), .A3(n1073), .A4(n1234), .ZN(n1202) );
INV_X1 U942 ( .A(n1072), .ZN(n1234) );
XOR2_X1 U943 ( .A(n1263), .B(n1102), .Z(n1072) );
NOR2_X1 U944 ( .A1(n1140), .A2(G902), .ZN(n1102) );
XOR2_X1 U945 ( .A(n1264), .B(n1265), .Z(n1140) );
XOR2_X1 U946 ( .A(G137), .B(n1266), .Z(n1265) );
NOR2_X1 U947 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
INV_X1 U948 ( .A(G221), .ZN(n1267) );
NAND2_X1 U949 ( .A1(n1269), .A2(KEYINPUT61), .ZN(n1264) );
XOR2_X1 U950 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U951 ( .A(n1272), .B(n1181), .Z(n1271) );
XNOR2_X1 U952 ( .A(n1259), .B(G140), .ZN(n1181) );
INV_X1 U953 ( .A(G110), .ZN(n1259) );
NOR2_X1 U954 ( .A1(KEYINPUT31), .A2(n1211), .ZN(n1272) );
XOR2_X1 U955 ( .A(n1273), .B(n1274), .Z(n1270) );
XOR2_X1 U956 ( .A(KEYINPUT43), .B(G125), .Z(n1274) );
NAND2_X1 U957 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND2_X1 U958 ( .A1(G128), .A2(n1248), .ZN(n1276) );
XOR2_X1 U959 ( .A(KEYINPUT53), .B(n1277), .Z(n1275) );
NOR2_X1 U960 ( .A1(G128), .A2(n1248), .ZN(n1277) );
NAND2_X1 U961 ( .A1(KEYINPUT14), .A2(n1141), .ZN(n1263) );
INV_X1 U962 ( .A(n1103), .ZN(n1141) );
NAND2_X1 U963 ( .A1(G217), .A2(n1278), .ZN(n1103) );
INV_X1 U964 ( .A(n1228), .ZN(n1073) );
XOR2_X1 U965 ( .A(n1090), .B(n1279), .Z(n1228) );
NOR2_X1 U966 ( .A1(KEYINPUT2), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U967 ( .A(G472), .B(KEYINPUT36), .ZN(n1280) );
NAND2_X1 U968 ( .A1(n1281), .A2(n1282), .ZN(n1090) );
XOR2_X1 U969 ( .A(n1283), .B(n1162), .Z(n1281) );
XOR2_X1 U970 ( .A(n1284), .B(n1285), .Z(n1162) );
XOR2_X1 U971 ( .A(n1286), .B(n1235), .Z(n1285) );
INV_X1 U972 ( .A(G101), .ZN(n1235) );
NAND2_X1 U973 ( .A1(n1287), .A2(G210), .ZN(n1286) );
XOR2_X1 U974 ( .A(n1175), .B(n1288), .Z(n1284) );
NOR2_X1 U975 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U976 ( .A(KEYINPUT0), .B(n1291), .Z(n1290) );
AND2_X1 U977 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NOR2_X1 U978 ( .A1(n1293), .A2(n1292), .ZN(n1289) );
XOR2_X1 U979 ( .A(G113), .B(KEYINPUT45), .Z(n1292) );
XNOR2_X1 U980 ( .A(KEYINPUT29), .B(n1294), .ZN(n1283) );
NOR2_X1 U981 ( .A1(KEYINPUT60), .A2(n1164), .ZN(n1294) );
AND3_X1 U982 ( .A1(n1251), .A2(n1252), .A3(n1231), .ZN(n1205) );
NOR2_X1 U983 ( .A1(n1077), .A2(n1095), .ZN(n1231) );
INV_X1 U984 ( .A(n1078), .ZN(n1095) );
NAND2_X1 U985 ( .A1(G221), .A2(n1278), .ZN(n1078) );
NAND2_X1 U986 ( .A1(G234), .A2(n1282), .ZN(n1278) );
XOR2_X1 U987 ( .A(n1091), .B(G469), .Z(n1077) );
NAND2_X1 U988 ( .A1(n1295), .A2(n1282), .ZN(n1091) );
XOR2_X1 U989 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U990 ( .A(n1298), .B(n1299), .Z(n1297) );
XNOR2_X1 U991 ( .A(n1300), .B(n1301), .ZN(n1299) );
NOR2_X1 U992 ( .A1(KEYINPUT42), .A2(n1175), .ZN(n1301) );
AND2_X1 U993 ( .A1(n1302), .A2(n1303), .ZN(n1175) );
NAND2_X1 U994 ( .A1(n1304), .A2(G137), .ZN(n1303) );
NAND2_X1 U995 ( .A1(n1305), .A2(n1227), .ZN(n1302) );
INV_X1 U996 ( .A(G137), .ZN(n1227) );
XNOR2_X1 U997 ( .A(n1304), .B(KEYINPUT10), .ZN(n1305) );
XNOR2_X1 U998 ( .A(n1306), .B(G134), .ZN(n1304) );
NAND2_X1 U999 ( .A1(KEYINPUT27), .A2(n1307), .ZN(n1306) );
INV_X1 U1000 ( .A(G131), .ZN(n1307) );
NAND2_X1 U1001 ( .A1(KEYINPUT1), .A2(n1171), .ZN(n1300) );
NOR2_X1 U1002 ( .A1(n1110), .A2(G953), .ZN(n1171) );
INV_X1 U1003 ( .A(G227), .ZN(n1110) );
XNOR2_X1 U1004 ( .A(n1122), .B(n1178), .ZN(n1296) );
XOR2_X1 U1005 ( .A(G104), .B(n1308), .Z(n1178) );
XOR2_X1 U1006 ( .A(G140), .B(n1180), .Z(n1122) );
XNOR2_X1 U1007 ( .A(n1309), .B(n1310), .ZN(n1180) );
XOR2_X1 U1008 ( .A(n1211), .B(KEYINPUT32), .Z(n1309) );
NAND2_X1 U1009 ( .A1(n1311), .A2(n1312), .ZN(n1252) );
NAND3_X1 U1010 ( .A1(n1134), .A2(n1238), .A3(G902), .ZN(n1312) );
NOR2_X1 U1011 ( .A1(n1126), .A2(G898), .ZN(n1134) );
XOR2_X1 U1012 ( .A(n1053), .B(KEYINPUT38), .Z(n1311) );
NAND3_X1 U1013 ( .A1(n1238), .A2(n1126), .A3(G952), .ZN(n1053) );
NAND2_X1 U1014 ( .A1(G237), .A2(G234), .ZN(n1238) );
NOR2_X1 U1015 ( .A1(n1066), .A2(n1067), .ZN(n1251) );
INV_X1 U1016 ( .A(n1233), .ZN(n1067) );
NAND2_X1 U1017 ( .A1(G214), .A2(n1313), .ZN(n1233) );
NOR2_X1 U1018 ( .A1(n1314), .A2(n1096), .ZN(n1066) );
NOR2_X1 U1019 ( .A1(n1098), .A2(n1315), .ZN(n1096) );
AND2_X1 U1020 ( .A1(n1316), .A2(n1098), .ZN(n1314) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1313), .ZN(n1098) );
NAND2_X1 U1022 ( .A1(n1317), .A2(n1282), .ZN(n1313) );
XOR2_X1 U1023 ( .A(KEYINPUT37), .B(G237), .Z(n1317) );
XNOR2_X1 U1024 ( .A(n1315), .B(KEYINPUT55), .ZN(n1316) );
INV_X1 U1025 ( .A(n1099), .ZN(n1315) );
NAND2_X1 U1026 ( .A1(n1318), .A2(n1282), .ZN(n1099) );
XOR2_X1 U1027 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1028 ( .A(n1185), .B(KEYINPUT4), .ZN(n1320) );
XOR2_X1 U1029 ( .A(n1132), .B(n1321), .Z(n1185) );
AND2_X1 U1030 ( .A1(n1126), .A2(G224), .ZN(n1321) );
XNOR2_X1 U1031 ( .A(n1322), .B(n1323), .ZN(n1132) );
XOR2_X1 U1032 ( .A(n1241), .B(n1324), .Z(n1323) );
NAND2_X1 U1033 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1034 ( .A1(n1327), .A2(n1293), .ZN(n1326) );
XOR2_X1 U1035 ( .A(KEYINPUT56), .B(n1328), .Z(n1325) );
NOR2_X1 U1036 ( .A1(n1293), .A2(n1327), .ZN(n1328) );
XNOR2_X1 U1037 ( .A(KEYINPUT17), .B(G113), .ZN(n1327) );
XOR2_X1 U1038 ( .A(G116), .B(n1248), .Z(n1293) );
INV_X1 U1039 ( .A(G119), .ZN(n1248) );
INV_X1 U1040 ( .A(G122), .ZN(n1241) );
XOR2_X1 U1041 ( .A(n1329), .B(n1298), .Z(n1322) );
XOR2_X1 U1042 ( .A(G101), .B(G110), .Z(n1298) );
NAND2_X1 U1043 ( .A1(n1330), .A2(KEYINPUT8), .ZN(n1329) );
XOR2_X1 U1044 ( .A(n1157), .B(n1331), .Z(n1330) );
NOR2_X1 U1045 ( .A1(KEYINPUT57), .A2(n1308), .ZN(n1331) );
INV_X1 U1046 ( .A(G104), .ZN(n1157) );
NAND2_X1 U1047 ( .A1(n1332), .A2(n1333), .ZN(n1319) );
OR3_X1 U1048 ( .A1(n1123), .A2(n1164), .A3(KEYINPUT59), .ZN(n1333) );
NAND2_X1 U1049 ( .A1(n1186), .A2(KEYINPUT59), .ZN(n1332) );
XOR2_X1 U1050 ( .A(n1123), .B(n1164), .Z(n1186) );
XOR2_X1 U1051 ( .A(n1334), .B(n1335), .Z(n1164) );
XOR2_X1 U1052 ( .A(KEYINPUT20), .B(G128), .Z(n1335) );
NAND2_X1 U1053 ( .A1(n1336), .A2(n1337), .ZN(n1334) );
OR2_X1 U1054 ( .A1(n1211), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1055 ( .A(n1339), .B(KEYINPUT3), .Z(n1336) );
NAND2_X1 U1056 ( .A1(n1338), .A2(n1211), .ZN(n1339) );
INV_X1 U1057 ( .A(n1056), .ZN(n1229) );
NAND2_X1 U1058 ( .A1(n1340), .A2(n1247), .ZN(n1056) );
XOR2_X1 U1059 ( .A(n1341), .B(G478), .Z(n1247) );
NAND2_X1 U1060 ( .A1(n1147), .A2(n1282), .ZN(n1341) );
INV_X1 U1061 ( .A(G902), .ZN(n1282) );
XNOR2_X1 U1062 ( .A(n1342), .B(n1343), .ZN(n1147) );
XOR2_X1 U1063 ( .A(n1344), .B(n1310), .Z(n1343) );
XOR2_X1 U1064 ( .A(G128), .B(n1338), .Z(n1310) );
NOR2_X1 U1065 ( .A1(n1268), .A2(n1345), .ZN(n1344) );
INV_X1 U1066 ( .A(G217), .ZN(n1345) );
NAND2_X1 U1067 ( .A1(n1346), .A2(n1126), .ZN(n1268) );
INV_X1 U1068 ( .A(G953), .ZN(n1126) );
XNOR2_X1 U1069 ( .A(G234), .B(KEYINPUT48), .ZN(n1346) );
XOR2_X1 U1070 ( .A(n1347), .B(G134), .Z(n1342) );
NAND3_X1 U1071 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1347) );
NAND2_X1 U1072 ( .A1(KEYINPUT47), .A2(n1351), .ZN(n1350) );
OR3_X1 U1073 ( .A1(n1351), .A2(KEYINPUT47), .A3(n1308), .ZN(n1349) );
NAND2_X1 U1074 ( .A1(n1308), .A2(n1352), .ZN(n1348) );
NAND2_X1 U1075 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
INV_X1 U1076 ( .A(KEYINPUT47), .ZN(n1354) );
XNOR2_X1 U1077 ( .A(n1351), .B(KEYINPUT26), .ZN(n1353) );
XNOR2_X1 U1078 ( .A(n1355), .B(G122), .ZN(n1351) );
NAND2_X1 U1079 ( .A1(KEYINPUT13), .A2(n1250), .ZN(n1355) );
INV_X1 U1080 ( .A(G116), .ZN(n1250) );
XOR2_X1 U1081 ( .A(G107), .B(KEYINPUT11), .Z(n1308) );
XOR2_X1 U1082 ( .A(n1094), .B(KEYINPUT54), .Z(n1340) );
XNOR2_X1 U1083 ( .A(G475), .B(n1356), .ZN(n1094) );
NOR2_X1 U1084 ( .A1(G902), .A2(n1156), .ZN(n1356) );
NAND3_X1 U1085 ( .A1(n1357), .A2(n1358), .A3(n1359), .ZN(n1156) );
NAND2_X1 U1086 ( .A1(KEYINPUT33), .A2(n1360), .ZN(n1359) );
NAND3_X1 U1087 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1358) );
INV_X1 U1088 ( .A(KEYINPUT33), .ZN(n1362) );
OR2_X1 U1089 ( .A1(n1363), .A2(n1361), .ZN(n1357) );
NOR2_X1 U1090 ( .A1(KEYINPUT35), .A2(n1360), .ZN(n1361) );
XOR2_X1 U1091 ( .A(G104), .B(n1364), .Z(n1360) );
XOR2_X1 U1092 ( .A(G122), .B(G113), .Z(n1364) );
XNOR2_X1 U1093 ( .A(n1365), .B(n1366), .ZN(n1363) );
XNOR2_X1 U1094 ( .A(n1367), .B(n1338), .ZN(n1366) );
XOR2_X1 U1095 ( .A(G143), .B(KEYINPUT51), .Z(n1338) );
NAND2_X1 U1096 ( .A1(n1287), .A2(G214), .ZN(n1367) );
NOR2_X1 U1097 ( .A1(G953), .A2(G237), .ZN(n1287) );
XOR2_X1 U1098 ( .A(n1368), .B(G131), .Z(n1365) );
NAND2_X1 U1099 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
NAND2_X1 U1100 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
NAND2_X1 U1101 ( .A1(KEYINPUT9), .A2(n1373), .ZN(n1372) );
NAND2_X1 U1102 ( .A1(KEYINPUT39), .A2(G146), .ZN(n1373) );
NAND2_X1 U1103 ( .A1(n1374), .A2(n1211), .ZN(n1369) );
INV_X1 U1104 ( .A(G146), .ZN(n1211) );
NAND2_X1 U1105 ( .A1(KEYINPUT39), .A2(n1375), .ZN(n1374) );
NAND2_X1 U1106 ( .A1(KEYINPUT9), .A2(n1376), .ZN(n1375) );
INV_X1 U1107 ( .A(n1371), .ZN(n1376) );
XOR2_X1 U1108 ( .A(n1123), .B(G140), .Z(n1371) );
INV_X1 U1109 ( .A(G125), .ZN(n1123) );
endmodule


