//Key = 1011100000001101101011011111000010000101110111111011101110110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375;

NAND3_X1 U762 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(G9) );
OR2_X1 U763 ( .A1(n1052), .A2(G107), .ZN(n1051) );
NAND2_X1 U764 ( .A1(KEYINPUT5), .A2(n1053), .ZN(n1050) );
NAND2_X1 U765 ( .A1(G107), .A2(n1054), .ZN(n1053) );
XNOR2_X1 U766 ( .A(KEYINPUT52), .B(n1052), .ZN(n1054) );
NAND2_X1 U767 ( .A1(n1055), .A2(n1056), .ZN(n1049) );
INV_X1 U768 ( .A(KEYINPUT5), .ZN(n1056) );
NAND2_X1 U769 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND3_X1 U770 ( .A1(KEYINPUT52), .A2(G107), .A3(n1052), .ZN(n1058) );
OR2_X1 U771 ( .A1(n1052), .A2(KEYINPUT52), .ZN(n1057) );
NOR2_X1 U772 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR4_X1 U773 ( .A1(G953), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1060) );
NOR2_X1 U774 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U775 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR3_X1 U776 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NOR2_X1 U777 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U778 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U779 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR2_X1 U780 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U781 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR2_X1 U782 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR2_X1 U783 ( .A1(n1083), .A2(n1084), .ZN(n1075) );
NOR2_X1 U784 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR2_X1 U785 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR3_X1 U786 ( .A1(n1084), .A2(n1089), .A3(n1078), .ZN(n1071) );
NOR2_X1 U787 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR3_X1 U788 ( .A1(n1084), .A2(n1092), .A3(n1078), .ZN(n1066) );
INV_X1 U789 ( .A(n1093), .ZN(n1078) );
NOR2_X1 U790 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR3_X1 U791 ( .A1(n1096), .A2(n1074), .A3(n1068), .ZN(n1094) );
INV_X1 U792 ( .A(n1097), .ZN(n1074) );
NOR3_X1 U793 ( .A1(n1061), .A2(G953), .A3(G952), .ZN(n1059) );
AND4_X1 U794 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1061) );
NOR4_X1 U795 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1101) );
NAND3_X1 U796 ( .A1(n1096), .A2(n1106), .A3(n1082), .ZN(n1102) );
NOR3_X1 U797 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1100) );
AND2_X1 U798 ( .A1(n1110), .A2(G472), .ZN(n1109) );
XOR2_X1 U799 ( .A(n1111), .B(KEYINPUT60), .Z(n1107) );
NAND2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U801 ( .A1(G475), .A2(n1114), .ZN(n1113) );
XOR2_X1 U802 ( .A(KEYINPUT12), .B(n1115), .Z(n1112) );
XNOR2_X1 U803 ( .A(KEYINPUT15), .B(n1116), .ZN(n1099) );
XNOR2_X1 U804 ( .A(n1117), .B(KEYINPUT29), .ZN(n1098) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(G72) );
NOR2_X1 U806 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U807 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NAND2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1118) );
NAND2_X1 U809 ( .A1(n1126), .A2(n1121), .ZN(n1125) );
XNOR2_X1 U810 ( .A(n1127), .B(n1128), .ZN(n1126) );
NAND3_X1 U811 ( .A1(G900), .A2(n1128), .A3(G953), .ZN(n1124) );
XNOR2_X1 U812 ( .A(n1129), .B(n1130), .ZN(n1128) );
XNOR2_X1 U813 ( .A(n1131), .B(n1132), .ZN(n1130) );
NAND2_X1 U814 ( .A1(n1133), .A2(KEYINPUT55), .ZN(n1131) );
XNOR2_X1 U815 ( .A(G125), .B(G140), .ZN(n1133) );
XOR2_X1 U816 ( .A(n1134), .B(n1135), .Z(n1129) );
NOR2_X1 U817 ( .A1(KEYINPUT8), .A2(n1136), .ZN(n1135) );
XNOR2_X1 U818 ( .A(KEYINPUT63), .B(n1137), .ZN(n1136) );
XNOR2_X1 U819 ( .A(G131), .B(G137), .ZN(n1134) );
NAND2_X1 U820 ( .A1(n1138), .A2(n1139), .ZN(G69) );
NAND2_X1 U821 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U822 ( .A1(G953), .A2(n1142), .ZN(n1141) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1142) );
NAND2_X1 U824 ( .A1(n1143), .A2(n1144), .ZN(n1138) );
NAND2_X1 U825 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U826 ( .A1(G953), .A2(n1147), .ZN(n1146) );
INV_X1 U827 ( .A(n1140), .ZN(n1143) );
XNOR2_X1 U828 ( .A(n1148), .B(n1149), .ZN(n1140) );
NOR2_X1 U829 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XNOR2_X1 U830 ( .A(G953), .B(KEYINPUT21), .ZN(n1151) );
NAND3_X1 U831 ( .A1(n1152), .A2(n1153), .A3(n1145), .ZN(n1148) );
INV_X1 U832 ( .A(n1154), .ZN(n1145) );
NAND2_X1 U833 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
INV_X1 U834 ( .A(n1157), .ZN(n1156) );
NAND2_X1 U835 ( .A1(n1158), .A2(n1157), .ZN(n1152) );
XNOR2_X1 U836 ( .A(KEYINPUT33), .B(n1155), .ZN(n1158) );
NOR2_X1 U837 ( .A1(n1159), .A2(n1160), .ZN(G66) );
NOR2_X1 U838 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(n1161) );
XOR2_X1 U841 ( .A(KEYINPUT23), .B(n1164), .Z(n1166) );
XNOR2_X1 U842 ( .A(n1163), .B(KEYINPUT17), .ZN(n1165) );
AND2_X1 U843 ( .A1(n1167), .A2(n1168), .ZN(n1163) );
NOR2_X1 U844 ( .A1(n1159), .A2(n1169), .ZN(G63) );
XOR2_X1 U845 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U846 ( .A(n1172), .B(KEYINPUT31), .Z(n1171) );
NAND2_X1 U847 ( .A1(n1167), .A2(G478), .ZN(n1172) );
NOR2_X1 U848 ( .A1(n1159), .A2(n1173), .ZN(G60) );
XOR2_X1 U849 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U850 ( .A1(n1167), .A2(G475), .ZN(n1174) );
XOR2_X1 U851 ( .A(G104), .B(n1176), .Z(G6) );
NOR2_X1 U852 ( .A1(n1159), .A2(n1177), .ZN(G57) );
XOR2_X1 U853 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U854 ( .A(n1180), .B(n1181), .ZN(n1179) );
NAND2_X1 U855 ( .A1(n1182), .A2(KEYINPUT27), .ZN(n1180) );
XOR2_X1 U856 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR3_X1 U857 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NOR2_X1 U858 ( .A1(KEYINPUT39), .A2(n1188), .ZN(n1187) );
NOR2_X1 U859 ( .A1(n1189), .A2(n1063), .ZN(n1188) );
NOR2_X1 U860 ( .A1(n1167), .A2(n1190), .ZN(n1186) );
INV_X1 U861 ( .A(KEYINPUT39), .ZN(n1190) );
INV_X1 U862 ( .A(G472), .ZN(n1185) );
NAND2_X1 U863 ( .A1(n1191), .A2(KEYINPUT4), .ZN(n1183) );
XOR2_X1 U864 ( .A(n1192), .B(n1193), .Z(n1191) );
XNOR2_X1 U865 ( .A(n1194), .B(n1195), .ZN(n1192) );
NOR2_X1 U866 ( .A1(KEYINPUT6), .A2(n1196), .ZN(n1195) );
INV_X1 U867 ( .A(n1197), .ZN(n1196) );
XNOR2_X1 U868 ( .A(G101), .B(KEYINPUT49), .ZN(n1178) );
NOR3_X1 U869 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(G54) );
AND2_X1 U870 ( .A1(KEYINPUT3), .A2(n1159), .ZN(n1200) );
NOR3_X1 U871 ( .A1(KEYINPUT3), .A2(n1121), .A3(n1201), .ZN(n1199) );
INV_X1 U872 ( .A(G952), .ZN(n1201) );
XOR2_X1 U873 ( .A(n1202), .B(n1203), .Z(n1198) );
XOR2_X1 U874 ( .A(n1204), .B(n1205), .Z(n1203) );
NOR2_X1 U875 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XOR2_X1 U876 ( .A(KEYINPUT30), .B(n1208), .Z(n1207) );
NAND2_X1 U877 ( .A1(KEYINPUT20), .A2(n1209), .ZN(n1204) );
XNOR2_X1 U878 ( .A(n1210), .B(n1211), .ZN(n1209) );
NAND2_X1 U879 ( .A1(n1167), .A2(G469), .ZN(n1202) );
NOR2_X1 U880 ( .A1(n1159), .A2(n1212), .ZN(G51) );
NOR2_X1 U881 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U882 ( .A(n1215), .B(KEYINPUT51), .Z(n1214) );
NAND2_X1 U883 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XNOR2_X1 U884 ( .A(n1218), .B(KEYINPUT7), .ZN(n1216) );
NOR2_X1 U885 ( .A1(n1217), .A2(n1219), .ZN(n1213) );
AND2_X1 U886 ( .A1(n1167), .A2(n1220), .ZN(n1217) );
AND2_X1 U887 ( .A1(G902), .A2(n1063), .ZN(n1167) );
NAND2_X1 U888 ( .A1(n1127), .A2(n1150), .ZN(n1063) );
AND4_X1 U889 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1150) );
NOR4_X1 U890 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1176), .ZN(n1224) );
AND4_X1 U891 ( .A1(n1091), .A2(n1093), .A3(n1228), .A4(n1229), .ZN(n1176) );
NOR2_X1 U892 ( .A1(n1230), .A2(n1231), .ZN(n1223) );
INV_X1 U893 ( .A(n1052), .ZN(n1230) );
NAND4_X1 U894 ( .A1(n1090), .A2(n1093), .A3(n1228), .A4(n1229), .ZN(n1052) );
NAND3_X1 U895 ( .A1(n1086), .A2(n1229), .A3(n1095), .ZN(n1221) );
AND4_X1 U896 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1127) );
AND4_X1 U897 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NAND2_X1 U898 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
XOR2_X1 U899 ( .A(n1242), .B(KEYINPUT25), .Z(n1240) );
NAND3_X1 U900 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1232) );
NAND2_X1 U901 ( .A1(n1246), .A2(n1247), .ZN(n1244) );
NAND3_X1 U902 ( .A1(n1248), .A2(n1090), .A3(KEYINPUT11), .ZN(n1246) );
NAND3_X1 U903 ( .A1(n1249), .A2(n1250), .A3(n1080), .ZN(n1243) );
NAND3_X1 U904 ( .A1(n1090), .A2(n1251), .A3(n1248), .ZN(n1250) );
INV_X1 U905 ( .A(KEYINPUT11), .ZN(n1251) );
NAND2_X1 U906 ( .A1(n1091), .A2(n1252), .ZN(n1249) );
XOR2_X1 U907 ( .A(KEYINPUT22), .B(n1248), .Z(n1252) );
NOR2_X1 U908 ( .A1(n1121), .A2(G952), .ZN(n1159) );
XNOR2_X1 U909 ( .A(n1253), .B(n1254), .ZN(G48) );
NOR2_X1 U910 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U911 ( .A(G143), .B(n1257), .Z(G45) );
NOR2_X1 U912 ( .A1(n1258), .A2(n1233), .ZN(n1257) );
NAND3_X1 U913 ( .A1(n1086), .A2(n1245), .A3(n1259), .ZN(n1233) );
NOR3_X1 U914 ( .A1(n1247), .A2(n1260), .A3(n1261), .ZN(n1259) );
XNOR2_X1 U915 ( .A(KEYINPUT38), .B(KEYINPUT16), .ZN(n1258) );
XNOR2_X1 U916 ( .A(G140), .B(n1239), .ZN(G42) );
NAND2_X1 U917 ( .A1(n1262), .A2(n1263), .ZN(n1239) );
XNOR2_X1 U918 ( .A(G137), .B(n1238), .ZN(G39) );
NAND3_X1 U919 ( .A1(n1248), .A2(n1262), .A3(n1097), .ZN(n1238) );
XNOR2_X1 U920 ( .A(G134), .B(n1237), .ZN(G36) );
NAND3_X1 U921 ( .A1(n1262), .A2(n1090), .A3(n1086), .ZN(n1237) );
AND2_X1 U922 ( .A1(n1245), .A2(n1241), .ZN(n1262) );
INV_X1 U923 ( .A(n1084), .ZN(n1241) );
XOR2_X1 U924 ( .A(G131), .B(n1264), .Z(G33) );
NOR2_X1 U925 ( .A1(n1084), .A2(n1242), .ZN(n1264) );
NAND3_X1 U926 ( .A1(n1245), .A2(n1091), .A3(n1086), .ZN(n1242) );
NAND2_X1 U927 ( .A1(n1265), .A2(n1082), .ZN(n1084) );
XOR2_X1 U928 ( .A(G128), .B(n1266), .Z(G30) );
NOR2_X1 U929 ( .A1(n1267), .A2(n1256), .ZN(n1266) );
NAND3_X1 U930 ( .A1(n1245), .A2(n1080), .A3(n1248), .ZN(n1256) );
AND2_X1 U931 ( .A1(n1228), .A2(n1268), .ZN(n1245) );
INV_X1 U932 ( .A(n1090), .ZN(n1267) );
XNOR2_X1 U933 ( .A(n1269), .B(n1270), .ZN(G3) );
NAND2_X1 U934 ( .A1(KEYINPUT26), .A2(n1271), .ZN(n1269) );
NAND4_X1 U935 ( .A1(n1272), .A2(n1095), .A3(n1086), .A4(n1273), .ZN(n1271) );
XNOR2_X1 U936 ( .A(n1080), .B(KEYINPUT59), .ZN(n1272) );
XNOR2_X1 U937 ( .A(G125), .B(n1236), .ZN(G27) );
NAND3_X1 U938 ( .A1(n1274), .A2(n1263), .A3(n1275), .ZN(n1236) );
AND3_X1 U939 ( .A1(n1080), .A2(n1268), .A3(n1096), .ZN(n1275) );
NAND2_X1 U940 ( .A1(n1276), .A2(n1065), .ZN(n1268) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1277), .A4(n1123), .ZN(n1276) );
INV_X1 U942 ( .A(G900), .ZN(n1123) );
NOR3_X1 U943 ( .A1(n1088), .A2(n1087), .A3(n1255), .ZN(n1263) );
INV_X1 U944 ( .A(n1091), .ZN(n1255) );
XOR2_X1 U945 ( .A(n1222), .B(n1278), .Z(G24) );
XOR2_X1 U946 ( .A(KEYINPUT61), .B(G122), .Z(n1278) );
NAND4_X1 U947 ( .A1(n1279), .A2(n1093), .A3(n1117), .A4(n1280), .ZN(n1222) );
NOR2_X1 U948 ( .A1(n1088), .A2(n1281), .ZN(n1093) );
XOR2_X1 U949 ( .A(n1282), .B(n1231), .Z(G21) );
AND3_X1 U950 ( .A1(n1097), .A2(n1248), .A3(n1279), .ZN(n1231) );
NOR2_X1 U951 ( .A1(n1087), .A2(n1283), .ZN(n1248) );
INV_X1 U952 ( .A(n1281), .ZN(n1087) );
NAND2_X1 U953 ( .A1(n1284), .A2(KEYINPUT37), .ZN(n1282) );
XNOR2_X1 U954 ( .A(G119), .B(KEYINPUT1), .ZN(n1284) );
XOR2_X1 U955 ( .A(G116), .B(n1227), .Z(G18) );
AND3_X1 U956 ( .A1(n1086), .A2(n1090), .A3(n1279), .ZN(n1227) );
NOR2_X1 U957 ( .A1(n1280), .A2(n1261), .ZN(n1090) );
INV_X1 U958 ( .A(n1117), .ZN(n1261) );
XOR2_X1 U959 ( .A(G113), .B(n1226), .Z(G15) );
AND3_X1 U960 ( .A1(n1086), .A2(n1091), .A3(n1279), .ZN(n1226) );
AND3_X1 U961 ( .A1(n1229), .A2(n1096), .A3(n1274), .ZN(n1279) );
INV_X1 U962 ( .A(n1068), .ZN(n1274) );
XOR2_X1 U963 ( .A(n1285), .B(KEYINPUT42), .Z(n1068) );
NOR2_X1 U964 ( .A1(n1117), .A2(n1260), .ZN(n1091) );
NOR2_X1 U965 ( .A1(n1281), .A2(n1283), .ZN(n1086) );
XOR2_X1 U966 ( .A(G110), .B(n1225), .Z(G12) );
AND4_X1 U967 ( .A1(n1095), .A2(n1229), .A3(n1283), .A4(n1281), .ZN(n1225) );
NAND2_X1 U968 ( .A1(n1286), .A2(n1106), .ZN(n1281) );
NAND2_X1 U969 ( .A1(n1168), .A2(n1287), .ZN(n1106) );
OR2_X1 U970 ( .A1(n1164), .A2(G902), .ZN(n1287) );
XNOR2_X1 U971 ( .A(n1104), .B(KEYINPUT14), .ZN(n1286) );
NOR3_X1 U972 ( .A1(n1168), .A2(G902), .A3(n1164), .ZN(n1104) );
XNOR2_X1 U973 ( .A(n1288), .B(n1289), .ZN(n1164) );
XOR2_X1 U974 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U975 ( .A(G125), .B(G119), .Z(n1291) );
XOR2_X1 U976 ( .A(KEYINPUT44), .B(G137), .Z(n1290) );
XOR2_X1 U977 ( .A(n1292), .B(n1293), .Z(n1288) );
XOR2_X1 U978 ( .A(n1294), .B(n1295), .Z(n1293) );
NAND3_X1 U979 ( .A1(n1296), .A2(n1121), .A3(G221), .ZN(n1295) );
NAND2_X1 U980 ( .A1(KEYINPUT45), .A2(n1253), .ZN(n1294) );
INV_X1 U981 ( .A(G146), .ZN(n1253) );
XNOR2_X1 U982 ( .A(n1297), .B(n1298), .ZN(n1292) );
AND2_X1 U983 ( .A1(G217), .A2(n1299), .ZN(n1168) );
INV_X1 U984 ( .A(n1088), .ZN(n1283) );
NAND3_X1 U985 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1088) );
INV_X1 U986 ( .A(n1103), .ZN(n1302) );
NOR2_X1 U987 ( .A1(n1110), .A2(G472), .ZN(n1103) );
NAND3_X1 U988 ( .A1(KEYINPUT48), .A2(G472), .A3(n1110), .ZN(n1301) );
OR2_X1 U989 ( .A1(n1110), .A2(KEYINPUT48), .ZN(n1300) );
NAND2_X1 U990 ( .A1(n1303), .A2(n1189), .ZN(n1110) );
XOR2_X1 U991 ( .A(n1304), .B(n1193), .Z(n1303) );
XNOR2_X1 U992 ( .A(n1305), .B(n1306), .ZN(n1193) );
XNOR2_X1 U993 ( .A(KEYINPUT57), .B(KEYINPUT46), .ZN(n1305) );
XOR2_X1 U994 ( .A(n1307), .B(n1211), .Z(n1304) );
XOR2_X1 U995 ( .A(n1197), .B(n1194), .Z(n1211) );
NAND2_X1 U996 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U997 ( .A1(n1181), .A2(n1270), .ZN(n1309) );
XOR2_X1 U998 ( .A(KEYINPUT50), .B(n1310), .Z(n1308) );
NOR2_X1 U999 ( .A1(n1181), .A2(n1270), .ZN(n1310) );
NAND3_X1 U1000 ( .A1(n1311), .A2(n1121), .A3(G210), .ZN(n1181) );
AND2_X1 U1001 ( .A1(n1080), .A2(n1273), .ZN(n1229) );
NAND2_X1 U1002 ( .A1(n1065), .A2(n1312), .ZN(n1273) );
NAND3_X1 U1003 ( .A1(G902), .A2(n1277), .A3(n1154), .ZN(n1312) );
NOR2_X1 U1004 ( .A1(n1121), .A2(G898), .ZN(n1154) );
NAND3_X1 U1005 ( .A1(n1277), .A2(n1121), .A3(G952), .ZN(n1065) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1277) );
INV_X1 U1007 ( .A(n1247), .ZN(n1080) );
NAND2_X1 U1008 ( .A1(n1082), .A2(n1081), .ZN(n1247) );
INV_X1 U1009 ( .A(n1265), .ZN(n1081) );
NOR2_X1 U1010 ( .A1(n1313), .A2(n1105), .ZN(n1265) );
NOR3_X1 U1011 ( .A1(n1220), .A2(G902), .A3(n1219), .ZN(n1105) );
INV_X1 U1012 ( .A(n1218), .ZN(n1219) );
XOR2_X1 U1013 ( .A(n1108), .B(KEYINPUT53), .Z(n1313) );
AND2_X1 U1014 ( .A1(n1220), .A2(n1314), .ZN(n1108) );
NAND2_X1 U1015 ( .A1(n1218), .A2(n1189), .ZN(n1314) );
XNOR2_X1 U1016 ( .A(n1315), .B(n1316), .ZN(n1218) );
XNOR2_X1 U1017 ( .A(n1157), .B(n1155), .ZN(n1316) );
XOR2_X1 U1018 ( .A(n1317), .B(n1306), .Z(n1155) );
XNOR2_X1 U1019 ( .A(n1318), .B(n1319), .ZN(n1306) );
XOR2_X1 U1020 ( .A(G116), .B(G113), .Z(n1319) );
XOR2_X1 U1021 ( .A(n1320), .B(G119), .Z(n1318) );
XNOR2_X1 U1022 ( .A(KEYINPUT28), .B(KEYINPUT0), .ZN(n1320) );
XNOR2_X1 U1023 ( .A(G110), .B(G122), .ZN(n1317) );
XNOR2_X1 U1024 ( .A(n1321), .B(n1322), .ZN(n1157) );
XNOR2_X1 U1025 ( .A(G101), .B(KEYINPUT62), .ZN(n1321) );
XNOR2_X1 U1026 ( .A(n1323), .B(n1137), .ZN(n1315) );
XNOR2_X1 U1027 ( .A(G125), .B(n1324), .ZN(n1323) );
NOR2_X1 U1028 ( .A1(G953), .A2(n1147), .ZN(n1324) );
INV_X1 U1029 ( .A(G224), .ZN(n1147) );
AND2_X1 U1030 ( .A1(G210), .A2(n1325), .ZN(n1220) );
NAND2_X1 U1031 ( .A1(G214), .A2(n1325), .ZN(n1082) );
NAND2_X1 U1032 ( .A1(n1311), .A2(n1189), .ZN(n1325) );
AND2_X1 U1033 ( .A1(n1097), .A2(n1228), .ZN(n1095) );
NOR2_X1 U1034 ( .A1(n1116), .A2(n1069), .ZN(n1228) );
INV_X1 U1035 ( .A(n1096), .ZN(n1069) );
NAND2_X1 U1036 ( .A1(G221), .A2(n1299), .ZN(n1096) );
NAND2_X1 U1037 ( .A1(G234), .A2(n1189), .ZN(n1299) );
INV_X1 U1038 ( .A(n1285), .ZN(n1116) );
XNOR2_X1 U1039 ( .A(n1326), .B(G469), .ZN(n1285) );
NAND2_X1 U1040 ( .A1(n1327), .A2(n1189), .ZN(n1326) );
XOR2_X1 U1041 ( .A(n1328), .B(n1329), .Z(n1327) );
NOR2_X1 U1042 ( .A1(n1208), .A2(n1206), .ZN(n1329) );
NOR3_X1 U1043 ( .A1(n1297), .A2(G953), .A3(n1122), .ZN(n1206) );
INV_X1 U1044 ( .A(G227), .ZN(n1122) );
AND2_X1 U1045 ( .A1(n1297), .A2(n1330), .ZN(n1208) );
NAND2_X1 U1046 ( .A1(G227), .A2(n1121), .ZN(n1330) );
XNOR2_X1 U1047 ( .A(G110), .B(n1331), .ZN(n1297) );
INV_X1 U1048 ( .A(G140), .ZN(n1331) );
XOR2_X1 U1049 ( .A(n1332), .B(n1333), .Z(n1328) );
NOR2_X1 U1050 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1051 ( .A(KEYINPUT10), .B(n1336), .Z(n1335) );
NOR2_X1 U1052 ( .A1(n1337), .A2(n1194), .ZN(n1336) );
INV_X1 U1053 ( .A(n1137), .ZN(n1194) );
XOR2_X1 U1054 ( .A(n1210), .B(KEYINPUT18), .Z(n1337) );
NOR2_X1 U1055 ( .A1(n1137), .A2(n1210), .ZN(n1334) );
NAND3_X1 U1056 ( .A1(n1338), .A2(n1339), .A3(n1340), .ZN(n1210) );
NAND2_X1 U1057 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1058 ( .A(KEYINPUT47), .B(n1322), .Z(n1342) );
XNOR2_X1 U1059 ( .A(KEYINPUT2), .B(KEYINPUT9), .ZN(n1341) );
NAND2_X1 U1060 ( .A1(G101), .A2(n1343), .ZN(n1339) );
NAND3_X1 U1061 ( .A1(n1344), .A2(n1270), .A3(n1345), .ZN(n1338) );
INV_X1 U1062 ( .A(n1343), .ZN(n1345) );
NAND2_X1 U1063 ( .A1(n1346), .A2(KEYINPUT54), .ZN(n1343) );
XNOR2_X1 U1064 ( .A(KEYINPUT47), .B(n1322), .ZN(n1346) );
XOR2_X1 U1065 ( .A(G104), .B(G107), .Z(n1322) );
INV_X1 U1066 ( .A(G101), .ZN(n1270) );
XOR2_X1 U1067 ( .A(KEYINPUT9), .B(KEYINPUT2), .Z(n1344) );
XOR2_X1 U1068 ( .A(G146), .B(n1347), .Z(n1137) );
NAND2_X1 U1069 ( .A1(KEYINPUT32), .A2(n1197), .ZN(n1332) );
XNOR2_X1 U1070 ( .A(n1348), .B(n1349), .ZN(n1197) );
XOR2_X1 U1071 ( .A(G137), .B(G131), .Z(n1349) );
NAND2_X1 U1072 ( .A1(KEYINPUT13), .A2(n1350), .ZN(n1348) );
NOR2_X1 U1073 ( .A1(n1117), .A2(n1280), .ZN(n1097) );
INV_X1 U1074 ( .A(n1260), .ZN(n1280) );
NOR2_X1 U1075 ( .A1(n1115), .A2(n1351), .ZN(n1260) );
AND2_X1 U1076 ( .A1(G475), .A2(n1114), .ZN(n1351) );
NOR2_X1 U1077 ( .A1(n1114), .A2(G475), .ZN(n1115) );
NAND2_X1 U1078 ( .A1(n1175), .A2(n1189), .ZN(n1114) );
XNOR2_X1 U1079 ( .A(n1352), .B(n1353), .ZN(n1175) );
XOR2_X1 U1080 ( .A(G113), .B(n1354), .Z(n1353) );
XOR2_X1 U1081 ( .A(KEYINPUT34), .B(G122), .Z(n1354) );
XOR2_X1 U1082 ( .A(n1355), .B(G104), .Z(n1352) );
NAND2_X1 U1083 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1084 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1085 ( .A(KEYINPUT41), .B(n1360), .Z(n1356) );
NOR2_X1 U1086 ( .A1(n1359), .A2(n1358), .ZN(n1360) );
XOR2_X1 U1087 ( .A(n1361), .B(n1362), .Z(n1358) );
XNOR2_X1 U1088 ( .A(G140), .B(n1363), .ZN(n1362) );
NOR2_X1 U1089 ( .A1(G125), .A2(KEYINPUT36), .ZN(n1363) );
OR2_X1 U1090 ( .A1(G146), .A2(KEYINPUT19), .ZN(n1361) );
XNOR2_X1 U1091 ( .A(n1364), .B(n1365), .ZN(n1359) );
AND3_X1 U1092 ( .A1(G214), .A2(n1121), .A3(n1311), .ZN(n1365) );
INV_X1 U1093 ( .A(G237), .ZN(n1311) );
INV_X1 U1094 ( .A(G953), .ZN(n1121) );
XNOR2_X1 U1095 ( .A(G143), .B(G131), .ZN(n1364) );
XNOR2_X1 U1096 ( .A(n1366), .B(G478), .ZN(n1117) );
NAND2_X1 U1097 ( .A1(n1170), .A2(n1367), .ZN(n1366) );
XNOR2_X1 U1098 ( .A(KEYINPUT24), .B(n1189), .ZN(n1367) );
INV_X1 U1099 ( .A(G902), .ZN(n1189) );
XOR2_X1 U1100 ( .A(n1368), .B(n1369), .Z(n1170) );
XOR2_X1 U1101 ( .A(G107), .B(n1370), .Z(n1369) );
XOR2_X1 U1102 ( .A(G122), .B(G116), .Z(n1370) );
XNOR2_X1 U1103 ( .A(n1371), .B(n1350), .ZN(n1368) );
INV_X1 U1104 ( .A(n1132), .ZN(n1350) );
XOR2_X1 U1105 ( .A(G134), .B(KEYINPUT43), .Z(n1132) );
XOR2_X1 U1106 ( .A(n1372), .B(n1373), .Z(n1371) );
NOR3_X1 U1107 ( .A1(n1374), .A2(G953), .A3(n1375), .ZN(n1373) );
INV_X1 U1108 ( .A(n1296), .ZN(n1375) );
XOR2_X1 U1109 ( .A(G234), .B(KEYINPUT35), .Z(n1296) );
XOR2_X1 U1110 ( .A(KEYINPUT56), .B(G217), .Z(n1374) );
NAND2_X1 U1111 ( .A1(KEYINPUT40), .A2(n1347), .ZN(n1372) );
XNOR2_X1 U1112 ( .A(G143), .B(n1298), .ZN(n1347) );
XOR2_X1 U1113 ( .A(G128), .B(KEYINPUT58), .Z(n1298) );
endmodule


