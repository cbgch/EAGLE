//Key = 0000001001011011011111100111100001111000100111100001100100010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411;

XNOR2_X1 U775 ( .A(n1081), .B(n1082), .ZN(G9) );
NOR2_X1 U776 ( .A1(n1083), .A2(n1084), .ZN(G75) );
AND4_X1 U777 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
NAND3_X1 U778 ( .A1(n1089), .A2(n1090), .A3(KEYINPUT12), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NAND4_X1 U780 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NAND2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U783 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1097) );
NAND2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U786 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND3_X1 U787 ( .A1(n1099), .A2(n1109), .A3(n1103), .ZN(n1091) );
NAND2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND3_X1 U789 ( .A1(n1112), .A2(n1113), .A3(n1093), .ZN(n1111) );
NAND2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND3_X1 U791 ( .A1(n1116), .A2(n1117), .A3(n1096), .ZN(n1112) );
NAND2_X1 U792 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NAND2_X1 U793 ( .A1(n1094), .A2(n1120), .ZN(n1110) );
NOR3_X1 U794 ( .A1(n1121), .A2(G953), .A3(G952), .ZN(n1083) );
INV_X1 U795 ( .A(n1087), .ZN(n1121) );
NAND4_X1 U796 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1087) );
NOR4_X1 U797 ( .A1(n1114), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1125) );
XOR2_X1 U798 ( .A(KEYINPUT34), .B(n1129), .Z(n1128) );
NOR2_X1 U799 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U800 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
INV_X1 U801 ( .A(n1134), .ZN(n1133) );
XNOR2_X1 U802 ( .A(KEYINPUT5), .B(n1135), .ZN(n1132) );
NOR2_X1 U803 ( .A1(n1134), .A2(n1135), .ZN(n1130) );
XOR2_X1 U804 ( .A(n1136), .B(n1137), .Z(n1127) );
XOR2_X1 U805 ( .A(KEYINPUT50), .B(n1138), .Z(n1137) );
NAND2_X1 U806 ( .A1(KEYINPUT14), .A2(n1139), .ZN(n1136) );
NOR2_X1 U807 ( .A1(n1140), .A2(n1141), .ZN(n1126) );
AND2_X1 U808 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
AND2_X1 U809 ( .A1(n1099), .A2(n1118), .ZN(n1124) );
XOR2_X1 U810 ( .A(n1144), .B(G475), .Z(n1123) );
XOR2_X1 U811 ( .A(n1145), .B(KEYINPUT4), .Z(n1122) );
XOR2_X1 U812 ( .A(n1146), .B(n1147), .Z(G72) );
NOR2_X1 U813 ( .A1(n1148), .A2(n1088), .ZN(n1147) );
NOR2_X1 U814 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U815 ( .A1(KEYINPUT53), .A2(n1151), .ZN(n1146) );
NOR3_X1 U816 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
NOR2_X1 U817 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U818 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
INV_X1 U819 ( .A(KEYINPUT52), .ZN(n1158) );
XOR2_X1 U820 ( .A(n1159), .B(KEYINPUT40), .Z(n1157) );
AND3_X1 U821 ( .A1(n1156), .A2(n1159), .A3(KEYINPUT52), .ZN(n1153) );
AND2_X1 U822 ( .A1(n1088), .A2(n1160), .ZN(n1156) );
NOR2_X1 U823 ( .A1(KEYINPUT52), .A2(n1159), .ZN(n1152) );
NAND2_X1 U824 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
NAND2_X1 U825 ( .A1(n1163), .A2(n1150), .ZN(n1162) );
XOR2_X1 U826 ( .A(n1164), .B(n1165), .Z(n1161) );
XNOR2_X1 U827 ( .A(n1166), .B(n1167), .ZN(n1165) );
XOR2_X1 U828 ( .A(n1168), .B(n1169), .Z(n1164) );
XNOR2_X1 U829 ( .A(n1170), .B(G125), .ZN(n1169) );
NAND2_X1 U830 ( .A1(KEYINPUT61), .A2(n1171), .ZN(n1168) );
XOR2_X1 U831 ( .A(KEYINPUT42), .B(G140), .Z(n1171) );
NAND2_X1 U832 ( .A1(n1172), .A2(n1173), .ZN(G69) );
NAND2_X1 U833 ( .A1(n1174), .A2(n1088), .ZN(n1173) );
XOR2_X1 U834 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U835 ( .A1(KEYINPUT11), .A2(n1177), .ZN(n1176) );
NAND2_X1 U836 ( .A1(n1178), .A2(G953), .ZN(n1172) );
XOR2_X1 U837 ( .A(n1175), .B(n1179), .Z(n1178) );
NOR2_X1 U838 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND2_X1 U839 ( .A1(n1182), .A2(n1183), .ZN(n1175) );
NAND2_X1 U840 ( .A1(n1163), .A2(n1181), .ZN(n1183) );
XNOR2_X1 U841 ( .A(n1184), .B(n1185), .ZN(n1182) );
XNOR2_X1 U842 ( .A(KEYINPUT32), .B(n1186), .ZN(n1185) );
NOR2_X1 U843 ( .A1(KEYINPUT30), .A2(n1187), .ZN(n1186) );
NOR2_X1 U844 ( .A1(n1188), .A2(n1189), .ZN(G66) );
XOR2_X1 U845 ( .A(n1190), .B(n1143), .Z(n1189) );
NAND2_X1 U846 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U847 ( .A1(n1188), .A2(n1193), .ZN(G63) );
NOR3_X1 U848 ( .A1(n1134), .A2(n1194), .A3(n1195), .ZN(n1193) );
AND3_X1 U849 ( .A1(n1196), .A2(G478), .A3(n1191), .ZN(n1195) );
NOR2_X1 U850 ( .A1(n1197), .A2(n1196), .ZN(n1194) );
NOR2_X1 U851 ( .A1(n1085), .A2(n1135), .ZN(n1197) );
INV_X1 U852 ( .A(G478), .ZN(n1135) );
NOR2_X1 U853 ( .A1(n1188), .A2(n1198), .ZN(G60) );
NOR2_X1 U854 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U855 ( .A(n1201), .B(KEYINPUT21), .Z(n1200) );
NAND2_X1 U856 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U857 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
INV_X1 U858 ( .A(n1204), .ZN(n1203) );
AND2_X1 U859 ( .A1(n1191), .A2(G475), .ZN(n1202) );
XNOR2_X1 U860 ( .A(G104), .B(n1205), .ZN(G6) );
NAND4_X1 U861 ( .A1(n1206), .A2(n1094), .A3(n1207), .A4(n1208), .ZN(n1205) );
OR2_X1 U862 ( .A1(n1209), .A2(KEYINPUT47), .ZN(n1208) );
NAND2_X1 U863 ( .A1(KEYINPUT47), .A2(n1210), .ZN(n1207) );
NAND3_X1 U864 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
NOR2_X1 U865 ( .A1(n1188), .A2(n1214), .ZN(G57) );
XOR2_X1 U866 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR2_X1 U867 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
NOR2_X1 U868 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NOR2_X1 U869 ( .A1(n1221), .A2(KEYINPUT8), .ZN(n1219) );
NOR2_X1 U870 ( .A1(KEYINPUT3), .A2(n1222), .ZN(n1221) );
NOR2_X1 U871 ( .A1(n1223), .A2(n1224), .ZN(n1217) );
NOR2_X1 U872 ( .A1(n1225), .A2(KEYINPUT3), .ZN(n1224) );
NOR2_X1 U873 ( .A1(KEYINPUT8), .A2(n1226), .ZN(n1225) );
INV_X1 U874 ( .A(n1220), .ZN(n1226) );
XNOR2_X1 U875 ( .A(n1227), .B(n1228), .ZN(n1220) );
XOR2_X1 U876 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U877 ( .A1(KEYINPUT25), .A2(n1231), .ZN(n1229) );
INV_X1 U878 ( .A(n1222), .ZN(n1223) );
NAND2_X1 U879 ( .A1(n1191), .A2(G472), .ZN(n1222) );
NOR3_X1 U880 ( .A1(n1188), .A2(n1232), .A3(n1233), .ZN(G54) );
NOR2_X1 U881 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U882 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND2_X1 U883 ( .A1(KEYINPUT43), .A2(n1238), .ZN(n1236) );
NOR2_X1 U884 ( .A1(n1231), .A2(n1239), .ZN(n1232) );
XOR2_X1 U885 ( .A(n1240), .B(n1237), .Z(n1239) );
XOR2_X1 U886 ( .A(n1241), .B(n1242), .Z(n1237) );
XNOR2_X1 U887 ( .A(n1243), .B(n1244), .ZN(n1242) );
XOR2_X1 U888 ( .A(n1245), .B(n1246), .Z(n1241) );
NOR2_X1 U889 ( .A1(G140), .A2(KEYINPUT16), .ZN(n1246) );
NAND2_X1 U890 ( .A1(n1191), .A2(G469), .ZN(n1245) );
NAND2_X1 U891 ( .A1(KEYINPUT43), .A2(n1247), .ZN(n1240) );
NOR2_X1 U892 ( .A1(n1188), .A2(n1248), .ZN(G51) );
XOR2_X1 U893 ( .A(n1249), .B(n1250), .Z(n1248) );
AND2_X1 U894 ( .A1(G210), .A2(n1191), .ZN(n1250) );
NOR2_X1 U895 ( .A1(n1142), .A2(n1085), .ZN(n1191) );
NOR2_X1 U896 ( .A1(n1160), .A2(n1177), .ZN(n1085) );
NAND4_X1 U897 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1177) );
NOR4_X1 U898 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
NOR2_X1 U899 ( .A1(n1212), .A2(n1259), .ZN(n1258) );
NOR3_X1 U900 ( .A1(n1101), .A2(n1260), .A3(n1115), .ZN(n1257) );
NOR2_X1 U901 ( .A1(n1261), .A2(n1082), .ZN(n1253) );
NOR3_X1 U902 ( .A1(n1115), .A2(n1260), .A3(n1102), .ZN(n1082) );
INV_X1 U903 ( .A(n1209), .ZN(n1260) );
INV_X1 U904 ( .A(n1094), .ZN(n1115) );
NAND4_X1 U905 ( .A1(n1262), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(n1160) );
AND4_X1 U906 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1269), .ZN(n1265) );
NOR3_X1 U907 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1264) );
NOR2_X1 U908 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
INV_X1 U909 ( .A(KEYINPUT19), .ZN(n1273) );
NOR4_X1 U910 ( .A1(KEYINPUT19), .A2(n1275), .A3(n1213), .A4(n1118), .ZN(n1271) );
NAND2_X1 U911 ( .A1(n1206), .A2(n1276), .ZN(n1275) );
NOR3_X1 U912 ( .A1(n1277), .A2(n1102), .A3(n1278), .ZN(n1270) );
INV_X1 U913 ( .A(n1279), .ZN(n1102) );
XNOR2_X1 U914 ( .A(KEYINPUT15), .B(n1117), .ZN(n1277) );
INV_X1 U915 ( .A(n1280), .ZN(n1117) );
NOR2_X1 U916 ( .A1(KEYINPUT10), .A2(n1281), .ZN(n1249) );
XOR2_X1 U917 ( .A(n1282), .B(KEYINPUT27), .Z(n1281) );
AND2_X1 U918 ( .A1(n1283), .A2(G953), .ZN(n1188) );
XNOR2_X1 U919 ( .A(G952), .B(KEYINPUT1), .ZN(n1283) );
XNOR2_X1 U920 ( .A(G146), .B(n1274), .ZN(G48) );
NAND4_X1 U921 ( .A1(n1206), .A2(n1276), .A3(n1213), .A4(n1284), .ZN(n1274) );
XNOR2_X1 U922 ( .A(G143), .B(n1266), .ZN(G45) );
NAND4_X1 U923 ( .A1(n1285), .A2(n1213), .A3(n1280), .A4(n1286), .ZN(n1266) );
NOR3_X1 U924 ( .A1(n1212), .A2(n1287), .A3(n1288), .ZN(n1286) );
XNOR2_X1 U925 ( .A(G140), .B(n1262), .ZN(G42) );
NAND4_X1 U926 ( .A1(n1289), .A2(n1206), .A3(n1118), .A4(n1119), .ZN(n1262) );
XNOR2_X1 U927 ( .A(G137), .B(n1263), .ZN(G39) );
NAND2_X1 U928 ( .A1(n1290), .A2(n1289), .ZN(n1263) );
XNOR2_X1 U929 ( .A(G134), .B(n1291), .ZN(G36) );
NAND4_X1 U930 ( .A1(n1292), .A2(n1293), .A3(n1280), .A4(n1279), .ZN(n1291) );
XNOR2_X1 U931 ( .A(n1287), .B(KEYINPUT7), .ZN(n1292) );
INV_X1 U932 ( .A(n1294), .ZN(n1287) );
XOR2_X1 U933 ( .A(n1269), .B(n1295), .Z(G33) );
NAND2_X1 U934 ( .A1(n1296), .A2(KEYINPUT26), .ZN(n1295) );
XNOR2_X1 U935 ( .A(G131), .B(KEYINPUT33), .ZN(n1296) );
NAND3_X1 U936 ( .A1(n1206), .A2(n1280), .A3(n1289), .ZN(n1269) );
INV_X1 U937 ( .A(n1278), .ZN(n1289) );
NAND2_X1 U938 ( .A1(n1293), .A2(n1294), .ZN(n1278) );
NOR3_X1 U939 ( .A1(n1105), .A2(n1114), .A3(n1297), .ZN(n1293) );
XNOR2_X1 U940 ( .A(G128), .B(n1268), .ZN(G30) );
NAND4_X1 U941 ( .A1(n1276), .A2(n1279), .A3(n1213), .A4(n1284), .ZN(n1268) );
INV_X1 U942 ( .A(n1105), .ZN(n1213) );
XOR2_X1 U943 ( .A(n1261), .B(n1298), .Z(G3) );
NOR2_X1 U944 ( .A1(KEYINPUT38), .A2(n1299), .ZN(n1298) );
AND3_X1 U945 ( .A1(n1280), .A2(n1209), .A3(n1103), .ZN(n1261) );
XNOR2_X1 U946 ( .A(G125), .B(n1267), .ZN(G27) );
NAND4_X1 U947 ( .A1(n1206), .A2(n1276), .A3(n1118), .A4(n1099), .ZN(n1267) );
AND3_X1 U948 ( .A1(n1294), .A2(n1119), .A3(n1120), .ZN(n1276) );
NAND2_X1 U949 ( .A1(n1300), .A2(n1301), .ZN(n1294) );
NAND2_X1 U950 ( .A1(n1302), .A2(n1150), .ZN(n1301) );
INV_X1 U951 ( .A(G900), .ZN(n1150) );
XOR2_X1 U952 ( .A(n1256), .B(n1303), .Z(G24) );
NOR2_X1 U953 ( .A1(KEYINPUT37), .A2(n1304), .ZN(n1303) );
AND4_X1 U954 ( .A1(n1285), .A2(n1099), .A3(n1305), .A4(n1094), .ZN(n1256) );
NOR2_X1 U955 ( .A1(n1119), .A2(n1284), .ZN(n1094) );
NOR2_X1 U956 ( .A1(n1288), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U957 ( .A(n1307), .B(KEYINPUT59), .ZN(n1288) );
XNOR2_X1 U958 ( .A(n1255), .B(n1308), .ZN(G21) );
XNOR2_X1 U959 ( .A(KEYINPUT51), .B(n1309), .ZN(n1308) );
AND3_X1 U960 ( .A1(n1099), .A2(n1310), .A3(n1290), .ZN(n1255) );
AND3_X1 U961 ( .A1(n1284), .A2(n1119), .A3(n1103), .ZN(n1290) );
XNOR2_X1 U962 ( .A(G116), .B(n1251), .ZN(G18) );
NAND4_X1 U963 ( .A1(n1280), .A2(n1099), .A3(n1279), .A4(n1310), .ZN(n1251) );
INV_X1 U964 ( .A(n1306), .ZN(n1310) );
NOR2_X1 U965 ( .A1(n1307), .A2(n1285), .ZN(n1279) );
XOR2_X1 U966 ( .A(n1311), .B(n1312), .Z(G15) );
NOR2_X1 U967 ( .A1(KEYINPUT60), .A2(n1313), .ZN(n1312) );
INV_X1 U968 ( .A(G113), .ZN(n1313) );
NOR2_X1 U969 ( .A1(n1314), .A2(n1212), .ZN(n1311) );
INV_X1 U970 ( .A(n1120), .ZN(n1212) );
XOR2_X1 U971 ( .A(n1259), .B(KEYINPUT29), .Z(n1314) );
NAND4_X1 U972 ( .A1(n1206), .A2(n1280), .A3(n1099), .A4(n1211), .ZN(n1259) );
NOR2_X1 U973 ( .A1(n1315), .A2(n1107), .ZN(n1099) );
INV_X1 U974 ( .A(n1316), .ZN(n1107) );
NOR2_X1 U975 ( .A1(n1119), .A2(n1118), .ZN(n1280) );
INV_X1 U976 ( .A(n1101), .ZN(n1206) );
NAND2_X1 U977 ( .A1(n1285), .A2(n1317), .ZN(n1101) );
XNOR2_X1 U978 ( .A(KEYINPUT24), .B(n1318), .ZN(n1317) );
XNOR2_X1 U979 ( .A(G110), .B(n1252), .ZN(G12) );
NAND4_X1 U980 ( .A1(n1103), .A2(n1209), .A3(n1118), .A4(n1119), .ZN(n1252) );
NAND2_X1 U981 ( .A1(n1319), .A2(n1145), .ZN(n1119) );
NAND3_X1 U982 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1145) );
NAND2_X1 U983 ( .A1(n1192), .A2(n1320), .ZN(n1319) );
NAND2_X1 U984 ( .A1(n1143), .A2(n1142), .ZN(n1320) );
XNOR2_X1 U985 ( .A(n1321), .B(n1322), .ZN(n1143) );
XNOR2_X1 U986 ( .A(n1323), .B(n1324), .ZN(n1322) );
NAND2_X1 U987 ( .A1(G221), .A2(n1325), .ZN(n1323) );
XOR2_X1 U988 ( .A(n1326), .B(n1327), .Z(n1321) );
NOR2_X1 U989 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U990 ( .A(n1330), .B(KEYINPUT9), .Z(n1329) );
NAND2_X1 U991 ( .A1(n1331), .A2(n1243), .ZN(n1330) );
NOR2_X1 U992 ( .A1(n1243), .A2(n1331), .ZN(n1328) );
XNOR2_X1 U993 ( .A(n1332), .B(n1333), .ZN(n1331) );
XNOR2_X1 U994 ( .A(n1334), .B(KEYINPUT28), .ZN(n1333) );
NAND2_X1 U995 ( .A1(KEYINPUT22), .A2(n1309), .ZN(n1334) );
XNOR2_X1 U996 ( .A(G137), .B(G146), .ZN(n1326) );
INV_X1 U997 ( .A(n1141), .ZN(n1192) );
NAND2_X1 U998 ( .A1(G217), .A2(n1335), .ZN(n1141) );
INV_X1 U999 ( .A(n1284), .ZN(n1118) );
XNOR2_X1 U1000 ( .A(n1336), .B(G472), .ZN(n1284) );
NAND2_X1 U1001 ( .A1(n1337), .A2(n1142), .ZN(n1336) );
XOR2_X1 U1002 ( .A(n1338), .B(n1216), .Z(n1337) );
XNOR2_X1 U1003 ( .A(n1339), .B(G101), .ZN(n1216) );
NAND2_X1 U1004 ( .A1(G210), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1005 ( .A(n1341), .B(KEYINPUT63), .Z(n1338) );
NAND2_X1 U1006 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1007 ( .A1(KEYINPUT57), .A2(n1344), .ZN(n1343) );
XNOR2_X1 U1008 ( .A(n1231), .B(n1345), .ZN(n1342) );
XOR2_X1 U1009 ( .A(n1346), .B(n1230), .Z(n1345) );
OR2_X1 U1010 ( .A1(n1344), .A2(KEYINPUT57), .ZN(n1346) );
XOR2_X1 U1011 ( .A(n1227), .B(KEYINPUT20), .Z(n1344) );
XOR2_X1 U1012 ( .A(n1187), .B(KEYINPUT41), .Z(n1227) );
NOR2_X1 U1013 ( .A1(n1105), .A2(n1306), .ZN(n1209) );
NAND2_X1 U1014 ( .A1(n1120), .A2(n1211), .ZN(n1306) );
NAND2_X1 U1015 ( .A1(n1300), .A2(n1347), .ZN(n1211) );
NAND2_X1 U1016 ( .A1(n1302), .A2(n1181), .ZN(n1347) );
INV_X1 U1017 ( .A(G898), .ZN(n1181) );
AND3_X1 U1018 ( .A1(G902), .A2(n1090), .A3(n1163), .ZN(n1302) );
XNOR2_X1 U1019 ( .A(G953), .B(KEYINPUT6), .ZN(n1163) );
NAND3_X1 U1020 ( .A1(n1090), .A2(n1088), .A3(G952), .ZN(n1300) );
NAND2_X1 U1021 ( .A1(G237), .A2(G234), .ZN(n1090) );
NOR2_X1 U1022 ( .A1(n1093), .A2(n1114), .ZN(n1120) );
INV_X1 U1023 ( .A(n1096), .ZN(n1114) );
NAND2_X1 U1024 ( .A1(G214), .A2(n1348), .ZN(n1096) );
INV_X1 U1025 ( .A(n1297), .ZN(n1093) );
XNOR2_X1 U1026 ( .A(n1138), .B(n1139), .ZN(n1297) );
NAND2_X1 U1027 ( .A1(n1349), .A2(n1348), .ZN(n1139) );
NAND2_X1 U1028 ( .A1(n1350), .A2(n1142), .ZN(n1348) );
INV_X1 U1029 ( .A(G237), .ZN(n1350) );
XNOR2_X1 U1030 ( .A(G210), .B(KEYINPUT55), .ZN(n1349) );
NOR2_X1 U1031 ( .A1(n1282), .A2(G902), .ZN(n1138) );
XOR2_X1 U1032 ( .A(n1351), .B(n1352), .Z(n1282) );
XOR2_X1 U1033 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1034 ( .A(G125), .B(n1355), .ZN(n1354) );
NOR2_X1 U1035 ( .A1(G953), .A2(n1180), .ZN(n1355) );
INV_X1 U1036 ( .A(G224), .ZN(n1180) );
NAND2_X1 U1037 ( .A1(KEYINPUT44), .A2(n1187), .ZN(n1353) );
XNOR2_X1 U1038 ( .A(G113), .B(n1356), .ZN(n1187) );
XNOR2_X1 U1039 ( .A(n1309), .B(G116), .ZN(n1356) );
INV_X1 U1040 ( .A(G119), .ZN(n1309) );
XNOR2_X1 U1041 ( .A(n1230), .B(n1357), .ZN(n1351) );
INV_X1 U1042 ( .A(n1184), .ZN(n1357) );
XNOR2_X1 U1043 ( .A(n1358), .B(n1359), .ZN(n1184) );
XNOR2_X1 U1044 ( .A(n1299), .B(n1360), .ZN(n1359) );
NOR2_X1 U1045 ( .A1(G107), .A2(KEYINPUT2), .ZN(n1360) );
XNOR2_X1 U1046 ( .A(G104), .B(n1361), .ZN(n1358) );
XNOR2_X1 U1047 ( .A(n1304), .B(G110), .ZN(n1361) );
XNOR2_X1 U1048 ( .A(n1362), .B(n1332), .ZN(n1230) );
XNOR2_X1 U1049 ( .A(n1363), .B(n1364), .ZN(n1362) );
NAND2_X1 U1050 ( .A1(KEYINPUT35), .A2(n1365), .ZN(n1363) );
NAND2_X1 U1051 ( .A1(n1366), .A2(n1316), .ZN(n1105) );
NAND2_X1 U1052 ( .A1(G221), .A2(n1335), .ZN(n1316) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1142), .ZN(n1335) );
XNOR2_X1 U1054 ( .A(KEYINPUT49), .B(n1108), .ZN(n1366) );
INV_X1 U1055 ( .A(n1315), .ZN(n1108) );
XNOR2_X1 U1056 ( .A(n1367), .B(G469), .ZN(n1315) );
NAND2_X1 U1057 ( .A1(n1368), .A2(n1142), .ZN(n1367) );
INV_X1 U1058 ( .A(G902), .ZN(n1142) );
XOR2_X1 U1059 ( .A(n1369), .B(n1370), .Z(n1368) );
XNOR2_X1 U1060 ( .A(n1238), .B(n1371), .ZN(n1370) );
NOR2_X1 U1061 ( .A1(KEYINPUT39), .A2(n1234), .ZN(n1371) );
INV_X1 U1062 ( .A(n1231), .ZN(n1234) );
XOR2_X1 U1063 ( .A(G131), .B(n1372), .Z(n1231) );
NOR2_X1 U1064 ( .A1(KEYINPUT56), .A2(n1167), .ZN(n1372) );
XNOR2_X1 U1065 ( .A(G134), .B(G137), .ZN(n1167) );
INV_X1 U1066 ( .A(n1247), .ZN(n1238) );
NAND2_X1 U1067 ( .A1(n1373), .A2(n1374), .ZN(n1247) );
NAND2_X1 U1068 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
XNOR2_X1 U1069 ( .A(G104), .B(G107), .ZN(n1375) );
NAND2_X1 U1070 ( .A1(n1377), .A2(n1378), .ZN(n1373) );
XNOR2_X1 U1071 ( .A(n1081), .B(G104), .ZN(n1378) );
XNOR2_X1 U1072 ( .A(n1376), .B(KEYINPUT0), .ZN(n1377) );
XOR2_X1 U1073 ( .A(n1166), .B(n1299), .Z(n1376) );
INV_X1 U1074 ( .A(G101), .ZN(n1299) );
XNOR2_X1 U1075 ( .A(n1379), .B(n1380), .ZN(n1166) );
NOR2_X1 U1076 ( .A1(KEYINPUT48), .A2(n1381), .ZN(n1380) );
XOR2_X1 U1077 ( .A(n1382), .B(n1365), .Z(n1381) );
XNOR2_X1 U1078 ( .A(n1383), .B(KEYINPUT46), .ZN(n1365) );
NAND2_X1 U1079 ( .A1(KEYINPUT18), .A2(n1364), .ZN(n1382) );
XNOR2_X1 U1080 ( .A(n1244), .B(n1384), .ZN(n1369) );
XNOR2_X1 U1081 ( .A(G140), .B(n1243), .ZN(n1384) );
INV_X1 U1082 ( .A(G110), .ZN(n1243) );
NOR2_X1 U1083 ( .A1(n1149), .A2(G953), .ZN(n1244) );
INV_X1 U1084 ( .A(G227), .ZN(n1149) );
NOR2_X1 U1085 ( .A1(n1318), .A2(n1285), .ZN(n1103) );
XOR2_X1 U1086 ( .A(n1385), .B(G475), .Z(n1285) );
NAND2_X1 U1087 ( .A1(KEYINPUT17), .A2(n1144), .ZN(n1385) );
NAND2_X1 U1088 ( .A1(n1386), .A2(n1204), .ZN(n1144) );
XNOR2_X1 U1089 ( .A(n1387), .B(n1388), .ZN(n1204) );
XOR2_X1 U1090 ( .A(n1389), .B(n1390), .Z(n1388) );
XOR2_X1 U1091 ( .A(n1391), .B(n1392), .Z(n1390) );
AND2_X1 U1092 ( .A1(n1340), .A2(G214), .ZN(n1392) );
NOR2_X1 U1093 ( .A1(G953), .A2(G237), .ZN(n1340) );
NAND2_X1 U1094 ( .A1(n1393), .A2(n1394), .ZN(n1391) );
NAND2_X1 U1095 ( .A1(n1324), .A2(n1395), .ZN(n1394) );
NAND2_X1 U1096 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
NAND2_X1 U1097 ( .A1(n1364), .A2(n1398), .ZN(n1397) );
INV_X1 U1098 ( .A(G146), .ZN(n1364) );
INV_X1 U1099 ( .A(KEYINPUT13), .ZN(n1396) );
NAND2_X1 U1100 ( .A1(G146), .A2(n1399), .ZN(n1393) );
NAND2_X1 U1101 ( .A1(n1398), .A2(n1400), .ZN(n1399) );
OR2_X1 U1102 ( .A1(n1324), .A2(KEYINPUT13), .ZN(n1400) );
XOR2_X1 U1103 ( .A(G125), .B(G140), .Z(n1324) );
INV_X1 U1104 ( .A(KEYINPUT23), .ZN(n1398) );
NAND2_X1 U1105 ( .A1(KEYINPUT62), .A2(n1170), .ZN(n1389) );
INV_X1 U1106 ( .A(G131), .ZN(n1170) );
XOR2_X1 U1107 ( .A(n1401), .B(n1402), .Z(n1387) );
XNOR2_X1 U1108 ( .A(n1383), .B(G122), .ZN(n1402) );
INV_X1 U1109 ( .A(G143), .ZN(n1383) );
XNOR2_X1 U1110 ( .A(G113), .B(G104), .ZN(n1401) );
XNOR2_X1 U1111 ( .A(G902), .B(KEYINPUT54), .ZN(n1386) );
INV_X1 U1112 ( .A(n1307), .ZN(n1318) );
XOR2_X1 U1113 ( .A(G478), .B(n1403), .Z(n1307) );
NOR2_X1 U1114 ( .A1(n1134), .A2(KEYINPUT31), .ZN(n1403) );
NOR2_X1 U1115 ( .A1(n1196), .A2(G902), .ZN(n1134) );
XOR2_X1 U1116 ( .A(n1404), .B(n1405), .Z(n1196) );
XNOR2_X1 U1117 ( .A(n1406), .B(n1332), .ZN(n1405) );
INV_X1 U1118 ( .A(n1379), .ZN(n1332) );
XOR2_X1 U1119 ( .A(G128), .B(KEYINPUT36), .Z(n1379) );
AND2_X1 U1120 ( .A1(n1325), .A2(G217), .ZN(n1406) );
AND2_X1 U1121 ( .A1(G234), .A2(n1088), .ZN(n1325) );
INV_X1 U1122 ( .A(G953), .ZN(n1088) );
XOR2_X1 U1123 ( .A(n1407), .B(n1408), .Z(n1404) );
NOR2_X1 U1124 ( .A1(KEYINPUT58), .A2(n1409), .ZN(n1408) );
XOR2_X1 U1125 ( .A(n1410), .B(n1411), .Z(n1409) );
XNOR2_X1 U1126 ( .A(n1304), .B(G116), .ZN(n1411) );
INV_X1 U1127 ( .A(G122), .ZN(n1304) );
NAND2_X1 U1128 ( .A1(KEYINPUT45), .A2(n1081), .ZN(n1410) );
INV_X1 U1129 ( .A(G107), .ZN(n1081) );
XNOR2_X1 U1130 ( .A(G134), .B(G143), .ZN(n1407) );
endmodule


