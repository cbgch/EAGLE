//Key = 1011001101111010010000010100110011100000110100010011110100011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;

XOR2_X1 U680 ( .A(G107), .B(n934), .Z(G9) );
NOR2_X1 U681 ( .A1(n935), .A2(n936), .ZN(G75) );
NOR3_X1 U682 ( .A1(n937), .A2(n938), .A3(n939), .ZN(n936) );
INV_X1 U683 ( .A(G952), .ZN(n938) );
NAND3_X1 U684 ( .A1(n940), .A2(n941), .A3(n942), .ZN(n937) );
NAND2_X1 U685 ( .A1(n943), .A2(n944), .ZN(n942) );
NAND2_X1 U686 ( .A1(n945), .A2(n946), .ZN(n944) );
NAND3_X1 U687 ( .A1(n947), .A2(n948), .A3(n949), .ZN(n946) );
NAND2_X1 U688 ( .A1(n950), .A2(n951), .ZN(n948) );
NAND2_X1 U689 ( .A1(n952), .A2(n953), .ZN(n951) );
NAND2_X1 U690 ( .A1(n954), .A2(n955), .ZN(n953) );
NAND2_X1 U691 ( .A1(n956), .A2(n957), .ZN(n955) );
NAND2_X1 U692 ( .A1(n958), .A2(n959), .ZN(n950) );
NAND2_X1 U693 ( .A1(n960), .A2(n961), .ZN(n959) );
XOR2_X1 U694 ( .A(KEYINPUT53), .B(n962), .Z(n960) );
NAND3_X1 U695 ( .A1(n952), .A2(n963), .A3(n958), .ZN(n945) );
NAND2_X1 U696 ( .A1(n964), .A2(n965), .ZN(n963) );
NAND2_X1 U697 ( .A1(n949), .A2(n966), .ZN(n965) );
NAND2_X1 U698 ( .A1(n967), .A2(n968), .ZN(n966) );
NAND2_X1 U699 ( .A1(n947), .A2(n969), .ZN(n964) );
NAND3_X1 U700 ( .A1(n970), .A2(n971), .A3(n972), .ZN(n969) );
NAND2_X1 U701 ( .A1(n949), .A2(n973), .ZN(n971) );
INV_X1 U702 ( .A(KEYINPUT61), .ZN(n973) );
NAND3_X1 U703 ( .A1(n974), .A2(n975), .A3(KEYINPUT61), .ZN(n970) );
INV_X1 U704 ( .A(n976), .ZN(n943) );
NOR3_X1 U705 ( .A1(n977), .A2(G953), .A3(n978), .ZN(n935) );
INV_X1 U706 ( .A(n940), .ZN(n978) );
NAND4_X1 U707 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(n940) );
NOR4_X1 U708 ( .A1(n956), .A2(n974), .A3(n983), .A4(n984), .ZN(n982) );
XNOR2_X1 U709 ( .A(n985), .B(KEYINPUT54), .ZN(n981) );
XNOR2_X1 U710 ( .A(n986), .B(n987), .ZN(n980) );
XNOR2_X1 U711 ( .A(n988), .B(KEYINPUT44), .ZN(n979) );
XNOR2_X1 U712 ( .A(G952), .B(KEYINPUT41), .ZN(n977) );
NAND2_X1 U713 ( .A1(n989), .A2(n990), .ZN(G72) );
NAND2_X1 U714 ( .A1(n991), .A2(n992), .ZN(n990) );
XOR2_X1 U715 ( .A(n993), .B(KEYINPUT48), .Z(n989) );
OR2_X1 U716 ( .A1(n992), .A2(n991), .ZN(n993) );
NAND2_X1 U717 ( .A1(G953), .A2(n994), .ZN(n991) );
NAND2_X1 U718 ( .A1(G900), .A2(G227), .ZN(n994) );
NAND2_X1 U719 ( .A1(n995), .A2(n996), .ZN(n992) );
NAND3_X1 U720 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
NAND2_X1 U721 ( .A1(n1000), .A2(n941), .ZN(n998) );
NAND2_X1 U722 ( .A1(n1001), .A2(G953), .ZN(n997) );
XOR2_X1 U723 ( .A(KEYINPUT43), .B(n1002), .Z(n995) );
NOR3_X1 U724 ( .A1(n999), .A2(G953), .A3(n1003), .ZN(n1002) );
AND2_X1 U725 ( .A1(n1004), .A2(n1005), .ZN(n999) );
NAND3_X1 U726 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1005) );
INV_X1 U727 ( .A(n1009), .ZN(n1008) );
XOR2_X1 U728 ( .A(n1010), .B(KEYINPUT45), .Z(n1004) );
NAND2_X1 U729 ( .A1(n1009), .A2(n1011), .ZN(n1010) );
NAND2_X1 U730 ( .A1(n1006), .A2(n1007), .ZN(n1011) );
INV_X1 U731 ( .A(n1012), .ZN(n1006) );
XOR2_X1 U732 ( .A(n1013), .B(n1014), .Z(n1009) );
XNOR2_X1 U733 ( .A(KEYINPUT35), .B(n1015), .ZN(n1014) );
XOR2_X1 U734 ( .A(n1016), .B(n1017), .Z(G69) );
NOR2_X1 U735 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR2_X1 U736 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
XOR2_X1 U737 ( .A(n1022), .B(KEYINPUT5), .Z(n1021) );
NAND2_X1 U738 ( .A1(n941), .A2(n1023), .ZN(n1022) );
NOR2_X1 U739 ( .A1(n1024), .A2(n1025), .ZN(n1020) );
NOR3_X1 U740 ( .A1(n1025), .A2(n1024), .A3(n1026), .ZN(n1018) );
AND2_X1 U741 ( .A1(n941), .A2(n1023), .ZN(n1026) );
NAND3_X1 U742 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1023) );
XNOR2_X1 U743 ( .A(KEYINPUT2), .B(n1030), .ZN(n1027) );
XNOR2_X1 U744 ( .A(n1031), .B(n1032), .ZN(n1025) );
NOR2_X1 U745 ( .A1(n1033), .A2(n1024), .ZN(n1016) );
NOR2_X1 U746 ( .A1(G224), .A2(n941), .ZN(n1033) );
NOR2_X1 U747 ( .A1(n1034), .A2(n1035), .ZN(G66) );
XNOR2_X1 U748 ( .A(n1036), .B(n1037), .ZN(n1035) );
XOR2_X1 U749 ( .A(KEYINPUT36), .B(n1038), .Z(n1037) );
NOR2_X1 U750 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U751 ( .A1(n1034), .A2(n1041), .ZN(G63) );
XOR2_X1 U752 ( .A(n1042), .B(n1043), .Z(n1041) );
XNOR2_X1 U753 ( .A(n1044), .B(KEYINPUT40), .ZN(n1043) );
NAND3_X1 U754 ( .A1(n1045), .A2(G478), .A3(KEYINPUT6), .ZN(n1044) );
NOR2_X1 U755 ( .A1(n1034), .A2(n1046), .ZN(G60) );
XOR2_X1 U756 ( .A(n1047), .B(n1048), .Z(n1046) );
AND2_X1 U757 ( .A1(G475), .A2(n1045), .ZN(n1048) );
NAND2_X1 U758 ( .A1(n1049), .A2(KEYINPUT9), .ZN(n1047) );
XNOR2_X1 U759 ( .A(n1050), .B(KEYINPUT11), .ZN(n1049) );
XNOR2_X1 U760 ( .A(G104), .B(n1051), .ZN(G6) );
NAND2_X1 U761 ( .A1(KEYINPUT59), .A2(n1052), .ZN(n1051) );
INV_X1 U762 ( .A(n1030), .ZN(n1052) );
NOR2_X1 U763 ( .A1(n1034), .A2(n1053), .ZN(G57) );
XOR2_X1 U764 ( .A(n1054), .B(n1055), .Z(n1053) );
AND2_X1 U765 ( .A1(G472), .A2(n1045), .ZN(n1054) );
INV_X1 U766 ( .A(n1040), .ZN(n1045) );
NOR2_X1 U767 ( .A1(n1034), .A2(n1056), .ZN(G54) );
XOR2_X1 U768 ( .A(n1057), .B(n1058), .Z(n1056) );
XOR2_X1 U769 ( .A(n1059), .B(n1060), .Z(n1058) );
XNOR2_X1 U770 ( .A(KEYINPUT27), .B(n1061), .ZN(n1060) );
XOR2_X1 U771 ( .A(n1062), .B(n1063), .Z(n1057) );
NOR3_X1 U772 ( .A1(n1040), .A2(KEYINPUT22), .A3(n1064), .ZN(n1063) );
XOR2_X1 U773 ( .A(n1065), .B(n1066), .Z(n1062) );
NOR2_X1 U774 ( .A1(G140), .A2(KEYINPUT56), .ZN(n1066) );
NAND2_X1 U775 ( .A1(KEYINPUT50), .A2(n1067), .ZN(n1065) );
XNOR2_X1 U776 ( .A(n1013), .B(n1068), .ZN(n1067) );
NOR2_X1 U777 ( .A1(n1034), .A2(n1069), .ZN(G51) );
XOR2_X1 U778 ( .A(n1070), .B(n1071), .Z(n1069) );
XOR2_X1 U779 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR3_X1 U780 ( .A1(n1040), .A2(KEYINPUT58), .A3(n987), .ZN(n1072) );
NAND2_X1 U781 ( .A1(n1074), .A2(n939), .ZN(n1040) );
NAND4_X1 U782 ( .A1(n1003), .A2(n1029), .A3(n1075), .A4(n1030), .ZN(n939) );
NAND3_X1 U783 ( .A1(n1076), .A2(n947), .A3(n1077), .ZN(n1030) );
XNOR2_X1 U784 ( .A(KEYINPUT23), .B(n1028), .ZN(n1075) );
AND4_X1 U785 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1029) );
NOR3_X1 U786 ( .A1(n1082), .A2(n1083), .A3(n934), .ZN(n1081) );
AND3_X1 U787 ( .A1(n962), .A2(n947), .A3(n1076), .ZN(n934) );
NAND4_X1 U788 ( .A1(n1084), .A2(n962), .A3(n1085), .A4(n1086), .ZN(n1080) );
OR2_X1 U789 ( .A1(n1087), .A2(KEYINPUT57), .ZN(n1086) );
NAND2_X1 U790 ( .A1(KEYINPUT57), .A2(n1088), .ZN(n1085) );
NAND3_X1 U791 ( .A1(n958), .A2(n1089), .A3(n1090), .ZN(n1088) );
INV_X1 U792 ( .A(n1000), .ZN(n1003) );
NAND4_X1 U793 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1000) );
AND4_X1 U794 ( .A1(n1095), .A2(n1096), .A3(n1097), .A4(n1098), .ZN(n1094) );
NOR3_X1 U795 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1093) );
NOR3_X1 U796 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
AND2_X1 U797 ( .A1(n1102), .A2(n1105), .ZN(n1100) );
INV_X1 U798 ( .A(KEYINPUT20), .ZN(n1102) );
XNOR2_X1 U799 ( .A(KEYINPUT46), .B(n1106), .ZN(n1074) );
XNOR2_X1 U800 ( .A(n1107), .B(n1108), .ZN(n1070) );
NOR2_X1 U801 ( .A1(KEYINPUT1), .A2(n1109), .ZN(n1108) );
XOR2_X1 U802 ( .A(n1110), .B(n1031), .Z(n1109) );
XOR2_X1 U803 ( .A(n1111), .B(n1112), .Z(n1031) );
NOR2_X1 U804 ( .A1(n941), .A2(G952), .ZN(n1034) );
XOR2_X1 U805 ( .A(n1096), .B(n1113), .Z(G48) );
XNOR2_X1 U806 ( .A(KEYINPUT10), .B(n1114), .ZN(n1113) );
NAND4_X1 U807 ( .A1(n1115), .A2(n1116), .A3(n1077), .A4(n1089), .ZN(n1096) );
XOR2_X1 U808 ( .A(n1117), .B(n1099), .Z(G45) );
AND3_X1 U809 ( .A1(n1084), .A2(n1116), .A3(n1118), .ZN(n1099) );
NOR3_X1 U810 ( .A1(n972), .A2(n1119), .A3(n1120), .ZN(n1118) );
NOR2_X1 U811 ( .A1(KEYINPUT63), .A2(n1121), .ZN(n1117) );
XNOR2_X1 U812 ( .A(KEYINPUT14), .B(n1122), .ZN(n1121) );
XNOR2_X1 U813 ( .A(G140), .B(n1091), .ZN(G42) );
NAND3_X1 U814 ( .A1(n1123), .A2(n1077), .A3(n1124), .ZN(n1091) );
XNOR2_X1 U815 ( .A(G137), .B(n1092), .ZN(G39) );
NAND3_X1 U816 ( .A1(n1115), .A2(n1123), .A3(n952), .ZN(n1092) );
XNOR2_X1 U817 ( .A(G134), .B(n1098), .ZN(G36) );
NAND3_X1 U818 ( .A1(n1123), .A2(n962), .A3(n1084), .ZN(n1098) );
XNOR2_X1 U819 ( .A(G131), .B(n1095), .ZN(G33) );
NAND3_X1 U820 ( .A1(n1123), .A2(n1077), .A3(n1084), .ZN(n1095) );
AND2_X1 U821 ( .A1(n1116), .A2(n949), .ZN(n1123) );
AND2_X1 U822 ( .A1(n975), .A2(n1125), .ZN(n949) );
XNOR2_X1 U823 ( .A(G128), .B(n1097), .ZN(G30) );
NAND4_X1 U824 ( .A1(n1115), .A2(n1116), .A3(n962), .A4(n1089), .ZN(n1097) );
NOR2_X1 U825 ( .A1(n954), .A2(n1126), .ZN(n1116) );
XNOR2_X1 U826 ( .A(G101), .B(n1127), .ZN(G3) );
NAND2_X1 U827 ( .A1(KEYINPUT17), .A2(n1128), .ZN(n1127) );
INV_X1 U828 ( .A(n1028), .ZN(n1128) );
NAND3_X1 U829 ( .A1(n1084), .A2(n1076), .A3(n952), .ZN(n1028) );
XOR2_X1 U830 ( .A(G125), .B(n1105), .Z(G27) );
NOR2_X1 U831 ( .A1(n1104), .A2(n1126), .ZN(n1105) );
INV_X1 U832 ( .A(n1103), .ZN(n1126) );
NAND2_X1 U833 ( .A1(n976), .A2(n1129), .ZN(n1103) );
NAND4_X1 U834 ( .A1(n1001), .A2(G902), .A3(G953), .A4(n1130), .ZN(n1129) );
XNOR2_X1 U835 ( .A(G900), .B(KEYINPUT37), .ZN(n1001) );
NAND4_X1 U836 ( .A1(n958), .A2(n1124), .A3(n1077), .A4(n1089), .ZN(n1104) );
XNOR2_X1 U837 ( .A(G122), .B(n1078), .ZN(G24) );
NAND4_X1 U838 ( .A1(n1087), .A2(n947), .A3(n988), .A4(n984), .ZN(n1078) );
INV_X1 U839 ( .A(n983), .ZN(n947) );
NAND2_X1 U840 ( .A1(n1131), .A2(n1132), .ZN(n983) );
XNOR2_X1 U841 ( .A(G119), .B(n1079), .ZN(G21) );
NAND3_X1 U842 ( .A1(n952), .A2(n1115), .A3(n1087), .ZN(n1079) );
AND2_X1 U843 ( .A1(n1133), .A2(n1134), .ZN(n1115) );
NAND2_X1 U844 ( .A1(n1135), .A2(n1136), .ZN(G18) );
NAND2_X1 U845 ( .A1(G116), .A2(n1137), .ZN(n1136) );
XOR2_X1 U846 ( .A(n1138), .B(KEYINPUT24), .Z(n1135) );
OR2_X1 U847 ( .A1(n1137), .A2(G116), .ZN(n1138) );
NAND3_X1 U848 ( .A1(n1084), .A2(n962), .A3(n1087), .ZN(n1137) );
INV_X1 U849 ( .A(n1139), .ZN(n1087) );
NOR2_X1 U850 ( .A1(n984), .A2(n1120), .ZN(n962) );
INV_X1 U851 ( .A(n988), .ZN(n1120) );
INV_X1 U852 ( .A(n967), .ZN(n1084) );
XNOR2_X1 U853 ( .A(n1083), .B(n1140), .ZN(G15) );
XNOR2_X1 U854 ( .A(G113), .B(KEYINPUT49), .ZN(n1140) );
NOR3_X1 U855 ( .A1(n967), .A2(n961), .A3(n1139), .ZN(n1083) );
NAND3_X1 U856 ( .A1(n1089), .A2(n1141), .A3(n958), .ZN(n1139) );
NOR2_X1 U857 ( .A1(n985), .A2(n956), .ZN(n958) );
INV_X1 U858 ( .A(n1077), .ZN(n961) );
NOR2_X1 U859 ( .A1(n988), .A2(n1119), .ZN(n1077) );
INV_X1 U860 ( .A(n984), .ZN(n1119) );
NAND2_X1 U861 ( .A1(n1131), .A2(n1133), .ZN(n967) );
XNOR2_X1 U862 ( .A(n1132), .B(KEYINPUT42), .ZN(n1133) );
INV_X1 U863 ( .A(n1134), .ZN(n1131) );
XNOR2_X1 U864 ( .A(n1061), .B(n1082), .ZN(G12) );
AND3_X1 U865 ( .A1(n952), .A2(n1076), .A3(n1124), .ZN(n1082) );
INV_X1 U866 ( .A(n968), .ZN(n1124) );
NAND2_X1 U867 ( .A1(n1132), .A2(n1134), .ZN(n968) );
XOR2_X1 U868 ( .A(n1142), .B(n1039), .Z(n1134) );
NAND2_X1 U869 ( .A1(G217), .A2(n1143), .ZN(n1039) );
NAND2_X1 U870 ( .A1(n1036), .A2(n1106), .ZN(n1142) );
XNOR2_X1 U871 ( .A(n1144), .B(n1145), .ZN(n1036) );
XNOR2_X1 U872 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U873 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U874 ( .A1(KEYINPUT15), .A2(n1114), .ZN(n1149) );
NAND3_X1 U875 ( .A1(n1150), .A2(n1151), .A3(n1007), .ZN(n1148) );
OR2_X1 U876 ( .A1(G140), .A2(KEYINPUT51), .ZN(n1151) );
NAND2_X1 U877 ( .A1(n1012), .A2(KEYINPUT51), .ZN(n1150) );
XOR2_X1 U878 ( .A(n1152), .B(n1153), .Z(n1144) );
XNOR2_X1 U879 ( .A(n1061), .B(n1154), .ZN(n1153) );
AND4_X1 U880 ( .A1(n1155), .A2(n941), .A3(G234), .A4(G221), .ZN(n1154) );
INV_X1 U881 ( .A(KEYINPUT4), .ZN(n1155) );
XNOR2_X1 U882 ( .A(G119), .B(KEYINPUT8), .ZN(n1152) );
XOR2_X1 U883 ( .A(n1156), .B(G472), .Z(n1132) );
NAND2_X1 U884 ( .A1(n1157), .A2(n1106), .ZN(n1156) );
XOR2_X1 U885 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U886 ( .A(KEYINPUT62), .B(KEYINPUT52), .Z(n1159) );
XNOR2_X1 U887 ( .A(n1055), .B(KEYINPUT0), .ZN(n1158) );
XNOR2_X1 U888 ( .A(n1160), .B(n1161), .ZN(n1055) );
XNOR2_X1 U889 ( .A(G143), .B(n1162), .ZN(n1161) );
NAND2_X1 U890 ( .A1(n1163), .A2(G210), .ZN(n1162) );
XNOR2_X1 U891 ( .A(n1164), .B(n1165), .ZN(n1160) );
INV_X1 U892 ( .A(n1013), .ZN(n1165) );
XOR2_X1 U893 ( .A(n1166), .B(n1146), .Z(n1013) );
XNOR2_X1 U894 ( .A(G137), .B(n1167), .ZN(n1146) );
NOR3_X1 U895 ( .A1(n954), .A2(n1090), .A3(n972), .ZN(n1076) );
INV_X1 U896 ( .A(n1089), .ZN(n972) );
NOR2_X1 U897 ( .A1(n975), .A2(n974), .ZN(n1089) );
INV_X1 U898 ( .A(n1125), .ZN(n974) );
NAND2_X1 U899 ( .A1(G214), .A2(n1168), .ZN(n1125) );
XNOR2_X1 U900 ( .A(n986), .B(n1169), .ZN(n975) );
NOR2_X1 U901 ( .A1(n1170), .A2(KEYINPUT13), .ZN(n1169) );
INV_X1 U902 ( .A(n987), .ZN(n1170) );
NAND2_X1 U903 ( .A1(G210), .A2(n1168), .ZN(n987) );
NAND2_X1 U904 ( .A1(n1171), .A2(n1106), .ZN(n1168) );
XNOR2_X1 U905 ( .A(G237), .B(KEYINPUT38), .ZN(n1171) );
NAND2_X1 U906 ( .A1(n1172), .A2(n1106), .ZN(n986) );
XOR2_X1 U907 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U908 ( .A(n1112), .B(n1073), .ZN(n1174) );
XNOR2_X1 U909 ( .A(n1175), .B(n1176), .ZN(n1073) );
XNOR2_X1 U910 ( .A(n1177), .B(n1178), .ZN(n1175) );
NAND2_X1 U911 ( .A1(G224), .A2(n941), .ZN(n1177) );
XOR2_X1 U912 ( .A(n1164), .B(n1110), .Z(n1173) );
AND2_X1 U913 ( .A1(KEYINPUT34), .A2(n1032), .ZN(n1110) );
XNOR2_X1 U914 ( .A(n1061), .B(n1179), .ZN(n1032) );
NOR2_X1 U915 ( .A1(KEYINPUT16), .A2(n1180), .ZN(n1179) );
XNOR2_X1 U916 ( .A(G122), .B(KEYINPUT55), .ZN(n1180) );
XOR2_X1 U917 ( .A(n1111), .B(n1107), .Z(n1164) );
NOR2_X1 U918 ( .A1(KEYINPUT30), .A2(n1114), .ZN(n1107) );
XOR2_X1 U919 ( .A(n1181), .B(n1182), .Z(n1111) );
XOR2_X1 U920 ( .A(G113), .B(G101), .Z(n1182) );
XNOR2_X1 U921 ( .A(G116), .B(n1183), .ZN(n1181) );
XNOR2_X1 U922 ( .A(KEYINPUT39), .B(n1184), .ZN(n1183) );
INV_X1 U923 ( .A(G119), .ZN(n1184) );
INV_X1 U924 ( .A(n1141), .ZN(n1090) );
NAND2_X1 U925 ( .A1(n976), .A2(n1185), .ZN(n1141) );
NAND3_X1 U926 ( .A1(n1024), .A2(n1130), .A3(G902), .ZN(n1185) );
NOR2_X1 U927 ( .A1(G898), .A2(n941), .ZN(n1024) );
NAND3_X1 U928 ( .A1(n1130), .A2(n941), .A3(G952), .ZN(n976) );
NAND2_X1 U929 ( .A1(G234), .A2(G237), .ZN(n1130) );
OR2_X1 U930 ( .A1(n957), .A2(n956), .ZN(n954) );
AND2_X1 U931 ( .A1(n1186), .A2(n1143), .ZN(n956) );
NAND2_X1 U932 ( .A1(G234), .A2(n1106), .ZN(n1143) );
XNOR2_X1 U933 ( .A(G221), .B(KEYINPUT60), .ZN(n1186) );
INV_X1 U934 ( .A(n985), .ZN(n957) );
XOR2_X1 U935 ( .A(n1187), .B(n1064), .Z(n985) );
INV_X1 U936 ( .A(G469), .ZN(n1064) );
NAND2_X1 U937 ( .A1(n1188), .A2(n1106), .ZN(n1187) );
XNOR2_X1 U938 ( .A(n1189), .B(n1167), .ZN(n1188) );
INV_X1 U939 ( .A(G128), .ZN(n1167) );
XOR2_X1 U940 ( .A(n1190), .B(n1191), .Z(n1189) );
XOR2_X1 U941 ( .A(n1192), .B(n1193), .Z(n1191) );
XNOR2_X1 U942 ( .A(KEYINPUT19), .B(n1194), .ZN(n1193) );
XOR2_X1 U943 ( .A(KEYINPUT47), .B(KEYINPUT26), .Z(n1192) );
XOR2_X1 U944 ( .A(n1195), .B(n1196), .Z(n1190) );
XOR2_X1 U945 ( .A(n1197), .B(n1068), .Z(n1196) );
XNOR2_X1 U946 ( .A(n1198), .B(n1112), .ZN(n1068) );
XNOR2_X1 U947 ( .A(G104), .B(G107), .ZN(n1112) );
XOR2_X1 U948 ( .A(n1015), .B(n1199), .Z(n1198) );
NOR2_X1 U949 ( .A1(KEYINPUT31), .A2(n1200), .ZN(n1199) );
XNOR2_X1 U950 ( .A(G101), .B(KEYINPUT32), .ZN(n1200) );
NAND2_X1 U951 ( .A1(n1201), .A2(n1202), .ZN(n1015) );
NAND2_X1 U952 ( .A1(G146), .A2(n1122), .ZN(n1202) );
XOR2_X1 U953 ( .A(KEYINPUT7), .B(n1203), .Z(n1201) );
NOR2_X1 U954 ( .A1(G146), .A2(n1122), .ZN(n1203) );
NAND2_X1 U955 ( .A1(KEYINPUT3), .A2(n1204), .ZN(n1197) );
XOR2_X1 U956 ( .A(n1166), .B(n1205), .Z(n1204) );
XNOR2_X1 U957 ( .A(KEYINPUT25), .B(n1206), .ZN(n1205) );
INV_X1 U958 ( .A(G137), .ZN(n1206) );
XOR2_X1 U959 ( .A(G131), .B(n1207), .Z(n1166) );
XNOR2_X1 U960 ( .A(G110), .B(n1059), .ZN(n1195) );
AND2_X1 U961 ( .A1(G227), .A2(n941), .ZN(n1059) );
NOR2_X1 U962 ( .A1(n988), .A2(n984), .ZN(n952) );
XNOR2_X1 U963 ( .A(n1208), .B(G475), .ZN(n984) );
NAND2_X1 U964 ( .A1(n1050), .A2(n1106), .ZN(n1208) );
XNOR2_X1 U965 ( .A(n1209), .B(G122), .ZN(n1050) );
XOR2_X1 U966 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U967 ( .A(n1212), .B(n1213), .Z(n1211) );
XOR2_X1 U968 ( .A(G131), .B(G113), .Z(n1213) );
XNOR2_X1 U969 ( .A(KEYINPUT33), .B(n1122), .ZN(n1212) );
XOR2_X1 U970 ( .A(n1214), .B(n1215), .Z(n1210) );
XOR2_X1 U971 ( .A(n1216), .B(n1217), .Z(n1215) );
NAND3_X1 U972 ( .A1(n1218), .A2(n1219), .A3(n1007), .ZN(n1217) );
NAND2_X1 U973 ( .A1(n1178), .A2(n1194), .ZN(n1007) );
OR2_X1 U974 ( .A1(G140), .A2(KEYINPUT28), .ZN(n1219) );
NAND2_X1 U975 ( .A1(KEYINPUT28), .A2(n1012), .ZN(n1218) );
NOR2_X1 U976 ( .A1(n1194), .A2(n1178), .ZN(n1012) );
XNOR2_X1 U977 ( .A(G125), .B(KEYINPUT18), .ZN(n1178) );
INV_X1 U978 ( .A(G140), .ZN(n1194) );
NAND2_X1 U979 ( .A1(KEYINPUT12), .A2(n1114), .ZN(n1216) );
INV_X1 U980 ( .A(G146), .ZN(n1114) );
XOR2_X1 U981 ( .A(n1220), .B(G104), .Z(n1214) );
NAND2_X1 U982 ( .A1(n1163), .A2(G214), .ZN(n1220) );
NOR2_X1 U983 ( .A1(G953), .A2(G237), .ZN(n1163) );
XNOR2_X1 U984 ( .A(n1221), .B(G478), .ZN(n988) );
NAND2_X1 U985 ( .A1(n1042), .A2(n1106), .ZN(n1221) );
INV_X1 U986 ( .A(G902), .ZN(n1106) );
XNOR2_X1 U987 ( .A(n1222), .B(n1223), .ZN(n1042) );
XOR2_X1 U988 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U989 ( .A(G116), .B(G107), .Z(n1225) );
AND3_X1 U990 ( .A1(G217), .A2(n941), .A3(G234), .ZN(n1224) );
INV_X1 U991 ( .A(G953), .ZN(n941) );
XNOR2_X1 U992 ( .A(n1176), .B(n1226), .ZN(n1222) );
XOR2_X1 U993 ( .A(n1227), .B(n1207), .Z(n1226) );
XOR2_X1 U994 ( .A(G134), .B(KEYINPUT29), .Z(n1207) );
NOR2_X1 U995 ( .A1(G122), .A2(KEYINPUT21), .ZN(n1227) );
XNOR2_X1 U996 ( .A(G128), .B(n1122), .ZN(n1176) );
INV_X1 U997 ( .A(G143), .ZN(n1122) );
INV_X1 U998 ( .A(G110), .ZN(n1061) );
endmodule


