//Key = 11011000011011111010001101011101000101111010001001100000000110111101100101010110100101111000101100001110001010111111000011101001
module c5315 ( G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, 
        G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, 
        G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, 
        G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, 
        G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, 
        G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, 
        G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, 
        G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, 
        G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, 
        G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, 
        G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, 
        G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, 
        G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, 
        G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, 
        G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, 
        G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, 
        G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, 
        G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, 
        G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, 
        G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, 
        G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, 
        G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, 
        G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, 
        G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, 
        G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, 
        G767, G807, G658, G690, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, 
        KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, 
        KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, 
        KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, 
        KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, 
        KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, 
        KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, 
        KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, 
        KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, 
        KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, 
        KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, 
        KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, 
        KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, 
        KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, 
        KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, 
        KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, 
        KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, 
        KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, 
        KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, 
        KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, 
        KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, 
        KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, 
        KEYINPUT125, KEYINPUT126, KEYINPUT127 );
  
input G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
         G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
         G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
         G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
         G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136,
         G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164,
         G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197,
         G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234,
         G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273,
         G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315,
         G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358,
         G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422,
         G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545,
         G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694,
         G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724,
         G4087, G4088, G4089, G4090, G4091, G4092, G4115, KEYINPUT0, KEYINPUT1,
         KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
         KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
         KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
         KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
         KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
         KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33,
         KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
         KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
         KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
         KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
         KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
         KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63,
         KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
         KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73,
         KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78,
         KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
         KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
         KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
         KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
         KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
         KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
         KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
         KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
         KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
         KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
         G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926,
         G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939,
         G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598,
         G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629,
         G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873,
         G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757,
         G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696,
         G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865,
         G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645,
         G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807,
         G658, G690;

  wire   n4175, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541;

  NOR2_X2 U2946 ( .A1(n4202), .A2(G4091), .ZN(n4504) );
  NOR2_X2 U2947 ( .A1(G4091), .A2(G4092), .ZN(n4255) );
  INV_X1 U2948 ( .A(G1), .ZN(n4175) );
  INV_X1 U2949 ( .A(n4175), .ZN(G939) );
  INV_X1 U2950 ( .A(n4175), .ZN(G921) );
  INV_X1 U2951 ( .A(n4175), .ZN(G949) );
  INV_X1 U2952 ( .A(n4175), .ZN(G993) );
  INV_X1 U2953 ( .A(n4175), .ZN(G978) );
  BUF_X1 U2954 ( .A(G137), .Z(G926) );
  BUF_X1 U2955 ( .A(G141), .Z(G923) );
  BUF_X1 U2956 ( .A(G141), .Z(G144) );
  BUF_X1 U2957 ( .A(G293), .Z(G298) );
  BUF_X1 U2958 ( .A(G299), .Z(G889) );
  BUF_X1 U2959 ( .A(G299), .Z(G887) );
  BUF_X1 U2960 ( .A(G549), .Z(G892) );
  BUF_X1 U2961 ( .A(G3173), .Z(G973) );
  BUF_X1 U2962 ( .A(G594), .Z(G604) );
  BUF_X1 U2963 ( .A(G594), .Z(G603) );
  BUF_X1 U2964 ( .A(G606), .Z(G602) );
  BUF_X1 U2965 ( .A(G717), .Z(G704) );
  NAND3_X1 U2966 ( .A1(n4193), .A2(n4194), .A3(n4195), .ZN(G882) );
  NAND2_X1 U2967 ( .A1(G4092), .A2(G118), .ZN(n4195) );
  NAND3_X1 U2968 ( .A1(n4196), .A2(n4197), .A3(n4198), .ZN(n4194) );
  INV_X1 U2969 ( .A(KEYINPUT48), .ZN(n4197) );
  NAND2_X1 U2970 ( .A1(n4199), .A2(n4200), .ZN(n4193) );
  NAND3_X1 U2971 ( .A1(n4201), .A2(n4202), .A3(n4203), .ZN(n4200) );
  NAND2_X1 U2972 ( .A1(KEYINPUT48), .A2(n4196), .ZN(n4201) );
  XNOR2_X1 U2973 ( .A(KEYINPUT104), .B(n4204), .ZN(G875) );
  NAND4_X1 U2974 ( .A1(n4205), .A2(n4206), .A3(n4207), .A4(n4208), .ZN(G859) );
  NAND2_X1 U2975 ( .A1(G11), .A2(n4209), .ZN(n4208) );
  NAND2_X1 U2976 ( .A1(n4210), .A2(n4211), .ZN(n4207) );
  NAND2_X1 U2977 ( .A1(n4212), .A2(n4213), .ZN(n4206) );
  XOR2_X1 U2978 ( .A(n4214), .B(KEYINPUT57), .Z(n4205) );
  NAND2_X1 U2979 ( .A1(G61), .A2(n4215), .ZN(n4214) );
  NOR4_X1 U2980 ( .A1(n4216), .A2(n4217), .A3(G1002), .A4(G1000), .ZN(G854) );
  OR3_X1 U2981 ( .A1(G848), .A2(G851), .A3(G998), .ZN(n4217) );
  XOR2_X1 U2982 ( .A(n4218), .B(n4219), .Z(G998) );
  NOR4_X1 U2983 ( .A1(n4220), .A2(n4221), .A3(n4222), .A4(n4223), .ZN(n4219) );
  NOR3_X1 U2984 ( .A1(n4224), .A2(n4225), .A3(n4226), .ZN(n4223) );
  NOR3_X1 U2985 ( .A1(n4227), .A2(n4226), .A3(n4228), .ZN(n4222) );
  INV_X1 U2986 ( .A(n4229), .ZN(n4226) );
  NOR3_X1 U2987 ( .A1(n4227), .A2(n4225), .A3(n4229), .ZN(n4221) );
  INV_X1 U2988 ( .A(n4224), .ZN(n4227) );
  NOR3_X1 U2989 ( .A1(n4224), .A2(n4229), .A3(n4228), .ZN(n4220) );
  INV_X1 U2990 ( .A(n4225), .ZN(n4228) );
  XOR2_X1 U2991 ( .A(n4230), .B(n4231), .Z(n4225) );
  XNOR2_X1 U2992 ( .A(n4232), .B(n4233), .ZN(n4229) );
  XOR2_X1 U2993 ( .A(n4234), .B(n4235), .Z(n4224) );
  NAND2_X1 U2994 ( .A1(n4236), .A2(n4237), .ZN(n4234) );
  NAND2_X1 U2995 ( .A1(G369), .A2(n4238), .ZN(n4237) );
  NAND2_X1 U2996 ( .A1(G372), .A2(G332), .ZN(n4236) );
  NAND2_X1 U2997 ( .A1(KEYINPUT38), .A2(n4239), .ZN(n4218) );
  XOR2_X1 U2998 ( .A(n4240), .B(n4241), .Z(n4239) );
  XNOR2_X1 U2999 ( .A(n4242), .B(n4243), .ZN(n4241) );
  XNOR2_X1 U3000 ( .A(n4244), .B(n4245), .ZN(n4240) );
  NOR2_X1 U3001 ( .A1(KEYINPUT52), .A2(n4246), .ZN(n4245) );
  NAND4_X1 U3002 ( .A1(G556), .A2(G386), .A3(G601), .A4(n4247), .ZN(n4216) );
  INV_X1 U3003 ( .A(G559), .ZN(G851) );
  INV_X1 U3004 ( .A(G245), .ZN(G848) );
  NAND2_X1 U3005 ( .A1(n4248), .A2(G386), .ZN(G847) );
  XNOR2_X1 U3006 ( .A(G556), .B(KEYINPUT95), .ZN(n4248) );
  NAND2_X1 U3007 ( .A1(n4249), .A2(G27), .ZN(G845) );
  INV_X1 U3008 ( .A(G2824), .ZN(n4249) );
  NAND3_X1 U3009 ( .A1(n4250), .A2(n4251), .A3(n4252), .ZN(G843) );
  NAND2_X1 U3010 ( .A1(G4091), .A2(n4253), .ZN(n4252) );
  NAND2_X1 U3011 ( .A1(n4254), .A2(n4255), .ZN(n4251) );
  XNOR2_X1 U3012 ( .A(n4256), .B(n4257), .ZN(n4254) );
  OR2_X1 U3013 ( .A1(n4258), .A2(n4202), .ZN(n4250) );
  NOR2_X1 U3014 ( .A1(G120), .A2(G4091), .ZN(n4258) );
  NAND2_X1 U3015 ( .A1(G83), .A2(n4259), .ZN(G820) );
  AND3_X1 U3016 ( .A1(n4260), .A2(n4261), .A3(n4262), .ZN(G818) );
  NAND2_X1 U3017 ( .A1(G4115), .A2(G135), .ZN(n4262) );
  NAND2_X1 U3018 ( .A1(n4263), .A2(n4264), .ZN(n4261) );
  INV_X1 U3019 ( .A(G3724), .ZN(n4264) );
  NAND2_X1 U3020 ( .A1(n4265), .A2(n4266), .ZN(n4263) );
  OR2_X1 U3021 ( .A1(n4267), .A2(G123), .ZN(n4266) );
  NAND2_X1 U3022 ( .A1(n4268), .A2(n4267), .ZN(n4265) );
  NAND2_X1 U3023 ( .A1(n4269), .A2(n4270), .ZN(n4268) );
  INV_X1 U3024 ( .A(KEYINPUT58), .ZN(n4270) );
  NAND2_X1 U3025 ( .A1(G3724), .A2(n4271), .ZN(n4260) );
  NAND2_X1 U3026 ( .A1(n4272), .A2(n4273), .ZN(n4271) );
  NAND2_X1 U3027 ( .A1(G3717), .A2(G623), .ZN(n4273) );
  NAND3_X1 U3028 ( .A1(n4274), .A2(n4275), .A3(n4267), .ZN(n4272) );
  INV_X1 U3029 ( .A(G3717), .ZN(n4267) );
  NAND2_X1 U3030 ( .A1(KEYINPUT58), .A2(n4269), .ZN(n4275) );
  XNOR2_X1 U3031 ( .A(n4246), .B(G132), .ZN(n4274) );
  NOR2_X1 U3032 ( .A1(G3173), .A2(n4276), .ZN(G815) );
  INV_X1 U3033 ( .A(G136), .ZN(n4276) );
  XOR2_X1 U3034 ( .A(n4277), .B(G132), .Z(G813) );
  AND2_X1 U3035 ( .A1(G141), .A2(G145), .ZN(G810) );
  NAND4_X1 U3036 ( .A1(n4278), .A2(n4279), .A3(n4280), .A4(n4281), .ZN(G807) );
  NAND2_X1 U3037 ( .A1(G64), .A2(n4215), .ZN(n4281) );
  NAND2_X1 U3038 ( .A1(G14), .A2(n4209), .ZN(n4280) );
  NAND2_X1 U3039 ( .A1(n4210), .A2(n4282), .ZN(n4279) );
  NAND2_X1 U3040 ( .A1(n4212), .A2(n4283), .ZN(n4278) );
  NAND4_X1 U3041 ( .A1(n4284), .A2(n4285), .A3(n4286), .A4(n4287), .ZN(G802) );
  NAND2_X1 U3042 ( .A1(G70), .A2(n4215), .ZN(n4287) );
  NAND2_X1 U3043 ( .A1(G67), .A2(n4209), .ZN(n4286) );
  NAND2_X1 U3044 ( .A1(n4210), .A2(n4288), .ZN(n4285) );
  NAND2_X1 U3045 ( .A1(n4212), .A2(n4289), .ZN(n4284) );
  NAND4_X1 U3046 ( .A1(n4290), .A2(n4291), .A3(n4292), .A4(n4293), .ZN(G797) );
  NAND2_X1 U3047 ( .A1(G17), .A2(n4215), .ZN(n4293) );
  NAND2_X1 U3048 ( .A1(G73), .A2(n4209), .ZN(n4292) );
  NAND2_X1 U3049 ( .A1(n4210), .A2(n4294), .ZN(n4291) );
  NAND2_X1 U3050 ( .A1(n4212), .A2(n4204), .ZN(n4290) );
  NAND4_X1 U3051 ( .A1(n4295), .A2(n4296), .A3(n4297), .A4(n4298), .ZN(G792) );
  NAND2_X1 U3052 ( .A1(G20), .A2(n4215), .ZN(n4298) );
  NOR2_X1 U3053 ( .A1(n4299), .A2(n4300), .ZN(n4215) );
  NAND2_X1 U3054 ( .A1(G76), .A2(n4209), .ZN(n4297) );
  NOR2_X1 U3055 ( .A1(n4300), .A2(G4089), .ZN(n4209) );
  NAND2_X1 U3056 ( .A1(n4210), .A2(n4301), .ZN(n4296) );
  NOR2_X1 U3057 ( .A1(n4302), .A2(G4089), .ZN(n4210) );
  NAND2_X1 U3058 ( .A1(n4212), .A2(n4303), .ZN(n4295) );
  NOR2_X1 U3059 ( .A1(n4299), .A2(n4302), .ZN(n4212) );
  INV_X1 U3060 ( .A(n4300), .ZN(n4302) );
  XOR2_X1 U3061 ( .A(G4090), .B(KEYINPUT83), .Z(n4300) );
  NAND4_X1 U3062 ( .A1(n4304), .A2(n4305), .A3(n4306), .A4(n4307), .ZN(G787) );
  NAND2_X1 U3063 ( .A1(G43), .A2(n4308), .ZN(n4307) );
  NAND2_X1 U3064 ( .A1(n4309), .A2(n4310), .ZN(n4306) );
  NAND2_X1 U3065 ( .A1(n4311), .A2(n4312), .ZN(n4305) );
  NAND2_X1 U3066 ( .A1(G37), .A2(n4313), .ZN(n4304) );
  NAND4_X1 U3067 ( .A1(n4314), .A2(n4315), .A3(n4316), .A4(n4317), .ZN(G782) );
  NAND2_X1 U3068 ( .A1(G91), .A2(n4308), .ZN(n4317) );
  NAND2_X1 U3069 ( .A1(n4309), .A2(n4318), .ZN(n4316) );
  NAND2_X1 U3070 ( .A1(n4311), .A2(n4319), .ZN(n4315) );
  NAND2_X1 U3071 ( .A1(G40), .A2(n4313), .ZN(n4314) );
  NAND4_X1 U3072 ( .A1(n4320), .A2(n4321), .A3(n4322), .A4(n4323), .ZN(G777) );
  NAND2_X1 U3073 ( .A1(n4309), .A2(n4324), .ZN(n4323) );
  NAND2_X1 U3074 ( .A1(n4311), .A2(n4325), .ZN(n4322) );
  NAND2_X1 U3075 ( .A1(G103), .A2(n4313), .ZN(n4321) );
  XOR2_X1 U3076 ( .A(n4326), .B(KEYINPUT99), .Z(n4320) );
  NAND2_X1 U3077 ( .A1(G100), .A2(n4308), .ZN(n4326) );
  NAND4_X1 U3078 ( .A1(n4327), .A2(n4328), .A3(n4329), .A4(n4330), .ZN(G772) );
  NAND2_X1 U3079 ( .A1(n4311), .A2(n4331), .ZN(n4330) );
  XNOR2_X1 U3080 ( .A(KEYINPUT67), .B(n4332), .ZN(n4331) );
  NAND2_X1 U3081 ( .A1(G46), .A2(n4308), .ZN(n4329) );
  NAND2_X1 U3082 ( .A1(n4309), .A2(n4333), .ZN(n4328) );
  NAND2_X1 U3083 ( .A1(G49), .A2(n4313), .ZN(n4327) );
  NAND4_X1 U3084 ( .A1(n4334), .A2(n4335), .A3(n4336), .A4(n4337), .ZN(G767) );
  NAND2_X1 U3085 ( .A1(n4338), .A2(n4282), .ZN(n4337) );
  NAND2_X1 U3086 ( .A1(n4339), .A2(G14), .ZN(n4336) );
  NAND2_X1 U3087 ( .A1(n4340), .A2(n4283), .ZN(n4335) );
  NAND2_X1 U3088 ( .A1(n4341), .A2(G64), .ZN(n4334) );
  NAND4_X1 U3089 ( .A1(n4342), .A2(n4343), .A3(n4344), .A4(n4345), .ZN(G762) );
  NAND2_X1 U3090 ( .A1(n4338), .A2(n4288), .ZN(n4345) );
  NAND2_X1 U3091 ( .A1(n4339), .A2(G67), .ZN(n4344) );
  NAND2_X1 U3092 ( .A1(n4340), .A2(n4289), .ZN(n4343) );
  NAND2_X1 U3093 ( .A1(n4341), .A2(G70), .ZN(n4342) );
  NAND3_X1 U3094 ( .A1(n4346), .A2(n4347), .A3(n4348), .ZN(G757) );
  NAND2_X1 U3095 ( .A1(n4340), .A2(n4204), .ZN(n4348) );
  NAND3_X1 U3096 ( .A1(G17), .A2(n4349), .A3(n4341), .ZN(n4347) );
  INV_X1 U3097 ( .A(KEYINPUT103), .ZN(n4349) );
  NAND3_X1 U3098 ( .A1(n4350), .A2(n4351), .A3(n4352), .ZN(n4346) );
  NAND2_X1 U3099 ( .A1(G836), .A2(n4353), .ZN(n4351) );
  NAND3_X1 U3100 ( .A1(n4354), .A2(n4355), .A3(G4087), .ZN(n4350) );
  INV_X1 U3101 ( .A(G73), .ZN(n4355) );
  NAND2_X1 U3102 ( .A1(KEYINPUT103), .A2(G17), .ZN(n4354) );
  NAND4_X1 U3103 ( .A1(n4356), .A2(n4357), .A3(n4358), .A4(n4359), .ZN(G752) );
  NAND2_X1 U3104 ( .A1(n4338), .A2(n4301), .ZN(n4359) );
  NAND2_X1 U3105 ( .A1(n4339), .A2(G76), .ZN(n4358) );
  NAND2_X1 U3106 ( .A1(n4340), .A2(n4303), .ZN(n4357) );
  NAND2_X1 U3107 ( .A1(n4341), .A2(G20), .ZN(n4356) );
  NAND4_X1 U3108 ( .A1(n4360), .A2(n4361), .A3(n4362), .A4(n4363), .ZN(G747) );
  NAND2_X1 U3109 ( .A1(n4364), .A2(G43), .ZN(n4363) );
  NAND2_X1 U3110 ( .A1(n4365), .A2(n4312), .ZN(n4362) );
  NAND2_X1 U3111 ( .A1(n4366), .A2(G37), .ZN(n4361) );
  XOR2_X1 U3112 ( .A(KEYINPUT73), .B(n4367), .Z(n4360) );
  AND2_X1 U3113 ( .A1(n4310), .A2(n4368), .ZN(n4367) );
  NAND4_X1 U3114 ( .A1(n4369), .A2(n4370), .A3(n4371), .A4(n4372), .ZN(G742) );
  NAND2_X1 U3115 ( .A1(n4368), .A2(n4373), .ZN(n4372) );
  XNOR2_X1 U3116 ( .A(KEYINPUT49), .B(n4318), .ZN(n4373) );
  NAND2_X1 U3117 ( .A1(n4364), .A2(G91), .ZN(n4371) );
  NAND2_X1 U3118 ( .A1(n4365), .A2(n4319), .ZN(n4370) );
  NAND2_X1 U3119 ( .A1(n4366), .A2(G40), .ZN(n4369) );
  NAND4_X1 U3120 ( .A1(n4374), .A2(n4375), .A3(n4376), .A4(n4377), .ZN(G737) );
  NAND2_X1 U3121 ( .A1(n4368), .A2(n4324), .ZN(n4377) );
  NAND2_X1 U3122 ( .A1(n4364), .A2(G100), .ZN(n4376) );
  NAND2_X1 U3123 ( .A1(n4365), .A2(n4325), .ZN(n4375) );
  NAND2_X1 U3124 ( .A1(n4366), .A2(G103), .ZN(n4374) );
  NAND4_X1 U3125 ( .A1(n4378), .A2(n4379), .A3(n4380), .A4(n4381), .ZN(G732) );
  NAND2_X1 U3126 ( .A1(n4368), .A2(n4333), .ZN(n4381) );
  NAND2_X1 U3127 ( .A1(n4364), .A2(G46), .ZN(n4380) );
  NAND2_X1 U3128 ( .A1(n4365), .A2(n4332), .ZN(n4379) );
  NAND2_X1 U3129 ( .A1(n4366), .A2(G49), .ZN(n4378) );
  NAND4_X1 U3130 ( .A1(n4382), .A2(n4383), .A3(n4384), .A4(n4385), .ZN(G727) );
  NAND2_X1 U3131 ( .A1(n4368), .A2(n4386), .ZN(n4385) );
  NOR2_X1 U3132 ( .A1(n4387), .A2(G4088), .ZN(n4368) );
  NAND2_X1 U3133 ( .A1(G109), .A2(n4364), .ZN(n4384) );
  NOR2_X1 U3134 ( .A1(n4388), .A2(G4088), .ZN(n4364) );
  NAND2_X1 U3135 ( .A1(n4365), .A2(n4389), .ZN(n4383) );
  NOR2_X1 U3136 ( .A1(n4387), .A2(n4352), .ZN(n4365) );
  NAND2_X1 U3137 ( .A1(G106), .A2(n4366), .ZN(n4382) );
  NOR2_X1 U3138 ( .A1(n4352), .A2(n4388), .ZN(n4366) );
  INV_X1 U3139 ( .A(n4387), .ZN(n4388) );
  XOR2_X1 U3140 ( .A(G4087), .B(KEYINPUT20), .Z(n4387) );
  NAND4_X1 U3141 ( .A1(n4390), .A2(n4391), .A3(n4392), .A4(n4393), .ZN(G722) );
  NAND2_X1 U3142 ( .A1(n4338), .A2(n4211), .ZN(n4393) );
  NOR2_X1 U3143 ( .A1(G4087), .A2(G4088), .ZN(n4338) );
  NAND2_X1 U3144 ( .A1(n4339), .A2(G11), .ZN(n4392) );
  NOR2_X1 U3145 ( .A1(n4353), .A2(G4088), .ZN(n4339) );
  NAND2_X1 U3146 ( .A1(n4340), .A2(n4213), .ZN(n4391) );
  NOR2_X1 U3147 ( .A1(n4352), .A2(G4087), .ZN(n4340) );
  NAND2_X1 U3148 ( .A1(n4341), .A2(G61), .ZN(n4390) );
  NOR2_X1 U3149 ( .A1(n4352), .A2(n4353), .ZN(n4341) );
  INV_X1 U3150 ( .A(G4087), .ZN(n4353) );
  INV_X1 U3151 ( .A(G4088), .ZN(n4352) );
  OR3_X1 U3152 ( .A1(n4394), .A2(n4395), .A3(G809), .ZN(G717) );
  NOR2_X1 U3153 ( .A1(G88), .A2(G2358), .ZN(n4395) );
  NOR2_X1 U3154 ( .A1(G34), .A2(n4396), .ZN(n4394) );
  AND2_X1 U3155 ( .A1(G141), .A2(n4397), .ZN(G715) );
  NAND3_X1 U3156 ( .A1(n4398), .A2(n4399), .A3(n4259), .ZN(n4397) );
  NAND2_X1 U3157 ( .A1(G82), .A2(n4396), .ZN(n4399) );
  NAND2_X1 U3158 ( .A1(G80), .A2(G2358), .ZN(n4398) );
  NAND4_X1 U3159 ( .A1(n4400), .A2(n4401), .A3(n4402), .A4(n4403), .ZN(G712) );
  NAND2_X1 U3160 ( .A1(G109), .A2(n4308), .ZN(n4403) );
  NOR2_X1 U3161 ( .A1(n4404), .A2(G4089), .ZN(n4308) );
  NAND2_X1 U3162 ( .A1(n4309), .A2(n4386), .ZN(n4402) );
  NOR2_X1 U3163 ( .A1(G4089), .A2(G4090), .ZN(n4309) );
  NAND2_X1 U3164 ( .A1(n4311), .A2(n4389), .ZN(n4401) );
  NOR2_X1 U3165 ( .A1(n4299), .A2(G4090), .ZN(n4311) );
  NAND2_X1 U3166 ( .A1(G106), .A2(n4313), .ZN(n4400) );
  NOR2_X1 U3167 ( .A1(n4299), .A2(n4404), .ZN(n4313) );
  INV_X1 U3168 ( .A(G4090), .ZN(n4404) );
  INV_X1 U3169 ( .A(G4089), .ZN(n4299) );
  AND2_X1 U3170 ( .A1(G141), .A2(n4405), .ZN(G707) );
  NAND3_X1 U3171 ( .A1(n4406), .A2(n4407), .A3(n4259), .ZN(n4405) );
  NAND2_X1 U3172 ( .A1(G79), .A2(n4396), .ZN(n4407) );
  NAND2_X1 U3173 ( .A1(G23), .A2(G2358), .ZN(n4406) );
  NOR2_X1 U3174 ( .A1(n4408), .A2(n4409), .ZN(G702) );
  XNOR2_X1 U3175 ( .A(KEYINPUT53), .B(n4410), .ZN(n4409) );
  NOR4_X1 U3176 ( .A1(n4411), .A2(n4412), .A3(n4413), .A4(n4414), .ZN(n4408) );
  NOR2_X1 U3177 ( .A1(G834), .A2(n4415), .ZN(n4414) );
  INV_X1 U3178 ( .A(n4301), .ZN(G834) );
  NOR2_X1 U3179 ( .A1(G873), .A2(n4416), .ZN(n4413) );
  INV_X1 U3180 ( .A(n4303), .ZN(G873) );
  AND2_X1 U3181 ( .A1(n4417), .A2(G149), .ZN(n4412) );
  NOR2_X1 U3182 ( .A1(n4418), .A2(n4419), .ZN(n4411) );
  INV_X1 U3183 ( .A(G146), .ZN(n4419) );
  NOR2_X1 U3184 ( .A1(n4420), .A2(n4421), .ZN(G699) );
  NOR4_X1 U3185 ( .A1(n4422), .A2(n4423), .A3(n4424), .A4(n4425), .ZN(n4420) );
  NOR2_X1 U3186 ( .A1(G836), .A2(n4415), .ZN(n4425) );
  INV_X1 U3187 ( .A(n4294), .ZN(G836) );
  NOR2_X1 U3188 ( .A1(n4426), .A2(n4416), .ZN(n4424) );
  INV_X1 U3189 ( .A(n4204), .ZN(n4426) );
  AND2_X1 U3190 ( .A1(n4417), .A2(G155), .ZN(n4423) );
  NOR2_X1 U3191 ( .A1(n4418), .A2(n4427), .ZN(n4422) );
  INV_X1 U3192 ( .A(G152), .ZN(n4427) );
  NOR2_X1 U3193 ( .A1(n4428), .A2(n4421), .ZN(G696) );
  NOR4_X1 U3194 ( .A1(n4429), .A2(n4430), .A3(n4431), .A4(n4432), .ZN(n4428) );
  NOR2_X1 U3195 ( .A1(G838), .A2(n4415), .ZN(n4432) );
  NOR2_X1 U3196 ( .A1(G877), .A2(n4416), .ZN(n4431) );
  INV_X1 U3197 ( .A(n4289), .ZN(G877) );
  AND2_X1 U3198 ( .A1(n4417), .A2(G188), .ZN(n4430) );
  NOR2_X1 U3199 ( .A1(n4418), .A2(n4433), .ZN(n4429) );
  INV_X1 U3200 ( .A(G158), .ZN(n4433) );
  NOR2_X1 U3201 ( .A1(n4434), .A2(n4421), .ZN(G693) );
  NOR4_X1 U3202 ( .A1(n4435), .A2(n4436), .A3(n4437), .A4(n4438), .ZN(n4434) );
  NOR2_X1 U3203 ( .A1(G822), .A2(n4415), .ZN(n4438) );
  INV_X1 U3204 ( .A(n4211), .ZN(G822) );
  NOR2_X1 U3205 ( .A1(G861), .A2(n4416), .ZN(n4437) );
  INV_X1 U3206 ( .A(n4213), .ZN(G861) );
  AND2_X1 U3207 ( .A1(n4417), .A2(G182), .ZN(n4436) );
  NOR2_X1 U3208 ( .A1(n4418), .A2(n4439), .ZN(n4435) );
  INV_X1 U3209 ( .A(G185), .ZN(n4439) );
  NAND3_X1 U3210 ( .A1(n4410), .A2(n4440), .A3(n4441), .ZN(G690) );
  NOR3_X1 U3211 ( .A1(n4442), .A2(n4443), .A3(n4444), .ZN(n4441) );
  NOR2_X1 U3212 ( .A1(G176), .A2(n4445), .ZN(n4444) );
  NOR2_X1 U3213 ( .A1(G179), .A2(n4418), .ZN(n4443) );
  NOR2_X1 U3214 ( .A1(n4416), .A2(n4283), .ZN(n4442) );
  NAND2_X1 U3215 ( .A1(n4446), .A2(n4447), .ZN(n4440) );
  INV_X1 U3216 ( .A(n4421), .ZN(n4410) );
  XOR2_X1 U3217 ( .A(G137), .B(KEYINPUT127), .Z(n4421) );
  NOR2_X1 U3218 ( .A1(n4448), .A2(n4449), .ZN(G688) );
  NOR4_X1 U3219 ( .A1(n4450), .A2(n4451), .A3(n4452), .A4(n4453), .ZN(n4448) );
  NOR2_X1 U3220 ( .A1(G863), .A2(n4416), .ZN(n4453) );
  INV_X1 U3221 ( .A(n4389), .ZN(G863) );
  AND2_X1 U3222 ( .A1(n4417), .A2(G191), .ZN(n4452) );
  NOR2_X1 U3223 ( .A1(n4418), .A2(n4454), .ZN(n4451) );
  INV_X1 U3224 ( .A(G161), .ZN(n4454) );
  NOR3_X1 U3225 ( .A1(G824), .A2(n4455), .A3(n4456), .ZN(n4450) );
  AND2_X1 U3226 ( .A1(n4416), .A2(KEYINPUT54), .ZN(n4456) );
  NOR2_X1 U3227 ( .A1(KEYINPUT54), .A2(n4447), .ZN(n4455) );
  INV_X1 U3228 ( .A(n4386), .ZN(G824) );
  NOR2_X1 U3229 ( .A1(n4457), .A2(n4449), .ZN(G685) );
  NOR4_X1 U3230 ( .A1(n4458), .A2(n4459), .A3(n4460), .A4(n4461), .ZN(n4457) );
  NOR2_X1 U3231 ( .A1(G865), .A2(n4416), .ZN(n4461) );
  NOR2_X1 U3232 ( .A1(n4445), .A2(n4462), .ZN(n4460) );
  NOR2_X1 U3233 ( .A1(n4418), .A2(n4463), .ZN(n4459) );
  NOR3_X1 U3234 ( .A1(G826), .A2(n4464), .A3(n4465), .ZN(n4458) );
  NOR2_X1 U3235 ( .A1(KEYINPUT108), .A2(n4417), .ZN(n4465) );
  AND2_X1 U3236 ( .A1(n4415), .A2(KEYINPUT108), .ZN(n4464) );
  NOR2_X1 U3237 ( .A1(n4466), .A2(n4449), .ZN(G682) );
  NOR4_X1 U3238 ( .A1(n4467), .A2(n4468), .A3(n4469), .A4(n4470), .ZN(n4466) );
  NOR2_X1 U3239 ( .A1(G828), .A2(n4415), .ZN(n4470) );
  NOR2_X1 U3240 ( .A1(G867), .A2(n4416), .ZN(n4469) );
  INV_X1 U3241 ( .A(n4325), .ZN(G867) );
  AND2_X1 U3242 ( .A1(n4417), .A2(G197), .ZN(n4468) );
  NOR2_X1 U3243 ( .A1(n4418), .A2(n4471), .ZN(n4467) );
  INV_X1 U3244 ( .A(G167), .ZN(n4471) );
  NOR2_X1 U3245 ( .A1(n4472), .A2(n4449), .ZN(G679) );
  NOR4_X1 U3246 ( .A1(n4473), .A2(n4474), .A3(n4475), .A4(n4476), .ZN(n4472) );
  NOR2_X1 U3247 ( .A1(G830), .A2(n4415), .ZN(n4476) );
  INV_X1 U3248 ( .A(n4318), .ZN(G830) );
  NOR2_X1 U3249 ( .A1(G869), .A2(n4416), .ZN(n4475) );
  INV_X1 U3250 ( .A(n4319), .ZN(G869) );
  AND2_X1 U3251 ( .A1(n4417), .A2(G203), .ZN(n4474) );
  NOR2_X1 U3252 ( .A1(n4418), .A2(n4477), .ZN(n4473) );
  INV_X1 U3253 ( .A(G173), .ZN(n4477) );
  NOR2_X1 U3254 ( .A1(n4478), .A2(n4449), .ZN(G676) );
  NOR4_X1 U3255 ( .A1(n4479), .A2(n4480), .A3(n4481), .A4(n4482), .ZN(n4478) );
  NOR2_X1 U3256 ( .A1(G832), .A2(n4415), .ZN(n4482) );
  INV_X1 U3257 ( .A(n4447), .ZN(n4415) );
  NOR2_X1 U3258 ( .A1(G1691), .A2(G1694), .ZN(n4447) );
  INV_X1 U3259 ( .A(n4310), .ZN(G832) );
  NOR2_X1 U3260 ( .A1(G871), .A2(n4416), .ZN(n4481) );
  OR2_X1 U3261 ( .A1(n4483), .A2(G1694), .ZN(n4416) );
  INV_X1 U3262 ( .A(n4312), .ZN(G871) );
  AND2_X1 U3263 ( .A1(n4417), .A2(G200), .ZN(n4480) );
  INV_X1 U3264 ( .A(n4445), .ZN(n4417) );
  NAND2_X1 U3265 ( .A1(G1694), .A2(n4483), .ZN(n4445) );
  INV_X1 U3266 ( .A(G1691), .ZN(n4483) );
  NOR2_X1 U3267 ( .A1(n4418), .A2(n4484), .ZN(n4479) );
  INV_X1 U3268 ( .A(G170), .ZN(n4484) );
  NAND2_X1 U3269 ( .A1(G1694), .A2(G1691), .ZN(n4418) );
  AND2_X1 U3270 ( .A1(G141), .A2(n4485), .ZN(G673) );
  NAND3_X1 U3271 ( .A1(n4486), .A2(n4487), .A3(n4259), .ZN(n4485) );
  NAND2_X1 U3272 ( .A1(G26), .A2(n4396), .ZN(n4487) );
  NAND2_X1 U3273 ( .A1(G81), .A2(G2358), .ZN(n4486) );
  NAND4_X1 U3274 ( .A1(n4488), .A2(n4489), .A3(n4490), .A4(n4491), .ZN(G670) );
  NAND2_X1 U3275 ( .A1(n4492), .A2(n4303), .ZN(n4491) );
  NAND3_X1 U3276 ( .A1(n4493), .A2(n4494), .A3(n4495), .ZN(n4303) );
  NAND2_X1 U3277 ( .A1(n4496), .A2(n4198), .ZN(n4495) );
  NAND2_X1 U3278 ( .A1(n4497), .A2(n4498), .ZN(n4494) );
  NAND2_X1 U3279 ( .A1(G128), .A2(n4499), .ZN(n4493) );
  NAND2_X1 U3280 ( .A1(n4500), .A2(n4301), .ZN(n4490) );
  NAND3_X1 U3281 ( .A1(n4501), .A2(n4502), .A3(n4503), .ZN(n4301) );
  NAND2_X1 U3282 ( .A1(G130), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U3283 ( .A1(n4255), .A2(n4505), .ZN(n4502) );
  NAND2_X1 U3284 ( .A1(n4506), .A2(n4507), .ZN(n4501) );
  NAND2_X1 U3285 ( .A1(n4508), .A2(G149), .ZN(n4489) );
  NAND2_X1 U3286 ( .A1(n4509), .A2(G146), .ZN(n4488) );
  NAND4_X1 U3287 ( .A1(n4510), .A2(n4511), .A3(n4512), .A4(n4513), .ZN(G667) );
  NOR2_X1 U3288 ( .A1(n4514), .A2(n4515), .ZN(n4513) );
  AND2_X1 U3289 ( .A1(G155), .A2(n4508), .ZN(n4515) );
  AND2_X1 U3290 ( .A1(n4204), .A2(n4492), .ZN(n4514) );
  NAND3_X1 U3291 ( .A1(n4516), .A2(n4517), .A3(n4518), .ZN(n4204) );
  NAND2_X1 U3292 ( .A1(n4519), .A2(n4198), .ZN(n4518) );
  INV_X1 U3293 ( .A(n4520), .ZN(n4519) );
  NAND2_X1 U3294 ( .A1(n4521), .A2(n4497), .ZN(n4517) );
  NAND2_X1 U3295 ( .A1(G127), .A2(n4499), .ZN(n4516) );
  NAND2_X1 U3296 ( .A1(n4509), .A2(G152), .ZN(n4512) );
  NAND3_X1 U3297 ( .A1(G137), .A2(n4522), .A3(n4523), .ZN(n4511) );
  INV_X1 U3298 ( .A(KEYINPUT10), .ZN(n4523) );
  NAND2_X1 U3299 ( .A1(n4524), .A2(n4294), .ZN(n4522) );
  NAND3_X1 U3300 ( .A1(n4500), .A2(n4294), .A3(KEYINPUT10), .ZN(n4510) );
  NAND3_X1 U3301 ( .A1(n4525), .A2(n4526), .A3(n4527), .ZN(n4294) );
  NAND2_X1 U3302 ( .A1(n4528), .A2(n4255), .ZN(n4527) );
  NAND2_X1 U3303 ( .A1(n4529), .A2(n4506), .ZN(n4526) );
  NAND2_X1 U3304 ( .A1(G119), .A2(n4504), .ZN(n4525) );
  NAND4_X1 U3305 ( .A1(n4530), .A2(n4531), .A3(n4532), .A4(n4533), .ZN(G664) );
  NAND3_X1 U3306 ( .A1(n4289), .A2(n4534), .A3(n4492), .ZN(n4533) );
  INV_X1 U3307 ( .A(KEYINPUT6), .ZN(n4534) );
  NAND2_X1 U3308 ( .A1(n4500), .A2(n4535), .ZN(n4532) );
  NAND2_X1 U3309 ( .A1(G838), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U3310 ( .A1(KEYINPUT6), .A2(n4289), .ZN(n4536) );
  NAND3_X1 U3311 ( .A1(n4537), .A2(n4538), .A3(n4539), .ZN(n4289) );
  NAND2_X1 U3312 ( .A1(n4540), .A2(n4198), .ZN(n4539) );
  INV_X1 U3313 ( .A(n4541), .ZN(n4540) );
  NAND4_X1 U3314 ( .A1(n4497), .A2(n4542), .A3(n4543), .A4(n4544), .ZN(n4538) );
  NAND2_X1 U3315 ( .A1(G126), .A2(n4499), .ZN(n4537) );
  INV_X1 U3316 ( .A(n4288), .ZN(G838) );
  NAND3_X1 U3317 ( .A1(n4545), .A2(n4546), .A3(n4547), .ZN(n4288) );
  NAND2_X1 U3318 ( .A1(n4506), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U3319 ( .A1(G129), .A2(n4504), .ZN(n4546) );
  NAND2_X1 U3320 ( .A1(n4549), .A2(n4255), .ZN(n4545) );
  NAND2_X1 U3321 ( .A1(n4508), .A2(G188), .ZN(n4531) );
  NAND2_X1 U3322 ( .A1(n4509), .A2(G158), .ZN(n4530) );
  NAND4_X1 U3323 ( .A1(n4550), .A2(n4551), .A3(n4552), .A4(n4553), .ZN(G661) );
  NAND2_X1 U3324 ( .A1(n4492), .A2(n4213), .ZN(n4553) );
  NAND3_X1 U3325 ( .A1(n4554), .A2(n4555), .A3(n4556), .ZN(n4213) );
  NAND2_X1 U3326 ( .A1(n4557), .A2(n4198), .ZN(n4556) );
  NOR2_X1 U3327 ( .A1(n4199), .A2(G4092), .ZN(n4198) );
  INV_X1 U3328 ( .A(n4558), .ZN(n4557) );
  NAND2_X1 U3329 ( .A1(n4497), .A2(n4559), .ZN(n4555) );
  AND2_X1 U3330 ( .A1(n4199), .A2(n4202), .ZN(n4497) );
  NAND2_X1 U3331 ( .A1(G117), .A2(n4499), .ZN(n4554) );
  NOR2_X1 U3332 ( .A1(n4202), .A2(n4199), .ZN(n4499) );
  XOR2_X1 U3333 ( .A(G4091), .B(KEYINPUT126), .Z(n4199) );
  NAND2_X1 U3334 ( .A1(n4500), .A2(n4211), .ZN(n4552) );
  NAND3_X1 U3335 ( .A1(n4560), .A2(n4561), .A3(n4562), .ZN(n4211) );
  NAND2_X1 U3336 ( .A1(n4563), .A2(n4255), .ZN(n4562) );
  NAND2_X1 U3337 ( .A1(n4506), .A2(n4564), .ZN(n4561) );
  NAND2_X1 U3338 ( .A1(G131), .A2(n4504), .ZN(n4560) );
  NAND2_X1 U3339 ( .A1(n4508), .A2(G182), .ZN(n4551) );
  NAND2_X1 U3340 ( .A1(n4509), .A2(G185), .ZN(n4550) );
  NAND4_X1 U3341 ( .A1(n4565), .A2(n4566), .A3(n4567), .A4(n4568), .ZN(G658) );
  NOR2_X1 U3342 ( .A1(n4569), .A2(n4449), .ZN(n4568) );
  NOR2_X1 U3343 ( .A1(G179), .A2(n4570), .ZN(n4569) );
  OR2_X1 U3344 ( .A1(n4571), .A2(n4283), .ZN(n4567) );
  NAND3_X1 U3345 ( .A1(n4572), .A2(n4573), .A3(n4574), .ZN(n4283) );
  NAND2_X1 U3346 ( .A1(G97), .A2(G4092), .ZN(n4574) );
  NAND2_X1 U3347 ( .A1(n4506), .A2(n4203), .ZN(n4573) );
  XOR2_X1 U3348 ( .A(n4575), .B(n4576), .Z(n4203) );
  AND2_X1 U3349 ( .A1(n4577), .A2(n4578), .ZN(n4576) );
  NAND3_X1 U3350 ( .A1(n4579), .A2(n4580), .A3(n4581), .ZN(n4578) );
  XOR2_X1 U3351 ( .A(n4582), .B(n4583), .Z(n4581) );
  NOR3_X1 U3352 ( .A1(n4584), .A2(n4585), .A3(n4586), .ZN(n4583) );
  NOR2_X1 U3353 ( .A1(n4587), .A2(n4588), .ZN(n4586) );
  NOR3_X1 U3354 ( .A1(n4589), .A2(n4590), .A3(n4591), .ZN(n4585) );
  NOR2_X1 U3355 ( .A1(n4592), .A2(n4593), .ZN(n4584) );
  XNOR2_X1 U3356 ( .A(n4590), .B(n4589), .ZN(n4593) );
  XNOR2_X1 U3357 ( .A(n4594), .B(n4595), .ZN(n4582) );
  NAND2_X1 U3358 ( .A1(KEYINPUT23), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U3359 ( .A1(n4597), .A2(KEYINPUT78), .ZN(n4594) );
  XOR2_X1 U3360 ( .A(n4598), .B(n4599), .Z(n4597) );
  NOR3_X1 U3361 ( .A1(n4600), .A2(n4601), .A3(n4602), .ZN(n4599) );
  NAND3_X1 U3362 ( .A1(n4603), .A2(n4604), .A3(n4605), .ZN(n4600) );
  XNOR2_X1 U3363 ( .A(KEYINPUT64), .B(n4606), .ZN(n4605) );
  OR3_X1 U3364 ( .A1(n4607), .A2(n4608), .A3(KEYINPUT116), .ZN(n4604) );
  NAND3_X1 U3365 ( .A1(n4609), .A2(n4608), .A3(KEYINPUT116), .ZN(n4603) );
  INV_X1 U3366 ( .A(n4607), .ZN(n4609) );
  NAND2_X1 U3367 ( .A1(n4610), .A2(KEYINPUT60), .ZN(n4598) );
  XNOR2_X1 U3368 ( .A(n4611), .B(n4612), .ZN(n4610) );
  NOR2_X1 U3369 ( .A1(n4613), .A2(n4614), .ZN(n4612) );
  NAND2_X1 U3370 ( .A1(n4615), .A2(n4616), .ZN(n4580) );
  NAND2_X1 U3371 ( .A1(G1497), .A2(n4617), .ZN(n4616) );
  XNOR2_X1 U3372 ( .A(KEYINPUT5), .B(n4618), .ZN(n4617) );
  NAND3_X1 U3373 ( .A1(KEYINPUT5), .A2(G1497), .A3(n4619), .ZN(n4579) );
  NAND3_X1 U3374 ( .A1(n4620), .A2(n4621), .A3(n4615), .ZN(n4577) );
  INV_X1 U3375 ( .A(n4619), .ZN(n4615) );
  OR2_X1 U3376 ( .A1(n4618), .A2(n4622), .ZN(n4621) );
  XOR2_X1 U3377 ( .A(n4623), .B(n4624), .Z(n4620) );
  XOR2_X1 U3378 ( .A(n4625), .B(n4626), .Z(n4624) );
  XNOR2_X1 U3379 ( .A(n4627), .B(n4628), .ZN(n4626) );
  NOR2_X1 U3380 ( .A1(KEYINPUT97), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U3381 ( .A1(n4630), .A2(n4631), .ZN(n4625) );
  OR2_X1 U3382 ( .A1(n4632), .A2(n4596), .ZN(n4631) );
  NAND3_X1 U3383 ( .A1(n4632), .A2(n4607), .A3(n4596), .ZN(n4630) );
  NOR2_X1 U3384 ( .A1(n4633), .A2(n4601), .ZN(n4632) );
  NOR3_X1 U3385 ( .A1(n4608), .A2(n4591), .A3(n4634), .ZN(n4601) );
  INV_X1 U3386 ( .A(n4606), .ZN(n4633) );
  XNOR2_X1 U3387 ( .A(n4589), .B(n4635), .ZN(n4623) );
  XNOR2_X1 U3388 ( .A(KEYINPUT111), .B(n4614), .ZN(n4635) );
  NAND2_X1 U3389 ( .A1(n4636), .A2(n4637), .ZN(n4575) );
  NAND2_X1 U3390 ( .A1(n4638), .A2(n4622), .ZN(n4637) );
  INV_X1 U3391 ( .A(G1497), .ZN(n4622) );
  NAND2_X1 U3392 ( .A1(n4639), .A2(n4640), .ZN(n4638) );
  NAND3_X1 U3393 ( .A1(n4641), .A2(n4642), .A3(n4643), .ZN(n4640) );
  INV_X1 U3394 ( .A(KEYINPUT42), .ZN(n4643) );
  NAND2_X1 U3395 ( .A1(n4644), .A2(KEYINPUT42), .ZN(n4639) );
  XNOR2_X1 U3396 ( .A(n4642), .B(n4645), .ZN(n4644) );
  XNOR2_X1 U3397 ( .A(n4646), .B(n4647), .ZN(n4642) );
  NAND2_X1 U3398 ( .A1(KEYINPUT63), .A2(n4648), .ZN(n4646) );
  XOR2_X1 U3399 ( .A(n4649), .B(n4650), .Z(n4648) );
  XOR2_X1 U3400 ( .A(n4651), .B(n4652), .Z(n4650) );
  NAND2_X1 U3401 ( .A1(n4653), .A2(n4654), .ZN(n4652) );
  NAND2_X1 U3402 ( .A1(n4655), .A2(n4656), .ZN(n4654) );
  INV_X1 U3403 ( .A(n4657), .ZN(n4655) );
  NAND2_X1 U3404 ( .A1(n4658), .A2(n4657), .ZN(n4653) );
  XNOR2_X1 U3405 ( .A(n4659), .B(n4660), .ZN(n4657) );
  NOR2_X1 U3406 ( .A1(KEYINPUT41), .A2(n4661), .ZN(n4660) );
  XOR2_X1 U3407 ( .A(n4662), .B(n4663), .Z(n4649) );
  NAND2_X1 U3408 ( .A1(n4664), .A2(G1497), .ZN(n4636) );
  XOR2_X1 U3409 ( .A(n4665), .B(n4666), .Z(n4664) );
  XNOR2_X1 U3410 ( .A(n4641), .B(n4667), .ZN(n4666) );
  NAND2_X1 U3411 ( .A1(n4668), .A2(n4669), .ZN(n4667) );
  NAND2_X1 U3412 ( .A1(n4670), .A2(n4656), .ZN(n4669) );
  NAND2_X1 U3413 ( .A1(n4671), .A2(n4672), .ZN(n4656) );
  NAND2_X1 U3414 ( .A1(n4673), .A2(n4674), .ZN(n4672) );
  INV_X1 U3415 ( .A(n4675), .ZN(n4670) );
  NAND2_X1 U3416 ( .A1(n4658), .A2(n4675), .ZN(n4668) );
  NAND3_X1 U3417 ( .A1(n4676), .A2(n4677), .A3(n4678), .ZN(n4675) );
  NAND2_X1 U3418 ( .A1(n4679), .A2(n4680), .ZN(n4678) );
  OR3_X1 U3419 ( .A1(n4680), .A2(n4679), .A3(KEYINPUT32), .ZN(n4677) );
  XNOR2_X1 U3420 ( .A(n4681), .B(n4682), .ZN(n4679) );
  NOR2_X1 U3421 ( .A1(n4683), .A2(n4662), .ZN(n4682) );
  NAND2_X1 U3422 ( .A1(n4684), .A2(KEYINPUT31), .ZN(n4681) );
  XOR2_X1 U3423 ( .A(n4685), .B(n4686), .Z(n4684) );
  NOR2_X1 U3424 ( .A1(n4687), .A2(n4659), .ZN(n4686) );
  NOR2_X1 U3425 ( .A1(n4647), .A2(n4671), .ZN(n4687) );
  NAND2_X1 U3426 ( .A1(KEYINPUT4), .A2(n4688), .ZN(n4680) );
  INV_X1 U3427 ( .A(n4689), .ZN(n4688) );
  NAND2_X1 U3428 ( .A1(n4689), .A2(KEYINPUT32), .ZN(n4676) );
  NOR2_X1 U3429 ( .A1(n4651), .A2(n4690), .ZN(n4689) );
  NOR3_X1 U3430 ( .A1(n4647), .A2(n4641), .A3(n4671), .ZN(n4690) );
  INV_X1 U3431 ( .A(n4683), .ZN(n4671) );
  NAND2_X1 U3432 ( .A1(n4691), .A2(n4692), .ZN(n4651) );
  NAND2_X1 U3433 ( .A1(n4645), .A2(n4659), .ZN(n4692) );
  NAND2_X1 U3434 ( .A1(n4693), .A2(n4694), .ZN(n4659) );
  XNOR2_X1 U3435 ( .A(n4695), .B(n4673), .ZN(n4658) );
  INV_X1 U3436 ( .A(n4645), .ZN(n4641) );
  XNOR2_X1 U3437 ( .A(n4696), .B(n4697), .ZN(n4665) );
  NAND2_X1 U3438 ( .A1(KEYINPUT114), .A2(n4663), .ZN(n4697) );
  NAND2_X1 U3439 ( .A1(n4698), .A2(n4255), .ZN(n4572) );
  INV_X1 U3440 ( .A(n4196), .ZN(n4698) );
  XNOR2_X1 U3441 ( .A(n4699), .B(n4700), .ZN(n4196) );
  NOR2_X1 U3442 ( .A1(n4701), .A2(n4702), .ZN(n4700) );
  NOR2_X1 U3443 ( .A1(n4703), .A2(n4704), .ZN(n4702) );
  NOR2_X1 U3444 ( .A1(n4705), .A2(n4706), .ZN(n4704) );
  NOR2_X1 U3445 ( .A1(n4707), .A2(n4708), .ZN(n4706) );
  NOR2_X1 U3446 ( .A1(G257), .A2(n4709), .ZN(n4705) );
  NOR2_X1 U3447 ( .A1(G389), .A2(n4710), .ZN(n4701) );
  NOR2_X1 U3448 ( .A1(n4711), .A2(n4712), .ZN(n4710) );
  NOR2_X1 U3449 ( .A1(n4713), .A2(n4708), .ZN(n4712) );
  NOR2_X1 U3450 ( .A1(G257), .A2(G254), .ZN(n4711) );
  XOR2_X1 U3451 ( .A(n4714), .B(n4715), .Z(n4699) );
  XOR2_X1 U3452 ( .A(n4716), .B(n4717), .Z(n4715) );
  XOR2_X1 U3453 ( .A(n4718), .B(n4719), .Z(n4717) );
  NOR2_X1 U3454 ( .A1(n4720), .A2(n4721), .ZN(n4719) );
  NOR2_X1 U3455 ( .A1(n4722), .A2(n4723), .ZN(n4721) );
  NOR2_X1 U3456 ( .A1(n4724), .A2(n4725), .ZN(n4723) );
  NOR2_X1 U3457 ( .A1(n4726), .A2(n4727), .ZN(n4725) );
  INV_X1 U3458 ( .A(KEYINPUT40), .ZN(n4727) );
  NOR2_X1 U3459 ( .A1(n4728), .A2(n4729), .ZN(n4726) );
  NOR2_X1 U3460 ( .A1(n4707), .A2(n4730), .ZN(n4729) );
  NOR2_X1 U3461 ( .A1(G265), .A2(n4709), .ZN(n4728) );
  NOR2_X1 U3462 ( .A1(KEYINPUT40), .A2(n4731), .ZN(n4724) );
  NOR2_X1 U3463 ( .A1(n4732), .A2(n4733), .ZN(n4731) );
  NOR2_X1 U3464 ( .A1(n4709), .A2(n4730), .ZN(n4733) );
  NOR2_X1 U3465 ( .A1(G265), .A2(n4707), .ZN(n4732) );
  NOR2_X1 U3466 ( .A1(G400), .A2(n4734), .ZN(n4720) );
  NOR2_X1 U3467 ( .A1(n4735), .A2(n4736), .ZN(n4734) );
  NOR2_X1 U3468 ( .A1(n4730), .A2(n4713), .ZN(n4736) );
  NOR2_X1 U3469 ( .A1(G265), .A2(G254), .ZN(n4735) );
  NAND2_X1 U3470 ( .A1(n4737), .A2(n4738), .ZN(n4718) );
  NAND2_X1 U3471 ( .A1(n4739), .A2(n4740), .ZN(n4738) );
  NAND2_X1 U3472 ( .A1(n4741), .A2(n4742), .ZN(n4739) );
  NAND2_X1 U3473 ( .A1(n4743), .A2(n4744), .ZN(n4742) );
  INV_X1 U3474 ( .A(KEYINPUT11), .ZN(n4744) );
  NAND2_X1 U3475 ( .A1(n4745), .A2(n4746), .ZN(n4743) );
  NAND2_X1 U3476 ( .A1(n4747), .A2(n4748), .ZN(n4746) );
  NAND2_X1 U3477 ( .A1(G226), .A2(n4749), .ZN(n4745) );
  NAND2_X1 U3478 ( .A1(KEYINPUT11), .A2(n4750), .ZN(n4741) );
  NAND2_X1 U3479 ( .A1(n4751), .A2(n4752), .ZN(n4750) );
  NAND2_X1 U3480 ( .A1(G226), .A2(n4748), .ZN(n4752) );
  NAND2_X1 U3481 ( .A1(n4749), .A2(n4747), .ZN(n4751) );
  NAND2_X1 U3482 ( .A1(n4753), .A2(G422), .ZN(n4737) );
  NAND2_X1 U3483 ( .A1(n4754), .A2(n4755), .ZN(n4753) );
  NAND2_X1 U3484 ( .A1(G251), .A2(n4747), .ZN(n4755) );
  NAND2_X1 U3485 ( .A1(G226), .A2(G248), .ZN(n4754) );
  XOR2_X1 U3486 ( .A(n4756), .B(n4757), .Z(n4716) );
  NOR2_X1 U3487 ( .A1(n4758), .A2(n4759), .ZN(n4757) );
  NOR2_X1 U3488 ( .A1(n4760), .A2(n4761), .ZN(n4759) );
  NOR2_X1 U3489 ( .A1(n4762), .A2(n4763), .ZN(n4761) );
  NOR2_X1 U3490 ( .A1(n4707), .A2(n4764), .ZN(n4763) );
  NOR2_X1 U3491 ( .A1(G273), .A2(n4709), .ZN(n4762) );
  NOR2_X1 U3492 ( .A1(G411), .A2(n4765), .ZN(n4758) );
  NOR2_X1 U3493 ( .A1(n4766), .A2(n4767), .ZN(n4765) );
  NOR3_X1 U3494 ( .A1(n4764), .A2(n4768), .A3(n4713), .ZN(n4767) );
  AND2_X1 U3495 ( .A1(G254), .A2(KEYINPUT98), .ZN(n4768) );
  NOR2_X1 U3496 ( .A1(G273), .A2(n4769), .ZN(n4766) );
  NOR2_X1 U3497 ( .A1(KEYINPUT98), .A2(n4748), .ZN(n4769) );
  NAND2_X1 U3498 ( .A1(n4770), .A2(n4771), .ZN(n4756) );
  NAND2_X1 U3499 ( .A1(n4772), .A2(n4773), .ZN(n4771) );
  NAND2_X1 U3500 ( .A1(n4774), .A2(n4775), .ZN(n4772) );
  NAND2_X1 U3501 ( .A1(n4776), .A2(n4777), .ZN(n4775) );
  INV_X1 U3502 ( .A(KEYINPUT118), .ZN(n4777) );
  NAND2_X1 U3503 ( .A1(n4778), .A2(n4779), .ZN(n4776) );
  NAND2_X1 U3504 ( .A1(n4780), .A2(n4748), .ZN(n4779) );
  NAND2_X1 U3505 ( .A1(G218), .A2(n4749), .ZN(n4778) );
  NAND2_X1 U3506 ( .A1(KEYINPUT118), .A2(n4781), .ZN(n4774) );
  NAND2_X1 U3507 ( .A1(n4782), .A2(n4783), .ZN(n4781) );
  NAND2_X1 U3508 ( .A1(G218), .A2(n4748), .ZN(n4783) );
  NAND2_X1 U3509 ( .A1(n4749), .A2(n4780), .ZN(n4782) );
  NAND2_X1 U3510 ( .A1(n4784), .A2(G468), .ZN(n4770) );
  NAND2_X1 U3511 ( .A1(n4785), .A2(n4786), .ZN(n4784) );
  NAND2_X1 U3512 ( .A1(G251), .A2(n4780), .ZN(n4786) );
  NAND2_X1 U3513 ( .A1(G218), .A2(G248), .ZN(n4785) );
  XOR2_X1 U3514 ( .A(n4787), .B(n4788), .Z(n4714) );
  XOR2_X1 U3515 ( .A(n4789), .B(n4790), .Z(n4788) );
  NAND2_X1 U3516 ( .A1(n4791), .A2(n4792), .ZN(n4790) );
  NAND2_X1 U3517 ( .A1(G435), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U3518 ( .A1(n4794), .A2(n4795), .ZN(n4793) );
  NAND2_X1 U3519 ( .A1(G251), .A2(n4796), .ZN(n4795) );
  XNOR2_X1 U3520 ( .A(KEYINPUT68), .B(n4797), .ZN(n4796) );
  NAND2_X1 U3521 ( .A1(G234), .A2(G248), .ZN(n4794) );
  NAND2_X1 U3522 ( .A1(n4798), .A2(n4799), .ZN(n4791) );
  NAND2_X1 U3523 ( .A1(n4800), .A2(n4801), .ZN(n4798) );
  NAND2_X1 U3524 ( .A1(n4802), .A2(n4803), .ZN(n4801) );
  INV_X1 U3525 ( .A(KEYINPUT28), .ZN(n4803) );
  NAND2_X1 U3526 ( .A1(n4804), .A2(n4805), .ZN(n4802) );
  NAND2_X1 U3527 ( .A1(G234), .A2(n4748), .ZN(n4805) );
  NAND2_X1 U3528 ( .A1(n4749), .A2(n4797), .ZN(n4804) );
  NAND2_X1 U3529 ( .A1(KEYINPUT28), .A2(n4806), .ZN(n4800) );
  NAND2_X1 U3530 ( .A1(n4807), .A2(n4808), .ZN(n4806) );
  NAND2_X1 U3531 ( .A1(n4797), .A2(n4748), .ZN(n4808) );
  NAND2_X1 U3532 ( .A1(n4749), .A2(G234), .ZN(n4807) );
  NAND2_X1 U3533 ( .A1(n4809), .A2(n4810), .ZN(n4789) );
  NAND3_X1 U3534 ( .A1(n4811), .A2(n4812), .A3(n4813), .ZN(n4810) );
  NAND2_X1 U3535 ( .A1(n4814), .A2(n4815), .ZN(n4812) );
  INV_X1 U3536 ( .A(KEYINPUT21), .ZN(n4815) );
  NAND2_X1 U3537 ( .A1(n4816), .A2(n4817), .ZN(n4814) );
  NAND2_X1 U3538 ( .A1(G254), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U3539 ( .A1(G281), .A2(n4713), .ZN(n4816) );
  NAND2_X1 U3540 ( .A1(KEYINPUT21), .A2(n4819), .ZN(n4811) );
  NAND2_X1 U3541 ( .A1(n4820), .A2(n4821), .ZN(n4819) );
  NAND2_X1 U3542 ( .A1(n4713), .A2(n4818), .ZN(n4821) );
  NAND2_X1 U3543 ( .A1(G281), .A2(G254), .ZN(n4820) );
  XOR2_X1 U3544 ( .A(KEYINPUT101), .B(n4822), .Z(n4809) );
  NOR3_X1 U3545 ( .A1(n4813), .A2(n4823), .A3(n4824), .ZN(n4822) );
  NOR3_X1 U3546 ( .A1(n4818), .A2(G248), .A3(n4825), .ZN(n4824) );
  AND2_X1 U3547 ( .A1(G251), .A2(KEYINPUT123), .ZN(n4825) );
  NOR2_X1 U3548 ( .A1(G281), .A2(n4826), .ZN(n4823) );
  NOR2_X1 U3549 ( .A1(KEYINPUT123), .A2(n4709), .ZN(n4826) );
  XOR2_X1 U3550 ( .A(n4827), .B(n4828), .Z(n4787) );
  NOR3_X1 U3551 ( .A1(n4829), .A2(KEYINPUT105), .A3(n4830), .ZN(n4828) );
  NOR3_X1 U3552 ( .A1(n4831), .A2(n4832), .A3(n4833), .ZN(n4830) );
  NOR2_X1 U3553 ( .A1(G210), .A2(n4834), .ZN(n4833) );
  XNOR2_X1 U3554 ( .A(KEYINPUT0), .B(n4748), .ZN(n4834) );
  NOR2_X1 U3555 ( .A1(n4749), .A2(n4835), .ZN(n4832) );
  XNOR2_X1 U3556 ( .A(KEYINPUT61), .B(n4836), .ZN(n4831) );
  NOR3_X1 U3557 ( .A1(n4836), .A2(n4837), .A3(n4838), .ZN(n4829) );
  NOR2_X1 U3558 ( .A1(G251), .A2(G210), .ZN(n4838) );
  NOR2_X1 U3559 ( .A1(G248), .A2(n4835), .ZN(n4837) );
  OR3_X1 U3560 ( .A1(G1689), .A2(G176), .A3(n4839), .ZN(n4566) );
  NAND2_X1 U3561 ( .A1(n4524), .A2(n4446), .ZN(n4565) );
  INV_X1 U3562 ( .A(n4282), .ZN(n4446) );
  NAND3_X1 U3563 ( .A1(n4840), .A2(n4841), .A3(n4842), .ZN(n4282) );
  NAND2_X1 U3564 ( .A1(G94), .A2(G4092), .ZN(n4842) );
  NAND2_X1 U3565 ( .A1(n4255), .A2(n4843), .ZN(n4841) );
  XOR2_X1 U3566 ( .A(n4256), .B(n4257), .Z(n4843) );
  NAND3_X1 U3567 ( .A1(n4844), .A2(n4845), .A3(KEYINPUT15), .ZN(n4257) );
  NAND2_X1 U3568 ( .A1(n4846), .A2(n4847), .ZN(n4845) );
  XOR2_X1 U3569 ( .A(KEYINPUT25), .B(n4848), .Z(n4844) );
  NOR2_X1 U3570 ( .A1(n4847), .A2(n4846), .ZN(n4848) );
  XNOR2_X1 U3571 ( .A(n4849), .B(n4850), .ZN(n4846) );
  NAND2_X1 U3572 ( .A1(n4851), .A2(n4852), .ZN(n4849) );
  NAND2_X1 U3573 ( .A1(G254), .A2(n4853), .ZN(n4852) );
  XOR2_X1 U3574 ( .A(KEYINPUT122), .B(n4854), .Z(n4851) );
  NOR2_X1 U3575 ( .A1(n4855), .A2(n4853), .ZN(n4854) );
  XOR2_X1 U3576 ( .A(KEYINPUT22), .B(G293), .Z(n4853) );
  XNOR2_X1 U3577 ( .A(n4856), .B(n4857), .ZN(n4847) );
  NOR3_X1 U3578 ( .A1(n4858), .A2(n4859), .A3(n4860), .ZN(n4857) );
  NOR3_X1 U3579 ( .A1(n4861), .A2(n4862), .A3(n4709), .ZN(n4860) );
  XNOR2_X1 U3580 ( .A(G308), .B(KEYINPUT18), .ZN(n4862) );
  NOR2_X1 U3581 ( .A1(G479), .A2(n4863), .ZN(n4859) );
  NOR2_X1 U3582 ( .A1(n4864), .A2(n4865), .ZN(n4863) );
  NOR2_X1 U3583 ( .A1(G242), .A2(n4866), .ZN(n4865) );
  NOR2_X1 U3584 ( .A1(G308), .A2(G254), .ZN(n4864) );
  XOR2_X1 U3585 ( .A(n4867), .B(KEYINPUT80), .Z(n4858) );
  NAND2_X1 U3586 ( .A1(n4868), .A2(n4869), .ZN(n4856) );
  NAND3_X1 U3587 ( .A1(n4870), .A2(n4871), .A3(n4872), .ZN(n4869) );
  NAND2_X1 U3588 ( .A1(G254), .A2(n4873), .ZN(n4871) );
  NAND2_X1 U3589 ( .A1(G316), .A2(G242), .ZN(n4870) );
  NAND4_X1 U3590 ( .A1(n4874), .A2(n4875), .A3(n4876), .A4(n4877), .ZN(n4256) );
  NAND3_X1 U3591 ( .A1(n4563), .A2(n4878), .A3(n4879), .ZN(n4877) );
  NAND3_X1 U3592 ( .A1(n4880), .A2(n4878), .A3(n4881), .ZN(n4876) );
  INV_X1 U3593 ( .A(n4882), .ZN(n4878) );
  XNOR2_X1 U3594 ( .A(KEYINPUT71), .B(n4883), .ZN(n4880) );
  NAND3_X1 U3595 ( .A1(n4882), .A2(n4884), .A3(n4563), .ZN(n4875) );
  XNOR2_X1 U3596 ( .A(n4879), .B(KEYINPUT72), .ZN(n4884) );
  NAND3_X1 U3597 ( .A1(n4882), .A2(n4879), .A3(n4883), .ZN(n4874) );
  INV_X1 U3598 ( .A(n4881), .ZN(n4879) );
  NAND2_X1 U3599 ( .A1(n4885), .A2(n4886), .ZN(n4881) );
  NAND2_X1 U3600 ( .A1(n4887), .A2(n4888), .ZN(n4886) );
  XNOR2_X1 U3601 ( .A(n4889), .B(n4855), .ZN(n4887) );
  NAND2_X1 U3602 ( .A1(n4890), .A2(G514), .ZN(n4885) );
  XNOR2_X1 U3603 ( .A(G248), .B(n4889), .ZN(n4890) );
  NAND2_X1 U3604 ( .A1(n4891), .A2(n4892), .ZN(n4889) );
  NAND2_X1 U3605 ( .A1(n4893), .A2(n4894), .ZN(n4892) );
  NAND2_X1 U3606 ( .A1(n4895), .A2(n4896), .ZN(n4893) );
  NAND2_X1 U3607 ( .A1(n4748), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U3608 ( .A1(G324), .A2(n4855), .ZN(n4895) );
  NAND2_X1 U3609 ( .A1(n4898), .A2(G503), .ZN(n4891) );
  NAND2_X1 U3610 ( .A1(n4899), .A2(n4900), .ZN(n4898) );
  NAND2_X1 U3611 ( .A1(G251), .A2(n4897), .ZN(n4900) );
  NAND2_X1 U3612 ( .A1(G324), .A2(G248), .ZN(n4899) );
  XNOR2_X1 U3613 ( .A(n4901), .B(n4902), .ZN(n4882) );
  NOR2_X1 U3614 ( .A1(n4903), .A2(n4904), .ZN(n4902) );
  NOR2_X1 U3615 ( .A1(n4905), .A2(n4906), .ZN(n4904) );
  NOR2_X1 U3616 ( .A1(n4907), .A2(n4908), .ZN(n4906) );
  NOR2_X1 U3617 ( .A1(n4909), .A2(n4707), .ZN(n4908) );
  NOR2_X1 U3618 ( .A1(G351), .A2(n4709), .ZN(n4907) );
  NOR2_X1 U3619 ( .A1(G534), .A2(n4910), .ZN(n4903) );
  NOR2_X1 U3620 ( .A1(n4911), .A2(n4912), .ZN(n4910) );
  NOR2_X1 U3621 ( .A1(G242), .A2(n4909), .ZN(n4912) );
  NOR2_X1 U3622 ( .A1(G351), .A2(G254), .ZN(n4911) );
  NAND2_X1 U3623 ( .A1(n4913), .A2(n4914), .ZN(n4901) );
  NAND3_X1 U3624 ( .A1(n4915), .A2(n4916), .A3(G523), .ZN(n4914) );
  NAND2_X1 U3625 ( .A1(n4709), .A2(n4917), .ZN(n4916) );
  NAND2_X1 U3626 ( .A1(n4918), .A2(G341), .ZN(n4915) );
  XNOR2_X1 U3627 ( .A(G248), .B(KEYINPUT43), .ZN(n4918) );
  XOR2_X1 U3628 ( .A(n4919), .B(KEYINPUT8), .Z(n4913) );
  NAND3_X1 U3629 ( .A1(n4920), .A2(n4921), .A3(n4922), .ZN(n4919) );
  NAND2_X1 U3630 ( .A1(G254), .A2(n4917), .ZN(n4921) );
  NAND2_X1 U3631 ( .A1(G242), .A2(G341), .ZN(n4920) );
  NAND2_X1 U3632 ( .A1(n4506), .A2(n4923), .ZN(n4840) );
  XOR2_X1 U3633 ( .A(KEYINPUT100), .B(n4253), .Z(n4923) );
  XNOR2_X1 U3634 ( .A(n4924), .B(n4925), .ZN(n4253) );
  NOR2_X1 U3635 ( .A1(n4926), .A2(n4927), .ZN(n4925) );
  NOR2_X1 U3636 ( .A1(n4928), .A2(n4929), .ZN(n4927) );
  XOR2_X1 U3637 ( .A(n4930), .B(n4931), .Z(n4929) );
  XOR2_X1 U3638 ( .A(n4932), .B(n4933), .Z(n4931) );
  XNOR2_X1 U3639 ( .A(n4934), .B(n4235), .ZN(n4933) );
  NOR3_X1 U3640 ( .A1(n4935), .A2(n4936), .A3(n4937), .ZN(n4932) );
  XOR2_X1 U3641 ( .A(n4938), .B(n4939), .Z(n4930) );
  NOR3_X1 U3642 ( .A1(n4940), .A2(n4941), .A3(n4942), .ZN(n4939) );
  NOR2_X1 U3643 ( .A1(n4943), .A2(n4944), .ZN(n4942) );
  NOR3_X1 U3644 ( .A1(n4945), .A2(n4946), .A3(n4947), .ZN(n4941) );
  NOR2_X1 U3645 ( .A1(n4948), .A2(n4949), .ZN(n4940) );
  XNOR2_X1 U3646 ( .A(n4946), .B(n4945), .ZN(n4949) );
  NAND2_X1 U3647 ( .A1(n4950), .A2(n4951), .ZN(n4938) );
  NAND3_X1 U3648 ( .A1(n4952), .A2(n4953), .A3(n4954), .ZN(n4951) );
  NAND2_X1 U3649 ( .A1(n4955), .A2(n4956), .ZN(n4952) );
  NAND2_X1 U3650 ( .A1(n4957), .A2(n4944), .ZN(n4956) );
  NAND2_X1 U3651 ( .A1(n4948), .A2(n4958), .ZN(n4955) );
  NAND3_X1 U3652 ( .A1(n4959), .A2(n4947), .A3(n4960), .ZN(n4950) );
  INV_X1 U3653 ( .A(G2174), .ZN(n4928) );
  NOR2_X1 U3654 ( .A1(n4961), .A2(n4962), .ZN(n4926) );
  XOR2_X1 U3655 ( .A(n4963), .B(n4964), .Z(n4962) );
  NAND2_X1 U3656 ( .A1(KEYINPUT106), .A2(n4943), .ZN(n4964) );
  NAND3_X1 U3657 ( .A1(n4965), .A2(n4966), .A3(n4967), .ZN(n4963) );
  OR2_X1 U3658 ( .A1(n4968), .A2(n4969), .ZN(n4967) );
  NAND3_X1 U3659 ( .A1(n4969), .A2(n4968), .A3(KEYINPUT86), .ZN(n4966) );
  XNOR2_X1 U3660 ( .A(n4970), .B(n4971), .ZN(n4968) );
  XNOR2_X1 U3661 ( .A(n4957), .B(n4972), .ZN(n4971) );
  XOR2_X1 U3662 ( .A(n4973), .B(n4974), .Z(n4972) );
  NOR3_X1 U3663 ( .A1(n4935), .A2(n4975), .A3(n4976), .ZN(n4974) );
  AND3_X1 U3664 ( .A1(KEYINPUT19), .A2(n4945), .A3(n4960), .ZN(n4976) );
  NOR2_X1 U3665 ( .A1(KEYINPUT19), .A2(n4977), .ZN(n4975) );
  NAND2_X1 U3666 ( .A1(n4978), .A2(n4979), .ZN(n4935) );
  NAND2_X1 U3667 ( .A1(n4943), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U3668 ( .A1(n4953), .A2(n4981), .ZN(n4980) );
  INV_X1 U3669 ( .A(n4982), .ZN(n4981) );
  NOR3_X1 U3670 ( .A1(n4983), .A2(n4960), .A3(n4982), .ZN(n4973) );
  NOR2_X1 U3671 ( .A1(n4944), .A2(n4984), .ZN(n4982) );
  XNOR2_X1 U3672 ( .A(KEYINPUT7), .B(n4953), .ZN(n4983) );
  NAND3_X1 U3673 ( .A1(G534), .A2(n4233), .A3(n4946), .ZN(n4953) );
  XNOR2_X1 U3674 ( .A(n4985), .B(n4948), .ZN(n4970) );
  NAND2_X1 U3675 ( .A1(KEYINPUT115), .A2(n4934), .ZN(n4985) );
  AND2_X1 U3676 ( .A1(KEYINPUT94), .A2(n4946), .ZN(n4969) );
  OR2_X1 U3677 ( .A1(n4946), .A2(KEYINPUT86), .ZN(n4965) );
  NAND3_X1 U3678 ( .A1(n4986), .A2(n4987), .A3(n4988), .ZN(n4924) );
  NAND2_X1 U3679 ( .A1(KEYINPUT33), .A2(n4989), .ZN(n4988) );
  OR3_X1 U3680 ( .A1(n4990), .A2(n4991), .A3(n4961), .ZN(n4989) );
  NAND3_X1 U3681 ( .A1(n4992), .A2(n4993), .A3(n4994), .ZN(n4987) );
  INV_X1 U3682 ( .A(n4961), .ZN(n4994) );
  XOR2_X1 U3683 ( .A(G2174), .B(KEYINPUT24), .Z(n4961) );
  NAND2_X1 U3684 ( .A1(n4991), .A2(n4995), .ZN(n4993) );
  NAND2_X1 U3685 ( .A1(KEYINPUT121), .A2(n4996), .ZN(n4995) );
  NAND3_X1 U3686 ( .A1(n4997), .A2(n4998), .A3(n4999), .ZN(n4992) );
  NAND2_X1 U3687 ( .A1(n4996), .A2(n5000), .ZN(n4998) );
  INV_X1 U3688 ( .A(KEYINPUT121), .ZN(n5000) );
  OR2_X1 U3689 ( .A1(n4990), .A2(KEYINPUT33), .ZN(n4997) );
  NAND3_X1 U3690 ( .A1(n5001), .A2(n5002), .A3(G2174), .ZN(n4986) );
  NAND2_X1 U3691 ( .A1(n4990), .A2(n5003), .ZN(n5002) );
  XNOR2_X1 U3692 ( .A(n5004), .B(n5005), .ZN(n4990) );
  XNOR2_X1 U3693 ( .A(n5006), .B(n5007), .ZN(n5005) );
  XNOR2_X1 U3694 ( .A(n4246), .B(n5008), .ZN(n5007) );
  XOR2_X1 U3695 ( .A(n5009), .B(n5010), .Z(n5004) );
  XNOR2_X1 U3696 ( .A(n5011), .B(n5012), .ZN(n5010) );
  NOR2_X1 U3697 ( .A1(KEYINPUT89), .A2(n5013), .ZN(n5012) );
  NAND2_X1 U3698 ( .A1(KEYINPUT110), .A2(n5014), .ZN(n5011) );
  NAND2_X1 U3699 ( .A1(n5015), .A2(n5008), .ZN(n5014) );
  XNOR2_X1 U3700 ( .A(n5015), .B(n5016), .ZN(n5009) );
  NOR2_X1 U3701 ( .A1(n5017), .A2(KEYINPUT66), .ZN(n5016) );
  AND2_X1 U3702 ( .A1(n5018), .A2(n5019), .ZN(n5015) );
  NAND2_X1 U3703 ( .A1(n5006), .A2(n5013), .ZN(n5019) );
  NAND2_X1 U3704 ( .A1(n5020), .A2(n5021), .ZN(n5001) );
  INV_X1 U3705 ( .A(n5003), .ZN(n5021) );
  NAND2_X1 U3706 ( .A1(n4991), .A2(n5022), .ZN(n5003) );
  XNOR2_X1 U3707 ( .A(KEYINPUT12), .B(n5023), .ZN(n5022) );
  INV_X1 U3708 ( .A(n4999), .ZN(n4991) );
  XOR2_X1 U3709 ( .A(n4996), .B(KEYINPUT124), .Z(n5020) );
  XNOR2_X1 U3710 ( .A(n5024), .B(n4243), .ZN(n4996) );
  NAND2_X1 U3711 ( .A1(n5025), .A2(n5026), .ZN(n5024) );
  NAND2_X1 U3712 ( .A1(n5027), .A2(n4246), .ZN(n5026) );
  XOR2_X1 U3713 ( .A(KEYINPUT85), .B(n5028), .Z(n5025) );
  NOR2_X1 U3714 ( .A1(n4246), .A2(n5027), .ZN(n5028) );
  XOR2_X1 U3715 ( .A(n5029), .B(n5030), .Z(n5027) );
  XNOR2_X1 U3716 ( .A(n5013), .B(n5031), .ZN(n5030) );
  XOR2_X1 U3717 ( .A(n5032), .B(n5018), .Z(n5031) );
  XNOR2_X1 U3718 ( .A(n5033), .B(n5034), .ZN(n5029) );
  NAND2_X1 U3719 ( .A1(KEYINPUT29), .A2(n5006), .ZN(n5033) );
  NAND2_X1 U3720 ( .A1(G140), .A2(n4259), .ZN(G656) );
  NAND4_X1 U3721 ( .A1(n5035), .A2(n5036), .A3(n5037), .A4(n5038), .ZN(G654) );
  NAND2_X1 U3722 ( .A1(n4492), .A2(n4389), .ZN(n5038) );
  NAND3_X1 U3723 ( .A1(n5039), .A2(n5040), .A3(n5041), .ZN(n4389) );
  NAND2_X1 U3724 ( .A1(n4506), .A2(n5042), .ZN(n5041) );
  NAND3_X1 U3725 ( .A1(n5043), .A2(n5044), .A3(n4255), .ZN(n5040) );
  NAND3_X1 U3726 ( .A1(G446), .A2(G251), .A3(n5045), .ZN(n5044) );
  XNOR2_X1 U3727 ( .A(G206), .B(KEYINPUT79), .ZN(n5045) );
  NAND2_X1 U3728 ( .A1(G115), .A2(n4504), .ZN(n5039) );
  NAND2_X1 U3729 ( .A1(n4500), .A2(n4386), .ZN(n5037) );
  NAND3_X1 U3730 ( .A1(n5046), .A2(n5047), .A3(n5048), .ZN(n4386) );
  NAND2_X1 U3731 ( .A1(n4506), .A2(n5049), .ZN(n5048) );
  NAND2_X1 U3732 ( .A1(G123), .A2(n4504), .ZN(n5047) );
  NAND2_X1 U3733 ( .A1(n4255), .A2(n4269), .ZN(n5046) );
  NAND2_X1 U3734 ( .A1(n4508), .A2(G191), .ZN(n5036) );
  NAND2_X1 U3735 ( .A1(n4509), .A2(G161), .ZN(n5035) );
  NOR2_X1 U3736 ( .A1(n4449), .A2(n5050), .ZN(G651) );
  XOR2_X1 U3737 ( .A(KEYINPUT70), .B(n5051), .Z(n5050) );
  NOR4_X1 U3738 ( .A1(n5052), .A2(n5053), .A3(n5054), .A4(n5055), .ZN(n5051) );
  NOR3_X1 U3739 ( .A1(n4839), .A2(G1689), .A3(n4462), .ZN(n5055) );
  INV_X1 U3740 ( .A(G194), .ZN(n4462) );
  NOR2_X1 U3741 ( .A1(G826), .A2(n5056), .ZN(n5054) );
  INV_X1 U3742 ( .A(n4333), .ZN(G826) );
  NAND3_X1 U3743 ( .A1(n5057), .A2(n5058), .A3(n5059), .ZN(n4333) );
  NAND2_X1 U3744 ( .A1(n4255), .A2(n4850), .ZN(n5059) );
  NAND2_X1 U3745 ( .A1(n5060), .A2(n4506), .ZN(n5058) );
  NAND2_X1 U3746 ( .A1(G121), .A2(n4504), .ZN(n5057) );
  NOR2_X1 U3747 ( .A1(G865), .A2(n4571), .ZN(n5053) );
  INV_X1 U3748 ( .A(n4332), .ZN(G865) );
  NAND3_X1 U3749 ( .A1(n5061), .A2(n5062), .A3(n5063), .ZN(n4332) );
  NAND2_X1 U3750 ( .A1(n5064), .A2(n4255), .ZN(n5063) );
  INV_X1 U3751 ( .A(n5065), .ZN(n5064) );
  NAND3_X1 U3752 ( .A1(n5066), .A2(n5067), .A3(n4506), .ZN(n5062) );
  NAND2_X1 U3753 ( .A1(G114), .A2(n4504), .ZN(n5061) );
  NOR2_X1 U3754 ( .A1(n4463), .A2(n4570), .ZN(n5052) );
  INV_X1 U3755 ( .A(G164), .ZN(n4463) );
  NAND4_X1 U3756 ( .A1(n5068), .A2(n5069), .A3(n5070), .A4(n5071), .ZN(G648) );
  NAND2_X1 U3757 ( .A1(n5072), .A2(n4500), .ZN(n5071) );
  XNOR2_X1 U3758 ( .A(G828), .B(KEYINPUT81), .ZN(n5072) );
  INV_X1 U3759 ( .A(n4324), .ZN(G828) );
  NAND3_X1 U3760 ( .A1(n5073), .A2(n5074), .A3(n5075), .ZN(n4324) );
  NAND2_X1 U3761 ( .A1(n4506), .A2(n5076), .ZN(n5075) );
  NAND2_X1 U3762 ( .A1(G116), .A2(n4504), .ZN(n5074) );
  NAND2_X1 U3763 ( .A1(n5077), .A2(n4255), .ZN(n5073) );
  INV_X1 U3764 ( .A(n5078), .ZN(n5077) );
  NAND2_X1 U3765 ( .A1(n4492), .A2(n4325), .ZN(n5070) );
  NAND3_X1 U3766 ( .A1(n5079), .A2(n5080), .A3(n5081), .ZN(n4325) );
  NAND2_X1 U3767 ( .A1(n4506), .A2(n5082), .ZN(n5081) );
  NAND2_X1 U3768 ( .A1(G53), .A2(n4504), .ZN(n5080) );
  NAND2_X1 U3769 ( .A1(n5083), .A2(n4255), .ZN(n5079) );
  INV_X1 U3770 ( .A(n5084), .ZN(n5083) );
  NAND2_X1 U3771 ( .A1(n4508), .A2(G197), .ZN(n5069) );
  NAND2_X1 U3772 ( .A1(n4509), .A2(G167), .ZN(n5068) );
  NAND4_X1 U3773 ( .A1(n5085), .A2(n5086), .A3(n5087), .A4(n5088), .ZN(G645) );
  NAND2_X1 U3774 ( .A1(n4492), .A2(n4319), .ZN(n5088) );
  NAND3_X1 U3775 ( .A1(n5089), .A2(n5090), .A3(n5091), .ZN(n4319) );
  NAND2_X1 U3776 ( .A1(n5092), .A2(n4506), .ZN(n5091) );
  NAND2_X1 U3777 ( .A1(G113), .A2(n4504), .ZN(n5090) );
  NAND2_X1 U3778 ( .A1(n5093), .A2(n4255), .ZN(n5089) );
  INV_X1 U3779 ( .A(n5094), .ZN(n5093) );
  NAND2_X1 U3780 ( .A1(n4500), .A2(n4318), .ZN(n5087) );
  NAND3_X1 U3781 ( .A1(n5095), .A2(n5096), .A3(n5097), .ZN(n4318) );
  NAND2_X1 U3782 ( .A1(n5098), .A2(n4255), .ZN(n5097) );
  INV_X1 U3783 ( .A(n5099), .ZN(n5098) );
  NAND2_X1 U3784 ( .A1(n5100), .A2(n4506), .ZN(n5096) );
  NAND2_X1 U3785 ( .A1(G112), .A2(n4504), .ZN(n5095) );
  NAND2_X1 U3786 ( .A1(n4508), .A2(G203), .ZN(n5086) );
  NAND2_X1 U3787 ( .A1(n4509), .A2(G173), .ZN(n5085) );
  NAND4_X1 U3788 ( .A1(n5101), .A2(n5102), .A3(n5103), .A4(n5104), .ZN(G642) );
  NAND2_X1 U3789 ( .A1(n4508), .A2(G200), .ZN(n5104) );
  NOR3_X1 U3790 ( .A1(n4449), .A2(G1689), .A3(n4839), .ZN(n4508) );
  NAND2_X1 U3791 ( .A1(n4509), .A2(G170), .ZN(n5103) );
  NOR2_X1 U3792 ( .A1(n4570), .A2(n4449), .ZN(n4509) );
  NAND2_X1 U3793 ( .A1(G1690), .A2(G1689), .ZN(n4570) );
  NAND2_X1 U3794 ( .A1(n4492), .A2(n4312), .ZN(n5102) );
  NAND3_X1 U3795 ( .A1(n5105), .A2(n5106), .A3(n5107), .ZN(n4312) );
  NAND2_X1 U3796 ( .A1(n4506), .A2(n5108), .ZN(n5107) );
  NAND2_X1 U3797 ( .A1(G122), .A2(n4504), .ZN(n5106) );
  NAND2_X1 U3798 ( .A1(n4255), .A2(n5109), .ZN(n5105) );
  NOR2_X1 U3799 ( .A1(n4571), .A2(n4449), .ZN(n4492) );
  NAND2_X1 U3800 ( .A1(G1689), .A2(n4839), .ZN(n4571) );
  INV_X1 U3801 ( .A(G1690), .ZN(n4839) );
  NAND2_X1 U3802 ( .A1(n4500), .A2(n4310), .ZN(n5101) );
  NAND3_X1 U3803 ( .A1(n5110), .A2(n5111), .A3(n5112), .ZN(n4310) );
  NAND2_X1 U3804 ( .A1(n4506), .A2(n5113), .ZN(n5112) );
  AND2_X1 U3805 ( .A1(G4091), .A2(n4202), .ZN(n4506) );
  NAND3_X1 U3806 ( .A1(n5114), .A2(n5115), .A3(n4255), .ZN(n5111) );
  NAND2_X1 U3807 ( .A1(G52), .A2(n4504), .ZN(n5110) );
  INV_X1 U3808 ( .A(G4092), .ZN(n4202) );
  NOR2_X1 U3809 ( .A1(n5056), .A2(n4449), .ZN(n4500) );
  INV_X1 U3810 ( .A(G137), .ZN(n4449) );
  INV_X1 U3811 ( .A(n4524), .ZN(n5056) );
  NOR2_X1 U3812 ( .A1(G1689), .A2(G1690), .ZN(n4524) );
  AND2_X1 U3813 ( .A1(G141), .A2(n5116), .ZN(G639) );
  NAND3_X1 U3814 ( .A1(n5117), .A2(n5118), .A3(n4259), .ZN(n5116) );
  INV_X1 U3815 ( .A(G809), .ZN(n4259) );
  NAND2_X1 U3816 ( .A1(G24), .A2(n4396), .ZN(n5118) );
  NAND2_X1 U3817 ( .A1(G25), .A2(G2358), .ZN(n5117) );
  OR3_X1 U3818 ( .A1(n5119), .A2(n5120), .A3(G809), .ZN(G636) );
  NAND2_X1 U3819 ( .A1(G31), .A2(G27), .ZN(G809) );
  NOR2_X1 U3820 ( .A1(G86), .A2(G2358), .ZN(n5120) );
  NOR2_X1 U3821 ( .A1(G87), .A2(n4396), .ZN(n5119) );
  INV_X1 U3822 ( .A(G2358), .ZN(n4396) );
  AND2_X1 U3823 ( .A1(G1), .A2(G373), .ZN(G634) );
  NOR4_X1 U3824 ( .A1(n5121), .A2(n5122), .A3(n5123), .A4(n5124), .ZN(G632) );
  NAND3_X1 U3825 ( .A1(n5125), .A2(n4683), .A3(n5126), .ZN(n5121) );
  NAND3_X1 U3826 ( .A1(n5034), .A2(n5127), .A3(n4246), .ZN(G629) );
  NAND3_X1 U3827 ( .A1(n5013), .A2(n4999), .A3(n5006), .ZN(n5127) );
  NAND2_X1 U3828 ( .A1(n5128), .A2(n5129), .ZN(n4999) );
  NAND2_X1 U3829 ( .A1(n4934), .A2(n5130), .ZN(n5129) );
  NAND4_X1 U3830 ( .A1(n4978), .A2(n5131), .A3(n5132), .A4(n5133), .ZN(n5130) );
  OR3_X1 U3831 ( .A1(n4954), .A2(n4943), .A3(KEYINPUT112), .ZN(n5133) );
  NAND2_X1 U3832 ( .A1(KEYINPUT112), .A2(n4937), .ZN(n5132) );
  NAND2_X1 U3833 ( .A1(n5134), .A2(G514), .ZN(n4978) );
  XNOR2_X1 U3834 ( .A(n5135), .B(KEYINPUT107), .ZN(n5134) );
  INV_X1 U3835 ( .A(n4231), .ZN(n5135) );
  AND2_X1 U3836 ( .A1(n5018), .A2(n5008), .ZN(n5034) );
  AND3_X1 U3837 ( .A1(n5136), .A2(n5137), .A3(n5138), .ZN(n5018) );
  NAND2_X1 U3838 ( .A1(n5032), .A2(n5006), .ZN(n5138) );
  OR2_X1 U3839 ( .A1(n5139), .A2(KEYINPUT30), .ZN(n5137) );
  NAND3_X1 U3840 ( .A1(n5140), .A2(n4861), .A3(KEYINPUT30), .ZN(n5136) );
  NOR3_X1 U3841 ( .A1(n5141), .A2(n5023), .A3(n5142), .ZN(G626) );
  NAND4_X1 U3842 ( .A1(n5143), .A2(n4934), .A3(n5144), .A4(n4943), .ZN(n5023) );
  NOR2_X1 U3843 ( .A1(n4235), .A2(n4947), .ZN(n5144) );
  AND3_X1 U3844 ( .A1(n5145), .A2(n5146), .A3(n5128), .ZN(n4934) );
  OR3_X1 U3845 ( .A1(n4230), .A2(G503), .A3(KEYINPUT93), .ZN(n5146) );
  NAND2_X1 U3846 ( .A1(KEYINPUT93), .A2(n4230), .ZN(n5145) );
  XNOR2_X1 U3847 ( .A(n4946), .B(KEYINPUT35), .ZN(n5143) );
  NAND3_X1 U3848 ( .A1(n5008), .A2(n5013), .A3(n5006), .ZN(n5141) );
  AND2_X1 U3849 ( .A1(n5147), .A2(n5148), .ZN(n5006) );
  NAND2_X1 U3850 ( .A1(KEYINPUT87), .A2(n5149), .ZN(n5148) );
  NAND2_X1 U3851 ( .A1(n5150), .A2(n5151), .ZN(n5147) );
  INV_X1 U3852 ( .A(KEYINPUT87), .ZN(n5151) );
  XNOR2_X1 U3853 ( .A(G479), .B(n4244), .ZN(n5150) );
  NAND2_X1 U3854 ( .A1(n5152), .A2(n5153), .ZN(n5013) );
  NAND2_X1 U3855 ( .A1(KEYINPUT34), .A2(n5154), .ZN(n5153) );
  NAND2_X1 U3856 ( .A1(n5155), .A2(n5156), .ZN(n5152) );
  INV_X1 U3857 ( .A(KEYINPUT34), .ZN(n5156) );
  NAND2_X1 U3858 ( .A1(n5157), .A2(n5158), .ZN(G621) );
  NAND2_X1 U3859 ( .A1(n5159), .A2(n5160), .ZN(n5158) );
  NAND2_X1 U3860 ( .A1(n5161), .A2(n5162), .ZN(n5160) );
  NAND2_X1 U3861 ( .A1(n5126), .A2(n5163), .ZN(n5162) );
  INV_X1 U3862 ( .A(n5164), .ZN(n5161) );
  NAND3_X1 U3863 ( .A1(n4246), .A2(n5165), .A3(n5166), .ZN(G618) );
  XNOR2_X1 U3864 ( .A(KEYINPUT2), .B(n4243), .ZN(n5166) );
  NAND2_X1 U3865 ( .A1(n5167), .A2(n5168), .ZN(n5165) );
  NAND3_X1 U3866 ( .A1(n5169), .A2(n5170), .A3(n5171), .ZN(n5168) );
  XOR2_X1 U3867 ( .A(n5139), .B(KEYINPUT125), .Z(n5171) );
  NAND2_X1 U3868 ( .A1(n5172), .A2(n5173), .ZN(n5170) );
  INV_X1 U3869 ( .A(n5174), .ZN(n5172) );
  NOR3_X1 U3870 ( .A1(n5175), .A2(n5176), .A3(n5174), .ZN(G615) );
  INV_X1 U3871 ( .A(n4936), .ZN(n5176) );
  NAND3_X1 U3872 ( .A1(n5167), .A2(n5177), .A3(n4246), .ZN(n5175) );
  INV_X1 U3873 ( .A(n5142), .ZN(n4246) );
  INV_X1 U3874 ( .A(G358), .ZN(G612) );
  INV_X1 U3875 ( .A(G338), .ZN(G611) );
  NOR4_X1 U3876 ( .A1(n5178), .A2(n5179), .A3(n4496), .A4(n5109), .ZN(G610) );
  AND2_X1 U3877 ( .A1(n5180), .A2(n5181), .ZN(n5109) );
  NAND2_X1 U3878 ( .A1(n5182), .A2(n4799), .ZN(n5181) );
  NAND2_X1 U3879 ( .A1(n5183), .A2(n5184), .ZN(n5182) );
  NAND2_X1 U3880 ( .A1(G3546), .A2(G234), .ZN(n5184) );
  NAND2_X1 U3881 ( .A1(n5185), .A2(n4797), .ZN(n5183) );
  NAND2_X1 U3882 ( .A1(n5186), .A2(G435), .ZN(n5180) );
  NAND2_X1 U3883 ( .A1(n5187), .A2(n5188), .ZN(n5186) );
  NAND2_X1 U3884 ( .A1(n4797), .A2(n5189), .ZN(n5188) );
  INV_X1 U3885 ( .A(G234), .ZN(n4797) );
  NAND2_X1 U3886 ( .A1(G234), .A2(n5190), .ZN(n5187) );
  AND2_X1 U3887 ( .A1(n5191), .A2(n5192), .ZN(n4496) );
  NAND2_X1 U3888 ( .A1(n5193), .A2(n4703), .ZN(n5192) );
  NAND2_X1 U3889 ( .A1(n5194), .A2(n5195), .ZN(n5193) );
  NAND2_X1 U3890 ( .A1(G257), .A2(G3546), .ZN(n5195) );
  NAND2_X1 U3891 ( .A1(n5185), .A2(n4708), .ZN(n5194) );
  NAND2_X1 U3892 ( .A1(n5196), .A2(G389), .ZN(n5191) );
  NAND2_X1 U3893 ( .A1(n5197), .A2(n5198), .ZN(n5196) );
  NAND2_X1 U3894 ( .A1(n4708), .A2(n5189), .ZN(n5198) );
  NAND2_X1 U3895 ( .A1(G257), .A2(n5190), .ZN(n5197) );
  NAND3_X1 U3896 ( .A1(n4541), .A2(n4827), .A3(n4520), .ZN(n5179) );
  NAND2_X1 U3897 ( .A1(n5199), .A2(n5200), .ZN(n4520) );
  NAND2_X1 U3898 ( .A1(n5201), .A2(n4722), .ZN(n5200) );
  NAND2_X1 U3899 ( .A1(n5202), .A2(n5203), .ZN(n5201) );
  NAND2_X1 U3900 ( .A1(G3546), .A2(G265), .ZN(n5203) );
  NAND2_X1 U3901 ( .A1(n5185), .A2(n4730), .ZN(n5202) );
  NAND2_X1 U3902 ( .A1(n5204), .A2(G400), .ZN(n5199) );
  NAND2_X1 U3903 ( .A1(n5205), .A2(n5206), .ZN(n5204) );
  NAND2_X1 U3904 ( .A1(n4730), .A2(n5189), .ZN(n5206) );
  NAND2_X1 U3905 ( .A1(G265), .A2(n5190), .ZN(n5205) );
  NAND2_X1 U3906 ( .A1(n5043), .A2(n5207), .ZN(n4827) );
  NAND3_X1 U3907 ( .A1(G251), .A2(n5208), .A3(G446), .ZN(n5207) );
  AND2_X1 U3908 ( .A1(n5209), .A2(n5210), .ZN(n5043) );
  NAND2_X1 U3909 ( .A1(n5211), .A2(n5212), .ZN(n5210) );
  INV_X1 U3910 ( .A(G446), .ZN(n5212) );
  NAND2_X1 U3911 ( .A1(n5213), .A2(n5214), .ZN(n5211) );
  NAND2_X1 U3912 ( .A1(G206), .A2(n4855), .ZN(n5214) );
  INV_X1 U3913 ( .A(G242), .ZN(n4855) );
  NAND2_X1 U3914 ( .A1(n5208), .A2(n4748), .ZN(n5213) );
  INV_X1 U3915 ( .A(G206), .ZN(n5208) );
  NAND3_X1 U3916 ( .A1(G206), .A2(G248), .A3(G446), .ZN(n5209) );
  NAND2_X1 U3917 ( .A1(n5215), .A2(n5216), .ZN(n4541) );
  NAND2_X1 U3918 ( .A1(n5217), .A2(n4760), .ZN(n5216) );
  INV_X1 U3919 ( .A(G411), .ZN(n4760) );
  NAND2_X1 U3920 ( .A1(n5218), .A2(n5219), .ZN(n5217) );
  NAND2_X1 U3921 ( .A1(G3546), .A2(G273), .ZN(n5219) );
  NAND2_X1 U3922 ( .A1(n5185), .A2(n4764), .ZN(n5218) );
  NAND2_X1 U3923 ( .A1(n5220), .A2(G411), .ZN(n5215) );
  NAND2_X1 U3924 ( .A1(n5221), .A2(n5222), .ZN(n5220) );
  NAND2_X1 U3925 ( .A1(n4764), .A2(n5189), .ZN(n5222) );
  INV_X1 U3926 ( .A(G273), .ZN(n4764) );
  NAND2_X1 U3927 ( .A1(G273), .A2(n5190), .ZN(n5221) );
  NAND4_X1 U3928 ( .A1(n4558), .A2(n5065), .A3(n5084), .A4(n5094), .ZN(n5178) );
  NAND2_X1 U3929 ( .A1(n5223), .A2(n5224), .ZN(n5094) );
  NAND2_X1 U3930 ( .A1(n5225), .A2(n4740), .ZN(n5224) );
  INV_X1 U3931 ( .A(G422), .ZN(n4740) );
  NAND2_X1 U3932 ( .A1(n5226), .A2(n5227), .ZN(n5225) );
  NAND2_X1 U3933 ( .A1(G226), .A2(G3546), .ZN(n5227) );
  NAND2_X1 U3934 ( .A1(n5185), .A2(n4747), .ZN(n5226) );
  NAND2_X1 U3935 ( .A1(n5228), .A2(G422), .ZN(n5223) );
  NAND2_X1 U3936 ( .A1(n5229), .A2(n5230), .ZN(n5228) );
  NAND2_X1 U3937 ( .A1(n4747), .A2(n5189), .ZN(n5230) );
  NAND2_X1 U3938 ( .A1(G226), .A2(n5190), .ZN(n5229) );
  NAND2_X1 U3939 ( .A1(n5231), .A2(n5232), .ZN(n5084) );
  NAND2_X1 U3940 ( .A1(n5233), .A2(n4773), .ZN(n5232) );
  INV_X1 U3941 ( .A(G468), .ZN(n4773) );
  NAND2_X1 U3942 ( .A1(n5234), .A2(n5235), .ZN(n5233) );
  NAND2_X1 U3943 ( .A1(G218), .A2(G3546), .ZN(n5235) );
  NAND2_X1 U3944 ( .A1(n5236), .A2(n4780), .ZN(n5234) );
  NAND2_X1 U3945 ( .A1(n5237), .A2(n5238), .ZN(n5236) );
  OR2_X1 U3946 ( .A1(G3550), .A2(KEYINPUT46), .ZN(n5238) );
  NAND2_X1 U3947 ( .A1(n5239), .A2(G468), .ZN(n5231) );
  NAND2_X1 U3948 ( .A1(n5240), .A2(n5241), .ZN(n5239) );
  NAND3_X1 U3949 ( .A1(KEYINPUT46), .A2(n5189), .A3(n4780), .ZN(n5241) );
  INV_X1 U3950 ( .A(G218), .ZN(n4780) );
  NAND2_X1 U3951 ( .A1(G218), .A2(n5190), .ZN(n5240) );
  NAND2_X1 U3952 ( .A1(n5242), .A2(n5243), .ZN(n5065) );
  NAND2_X1 U3953 ( .A1(n5244), .A2(n4836), .ZN(n5243) );
  NAND2_X1 U3954 ( .A1(n5245), .A2(n5246), .ZN(n5244) );
  NAND2_X1 U3955 ( .A1(G210), .A2(G3546), .ZN(n5246) );
  NAND2_X1 U3956 ( .A1(n5185), .A2(n4835), .ZN(n5245) );
  NAND2_X1 U3957 ( .A1(n5247), .A2(G457), .ZN(n5242) );
  NAND2_X1 U3958 ( .A1(n5248), .A2(n5249), .ZN(n5247) );
  NAND2_X1 U3959 ( .A1(n4835), .A2(n5189), .ZN(n5249) );
  INV_X1 U3960 ( .A(G210), .ZN(n4835) );
  NAND2_X1 U3961 ( .A1(G210), .A2(n5190), .ZN(n5248) );
  NAND2_X1 U3962 ( .A1(n5250), .A2(n5251), .ZN(n4558) );
  NAND2_X1 U3963 ( .A1(n5252), .A2(n4813), .ZN(n5251) );
  NAND2_X1 U3964 ( .A1(n5253), .A2(n5254), .ZN(n5252) );
  NAND2_X1 U3965 ( .A1(G3546), .A2(G281), .ZN(n5254) );
  NAND2_X1 U3966 ( .A1(n5185), .A2(n4818), .ZN(n5253) );
  NAND2_X1 U3967 ( .A1(n5255), .A2(G374), .ZN(n5250) );
  NAND2_X1 U3968 ( .A1(n5256), .A2(n5257), .ZN(n5255) );
  NAND2_X1 U3969 ( .A1(n4818), .A2(n5189), .ZN(n5257) );
  NAND2_X1 U3970 ( .A1(G281), .A2(n5190), .ZN(n5256) );
  INV_X1 U3971 ( .A(G549), .ZN(G606) );
  INV_X1 U3972 ( .A(G545), .ZN(G594) );
  NOR2_X1 U3973 ( .A1(G849), .A2(G850), .ZN(G601) );
  INV_X1 U3974 ( .A(G562), .ZN(G850) );
  INV_X1 U3975 ( .A(G552), .ZN(G849) );
  INV_X1 U3976 ( .A(G366), .ZN(G600) );
  INV_X1 U3977 ( .A(G348), .ZN(G599) );
  NOR4_X1 U3978 ( .A1(n5258), .A2(n5259), .A3(n4563), .A4(n4549), .ZN(G598) );
  AND2_X1 U3979 ( .A1(n5260), .A2(n5261), .ZN(n4549) );
  NAND2_X1 U3980 ( .A1(n5262), .A2(n4905), .ZN(n5261) );
  INV_X1 U3981 ( .A(G534), .ZN(n4905) );
  NAND2_X1 U3982 ( .A1(n5263), .A2(n5264), .ZN(n5262) );
  NAND2_X1 U3983 ( .A1(G3546), .A2(G351), .ZN(n5264) );
  NAND2_X1 U3984 ( .A1(n5185), .A2(n4909), .ZN(n5263) );
  NAND2_X1 U3985 ( .A1(n5265), .A2(G534), .ZN(n5260) );
  NAND2_X1 U3986 ( .A1(n5266), .A2(n5267), .ZN(n5265) );
  NAND2_X1 U3987 ( .A1(n4909), .A2(n5189), .ZN(n5267) );
  NAND2_X1 U3988 ( .A1(G351), .A2(n5190), .ZN(n5266) );
  INV_X1 U3989 ( .A(n4883), .ZN(n4563) );
  NAND2_X1 U3990 ( .A1(n5268), .A2(n5269), .ZN(n4883) );
  OR2_X1 U3991 ( .A1(n4709), .A2(G361), .ZN(n5269) );
  NAND2_X1 U3992 ( .A1(G248), .A2(G361), .ZN(n5268) );
  NAND3_X1 U3993 ( .A1(n5078), .A2(n5099), .A3(n5270), .ZN(n5259) );
  NAND2_X1 U3994 ( .A1(n5114), .A2(n5115), .ZN(n5270) );
  NAND3_X1 U3995 ( .A1(n5271), .A2(n5272), .A3(G503), .ZN(n5115) );
  NAND2_X1 U3996 ( .A1(G3550), .A2(n4897), .ZN(n5272) );
  NAND2_X1 U3997 ( .A1(G324), .A2(n5273), .ZN(n5271) );
  NAND3_X1 U3998 ( .A1(n5274), .A2(n5275), .A3(n4894), .ZN(n5114) );
  INV_X1 U3999 ( .A(G503), .ZN(n4894) );
  NAND2_X1 U4000 ( .A1(G324), .A2(n5276), .ZN(n5275) );
  NAND2_X1 U4001 ( .A1(n5237), .A2(n4897), .ZN(n5274) );
  NAND2_X1 U4002 ( .A1(n5277), .A2(n4868), .ZN(n5099) );
  NAND3_X1 U4003 ( .A1(n5278), .A2(n5279), .A3(G490), .ZN(n4868) );
  NAND2_X1 U4004 ( .A1(n4709), .A2(n4873), .ZN(n5279) );
  INV_X1 U4005 ( .A(G251), .ZN(n4709) );
  NAND2_X1 U4006 ( .A1(G316), .A2(n4707), .ZN(n5278) );
  NAND3_X1 U4007 ( .A1(n5280), .A2(n5281), .A3(n4872), .ZN(n5277) );
  NAND2_X1 U4008 ( .A1(n5282), .A2(n4873), .ZN(n5281) );
  NAND2_X1 U4009 ( .A1(n4748), .A2(n5283), .ZN(n5282) );
  OR2_X1 U4010 ( .A1(n4749), .A2(KEYINPUT65), .ZN(n5283) );
  NAND3_X1 U4011 ( .A1(KEYINPUT65), .A2(n4713), .A3(G316), .ZN(n5280) );
  NAND3_X1 U4012 ( .A1(n5284), .A2(n5285), .A3(n4867), .ZN(n5078) );
  NAND3_X1 U4013 ( .A1(G248), .A2(G308), .A3(G479), .ZN(n4867) );
  NAND2_X1 U4014 ( .A1(n5286), .A2(n4861), .ZN(n5285) );
  NAND2_X1 U4015 ( .A1(n5287), .A2(n5288), .ZN(n5286) );
  NAND2_X1 U4016 ( .A1(n4748), .A2(n4866), .ZN(n5288) );
  NAND2_X1 U4017 ( .A1(n4749), .A2(G308), .ZN(n5287) );
  INV_X1 U4018 ( .A(n4713), .ZN(n4749) );
  NAND3_X1 U4019 ( .A1(G251), .A2(n4866), .A3(G479), .ZN(n5284) );
  OR4_X1 U4020 ( .A1(n4269), .A2(n4505), .A3(n4850), .A4(n4528), .ZN(n5258) );
  AND2_X1 U4021 ( .A1(n5289), .A2(n5290), .ZN(n4528) );
  NAND2_X1 U4022 ( .A1(n5291), .A2(n4922), .ZN(n5290) );
  NAND2_X1 U4023 ( .A1(n5292), .A2(n5293), .ZN(n5291) );
  NAND2_X1 U4024 ( .A1(G3546), .A2(G341), .ZN(n5293) );
  NAND2_X1 U4025 ( .A1(n5185), .A2(n4917), .ZN(n5292) );
  INV_X1 U4026 ( .A(n5237), .ZN(n5185) );
  XOR2_X1 U4027 ( .A(KEYINPUT113), .B(G3548), .Z(n5237) );
  NAND2_X1 U4028 ( .A1(n5294), .A2(G523), .ZN(n5289) );
  NAND2_X1 U4029 ( .A1(n5295), .A2(n5296), .ZN(n5294) );
  NAND2_X1 U4030 ( .A1(n4917), .A2(n5189), .ZN(n5296) );
  INV_X1 U4031 ( .A(G3550), .ZN(n5189) );
  INV_X1 U4032 ( .A(G341), .ZN(n4917) );
  NAND2_X1 U4033 ( .A1(G341), .A2(n5190), .ZN(n5295) );
  NAND2_X1 U4034 ( .A1(n5297), .A2(n5298), .ZN(n4850) );
  OR2_X1 U4035 ( .A1(G251), .A2(G302), .ZN(n5298) );
  NAND2_X1 U4036 ( .A1(G302), .A2(n4707), .ZN(n5297) );
  INV_X1 U4037 ( .A(G248), .ZN(n4707) );
  NAND2_X1 U4038 ( .A1(n5299), .A2(n5300), .ZN(n4505) );
  NAND2_X1 U4039 ( .A1(n5276), .A2(n4888), .ZN(n5300) );
  INV_X1 U4040 ( .A(G3546), .ZN(n5276) );
  NAND2_X1 U4041 ( .A1(n5273), .A2(G514), .ZN(n5299) );
  INV_X1 U4042 ( .A(n5190), .ZN(n5273) );
  XOR2_X1 U4043 ( .A(KEYINPUT14), .B(G3552), .Z(n5190) );
  NAND2_X1 U4044 ( .A1(n5301), .A2(n5302), .ZN(n4269) );
  OR2_X1 U4045 ( .A1(n4748), .A2(G293), .ZN(n5302) );
  INV_X1 U4046 ( .A(G254), .ZN(n4748) );
  NAND2_X1 U4047 ( .A1(G293), .A2(n4713), .ZN(n5301) );
  XOR2_X1 U4048 ( .A(G242), .B(KEYINPUT74), .Z(n4713) );
  INV_X1 U4049 ( .A(G299), .ZN(G593) );
  NAND2_X1 U4050 ( .A1(n5157), .A2(n5303), .ZN(G591) );
  NAND2_X1 U4051 ( .A1(n4589), .A2(n5304), .ZN(n5303) );
  NAND3_X1 U4052 ( .A1(n5305), .A2(n4606), .A3(n5306), .ZN(n5304) );
  NAND2_X1 U4053 ( .A1(n4596), .A2(n4614), .ZN(n5306) );
  INV_X1 U4054 ( .A(n4608), .ZN(n4596) );
  NAND2_X1 U4055 ( .A1(n5307), .A2(n5308), .ZN(n4606) );
  XNOR2_X1 U4056 ( .A(KEYINPUT26), .B(n4836), .ZN(n5307) );
  NAND2_X1 U4057 ( .A1(n4602), .A2(n4619), .ZN(n5305) );
  NAND3_X1 U4058 ( .A1(n5309), .A2(n5310), .A3(n5311), .ZN(n4619) );
  NAND2_X1 U4059 ( .A1(n4663), .A2(n5312), .ZN(n5311) );
  NAND2_X1 U4060 ( .A1(n4691), .A2(n5313), .ZN(n5312) );
  NAND2_X1 U4061 ( .A1(n4645), .A2(n5314), .ZN(n5313) );
  NAND2_X1 U4062 ( .A1(n5315), .A2(n4694), .ZN(n5314) );
  NAND2_X1 U4063 ( .A1(n4696), .A2(n4662), .ZN(n4694) );
  NAND2_X1 U4064 ( .A1(KEYINPUT62), .A2(n5316), .ZN(n5315) );
  NAND2_X1 U4065 ( .A1(n5317), .A2(n5318), .ZN(n5309) );
  INV_X1 U4066 ( .A(KEYINPUT62), .ZN(n5318) );
  NAND2_X1 U4067 ( .A1(n5316), .A2(n5319), .ZN(n5317) );
  NOR3_X1 U4068 ( .A1(n5320), .A2(n4587), .A3(n4618), .ZN(G588) );
  NAND4_X1 U4069 ( .A1(n4696), .A2(n5319), .A3(n5321), .A4(n5322), .ZN(n4618) );
  XNOR2_X1 U4070 ( .A(KEYINPUT47), .B(n4674), .ZN(n5322) );
  AND2_X1 U4071 ( .A1(n4663), .A2(n4645), .ZN(n5319) );
  NAND2_X1 U4072 ( .A1(n5323), .A2(n5324), .ZN(n4645) );
  NAND2_X1 U4073 ( .A1(KEYINPUT17), .A2(n5325), .ZN(n5324) );
  NAND2_X1 U4074 ( .A1(n4691), .A2(n5326), .ZN(n5325) );
  NAND2_X1 U4075 ( .A1(n5327), .A2(n4703), .ZN(n5326) );
  NAND2_X1 U4076 ( .A1(n5328), .A2(n5329), .ZN(n5323) );
  INV_X1 U4077 ( .A(KEYINPUT17), .ZN(n5329) );
  XNOR2_X1 U4078 ( .A(n5327), .B(G389), .ZN(n5328) );
  AND2_X1 U4079 ( .A1(n5330), .A2(n5331), .ZN(n4663) );
  NAND2_X1 U4080 ( .A1(KEYINPUT1), .A2(n5332), .ZN(n5331) );
  NAND2_X1 U4081 ( .A1(n4799), .A2(n5333), .ZN(n5330) );
  NAND2_X1 U4082 ( .A1(KEYINPUT1), .A2(n5334), .ZN(n5333) );
  INV_X1 U4083 ( .A(n4647), .ZN(n4696) );
  INV_X1 U4084 ( .A(n4602), .ZN(n5320) );
  NOR2_X1 U4085 ( .A1(n4608), .A2(n4588), .ZN(n4602) );
  INV_X1 U4086 ( .A(n4613), .ZN(n4588) );
  NOR2_X1 U4087 ( .A1(n4591), .A2(n4629), .ZN(n4613) );
  INV_X1 U4088 ( .A(n4590), .ZN(n4629) );
  XOR2_X1 U4089 ( .A(n5335), .B(KEYINPUT119), .Z(n4590) );
  NAND3_X1 U4090 ( .A1(n5336), .A2(n5337), .A3(n5338), .ZN(n4608) );
  NAND3_X1 U4091 ( .A1(KEYINPUT39), .A2(n5339), .A3(n4836), .ZN(n5337) );
  INV_X1 U4092 ( .A(n5308), .ZN(n5339) );
  OR2_X1 U4093 ( .A1(n4836), .A2(KEYINPUT39), .ZN(n5336) );
  NOR4_X1 U4094 ( .A1(n5340), .A2(n5341), .A3(n5113), .A4(n5049), .ZN(G585) );
  INV_X1 U4095 ( .A(G623), .ZN(n5049) );
  XOR2_X1 U4096 ( .A(n4277), .B(n5142), .Z(G623) );
  NAND2_X1 U4097 ( .A1(n5342), .A2(n5343), .ZN(n5142) );
  NAND2_X1 U4098 ( .A1(G293), .A2(n5344), .ZN(n5343) );
  NAND2_X1 U4099 ( .A1(G332), .A2(G299), .ZN(n5342) );
  NAND2_X1 U4100 ( .A1(n5345), .A2(n5346), .ZN(n4277) );
  NAND2_X1 U4101 ( .A1(n5347), .A2(n5348), .ZN(n5346) );
  NAND2_X1 U4102 ( .A1(n5008), .A2(n5349), .ZN(n5348) );
  NAND2_X1 U4103 ( .A1(n5167), .A2(n5350), .ZN(n5349) );
  NAND2_X1 U4104 ( .A1(KEYINPUT77), .A2(n5351), .ZN(n5345) );
  NAND2_X1 U4105 ( .A1(n5008), .A2(n5352), .ZN(n5351) );
  NAND2_X1 U4106 ( .A1(n5167), .A2(n5353), .ZN(n5352) );
  XOR2_X1 U4107 ( .A(n5354), .B(n5177), .Z(n5113) );
  NAND2_X1 U4108 ( .A1(n5355), .A2(n5356), .ZN(n5354) );
  NAND2_X1 U4109 ( .A1(n4943), .A2(n5357), .ZN(n5356) );
  OR3_X1 U4110 ( .A1(n5100), .A2(n4529), .A3(n5060), .ZN(n5341) );
  XOR2_X1 U4111 ( .A(n5167), .B(n5353), .Z(n5060) );
  OR2_X1 U4112 ( .A1(n5350), .A2(n5358), .ZN(n5353) );
  NOR2_X1 U4113 ( .A1(n5174), .A2(n5347), .ZN(n5358) );
  NAND2_X1 U4114 ( .A1(n5359), .A2(n5360), .ZN(n5174) );
  NAND2_X1 U4115 ( .A1(n5139), .A2(n5169), .ZN(n5350) );
  NAND2_X1 U4116 ( .A1(n5359), .A2(n5032), .ZN(n5169) );
  XNOR2_X1 U4117 ( .A(n5008), .B(KEYINPUT37), .ZN(n5167) );
  INV_X1 U4118 ( .A(n4243), .ZN(n5008) );
  NAND2_X1 U4119 ( .A1(n5361), .A2(n5362), .ZN(n4243) );
  NAND2_X1 U4120 ( .A1(G302), .A2(n5344), .ZN(n5362) );
  NAND2_X1 U4121 ( .A1(G307), .A2(G332), .ZN(n5361) );
  XOR2_X1 U4122 ( .A(n5363), .B(n4946), .Z(n4529) );
  NAND3_X1 U4123 ( .A1(n4959), .A2(n5364), .A3(KEYINPUT102), .ZN(n5363) );
  NAND2_X1 U4124 ( .A1(n4948), .A2(G54), .ZN(n5364) );
  INV_X1 U4125 ( .A(n4957), .ZN(n4959) );
  XOR2_X1 U4126 ( .A(n5360), .B(n5365), .Z(n5100) );
  NAND2_X1 U4127 ( .A1(n5366), .A2(n5367), .ZN(n5360) );
  NAND2_X1 U4128 ( .A1(KEYINPUT36), .A2(n5154), .ZN(n5367) );
  OR2_X1 U4129 ( .A1(n5032), .A2(n5017), .ZN(n5154) );
  NAND2_X1 U4130 ( .A1(n5155), .A2(n5368), .ZN(n5366) );
  INV_X1 U4131 ( .A(KEYINPUT36), .ZN(n5368) );
  XNOR2_X1 U4132 ( .A(G490), .B(n4242), .ZN(n5155) );
  OR4_X1 U4133 ( .A1(n4564), .A2(n5076), .A3(n4507), .A4(n4548), .ZN(n5340) );
  XOR2_X1 U4134 ( .A(n5369), .B(n4948), .Z(n4548) );
  XOR2_X1 U4135 ( .A(n5357), .B(n4943), .Z(n4507) );
  NAND3_X1 U4136 ( .A1(n5370), .A2(n4954), .A3(n5371), .ZN(n5357) );
  NAND2_X1 U4137 ( .A1(n4946), .A2(n4957), .ZN(n5371) );
  NAND2_X1 U4138 ( .A1(n5372), .A2(G54), .ZN(n5370) );
  NAND2_X1 U4139 ( .A1(n5373), .A2(n5374), .ZN(n5076) );
  NAND2_X1 U4140 ( .A1(n5375), .A2(n5365), .ZN(n5374) );
  XNOR2_X1 U4141 ( .A(n5359), .B(n5017), .ZN(n5375) );
  NOR2_X1 U4142 ( .A1(n5376), .A2(G490), .ZN(n5017) );
  XOR2_X1 U4143 ( .A(KEYINPUT92), .B(n5377), .Z(n5373) );
  NOR2_X1 U4144 ( .A1(n5378), .A2(n5365), .ZN(n5377) );
  INV_X1 U4145 ( .A(n5347), .ZN(n5365) );
  NOR2_X1 U4146 ( .A1(n5173), .A2(n5379), .ZN(n5347) );
  AND3_X1 U4147 ( .A1(G54), .A2(n5177), .A3(n4936), .ZN(n5379) );
  NOR3_X1 U4148 ( .A1(n4944), .A2(n4235), .A3(n4945), .ZN(n4936) );
  INV_X1 U4149 ( .A(n5372), .ZN(n4944) );
  NOR2_X1 U4150 ( .A1(n4947), .A2(n4958), .ZN(n5372) );
  INV_X1 U4151 ( .A(n4948), .ZN(n4947) );
  NAND2_X1 U4152 ( .A1(n5128), .A2(n5380), .ZN(n5173) );
  NAND2_X1 U4153 ( .A1(n5381), .A2(n5177), .ZN(n5380) );
  NAND2_X1 U4154 ( .A1(n5382), .A2(n5383), .ZN(n5177) );
  NAND3_X1 U4155 ( .A1(n4230), .A2(n5128), .A3(KEYINPUT16), .ZN(n5383) );
  NAND2_X1 U4156 ( .A1(G503), .A2(n5384), .ZN(n5382) );
  NAND2_X1 U4157 ( .A1(n5385), .A2(KEYINPUT16), .ZN(n5384) );
  INV_X1 U4158 ( .A(n5128), .ZN(n5385) );
  NAND3_X1 U4159 ( .A1(n5131), .A2(n4977), .A3(n5355), .ZN(n5381) );
  NAND2_X1 U4160 ( .A1(n5386), .A2(n4231), .ZN(n5355) );
  XNOR2_X1 U4161 ( .A(KEYINPUT84), .B(n4888), .ZN(n5386) );
  INV_X1 U4162 ( .A(G514), .ZN(n4888) );
  INV_X1 U4163 ( .A(n4937), .ZN(n4977) );
  NOR2_X1 U4164 ( .A1(n4954), .A2(n4945), .ZN(n4937) );
  NAND3_X1 U4165 ( .A1(n4946), .A2(n4957), .A3(n4943), .ZN(n5131) );
  INV_X1 U4166 ( .A(n4945), .ZN(n4943) );
  XNOR2_X1 U4167 ( .A(G514), .B(n4231), .ZN(n4945) );
  NAND2_X1 U4168 ( .A1(n5387), .A2(n5388), .ZN(n4231) );
  NAND2_X1 U4169 ( .A1(G332), .A2(G338), .ZN(n5388) );
  NAND2_X1 U4170 ( .A1(n5389), .A2(n5390), .ZN(n4957) );
  NAND2_X1 U4171 ( .A1(n4948), .A2(n4235), .ZN(n5390) );
  XOR2_X1 U4172 ( .A(G534), .B(n4233), .Z(n4948) );
  NAND2_X1 U4173 ( .A1(G534), .A2(n4233), .ZN(n5389) );
  NAND2_X1 U4174 ( .A1(n5391), .A2(n5392), .ZN(n4233) );
  NAND2_X1 U4175 ( .A1(G332), .A2(G358), .ZN(n5392) );
  XOR2_X1 U4176 ( .A(KEYINPUT50), .B(n5393), .Z(n5391) );
  NOR2_X1 U4177 ( .A1(n5387), .A2(n4909), .ZN(n5393) );
  INV_X1 U4178 ( .A(n4958), .ZN(n4946) );
  NAND2_X1 U4179 ( .A1(n4954), .A2(n5394), .ZN(n4958) );
  NAND2_X1 U4180 ( .A1(n4232), .A2(n4922), .ZN(n5394) );
  INV_X1 U4181 ( .A(n4960), .ZN(n4954) );
  NOR2_X1 U4182 ( .A1(n4922), .A2(n4232), .ZN(n4960) );
  AND2_X1 U4183 ( .A1(n5395), .A2(n5396), .ZN(n4232) );
  NAND2_X1 U4184 ( .A1(G341), .A2(n4238), .ZN(n5396) );
  NAND2_X1 U4185 ( .A1(G332), .A2(G348), .ZN(n5395) );
  INV_X1 U4186 ( .A(G523), .ZN(n4922) );
  NAND2_X1 U4187 ( .A1(G503), .A2(n4230), .ZN(n5128) );
  NAND2_X1 U4188 ( .A1(n5397), .A2(n5398), .ZN(n4230) );
  NAND2_X1 U4189 ( .A1(G324), .A2(n5344), .ZN(n5398) );
  NAND2_X1 U4190 ( .A1(G331), .A2(G332), .ZN(n5397) );
  XNOR2_X1 U4191 ( .A(n5359), .B(n5032), .ZN(n5378) );
  NOR2_X1 U4192 ( .A1(n4872), .A2(n4242), .ZN(n5032) );
  INV_X1 U4193 ( .A(n5376), .ZN(n4242) );
  NAND2_X1 U4194 ( .A1(n5399), .A2(n5400), .ZN(n5376) );
  NAND2_X1 U4195 ( .A1(G316), .A2(n5344), .ZN(n5400) );
  NAND2_X1 U4196 ( .A1(G323), .A2(G332), .ZN(n5399) );
  INV_X1 U4197 ( .A(G490), .ZN(n4872) );
  INV_X1 U4198 ( .A(n5149), .ZN(n5359) );
  NAND2_X1 U4199 ( .A1(n5139), .A2(n5401), .ZN(n5149) );
  NAND2_X1 U4200 ( .A1(n4244), .A2(n4861), .ZN(n5401) );
  INV_X1 U4201 ( .A(G479), .ZN(n4861) );
  INV_X1 U4202 ( .A(n5140), .ZN(n4244) );
  NAND2_X1 U4203 ( .A1(G479), .A2(n5140), .ZN(n5139) );
  NAND2_X1 U4204 ( .A1(n5402), .A2(n5403), .ZN(n5140) );
  NAND2_X1 U4205 ( .A1(G308), .A2(n5344), .ZN(n5403) );
  INV_X1 U4206 ( .A(G332), .ZN(n5344) );
  NAND2_X1 U4207 ( .A1(G315), .A2(G332), .ZN(n5402) );
  NAND2_X1 U4208 ( .A1(n5404), .A2(n5369), .ZN(n4564) );
  NAND2_X1 U4209 ( .A1(n4984), .A2(n5405), .ZN(n5369) );
  INV_X1 U4210 ( .A(G54), .ZN(n5405) );
  INV_X1 U4211 ( .A(n4235), .ZN(n4984) );
  XOR2_X1 U4212 ( .A(n5406), .B(KEYINPUT90), .Z(n5404) );
  NAND2_X1 U4213 ( .A1(G54), .A2(n4235), .ZN(n5406) );
  NAND2_X1 U4214 ( .A1(n5407), .A2(n5408), .ZN(n4235) );
  NAND2_X1 U4215 ( .A1(G361), .A2(n5409), .ZN(n5408) );
  XNOR2_X1 U4216 ( .A(KEYINPUT69), .B(n5387), .ZN(n5409) );
  INV_X1 U4217 ( .A(n4238), .ZN(n5387) );
  XOR2_X1 U4218 ( .A(G332), .B(KEYINPUT9), .Z(n4238) );
  NAND2_X1 U4219 ( .A1(G332), .A2(G366), .ZN(n5407) );
  NOR4_X1 U4220 ( .A1(n5410), .A2(n5411), .A3(n4559), .A4(n5042), .ZN(G575) );
  NAND2_X1 U4221 ( .A1(n5412), .A2(n5413), .ZN(n5042) );
  NAND2_X1 U4222 ( .A1(n5414), .A2(n5415), .ZN(n5413) );
  XNOR2_X1 U4223 ( .A(n5159), .B(n5416), .ZN(n5414) );
  NOR2_X1 U4224 ( .A1(n5126), .A2(n5164), .ZN(n5416) );
  AND3_X1 U4225 ( .A1(n5417), .A2(n5335), .A3(n4592), .ZN(n5126) );
  NAND2_X1 U4226 ( .A1(n5418), .A2(n5419), .ZN(n5412) );
  XNOR2_X1 U4227 ( .A(n5420), .B(n5164), .ZN(n5418) );
  NAND2_X1 U4228 ( .A1(n5421), .A2(n5338), .ZN(n5164) );
  NAND2_X1 U4229 ( .A1(G457), .A2(n5308), .ZN(n5338) );
  NAND2_X1 U4230 ( .A1(n5417), .A2(n4614), .ZN(n5421) );
  NAND2_X1 U4231 ( .A1(KEYINPUT27), .A2(n5422), .ZN(n5420) );
  XNOR2_X1 U4232 ( .A(KEYINPUT91), .B(n5122), .ZN(n5422) );
  INV_X1 U4233 ( .A(n5159), .ZN(n5122) );
  XOR2_X1 U4234 ( .A(n4589), .B(KEYINPUT56), .Z(n5159) );
  INV_X1 U4235 ( .A(n4587), .ZN(n4589) );
  NAND2_X1 U4236 ( .A1(n5157), .A2(n5423), .ZN(n4587) );
  OR2_X1 U4237 ( .A1(n5424), .A2(G446), .ZN(n5423) );
  NAND2_X1 U4238 ( .A1(G446), .A2(n5424), .ZN(n5157) );
  XNOR2_X1 U4239 ( .A(n4674), .B(G4), .ZN(n4559) );
  NAND3_X1 U4240 ( .A1(n5425), .A2(n5426), .A3(n5427), .ZN(n5411) );
  INV_X1 U4241 ( .A(n4521), .ZN(n5427) );
  XOR2_X1 U4242 ( .A(n5428), .B(n5429), .Z(n4521) );
  OR2_X1 U4243 ( .A1(n4662), .A2(n5430), .ZN(n5428) );
  NAND3_X1 U4244 ( .A1(n4543), .A2(n4544), .A3(n4542), .ZN(n5426) );
  NAND3_X1 U4245 ( .A1(n5431), .A2(n4661), .A3(n4673), .ZN(n4542) );
  NAND2_X1 U4246 ( .A1(G4), .A2(n4695), .ZN(n5431) );
  INV_X1 U4247 ( .A(n4674), .ZN(n4695) );
  NAND2_X1 U4248 ( .A1(n5066), .A2(n5067), .ZN(n5425) );
  NAND2_X1 U4249 ( .A1(n5432), .A2(n5415), .ZN(n5067) );
  XNOR2_X1 U4250 ( .A(n5433), .B(n5417), .ZN(n5432) );
  NOR2_X1 U4251 ( .A1(KEYINPUT96), .A2(n5434), .ZN(n5433) );
  NOR2_X1 U4252 ( .A1(n5435), .A2(n4614), .ZN(n5434) );
  AND2_X1 U4253 ( .A1(n5335), .A2(n4592), .ZN(n5435) );
  NAND2_X1 U4254 ( .A1(n5419), .A2(n5436), .ZN(n5066) );
  XNOR2_X1 U4255 ( .A(n5417), .B(n4614), .ZN(n5436) );
  NAND2_X1 U4256 ( .A1(n4607), .A2(n5437), .ZN(n4614) );
  NAND2_X1 U4257 ( .A1(n5438), .A2(n4592), .ZN(n5437) );
  XNOR2_X1 U4258 ( .A(n4836), .B(n5308), .ZN(n5417) );
  INV_X1 U4259 ( .A(G457), .ZN(n4836) );
  OR4_X1 U4260 ( .A1(n5439), .A2(n4498), .A3(n5108), .A4(n5082), .ZN(n5410) );
  NAND2_X1 U4261 ( .A1(n5440), .A2(n5441), .ZN(n5082) );
  NAND2_X1 U4262 ( .A1(n5419), .A2(n4627), .ZN(n5441) );
  XNOR2_X1 U4263 ( .A(n4592), .B(n4634), .ZN(n4627) );
  XOR2_X1 U4264 ( .A(n5442), .B(KEYINPUT117), .Z(n5440) );
  NAND2_X1 U4265 ( .A1(n5443), .A2(n5415), .ZN(n5442) );
  INV_X1 U4266 ( .A(n5419), .ZN(n5415) );
  XNOR2_X1 U4267 ( .A(n4592), .B(n4611), .ZN(n5443) );
  INV_X1 U4268 ( .A(n4591), .ZN(n4592) );
  NAND2_X1 U4269 ( .A1(n4607), .A2(n5444), .ZN(n4591) );
  OR2_X1 U4270 ( .A1(n5445), .A2(G468), .ZN(n5444) );
  NAND2_X1 U4271 ( .A1(G468), .A2(n5445), .ZN(n4607) );
  NAND2_X1 U4272 ( .A1(n5446), .A2(n5447), .ZN(n5108) );
  NAND2_X1 U4273 ( .A1(n5448), .A2(n5449), .ZN(n5447) );
  XNOR2_X1 U4274 ( .A(KEYINPUT88), .B(n5450), .ZN(n5448) );
  NAND2_X1 U4275 ( .A1(n5451), .A2(n5125), .ZN(n5446) );
  XOR2_X1 U4276 ( .A(n5450), .B(KEYINPUT59), .Z(n5451) );
  NAND2_X1 U4277 ( .A1(n4691), .A2(n5452), .ZN(n5450) );
  NAND2_X1 U4278 ( .A1(n5453), .A2(n5454), .ZN(n5452) );
  NAND2_X1 U4279 ( .A1(n5455), .A2(n5456), .ZN(n4498) );
  NAND2_X1 U4280 ( .A1(n5123), .A2(n5453), .ZN(n5456) );
  XOR2_X1 U4281 ( .A(KEYINPUT13), .B(n5457), .Z(n5455) );
  NOR2_X1 U4282 ( .A1(n5123), .A2(n5453), .ZN(n5457) );
  NAND2_X1 U4283 ( .A1(n5458), .A2(n5459), .ZN(n5453) );
  NAND2_X1 U4284 ( .A1(n5430), .A2(n5429), .ZN(n5459) );
  INV_X1 U4285 ( .A(n4543), .ZN(n5430) );
  INV_X1 U4286 ( .A(n5460), .ZN(n5458) );
  XNOR2_X1 U4287 ( .A(n5092), .B(KEYINPUT75), .ZN(n5439) );
  XNOR2_X1 U4288 ( .A(n5335), .B(n5419), .ZN(n5092) );
  NOR2_X1 U4289 ( .A1(n5163), .A2(n5461), .ZN(n5419) );
  NOR4_X1 U4290 ( .A1(n5449), .A2(n4543), .A3(n5124), .A4(n5123), .ZN(n5461) );
  INV_X1 U4291 ( .A(n5454), .ZN(n5123) );
  INV_X1 U4292 ( .A(n5429), .ZN(n5124) );
  NAND2_X1 U4293 ( .A1(G4), .A2(n4683), .ZN(n4543) );
  NOR2_X1 U4294 ( .A1(n4674), .A2(n4673), .ZN(n4683) );
  INV_X1 U4295 ( .A(n5321), .ZN(n4673) );
  NAND2_X1 U4296 ( .A1(n4661), .A2(n4685), .ZN(n4674) );
  NAND2_X1 U4297 ( .A1(n5462), .A2(n4813), .ZN(n4685) );
  INV_X1 U4298 ( .A(n5463), .ZN(n4661) );
  NAND2_X1 U4299 ( .A1(n5310), .A2(n5464), .ZN(n5163) );
  NAND2_X1 U4300 ( .A1(n5125), .A2(n5465), .ZN(n5464) );
  NAND2_X1 U4301 ( .A1(n4691), .A2(n5466), .ZN(n5465) );
  NAND2_X1 U4302 ( .A1(n5460), .A2(n5454), .ZN(n5466) );
  NAND2_X1 U4303 ( .A1(n5467), .A2(n5468), .ZN(n5454) );
  NAND2_X1 U4304 ( .A1(n5469), .A2(n4703), .ZN(n5468) );
  INV_X1 U4305 ( .A(G389), .ZN(n4703) );
  XOR2_X1 U4306 ( .A(n5470), .B(KEYINPUT51), .Z(n5467) );
  NAND2_X1 U4307 ( .A1(n5327), .A2(G389), .ZN(n5470) );
  INV_X1 U4308 ( .A(n5469), .ZN(n5327) );
  NAND2_X1 U4309 ( .A1(n4693), .A2(n5471), .ZN(n5460) );
  NAND2_X1 U4310 ( .A1(n5429), .A2(n4662), .ZN(n5471) );
  NAND2_X1 U4311 ( .A1(n4544), .A2(n5472), .ZN(n4662) );
  NAND2_X1 U4312 ( .A1(G411), .A2(n5473), .ZN(n5472) );
  NAND2_X1 U4313 ( .A1(n5463), .A2(n5321), .ZN(n4544) );
  XOR2_X1 U4314 ( .A(G411), .B(n5473), .Z(n5321) );
  NOR2_X1 U4315 ( .A1(n5462), .A2(n4813), .ZN(n5463) );
  INV_X1 U4316 ( .A(G374), .ZN(n4813) );
  NAND2_X1 U4317 ( .A1(n5474), .A2(n5475), .ZN(n5429) );
  NAND2_X1 U4318 ( .A1(KEYINPUT82), .A2(n4647), .ZN(n5475) );
  NAND2_X1 U4319 ( .A1(n4693), .A2(n5476), .ZN(n4647) );
  NAND2_X1 U4320 ( .A1(n5477), .A2(n4722), .ZN(n5476) );
  NAND2_X1 U4321 ( .A1(n5478), .A2(n5479), .ZN(n5474) );
  INV_X1 U4322 ( .A(KEYINPUT82), .ZN(n5479) );
  XNOR2_X1 U4323 ( .A(G400), .B(n5477), .ZN(n5478) );
  INV_X1 U4324 ( .A(n5316), .ZN(n4693) );
  NOR2_X1 U4325 ( .A1(n5477), .A2(n4722), .ZN(n5316) );
  INV_X1 U4326 ( .A(G400), .ZN(n4722) );
  NAND2_X1 U4327 ( .A1(G389), .A2(n5469), .ZN(n4691) );
  INV_X1 U4328 ( .A(n5449), .ZN(n5125) );
  NAND2_X1 U4329 ( .A1(n5310), .A2(n5480), .ZN(n5449) );
  NAND2_X1 U4330 ( .A1(n5481), .A2(n4799), .ZN(n5480) );
  INV_X1 U4331 ( .A(n5332), .ZN(n5310) );
  NOR2_X1 U4332 ( .A1(n4799), .A2(n5481), .ZN(n5332) );
  INV_X1 U4333 ( .A(G435), .ZN(n4799) );
  NOR2_X1 U4334 ( .A1(n4611), .A2(n5438), .ZN(n5335) );
  INV_X1 U4335 ( .A(n4634), .ZN(n5438) );
  NAND2_X1 U4336 ( .A1(G422), .A2(n5482), .ZN(n4634) );
  NOR2_X1 U4337 ( .A1(n5482), .A2(G422), .ZN(n4611) );
  XNOR2_X1 U4338 ( .A(n4247), .B(KEYINPUT109), .ZN(G1004) );
  AND2_X1 U4339 ( .A1(n5483), .A2(n5484), .ZN(n4247) );
  NAND2_X1 U4340 ( .A1(n5485), .A2(n5486), .ZN(n5484) );
  XNOR2_X1 U4341 ( .A(n5487), .B(n5488), .ZN(n5485) );
  XOR2_X1 U4342 ( .A(n5489), .B(KEYINPUT55), .Z(n5483) );
  NAND2_X1 U4343 ( .A1(n5490), .A2(n5491), .ZN(n5489) );
  INV_X1 U4344 ( .A(n5486), .ZN(n5491) );
  XNOR2_X1 U4345 ( .A(n5492), .B(n5493), .ZN(n5486) );
  XNOR2_X1 U4346 ( .A(n4747), .B(G218), .ZN(n5493) );
  INV_X1 U4347 ( .A(G226), .ZN(n4747) );
  XNOR2_X1 U4348 ( .A(G206), .B(G210), .ZN(n5492) );
  XNOR2_X1 U4349 ( .A(n5488), .B(n5494), .ZN(n5490) );
  INV_X1 U4350 ( .A(n5487), .ZN(n5494) );
  XNOR2_X1 U4351 ( .A(n5495), .B(n5496), .ZN(n5487) );
  XNOR2_X1 U4352 ( .A(n4708), .B(G234), .ZN(n5496) );
  INV_X1 U4353 ( .A(G257), .ZN(n4708) );
  NAND2_X1 U4354 ( .A1(n5497), .A2(n5498), .ZN(n5495) );
  NAND2_X1 U4355 ( .A1(G273), .A2(n4730), .ZN(n5498) );
  XOR2_X1 U4356 ( .A(KEYINPUT120), .B(n5499), .Z(n5497) );
  NOR2_X1 U4357 ( .A1(G273), .A2(n4730), .ZN(n5499) );
  XNOR2_X1 U4358 ( .A(G289), .B(G281), .ZN(n5488) );
  XOR2_X1 U4359 ( .A(n5500), .B(n5501), .Z(G1002) );
  XNOR2_X1 U4360 ( .A(n4909), .B(G341), .ZN(n5501) );
  INV_X1 U4361 ( .A(G351), .ZN(n4909) );
  XOR2_X1 U4362 ( .A(n5502), .B(G302), .Z(n5500) );
  XOR2_X1 U4363 ( .A(n5503), .B(n5504), .Z(n5502) );
  XNOR2_X1 U4364 ( .A(n4897), .B(n5505), .ZN(n5504) );
  XOR2_X1 U4365 ( .A(G369), .B(G361), .Z(n5505) );
  INV_X1 U4366 ( .A(G324), .ZN(n4897) );
  XOR2_X1 U4367 ( .A(n5506), .B(n5507), .Z(n5503) );
  XNOR2_X1 U4368 ( .A(n4866), .B(G293), .ZN(n5507) );
  INV_X1 U4369 ( .A(G308), .ZN(n4866) );
  NAND2_X1 U4370 ( .A1(KEYINPUT3), .A2(n5508), .ZN(n5506) );
  XNOR2_X1 U4371 ( .A(KEYINPUT76), .B(n4873), .ZN(n5508) );
  INV_X1 U4372 ( .A(G316), .ZN(n4873) );
  XNOR2_X1 U4373 ( .A(n5509), .B(n5510), .ZN(G1000) );
  XOR2_X1 U4374 ( .A(n5511), .B(n5512), .Z(n5510) );
  XOR2_X1 U4375 ( .A(n5477), .B(n5473), .Z(n5512) );
  NAND2_X1 U4376 ( .A1(n5513), .A2(n5514), .ZN(n5473) );
  NAND2_X1 U4377 ( .A1(G273), .A2(n5515), .ZN(n5514) );
  NAND2_X1 U4378 ( .A1(G280), .A2(G335), .ZN(n5513) );
  NAND2_X1 U4379 ( .A1(n5516), .A2(n5517), .ZN(n5477) );
  OR2_X1 U4380 ( .A1(G272), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U4381 ( .A1(n4730), .A2(n5515), .ZN(n5516) );
  INV_X1 U4382 ( .A(G265), .ZN(n4730) );
  XNOR2_X1 U4383 ( .A(n5481), .B(n5469), .ZN(n5511) );
  NAND2_X1 U4384 ( .A1(n5518), .A2(n5519), .ZN(n5469) );
  NAND2_X1 U4385 ( .A1(G257), .A2(n5515), .ZN(n5519) );
  NAND2_X1 U4386 ( .A1(G264), .A2(G335), .ZN(n5518) );
  INV_X1 U4387 ( .A(n5334), .ZN(n5481) );
  NAND2_X1 U4388 ( .A1(n5520), .A2(n5521), .ZN(n5334) );
  NAND2_X1 U4389 ( .A1(G234), .A2(n5515), .ZN(n5521) );
  XOR2_X1 U4390 ( .A(n5522), .B(KEYINPUT44), .Z(n5520) );
  NAND2_X1 U4391 ( .A1(G241), .A2(G335), .ZN(n5522) );
  XOR2_X1 U4392 ( .A(n5523), .B(n5524), .Z(n5509) );
  XOR2_X1 U4393 ( .A(n5462), .B(n5482), .Z(n5524) );
  NAND2_X1 U4394 ( .A1(n5525), .A2(n5526), .ZN(n5482) );
  NAND2_X1 U4395 ( .A1(G226), .A2(n5515), .ZN(n5526) );
  NAND2_X1 U4396 ( .A1(G233), .A2(G335), .ZN(n5525) );
  NAND2_X1 U4397 ( .A1(n5527), .A2(n5528), .ZN(n5462) );
  OR2_X1 U4398 ( .A1(G288), .A2(n5515), .ZN(n5528) );
  NAND2_X1 U4399 ( .A1(n4818), .A2(n5515), .ZN(n5527) );
  INV_X1 U4400 ( .A(G281), .ZN(n4818) );
  XNOR2_X1 U4401 ( .A(n5529), .B(n5308), .ZN(n5523) );
  NAND2_X1 U4402 ( .A1(n5530), .A2(n5531), .ZN(n5308) );
  NAND2_X1 U4403 ( .A1(G210), .A2(n5515), .ZN(n5531) );
  NAND2_X1 U4404 ( .A1(G217), .A2(G335), .ZN(n5530) );
  NAND2_X1 U4405 ( .A1(n5532), .A2(n5533), .ZN(n5529) );
  NAND2_X1 U4406 ( .A1(n5534), .A2(n5515), .ZN(n5533) );
  XOR2_X1 U4407 ( .A(G289), .B(n5535), .Z(n5534) );
  NAND2_X1 U4408 ( .A1(n5536), .A2(G335), .ZN(n5532) );
  XOR2_X1 U4409 ( .A(G292), .B(n5535), .Z(n5536) );
  XNOR2_X1 U4410 ( .A(n5445), .B(n5537), .ZN(n5535) );
  NOR2_X1 U4411 ( .A1(KEYINPUT45), .A2(n5424), .ZN(n5537) );
  NAND2_X1 U4412 ( .A1(n5538), .A2(n5539), .ZN(n5424) );
  NAND2_X1 U4413 ( .A1(G206), .A2(n5515), .ZN(n5539) );
  NAND2_X1 U4414 ( .A1(G209), .A2(G335), .ZN(n5538) );
  NAND2_X1 U4415 ( .A1(n5540), .A2(n5541), .ZN(n5445) );
  NAND2_X1 U4416 ( .A1(G218), .A2(n5515), .ZN(n5541) );
  INV_X1 U4417 ( .A(G335), .ZN(n5515) );
  NAND2_X1 U4418 ( .A1(G225), .A2(G335), .ZN(n5540) );
endmodule

