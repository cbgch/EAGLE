//Key = 0100001100011001011001011011001100001011101001000101101111110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;

XNOR2_X1 U751 ( .A(G107), .B(n1043), .ZN(G9) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
AND4_X1 U754 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1048) );
OR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
NOR2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR3_X1 U757 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
AND2_X1 U758 ( .A1(n1061), .A2(KEYINPUT4), .ZN(n1060) );
NOR2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1058) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1054) );
INV_X1 U761 ( .A(n1061), .ZN(n1065) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR3_X1 U763 ( .A1(n1068), .A2(KEYINPUT4), .A3(n1069), .ZN(n1066) );
NAND3_X1 U764 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1046) );
NAND4_X1 U765 ( .A1(n1061), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1072) );
NAND2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND3_X1 U767 ( .A1(n1052), .A2(n1078), .A3(KEYINPUT34), .ZN(n1076) );
NAND3_X1 U768 ( .A1(n1079), .A2(n1080), .A3(n1053), .ZN(n1074) );
INV_X1 U769 ( .A(n1077), .ZN(n1053) );
NAND2_X1 U770 ( .A1(n1051), .A2(n1081), .ZN(n1080) );
OR2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1052), .A2(n1084), .ZN(n1079) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
OR2_X1 U774 ( .A1(n1087), .A2(KEYINPUT34), .ZN(n1086) );
AND3_X1 U775 ( .A1(n1070), .A2(n1071), .A3(n1088), .ZN(n1044) );
NAND4_X1 U776 ( .A1(n1089), .A2(n1073), .A3(n1090), .A4(n1091), .ZN(n1070) );
NOR4_X1 U777 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
XOR2_X1 U778 ( .A(n1096), .B(KEYINPUT30), .Z(n1094) );
NAND2_X1 U779 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U780 ( .A1(n1097), .A2(n1098), .ZN(n1093) );
XOR2_X1 U781 ( .A(n1099), .B(KEYINPUT28), .Z(n1098) );
XOR2_X1 U782 ( .A(G478), .B(KEYINPUT57), .Z(n1097) );
NOR2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1090) );
XNOR2_X1 U784 ( .A(n1102), .B(n1103), .ZN(n1089) );
XOR2_X1 U785 ( .A(n1104), .B(n1105), .Z(G72) );
NOR2_X1 U786 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U787 ( .A(KEYINPUT20), .B(n1108), .Z(n1107) );
NOR3_X1 U788 ( .A1(n1109), .A2(n1110), .A3(n1047), .ZN(n1108) );
NOR2_X1 U789 ( .A1(G900), .A2(n1071), .ZN(n1110) );
AND3_X1 U790 ( .A1(n1109), .A2(n1071), .A3(n1047), .ZN(n1106) );
XNOR2_X1 U791 ( .A(n1111), .B(n1112), .ZN(n1109) );
NAND2_X1 U792 ( .A1(G953), .A2(n1113), .ZN(n1104) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1114), .A2(n1115), .ZN(G69) );
NAND2_X1 U795 ( .A1(n1116), .A2(n1071), .ZN(n1115) );
XNOR2_X1 U796 ( .A(n1049), .B(n1117), .ZN(n1116) );
NAND2_X1 U797 ( .A1(n1118), .A2(G953), .ZN(n1114) );
NAND2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U799 ( .A1(n1117), .A2(n1121), .ZN(n1120) );
NAND2_X1 U800 ( .A1(G224), .A2(n1122), .ZN(n1119) );
NAND2_X1 U801 ( .A1(G898), .A2(n1117), .ZN(n1122) );
NAND3_X1 U802 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1117) );
XOR2_X1 U803 ( .A(n1126), .B(KEYINPUT14), .Z(n1125) );
OR2_X1 U804 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U805 ( .A1(n1128), .A2(n1127), .ZN(n1124) );
NAND2_X1 U806 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
XNOR2_X1 U807 ( .A(KEYINPUT62), .B(n1131), .ZN(n1129) );
NAND2_X1 U808 ( .A1(G953), .A2(n1132), .ZN(n1123) );
NOR3_X1 U809 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1136), .A2(n1071), .A3(n1088), .ZN(n1135) );
INV_X1 U811 ( .A(G952), .ZN(n1088) );
AND2_X1 U812 ( .A1(n1136), .A2(n1137), .ZN(n1134) );
INV_X1 U813 ( .A(KEYINPUT32), .ZN(n1136) );
XOR2_X1 U814 ( .A(n1138), .B(n1139), .Z(n1133) );
NAND2_X1 U815 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NOR2_X1 U816 ( .A1(n1137), .A2(n1142), .ZN(G63) );
NOR3_X1 U817 ( .A1(n1099), .A2(n1143), .A3(n1144), .ZN(n1142) );
NOR3_X1 U818 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
AND2_X1 U819 ( .A1(n1145), .A2(n1147), .ZN(n1143) );
NAND3_X1 U820 ( .A1(G478), .A2(n1148), .A3(KEYINPUT54), .ZN(n1147) );
NOR3_X1 U821 ( .A1(n1149), .A2(n1137), .A3(n1150), .ZN(G60) );
NOR4_X1 U822 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
NOR2_X1 U823 ( .A1(KEYINPUT6), .A2(n1155), .ZN(n1152) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
INV_X1 U825 ( .A(KEYINPUT6), .ZN(n1157) );
NOR2_X1 U826 ( .A1(n1158), .A2(n1156), .ZN(n1149) );
NOR2_X1 U827 ( .A1(KEYINPUT61), .A2(n1155), .ZN(n1156) );
NOR2_X1 U828 ( .A1(n1153), .A2(n1154), .ZN(n1158) );
XNOR2_X1 U829 ( .A(n1159), .B(n1160), .ZN(G6) );
NOR3_X1 U830 ( .A1(n1161), .A2(KEYINPUT5), .A3(n1162), .ZN(n1160) );
NOR2_X1 U831 ( .A1(n1137), .A2(n1163), .ZN(G57) );
XOR2_X1 U832 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U833 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
NAND3_X1 U834 ( .A1(n1168), .A2(G472), .A3(n1140), .ZN(n1167) );
XOR2_X1 U835 ( .A(n1169), .B(KEYINPUT53), .Z(n1166) );
NAND2_X1 U836 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U837 ( .A(n1172), .B(KEYINPUT25), .Z(n1171) );
NAND2_X1 U838 ( .A1(n1140), .A2(G472), .ZN(n1172) );
XNOR2_X1 U839 ( .A(KEYINPUT22), .B(n1168), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1137), .A2(n1173), .ZN(G54) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U842 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U843 ( .A1(n1140), .A2(G469), .ZN(n1177) );
NAND2_X1 U844 ( .A1(KEYINPUT49), .A2(n1178), .ZN(n1176) );
XOR2_X1 U845 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U846 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U847 ( .A1(KEYINPUT0), .A2(n1183), .ZN(n1182) );
XNOR2_X1 U848 ( .A(KEYINPUT9), .B(n1184), .ZN(n1183) );
XNOR2_X1 U849 ( .A(KEYINPUT16), .B(n1185), .ZN(n1179) );
INV_X1 U850 ( .A(G110), .ZN(n1185) );
NOR2_X1 U851 ( .A1(n1137), .A2(n1186), .ZN(G51) );
XOR2_X1 U852 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U853 ( .A(n1189), .B(KEYINPUT47), .Z(n1188) );
NAND2_X1 U854 ( .A1(n1140), .A2(G210), .ZN(n1189) );
INV_X1 U855 ( .A(n1154), .ZN(n1140) );
NAND2_X1 U856 ( .A1(G902), .A2(n1148), .ZN(n1154) );
NAND2_X1 U857 ( .A1(n1190), .A2(n1191), .ZN(n1148) );
INV_X1 U858 ( .A(n1049), .ZN(n1191) );
NAND4_X1 U859 ( .A1(n1192), .A2(n1043), .A3(n1193), .A4(n1194), .ZN(n1049) );
NOR3_X1 U860 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
NOR2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR2_X1 U862 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
NOR2_X1 U863 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U864 ( .A(n1078), .B(KEYINPUT33), .ZN(n1202) );
NOR2_X1 U865 ( .A1(n1204), .A2(n1205), .ZN(n1200) );
XOR2_X1 U866 ( .A(n1051), .B(KEYINPUT36), .Z(n1205) );
INV_X1 U867 ( .A(n1206), .ZN(n1196) );
NOR2_X1 U868 ( .A1(n1207), .A2(n1162), .ZN(n1195) );
NOR2_X1 U869 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XNOR2_X1 U870 ( .A(KEYINPUT37), .B(n1161), .ZN(n1209) );
NAND3_X1 U871 ( .A1(n1210), .A2(n1051), .A3(n1082), .ZN(n1161) );
NAND4_X1 U872 ( .A1(n1067), .A2(n1083), .A3(n1210), .A4(n1051), .ZN(n1043) );
INV_X1 U873 ( .A(n1047), .ZN(n1190) );
NAND4_X1 U874 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1047) );
NOR3_X1 U875 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
INV_X1 U876 ( .A(n1218), .ZN(n1216) );
NOR2_X1 U877 ( .A1(n1219), .A2(n1220), .ZN(n1215) );
NOR2_X1 U878 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
NOR2_X1 U879 ( .A1(n1223), .A2(n1087), .ZN(n1222) );
NOR2_X1 U880 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NOR2_X1 U881 ( .A1(n1203), .A2(n1057), .ZN(n1225) );
NOR2_X1 U882 ( .A1(n1226), .A2(n1204), .ZN(n1224) );
XNOR2_X1 U883 ( .A(n1067), .B(KEYINPUT50), .ZN(n1226) );
NOR3_X1 U884 ( .A1(n1227), .A2(n1057), .A3(n1085), .ZN(n1221) );
INV_X1 U885 ( .A(n1073), .ZN(n1057) );
XOR2_X1 U886 ( .A(KEYINPUT1), .B(n1082), .Z(n1227) );
NOR2_X1 U887 ( .A1(n1071), .A2(G952), .ZN(n1137) );
NAND2_X1 U888 ( .A1(n1228), .A2(n1229), .ZN(G48) );
NAND2_X1 U889 ( .A1(G146), .A2(n1230), .ZN(n1229) );
XOR2_X1 U890 ( .A(n1231), .B(KEYINPUT2), .Z(n1228) );
NAND2_X1 U891 ( .A1(n1217), .A2(n1232), .ZN(n1231) );
INV_X1 U892 ( .A(n1230), .ZN(n1217) );
NAND3_X1 U893 ( .A1(n1082), .A2(n1067), .A3(n1233), .ZN(n1230) );
XNOR2_X1 U894 ( .A(G143), .B(n1234), .ZN(G45) );
NAND4_X1 U895 ( .A1(n1235), .A2(n1236), .A3(n1067), .A4(n1078), .ZN(n1234) );
XNOR2_X1 U896 ( .A(G140), .B(n1237), .ZN(G42) );
NAND4_X1 U897 ( .A1(n1238), .A2(n1236), .A3(n1082), .A4(n1239), .ZN(n1237) );
XNOR2_X1 U898 ( .A(n1073), .B(KEYINPUT56), .ZN(n1238) );
NAND2_X1 U899 ( .A1(n1240), .A2(n1241), .ZN(G39) );
NAND2_X1 U900 ( .A1(G137), .A2(n1218), .ZN(n1241) );
XOR2_X1 U901 ( .A(n1242), .B(KEYINPUT60), .Z(n1240) );
OR2_X1 U902 ( .A1(n1218), .A2(G137), .ZN(n1242) );
NAND3_X1 U903 ( .A1(n1233), .A2(n1073), .A3(n1052), .ZN(n1218) );
XNOR2_X1 U904 ( .A(G134), .B(n1243), .ZN(G36) );
NAND3_X1 U905 ( .A1(n1244), .A2(n1073), .A3(n1245), .ZN(n1243) );
NOR3_X1 U906 ( .A1(n1203), .A2(n1246), .A3(n1087), .ZN(n1245) );
XNOR2_X1 U907 ( .A(n1059), .B(KEYINPUT27), .ZN(n1244) );
XNOR2_X1 U908 ( .A(G131), .B(n1213), .ZN(G33) );
NAND4_X1 U909 ( .A1(n1236), .A2(n1082), .A3(n1073), .A4(n1078), .ZN(n1213) );
NOR2_X1 U910 ( .A1(n1069), .A2(n1247), .ZN(n1073) );
INV_X1 U911 ( .A(n1068), .ZN(n1247) );
XNOR2_X1 U912 ( .A(G128), .B(n1211), .ZN(G30) );
NAND3_X1 U913 ( .A1(n1067), .A2(n1083), .A3(n1233), .ZN(n1211) );
NOR3_X1 U914 ( .A1(n1248), .A2(n1249), .A3(n1220), .ZN(n1233) );
INV_X1 U915 ( .A(n1236), .ZN(n1220) );
NOR2_X1 U916 ( .A1(n1250), .A2(n1246), .ZN(n1236) );
XNOR2_X1 U917 ( .A(G101), .B(n1206), .ZN(G3) );
NAND4_X1 U918 ( .A1(n1052), .A2(n1067), .A3(n1210), .A4(n1078), .ZN(n1206) );
XNOR2_X1 U919 ( .A(n1251), .B(n1252), .ZN(G27) );
NAND2_X1 U920 ( .A1(KEYINPUT38), .A2(n1212), .ZN(n1251) );
NAND4_X1 U921 ( .A1(n1082), .A2(n1061), .A3(n1253), .A4(n1239), .ZN(n1212) );
NOR2_X1 U922 ( .A1(n1246), .A2(n1162), .ZN(n1253) );
AND2_X1 U923 ( .A1(n1254), .A2(n1077), .ZN(n1246) );
NAND4_X1 U924 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1256), .ZN(n1254) );
INV_X1 U925 ( .A(G900), .ZN(n1256) );
XNOR2_X1 U926 ( .A(G122), .B(n1257), .ZN(G24) );
NAND3_X1 U927 ( .A1(n1235), .A2(n1051), .A3(n1258), .ZN(n1257) );
NAND2_X1 U928 ( .A1(n1259), .A2(n1260), .ZN(n1051) );
OR3_X1 U929 ( .A1(n1261), .A2(n1100), .A3(KEYINPUT8), .ZN(n1260) );
NAND2_X1 U930 ( .A1(KEYINPUT8), .A2(n1078), .ZN(n1259) );
INV_X1 U931 ( .A(n1204), .ZN(n1235) );
NAND2_X1 U932 ( .A1(n1262), .A2(n1263), .ZN(n1204) );
XNOR2_X1 U933 ( .A(G119), .B(n1193), .ZN(G21) );
NAND4_X1 U934 ( .A1(n1258), .A2(n1052), .A3(n1261), .A4(n1100), .ZN(n1193) );
INV_X1 U935 ( .A(n1199), .ZN(n1258) );
XOR2_X1 U936 ( .A(n1264), .B(n1265), .Z(G18) );
NAND2_X1 U937 ( .A1(n1266), .A2(n1083), .ZN(n1265) );
INV_X1 U938 ( .A(n1203), .ZN(n1083) );
NAND2_X1 U939 ( .A1(n1263), .A2(n1267), .ZN(n1203) );
NAND2_X1 U940 ( .A1(KEYINPUT51), .A2(G116), .ZN(n1264) );
XNOR2_X1 U941 ( .A(n1268), .B(n1192), .ZN(G15) );
NAND2_X1 U942 ( .A1(n1266), .A2(n1082), .ZN(n1192) );
NOR2_X1 U943 ( .A1(n1267), .A2(n1263), .ZN(n1082) );
NOR2_X1 U944 ( .A1(n1199), .A2(n1087), .ZN(n1266) );
INV_X1 U945 ( .A(n1078), .ZN(n1087) );
NOR2_X1 U946 ( .A1(n1261), .A2(n1249), .ZN(n1078) );
INV_X1 U947 ( .A(n1100), .ZN(n1249) );
NAND3_X1 U948 ( .A1(n1067), .A2(n1269), .A3(n1061), .ZN(n1199) );
NOR2_X1 U949 ( .A1(n1062), .A2(n1092), .ZN(n1061) );
INV_X1 U950 ( .A(n1063), .ZN(n1092) );
XNOR2_X1 U951 ( .A(G113), .B(KEYINPUT17), .ZN(n1268) );
XNOR2_X1 U952 ( .A(G110), .B(n1270), .ZN(G12) );
NAND2_X1 U953 ( .A1(n1271), .A2(n1067), .ZN(n1270) );
INV_X1 U954 ( .A(n1162), .ZN(n1067) );
NAND2_X1 U955 ( .A1(n1069), .A2(n1068), .ZN(n1162) );
NAND2_X1 U956 ( .A1(G214), .A2(n1272), .ZN(n1068) );
NAND2_X1 U957 ( .A1(n1273), .A2(n1146), .ZN(n1272) );
NAND2_X1 U958 ( .A1(n1274), .A2(n1275), .ZN(n1069) );
NAND2_X1 U959 ( .A1(G210), .A2(n1276), .ZN(n1275) );
NAND2_X1 U960 ( .A1(n1146), .A2(n1277), .ZN(n1276) );
OR2_X1 U961 ( .A1(n1273), .A2(n1278), .ZN(n1277) );
INV_X1 U962 ( .A(G237), .ZN(n1273) );
NAND3_X1 U963 ( .A1(n1279), .A2(n1146), .A3(n1278), .ZN(n1274) );
XNOR2_X1 U964 ( .A(n1187), .B(KEYINPUT21), .ZN(n1278) );
XOR2_X1 U965 ( .A(n1280), .B(n1281), .Z(n1187) );
XNOR2_X1 U966 ( .A(n1252), .B(n1282), .ZN(n1281) );
NOR2_X1 U967 ( .A1(G953), .A2(n1121), .ZN(n1282) );
INV_X1 U968 ( .A(G224), .ZN(n1121) );
INV_X1 U969 ( .A(G125), .ZN(n1252) );
XNOR2_X1 U970 ( .A(n1283), .B(n1284), .ZN(n1280) );
NAND2_X1 U971 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
NAND2_X1 U972 ( .A1(n1128), .A2(n1287), .ZN(n1286) );
NAND2_X1 U973 ( .A1(n1130), .A2(n1131), .ZN(n1287) );
NAND2_X1 U974 ( .A1(n1288), .A2(n1289), .ZN(n1131) );
OR2_X1 U975 ( .A1(n1289), .A2(n1288), .ZN(n1130) );
INV_X1 U976 ( .A(n1290), .ZN(n1128) );
NAND2_X1 U977 ( .A1(n1291), .A2(n1290), .ZN(n1285) );
XOR2_X1 U978 ( .A(G110), .B(n1292), .Z(n1290) );
XOR2_X1 U979 ( .A(KEYINPUT7), .B(G122), .Z(n1292) );
XOR2_X1 U980 ( .A(n1289), .B(n1288), .Z(n1291) );
NAND2_X1 U981 ( .A1(n1293), .A2(n1294), .ZN(n1288) );
NAND2_X1 U982 ( .A1(G107), .A2(n1295), .ZN(n1294) );
NAND2_X1 U983 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
XOR2_X1 U984 ( .A(n1295), .B(KEYINPUT42), .Z(n1296) );
XNOR2_X1 U985 ( .A(G101), .B(n1298), .ZN(n1295) );
XNOR2_X1 U986 ( .A(KEYINPUT18), .B(n1159), .ZN(n1298) );
NAND3_X1 U987 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1289) );
NAND2_X1 U988 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U989 ( .A1(n1304), .A2(n1305), .ZN(n1300) );
INV_X1 U990 ( .A(KEYINPUT52), .ZN(n1305) );
NAND2_X1 U991 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
XNOR2_X1 U992 ( .A(KEYINPUT13), .B(n1303), .ZN(n1306) );
NAND2_X1 U993 ( .A1(KEYINPUT52), .A2(n1308), .ZN(n1299) );
NAND2_X1 U994 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
OR3_X1 U995 ( .A1(n1303), .A2(n1302), .A3(KEYINPUT13), .ZN(n1310) );
INV_X1 U996 ( .A(n1307), .ZN(n1302) );
XOR2_X1 U997 ( .A(G116), .B(G119), .Z(n1307) );
NAND2_X1 U998 ( .A1(KEYINPUT13), .A2(n1303), .ZN(n1309) );
NAND2_X1 U999 ( .A1(G210), .A2(G237), .ZN(n1279) );
XNOR2_X1 U1000 ( .A(n1208), .B(KEYINPUT40), .ZN(n1271) );
AND3_X1 U1001 ( .A1(n1239), .A2(n1210), .A3(n1052), .ZN(n1208) );
NOR2_X1 U1002 ( .A1(n1263), .A2(n1262), .ZN(n1052) );
INV_X1 U1003 ( .A(n1267), .ZN(n1262) );
XOR2_X1 U1004 ( .A(n1095), .B(KEYINPUT23), .Z(n1267) );
XOR2_X1 U1005 ( .A(n1311), .B(n1153), .Z(n1095) );
INV_X1 U1006 ( .A(G475), .ZN(n1153) );
OR2_X1 U1007 ( .A1(n1155), .A2(G902), .ZN(n1311) );
XOR2_X1 U1008 ( .A(n1312), .B(n1313), .Z(n1155) );
XOR2_X1 U1009 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1010 ( .A(G143), .B(G131), .Z(n1315) );
XOR2_X1 U1011 ( .A(KEYINPUT59), .B(KEYINPUT58), .Z(n1314) );
XOR2_X1 U1012 ( .A(n1316), .B(n1317), .Z(n1312) );
XOR2_X1 U1013 ( .A(n1318), .B(n1319), .Z(n1317) );
NAND2_X1 U1014 ( .A1(n1320), .A2(G214), .ZN(n1319) );
NAND2_X1 U1015 ( .A1(KEYINPUT55), .A2(n1321), .ZN(n1318) );
XNOR2_X1 U1016 ( .A(n1159), .B(n1322), .ZN(n1321) );
XNOR2_X1 U1017 ( .A(G122), .B(n1303), .ZN(n1322) );
INV_X1 U1018 ( .A(G113), .ZN(n1303) );
XNOR2_X1 U1019 ( .A(n1112), .B(n1323), .ZN(n1316) );
XNOR2_X1 U1020 ( .A(G125), .B(n1184), .ZN(n1112) );
XOR2_X1 U1021 ( .A(n1099), .B(n1324), .Z(n1263) );
XOR2_X1 U1022 ( .A(KEYINPUT35), .B(G478), .Z(n1324) );
AND2_X1 U1023 ( .A1(n1145), .A2(n1146), .ZN(n1099) );
NAND2_X1 U1024 ( .A1(n1325), .A2(n1326), .ZN(n1145) );
NAND3_X1 U1025 ( .A1(n1327), .A2(n1328), .A3(G217), .ZN(n1326) );
NAND2_X1 U1026 ( .A1(n1329), .A2(n1330), .ZN(n1325) );
NAND2_X1 U1027 ( .A1(G217), .A2(n1328), .ZN(n1330) );
XNOR2_X1 U1028 ( .A(KEYINPUT29), .B(n1327), .ZN(n1329) );
XOR2_X1 U1029 ( .A(n1331), .B(n1332), .Z(n1327) );
XOR2_X1 U1030 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1031 ( .A(n1335), .B(G107), .ZN(n1334) );
NOR2_X1 U1032 ( .A1(G143), .A2(KEYINPUT43), .ZN(n1333) );
XOR2_X1 U1033 ( .A(n1336), .B(n1337), .Z(n1331) );
XNOR2_X1 U1034 ( .A(n1338), .B(G122), .ZN(n1337) );
XNOR2_X1 U1035 ( .A(G134), .B(KEYINPUT31), .ZN(n1336) );
AND2_X1 U1036 ( .A1(n1059), .A2(n1269), .ZN(n1210) );
NAND2_X1 U1037 ( .A1(n1077), .A2(n1339), .ZN(n1269) );
NAND4_X1 U1038 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1132), .ZN(n1339) );
INV_X1 U1039 ( .A(G898), .ZN(n1132) );
NAND3_X1 U1040 ( .A1(n1255), .A2(n1071), .A3(G952), .ZN(n1077) );
NAND2_X1 U1041 ( .A1(G234), .A2(G237), .ZN(n1255) );
INV_X1 U1042 ( .A(n1250), .ZN(n1059) );
NAND2_X1 U1043 ( .A1(n1062), .A2(n1063), .ZN(n1250) );
NAND2_X1 U1044 ( .A1(G221), .A2(n1340), .ZN(n1063) );
XNOR2_X1 U1045 ( .A(n1341), .B(n1102), .ZN(n1062) );
NAND2_X1 U1046 ( .A1(n1342), .A2(n1146), .ZN(n1102) );
XOR2_X1 U1047 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1048 ( .A(KEYINPUT63), .B(n1181), .Z(n1344) );
AND2_X1 U1049 ( .A1(G227), .A2(n1071), .ZN(n1181) );
XNOR2_X1 U1050 ( .A(n1174), .B(n1345), .ZN(n1343) );
XNOR2_X1 U1051 ( .A(n1346), .B(n1347), .ZN(n1174) );
XNOR2_X1 U1052 ( .A(n1348), .B(n1349), .ZN(n1347) );
XNOR2_X1 U1053 ( .A(KEYINPUT10), .B(n1297), .ZN(n1349) );
INV_X1 U1054 ( .A(G107), .ZN(n1297) );
XOR2_X1 U1055 ( .A(n1111), .B(n1350), .Z(n1346) );
NOR2_X1 U1056 ( .A1(KEYINPUT46), .A2(n1159), .ZN(n1350) );
INV_X1 U1057 ( .A(G104), .ZN(n1159) );
XOR2_X1 U1058 ( .A(n1351), .B(n1352), .Z(n1111) );
XNOR2_X1 U1059 ( .A(n1353), .B(G146), .ZN(n1351) );
NAND2_X1 U1060 ( .A1(KEYINPUT26), .A2(n1103), .ZN(n1341) );
XNOR2_X1 U1061 ( .A(G469), .B(KEYINPUT3), .ZN(n1103) );
INV_X1 U1062 ( .A(n1085), .ZN(n1239) );
NAND2_X1 U1063 ( .A1(n1354), .A2(n1261), .ZN(n1085) );
INV_X1 U1064 ( .A(n1248), .ZN(n1261) );
XOR2_X1 U1065 ( .A(n1101), .B(KEYINPUT24), .Z(n1248) );
XNOR2_X1 U1066 ( .A(n1355), .B(n1141), .ZN(n1101) );
AND2_X1 U1067 ( .A1(G217), .A2(n1340), .ZN(n1141) );
NAND2_X1 U1068 ( .A1(G234), .A2(n1146), .ZN(n1340) );
NAND2_X1 U1069 ( .A1(n1139), .A2(n1146), .ZN(n1355) );
XNOR2_X1 U1070 ( .A(n1356), .B(n1357), .ZN(n1139) );
NOR2_X1 U1071 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1072 ( .A(n1360), .B(KEYINPUT45), .Z(n1359) );
NAND3_X1 U1073 ( .A1(G221), .A2(n1328), .A3(G137), .ZN(n1360) );
NOR2_X1 U1074 ( .A1(n1361), .A2(G137), .ZN(n1358) );
AND2_X1 U1075 ( .A1(n1328), .A2(G221), .ZN(n1361) );
AND2_X1 U1076 ( .A1(G234), .A2(n1071), .ZN(n1328) );
INV_X1 U1077 ( .A(G953), .ZN(n1071) );
NAND2_X1 U1078 ( .A1(KEYINPUT11), .A2(n1362), .ZN(n1356) );
XOR2_X1 U1079 ( .A(n1363), .B(n1364), .Z(n1362) );
XNOR2_X1 U1080 ( .A(n1345), .B(n1323), .ZN(n1364) );
XNOR2_X1 U1081 ( .A(n1232), .B(KEYINPUT48), .ZN(n1323) );
XNOR2_X1 U1082 ( .A(G110), .B(n1184), .ZN(n1345) );
INV_X1 U1083 ( .A(G140), .ZN(n1184) );
XOR2_X1 U1084 ( .A(n1365), .B(n1366), .Z(n1363) );
NOR2_X1 U1085 ( .A1(G125), .A2(KEYINPUT44), .ZN(n1366) );
XOR2_X1 U1086 ( .A(n1367), .B(KEYINPUT41), .Z(n1365) );
NAND2_X1 U1087 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
NAND2_X1 U1088 ( .A1(G119), .A2(n1338), .ZN(n1369) );
XOR2_X1 U1089 ( .A(KEYINPUT15), .B(n1370), .Z(n1368) );
NOR2_X1 U1090 ( .A1(G119), .A2(n1338), .ZN(n1370) );
XNOR2_X1 U1091 ( .A(n1100), .B(KEYINPUT8), .ZN(n1354) );
XNOR2_X1 U1092 ( .A(n1371), .B(G472), .ZN(n1100) );
NAND2_X1 U1093 ( .A1(n1372), .A2(n1146), .ZN(n1371) );
INV_X1 U1094 ( .A(G902), .ZN(n1146) );
XNOR2_X1 U1095 ( .A(n1165), .B(n1373), .ZN(n1372) );
NOR2_X1 U1096 ( .A1(KEYINPUT19), .A2(n1168), .ZN(n1373) );
XOR2_X1 U1097 ( .A(n1374), .B(n1375), .Z(n1168) );
XOR2_X1 U1098 ( .A(n1376), .B(n1377), .Z(n1375) );
XNOR2_X1 U1099 ( .A(G119), .B(G113), .ZN(n1377) );
NAND2_X1 U1100 ( .A1(KEYINPUT39), .A2(n1335), .ZN(n1376) );
INV_X1 U1101 ( .A(G116), .ZN(n1335) );
XOR2_X1 U1102 ( .A(n1284), .B(n1353), .Z(n1374) );
XOR2_X1 U1103 ( .A(G131), .B(n1378), .Z(n1353) );
XOR2_X1 U1104 ( .A(G137), .B(G134), .Z(n1378) );
NAND2_X1 U1105 ( .A1(n1379), .A2(n1380), .ZN(n1284) );
NAND2_X1 U1106 ( .A1(n1381), .A2(n1232), .ZN(n1380) );
INV_X1 U1107 ( .A(G146), .ZN(n1232) );
XOR2_X1 U1108 ( .A(KEYINPUT12), .B(n1352), .Z(n1381) );
NAND2_X1 U1109 ( .A1(n1352), .A2(G146), .ZN(n1379) );
XNOR2_X1 U1110 ( .A(n1338), .B(G143), .ZN(n1352) );
INV_X1 U1111 ( .A(G128), .ZN(n1338) );
XOR2_X1 U1112 ( .A(n1382), .B(n1348), .Z(n1165) );
INV_X1 U1113 ( .A(G101), .ZN(n1348) );
NAND2_X1 U1114 ( .A1(n1320), .A2(G210), .ZN(n1382) );
NOR2_X1 U1115 ( .A1(G953), .A2(G237), .ZN(n1320) );
endmodule


