//Key = 0111100010100111110001111000000101000010110100010010111000000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367;

XNOR2_X1 U749 ( .A(G107), .B(n1045), .ZN(G9) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(G75) );
XOR2_X1 U751 ( .A(n1048), .B(KEYINPUT54), .Z(n1047) );
NAND4_X1 U752 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
NAND3_X1 U753 ( .A1(n1053), .A2(n1054), .A3(KEYINPUT39), .ZN(n1052) );
NAND4_X1 U754 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NAND2_X1 U755 ( .A1(n1055), .A2(n1059), .ZN(n1051) );
NAND2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U757 ( .A1(n1062), .A2(n1063), .A3(n1058), .ZN(n1061) );
NAND2_X1 U758 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND3_X1 U759 ( .A1(n1057), .A2(n1066), .A3(KEYINPUT9), .ZN(n1064) );
NAND3_X1 U760 ( .A1(n1067), .A2(n1068), .A3(n1053), .ZN(n1062) );
NAND2_X1 U761 ( .A1(n1057), .A2(n1069), .ZN(n1068) );
NAND2_X1 U762 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1072), .ZN(n1071) );
INV_X1 U764 ( .A(KEYINPUT9), .ZN(n1072) );
OR2_X1 U765 ( .A1(n1073), .A2(KEYINPUT39), .ZN(n1070) );
NAND2_X1 U766 ( .A1(n1074), .A2(n1075), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U768 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
INV_X1 U769 ( .A(n1080), .ZN(n1076) );
NAND3_X1 U770 ( .A1(n1074), .A2(n1081), .A3(n1057), .ZN(n1060) );
NAND2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1053), .A2(n1084), .ZN(n1083) );
NAND2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U775 ( .A1(n1058), .A2(n1089), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U777 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
INV_X1 U778 ( .A(n1094), .ZN(n1090) );
INV_X1 U779 ( .A(n1095), .ZN(n1055) );
INV_X1 U780 ( .A(n1096), .ZN(n1050) );
NOR2_X1 U781 ( .A1(G952), .A2(n1096), .ZN(n1046) );
NAND2_X1 U782 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND4_X1 U783 ( .A1(n1099), .A2(n1074), .A3(n1100), .A4(n1101), .ZN(n1098) );
NOR4_X1 U784 ( .A1(n1092), .A2(n1078), .A3(n1102), .A4(n1103), .ZN(n1101) );
XOR2_X1 U785 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U786 ( .A1(n1106), .A2(KEYINPUT46), .ZN(n1105) );
XNOR2_X1 U787 ( .A(n1107), .B(n1108), .ZN(n1102) );
NAND2_X1 U788 ( .A1(KEYINPUT40), .A2(n1109), .ZN(n1107) );
NOR2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U791 ( .A(n1114), .B(KEYINPUT53), .Z(n1113) );
NOR2_X1 U792 ( .A1(n1115), .A2(n1116), .ZN(n1110) );
XOR2_X1 U793 ( .A(KEYINPUT24), .B(n1117), .Z(n1116) );
XOR2_X1 U794 ( .A(n1118), .B(n1119), .Z(n1099) );
XOR2_X1 U795 ( .A(n1120), .B(n1121), .Z(G72) );
NOR2_X1 U796 ( .A1(n1122), .A2(n1097), .ZN(n1121) );
AND2_X1 U797 ( .A1(G227), .A2(G900), .ZN(n1122) );
NOR2_X1 U798 ( .A1(KEYINPUT18), .A2(n1123), .ZN(n1120) );
XOR2_X1 U799 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U800 ( .A1(n1126), .A2(G953), .ZN(n1125) );
AND3_X1 U801 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
NAND2_X1 U802 ( .A1(n1130), .A2(n1131), .ZN(n1124) );
INV_X1 U803 ( .A(n1132), .ZN(n1131) );
XOR2_X1 U804 ( .A(n1133), .B(n1134), .Z(n1130) );
XOR2_X1 U805 ( .A(G125), .B(n1135), .Z(n1134) );
XOR2_X1 U806 ( .A(KEYINPUT26), .B(G131), .Z(n1135) );
XOR2_X1 U807 ( .A(n1136), .B(n1137), .Z(n1133) );
XOR2_X1 U808 ( .A(n1138), .B(n1139), .Z(n1136) );
NOR2_X1 U809 ( .A1(G137), .A2(KEYINPUT35), .ZN(n1139) );
XOR2_X1 U810 ( .A(n1140), .B(n1141), .Z(G69) );
XOR2_X1 U811 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U812 ( .A1(G953), .A2(n1144), .ZN(n1143) );
NAND2_X1 U813 ( .A1(G898), .A2(G224), .ZN(n1144) );
NAND4_X1 U814 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1142) );
NAND2_X1 U815 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
INV_X1 U816 ( .A(KEYINPUT62), .ZN(n1150) );
NAND2_X1 U817 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
NAND2_X1 U818 ( .A1(n1153), .A2(KEYINPUT62), .ZN(n1147) );
XOR2_X1 U819 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U820 ( .A1(G953), .A2(n1156), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1157), .A2(G953), .ZN(n1140) );
NOR2_X1 U822 ( .A1(n1158), .A2(n1159), .ZN(G66) );
XNOR2_X1 U823 ( .A(n1160), .B(n1161), .ZN(n1159) );
NOR2_X1 U824 ( .A1(n1118), .A2(n1162), .ZN(n1161) );
NOR3_X1 U825 ( .A1(n1158), .A2(n1163), .A3(n1164), .ZN(G63) );
AND4_X1 U826 ( .A1(n1165), .A2(KEYINPUT22), .A3(G478), .A4(n1166), .ZN(n1164) );
NOR2_X1 U827 ( .A1(n1165), .A2(n1167), .ZN(n1163) );
NOR3_X1 U828 ( .A1(n1162), .A2(n1168), .A3(n1169), .ZN(n1167) );
NOR2_X1 U829 ( .A1(KEYINPUT22), .A2(n1170), .ZN(n1168) );
NOR2_X1 U830 ( .A1(n1171), .A2(KEYINPUT20), .ZN(n1165) );
NOR2_X1 U831 ( .A1(n1158), .A2(n1172), .ZN(G60) );
XOR2_X1 U832 ( .A(n1173), .B(n1174), .Z(n1172) );
AND2_X1 U833 ( .A1(G475), .A2(n1166), .ZN(n1173) );
XOR2_X1 U834 ( .A(G104), .B(n1175), .Z(G6) );
NOR2_X1 U835 ( .A1(n1158), .A2(n1176), .ZN(G57) );
XOR2_X1 U836 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U837 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U838 ( .A(n1181), .B(n1182), .Z(n1177) );
XOR2_X1 U839 ( .A(KEYINPUT41), .B(G101), .Z(n1182) );
NOR2_X1 U840 ( .A1(n1104), .A2(n1162), .ZN(n1181) );
INV_X1 U841 ( .A(G472), .ZN(n1104) );
NOR2_X1 U842 ( .A1(n1158), .A2(n1183), .ZN(G54) );
NOR2_X1 U843 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U844 ( .A(n1186), .B(KEYINPUT43), .Z(n1185) );
NAND2_X1 U845 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NOR2_X1 U846 ( .A1(n1187), .A2(n1188), .ZN(n1184) );
XOR2_X1 U847 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U848 ( .A1(KEYINPUT0), .A2(n1191), .ZN(n1190) );
NOR2_X1 U849 ( .A1(n1162), .A2(n1109), .ZN(n1187) );
INV_X1 U850 ( .A(G469), .ZN(n1109) );
INV_X1 U851 ( .A(n1166), .ZN(n1162) );
NOR2_X1 U852 ( .A1(n1158), .A2(n1192), .ZN(G51) );
XOR2_X1 U853 ( .A(n1193), .B(n1194), .Z(n1192) );
NAND3_X1 U854 ( .A1(n1166), .A2(n1117), .A3(KEYINPUT3), .ZN(n1194) );
INV_X1 U855 ( .A(n1114), .ZN(n1117) );
NOR2_X1 U856 ( .A1(n1195), .A2(n1049), .ZN(n1166) );
AND4_X1 U857 ( .A1(n1157), .A2(n1127), .A3(n1196), .A4(n1128), .ZN(n1049) );
XNOR2_X1 U858 ( .A(KEYINPUT38), .B(n1129), .ZN(n1196) );
AND4_X1 U859 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1127) );
AND3_X1 U860 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
AND4_X1 U861 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1157) );
AND4_X1 U862 ( .A1(n1045), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1207) );
NAND3_X1 U863 ( .A1(n1066), .A2(n1058), .A3(n1211), .ZN(n1045) );
NOR2_X1 U864 ( .A1(n1175), .A2(n1212), .ZN(n1206) );
NOR2_X1 U865 ( .A1(n1213), .A2(n1085), .ZN(n1212) );
INV_X1 U866 ( .A(n1214), .ZN(n1085) );
AND3_X1 U867 ( .A1(n1211), .A2(n1058), .A3(n1056), .ZN(n1175) );
NAND2_X1 U868 ( .A1(n1215), .A2(n1216), .ZN(n1193) );
NAND2_X1 U869 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U870 ( .A(n1219), .B(KEYINPUT42), .Z(n1215) );
OR2_X1 U871 ( .A1(n1218), .A2(n1217), .ZN(n1219) );
NAND2_X1 U872 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
NAND2_X1 U873 ( .A1(KEYINPUT28), .A2(n1222), .ZN(n1221) );
XOR2_X1 U874 ( .A(n1223), .B(n1224), .Z(n1220) );
OR2_X1 U875 ( .A1(n1222), .A2(KEYINPUT28), .ZN(n1223) );
XNOR2_X1 U876 ( .A(n1225), .B(G125), .ZN(n1222) );
AND2_X1 U877 ( .A1(G953), .A2(n1226), .ZN(n1158) );
XOR2_X1 U878 ( .A(KEYINPUT8), .B(G952), .Z(n1226) );
XOR2_X1 U879 ( .A(G146), .B(n1227), .Z(G48) );
NOR2_X1 U880 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
AND2_X1 U881 ( .A1(KEYINPUT31), .A2(n1199), .ZN(n1229) );
NOR2_X1 U882 ( .A1(KEYINPUT13), .A2(n1199), .ZN(n1228) );
NAND2_X1 U883 ( .A1(n1230), .A2(n1056), .ZN(n1199) );
XNOR2_X1 U884 ( .A(G143), .B(n1129), .ZN(G45) );
NAND4_X1 U885 ( .A1(n1231), .A2(n1094), .A3(n1232), .A4(n1233), .ZN(n1129) );
XOR2_X1 U886 ( .A(n1234), .B(G140), .Z(G42) );
NAND2_X1 U887 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
OR2_X1 U888 ( .A1(n1128), .A2(KEYINPUT5), .ZN(n1236) );
NAND2_X1 U889 ( .A1(n1237), .A2(n1053), .ZN(n1128) );
NAND3_X1 U890 ( .A1(n1237), .A2(n1065), .A3(KEYINPUT5), .ZN(n1235) );
AND3_X1 U891 ( .A1(n1087), .A2(n1056), .A3(n1238), .ZN(n1237) );
XNOR2_X1 U892 ( .A(G137), .B(n1197), .ZN(G39) );
NAND4_X1 U893 ( .A1(n1053), .A2(n1238), .A3(n1074), .A4(n1239), .ZN(n1197) );
XNOR2_X1 U894 ( .A(G134), .B(n1198), .ZN(G36) );
NAND3_X1 U895 ( .A1(n1053), .A2(n1066), .A3(n1231), .ZN(n1198) );
XOR2_X1 U896 ( .A(G131), .B(n1240), .Z(G33) );
NOR2_X1 U897 ( .A1(KEYINPUT25), .A2(n1201), .ZN(n1240) );
NAND3_X1 U898 ( .A1(n1053), .A2(n1056), .A3(n1231), .ZN(n1201) );
AND3_X1 U899 ( .A1(n1080), .A2(n1241), .A3(n1214), .ZN(n1231) );
INV_X1 U900 ( .A(n1065), .ZN(n1053) );
NAND2_X1 U901 ( .A1(n1093), .A2(n1242), .ZN(n1065) );
XNOR2_X1 U902 ( .A(n1243), .B(KEYINPUT52), .ZN(n1093) );
XOR2_X1 U903 ( .A(n1244), .B(n1203), .Z(G30) );
NAND2_X1 U904 ( .A1(n1230), .A2(n1066), .ZN(n1203) );
AND3_X1 U905 ( .A1(n1094), .A2(n1239), .A3(n1238), .ZN(n1230) );
AND3_X1 U906 ( .A1(n1088), .A2(n1241), .A3(n1080), .ZN(n1238) );
NAND2_X1 U907 ( .A1(n1245), .A2(n1246), .ZN(G3) );
NAND3_X1 U908 ( .A1(KEYINPUT21), .A2(n1247), .A3(n1248), .ZN(n1246) );
NAND2_X1 U909 ( .A1(n1249), .A2(G101), .ZN(n1245) );
NAND2_X1 U910 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND2_X1 U911 ( .A1(n1247), .A2(n1252), .ZN(n1251) );
INV_X1 U912 ( .A(KEYINPUT2), .ZN(n1252) );
NAND2_X1 U913 ( .A1(KEYINPUT2), .A2(n1253), .ZN(n1250) );
NAND2_X1 U914 ( .A1(KEYINPUT21), .A2(n1247), .ZN(n1253) );
AND2_X1 U915 ( .A1(n1254), .A2(n1255), .ZN(n1247) );
XOR2_X1 U916 ( .A(KEYINPUT7), .B(n1214), .Z(n1255) );
XOR2_X1 U917 ( .A(n1256), .B(n1202), .Z(G27) );
NAND4_X1 U918 ( .A1(n1088), .A2(n1241), .A3(n1094), .A4(n1257), .ZN(n1202) );
NOR3_X1 U919 ( .A1(n1073), .A2(n1258), .A3(n1239), .ZN(n1257) );
NAND2_X1 U920 ( .A1(n1095), .A2(n1259), .ZN(n1241) );
NAND3_X1 U921 ( .A1(G902), .A2(n1260), .A3(n1132), .ZN(n1259) );
NOR2_X1 U922 ( .A1(n1097), .A2(G900), .ZN(n1132) );
XNOR2_X1 U923 ( .A(G122), .B(n1204), .ZN(G24) );
NAND4_X1 U924 ( .A1(n1261), .A2(n1058), .A3(n1232), .A4(n1233), .ZN(n1204) );
NOR2_X1 U925 ( .A1(n1239), .A2(n1262), .ZN(n1058) );
XOR2_X1 U926 ( .A(n1263), .B(n1205), .Z(G21) );
NAND4_X1 U927 ( .A1(n1261), .A2(n1074), .A3(n1088), .A4(n1239), .ZN(n1205) );
XNOR2_X1 U928 ( .A(G116), .B(n1210), .ZN(G18) );
NAND3_X1 U929 ( .A1(n1214), .A2(n1066), .A3(n1261), .ZN(n1210) );
NOR2_X1 U930 ( .A1(n1232), .A2(n1264), .ZN(n1066) );
NAND2_X1 U931 ( .A1(n1265), .A2(n1266), .ZN(G15) );
NAND2_X1 U932 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XOR2_X1 U933 ( .A(n1209), .B(KEYINPUT16), .Z(n1267) );
NAND2_X1 U934 ( .A1(n1269), .A2(G113), .ZN(n1265) );
XNOR2_X1 U935 ( .A(KEYINPUT17), .B(n1209), .ZN(n1269) );
NAND3_X1 U936 ( .A1(n1214), .A2(n1056), .A3(n1261), .ZN(n1209) );
AND3_X1 U937 ( .A1(n1094), .A2(n1270), .A3(n1057), .ZN(n1261) );
INV_X1 U938 ( .A(n1258), .ZN(n1057) );
NAND2_X1 U939 ( .A1(n1079), .A2(n1271), .ZN(n1258) );
INV_X1 U940 ( .A(n1073), .ZN(n1056) );
NAND2_X1 U941 ( .A1(n1264), .A2(n1232), .ZN(n1073) );
NOR2_X1 U942 ( .A1(n1087), .A2(n1262), .ZN(n1214) );
XNOR2_X1 U943 ( .A(G110), .B(n1208), .ZN(G12) );
NAND3_X1 U944 ( .A1(n1087), .A2(n1088), .A3(n1254), .ZN(n1208) );
INV_X1 U945 ( .A(n1213), .ZN(n1254) );
NAND2_X1 U946 ( .A1(n1074), .A2(n1211), .ZN(n1213) );
AND3_X1 U947 ( .A1(n1080), .A2(n1270), .A3(n1094), .ZN(n1211) );
NOR2_X1 U948 ( .A1(n1243), .A2(n1092), .ZN(n1094) );
INV_X1 U949 ( .A(n1242), .ZN(n1092) );
NAND2_X1 U950 ( .A1(G214), .A2(n1272), .ZN(n1242) );
XOR2_X1 U951 ( .A(n1115), .B(n1114), .Z(n1243) );
NAND2_X1 U952 ( .A1(G210), .A2(n1272), .ZN(n1114) );
NAND2_X1 U953 ( .A1(n1273), .A2(n1195), .ZN(n1272) );
INV_X1 U954 ( .A(G237), .ZN(n1273) );
INV_X1 U955 ( .A(n1112), .ZN(n1115) );
NAND2_X1 U956 ( .A1(n1274), .A2(n1195), .ZN(n1112) );
XOR2_X1 U957 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U958 ( .A(KEYINPUT59), .B(n1224), .Z(n1276) );
AND2_X1 U959 ( .A1(G224), .A2(n1097), .ZN(n1224) );
XOR2_X1 U960 ( .A(n1277), .B(n1278), .Z(n1275) );
NOR2_X1 U961 ( .A1(n1217), .A2(KEYINPUT48), .ZN(n1278) );
AND3_X1 U962 ( .A1(n1152), .A2(n1151), .A3(n1146), .ZN(n1217) );
NAND3_X1 U963 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1146) );
NAND3_X1 U964 ( .A1(n1282), .A2(n1154), .A3(n1155), .ZN(n1151) );
INV_X1 U965 ( .A(n1283), .ZN(n1154) );
NAND2_X1 U966 ( .A1(n1281), .A2(n1279), .ZN(n1282) );
NAND2_X1 U967 ( .A1(n1283), .A2(n1280), .ZN(n1152) );
INV_X1 U968 ( .A(n1155), .ZN(n1280) );
XNOR2_X1 U969 ( .A(G122), .B(n1284), .ZN(n1155) );
NOR2_X1 U970 ( .A1(n1279), .A2(n1281), .ZN(n1283) );
XOR2_X1 U971 ( .A(n1285), .B(n1286), .Z(n1281) );
NOR2_X1 U972 ( .A1(G104), .A2(KEYINPUT37), .ZN(n1286) );
XNOR2_X1 U973 ( .A(n1287), .B(n1288), .ZN(n1279) );
XOR2_X1 U974 ( .A(KEYINPUT60), .B(G119), .Z(n1288) );
XNOR2_X1 U975 ( .A(G116), .B(n1289), .ZN(n1287) );
NAND2_X1 U976 ( .A1(n1290), .A2(n1291), .ZN(n1277) );
NAND2_X1 U977 ( .A1(n1292), .A2(n1256), .ZN(n1291) );
XOR2_X1 U978 ( .A(n1225), .B(KEYINPUT56), .Z(n1292) );
OR2_X1 U979 ( .A1(n1256), .A2(n1225), .ZN(n1290) );
NAND2_X1 U980 ( .A1(n1095), .A2(n1293), .ZN(n1270) );
NAND4_X1 U981 ( .A1(G953), .A2(G902), .A3(n1260), .A4(n1156), .ZN(n1293) );
INV_X1 U982 ( .A(G898), .ZN(n1156) );
NAND3_X1 U983 ( .A1(n1260), .A2(n1097), .A3(G952), .ZN(n1095) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1260) );
NOR2_X1 U985 ( .A1(n1079), .A2(n1078), .ZN(n1080) );
INV_X1 U986 ( .A(n1271), .ZN(n1078) );
NAND2_X1 U987 ( .A1(n1294), .A2(n1295), .ZN(n1271) );
XNOR2_X1 U988 ( .A(G221), .B(KEYINPUT61), .ZN(n1294) );
XNOR2_X1 U989 ( .A(n1108), .B(n1296), .ZN(n1079) );
XOR2_X1 U990 ( .A(KEYINPUT4), .B(G469), .Z(n1296) );
NAND2_X1 U991 ( .A1(n1297), .A2(n1195), .ZN(n1108) );
XOR2_X1 U992 ( .A(n1191), .B(n1298), .Z(n1297) );
XOR2_X1 U993 ( .A(n1189), .B(KEYINPUT36), .Z(n1298) );
XOR2_X1 U994 ( .A(n1299), .B(n1300), .Z(n1189) );
XOR2_X1 U995 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U996 ( .A(G104), .B(KEYINPUT57), .ZN(n1302) );
XOR2_X1 U997 ( .A(n1285), .B(n1137), .Z(n1299) );
XNOR2_X1 U998 ( .A(n1303), .B(n1304), .ZN(n1137) );
XOR2_X1 U999 ( .A(G107), .B(n1248), .Z(n1285) );
XOR2_X1 U1000 ( .A(n1305), .B(n1284), .Z(n1191) );
XOR2_X1 U1001 ( .A(n1306), .B(n1307), .Z(n1305) );
INV_X1 U1002 ( .A(n1138), .ZN(n1307) );
NAND2_X1 U1003 ( .A1(G227), .A2(n1097), .ZN(n1306) );
NOR2_X1 U1004 ( .A1(n1233), .A2(n1232), .ZN(n1074) );
XNOR2_X1 U1005 ( .A(n1308), .B(G475), .ZN(n1232) );
OR2_X1 U1006 ( .A1(n1174), .A2(G902), .ZN(n1308) );
XNOR2_X1 U1007 ( .A(n1309), .B(n1310), .ZN(n1174) );
XNOR2_X1 U1008 ( .A(n1289), .B(n1311), .ZN(n1310) );
XOR2_X1 U1009 ( .A(n1312), .B(n1313), .Z(n1311) );
NOR2_X1 U1010 ( .A1(G125), .A2(KEYINPUT45), .ZN(n1313) );
XOR2_X1 U1011 ( .A(n1314), .B(n1315), .Z(n1309) );
NOR2_X1 U1012 ( .A1(G122), .A2(KEYINPUT12), .ZN(n1315) );
XOR2_X1 U1013 ( .A(n1316), .B(G104), .Z(n1314) );
NAND2_X1 U1014 ( .A1(KEYINPUT15), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1015 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1016 ( .A(G131), .B(n1320), .Z(n1319) );
AND3_X1 U1017 ( .A1(n1321), .A2(n1322), .A3(G214), .ZN(n1320) );
INV_X1 U1018 ( .A(KEYINPUT34), .ZN(n1322) );
XOR2_X1 U1019 ( .A(KEYINPUT29), .B(G143), .Z(n1318) );
INV_X1 U1020 ( .A(n1264), .ZN(n1233) );
XOR2_X1 U1021 ( .A(n1169), .B(n1323), .Z(n1264) );
NOR2_X1 U1022 ( .A1(n1171), .A2(G902), .ZN(n1323) );
INV_X1 U1023 ( .A(n1170), .ZN(n1171) );
NAND2_X1 U1024 ( .A1(n1324), .A2(n1325), .ZN(n1170) );
NAND2_X1 U1025 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1027 ( .A(KEYINPUT1), .B(n1329), .Z(n1324) );
NOR3_X1 U1028 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1329) );
INV_X1 U1029 ( .A(G217), .ZN(n1332) );
XNOR2_X1 U1030 ( .A(KEYINPUT10), .B(n1326), .ZN(n1330) );
XOR2_X1 U1031 ( .A(n1333), .B(n1334), .Z(n1326) );
XNOR2_X1 U1032 ( .A(n1335), .B(n1303), .ZN(n1334) );
XOR2_X1 U1033 ( .A(G134), .B(n1244), .Z(n1303) );
INV_X1 U1034 ( .A(G128), .ZN(n1244) );
NOR2_X1 U1035 ( .A1(G143), .A2(KEYINPUT49), .ZN(n1335) );
XNOR2_X1 U1036 ( .A(G107), .B(n1336), .ZN(n1333) );
XOR2_X1 U1037 ( .A(G122), .B(G116), .Z(n1336) );
INV_X1 U1038 ( .A(G478), .ZN(n1169) );
XNOR2_X1 U1039 ( .A(n1262), .B(KEYINPUT33), .ZN(n1088) );
XNOR2_X1 U1040 ( .A(n1119), .B(n1337), .ZN(n1262) );
NOR2_X1 U1041 ( .A1(n1338), .A2(KEYINPUT51), .ZN(n1337) );
INV_X1 U1042 ( .A(n1118), .ZN(n1338) );
NAND2_X1 U1043 ( .A1(G217), .A2(n1295), .ZN(n1118) );
NAND2_X1 U1044 ( .A1(n1339), .A2(G234), .ZN(n1295) );
XOR2_X1 U1045 ( .A(n1195), .B(KEYINPUT30), .Z(n1339) );
AND2_X1 U1046 ( .A1(n1340), .A2(n1160), .ZN(n1119) );
XNOR2_X1 U1047 ( .A(n1341), .B(n1342), .ZN(n1160) );
XOR2_X1 U1048 ( .A(G137), .B(n1343), .Z(n1342) );
NOR2_X1 U1049 ( .A1(KEYINPUT32), .A2(n1344), .ZN(n1343) );
XOR2_X1 U1050 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1051 ( .A(n1347), .B(n1348), .Z(n1346) );
XOR2_X1 U1052 ( .A(n1256), .B(KEYINPUT58), .Z(n1348) );
INV_X1 U1053 ( .A(G125), .ZN(n1256) );
NAND2_X1 U1054 ( .A1(n1349), .A2(n1350), .ZN(n1347) );
NAND2_X1 U1055 ( .A1(G128), .A2(n1263), .ZN(n1350) );
XOR2_X1 U1056 ( .A(KEYINPUT50), .B(n1351), .Z(n1349) );
NOR2_X1 U1057 ( .A1(G128), .A2(n1263), .ZN(n1351) );
INV_X1 U1058 ( .A(G119), .ZN(n1263) );
XOR2_X1 U1059 ( .A(n1312), .B(n1284), .Z(n1345) );
XOR2_X1 U1060 ( .A(G110), .B(KEYINPUT27), .Z(n1284) );
XOR2_X1 U1061 ( .A(G146), .B(n1138), .Z(n1312) );
XNOR2_X1 U1062 ( .A(G140), .B(KEYINPUT14), .ZN(n1138) );
NAND2_X1 U1063 ( .A1(n1328), .A2(G221), .ZN(n1341) );
INV_X1 U1064 ( .A(n1331), .ZN(n1328) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1097), .ZN(n1331) );
INV_X1 U1066 ( .A(G953), .ZN(n1097) );
XOR2_X1 U1067 ( .A(n1195), .B(KEYINPUT6), .Z(n1340) );
INV_X1 U1068 ( .A(n1239), .ZN(n1087) );
XOR2_X1 U1069 ( .A(n1106), .B(G472), .Z(n1239) );
AND2_X1 U1070 ( .A1(n1352), .A2(n1195), .ZN(n1106) );
INV_X1 U1071 ( .A(G902), .ZN(n1195) );
XOR2_X1 U1072 ( .A(n1353), .B(n1179), .Z(n1352) );
XNOR2_X1 U1073 ( .A(n1354), .B(n1289), .ZN(n1179) );
XNOR2_X1 U1074 ( .A(n1268), .B(KEYINPUT19), .ZN(n1289) );
INV_X1 U1075 ( .A(G113), .ZN(n1268) );
XOR2_X1 U1076 ( .A(n1355), .B(n1356), .Z(n1354) );
NOR2_X1 U1077 ( .A1(KEYINPUT11), .A2(n1357), .ZN(n1356) );
XOR2_X1 U1078 ( .A(n1358), .B(G116), .Z(n1357) );
NAND2_X1 U1079 ( .A1(KEYINPUT23), .A2(G119), .ZN(n1358) );
NAND2_X1 U1080 ( .A1(n1321), .A2(G210), .ZN(n1355) );
NOR2_X1 U1081 ( .A1(G953), .A2(G237), .ZN(n1321) );
XNOR2_X1 U1082 ( .A(n1359), .B(n1360), .ZN(n1353) );
NOR2_X1 U1083 ( .A1(KEYINPUT55), .A2(n1248), .ZN(n1360) );
INV_X1 U1084 ( .A(G101), .ZN(n1248) );
NOR2_X1 U1085 ( .A1(KEYINPUT44), .A2(n1180), .ZN(n1359) );
XNOR2_X1 U1086 ( .A(n1225), .B(n1361), .ZN(n1180) );
XNOR2_X1 U1087 ( .A(G134), .B(n1301), .ZN(n1361) );
XOR2_X1 U1088 ( .A(n1362), .B(G137), .Z(n1301) );
NAND2_X1 U1089 ( .A1(KEYINPUT47), .A2(n1363), .ZN(n1362) );
INV_X1 U1090 ( .A(G131), .ZN(n1363) );
NAND2_X1 U1091 ( .A1(n1364), .A2(n1365), .ZN(n1225) );
NAND3_X1 U1092 ( .A1(G128), .A2(n1304), .A3(n1366), .ZN(n1365) );
INV_X1 U1093 ( .A(KEYINPUT63), .ZN(n1366) );
NAND2_X1 U1094 ( .A1(n1367), .A2(KEYINPUT63), .ZN(n1364) );
XOR2_X1 U1095 ( .A(G128), .B(n1304), .Z(n1367) );
XOR2_X1 U1096 ( .A(G146), .B(G143), .Z(n1304) );
endmodule


