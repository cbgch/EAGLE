//Key = 1111011011111110011011000010111111010100100101001111111110010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400;

XNOR2_X1 U770 ( .A(G107), .B(n1066), .ZN(G9) );
NAND4_X1 U771 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
XOR2_X1 U772 ( .A(n1071), .B(KEYINPUT55), .Z(n1067) );
NOR2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(G75) );
NOR4_X1 U774 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
INV_X1 U775 ( .A(G952), .ZN(n1076) );
NAND4_X1 U776 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1074) );
NAND4_X1 U777 ( .A1(n1082), .A2(n1083), .A3(n1070), .A4(n1084), .ZN(n1079) );
NAND3_X1 U778 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND3_X1 U780 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1085) );
NAND3_X1 U781 ( .A1(n1088), .A2(n1093), .A3(n1090), .ZN(n1078) );
NAND2_X1 U782 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND3_X1 U783 ( .A1(n1083), .A2(n1096), .A3(n1097), .ZN(n1095) );
XNOR2_X1 U784 ( .A(n1082), .B(KEYINPUT35), .ZN(n1097) );
NAND2_X1 U785 ( .A1(n1082), .A2(n1098), .ZN(n1094) );
NAND3_X1 U786 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NAND2_X1 U787 ( .A1(n1070), .A2(n1102), .ZN(n1101) );
NAND3_X1 U788 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1100) );
XOR2_X1 U789 ( .A(KEYINPUT48), .B(n1106), .Z(n1104) );
XOR2_X1 U790 ( .A(KEYINPUT44), .B(n1070), .Z(n1103) );
NAND2_X1 U791 ( .A1(n1083), .A2(n1107), .ZN(n1099) );
AND2_X1 U792 ( .A1(KEYINPUT40), .A2(n1108), .ZN(n1082) );
NOR3_X1 U793 ( .A1(n1109), .A2(G953), .A3(n1110), .ZN(n1072) );
INV_X1 U794 ( .A(n1080), .ZN(n1110) );
NAND2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1080) );
NOR4_X1 U796 ( .A1(n1105), .A2(n1092), .A3(n1113), .A4(n1114), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U798 ( .A(KEYINPUT42), .B(KEYINPUT11), .Z(n1116) );
XOR2_X1 U799 ( .A(n1117), .B(n1118), .Z(n1113) );
NOR2_X1 U800 ( .A1(n1119), .A2(KEYINPUT27), .ZN(n1118) );
NOR4_X1 U801 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1111) );
XNOR2_X1 U802 ( .A(n1124), .B(n1125), .ZN(n1123) );
XOR2_X1 U803 ( .A(G478), .B(n1126), .Z(n1122) );
XOR2_X1 U804 ( .A(n1127), .B(n1128), .Z(n1121) );
XOR2_X1 U805 ( .A(n1129), .B(n1130), .Z(n1120) );
XOR2_X1 U806 ( .A(KEYINPUT16), .B(G952), .Z(n1109) );
XOR2_X1 U807 ( .A(n1131), .B(n1132), .Z(G72) );
XOR2_X1 U808 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U810 ( .A1(G953), .A2(n1137), .ZN(n1136) );
XOR2_X1 U811 ( .A(n1138), .B(n1139), .Z(n1135) );
XOR2_X1 U812 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U813 ( .A1(KEYINPUT25), .A2(n1142), .ZN(n1141) );
XOR2_X1 U814 ( .A(n1143), .B(n1144), .Z(n1138) );
NAND2_X1 U815 ( .A1(KEYINPUT59), .A2(n1145), .ZN(n1133) );
NAND2_X1 U816 ( .A1(G953), .A2(n1146), .ZN(n1145) );
NAND2_X1 U817 ( .A1(n1147), .A2(G900), .ZN(n1146) );
XNOR2_X1 U818 ( .A(G227), .B(KEYINPUT2), .ZN(n1147) );
NOR2_X1 U819 ( .A1(n1148), .A2(KEYINPUT19), .ZN(n1131) );
AND2_X1 U820 ( .A1(n1081), .A2(n1077), .ZN(n1148) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(G69) );
XOR2_X1 U822 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND3_X1 U823 ( .A1(n1153), .A2(n1154), .A3(KEYINPUT54), .ZN(n1152) );
NAND2_X1 U824 ( .A1(G953), .A2(n1155), .ZN(n1153) );
NAND2_X1 U825 ( .A1(n1156), .A2(n1154), .ZN(n1151) );
INV_X1 U826 ( .A(n1157), .ZN(n1154) );
XOR2_X1 U827 ( .A(n1158), .B(KEYINPUT4), .Z(n1156) );
NAND2_X1 U828 ( .A1(n1081), .A2(n1075), .ZN(n1149) );
NOR2_X1 U829 ( .A1(n1159), .A2(n1160), .ZN(G66) );
XNOR2_X1 U830 ( .A(n1161), .B(KEYINPUT43), .ZN(n1160) );
NOR3_X1 U831 ( .A1(n1124), .A2(n1162), .A3(n1163), .ZN(n1159) );
NOR3_X1 U832 ( .A1(n1164), .A2(n1125), .A3(n1165), .ZN(n1163) );
NOR2_X1 U833 ( .A1(n1166), .A2(n1167), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1168), .A2(n1125), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1161), .A2(n1169), .ZN(G63) );
NOR3_X1 U836 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1169) );
AND2_X1 U837 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U838 ( .A1(n1175), .A2(n1173), .ZN(n1171) );
NOR2_X1 U839 ( .A1(n1176), .A2(n1126), .ZN(n1175) );
NOR2_X1 U840 ( .A1(n1177), .A2(n1174), .ZN(n1176) );
NOR2_X1 U841 ( .A1(n1168), .A2(n1178), .ZN(n1177) );
NOR3_X1 U842 ( .A1(n1165), .A2(n1179), .A3(n1178), .ZN(n1170) );
NOR2_X1 U843 ( .A1(n1174), .A2(n1173), .ZN(n1179) );
INV_X1 U844 ( .A(KEYINPUT5), .ZN(n1173) );
NOR2_X1 U845 ( .A1(n1161), .A2(n1180), .ZN(G60) );
XOR2_X1 U846 ( .A(n1181), .B(n1182), .Z(n1180) );
AND2_X1 U847 ( .A1(G475), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U848 ( .A(G104), .B(n1184), .ZN(G6) );
NAND4_X1 U849 ( .A1(n1185), .A2(n1068), .A3(n1186), .A4(n1070), .ZN(n1184) );
NOR2_X1 U850 ( .A1(KEYINPUT36), .A2(n1071), .ZN(n1186) );
NOR2_X1 U851 ( .A1(n1161), .A2(n1187), .ZN(G57) );
XOR2_X1 U852 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U853 ( .A(n1190), .B(n1191), .Z(n1188) );
AND2_X1 U854 ( .A1(G472), .A2(n1183), .ZN(n1191) );
NAND3_X1 U855 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1190) );
NAND3_X1 U856 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1193) );
INV_X1 U857 ( .A(n1198), .ZN(n1196) );
OR2_X1 U858 ( .A1(n1197), .A2(n1195), .ZN(n1192) );
INV_X1 U859 ( .A(n1199), .ZN(n1195) );
NAND2_X1 U860 ( .A1(n1200), .A2(n1201), .ZN(n1197) );
XOR2_X1 U861 ( .A(KEYINPUT3), .B(n1202), .Z(n1201) );
NOR2_X1 U862 ( .A1(n1161), .A2(n1203), .ZN(G54) );
XOR2_X1 U863 ( .A(n1204), .B(n1205), .Z(n1203) );
XNOR2_X1 U864 ( .A(n1206), .B(n1207), .ZN(n1205) );
XOR2_X1 U865 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR3_X1 U866 ( .A1(n1210), .A2(n1127), .A3(n1165), .ZN(n1209) );
INV_X1 U867 ( .A(G469), .ZN(n1127) );
XOR2_X1 U868 ( .A(KEYINPUT28), .B(KEYINPUT12), .Z(n1210) );
NAND2_X1 U869 ( .A1(n1211), .A2(KEYINPUT45), .ZN(n1208) );
XOR2_X1 U870 ( .A(n1212), .B(KEYINPUT49), .Z(n1211) );
XOR2_X1 U871 ( .A(n1213), .B(n1214), .Z(n1204) );
NOR2_X1 U872 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U873 ( .A(n1217), .B(KEYINPUT21), .Z(n1216) );
NAND2_X1 U874 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U875 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
OR2_X1 U876 ( .A1(n1222), .A2(KEYINPUT39), .ZN(n1220) );
NOR3_X1 U877 ( .A1(n1218), .A2(n1223), .A3(n1224), .ZN(n1215) );
NOR2_X1 U878 ( .A1(KEYINPUT39), .A2(n1222), .ZN(n1224) );
INV_X1 U879 ( .A(n1221), .ZN(n1223) );
NAND3_X1 U880 ( .A1(n1143), .A2(n1225), .A3(KEYINPUT39), .ZN(n1221) );
XNOR2_X1 U881 ( .A(KEYINPUT52), .B(KEYINPUT51), .ZN(n1213) );
NOR2_X1 U882 ( .A1(n1161), .A2(n1226), .ZN(G51) );
NOR2_X1 U883 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NOR2_X1 U884 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NOR2_X1 U885 ( .A1(n1231), .A2(n1232), .ZN(n1227) );
XOR2_X1 U886 ( .A(KEYINPUT20), .B(n1230), .Z(n1232) );
XNOR2_X1 U887 ( .A(n1233), .B(n1234), .ZN(n1230) );
NOR2_X1 U888 ( .A1(KEYINPUT41), .A2(n1158), .ZN(n1234) );
XOR2_X1 U889 ( .A(KEYINPUT0), .B(n1229), .Z(n1231) );
NOR2_X1 U890 ( .A1(n1165), .A2(n1117), .ZN(n1229) );
INV_X1 U891 ( .A(n1183), .ZN(n1165) );
NOR2_X1 U892 ( .A1(n1235), .A2(n1168), .ZN(n1183) );
NOR2_X1 U893 ( .A1(n1075), .A2(n1236), .ZN(n1168) );
XOR2_X1 U894 ( .A(KEYINPUT15), .B(n1077), .Z(n1236) );
NAND4_X1 U895 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1077) );
AND4_X1 U896 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1240) );
NOR2_X1 U897 ( .A1(n1245), .A2(n1246), .ZN(n1239) );
NAND4_X1 U898 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1075) );
NAND2_X1 U899 ( .A1(n1068), .A2(n1251), .ZN(n1247) );
NAND2_X1 U900 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U901 ( .A1(n1254), .A2(n1255), .ZN(n1252) );
NAND2_X1 U902 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U903 ( .A1(n1090), .A2(n1258), .ZN(n1257) );
NAND2_X1 U904 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND2_X1 U905 ( .A1(n1070), .A2(n1089), .ZN(n1256) );
OR2_X1 U906 ( .A1(n1185), .A2(n1069), .ZN(n1089) );
NOR2_X1 U907 ( .A1(n1081), .A2(G952), .ZN(n1161) );
XNOR2_X1 U908 ( .A(n1246), .B(n1261), .ZN(G48) );
NAND2_X1 U909 ( .A1(KEYINPUT30), .A2(G146), .ZN(n1261) );
AND3_X1 U910 ( .A1(n1185), .A2(n1102), .A3(n1262), .ZN(n1246) );
XOR2_X1 U911 ( .A(G143), .B(n1245), .Z(G45) );
AND4_X1 U912 ( .A1(n1263), .A2(n1102), .A3(n1264), .A4(n1265), .ZN(n1245) );
AND2_X1 U913 ( .A1(n1107), .A2(n1266), .ZN(n1265) );
NAND3_X1 U914 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(G42) );
NAND2_X1 U915 ( .A1(G140), .A2(n1237), .ZN(n1269) );
NAND2_X1 U916 ( .A1(KEYINPUT58), .A2(n1270), .ZN(n1268) );
NAND2_X1 U917 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U918 ( .A(KEYINPUT13), .B(G140), .Z(n1272) );
NAND2_X1 U919 ( .A1(n1273), .A2(n1274), .ZN(n1267) );
INV_X1 U920 ( .A(KEYINPUT58), .ZN(n1274) );
NAND2_X1 U921 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND3_X1 U922 ( .A1(KEYINPUT13), .A2(n1271), .A3(n1277), .ZN(n1276) );
INV_X1 U923 ( .A(n1237), .ZN(n1271) );
NAND4_X1 U924 ( .A1(n1083), .A2(n1266), .A3(n1096), .A4(n1185), .ZN(n1237) );
OR2_X1 U925 ( .A1(n1277), .A2(KEYINPUT13), .ZN(n1275) );
XOR2_X1 U926 ( .A(n1238), .B(n1278), .Z(G39) );
NAND2_X1 U927 ( .A1(KEYINPUT6), .A2(G137), .ZN(n1278) );
NAND3_X1 U928 ( .A1(n1262), .A2(n1090), .A3(n1083), .ZN(n1238) );
XNOR2_X1 U929 ( .A(G134), .B(n1244), .ZN(G36) );
NAND2_X1 U930 ( .A1(n1279), .A2(n1069), .ZN(n1244) );
XNOR2_X1 U931 ( .A(G131), .B(n1243), .ZN(G33) );
NAND2_X1 U932 ( .A1(n1279), .A2(n1185), .ZN(n1243) );
AND3_X1 U933 ( .A1(n1266), .A2(n1107), .A3(n1083), .ZN(n1279) );
NOR2_X1 U934 ( .A1(n1280), .A2(n1106), .ZN(n1083) );
XOR2_X1 U935 ( .A(n1105), .B(KEYINPUT63), .Z(n1280) );
XOR2_X1 U936 ( .A(n1281), .B(n1242), .Z(G30) );
NAND3_X1 U937 ( .A1(n1069), .A2(n1102), .A3(n1262), .ZN(n1242) );
AND3_X1 U938 ( .A1(n1282), .A2(n1283), .A3(n1266), .ZN(n1262) );
NOR2_X1 U939 ( .A1(n1071), .A2(n1284), .ZN(n1266) );
INV_X1 U940 ( .A(n1254), .ZN(n1071) );
XOR2_X1 U941 ( .A(G101), .B(n1285), .Z(G3) );
NOR4_X1 U942 ( .A1(n1286), .A2(n1287), .A3(n1259), .A4(n1086), .ZN(n1285) );
INV_X1 U943 ( .A(n1107), .ZN(n1259) );
NOR2_X1 U944 ( .A1(KEYINPUT1), .A2(n1288), .ZN(n1287) );
NOR2_X1 U945 ( .A1(n1068), .A2(n1289), .ZN(n1286) );
INV_X1 U946 ( .A(KEYINPUT1), .ZN(n1289) );
XNOR2_X1 U947 ( .A(G125), .B(n1241), .ZN(G27) );
NAND3_X1 U948 ( .A1(n1096), .A2(n1185), .A3(n1290), .ZN(n1241) );
NOR3_X1 U949 ( .A1(n1291), .A2(n1284), .A3(n1292), .ZN(n1290) );
AND2_X1 U950 ( .A1(n1293), .A2(n1294), .ZN(n1284) );
NAND4_X1 U951 ( .A1(G902), .A2(G953), .A3(n1108), .A4(n1137), .ZN(n1294) );
INV_X1 U952 ( .A(G900), .ZN(n1137) );
INV_X1 U953 ( .A(n1260), .ZN(n1096) );
XOR2_X1 U954 ( .A(G122), .B(n1295), .Z(G24) );
NOR3_X1 U955 ( .A1(n1253), .A2(n1296), .A3(n1297), .ZN(n1295) );
NOR2_X1 U956 ( .A1(n1288), .A2(n1298), .ZN(n1297) );
INV_X1 U957 ( .A(KEYINPUT7), .ZN(n1298) );
NOR2_X1 U958 ( .A1(n1299), .A2(n1102), .ZN(n1288) );
INV_X1 U959 ( .A(n1292), .ZN(n1102) );
NOR2_X1 U960 ( .A1(KEYINPUT7), .A2(n1068), .ZN(n1296) );
NAND4_X1 U961 ( .A1(n1264), .A2(n1088), .A3(n1263), .A4(n1070), .ZN(n1253) );
NOR2_X1 U962 ( .A1(n1283), .A2(n1282), .ZN(n1070) );
XNOR2_X1 U963 ( .A(G119), .B(n1248), .ZN(G21) );
NAND4_X1 U964 ( .A1(n1068), .A2(n1283), .A3(n1282), .A4(n1300), .ZN(n1248) );
AND2_X1 U965 ( .A1(n1088), .A2(n1090), .ZN(n1300) );
XOR2_X1 U966 ( .A(n1249), .B(n1301), .Z(G18) );
XNOR2_X1 U967 ( .A(G116), .B(KEYINPUT23), .ZN(n1301) );
NAND2_X1 U968 ( .A1(n1302), .A2(n1069), .ZN(n1249) );
AND2_X1 U969 ( .A1(n1263), .A2(n1303), .ZN(n1069) );
XNOR2_X1 U970 ( .A(G113), .B(n1250), .ZN(G15) );
NAND2_X1 U971 ( .A1(n1185), .A2(n1302), .ZN(n1250) );
AND3_X1 U972 ( .A1(n1088), .A2(n1068), .A3(n1107), .ZN(n1302) );
NOR2_X1 U973 ( .A1(n1304), .A2(n1283), .ZN(n1107) );
INV_X1 U974 ( .A(n1291), .ZN(n1088) );
NAND2_X1 U975 ( .A1(n1305), .A2(n1091), .ZN(n1291) );
NOR2_X1 U976 ( .A1(n1303), .A2(n1263), .ZN(n1185) );
INV_X1 U977 ( .A(n1264), .ZN(n1303) );
XOR2_X1 U978 ( .A(G110), .B(n1306), .Z(G12) );
NOR4_X1 U979 ( .A1(n1307), .A2(n1308), .A3(n1260), .A4(n1086), .ZN(n1306) );
NAND2_X1 U980 ( .A1(n1090), .A2(n1254), .ZN(n1086) );
NOR2_X1 U981 ( .A1(n1091), .A2(n1092), .ZN(n1254) );
INV_X1 U982 ( .A(n1305), .ZN(n1092) );
NAND2_X1 U983 ( .A1(G221), .A2(n1309), .ZN(n1305) );
NAND3_X1 U984 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1091) );
NAND2_X1 U985 ( .A1(G469), .A2(n1313), .ZN(n1312) );
NAND2_X1 U986 ( .A1(n1314), .A2(n1128), .ZN(n1313) );
NAND3_X1 U987 ( .A1(n1315), .A2(n1128), .A3(n1316), .ZN(n1311) );
INV_X1 U988 ( .A(n1314), .ZN(n1315) );
XOR2_X1 U989 ( .A(n1317), .B(G469), .Z(n1314) );
XNOR2_X1 U990 ( .A(KEYINPUT60), .B(KEYINPUT29), .ZN(n1317) );
OR2_X1 U991 ( .A1(n1128), .A2(n1316), .ZN(n1310) );
INV_X1 U992 ( .A(KEYINPUT38), .ZN(n1316) );
NAND4_X1 U993 ( .A1(n1318), .A2(n1235), .A3(n1319), .A4(n1320), .ZN(n1128) );
OR2_X1 U994 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND4_X1 U995 ( .A1(n1323), .A2(n1321), .A3(KEYINPUT56), .A4(n1322), .ZN(n1319) );
INV_X1 U996 ( .A(KEYINPUT62), .ZN(n1321) );
XOR2_X1 U997 ( .A(n1222), .B(n1202), .Z(n1323) );
NAND2_X1 U998 ( .A1(n1324), .A2(n1325), .ZN(n1318) );
NAND2_X1 U999 ( .A1(KEYINPUT56), .A2(n1322), .ZN(n1325) );
XNOR2_X1 U1000 ( .A(n1212), .B(n1206), .ZN(n1322) );
XNOR2_X1 U1001 ( .A(n1326), .B(G140), .ZN(n1206) );
NAND2_X1 U1002 ( .A1(G227), .A2(n1081), .ZN(n1212) );
XOR2_X1 U1003 ( .A(n1218), .B(n1222), .Z(n1324) );
XOR2_X1 U1004 ( .A(n1143), .B(n1327), .Z(n1222) );
INV_X1 U1005 ( .A(n1225), .ZN(n1327) );
XOR2_X1 U1006 ( .A(n1328), .B(KEYINPUT61), .Z(n1143) );
NOR2_X1 U1007 ( .A1(n1264), .A2(n1263), .ZN(n1090) );
XOR2_X1 U1008 ( .A(n1329), .B(n1126), .Z(n1263) );
NOR2_X1 U1009 ( .A1(n1174), .A2(G902), .ZN(n1126) );
XNOR2_X1 U1010 ( .A(n1330), .B(n1331), .ZN(n1174) );
XOR2_X1 U1011 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1012 ( .A(G107), .B(n1334), .Z(n1333) );
AND3_X1 U1013 ( .A1(G217), .A2(n1081), .A3(G234), .ZN(n1334) );
XOR2_X1 U1014 ( .A(G143), .B(G116), .Z(n1332) );
XOR2_X1 U1015 ( .A(n1335), .B(n1336), .Z(n1330) );
XNOR2_X1 U1016 ( .A(n1337), .B(n1338), .ZN(n1336) );
NOR2_X1 U1017 ( .A1(G122), .A2(KEYINPUT57), .ZN(n1338) );
NAND2_X1 U1018 ( .A1(KEYINPUT33), .A2(n1339), .ZN(n1337) );
INV_X1 U1019 ( .A(n1142), .ZN(n1339) );
NAND2_X1 U1020 ( .A1(KEYINPUT53), .A2(n1281), .ZN(n1335) );
NAND2_X1 U1021 ( .A1(KEYINPUT50), .A2(n1178), .ZN(n1329) );
INV_X1 U1022 ( .A(G478), .ZN(n1178) );
XOR2_X1 U1023 ( .A(n1115), .B(KEYINPUT31), .Z(n1264) );
XOR2_X1 U1024 ( .A(n1340), .B(G475), .Z(n1115) );
OR2_X1 U1025 ( .A1(n1182), .A2(G902), .ZN(n1340) );
XNOR2_X1 U1026 ( .A(n1341), .B(n1342), .ZN(n1182) );
XOR2_X1 U1027 ( .A(n1343), .B(n1344), .Z(n1342) );
NAND2_X1 U1028 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1029 ( .A1(G146), .A2(n1347), .ZN(n1346) );
NAND2_X1 U1030 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XNOR2_X1 U1031 ( .A(KEYINPUT14), .B(n1350), .ZN(n1348) );
NAND2_X1 U1032 ( .A1(n1351), .A2(n1352), .ZN(n1345) );
NAND2_X1 U1033 ( .A1(n1353), .A2(n1354), .ZN(n1351) );
OR2_X1 U1034 ( .A1(n1350), .A2(KEYINPUT14), .ZN(n1354) );
NAND2_X1 U1035 ( .A1(n1140), .A2(KEYINPUT14), .ZN(n1353) );
INV_X1 U1036 ( .A(n1355), .ZN(n1140) );
NAND2_X1 U1037 ( .A1(n1356), .A2(KEYINPUT37), .ZN(n1343) );
XNOR2_X1 U1038 ( .A(G104), .B(n1357), .ZN(n1356) );
XOR2_X1 U1039 ( .A(n1358), .B(n1359), .Z(n1341) );
NOR4_X1 U1040 ( .A1(KEYINPUT22), .A2(G953), .A3(G237), .A4(n1360), .ZN(n1359) );
INV_X1 U1041 ( .A(G214), .ZN(n1360) );
XNOR2_X1 U1042 ( .A(G131), .B(G143), .ZN(n1358) );
NAND2_X1 U1043 ( .A1(n1304), .A2(n1283), .ZN(n1260) );
NAND2_X1 U1044 ( .A1(n1361), .A2(n1362), .ZN(n1283) );
NAND2_X1 U1045 ( .A1(n1363), .A2(n1125), .ZN(n1362) );
XOR2_X1 U1046 ( .A(KEYINPUT18), .B(n1364), .Z(n1361) );
NOR2_X1 U1047 ( .A1(n1363), .A2(n1125), .ZN(n1364) );
NAND2_X1 U1048 ( .A1(G217), .A2(n1309), .ZN(n1125) );
NAND2_X1 U1049 ( .A1(G234), .A2(n1235), .ZN(n1309) );
XNOR2_X1 U1050 ( .A(n1124), .B(KEYINPUT10), .ZN(n1363) );
NOR2_X1 U1051 ( .A1(n1167), .A2(G902), .ZN(n1124) );
INV_X1 U1052 ( .A(n1164), .ZN(n1167) );
XOR2_X1 U1053 ( .A(n1365), .B(n1366), .Z(n1164) );
AND3_X1 U1054 ( .A1(G221), .A2(n1081), .A3(G234), .ZN(n1366) );
XOR2_X1 U1055 ( .A(n1367), .B(G137), .Z(n1365) );
NAND2_X1 U1056 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
NAND2_X1 U1057 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1058 ( .A(n1372), .B(KEYINPUT46), .Z(n1368) );
OR2_X1 U1059 ( .A1(n1371), .A2(n1370), .ZN(n1372) );
XOR2_X1 U1060 ( .A(n1355), .B(n1352), .Z(n1370) );
INV_X1 U1061 ( .A(G146), .ZN(n1352) );
NAND2_X1 U1062 ( .A1(n1350), .A2(n1349), .ZN(n1355) );
NAND2_X1 U1063 ( .A1(G125), .A2(n1277), .ZN(n1349) );
OR2_X1 U1064 ( .A1(n1277), .A2(G125), .ZN(n1350) );
INV_X1 U1065 ( .A(G140), .ZN(n1277) );
XNOR2_X1 U1066 ( .A(n1326), .B(n1373), .ZN(n1371) );
XOR2_X1 U1067 ( .A(G128), .B(G119), .Z(n1373) );
INV_X1 U1068 ( .A(G110), .ZN(n1326) );
INV_X1 U1069 ( .A(n1282), .ZN(n1304) );
XOR2_X1 U1070 ( .A(n1374), .B(n1375), .Z(n1282) );
INV_X1 U1071 ( .A(n1129), .ZN(n1375) );
XNOR2_X1 U1072 ( .A(G472), .B(KEYINPUT8), .ZN(n1129) );
NAND2_X1 U1073 ( .A1(KEYINPUT26), .A2(n1130), .ZN(n1374) );
AND2_X1 U1074 ( .A1(n1376), .A2(n1235), .ZN(n1130) );
XNOR2_X1 U1075 ( .A(n1377), .B(n1189), .ZN(n1376) );
XNOR2_X1 U1076 ( .A(n1378), .B(G101), .ZN(n1189) );
NAND3_X1 U1077 ( .A1(n1379), .A2(n1081), .A3(G210), .ZN(n1378) );
NAND3_X1 U1078 ( .A1(n1380), .A2(n1381), .A3(n1194), .ZN(n1377) );
NAND2_X1 U1079 ( .A1(n1198), .A2(n1199), .ZN(n1194) );
NOR2_X1 U1080 ( .A1(n1200), .A2(n1218), .ZN(n1198) );
NAND2_X1 U1081 ( .A1(n1382), .A2(n1200), .ZN(n1381) );
XOR2_X1 U1082 ( .A(n1199), .B(n1202), .Z(n1382) );
OR3_X1 U1083 ( .A1(n1199), .A2(n1202), .A3(n1200), .ZN(n1380) );
INV_X1 U1084 ( .A(n1218), .ZN(n1202) );
XOR2_X1 U1085 ( .A(n1142), .B(n1144), .Z(n1218) );
XOR2_X1 U1086 ( .A(G131), .B(G137), .Z(n1144) );
XNOR2_X1 U1087 ( .A(G134), .B(KEYINPUT17), .ZN(n1142) );
XNOR2_X1 U1088 ( .A(G113), .B(n1383), .ZN(n1199) );
NOR2_X1 U1089 ( .A1(n1384), .A2(n1385), .ZN(n1308) );
INV_X1 U1090 ( .A(KEYINPUT47), .ZN(n1385) );
NOR2_X1 U1091 ( .A1(n1292), .A2(n1386), .ZN(n1384) );
NOR2_X1 U1092 ( .A1(KEYINPUT47), .A2(n1068), .ZN(n1307) );
NOR2_X1 U1093 ( .A1(n1292), .A2(n1299), .ZN(n1068) );
INV_X1 U1094 ( .A(n1386), .ZN(n1299) );
NAND2_X1 U1095 ( .A1(n1293), .A2(n1387), .ZN(n1386) );
NAND3_X1 U1096 ( .A1(n1157), .A2(n1108), .A3(G902), .ZN(n1387) );
NOR2_X1 U1097 ( .A1(G898), .A2(n1081), .ZN(n1157) );
NAND3_X1 U1098 ( .A1(n1108), .A2(n1081), .A3(G952), .ZN(n1293) );
INV_X1 U1099 ( .A(G953), .ZN(n1081) );
NAND2_X1 U1100 ( .A1(G234), .A2(G237), .ZN(n1108) );
NAND2_X1 U1101 ( .A1(n1388), .A2(n1106), .ZN(n1292) );
XNOR2_X1 U1102 ( .A(n1119), .B(n1117), .ZN(n1106) );
NAND2_X1 U1103 ( .A1(G210), .A2(n1389), .ZN(n1117) );
AND2_X1 U1104 ( .A1(n1390), .A2(n1235), .ZN(n1119) );
XOR2_X1 U1105 ( .A(n1233), .B(n1391), .Z(n1390) );
INV_X1 U1106 ( .A(n1158), .ZN(n1391) );
XOR2_X1 U1107 ( .A(n1392), .B(n1393), .Z(n1158) );
XOR2_X1 U1108 ( .A(n1394), .B(n1395), .Z(n1393) );
XOR2_X1 U1109 ( .A(KEYINPUT9), .B(G110), .Z(n1395) );
NOR2_X1 U1110 ( .A1(KEYINPUT24), .A2(n1383), .ZN(n1394) );
XOR2_X1 U1111 ( .A(G116), .B(G119), .Z(n1383) );
XOR2_X1 U1112 ( .A(n1225), .B(n1357), .Z(n1392) );
XOR2_X1 U1113 ( .A(G113), .B(G122), .Z(n1357) );
XNOR2_X1 U1114 ( .A(G101), .B(n1396), .ZN(n1225) );
XOR2_X1 U1115 ( .A(G107), .B(G104), .Z(n1396) );
XOR2_X1 U1116 ( .A(n1200), .B(n1397), .Z(n1233) );
XOR2_X1 U1117 ( .A(G125), .B(n1398), .Z(n1397) );
NOR2_X1 U1118 ( .A1(G953), .A2(n1155), .ZN(n1398) );
INV_X1 U1119 ( .A(G224), .ZN(n1155) );
XOR2_X1 U1120 ( .A(n1328), .B(KEYINPUT32), .Z(n1200) );
XOR2_X1 U1121 ( .A(n1281), .B(n1399), .Z(n1328) );
XOR2_X1 U1122 ( .A(G146), .B(G143), .Z(n1399) );
INV_X1 U1123 ( .A(G128), .ZN(n1281) );
XNOR2_X1 U1124 ( .A(n1105), .B(KEYINPUT63), .ZN(n1388) );
AND2_X1 U1125 ( .A1(G214), .A2(n1389), .ZN(n1105) );
NAND2_X1 U1126 ( .A1(n1400), .A2(n1235), .ZN(n1389) );
INV_X1 U1127 ( .A(G902), .ZN(n1235) );
XOR2_X1 U1128 ( .A(n1379), .B(KEYINPUT34), .Z(n1400) );
INV_X1 U1129 ( .A(G237), .ZN(n1379) );
endmodule


