//Key = 0111010000100101010101001110011111101101010010110011000100001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;

XNOR2_X1 U736 ( .A(G107), .B(n1012), .ZN(G9) );
NOR2_X1 U737 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1014) );
NOR2_X1 U739 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
NOR2_X1 U740 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR3_X1 U741 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NOR2_X1 U742 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(n1026) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U746 ( .A1(n1034), .A2(n1028), .ZN(n1033) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1032) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR4_X1 U749 ( .A1(n1039), .A2(n1031), .A3(n1028), .A4(n1036), .ZN(n1021) );
NOR2_X1 U750 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1025), .ZN(n1041) );
INV_X1 U752 ( .A(n1043), .ZN(n1025) );
NOR3_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1042) );
AND3_X1 U754 ( .A1(KEYINPUT10), .A2(n1047), .A3(n1048), .ZN(n1046) );
NOR2_X1 U755 ( .A1(KEYINPUT10), .A2(n1023), .ZN(n1045) );
NOR2_X1 U756 ( .A1(n1049), .A2(n1023), .ZN(n1040) );
NOR2_X1 U757 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR3_X1 U759 ( .A1(n1018), .A2(G952), .A3(n1015), .ZN(n1013) );
AND4_X1 U760 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1015) );
NOR4_X1 U761 ( .A1(n1048), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1057) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
INV_X1 U763 ( .A(n1063), .ZN(n1059) );
NOR2_X1 U764 ( .A1(n1028), .A2(n1064), .ZN(n1056) );
XNOR2_X1 U765 ( .A(G472), .B(n1065), .ZN(n1064) );
XOR2_X1 U766 ( .A(n1066), .B(n1067), .Z(G72) );
NAND2_X1 U767 ( .A1(G953), .A2(n1068), .ZN(n1067) );
NAND2_X1 U768 ( .A1(G900), .A2(G227), .ZN(n1068) );
NAND3_X1 U769 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1066) );
NAND2_X1 U770 ( .A1(KEYINPUT27), .A2(n1072), .ZN(n1071) );
INV_X1 U771 ( .A(n1073), .ZN(n1072) );
OR3_X1 U772 ( .A1(n1074), .A2(KEYINPUT27), .A3(n1075), .ZN(n1070) );
NAND2_X1 U773 ( .A1(n1075), .A2(n1074), .ZN(n1069) );
NAND2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
XOR2_X1 U775 ( .A(KEYINPUT39), .B(n1078), .Z(n1077) );
XOR2_X1 U776 ( .A(n1079), .B(n1080), .Z(n1076) );
XNOR2_X1 U777 ( .A(n1081), .B(n1082), .ZN(n1080) );
NAND2_X1 U778 ( .A1(KEYINPUT32), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U779 ( .A(n1084), .B(n1085), .ZN(n1079) );
NAND2_X1 U780 ( .A1(KEYINPUT34), .A2(n1073), .ZN(n1075) );
NOR2_X1 U781 ( .A1(n1086), .A2(G953), .ZN(n1073) );
NAND2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(G69) );
NAND2_X1 U783 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(n1087) );
NAND2_X1 U785 ( .A1(n1093), .A2(n1090), .ZN(n1092) );
NAND2_X1 U786 ( .A1(G953), .A2(n1094), .ZN(n1090) );
INV_X1 U787 ( .A(n1089), .ZN(n1091) );
XNOR2_X1 U788 ( .A(n1095), .B(n1096), .ZN(n1089) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U790 ( .A(n1099), .B(n1100), .Z(n1098) );
XNOR2_X1 U791 ( .A(n1101), .B(n1102), .ZN(n1100) );
NAND2_X1 U792 ( .A1(KEYINPUT50), .A2(n1103), .ZN(n1101) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(n1095) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U795 ( .A(n1108), .B(KEYINPUT63), .Z(n1106) );
NOR2_X1 U796 ( .A1(n1109), .A2(n1110), .ZN(G66) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND3_X1 U798 ( .A1(G902), .A2(n1113), .A3(n1114), .ZN(n1112) );
XNOR2_X1 U799 ( .A(KEYINPUT17), .B(n1017), .ZN(n1113) );
NOR2_X1 U800 ( .A1(n1109), .A2(n1115), .ZN(G63) );
XOR2_X1 U801 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NOR3_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(G60) );
AND2_X1 U804 ( .A1(KEYINPUT46), .A2(n1109), .ZN(n1122) );
NOR3_X1 U805 ( .A1(KEYINPUT46), .A2(G953), .A3(G952), .ZN(n1121) );
XOR2_X1 U806 ( .A(n1123), .B(n1124), .Z(n1120) );
NOR2_X1 U807 ( .A1(n1125), .A2(n1119), .ZN(n1123) );
XNOR2_X1 U808 ( .A(G104), .B(n1126), .ZN(G6) );
NAND2_X1 U809 ( .A1(KEYINPUT47), .A2(n1127), .ZN(n1126) );
NOR2_X1 U810 ( .A1(n1109), .A2(n1128), .ZN(G57) );
XNOR2_X1 U811 ( .A(n1129), .B(n1130), .ZN(n1128) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1119), .ZN(n1131) );
NOR2_X1 U814 ( .A1(n1109), .A2(n1134), .ZN(G54) );
XOR2_X1 U815 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U816 ( .A(n1137), .B(n1138), .ZN(n1136) );
XOR2_X1 U817 ( .A(n1139), .B(n1140), .Z(n1135) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1119), .ZN(n1140) );
INV_X1 U819 ( .A(G469), .ZN(n1141) );
NAND2_X1 U820 ( .A1(KEYINPUT31), .A2(G110), .ZN(n1139) );
NOR2_X1 U821 ( .A1(n1109), .A2(n1142), .ZN(G51) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U823 ( .A(KEYINPUT2), .B(n1145), .Z(n1144) );
XOR2_X1 U824 ( .A(n1146), .B(n1147), .Z(n1143) );
NOR3_X1 U825 ( .A1(n1148), .A2(n1149), .A3(n1119), .ZN(n1147) );
NAND2_X1 U826 ( .A1(G902), .A2(n1017), .ZN(n1119) );
NAND3_X1 U827 ( .A1(n1086), .A2(n1108), .A3(n1107), .ZN(n1017) );
AND4_X1 U828 ( .A1(n1150), .A2(n1012), .A3(n1151), .A4(n1152), .ZN(n1107) );
NOR4_X1 U829 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1127), .ZN(n1152) );
AND3_X1 U830 ( .A1(n1156), .A2(n1051), .A3(n1038), .ZN(n1127) );
NAND3_X1 U831 ( .A1(n1156), .A2(n1051), .A3(n1037), .ZN(n1012) );
AND4_X1 U832 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1086) );
AND4_X1 U833 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
NAND2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(n1159) );
XNOR2_X1 U835 ( .A(KEYINPUT0), .B(n1167), .ZN(n1166) );
NAND3_X1 U836 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1157) );
NAND2_X1 U837 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
NAND3_X1 U838 ( .A1(n1173), .A2(n1174), .A3(n1044), .ZN(n1172) );
NAND2_X1 U839 ( .A1(n1165), .A2(n1037), .ZN(n1171) );
XOR2_X1 U840 ( .A(KEYINPUT18), .B(n1175), .Z(n1148) );
NOR2_X1 U841 ( .A1(n1104), .A2(G952), .ZN(n1109) );
NAND2_X1 U842 ( .A1(n1176), .A2(n1177), .ZN(G48) );
NAND2_X1 U843 ( .A1(G146), .A2(n1178), .ZN(n1177) );
NAND2_X1 U844 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
OR2_X1 U845 ( .A1(KEYINPUT38), .A2(KEYINPUT44), .ZN(n1180) );
NAND3_X1 U846 ( .A1(n1181), .A2(n1182), .A3(KEYINPUT44), .ZN(n1176) );
OR2_X1 U847 ( .A1(n1179), .A2(KEYINPUT38), .ZN(n1182) );
NAND2_X1 U848 ( .A1(n1179), .A2(n1183), .ZN(n1181) );
OR2_X1 U849 ( .A1(G146), .A2(KEYINPUT38), .ZN(n1183) );
INV_X1 U850 ( .A(n1158), .ZN(n1179) );
NAND3_X1 U851 ( .A1(n1038), .A2(n1044), .A3(n1184), .ZN(n1158) );
XNOR2_X1 U852 ( .A(G143), .B(n1185), .ZN(G45) );
NAND3_X1 U853 ( .A1(n1186), .A2(n1170), .A3(n1187), .ZN(n1185) );
AND3_X1 U854 ( .A1(n1044), .A2(n1174), .A3(n1173), .ZN(n1187) );
XNOR2_X1 U855 ( .A(n1168), .B(KEYINPUT19), .ZN(n1186) );
NAND2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(G42) );
NAND2_X1 U857 ( .A1(KEYINPUT23), .A2(G140), .ZN(n1189) );
XOR2_X1 U858 ( .A(n1190), .B(n1191), .Z(n1188) );
NOR2_X1 U859 ( .A1(n1023), .A2(n1167), .ZN(n1191) );
NAND2_X1 U860 ( .A1(n1170), .A2(n1192), .ZN(n1167) );
INV_X1 U861 ( .A(n1165), .ZN(n1023) );
NOR2_X1 U862 ( .A1(G140), .A2(KEYINPUT23), .ZN(n1190) );
XNOR2_X1 U863 ( .A(G137), .B(n1164), .ZN(G39) );
NAND3_X1 U864 ( .A1(n1184), .A2(n1193), .A3(n1165), .ZN(n1164) );
XNOR2_X1 U865 ( .A(G134), .B(n1194), .ZN(G36) );
NAND4_X1 U866 ( .A1(n1165), .A2(n1170), .A3(n1037), .A4(n1195), .ZN(n1194) );
XNOR2_X1 U867 ( .A(KEYINPUT16), .B(n1029), .ZN(n1195) );
INV_X1 U868 ( .A(n1168), .ZN(n1029) );
XNOR2_X1 U869 ( .A(G131), .B(n1163), .ZN(G33) );
NAND4_X1 U870 ( .A1(n1165), .A2(n1170), .A3(n1168), .A4(n1038), .ZN(n1163) );
NOR2_X1 U871 ( .A1(n1196), .A2(n1048), .ZN(n1165) );
XNOR2_X1 U872 ( .A(G128), .B(n1162), .ZN(G30) );
NAND3_X1 U873 ( .A1(n1037), .A2(n1044), .A3(n1184), .ZN(n1162) );
AND3_X1 U874 ( .A1(n1031), .A2(n1197), .A3(n1170), .ZN(n1184) );
AND2_X1 U875 ( .A1(n1051), .A2(n1198), .ZN(n1170) );
XOR2_X1 U876 ( .A(n1199), .B(n1155), .Z(G3) );
AND2_X1 U877 ( .A1(n1168), .A2(n1200), .ZN(n1155) );
XNOR2_X1 U878 ( .A(G101), .B(KEYINPUT15), .ZN(n1199) );
XNOR2_X1 U879 ( .A(G125), .B(n1161), .ZN(G27) );
NAND4_X1 U880 ( .A1(n1192), .A2(n1043), .A3(n1044), .A4(n1198), .ZN(n1161) );
NAND2_X1 U881 ( .A1(n1201), .A2(n1020), .ZN(n1198) );
XOR2_X1 U882 ( .A(n1202), .B(KEYINPUT9), .Z(n1201) );
NAND2_X1 U883 ( .A1(n1078), .A2(n1203), .ZN(n1202) );
INV_X1 U884 ( .A(n1204), .ZN(n1203) );
NOR2_X1 U885 ( .A1(n1104), .A2(G900), .ZN(n1078) );
AND3_X1 U886 ( .A1(n1197), .A2(n1205), .A3(n1038), .ZN(n1192) );
XOR2_X1 U887 ( .A(n1151), .B(n1206), .Z(G24) );
NAND2_X1 U888 ( .A1(KEYINPUT33), .A2(G122), .ZN(n1206) );
NAND4_X1 U889 ( .A1(n1156), .A2(n1043), .A3(n1173), .A4(n1174), .ZN(n1151) );
NOR3_X1 U890 ( .A1(n1036), .A2(n1031), .A3(n1207), .ZN(n1156) );
XNOR2_X1 U891 ( .A(G119), .B(n1150), .ZN(G21) );
NAND4_X1 U892 ( .A1(n1031), .A2(n1193), .A3(n1208), .A4(n1043), .ZN(n1150) );
NOR2_X1 U893 ( .A1(n1034), .A2(n1207), .ZN(n1208) );
INV_X1 U894 ( .A(n1197), .ZN(n1034) );
XNOR2_X1 U895 ( .A(G116), .B(n1108), .ZN(G18) );
NAND4_X1 U896 ( .A1(n1168), .A2(n1037), .A3(n1043), .A4(n1209), .ZN(n1108) );
AND2_X1 U897 ( .A1(n1210), .A2(n1173), .ZN(n1037) );
XOR2_X1 U898 ( .A(n1211), .B(KEYINPUT60), .Z(n1173) );
NAND2_X1 U899 ( .A1(n1212), .A2(n1213), .ZN(G15) );
NAND2_X1 U900 ( .A1(n1214), .A2(n1154), .ZN(n1213) );
XNOR2_X1 U901 ( .A(G113), .B(KEYINPUT43), .ZN(n1214) );
XOR2_X1 U902 ( .A(KEYINPUT55), .B(n1215), .Z(n1212) );
NOR2_X1 U903 ( .A1(n1154), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U904 ( .A(G113), .B(KEYINPUT57), .ZN(n1216) );
AND4_X1 U905 ( .A1(n1168), .A2(n1038), .A3(n1043), .A4(n1209), .ZN(n1154) );
AND2_X1 U906 ( .A1(n1211), .A2(n1174), .ZN(n1038) );
NOR2_X1 U907 ( .A1(n1217), .A2(n1036), .ZN(n1168) );
XOR2_X1 U908 ( .A(n1197), .B(KEYINPUT12), .Z(n1036) );
XNOR2_X1 U909 ( .A(n1031), .B(KEYINPUT58), .ZN(n1217) );
INV_X1 U910 ( .A(n1205), .ZN(n1031) );
XNOR2_X1 U911 ( .A(G110), .B(n1218), .ZN(G12) );
NAND2_X1 U912 ( .A1(KEYINPUT26), .A2(n1153), .ZN(n1218) );
AND3_X1 U913 ( .A1(n1197), .A2(n1205), .A3(n1200), .ZN(n1153) );
AND3_X1 U914 ( .A1(n1209), .A2(n1051), .A3(n1193), .ZN(n1200) );
INV_X1 U915 ( .A(n1028), .ZN(n1193) );
NAND2_X1 U916 ( .A1(n1210), .A2(n1211), .ZN(n1028) );
XNOR2_X1 U917 ( .A(n1219), .B(n1118), .ZN(n1211) );
INV_X1 U918 ( .A(G478), .ZN(n1118) );
OR2_X1 U919 ( .A1(n1117), .A2(G902), .ZN(n1219) );
XNOR2_X1 U920 ( .A(n1220), .B(n1221), .ZN(n1117) );
AND2_X1 U921 ( .A1(n1222), .A2(G217), .ZN(n1221) );
NAND2_X1 U922 ( .A1(n1223), .A2(n1224), .ZN(n1220) );
OR2_X1 U923 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U924 ( .A(n1227), .B(KEYINPUT62), .Z(n1223) );
NAND2_X1 U925 ( .A1(n1226), .A2(n1225), .ZN(n1227) );
XOR2_X1 U926 ( .A(G107), .B(n1228), .Z(n1225) );
XNOR2_X1 U927 ( .A(G122), .B(n1229), .ZN(n1228) );
XNOR2_X1 U928 ( .A(n1230), .B(n1231), .ZN(n1226) );
NOR2_X1 U929 ( .A1(G143), .A2(KEYINPUT49), .ZN(n1231) );
XNOR2_X1 U930 ( .A(G134), .B(G128), .ZN(n1230) );
INV_X1 U931 ( .A(n1174), .ZN(n1210) );
XOR2_X1 U932 ( .A(n1232), .B(n1125), .Z(n1174) );
INV_X1 U933 ( .A(G475), .ZN(n1125) );
OR2_X1 U934 ( .A1(n1124), .A2(G902), .ZN(n1232) );
XNOR2_X1 U935 ( .A(n1233), .B(n1234), .ZN(n1124) );
XNOR2_X1 U936 ( .A(n1235), .B(n1236), .ZN(n1234) );
XOR2_X1 U937 ( .A(n1237), .B(n1238), .Z(n1233) );
AND2_X1 U938 ( .A1(n1239), .A2(G214), .ZN(n1238) );
XNOR2_X1 U939 ( .A(n1240), .B(n1085), .ZN(n1237) );
INV_X1 U940 ( .A(G131), .ZN(n1085) );
NAND4_X1 U941 ( .A1(KEYINPUT36), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1240) );
NAND3_X1 U942 ( .A1(KEYINPUT30), .A2(n1244), .A3(n1245), .ZN(n1243) );
OR2_X1 U943 ( .A1(n1245), .A2(n1244), .ZN(n1242) );
NOR2_X1 U944 ( .A1(G104), .A2(KEYINPUT54), .ZN(n1244) );
XOR2_X1 U945 ( .A(G122), .B(n1246), .Z(n1245) );
OR2_X1 U946 ( .A1(n1247), .A2(KEYINPUT30), .ZN(n1241) );
INV_X1 U947 ( .A(G104), .ZN(n1247) );
NAND2_X1 U948 ( .A1(n1248), .A2(n1249), .ZN(n1051) );
OR3_X1 U949 ( .A1(n1250), .A2(n1251), .A3(KEYINPUT59), .ZN(n1249) );
INV_X1 U950 ( .A(n1052), .ZN(n1251) );
NAND2_X1 U951 ( .A1(KEYINPUT59), .A2(n1043), .ZN(n1248) );
NOR2_X1 U952 ( .A1(n1250), .A2(n1052), .ZN(n1043) );
XOR2_X1 U953 ( .A(n1055), .B(KEYINPUT5), .Z(n1052) );
XNOR2_X1 U954 ( .A(G469), .B(n1252), .ZN(n1055) );
NOR2_X1 U955 ( .A1(G902), .A2(n1253), .ZN(n1252) );
XOR2_X1 U956 ( .A(n1138), .B(n1254), .Z(n1253) );
XNOR2_X1 U957 ( .A(n1255), .B(n1256), .ZN(n1254) );
NOR2_X1 U958 ( .A1(KEYINPUT48), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U959 ( .A(KEYINPUT21), .B(n1258), .ZN(n1257) );
INV_X1 U960 ( .A(n1137), .ZN(n1258) );
XNOR2_X1 U961 ( .A(n1259), .B(n1260), .ZN(n1137) );
XNOR2_X1 U962 ( .A(G107), .B(n1261), .ZN(n1260) );
XOR2_X1 U963 ( .A(n1084), .B(n1262), .Z(n1259) );
NOR2_X1 U964 ( .A1(G104), .A2(KEYINPUT35), .ZN(n1262) );
NAND2_X1 U965 ( .A1(n1263), .A2(n1264), .ZN(n1084) );
NAND2_X1 U966 ( .A1(G128), .A2(n1235), .ZN(n1264) );
XOR2_X1 U967 ( .A(KEYINPUT25), .B(n1265), .Z(n1263) );
NOR2_X1 U968 ( .A1(G128), .A2(n1235), .ZN(n1265) );
XNOR2_X1 U969 ( .A(n1266), .B(n1267), .ZN(n1138) );
XOR2_X1 U970 ( .A(G140), .B(n1268), .Z(n1267) );
AND2_X1 U971 ( .A1(n1104), .A2(G227), .ZN(n1268) );
XOR2_X1 U972 ( .A(n1058), .B(KEYINPUT45), .Z(n1250) );
INV_X1 U973 ( .A(n1053), .ZN(n1058) );
NAND2_X1 U974 ( .A1(G221), .A2(n1269), .ZN(n1053) );
INV_X1 U975 ( .A(n1207), .ZN(n1209) );
NAND2_X1 U976 ( .A1(n1044), .A2(n1270), .ZN(n1207) );
NAND2_X1 U977 ( .A1(n1271), .A2(n1020), .ZN(n1270) );
NAND3_X1 U978 ( .A1(n1272), .A2(n1273), .A3(G952), .ZN(n1020) );
INV_X1 U979 ( .A(n1018), .ZN(n1272) );
XOR2_X1 U980 ( .A(G953), .B(KEYINPUT52), .Z(n1018) );
XOR2_X1 U981 ( .A(KEYINPUT13), .B(n1274), .Z(n1271) );
NOR2_X1 U982 ( .A1(n1204), .A2(n1093), .ZN(n1274) );
INV_X1 U983 ( .A(n1097), .ZN(n1093) );
NOR2_X1 U984 ( .A1(G898), .A2(n1104), .ZN(n1097) );
NAND2_X1 U985 ( .A1(G902), .A2(n1273), .ZN(n1204) );
NAND2_X1 U986 ( .A1(G237), .A2(G234), .ZN(n1273) );
NOR2_X1 U987 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NOR2_X1 U988 ( .A1(n1275), .A2(n1175), .ZN(n1048) );
INV_X1 U989 ( .A(G214), .ZN(n1275) );
INV_X1 U990 ( .A(n1196), .ZN(n1047) );
NAND3_X1 U991 ( .A1(n1276), .A2(n1277), .A3(n1063), .ZN(n1196) );
NAND2_X1 U992 ( .A1(n1061), .A2(n1062), .ZN(n1063) );
NAND2_X1 U993 ( .A1(KEYINPUT4), .A2(n1062), .ZN(n1277) );
OR3_X1 U994 ( .A1(n1061), .A2(KEYINPUT4), .A3(n1062), .ZN(n1276) );
NAND3_X1 U995 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1062) );
XOR2_X1 U996 ( .A(KEYINPUT29), .B(n1281), .Z(n1280) );
NOR2_X1 U997 ( .A1(n1145), .A2(n1146), .ZN(n1281) );
NAND2_X1 U998 ( .A1(n1145), .A2(n1146), .ZN(n1278) );
XOR2_X1 U999 ( .A(n1282), .B(n1283), .Z(n1146) );
XNOR2_X1 U1000 ( .A(n1284), .B(n1285), .ZN(n1283) );
NOR2_X1 U1001 ( .A1(G953), .A2(n1094), .ZN(n1285) );
INV_X1 U1002 ( .A(G224), .ZN(n1094) );
INV_X1 U1003 ( .A(G125), .ZN(n1284) );
AND2_X1 U1004 ( .A1(n1286), .A2(n1287), .ZN(n1145) );
NAND2_X1 U1005 ( .A1(n1288), .A2(n1099), .ZN(n1287) );
XNOR2_X1 U1006 ( .A(n1103), .B(n1102), .ZN(n1288) );
NAND2_X1 U1007 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
XNOR2_X1 U1008 ( .A(n1103), .B(n1291), .ZN(n1290) );
INV_X1 U1009 ( .A(n1102), .ZN(n1291) );
XOR2_X1 U1010 ( .A(n1246), .B(n1292), .Z(n1102) );
NOR3_X1 U1011 ( .A1(n1293), .A2(KEYINPUT8), .A3(n1294), .ZN(n1292) );
NOR2_X1 U1012 ( .A1(n1295), .A2(n1229), .ZN(n1293) );
INV_X1 U1013 ( .A(G116), .ZN(n1229) );
XNOR2_X1 U1014 ( .A(G119), .B(KEYINPUT51), .ZN(n1295) );
XNOR2_X1 U1015 ( .A(n1296), .B(n1297), .ZN(n1103) );
NOR2_X1 U1016 ( .A1(KEYINPUT40), .A2(n1261), .ZN(n1297) );
INV_X1 U1017 ( .A(G101), .ZN(n1261) );
XNOR2_X1 U1018 ( .A(G104), .B(G107), .ZN(n1296) );
XNOR2_X1 U1019 ( .A(KEYINPUT42), .B(n1099), .ZN(n1289) );
XOR2_X1 U1020 ( .A(G122), .B(n1255), .Z(n1099) );
NOR2_X1 U1021 ( .A1(n1149), .A2(n1175), .ZN(n1061) );
NOR2_X1 U1022 ( .A1(n1298), .A2(G237), .ZN(n1175) );
XNOR2_X1 U1023 ( .A(KEYINPUT6), .B(n1279), .ZN(n1298) );
INV_X1 U1024 ( .A(G210), .ZN(n1149) );
XOR2_X1 U1025 ( .A(n1299), .B(n1133), .Z(n1205) );
INV_X1 U1026 ( .A(G472), .ZN(n1133) );
NAND2_X1 U1027 ( .A1(KEYINPUT3), .A2(n1065), .ZN(n1299) );
NAND2_X1 U1028 ( .A1(n1300), .A2(n1279), .ZN(n1065) );
XOR2_X1 U1029 ( .A(n1301), .B(n1132), .Z(n1300) );
XNOR2_X1 U1030 ( .A(n1302), .B(G101), .ZN(n1132) );
NAND2_X1 U1031 ( .A1(G210), .A2(n1239), .ZN(n1302) );
NOR2_X1 U1032 ( .A1(G953), .A2(G237), .ZN(n1239) );
XNOR2_X1 U1033 ( .A(KEYINPUT28), .B(n1303), .ZN(n1301) );
NOR2_X1 U1034 ( .A1(KEYINPUT7), .A2(n1129), .ZN(n1303) );
XOR2_X1 U1035 ( .A(n1304), .B(n1305), .Z(n1129) );
XNOR2_X1 U1036 ( .A(n1282), .B(n1246), .ZN(n1305) );
XOR2_X1 U1037 ( .A(G113), .B(KEYINPUT56), .Z(n1246) );
XOR2_X1 U1038 ( .A(n1306), .B(n1235), .Z(n1282) );
XOR2_X1 U1039 ( .A(G143), .B(G146), .Z(n1235) );
NAND2_X1 U1040 ( .A1(KEYINPUT24), .A2(G128), .ZN(n1306) );
XOR2_X1 U1041 ( .A(n1266), .B(n1307), .Z(n1304) );
NOR2_X1 U1042 ( .A1(n1294), .A2(n1308), .ZN(n1307) );
NOR2_X1 U1043 ( .A1(G119), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1044 ( .A(G116), .B(KEYINPUT53), .ZN(n1309) );
NOR2_X1 U1045 ( .A1(n1310), .A2(G116), .ZN(n1294) );
INV_X1 U1046 ( .A(G119), .ZN(n1310) );
XNOR2_X1 U1047 ( .A(G131), .B(n1083), .ZN(n1266) );
XNOR2_X1 U1048 ( .A(G134), .B(n1311), .ZN(n1083) );
XNOR2_X1 U1049 ( .A(n1054), .B(KEYINPUT22), .ZN(n1197) );
XOR2_X1 U1050 ( .A(n1312), .B(n1114), .Z(n1054) );
AND2_X1 U1051 ( .A1(G217), .A2(n1269), .ZN(n1114) );
NAND2_X1 U1052 ( .A1(n1313), .A2(G234), .ZN(n1269) );
XNOR2_X1 U1053 ( .A(KEYINPUT6), .B(G902), .ZN(n1313) );
NAND2_X1 U1054 ( .A1(n1279), .A2(n1111), .ZN(n1312) );
NAND2_X1 U1055 ( .A1(n1314), .A2(n1315), .ZN(n1111) );
NAND3_X1 U1056 ( .A1(n1316), .A2(n1311), .A3(KEYINPUT37), .ZN(n1315) );
XOR2_X1 U1057 ( .A(n1317), .B(n1318), .Z(n1316) );
NOR2_X1 U1058 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NOR2_X1 U1059 ( .A1(KEYINPUT61), .A2(n1321), .ZN(n1320) );
NOR2_X1 U1060 ( .A1(KEYINPUT20), .A2(n1322), .ZN(n1319) );
NAND2_X1 U1061 ( .A1(n1323), .A2(n1324), .ZN(n1314) );
NAND2_X1 U1062 ( .A1(KEYINPUT37), .A2(n1311), .ZN(n1324) );
INV_X1 U1063 ( .A(G137), .ZN(n1311) );
XOR2_X1 U1064 ( .A(n1325), .B(n1317), .Z(n1323) );
XNOR2_X1 U1065 ( .A(n1326), .B(n1236), .ZN(n1317) );
INV_X1 U1066 ( .A(n1082), .ZN(n1236) );
XOR2_X1 U1067 ( .A(G125), .B(G140), .Z(n1082) );
XOR2_X1 U1068 ( .A(n1327), .B(G146), .Z(n1326) );
NAND3_X1 U1069 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1327) );
NAND2_X1 U1070 ( .A1(KEYINPUT14), .A2(n1331), .ZN(n1330) );
NAND3_X1 U1071 ( .A1(n1332), .A2(n1333), .A3(G110), .ZN(n1329) );
NAND2_X1 U1072 ( .A1(n1334), .A2(n1255), .ZN(n1328) );
INV_X1 U1073 ( .A(G110), .ZN(n1255) );
NAND2_X1 U1074 ( .A1(n1335), .A2(n1333), .ZN(n1334) );
INV_X1 U1075 ( .A(KEYINPUT14), .ZN(n1333) );
XNOR2_X1 U1076 ( .A(KEYINPUT1), .B(n1332), .ZN(n1335) );
INV_X1 U1077 ( .A(n1331), .ZN(n1332) );
XOR2_X1 U1078 ( .A(G128), .B(n1336), .Z(n1331) );
NOR2_X1 U1079 ( .A1(KEYINPUT11), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1080 ( .A(G119), .B(KEYINPUT41), .ZN(n1337) );
NAND2_X1 U1081 ( .A1(n1338), .A2(n1339), .ZN(n1325) );
NAND2_X1 U1082 ( .A1(KEYINPUT20), .A2(n1322), .ZN(n1339) );
NAND2_X1 U1083 ( .A1(n1321), .A2(KEYINPUT61), .ZN(n1338) );
INV_X1 U1084 ( .A(n1322), .ZN(n1321) );
NAND2_X1 U1085 ( .A1(G221), .A2(n1222), .ZN(n1322) );
AND2_X1 U1086 ( .A1(G234), .A2(n1104), .ZN(n1222) );
INV_X1 U1087 ( .A(G953), .ZN(n1104) );
INV_X1 U1088 ( .A(G902), .ZN(n1279) );
endmodule


