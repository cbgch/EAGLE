//Key = 00010110100011011000011011111010001101010011000000101110010010001011101010111101100101010110100101111000101100001110001010010011
module c7552 ( G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, 
        G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, 
        G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, 
        G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, 
        G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, 
        G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, 
        G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, 
        G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, 
        G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, 
        G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, 
        G239, G240, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, 
        G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, 
        G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, 
        G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, 
        G4432, G4437, G4526, G4528, G2, G3, G450, G448, G444, G442, G440, G438, 
        G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, 
        G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, 
        G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, 
        G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, 
        G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, 
        G412, G414, G416, G249, G295, G324, G252, G276, G310, G313, G316, G319, 
        G327, G330, G333, G336, G418, G273, G298, G301, G304, G307, G344, G422, 
        G469, G419, G471, G359, G362, G365, G368, G347, G350, G353, G356, G321, 
        G338, G370, G399, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, 
        KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, 
        KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, 
        KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, 
        KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, 
        KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, 
        KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, 
        KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, 
        KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, 
        KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, 
        KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, 
        KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, 
        KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, 
        KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, 
        KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, 
        KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, 
        KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, 
        KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, 
        KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, 
        KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, 
        KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, 
        KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, 
        KEYINPUT125, KEYINPUT126, KEYINPUT127 );

  input G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
         G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
         G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
         G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
         G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133,
         G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
         G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165,
         G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176,
         G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187,
         G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
         G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209,
         G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220,
         G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231,
         G232, G233, G234, G235, G236, G237, G238, G239, G240, G1197, G1455,
         G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211,
         G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701,
         G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394,
         G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528,
         KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
         KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
         KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
         KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
         KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
         KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
         KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
         KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
         KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
         KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
         KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
         KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
         KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65, KEYINPUT66,
         KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
         KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
         KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
         KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
         KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91,
         KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96,
         KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100, KEYINPUT101,
         KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105, KEYINPUT106,
         KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110, KEYINPUT111,
         KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115, KEYINPUT116,
         KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120, KEYINPUT121,
         KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125, KEYINPUT126,
         KEYINPUT127;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
         G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552,
         G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528,
         G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410,
         G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373,
         G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382,
         G385, G412, G414, G416, G249, G295, G324, G252, G276, G310, G313,
         G316, G319, G327, G330, G333, G336, G418, G273, G298, G301, G304,
         G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, G347,
         G350, G353, G356, G321, G338, G370, G399;

  wire   n4463, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947;

  INV_X4 U3097 ( .A(G18), .ZN(n4527) );
  INV_X1 U3098 ( .A(G1), .ZN(n4463) );
  INV_X1 U3099 ( .A(n4463), .ZN(G2) );
  INV_X1 U3100 ( .A(n4463), .ZN(G3) );
  INV_X1 U3101 ( .A(n4463), .ZN(G453) );
  INV_X1 U3102 ( .A(n4463), .ZN(G432) );
  BUF_X1 U3103 ( .A(G106), .Z(G446) );
  BUF_X1 U3104 ( .A(G1459), .Z(G450) );
  BUF_X1 U3105 ( .A(G1462), .Z(G436) );
  BUF_X1 U3106 ( .A(G1469), .Z(G448) );
  BUF_X1 U3107 ( .A(G1480), .Z(G444) );
  BUF_X1 U3108 ( .A(G1486), .Z(G442) );
  BUF_X1 U3109 ( .A(G1496), .Z(G438) );
  BUF_X1 U3110 ( .A(G2208), .Z(G496) );
  BUF_X1 U3111 ( .A(G2211), .Z(G478) );
  BUF_X1 U3112 ( .A(G2218), .Z(G494) );
  BUF_X1 U3113 ( .A(G2224), .Z(G492) );
  BUF_X1 U3114 ( .A(G2230), .Z(G490) );
  BUF_X1 U3115 ( .A(G2236), .Z(G488) );
  BUF_X1 U3116 ( .A(G2239), .Z(G486) );
  BUF_X1 U3117 ( .A(G2247), .Z(G484) );
  BUF_X1 U3118 ( .A(G2253), .Z(G482) );
  BUF_X1 U3119 ( .A(G2256), .Z(G480) );
  BUF_X1 U3120 ( .A(G3698), .Z(G560) );
  BUF_X1 U3121 ( .A(G3701), .Z(G542) );
  BUF_X1 U3122 ( .A(G3705), .Z(G558) );
  BUF_X1 U3123 ( .A(G3711), .Z(G556) );
  BUF_X1 U3124 ( .A(G3717), .Z(G554) );
  BUF_X1 U3125 ( .A(G3723), .Z(G552) );
  BUF_X1 U3126 ( .A(G3729), .Z(G550) );
  BUF_X1 U3127 ( .A(G3737), .Z(G548) );
  BUF_X1 U3128 ( .A(G3743), .Z(G546) );
  BUF_X1 U3129 ( .A(G3749), .Z(G544) );
  BUF_X1 U3130 ( .A(G4393), .Z(G540) );
  BUF_X1 U3131 ( .A(G4394), .Z(G522) );
  BUF_X1 U3132 ( .A(G4400), .Z(G538) );
  BUF_X1 U3133 ( .A(G4405), .Z(G536) );
  BUF_X1 U3134 ( .A(G4410), .Z(G534) );
  BUF_X1 U3135 ( .A(G4415), .Z(G532) );
  BUF_X1 U3136 ( .A(G4420), .Z(G530) );
  BUF_X1 U3137 ( .A(G4432), .Z(G526) );
  BUF_X1 U3138 ( .A(G4437), .Z(G524) );
  BUF_X1 U3139 ( .A(G341), .Z(G279) );
  BUF_X1 U3140 ( .A(G289), .Z(G284) );
  BUF_X1 U3141 ( .A(G264), .Z(G258) );
  BUF_X1 U3142 ( .A(G469), .Z(G422) );
  BUF_X1 U3143 ( .A(G471), .Z(G419) );
  BUF_X1 U3144 ( .A(G292), .Z(G281) );
  XNOR2_X1 U3145 ( .A(KEYINPUT40), .B(n4510), .ZN(G528) );
  XNOR2_X1 U3146 ( .A(n4511), .B(n4512), .ZN(G471) );
  XNOR2_X1 U3147 ( .A(n4513), .B(n4514), .ZN(G469) );
  NAND2_X1 U3148 ( .A1(n4515), .A2(n4516), .ZN(n4513) );
  NAND2_X1 U3149 ( .A1(n4517), .A2(n4512), .ZN(n4516) );
  NAND2_X1 U3150 ( .A1(KEYINPUT52), .A2(n4518), .ZN(n4517) );
  XNOR2_X1 U3151 ( .A(G1492), .B(KEYINPUT25), .ZN(G440) );
  OR4_X1 U3152 ( .A1(G406), .A2(G408), .A3(G404), .A4(n4519), .ZN(G418) );
  OR4_X1 U3153 ( .A1(G416), .A2(G414), .A3(G412), .A4(G410), .ZN(n4519) );
  NAND3_X1 U3154 ( .A1(n4520), .A2(n4521), .A3(n4522), .ZN(G416) );
  NOR3_X1 U3155 ( .A1(n4523), .A2(n4524), .A3(n4525), .ZN(n4522) );
  NOR3_X1 U3156 ( .A1(n4526), .A2(G165), .A3(n4527), .ZN(n4525) );
  NOR2_X1 U3157 ( .A1(n4528), .A2(n4529), .ZN(n4524) );
  INV_X1 U3158 ( .A(n4526), .ZN(n4529) );
  XNOR2_X1 U3159 ( .A(n4530), .B(n4531), .ZN(n4526) );
  XNOR2_X1 U3160 ( .A(n4532), .B(n4533), .ZN(n4531) );
  XNOR2_X1 U3161 ( .A(n4534), .B(n4535), .ZN(n4533) );
  NOR2_X1 U3162 ( .A1(G170), .A2(n4536), .ZN(n4534) );
  XOR2_X1 U3163 ( .A(n4537), .B(n4538), .Z(n4530) );
  XOR2_X1 U3164 ( .A(n4539), .B(n4540), .Z(n4538) );
  NAND2_X1 U3165 ( .A1(n4541), .A2(n4542), .ZN(n4537) );
  NAND2_X1 U3166 ( .A1(G164), .A2(n4543), .ZN(n4542) );
  NOR2_X1 U3167 ( .A1(n4544), .A2(n4545), .ZN(n4528) );
  AND2_X1 U3168 ( .A1(n4543), .A2(G165), .ZN(n4544) );
  XOR2_X1 U3169 ( .A(n4546), .B(n4547), .Z(n4523) );
  XOR2_X1 U3170 ( .A(n4548), .B(n4549), .Z(n4547) );
  XNOR2_X1 U3171 ( .A(n4550), .B(n4551), .ZN(n4549) );
  XOR2_X1 U3172 ( .A(n4552), .B(n4553), .Z(n4551) );
  XOR2_X1 U3173 ( .A(n4554), .B(n4555), .Z(n4553) );
  NOR2_X1 U3174 ( .A1(n4556), .A2(n4557), .ZN(n4552) );
  NOR2_X1 U3175 ( .A1(G18), .A2(G141), .ZN(n4557) );
  NOR2_X1 U3176 ( .A1(G181), .A2(n4527), .ZN(n4556) );
  XOR2_X1 U3177 ( .A(n4558), .B(n4559), .Z(n4548) );
  XOR2_X1 U3178 ( .A(n4560), .B(n4561), .Z(n4546) );
  XNOR2_X1 U3179 ( .A(n4562), .B(n4563), .ZN(n4561) );
  NAND2_X1 U3180 ( .A1(n4564), .A2(n4565), .ZN(n4562) );
  OR2_X1 U3181 ( .A1(n4566), .A2(n4567), .ZN(n4565) );
  XOR2_X1 U3182 ( .A(n4568), .B(KEYINPUT41), .Z(n4564) );
  NAND2_X1 U3183 ( .A1(n4567), .A2(n4566), .ZN(n4568) );
  XOR2_X1 U3184 ( .A(n4569), .B(KEYINPUT56), .Z(n4560) );
  NAND2_X1 U3185 ( .A1(KEYINPUT72), .A2(n4570), .ZN(n4569) );
  INV_X1 U3186 ( .A(n4571), .ZN(n4570) );
  XOR2_X1 U3187 ( .A(n4572), .B(n4573), .Z(n4521) );
  XOR2_X1 U3188 ( .A(n4574), .B(n4575), .Z(n4573) );
  XOR2_X1 U3189 ( .A(n4576), .B(n4577), .Z(n4575) );
  XNOR2_X1 U3190 ( .A(n4578), .B(n4579), .ZN(n4577) );
  NAND2_X1 U3191 ( .A1(n4580), .A2(n4581), .ZN(n4578) );
  NAND2_X1 U3192 ( .A1(n4582), .A2(n4583), .ZN(n4581) );
  XNOR2_X1 U3193 ( .A(G115), .B(n4584), .ZN(n4582) );
  NAND2_X1 U3194 ( .A1(n4585), .A2(n4586), .ZN(n4580) );
  XNOR2_X1 U3195 ( .A(G197), .B(n4584), .ZN(n4585) );
  XNOR2_X1 U3196 ( .A(n4587), .B(n4588), .ZN(n4576) );
  NAND2_X1 U3197 ( .A1(KEYINPUT13), .A2(n4589), .ZN(n4587) );
  INV_X1 U3198 ( .A(n4590), .ZN(n4589) );
  XOR2_X1 U3199 ( .A(n4591), .B(n4592), .Z(n4574) );
  XOR2_X1 U3200 ( .A(n4593), .B(n4594), .Z(n4592) );
  XNOR2_X1 U3201 ( .A(n4595), .B(n4596), .ZN(n4591) );
  XNOR2_X1 U3202 ( .A(n4597), .B(n4598), .ZN(n4520) );
  XOR2_X1 U3203 ( .A(n4599), .B(n4600), .Z(n4597) );
  XOR2_X1 U3204 ( .A(n4601), .B(n4602), .Z(n4600) );
  XOR2_X1 U3205 ( .A(n4603), .B(n4604), .Z(n4602) );
  NOR2_X1 U3206 ( .A1(n4605), .A2(n4606), .ZN(n4604) );
  XOR2_X1 U3207 ( .A(KEYINPUT11), .B(n4607), .Z(n4606) );
  NOR2_X1 U3208 ( .A1(n4608), .A2(n4609), .ZN(n4607) );
  AND2_X1 U3209 ( .A1(n4609), .A2(n4608), .ZN(n4605) );
  XOR2_X1 U3210 ( .A(n4610), .B(KEYINPUT43), .Z(n4601) );
  NAND3_X1 U3211 ( .A1(n4611), .A2(n4612), .A3(n4613), .ZN(n4610) );
  NAND2_X1 U3212 ( .A1(n4614), .A2(G18), .ZN(n4613) );
  XNOR2_X1 U3213 ( .A(G208), .B(n4615), .ZN(n4614) );
  OR3_X1 U3214 ( .A1(n4615), .A2(G18), .A3(G44), .ZN(n4612) );
  NAND2_X1 U3215 ( .A1(G44), .A2(n4616), .ZN(n4611) );
  XOR2_X1 U3216 ( .A(n4617), .B(n4618), .Z(n4599) );
  XNOR2_X1 U3217 ( .A(n4619), .B(n4620), .ZN(n4618) );
  XNOR2_X1 U3218 ( .A(n4621), .B(n4622), .ZN(n4617) );
  NAND4_X1 U3219 ( .A1(n4623), .A2(n4624), .A3(n4625), .A4(n4626), .ZN(G414) );
  NAND2_X1 U3220 ( .A1(G18), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U3221 ( .A1(n4628), .A2(n4629), .ZN(n4627) );
  XNOR2_X1 U3222 ( .A(n4630), .B(n4631), .ZN(n4629) );
  XNOR2_X1 U3223 ( .A(G1492), .B(n4632), .ZN(n4628) );
  NAND2_X1 U3224 ( .A1(n4633), .A2(n4527), .ZN(n4625) );
  NAND2_X1 U3225 ( .A1(n4634), .A2(n4635), .ZN(n4633) );
  XNOR2_X1 U3226 ( .A(G70), .B(n4631), .ZN(n4635) );
  XNOR2_X1 U3227 ( .A(n4636), .B(n4637), .ZN(n4631) );
  XOR2_X1 U3228 ( .A(n4638), .B(n4639), .Z(n4637) );
  XOR2_X1 U3229 ( .A(n4640), .B(n4641), .Z(n4638) );
  XOR2_X1 U3230 ( .A(n4642), .B(n4643), .Z(n4641) );
  XOR2_X1 U3231 ( .A(n4644), .B(n4645), .Z(n4643) );
  XNOR2_X1 U3232 ( .A(n4646), .B(n4647), .ZN(n4642) );
  XOR2_X1 U3233 ( .A(n4648), .B(n4649), .Z(n4640) );
  XOR2_X1 U3234 ( .A(n4650), .B(n4651), .Z(n4649) );
  XOR2_X1 U3235 ( .A(n4652), .B(KEYINPUT120), .Z(n4648) );
  NAND2_X1 U3236 ( .A1(n4653), .A2(n4654), .ZN(n4636) );
  OR2_X1 U3237 ( .A1(G3698), .A2(n4527), .ZN(n4654) );
  NAND2_X1 U3238 ( .A1(G69), .A2(n4527), .ZN(n4653) );
  XOR2_X1 U3239 ( .A(n4632), .B(G1455), .Z(n4634) );
  NAND2_X1 U3240 ( .A1(n4655), .A2(n4656), .ZN(n4632) );
  NAND2_X1 U3241 ( .A1(n4657), .A2(n4527), .ZN(n4656) );
  XNOR2_X1 U3242 ( .A(G2204), .B(n4658), .ZN(n4657) );
  NAND2_X1 U3243 ( .A1(n4659), .A2(G18), .ZN(n4655) );
  XOR2_X1 U3244 ( .A(G1496), .B(n4658), .Z(n4659) );
  XNOR2_X1 U3245 ( .A(n4660), .B(n4661), .ZN(n4658) );
  XOR2_X1 U3246 ( .A(n4662), .B(n4663), .Z(n4661) );
  NAND2_X1 U3247 ( .A1(n4664), .A2(n4665), .ZN(n4660) );
  NAND2_X1 U3248 ( .A1(n4666), .A2(n4667), .ZN(n4665) );
  NAND2_X1 U3249 ( .A1(KEYINPUT39), .A2(n4668), .ZN(n4667) );
  INV_X1 U3250 ( .A(n4669), .ZN(n4666) );
  NAND2_X1 U3251 ( .A1(n4668), .A2(n4669), .ZN(n4664) );
  NAND2_X1 U3252 ( .A1(n4670), .A2(n4671), .ZN(n4669) );
  NAND2_X1 U3253 ( .A1(n4672), .A2(n4673), .ZN(n4671) );
  XOR2_X1 U3254 ( .A(KEYINPUT114), .B(n4674), .Z(n4670) );
  NOR2_X1 U3255 ( .A1(n4672), .A2(n4673), .ZN(n4674) );
  INV_X1 U3256 ( .A(n4675), .ZN(n4672) );
  NAND2_X1 U3257 ( .A1(n4676), .A2(n4677), .ZN(n4668) );
  NAND2_X1 U3258 ( .A1(n4678), .A2(n4527), .ZN(n4677) );
  XNOR2_X1 U3259 ( .A(G114), .B(n4679), .ZN(n4678) );
  NAND2_X1 U3260 ( .A1(n4680), .A2(G18), .ZN(n4676) );
  XOR2_X1 U3261 ( .A(n4679), .B(G1459), .Z(n4680) );
  XOR2_X1 U3262 ( .A(n4681), .B(n4682), .Z(n4624) );
  XNOR2_X1 U3263 ( .A(n4683), .B(n4684), .ZN(n4682) );
  NOR2_X1 U3264 ( .A1(KEYINPUT84), .A2(n4685), .ZN(n4684) );
  XNOR2_X1 U3265 ( .A(n4686), .B(n4687), .ZN(n4685) );
  XOR2_X1 U3266 ( .A(n4688), .B(KEYINPUT48), .Z(n4686) );
  NAND3_X1 U3267 ( .A1(n4689), .A2(n4690), .A3(KEYINPUT66), .ZN(n4683) );
  NAND2_X1 U3268 ( .A1(n4691), .A2(n4527), .ZN(n4690) );
  XOR2_X1 U3269 ( .A(G82), .B(n4692), .Z(n4691) );
  NAND2_X1 U3270 ( .A1(n4693), .A2(G18), .ZN(n4689) );
  XNOR2_X1 U3271 ( .A(n4692), .B(G2208), .ZN(n4693) );
  XNOR2_X1 U3272 ( .A(n4694), .B(n4695), .ZN(n4692) );
  NOR2_X1 U3273 ( .A1(n4696), .A2(n4697), .ZN(n4695) );
  AND2_X1 U3274 ( .A1(n4698), .A2(n4699), .ZN(n4697) );
  NOR3_X1 U3275 ( .A1(n4698), .A2(KEYINPUT124), .A3(n4699), .ZN(n4696) );
  XOR2_X1 U3276 ( .A(n4700), .B(n4701), .Z(n4699) );
  XOR2_X1 U3277 ( .A(n4702), .B(n4703), .Z(n4698) );
  XOR2_X1 U3278 ( .A(n4704), .B(n4705), .Z(n4681) );
  XOR2_X1 U3279 ( .A(n4706), .B(n4707), .Z(n4623) );
  NOR4_X1 U3280 ( .A1(n4708), .A2(n4709), .A3(n4710), .A4(n4711), .ZN(n4707) );
  NOR3_X1 U3281 ( .A1(n4712), .A2(n4713), .A3(n4714), .ZN(n4711) );
  AND3_X1 U3282 ( .A1(n4712), .A2(n4715), .A3(n4713), .ZN(n4710) );
  NOR3_X1 U3283 ( .A1(n4713), .A2(n4716), .A3(n4715), .ZN(n4709) );
  INV_X1 U3284 ( .A(n4714), .ZN(n4715) );
  AND3_X1 U3285 ( .A1(n4713), .A2(n4714), .A3(n4716), .ZN(n4708) );
  XNOR2_X1 U3286 ( .A(n4712), .B(KEYINPUT62), .ZN(n4716) );
  XNOR2_X1 U3287 ( .A(n4717), .B(n4718), .ZN(n4712) );
  XNOR2_X1 U3288 ( .A(n4719), .B(n4720), .ZN(n4714) );
  NAND2_X1 U3289 ( .A1(n4721), .A2(n4722), .ZN(n4713) );
  NAND2_X1 U3290 ( .A1(n4723), .A2(n4527), .ZN(n4722) );
  XNOR2_X1 U3291 ( .A(G58), .B(n4724), .ZN(n4723) );
  NAND2_X1 U3292 ( .A1(n4725), .A2(G18), .ZN(n4721) );
  XOR2_X1 U3293 ( .A(n4724), .B(G4393), .Z(n4725) );
  NAND2_X1 U3294 ( .A1(KEYINPUT67), .A2(n4726), .ZN(n4706) );
  XOR2_X1 U3295 ( .A(n4727), .B(n4728), .Z(n4726) );
  XOR2_X1 U3296 ( .A(n4729), .B(n4730), .Z(n4728) );
  XOR2_X1 U3297 ( .A(n4731), .B(n4732), .Z(n4727) );
  NAND3_X1 U3298 ( .A1(n4733), .A2(n4734), .A3(n4735), .ZN(G412) );
  NOR3_X1 U3299 ( .A1(n4736), .A2(n4737), .A3(n4738), .ZN(n4735) );
  AND3_X1 U3300 ( .A1(G212), .A2(n4543), .A3(n4739), .ZN(n4738) );
  NOR3_X1 U3301 ( .A1(G212), .A2(n4739), .A3(n4527), .ZN(n4737) );
  XNOR2_X1 U3302 ( .A(n4740), .B(n4741), .ZN(n4739) );
  XOR2_X1 U3303 ( .A(n4742), .B(n4743), .Z(n4741) );
  XNOR2_X1 U3304 ( .A(n4744), .B(n4745), .ZN(n4743) );
  NOR3_X1 U3305 ( .A1(n4545), .A2(G209), .A3(n4746), .ZN(n4742) );
  XNOR2_X1 U3306 ( .A(n4747), .B(n4748), .ZN(n4740) );
  XOR2_X1 U3307 ( .A(n4749), .B(n4750), .Z(n4747) );
  NOR2_X1 U3308 ( .A1(n4545), .A2(n4751), .ZN(n4750) );
  NOR2_X1 U3309 ( .A1(n4746), .A2(n4752), .ZN(n4751) );
  XNOR2_X1 U3310 ( .A(KEYINPUT7), .B(G211), .ZN(n4752) );
  XOR2_X1 U3311 ( .A(n4753), .B(n4754), .Z(n4736) );
  XOR2_X1 U3312 ( .A(n4755), .B(n4756), .Z(n4754) );
  XOR2_X1 U3313 ( .A(n4757), .B(n4758), .Z(n4756) );
  NAND2_X1 U3314 ( .A1(n4759), .A2(n4760), .ZN(n4755) );
  NAND2_X1 U3315 ( .A1(n4761), .A2(n4527), .ZN(n4760) );
  XOR2_X1 U3316 ( .A(G115), .B(n4762), .Z(n4761) );
  NAND2_X1 U3317 ( .A1(n4763), .A2(G18), .ZN(n4759) );
  XOR2_X1 U3318 ( .A(G227), .B(n4762), .Z(n4763) );
  XNOR2_X1 U3319 ( .A(n4764), .B(n4765), .ZN(n4762) );
  XOR2_X1 U3320 ( .A(n4766), .B(n4767), .Z(n4753) );
  XOR2_X1 U3321 ( .A(n4768), .B(n4769), .Z(n4767) );
  XNOR2_X1 U3322 ( .A(n4770), .B(n4771), .ZN(n4766) );
  NAND4_X1 U3323 ( .A1(n4772), .A2(n4773), .A3(n4774), .A4(n4775), .ZN(n4770) );
  NAND3_X1 U3324 ( .A1(n4776), .A2(n4777), .A3(n4778), .ZN(n4775) );
  INV_X1 U3325 ( .A(KEYINPUT44), .ZN(n4778) );
  NAND2_X1 U3326 ( .A1(KEYINPUT126), .A2(n4779), .ZN(n4777) );
  NAND3_X1 U3327 ( .A1(n4780), .A2(n4781), .A3(KEYINPUT44), .ZN(n4774) );
  OR2_X1 U3328 ( .A1(n4782), .A2(KEYINPUT126), .ZN(n4781) );
  OR2_X1 U3329 ( .A1(n4779), .A2(KEYINPUT85), .ZN(n4773) );
  NAND3_X1 U3330 ( .A1(n4783), .A2(n4779), .A3(KEYINPUT85), .ZN(n4772) );
  XNOR2_X1 U3331 ( .A(KEYINPUT126), .B(n4780), .ZN(n4783) );
  XOR2_X1 U3332 ( .A(n4784), .B(n4785), .Z(n4734) );
  XNOR2_X1 U3333 ( .A(n4786), .B(n4787), .ZN(n4785) );
  XNOR2_X1 U3334 ( .A(n4788), .B(n4789), .ZN(n4784) );
  XNOR2_X1 U3335 ( .A(n4790), .B(n4791), .ZN(n4789) );
  NOR3_X1 U3336 ( .A1(KEYINPUT55), .A2(n4792), .A3(n4793), .ZN(n4791) );
  NOR2_X1 U3337 ( .A1(n4527), .A2(n4794), .ZN(n4793) );
  XOR2_X1 U3338 ( .A(n4795), .B(G239), .Z(n4794) );
  NOR2_X1 U3339 ( .A1(G18), .A2(n4796), .ZN(n4792) );
  XOR2_X1 U3340 ( .A(n4795), .B(G44), .Z(n4796) );
  XNOR2_X1 U3341 ( .A(n4797), .B(n4798), .ZN(n4795) );
  NAND2_X1 U3342 ( .A1(n4799), .A2(n4800), .ZN(n4797) );
  NAND2_X1 U3343 ( .A1(n4801), .A2(n4802), .ZN(n4800) );
  NAND2_X1 U3344 ( .A1(n4803), .A2(KEYINPUT12), .ZN(n4802) );
  XNOR2_X1 U3345 ( .A(n4804), .B(n4805), .ZN(n4801) );
  NAND2_X1 U3346 ( .A1(n4803), .A2(n4806), .ZN(n4799) );
  XNOR2_X1 U3347 ( .A(n4807), .B(n4804), .ZN(n4806) );
  XNOR2_X1 U3348 ( .A(n4808), .B(n4809), .ZN(n4803) );
  XOR2_X1 U3349 ( .A(n4810), .B(n4811), .Z(n4733) );
  XOR2_X1 U3350 ( .A(n4812), .B(n4813), .Z(n4811) );
  XNOR2_X1 U3351 ( .A(n4814), .B(n4815), .ZN(n4813) );
  NAND2_X1 U3352 ( .A1(n4816), .A2(n4817), .ZN(n4812) );
  NAND2_X1 U3353 ( .A1(n4818), .A2(n4527), .ZN(n4817) );
  XOR2_X1 U3354 ( .A(n4819), .B(G141), .Z(n4818) );
  NAND2_X1 U3355 ( .A1(n4820), .A2(G18), .ZN(n4816) );
  XOR2_X1 U3356 ( .A(n4819), .B(G161), .Z(n4820) );
  XNOR2_X1 U3357 ( .A(n4821), .B(n4822), .ZN(n4819) );
  XOR2_X1 U3358 ( .A(n4823), .B(n4824), .Z(n4810) );
  XNOR2_X1 U3359 ( .A(n4825), .B(n4826), .ZN(n4824) );
  NOR2_X1 U3360 ( .A1(KEYINPUT49), .A2(n4827), .ZN(n4826) );
  XOR2_X1 U3361 ( .A(n4828), .B(n4829), .Z(n4827) );
  NAND2_X1 U3362 ( .A1(KEYINPUT34), .A2(n4830), .ZN(n4828) );
  XNOR2_X1 U3363 ( .A(n4831), .B(n4832), .ZN(n4823) );
  NAND4_X1 U3364 ( .A1(G199), .A2(G188), .A3(G172), .A4(G162), .ZN(G410) );
  NAND4_X1 U3365 ( .A1(G186), .A2(G185), .A3(G183), .A4(G182), .ZN(G408) );
  NAND4_X1 U3366 ( .A1(G230), .A2(G218), .A3(G210), .A4(G152), .ZN(G406) );
  NAND4_X1 U3367 ( .A1(G240), .A2(G228), .A3(G184), .A4(G150), .ZN(G404) );
  OR2_X1 U3368 ( .A1(G5), .A2(G57), .ZN(G402) );
  XOR2_X1 U3369 ( .A(n4833), .B(n4834), .Z(G399) );
  NOR2_X1 U3370 ( .A1(n4835), .A2(n4836), .ZN(n4834) );
  NOR2_X1 U3371 ( .A1(G4526), .A2(n4837), .ZN(n4836) );
  NOR2_X1 U3372 ( .A1(n4838), .A2(n4839), .ZN(n4837) );
  AND2_X1 U3373 ( .A1(n4840), .A2(n4841), .ZN(n4839) );
  NOR2_X1 U3374 ( .A1(n4841), .A2(n4842), .ZN(n4838) );
  INV_X1 U3375 ( .A(n4843), .ZN(n4842) );
  NOR2_X1 U3376 ( .A1(KEYINPUT2), .A2(n4844), .ZN(n4841) );
  XOR2_X1 U3377 ( .A(n4845), .B(n4846), .Z(n4844) );
  XOR2_X1 U3378 ( .A(n4847), .B(n4848), .Z(n4845) );
  NOR2_X1 U3379 ( .A1(n4849), .A2(n4850), .ZN(n4848) );
  XNOR2_X1 U3380 ( .A(n4851), .B(n4852), .ZN(n4850) );
  NOR2_X1 U3381 ( .A1(n4853), .A2(n4854), .ZN(n4852) );
  NOR2_X1 U3382 ( .A1(n4855), .A2(n4856), .ZN(n4835) );
  XOR2_X1 U3383 ( .A(n4857), .B(n4858), .Z(n4856) );
  XOR2_X1 U3384 ( .A(n4859), .B(n4860), .Z(n4858) );
  NAND2_X1 U3385 ( .A1(KEYINPUT26), .A2(n4861), .ZN(n4860) );
  NAND4_X1 U3386 ( .A1(n4862), .A2(n4863), .A3(n4864), .A4(n4865), .ZN(n4859) );
  NOR2_X1 U3387 ( .A1(n4854), .A2(n4849), .ZN(n4865) );
  NOR3_X1 U3388 ( .A1(n4851), .A2(n4866), .A3(n4867), .ZN(n4849) );
  NAND2_X1 U3389 ( .A1(n4853), .A2(n4868), .ZN(n4864) );
  INV_X1 U3390 ( .A(KEYINPUT47), .ZN(n4868) );
  NOR2_X1 U3391 ( .A1(n4869), .A2(n4866), .ZN(n4853) );
  NAND3_X1 U3392 ( .A1(KEYINPUT47), .A2(n4870), .A3(n4866), .ZN(n4863) );
  NAND2_X1 U3393 ( .A1(n4871), .A2(n4872), .ZN(n4862) );
  XOR2_X1 U3394 ( .A(n4873), .B(n4847), .Z(n4857) );
  NAND3_X1 U3395 ( .A1(n4874), .A2(n4875), .A3(n4876), .ZN(n4847) );
  NAND2_X1 U3396 ( .A1(n4877), .A2(n4878), .ZN(n4876) );
  XNOR2_X1 U3397 ( .A(n4879), .B(n4880), .ZN(n4877) );
  NAND2_X1 U3398 ( .A1(n4881), .A2(n4871), .ZN(n4875) );
  NAND3_X1 U3399 ( .A1(n4882), .A2(n4867), .A3(n4880), .ZN(n4874) );
  NAND2_X1 U3400 ( .A1(n4883), .A2(n4884), .ZN(n4873) );
  NAND3_X1 U3401 ( .A1(n4885), .A2(n4886), .A3(n4843), .ZN(n4884) );
  NAND2_X1 U3402 ( .A1(n4887), .A2(n4888), .ZN(n4843) );
  NAND2_X1 U3403 ( .A1(n4889), .A2(n4866), .ZN(n4888) );
  NAND2_X1 U3404 ( .A1(n4871), .A2(n4890), .ZN(n4886) );
  NAND2_X1 U3405 ( .A1(n4891), .A2(n4887), .ZN(n4890) );
  INV_X1 U3406 ( .A(n4892), .ZN(n4887) );
  OR2_X1 U3407 ( .A1(n4846), .A2(n4871), .ZN(n4885) );
  XOR2_X1 U3408 ( .A(n4893), .B(n4894), .Z(n4846) );
  NAND2_X1 U3409 ( .A1(n4840), .A2(n4895), .ZN(n4883) );
  NAND3_X1 U3410 ( .A1(n4896), .A2(n4897), .A3(n4898), .ZN(n4895) );
  NAND2_X1 U3411 ( .A1(n4871), .A2(n4894), .ZN(n4898) );
  OR3_X1 U3412 ( .A1(n4893), .A2(n4871), .A3(n4894), .ZN(n4897) );
  NAND2_X1 U3413 ( .A1(n4893), .A2(n4894), .ZN(n4896) );
  INV_X1 U3414 ( .A(n4891), .ZN(n4894) );
  NOR2_X1 U3415 ( .A1(n4899), .A2(n4900), .ZN(n4891) );
  AND2_X1 U3416 ( .A1(n4892), .A2(n4893), .ZN(n4900) );
  NAND2_X1 U3417 ( .A1(n4869), .A2(n4901), .ZN(n4893) );
  NAND2_X1 U3418 ( .A1(n4879), .A2(n4902), .ZN(n4901) );
  XNOR2_X1 U3419 ( .A(n4872), .B(n4889), .ZN(n4840) );
  NAND2_X1 U3420 ( .A1(n4903), .A2(n4904), .ZN(n4833) );
  NAND2_X1 U3421 ( .A1(n4905), .A2(n4906), .ZN(n4904) );
  XOR2_X1 U3422 ( .A(n4907), .B(n4908), .Z(n4905) );
  XNOR2_X1 U3423 ( .A(n4909), .B(n4910), .ZN(n4908) );
  NAND3_X1 U3424 ( .A1(n4911), .A2(n4912), .A3(n4913), .ZN(n4909) );
  NAND2_X1 U3425 ( .A1(n4914), .A2(n4915), .ZN(n4913) );
  XNOR2_X1 U3426 ( .A(n4916), .B(n4917), .ZN(n4914) );
  OR3_X1 U3427 ( .A1(n4917), .A2(n4915), .A3(n4918), .ZN(n4912) );
  OR2_X1 U3428 ( .A1(n4919), .A2(n4916), .ZN(n4911) );
  XNOR2_X1 U3429 ( .A(n4920), .B(n4921), .ZN(n4907) );
  XNOR2_X1 U3430 ( .A(n4922), .B(n4923), .ZN(n4921) );
  NOR2_X1 U3431 ( .A1(KEYINPUT61), .A2(n4924), .ZN(n4922) );
  XNOR2_X1 U3432 ( .A(n4925), .B(KEYINPUT1), .ZN(n4924) );
  NAND2_X1 U3433 ( .A1(n4926), .A2(n4927), .ZN(n4903) );
  NAND3_X1 U3434 ( .A1(n4928), .A2(n4929), .A3(n4930), .ZN(n4927) );
  NAND2_X1 U3435 ( .A1(n4931), .A2(n4855), .ZN(n4929) );
  INV_X1 U3436 ( .A(G4526), .ZN(n4855) );
  NAND2_X1 U3437 ( .A1(n4932), .A2(G4526), .ZN(n4928) );
  XOR2_X1 U3438 ( .A(n4933), .B(n4934), .Z(n4926) );
  XOR2_X1 U3439 ( .A(n4935), .B(n4936), .Z(n4934) );
  NAND2_X1 U3440 ( .A1(n4937), .A2(n4938), .ZN(n4936) );
  NAND2_X1 U3441 ( .A1(n4920), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U3442 ( .A1(n4940), .A2(n4941), .ZN(n4937) );
  NAND2_X1 U3443 ( .A1(n4942), .A2(n4939), .ZN(n4941) );
  INV_X1 U3444 ( .A(n4920), .ZN(n4940) );
  NAND2_X1 U3445 ( .A1(n4943), .A2(n4944), .ZN(n4935) );
  NAND2_X1 U3446 ( .A1(n4917), .A2(n4923), .ZN(n4944) );
  OR3_X1 U3447 ( .A1(n4917), .A2(n4945), .A3(n4923), .ZN(n4943) );
  XNOR2_X1 U3448 ( .A(n4946), .B(n4942), .ZN(n4933) );
  XNOR2_X1 U3449 ( .A(n4947), .B(n4925), .ZN(n4946) );
  XNOR2_X1 U3450 ( .A(n4948), .B(n4949), .ZN(G397) );
  NAND2_X1 U3451 ( .A1(KEYINPUT42), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U3452 ( .A1(n4951), .A2(n4851), .ZN(n4950) );
  NAND2_X1 U3453 ( .A1(G4526), .A2(n4882), .ZN(n4951) );
  XNOR2_X1 U3454 ( .A(n4952), .B(n4866), .ZN(G394) );
  XNOR2_X1 U3455 ( .A(n4953), .B(n4889), .ZN(G391) );
  NAND2_X1 U3456 ( .A1(n4954), .A2(n4955), .ZN(n4953) );
  NAND2_X1 U3457 ( .A1(n4872), .A2(n4952), .ZN(n4955) );
  INV_X1 U3458 ( .A(n4866), .ZN(n4872) );
  XNOR2_X1 U3459 ( .A(n4956), .B(n4880), .ZN(G388) );
  NAND3_X1 U3460 ( .A1(n4957), .A2(n4958), .A3(n4959), .ZN(n4956) );
  NAND2_X1 U3461 ( .A1(n4960), .A2(n4961), .ZN(n4958) );
  XNOR2_X1 U3462 ( .A(KEYINPUT111), .B(n4954), .ZN(n4961) );
  NAND2_X1 U3463 ( .A1(n4892), .A2(n4952), .ZN(n4957) );
  NAND3_X1 U3464 ( .A1(n4869), .A2(n4962), .A3(n4963), .ZN(n4952) );
  NAND2_X1 U3465 ( .A1(n4902), .A2(n4948), .ZN(n4963) );
  XNOR2_X1 U3466 ( .A(n4964), .B(n4965), .ZN(G385) );
  NAND2_X1 U3467 ( .A1(KEYINPUT107), .A2(n4966), .ZN(n4965) );
  XNOR2_X1 U3468 ( .A(n4967), .B(n4968), .ZN(G382) );
  NOR2_X1 U3469 ( .A1(n4916), .A2(n4969), .ZN(n4967) );
  AND2_X1 U3470 ( .A1(n4939), .A2(n4966), .ZN(n4969) );
  XNOR2_X1 U3471 ( .A(n4970), .B(n4925), .ZN(G379) );
  NAND2_X1 U3472 ( .A1(n4971), .A2(n4972), .ZN(n4970) );
  NAND2_X1 U3473 ( .A1(KEYINPUT123), .A2(n4973), .ZN(n4972) );
  NAND2_X1 U3474 ( .A1(n4974), .A2(n4975), .ZN(n4973) );
  NAND3_X1 U3475 ( .A1(n4968), .A2(n4966), .A3(n4964), .ZN(n4975) );
  INV_X1 U3476 ( .A(n4976), .ZN(n4974) );
  NAND2_X1 U3477 ( .A1(n4977), .A2(n4976), .ZN(n4971) );
  NAND2_X1 U3478 ( .A1(n4978), .A2(n4979), .ZN(G376) );
  NAND2_X1 U3479 ( .A1(n4980), .A2(n4966), .ZN(n4979) );
  XOR2_X1 U3480 ( .A(n4981), .B(n4982), .Z(n4980) );
  NOR2_X1 U3481 ( .A1(n4983), .A2(n4984), .ZN(n4982) );
  NAND2_X1 U3482 ( .A1(KEYINPUT77), .A2(n4947), .ZN(n4981) );
  NAND2_X1 U3483 ( .A1(n4985), .A2(n4977), .ZN(n4978) );
  XNOR2_X1 U3484 ( .A(n4984), .B(n4915), .ZN(n4985) );
  XNOR2_X1 U3485 ( .A(G4526), .B(n4986), .ZN(G373) );
  NAND2_X1 U3486 ( .A1(KEYINPUT35), .A2(n4882), .ZN(n4986) );
  NAND2_X1 U3487 ( .A1(n4987), .A2(n4988), .ZN(G370) );
  NAND2_X1 U3488 ( .A1(n4989), .A2(n4990), .ZN(n4988) );
  XOR2_X1 U3489 ( .A(n4991), .B(n4992), .Z(n4989) );
  XOR2_X1 U3490 ( .A(n4993), .B(n4994), .Z(n4992) );
  XOR2_X1 U3491 ( .A(n4995), .B(n4996), .Z(n4994) );
  XNOR2_X1 U3492 ( .A(n4997), .B(n4998), .ZN(n4996) );
  NAND2_X1 U3493 ( .A1(KEYINPUT95), .A2(n4999), .ZN(n4997) );
  NAND2_X1 U3494 ( .A1(n5000), .A2(n5001), .ZN(n4999) );
  XOR2_X1 U3495 ( .A(n5002), .B(n5003), .Z(n4995) );
  XOR2_X1 U3496 ( .A(n5004), .B(n5005), .Z(n4993) );
  XOR2_X1 U3497 ( .A(n5006), .B(n5007), .Z(n5005) );
  NOR2_X1 U3498 ( .A1(KEYINPUT19), .A2(n5008), .ZN(n5007) );
  NOR2_X1 U3499 ( .A1(n5009), .A2(n5010), .ZN(n5006) );
  XOR2_X1 U3500 ( .A(n5011), .B(n5012), .Z(n5004) );
  NOR2_X1 U3501 ( .A1(n5013), .A2(n5014), .ZN(n5012) );
  NAND2_X1 U3502 ( .A1(n5015), .A2(n5016), .ZN(n4987) );
  INV_X1 U3503 ( .A(n4990), .ZN(n5016) );
  XOR2_X1 U3504 ( .A(n5017), .B(n5018), .Z(n5015) );
  XNOR2_X1 U3505 ( .A(n5019), .B(n5008), .ZN(n5018) );
  XOR2_X1 U3506 ( .A(n5020), .B(n5021), .Z(n5017) );
  XOR2_X1 U3507 ( .A(n5022), .B(n5023), .Z(n5021) );
  XNOR2_X1 U3508 ( .A(n5014), .B(n5024), .ZN(n5023) );
  XOR2_X1 U3509 ( .A(n5010), .B(KEYINPUT125), .Z(n5022) );
  NAND2_X1 U3510 ( .A1(n5025), .A2(n5026), .ZN(n5010) );
  NAND2_X1 U3511 ( .A1(n5027), .A2(n5028), .ZN(n5025) );
  XNOR2_X1 U3512 ( .A(n5019), .B(KEYINPUT98), .ZN(n5027) );
  XOR2_X1 U3513 ( .A(n5029), .B(n5030), .Z(n5020) );
  XNOR2_X1 U3514 ( .A(n5031), .B(n5003), .ZN(n5030) );
  XNOR2_X1 U3515 ( .A(n5028), .B(n5032), .ZN(n5003) );
  NAND2_X1 U3516 ( .A1(KEYINPUT30), .A2(n5002), .ZN(n5031) );
  XOR2_X1 U3517 ( .A(n4991), .B(n5033), .Z(n5029) );
  NOR2_X1 U3518 ( .A1(KEYINPUT122), .A2(n5034), .ZN(n5033) );
  NAND3_X1 U3519 ( .A1(n5035), .A2(n5036), .A3(n5037), .ZN(n4991) );
  NAND3_X1 U3520 ( .A1(n5038), .A2(n4990), .A3(n5039), .ZN(n5037) );
  XOR2_X1 U3521 ( .A(KEYINPUT87), .B(n5040), .Z(n5039) );
  NAND2_X1 U3522 ( .A1(n5041), .A2(n5042), .ZN(n5038) );
  OR3_X1 U3523 ( .A1(n4990), .A2(n5040), .A3(n5041), .ZN(n5036) );
  XNOR2_X1 U3524 ( .A(n5043), .B(n5044), .ZN(n5040) );
  NAND2_X1 U3525 ( .A1(KEYINPUT76), .A2(n5045), .ZN(n5043) );
  XOR2_X1 U3526 ( .A(n5046), .B(n5047), .Z(n5045) );
  XOR2_X1 U3527 ( .A(n5048), .B(n5049), .Z(n5047) );
  NAND3_X1 U3528 ( .A1(n5050), .A2(n5051), .A3(KEYINPUT106), .ZN(n5049) );
  NAND2_X1 U3529 ( .A1(n5052), .A2(n5053), .ZN(n5051) );
  OR3_X1 U3530 ( .A1(n5054), .A2(n5052), .A3(n5053), .ZN(n5050) );
  NOR2_X1 U3531 ( .A1(n5055), .A2(n5056), .ZN(n5046) );
  NAND3_X1 U3532 ( .A1(n5057), .A2(n5058), .A3(n5041), .ZN(n5035) );
  INV_X1 U3533 ( .A(n5059), .ZN(n5041) );
  NAND2_X1 U3534 ( .A1(n5060), .A2(n4990), .ZN(n5058) );
  NAND3_X1 U3535 ( .A1(n4919), .A2(n5061), .A3(n5062), .ZN(n4990) );
  NAND2_X1 U3536 ( .A1(n5063), .A2(n5064), .ZN(n5062) );
  INV_X1 U3537 ( .A(n4906), .ZN(n5064) );
  NOR2_X1 U3538 ( .A1(n4932), .A2(n5065), .ZN(n4906) );
  XNOR2_X1 U3539 ( .A(n4931), .B(KEYINPUT127), .ZN(n4932) );
  XNOR2_X1 U3540 ( .A(n5044), .B(n5066), .ZN(n5057) );
  XOR2_X1 U3541 ( .A(n5048), .B(n5067), .Z(n5066) );
  NAND2_X1 U3542 ( .A1(n5068), .A2(n5069), .ZN(n5067) );
  OR2_X1 U3543 ( .A1(n5056), .A2(n5070), .ZN(n5069) );
  XOR2_X1 U3544 ( .A(n5071), .B(KEYINPUT9), .Z(n5068) );
  NAND2_X1 U3545 ( .A1(n5070), .A2(n5056), .ZN(n5071) );
  XNOR2_X1 U3546 ( .A(n5053), .B(n5072), .ZN(n5070) );
  NAND2_X1 U3547 ( .A1(n5073), .A2(n5074), .ZN(n5048) );
  NAND2_X1 U3548 ( .A1(n5075), .A2(n5076), .ZN(n5074) );
  NAND2_X1 U3549 ( .A1(n5077), .A2(n5078), .ZN(n5076) );
  NAND2_X1 U3550 ( .A1(n5054), .A2(n5078), .ZN(n5073) );
  XOR2_X1 U3551 ( .A(n5079), .B(n5080), .Z(n5044) );
  XNOR2_X1 U3552 ( .A(n5081), .B(n5082), .ZN(G368) );
  XNOR2_X1 U3553 ( .A(n5083), .B(n4998), .ZN(G365) );
  NAND2_X1 U3554 ( .A1(KEYINPUT22), .A2(n5084), .ZN(n5083) );
  NAND2_X1 U3555 ( .A1(n5085), .A2(n5026), .ZN(n5084) );
  NAND2_X1 U3556 ( .A1(n5028), .A2(n5082), .ZN(n5085) );
  NAND2_X1 U3557 ( .A1(n5086), .A2(n5087), .ZN(n5082) );
  NAND2_X1 U3558 ( .A1(n5088), .A2(n5011), .ZN(n5087) );
  XNOR2_X1 U3559 ( .A(n5032), .B(n5089), .ZN(G362) );
  XNOR2_X1 U3560 ( .A(n5090), .B(n5008), .ZN(G359) );
  NAND2_X1 U3561 ( .A1(n5091), .A2(n5092), .ZN(n5090) );
  NAND2_X1 U3562 ( .A1(n5093), .A2(n5089), .ZN(n5092) );
  NAND2_X1 U3563 ( .A1(n5000), .A2(n5094), .ZN(n5089) );
  NAND3_X1 U3564 ( .A1(n5095), .A2(n5088), .A3(n5096), .ZN(n5094) );
  INV_X1 U3565 ( .A(n5024), .ZN(n5000) );
  XOR2_X1 U3566 ( .A(n5097), .B(KEYINPUT109), .Z(n5091) );
  NAND2_X1 U3567 ( .A1(n5098), .A2(n5099), .ZN(G356) );
  NAND2_X1 U3568 ( .A1(n5100), .A2(n5101), .ZN(n5099) );
  OR2_X1 U3569 ( .A1(n5102), .A2(n5100), .ZN(n5098) );
  NAND2_X1 U3570 ( .A1(n5103), .A2(n5104), .ZN(G353) );
  NAND2_X1 U3571 ( .A1(n5105), .A2(n5101), .ZN(n5104) );
  XNOR2_X1 U3572 ( .A(n5106), .B(n5078), .ZN(n5105) );
  NAND3_X1 U3573 ( .A1(n5107), .A2(n5108), .A3(n5109), .ZN(n5103) );
  NAND2_X1 U3574 ( .A1(KEYINPUT113), .A2(n5110), .ZN(n5108) );
  XNOR2_X1 U3575 ( .A(n5106), .B(n5077), .ZN(n5110) );
  NAND3_X1 U3576 ( .A1(n5111), .A2(n5112), .A3(n5113), .ZN(n5107) );
  INV_X1 U3577 ( .A(KEYINPUT113), .ZN(n5113) );
  NAND2_X1 U3578 ( .A1(n5077), .A2(n5106), .ZN(n5111) );
  NAND2_X1 U3579 ( .A1(n5114), .A2(n5115), .ZN(G350) );
  NAND2_X1 U3580 ( .A1(n5116), .A2(n5109), .ZN(n5115) );
  XOR2_X1 U3581 ( .A(n5117), .B(n5118), .Z(n5116) );
  NAND2_X1 U3582 ( .A1(n5119), .A2(n5101), .ZN(n5114) );
  XOR2_X1 U3583 ( .A(n5120), .B(n5121), .Z(n5119) );
  NOR2_X1 U3584 ( .A1(KEYINPUT38), .A2(n5117), .ZN(n5121) );
  NAND2_X1 U3585 ( .A1(n5118), .A2(n5122), .ZN(n5120) );
  NAND2_X1 U3586 ( .A1(n5123), .A2(n5124), .ZN(G347) );
  NAND2_X1 U3587 ( .A1(n5125), .A2(n5126), .ZN(n5124) );
  NAND2_X1 U3588 ( .A1(n5127), .A2(n5128), .ZN(n5125) );
  NAND2_X1 U3589 ( .A1(n5129), .A2(n5101), .ZN(n5128) );
  NAND3_X1 U3590 ( .A1(n5130), .A2(n5131), .A3(n5132), .ZN(n5129) );
  NAND2_X1 U3591 ( .A1(n5109), .A2(n5133), .ZN(n5127) );
  INV_X1 U3592 ( .A(n5102), .ZN(n5109) );
  NAND3_X1 U3593 ( .A1(n5132), .A2(n5134), .A3(n5079), .ZN(n5123) );
  NAND2_X1 U3594 ( .A1(n5102), .A2(n5135), .ZN(n5134) );
  NAND3_X1 U3595 ( .A1(n5130), .A2(n5131), .A3(n5101), .ZN(n5135) );
  INV_X1 U3596 ( .A(KEYINPUT101), .ZN(n5131) );
  INV_X1 U3597 ( .A(n5136), .ZN(n5130) );
  XNOR2_X1 U3598 ( .A(n5101), .B(KEYINPUT92), .ZN(n5102) );
  NAND2_X1 U3599 ( .A1(n5137), .A2(n5138), .ZN(n5101) );
  NAND2_X1 U3600 ( .A1(n5139), .A2(n5088), .ZN(n5138) );
  NAND2_X1 U3601 ( .A1(n5140), .A2(n5141), .ZN(G344) );
  NAND2_X1 U3602 ( .A1(n5142), .A2(n5096), .ZN(n5141) );
  XOR2_X1 U3603 ( .A(KEYINPUT3), .B(n5143), .Z(n5140) );
  NOR2_X1 U3604 ( .A1(n5142), .A2(n5096), .ZN(n5143) );
  INV_X1 U3605 ( .A(n5088), .ZN(n5142) );
  NAND2_X1 U3606 ( .A1(n5144), .A2(n5145), .ZN(n5088) );
  NAND2_X1 U3607 ( .A1(n5146), .A2(n4966), .ZN(n5145) );
  INV_X1 U3608 ( .A(n4977), .ZN(n4966) );
  NOR2_X1 U3609 ( .A1(n5147), .A2(n5148), .ZN(n4977) );
  INV_X1 U3610 ( .A(G15), .ZN(G341) );
  XOR2_X1 U3611 ( .A(n5149), .B(n5150), .Z(G338) );
  NAND2_X1 U3612 ( .A1(n5151), .A2(n5152), .ZN(n5150) );
  NAND2_X1 U3613 ( .A1(n5153), .A2(n5154), .ZN(n5152) );
  XOR2_X1 U3614 ( .A(n5155), .B(n5156), .Z(n5153) );
  XOR2_X1 U3615 ( .A(n5157), .B(n5158), .Z(n5156) );
  XOR2_X1 U3616 ( .A(n5159), .B(n5160), .Z(n5158) );
  NAND2_X1 U3617 ( .A1(n5161), .A2(n5162), .ZN(n5159) );
  INV_X1 U3618 ( .A(n5163), .ZN(n5161) );
  NOR2_X1 U3619 ( .A1(n5164), .A2(n5165), .ZN(n5157) );
  AND2_X1 U3620 ( .A1(n5166), .A2(n5167), .ZN(n5164) );
  XOR2_X1 U3621 ( .A(n5168), .B(n5169), .Z(n5155) );
  XNOR2_X1 U3622 ( .A(n5170), .B(n5171), .ZN(n5169) );
  XNOR2_X1 U3623 ( .A(n5172), .B(n5173), .ZN(n5168) );
  NOR2_X1 U3624 ( .A1(KEYINPUT73), .A2(n5174), .ZN(n5172) );
  NOR2_X1 U3625 ( .A1(n5167), .A2(n5175), .ZN(n5174) );
  NAND2_X1 U3626 ( .A1(n5176), .A2(n5177), .ZN(n5151) );
  XNOR2_X1 U3627 ( .A(n5171), .B(n5178), .ZN(n5177) );
  NOR2_X1 U3628 ( .A1(n5179), .A2(n5180), .ZN(n5178) );
  XOR2_X1 U3629 ( .A(n5181), .B(KEYINPUT83), .Z(n5180) );
  NAND2_X1 U3630 ( .A1(n5182), .A2(n5166), .ZN(n5181) );
  NOR2_X1 U3631 ( .A1(n5166), .A2(n5182), .ZN(n5179) );
  XNOR2_X1 U3632 ( .A(n5183), .B(n5184), .ZN(n5182) );
  XOR2_X1 U3633 ( .A(n5175), .B(n5160), .Z(n5184) );
  NAND3_X1 U3634 ( .A1(n5185), .A2(n5186), .A3(n5187), .ZN(n5160) );
  NAND2_X1 U3635 ( .A1(n5188), .A2(n5189), .ZN(n5187) );
  XNOR2_X1 U3636 ( .A(n5190), .B(n5191), .ZN(n5188) );
  NAND3_X1 U3637 ( .A1(n5192), .A2(n5190), .A3(n5193), .ZN(n5186) );
  NAND2_X1 U3638 ( .A1(n5167), .A2(n5191), .ZN(n5185) );
  NAND2_X1 U3639 ( .A1(n5194), .A2(n5195), .ZN(n5175) );
  XOR2_X1 U3640 ( .A(KEYINPUT8), .B(n5196), .Z(n5194) );
  NOR2_X1 U3641 ( .A1(n5197), .A2(n5190), .ZN(n5196) );
  XOR2_X1 U3642 ( .A(n5198), .B(n5199), .Z(n5183) );
  NOR3_X1 U3643 ( .A1(n5200), .A2(n5201), .A3(n5202), .ZN(n5199) );
  NOR2_X1 U3644 ( .A1(KEYINPUT74), .A2(n5203), .ZN(n5202) );
  NOR2_X1 U3645 ( .A1(n5204), .A2(n5205), .ZN(n5203) );
  NOR2_X1 U3646 ( .A1(n5206), .A2(n5204), .ZN(n5200) );
  NOR3_X1 U3647 ( .A1(n5207), .A2(n5208), .A3(n5209), .ZN(n5206) );
  NOR2_X1 U3648 ( .A1(n5205), .A2(n5210), .ZN(n5209) );
  INV_X1 U3649 ( .A(KEYINPUT74), .ZN(n5210) );
  NOR2_X1 U3650 ( .A1(n5173), .A2(n5195), .ZN(n5207) );
  NAND2_X1 U3651 ( .A1(n5211), .A2(n5212), .ZN(n5198) );
  NAND2_X1 U3652 ( .A1(n5213), .A2(n5197), .ZN(n5212) );
  NAND2_X1 U3653 ( .A1(n5214), .A2(n5215), .ZN(n5211) );
  INV_X1 U3654 ( .A(n5154), .ZN(n5176) );
  NAND2_X1 U3655 ( .A1(n5216), .A2(n5217), .ZN(n5149) );
  NAND3_X1 U3656 ( .A1(n5218), .A2(n5219), .A3(n5220), .ZN(n5217) );
  XOR2_X1 U3657 ( .A(n4515), .B(n5221), .Z(n5218) );
  XNOR2_X1 U3658 ( .A(n5222), .B(KEYINPUT110), .ZN(n5221) );
  NAND2_X1 U3659 ( .A1(n5223), .A2(n5224), .ZN(n5216) );
  NAND2_X1 U3660 ( .A1(n5220), .A2(n5219), .ZN(n5224) );
  NAND2_X1 U3661 ( .A1(n5225), .A2(n5154), .ZN(n5219) );
  INV_X1 U3662 ( .A(n5226), .ZN(n5220) );
  XOR2_X1 U3663 ( .A(n5227), .B(n5228), .Z(n5223) );
  XOR2_X1 U3664 ( .A(n5229), .B(n5222), .Z(n5228) );
  NOR2_X1 U3665 ( .A1(n5230), .A2(n5231), .ZN(n5222) );
  AND2_X1 U3666 ( .A1(n4514), .A2(n4511), .ZN(n5230) );
  NOR2_X1 U3667 ( .A1(n4518), .A2(n5232), .ZN(n5229) );
  NOR2_X1 U3668 ( .A1(n5227), .A2(KEYINPUT20), .ZN(n5232) );
  INV_X1 U3669 ( .A(n5233), .ZN(n4518) );
  NOR2_X1 U3670 ( .A1(n5231), .A2(n5234), .ZN(n5227) );
  NAND2_X1 U3671 ( .A1(n5235), .A2(n5236), .ZN(G336) );
  OR2_X1 U3672 ( .A1(n5237), .A2(n5238), .ZN(n5236) );
  XOR2_X1 U3673 ( .A(n5239), .B(KEYINPUT14), .Z(n5235) );
  NAND2_X1 U3674 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  XOR2_X1 U3675 ( .A(n5240), .B(KEYINPUT89), .Z(n5238) );
  XNOR2_X1 U3676 ( .A(n5166), .B(n5241), .ZN(G333) );
  NAND2_X1 U3677 ( .A1(KEYINPUT75), .A2(n5242), .ZN(n5241) );
  NAND2_X1 U3678 ( .A1(n5243), .A2(n5195), .ZN(n5242) );
  NAND2_X1 U3679 ( .A1(n5240), .A2(n5237), .ZN(n5243) );
  XNOR2_X1 U3680 ( .A(n5244), .B(n5245), .ZN(G330) );
  XOR2_X1 U3681 ( .A(n5246), .B(n5247), .Z(G327) );
  NAND2_X1 U3682 ( .A1(n5248), .A2(n5249), .ZN(n5247) );
  OR2_X1 U3683 ( .A1(n5245), .A2(n5250), .ZN(n5249) );
  NOR2_X1 U3684 ( .A1(n5213), .A2(n5251), .ZN(n5245) );
  AND3_X1 U3685 ( .A1(n5166), .A2(n5237), .A3(n5240), .ZN(n5251) );
  INV_X1 U3686 ( .A(n5252), .ZN(n5240) );
  NAND2_X1 U3687 ( .A1(n5197), .A2(n5253), .ZN(n5237) );
  NAND2_X1 U3688 ( .A1(n5192), .A2(n5254), .ZN(n5253) );
  NAND2_X1 U3689 ( .A1(KEYINPUT24), .A2(n5255), .ZN(n5246) );
  XNOR2_X1 U3690 ( .A(n5189), .B(n5254), .ZN(G324) );
  XOR2_X1 U3691 ( .A(n5256), .B(n5257), .Z(G321) );
  NOR2_X1 U3692 ( .A1(n5258), .A2(n5259), .ZN(n5257) );
  NOR2_X1 U3693 ( .A1(n5260), .A2(n5261), .ZN(n5259) );
  XOR2_X1 U3694 ( .A(n5262), .B(n5263), .Z(n5261) );
  XOR2_X1 U3695 ( .A(n5264), .B(n5265), .Z(n5263) );
  XNOR2_X1 U3696 ( .A(n5266), .B(n5267), .ZN(n5265) );
  XOR2_X1 U3697 ( .A(n5268), .B(n5269), .Z(n5264) );
  NOR2_X1 U3698 ( .A1(n5270), .A2(n5271), .ZN(n5269) );
  NOR2_X1 U3699 ( .A1(KEYINPUT91), .A2(n5272), .ZN(n5268) );
  XOR2_X1 U3700 ( .A(n5273), .B(n5274), .Z(n5262) );
  XOR2_X1 U3701 ( .A(n5275), .B(n5276), .Z(n5274) );
  XOR2_X1 U3702 ( .A(KEYINPUT68), .B(KEYINPUT17), .Z(n5273) );
  NOR2_X1 U3703 ( .A1(n5277), .A2(n5278), .ZN(n5258) );
  XNOR2_X1 U3704 ( .A(n5279), .B(n5267), .ZN(n5278) );
  XNOR2_X1 U3705 ( .A(n5280), .B(n5281), .ZN(n5267) );
  NAND2_X1 U3706 ( .A1(KEYINPUT112), .A2(n5282), .ZN(n5279) );
  XOR2_X1 U3707 ( .A(n5283), .B(n5284), .Z(n5282) );
  XOR2_X1 U3708 ( .A(n5285), .B(n5266), .Z(n5284) );
  XOR2_X1 U3709 ( .A(n5286), .B(n5287), .Z(n5266) );
  NOR2_X1 U3710 ( .A1(n5271), .A2(n4821), .ZN(n5285) );
  XOR2_X1 U3711 ( .A(n5288), .B(n5289), .Z(n5283) );
  XOR2_X1 U3712 ( .A(n5290), .B(n5291), .Z(n5289) );
  NOR2_X1 U3713 ( .A1(n5292), .A2(n5276), .ZN(n5291) );
  NAND2_X1 U3714 ( .A1(n5293), .A2(n5294), .ZN(n5276) );
  NAND2_X1 U3715 ( .A1(n5295), .A2(n5270), .ZN(n5294) );
  XNOR2_X1 U3716 ( .A(n5286), .B(KEYINPUT27), .ZN(n5295) );
  NOR2_X1 U3717 ( .A1(n5296), .A2(n5272), .ZN(n5290) );
  NOR2_X1 U3718 ( .A1(n5297), .A2(n5275), .ZN(n5288) );
  NAND2_X1 U3719 ( .A1(n5298), .A2(n5299), .ZN(n5256) );
  NAND2_X1 U3720 ( .A1(n5300), .A2(n5301), .ZN(n5299) );
  INV_X1 U3721 ( .A(n5302), .ZN(n5301) );
  XOR2_X1 U3722 ( .A(n5303), .B(n5304), .Z(n5300) );
  XNOR2_X1 U3723 ( .A(n5305), .B(n5306), .ZN(n5304) );
  NAND2_X1 U3724 ( .A1(n5307), .A2(n5308), .ZN(n5306) );
  NAND2_X1 U3725 ( .A1(n5309), .A2(n5310), .ZN(n5308) );
  NAND2_X1 U3726 ( .A1(n5311), .A2(n5312), .ZN(n5307) );
  XOR2_X1 U3727 ( .A(n5313), .B(n5314), .Z(n5303) );
  NAND2_X1 U3728 ( .A1(n5315), .A2(n5316), .ZN(n5314) );
  NAND2_X1 U3729 ( .A1(n5317), .A2(n5302), .ZN(n5298) );
  NOR2_X1 U3730 ( .A1(n5318), .A2(n5319), .ZN(n5302) );
  AND3_X1 U3731 ( .A1(n5287), .A2(n5260), .A3(n5296), .ZN(n5319) );
  XNOR2_X1 U3732 ( .A(n5305), .B(n5320), .ZN(n5317) );
  XNOR2_X1 U3733 ( .A(n5321), .B(n5313), .ZN(n5320) );
  NAND3_X1 U3734 ( .A1(n5322), .A2(n5323), .A3(n5316), .ZN(n5313) );
  INV_X1 U3735 ( .A(n5324), .ZN(n5316) );
  NAND2_X1 U3736 ( .A1(n5325), .A2(n5326), .ZN(n5323) );
  XNOR2_X1 U3737 ( .A(n5327), .B(n5328), .ZN(n5325) );
  NAND3_X1 U3738 ( .A1(n5328), .A2(n5329), .A3(n5330), .ZN(n5322) );
  NAND3_X1 U3739 ( .A1(n5331), .A2(n5332), .A3(n5333), .ZN(n5321) );
  NAND2_X1 U3740 ( .A1(KEYINPUT71), .A2(n5334), .ZN(n5333) );
  NAND2_X1 U3741 ( .A1(n5315), .A2(n5335), .ZN(n5334) );
  NAND2_X1 U3742 ( .A1(n5336), .A2(KEYINPUT116), .ZN(n5335) );
  NAND4_X1 U3743 ( .A1(n5337), .A2(n5338), .A3(n5315), .A4(n5336), .ZN(n5332) );
  INV_X1 U3744 ( .A(n5339), .ZN(n5336) );
  NAND2_X1 U3745 ( .A1(n5339), .A2(n5340), .ZN(n5331) );
  NAND3_X1 U3746 ( .A1(n5341), .A2(n5342), .A3(n5343), .ZN(n5340) );
  NAND2_X1 U3747 ( .A1(KEYINPUT71), .A2(n5337), .ZN(n5343) );
  INV_X1 U3748 ( .A(KEYINPUT116), .ZN(n5337) );
  NAND2_X1 U3749 ( .A1(KEYINPUT45), .A2(n5315), .ZN(n5342) );
  NAND2_X1 U3750 ( .A1(n5344), .A2(n5345), .ZN(n5341) );
  INV_X1 U3751 ( .A(KEYINPUT45), .ZN(n5345) );
  NAND2_X1 U3752 ( .A1(n5315), .A2(n5346), .ZN(n5344) );
  NAND2_X1 U3753 ( .A1(KEYINPUT116), .A2(n5338), .ZN(n5346) );
  INV_X1 U3754 ( .A(KEYINPUT71), .ZN(n5338) );
  AND2_X1 U3755 ( .A1(n5347), .A2(n5348), .ZN(n5315) );
  NAND2_X1 U3756 ( .A1(n5349), .A2(n5310), .ZN(n5348) );
  XNOR2_X1 U3757 ( .A(n5350), .B(n5310), .ZN(n5339) );
  XNOR2_X1 U3758 ( .A(n5351), .B(n5352), .ZN(G319) );
  NAND2_X1 U3759 ( .A1(n5353), .A2(n5354), .ZN(n5351) );
  NAND2_X1 U3760 ( .A1(n5271), .A2(n5355), .ZN(n5354) );
  XOR2_X1 U3761 ( .A(n5356), .B(n5281), .Z(G316) );
  NAND3_X1 U3762 ( .A1(n5357), .A2(n5358), .A3(KEYINPUT100), .ZN(n5356) );
  NAND3_X1 U3763 ( .A1(n5359), .A2(n5355), .A3(n5286), .ZN(n5358) );
  XOR2_X1 U3764 ( .A(KEYINPUT102), .B(n5271), .Z(n5359) );
  INV_X1 U3765 ( .A(n5360), .ZN(n5357) );
  XOR2_X1 U3766 ( .A(n5361), .B(n5362), .Z(G313) );
  XNOR2_X1 U3767 ( .A(n5363), .B(n5364), .ZN(G310) );
  NAND2_X1 U3768 ( .A1(n5365), .A2(n5366), .ZN(n5363) );
  NAND2_X1 U3769 ( .A1(n5362), .A2(n5361), .ZN(n5365) );
  OR2_X1 U3770 ( .A1(n5275), .A2(n5367), .ZN(n5361) );
  XNOR2_X1 U3771 ( .A(n5327), .B(n5368), .ZN(G307) );
  NAND2_X1 U3772 ( .A1(n5369), .A2(n5370), .ZN(G304) );
  NAND2_X1 U3773 ( .A1(n5371), .A2(n5372), .ZN(n5370) );
  XNOR2_X1 U3774 ( .A(n5330), .B(n5309), .ZN(n5371) );
  NAND2_X1 U3775 ( .A1(n5368), .A2(n5373), .ZN(n5369) );
  NAND2_X1 U3776 ( .A1(n5374), .A2(n5375), .ZN(n5373) );
  NAND2_X1 U3777 ( .A1(KEYINPUT115), .A2(n5376), .ZN(n5375) );
  NAND2_X1 U3778 ( .A1(n5377), .A2(n5378), .ZN(n5376) );
  OR2_X1 U3779 ( .A1(n5330), .A2(n5350), .ZN(n5378) );
  NAND2_X1 U3780 ( .A1(n5379), .A2(n5380), .ZN(n5374) );
  INV_X1 U3781 ( .A(KEYINPUT115), .ZN(n5380) );
  XNOR2_X1 U3782 ( .A(n5350), .B(n5326), .ZN(n5379) );
  XNOR2_X1 U3783 ( .A(n5381), .B(n5382), .ZN(G301) );
  NOR2_X1 U3784 ( .A1(n5383), .A2(n5310), .ZN(n5382) );
  NOR2_X1 U3785 ( .A1(n5368), .A2(n5311), .ZN(n5383) );
  NAND2_X1 U3786 ( .A1(n5384), .A2(n5385), .ZN(G298) );
  NAND2_X1 U3787 ( .A1(n5386), .A2(n5372), .ZN(n5385) );
  INV_X1 U3788 ( .A(n5368), .ZN(n5372) );
  XOR2_X1 U3789 ( .A(n5387), .B(KEYINPUT4), .Z(n5386) );
  NAND2_X1 U3790 ( .A1(n5388), .A2(n5389), .ZN(n5387) );
  NAND3_X1 U3791 ( .A1(n5390), .A2(n5347), .A3(n5391), .ZN(n5389) );
  XOR2_X1 U3792 ( .A(n5392), .B(KEYINPUT63), .Z(n5388) );
  NAND2_X1 U3793 ( .A1(n5393), .A2(n5394), .ZN(n5392) );
  NAND2_X1 U3794 ( .A1(n5390), .A2(n5347), .ZN(n5394) );
  OR2_X1 U3795 ( .A1(n5395), .A2(n5311), .ZN(n5390) );
  NOR2_X1 U3796 ( .A1(n5310), .A2(n5396), .ZN(n5311) );
  NOR2_X1 U3797 ( .A1(n5329), .A2(n5326), .ZN(n5396) );
  NAND2_X1 U3798 ( .A1(n5368), .A2(n5397), .ZN(n5384) );
  XNOR2_X1 U3799 ( .A(n5398), .B(n5393), .ZN(n5397) );
  NOR2_X1 U3800 ( .A1(n5399), .A2(n5400), .ZN(n5368) );
  AND3_X1 U3801 ( .A1(n5362), .A2(n5287), .A3(n5367), .ZN(n5400) );
  AND2_X1 U3802 ( .A1(n5297), .A2(n5355), .ZN(n5367) );
  XOR2_X1 U3803 ( .A(n5355), .B(n5271), .Z(G295) );
  NAND3_X1 U3804 ( .A1(G133), .A2(n5401), .A3(G134), .ZN(G292) );
  NAND2_X1 U3805 ( .A1(G1197), .A2(n5401), .ZN(G289) );
  INV_X1 U3806 ( .A(G5), .ZN(n5401) );
  XNOR2_X1 U3807 ( .A(G15), .B(KEYINPUT117), .ZN(G286) );
  AND2_X1 U3808 ( .A1(G1), .A2(G163), .ZN(G278) );
  NAND2_X1 U3809 ( .A1(n5402), .A2(n5403), .ZN(G276) );
  NAND2_X1 U3810 ( .A1(n5404), .A2(n5154), .ZN(n5403) );
  NAND2_X1 U3811 ( .A1(n5405), .A2(n5406), .ZN(n5154) );
  NAND2_X1 U3812 ( .A1(n5407), .A2(n5260), .ZN(n5406) );
  INV_X1 U3813 ( .A(n5277), .ZN(n5260) );
  NOR2_X1 U3814 ( .A1(n5408), .A2(n5409), .ZN(n5277) );
  AND4_X1 U3815 ( .A1(n5055), .A2(n5060), .A3(n5079), .A4(n5410), .ZN(n5409) );
  NAND2_X1 U3816 ( .A1(n5411), .A2(n5412), .ZN(n5410) );
  NAND2_X1 U3817 ( .A1(n5065), .A2(n5063), .ZN(n5412) );
  INV_X1 U3818 ( .A(n5413), .ZN(n5411) );
  NAND2_X1 U3819 ( .A1(n5414), .A2(n5415), .ZN(G273) );
  NAND2_X1 U3820 ( .A1(n5231), .A2(n4512), .ZN(n5415) );
  NAND2_X1 U3821 ( .A1(n5416), .A2(n5417), .ZN(n4512) );
  NAND2_X1 U3822 ( .A1(n5418), .A2(n5254), .ZN(n5417) );
  NAND3_X1 U3823 ( .A1(n5419), .A2(n5420), .A3(n5421), .ZN(n5254) );
  XOR2_X1 U3824 ( .A(n5422), .B(KEYINPUT29), .Z(n5421) );
  NAND2_X1 U3825 ( .A1(n5423), .A2(n5424), .ZN(n5422) );
  NAND2_X1 U3826 ( .A1(n5424), .A2(n5425), .ZN(n5420) );
  NAND3_X1 U3827 ( .A1(n5426), .A2(n5427), .A3(n5402), .ZN(G270) );
  AND2_X1 U3828 ( .A1(n5414), .A2(n5428), .ZN(n5402) );
  NAND2_X1 U3829 ( .A1(n5231), .A2(n5226), .ZN(n5428) );
  NAND2_X1 U3830 ( .A1(n5429), .A2(n5430), .ZN(n5226) );
  NAND2_X1 U3831 ( .A1(n5191), .A2(n5163), .ZN(n5430) );
  NAND2_X1 U3832 ( .A1(n5248), .A2(n5431), .ZN(n5163) );
  NAND2_X1 U3833 ( .A1(n5171), .A2(n5165), .ZN(n5431) );
  INV_X1 U3834 ( .A(n5214), .ZN(n5165) );
  NOR2_X1 U3835 ( .A1(n5213), .A2(n5208), .ZN(n5214) );
  NOR3_X1 U3836 ( .A1(n5197), .A2(n5173), .A3(n5190), .ZN(n5208) );
  NAND4_X1 U3837 ( .A1(n5079), .A2(n5432), .A3(n5060), .A4(n5433), .ZN(n5427) );
  NOR2_X1 U3838 ( .A1(n5434), .A2(n5435), .ZN(n5433) );
  INV_X1 U3839 ( .A(n5042), .ZN(n5060) );
  NAND2_X1 U3840 ( .A1(n5013), .A2(n5436), .ZN(n5042) );
  NOR2_X1 U3841 ( .A1(n5001), .A2(n5032), .ZN(n5013) );
  NAND2_X1 U3842 ( .A1(n5009), .A2(n4998), .ZN(n5001) );
  AND2_X1 U3843 ( .A1(n5028), .A2(n5002), .ZN(n5009) );
  NAND2_X1 U3844 ( .A1(n5437), .A2(n5438), .ZN(n5002) );
  NAND2_X1 U3845 ( .A1(n5096), .A2(n5439), .ZN(n5438) );
  INV_X1 U3846 ( .A(KEYINPUT94), .ZN(n5439) );
  NAND2_X1 U3847 ( .A1(KEYINPUT94), .A2(G4394), .ZN(n5437) );
  INV_X1 U3848 ( .A(n5081), .ZN(n5028) );
  NAND2_X1 U3849 ( .A1(n5440), .A2(n5441), .ZN(n5432) );
  NAND3_X1 U3850 ( .A1(n5063), .A2(n5442), .A3(n5065), .ZN(n5441) );
  INV_X1 U3851 ( .A(n4930), .ZN(n5065) );
  NAND3_X1 U3852 ( .A1(n5443), .A2(G4526), .A3(n4871), .ZN(n4930) );
  NOR2_X1 U3853 ( .A1(n4867), .A2(n4878), .ZN(n4871) );
  INV_X1 U3854 ( .A(n4882), .ZN(n4878) );
  XNOR2_X1 U3855 ( .A(KEYINPUT121), .B(n5444), .ZN(n5442) );
  NAND2_X1 U3856 ( .A1(n5445), .A2(n5413), .ZN(n5440) );
  NAND3_X1 U3857 ( .A1(n4919), .A2(n5061), .A3(n5446), .ZN(n5413) );
  NAND2_X1 U3858 ( .A1(n5063), .A2(n4931), .ZN(n5446) );
  NAND3_X1 U3859 ( .A1(n5447), .A2(n5448), .A3(n5449), .ZN(n4931) );
  XOR2_X1 U3860 ( .A(n5450), .B(KEYINPUT81), .Z(n5449) );
  NAND2_X1 U3861 ( .A1(n4879), .A2(n5451), .ZN(n5448) );
  INV_X1 U3862 ( .A(n4867), .ZN(n4879) );
  NAND3_X1 U3863 ( .A1(n5452), .A2(n5453), .A3(n4869), .ZN(n4867) );
  OR3_X1 U3864 ( .A1(n5454), .A2(n4805), .A3(KEYINPUT93), .ZN(n5453) );
  NAND2_X1 U3865 ( .A1(KEYINPUT93), .A2(n5454), .ZN(n5452) );
  AND3_X1 U3866 ( .A1(n4947), .A2(n4964), .A3(n4945), .ZN(n5063) );
  NOR2_X1 U3867 ( .A1(n4942), .A2(n4925), .ZN(n4945) );
  INV_X1 U3868 ( .A(n4910), .ZN(n4942) );
  INV_X1 U3869 ( .A(n4923), .ZN(n4964) );
  NAND2_X1 U3870 ( .A1(n4947), .A2(n4917), .ZN(n4919) );
  NAND2_X1 U3871 ( .A1(n5455), .A2(n5456), .ZN(n4917) );
  NAND2_X1 U3872 ( .A1(n5457), .A2(n4920), .ZN(n5456) );
  NAND2_X1 U3873 ( .A1(n5458), .A2(n5459), .ZN(n4920) );
  NAND2_X1 U3874 ( .A1(n4910), .A2(n4916), .ZN(n5459) );
  XOR2_X1 U3875 ( .A(n5460), .B(KEYINPUT80), .Z(n4910) );
  XNOR2_X1 U3876 ( .A(n5404), .B(KEYINPUT99), .ZN(n5445) );
  NAND2_X1 U3877 ( .A1(n5404), .A2(n5461), .ZN(n5426) );
  NAND2_X1 U3878 ( .A1(n5405), .A2(n5462), .ZN(n5461) );
  NAND2_X1 U3879 ( .A1(n5407), .A2(n5408), .ZN(n5462) );
  NAND2_X1 U3880 ( .A1(n5463), .A2(n5464), .ZN(n5408) );
  NAND2_X1 U3881 ( .A1(n5079), .A2(n5465), .ZN(n5464) );
  NAND2_X1 U3882 ( .A1(n5466), .A2(n5467), .ZN(n5465) );
  NAND2_X1 U3883 ( .A1(n5055), .A2(n5059), .ZN(n5467) );
  NAND2_X1 U3884 ( .A1(n5468), .A2(n5469), .ZN(n5059) );
  XOR2_X1 U3885 ( .A(n5470), .B(KEYINPUT32), .Z(n5468) );
  INV_X1 U3886 ( .A(n5434), .ZN(n5055) );
  NAND3_X1 U3887 ( .A1(n5080), .A2(n5078), .A3(n5054), .ZN(n5434) );
  NOR2_X1 U3888 ( .A1(n5072), .A2(n5075), .ZN(n5054) );
  INV_X1 U3889 ( .A(n5471), .ZN(n5075) );
  INV_X1 U3890 ( .A(n5052), .ZN(n5078) );
  NOR2_X1 U3891 ( .A1(n5472), .A2(n4780), .ZN(n5052) );
  INV_X1 U3892 ( .A(n5056), .ZN(n5466) );
  NAND3_X1 U3893 ( .A1(n5473), .A2(n5474), .A3(n5475), .ZN(n5056) );
  NAND2_X1 U3894 ( .A1(n5080), .A2(n5053), .ZN(n5475) );
  NAND2_X1 U3895 ( .A1(n5476), .A2(n5477), .ZN(n5053) );
  NAND2_X1 U3896 ( .A1(n5072), .A2(n5471), .ZN(n5477) );
  NAND3_X1 U3897 ( .A1(n5478), .A2(n5479), .A3(n5480), .ZN(n5471) );
  NAND2_X1 U3898 ( .A1(n4510), .A2(n5481), .ZN(n5480) );
  NAND2_X1 U3899 ( .A1(KEYINPUT69), .A2(n5482), .ZN(n5479) );
  NAND3_X1 U3900 ( .A1(n5483), .A2(n5484), .A3(n5476), .ZN(n5482) );
  NAND2_X1 U3901 ( .A1(n4779), .A2(n5481), .ZN(n5484) );
  NAND3_X1 U3902 ( .A1(G4427), .A2(n4782), .A3(KEYINPUT118), .ZN(n5483) );
  NAND2_X1 U3903 ( .A1(n5485), .A2(n5486), .ZN(n5478) );
  INV_X1 U3904 ( .A(KEYINPUT69), .ZN(n5486) );
  XNOR2_X1 U3905 ( .A(n5487), .B(n4779), .ZN(n5485) );
  NOR2_X1 U3906 ( .A1(n4510), .A2(n5481), .ZN(n5487) );
  INV_X1 U3907 ( .A(KEYINPUT118), .ZN(n5481) );
  AND2_X1 U3908 ( .A1(n5488), .A2(n5489), .ZN(n5080) );
  NAND2_X1 U3909 ( .A1(n5490), .A2(n5491), .ZN(n5489) );
  NAND2_X1 U3910 ( .A1(n5492), .A2(n5493), .ZN(n5488) );
  NAND2_X1 U3911 ( .A1(n4765), .A2(n5491), .ZN(n5493) );
  INV_X1 U3912 ( .A(KEYINPUT103), .ZN(n5491) );
  OR3_X1 U3913 ( .A1(n5492), .A2(n4765), .A3(KEYINPUT28), .ZN(n5474) );
  INV_X1 U3914 ( .A(n5494), .ZN(n5492) );
  NAND2_X1 U3915 ( .A1(KEYINPUT28), .A2(n5490), .ZN(n5473) );
  INV_X1 U3916 ( .A(n5495), .ZN(n5490) );
  INV_X1 U3917 ( .A(n5435), .ZN(n5407) );
  NAND4_X1 U3918 ( .A1(n5296), .A2(n5324), .A3(n5287), .A4(n5305), .ZN(n5435) );
  AND2_X1 U3919 ( .A1(n5297), .A2(n5280), .ZN(n5296) );
  AND2_X1 U3920 ( .A1(n5496), .A2(n5497), .ZN(n5405) );
  NAND2_X1 U3921 ( .A1(n5305), .A2(n5498), .ZN(n5497) );
  NAND4_X1 U3922 ( .A1(n5499), .A2(n5347), .A3(n5500), .A4(n5501), .ZN(n5498) );
  NAND2_X1 U3923 ( .A1(n5349), .A2(n5502), .ZN(n5501) );
  NAND2_X1 U3924 ( .A1(n5377), .A2(n5503), .ZN(n5502) );
  OR2_X1 U3925 ( .A1(n5504), .A2(KEYINPUT105), .ZN(n5503) );
  INV_X1 U3926 ( .A(n5328), .ZN(n5349) );
  NAND3_X1 U3927 ( .A1(KEYINPUT105), .A2(n5505), .A3(n5328), .ZN(n5500) );
  NAND2_X1 U3928 ( .A1(n5324), .A2(n5318), .ZN(n5499) );
  NAND2_X1 U3929 ( .A1(n5506), .A2(n5507), .ZN(n5318) );
  NAND2_X1 U3930 ( .A1(n5287), .A2(n5272), .ZN(n5507) );
  NAND2_X1 U3931 ( .A1(n5508), .A2(n5509), .ZN(n5272) );
  NAND2_X1 U3932 ( .A1(n5280), .A2(n5275), .ZN(n5509) );
  NAND2_X1 U3933 ( .A1(n5510), .A2(n5511), .ZN(n5280) );
  NAND2_X1 U3934 ( .A1(n5512), .A2(n5513), .ZN(n5511) );
  XOR2_X1 U3935 ( .A(KEYINPUT53), .B(n5514), .Z(n5510) );
  NOR2_X1 U3936 ( .A1(n5512), .A2(n5513), .ZN(n5514) );
  NAND2_X1 U3937 ( .A1(n4822), .A2(n5513), .ZN(n5508) );
  NOR3_X1 U3938 ( .A1(n5329), .A2(n5326), .A3(n5328), .ZN(n5324) );
  NAND2_X1 U3939 ( .A1(n5347), .A2(n5515), .ZN(n5328) );
  NAND2_X1 U3940 ( .A1(n5516), .A2(G2253), .ZN(n5515) );
  INV_X1 U3941 ( .A(n5444), .ZN(n5404) );
  NAND2_X1 U3942 ( .A1(n5231), .A2(n5225), .ZN(n5444) );
  NOR2_X1 U3943 ( .A1(n5162), .A2(n5193), .ZN(n5225) );
  INV_X1 U3944 ( .A(n5191), .ZN(n5193) );
  XOR2_X1 U3945 ( .A(n5517), .B(KEYINPUT78), .Z(n5191) );
  NAND3_X1 U3946 ( .A1(n5171), .A2(n5166), .A3(n5167), .ZN(n5162) );
  NOR2_X1 U3947 ( .A1(n5190), .A2(n5189), .ZN(n5167) );
  NAND2_X1 U3948 ( .A1(n5518), .A2(n5519), .ZN(n5190) );
  NAND2_X1 U3949 ( .A1(n4745), .A2(n5520), .ZN(n5519) );
  NAND2_X1 U3950 ( .A1(n5521), .A2(n5522), .ZN(n5520) );
  NAND2_X1 U3951 ( .A1(n5523), .A2(n5521), .ZN(n5518) );
  INV_X1 U3952 ( .A(KEYINPUT31), .ZN(n5521) );
  INV_X1 U3953 ( .A(n5204), .ZN(n5171) );
  NAND2_X1 U3954 ( .A1(n5524), .A2(n5525), .ZN(n5204) );
  NAND2_X1 U3955 ( .A1(G1480), .A2(n5526), .ZN(n5525) );
  NAND2_X1 U3956 ( .A1(KEYINPUT5), .A2(n4744), .ZN(n5526) );
  NAND2_X1 U3957 ( .A1(KEYINPUT5), .A2(n5201), .ZN(n5524) );
  NAND2_X1 U3958 ( .A1(n5527), .A2(n5528), .ZN(G264) );
  NAND2_X1 U3959 ( .A1(n5529), .A2(n5530), .ZN(n5528) );
  NAND2_X1 U3960 ( .A1(n5531), .A2(n5532), .ZN(G252) );
  NAND2_X1 U3961 ( .A1(n5533), .A2(n5534), .ZN(n5532) );
  NAND2_X1 U3962 ( .A1(n5535), .A2(n5536), .ZN(n5534) );
  NAND2_X1 U3963 ( .A1(KEYINPUT23), .A2(n5537), .ZN(n5536) );
  INV_X1 U3964 ( .A(n5538), .ZN(n5533) );
  NAND2_X1 U3965 ( .A1(n5539), .A2(n5540), .ZN(n5531) );
  INV_X1 U3966 ( .A(KEYINPUT23), .ZN(n5540) );
  NAND2_X1 U3967 ( .A1(n5527), .A2(n5541), .ZN(G249) );
  NAND2_X1 U3968 ( .A1(n5542), .A2(n5530), .ZN(n5541) );
  XOR2_X1 U3969 ( .A(n5529), .B(KEYINPUT86), .Z(n5542) );
  NAND2_X1 U3970 ( .A1(n5543), .A2(n5544), .ZN(n5529) );
  NAND2_X1 U3971 ( .A1(n5545), .A2(n5546), .ZN(n5544) );
  NAND2_X1 U3972 ( .A1(n5547), .A2(n5548), .ZN(n5546) );
  NAND2_X1 U3973 ( .A1(n4662), .A2(n5549), .ZN(n5548) );
  OR2_X1 U3974 ( .A1(n5550), .A2(n4539), .ZN(n5549) );
  NAND2_X1 U3975 ( .A1(n5550), .A2(n4539), .ZN(n5547) );
  NAND2_X1 U3976 ( .A1(n5551), .A2(n5552), .ZN(n5550) );
  NAND2_X1 U3977 ( .A1(n5553), .A2(n5554), .ZN(n5552) );
  INV_X1 U3978 ( .A(n5555), .ZN(n5553) );
  NAND2_X1 U3979 ( .A1(n4673), .A2(n4532), .ZN(n5551) );
  XOR2_X1 U3980 ( .A(n5556), .B(KEYINPUT82), .Z(n5543) );
  NAND2_X1 U3981 ( .A1(n4663), .A2(n4540), .ZN(n5556) );
  AND2_X1 U3982 ( .A1(n5557), .A2(n5558), .ZN(n5527) );
  NAND4_X1 U3983 ( .A1(n5559), .A2(n5530), .A3(n5560), .A4(n5561), .ZN(n5558) );
  NOR4_X1 U3984 ( .A1(n5554), .A2(n5562), .A3(n5555), .A4(n5563), .ZN(n5561) );
  XNOR2_X1 U3985 ( .A(n4662), .B(n4539), .ZN(n5563) );
  NAND2_X1 U3986 ( .A1(n4541), .A2(n5564), .ZN(n4539) );
  NAND2_X1 U3987 ( .A1(G167), .A2(n4543), .ZN(n5564) );
  NAND2_X1 U3988 ( .A1(n5565), .A2(n5566), .ZN(n4662) );
  NAND2_X1 U3989 ( .A1(G18), .A2(n5567), .ZN(n5566) );
  NAND2_X1 U3990 ( .A1(G112), .A2(n4527), .ZN(n5565) );
  NAND2_X1 U3991 ( .A1(n5568), .A2(n5569), .ZN(n5555) );
  OR2_X1 U3992 ( .A1(n4675), .A2(n4535), .ZN(n5569) );
  XOR2_X1 U3993 ( .A(n4532), .B(n4673), .Z(n5568) );
  NAND2_X1 U3994 ( .A1(n5570), .A2(n5571), .ZN(n4673) );
  OR2_X1 U3995 ( .A1(n4527), .A2(G106), .ZN(n5571) );
  NAND2_X1 U3996 ( .A1(G87), .A2(n4527), .ZN(n5570) );
  NAND2_X1 U3997 ( .A1(n5572), .A2(n5573), .ZN(n4532) );
  OR2_X1 U3998 ( .A1(n5574), .A2(n4536), .ZN(n5573) );
  NOR2_X1 U3999 ( .A1(G168), .A2(n5575), .ZN(n5574) );
  INV_X1 U4000 ( .A(KEYINPUT64), .ZN(n5575) );
  NAND2_X1 U4001 ( .A1(KEYINPUT64), .A2(n4545), .ZN(n5572) );
  INV_X1 U4002 ( .A(n5545), .ZN(n5562) );
  XOR2_X1 U4003 ( .A(n4663), .B(n4540), .Z(n5545) );
  NAND2_X1 U4004 ( .A1(n4541), .A2(n5576), .ZN(n4540) );
  NAND2_X1 U4005 ( .A1(G166), .A2(n4543), .ZN(n5576) );
  NAND2_X1 U4006 ( .A1(n5577), .A2(n5578), .ZN(n4663) );
  NAND2_X1 U4007 ( .A1(G88), .A2(n4527), .ZN(n5578) );
  NAND2_X1 U4008 ( .A1(n5579), .A2(G18), .ZN(n5577) );
  XOR2_X1 U4009 ( .A(KEYINPUT104), .B(G1486), .Z(n5579) );
  NAND2_X1 U4010 ( .A1(n5580), .A2(n5581), .ZN(n5554) );
  NAND2_X1 U4011 ( .A1(n4679), .A2(n4543), .ZN(n5581) );
  NAND2_X1 U4012 ( .A1(n4675), .A2(n4535), .ZN(n5580) );
  NAND2_X1 U4013 ( .A1(n4541), .A2(n5582), .ZN(n4535) );
  NAND2_X1 U4014 ( .A1(G169), .A2(n4543), .ZN(n5582) );
  NAND2_X1 U4015 ( .A1(n5583), .A2(n5584), .ZN(n4675) );
  NAND2_X1 U4016 ( .A1(G18), .A2(n5522), .ZN(n5584) );
  INV_X1 U4017 ( .A(G1469), .ZN(n5522) );
  NAND2_X1 U4018 ( .A1(G111), .A2(n4527), .ZN(n5583) );
  NOR2_X1 U4019 ( .A1(n5585), .A2(n5586), .ZN(n5560) );
  NOR2_X1 U4020 ( .A1(n4563), .A2(n4704), .ZN(n5586) );
  NOR2_X1 U4021 ( .A1(n4679), .A2(n4543), .ZN(n5585) );
  NAND2_X1 U4022 ( .A1(n5587), .A2(n5588), .ZN(n4679) );
  OR2_X1 U4023 ( .A1(n4527), .A2(G1462), .ZN(n5588) );
  NAND2_X1 U4024 ( .A1(G113), .A2(n4527), .ZN(n5587) );
  NAND3_X1 U4025 ( .A1(n5589), .A2(n5590), .A3(n5591), .ZN(n5530) );
  NAND2_X1 U4026 ( .A1(n5592), .A2(n5593), .ZN(n5591) );
  NAND2_X1 U4027 ( .A1(KEYINPUT46), .A2(n5594), .ZN(n5592) );
  NAND2_X1 U4028 ( .A1(G1455), .A2(n5595), .ZN(n5589) );
  NAND2_X1 U4029 ( .A1(n5594), .A2(n5596), .ZN(n5595) );
  NAND2_X1 U4030 ( .A1(KEYINPUT46), .A2(G4528), .ZN(n5596) );
  INV_X1 U4031 ( .A(G2204), .ZN(n5594) );
  NAND3_X1 U4032 ( .A1(n5597), .A2(n5598), .A3(n5599), .ZN(n5559) );
  NAND2_X1 U4033 ( .A1(n4705), .A2(n4554), .ZN(n5599) );
  NAND3_X1 U4034 ( .A1(n5600), .A2(n5601), .A3(n5602), .ZN(n5598) );
  OR2_X1 U4035 ( .A1(n4554), .A2(n4705), .ZN(n5602) );
  AND2_X1 U4036 ( .A1(n5603), .A2(n5604), .ZN(n4705) );
  NAND2_X1 U4037 ( .A1(G18), .A2(G2253), .ZN(n5604) );
  OR2_X1 U4038 ( .A1(G18), .A2(G109), .ZN(n5603) );
  NAND2_X1 U4039 ( .A1(n5605), .A2(n5606), .ZN(n4554) );
  NAND3_X1 U4040 ( .A1(n5607), .A2(n4543), .A3(n5608), .ZN(n5606) );
  OR2_X1 U4041 ( .A1(n4545), .A2(G174), .ZN(n5607) );
  OR3_X1 U4042 ( .A1(n4536), .A2(G174), .A3(n5608), .ZN(n5605) );
  INV_X1 U4043 ( .A(KEYINPUT0), .ZN(n5608) );
  NAND3_X1 U4044 ( .A1(n5609), .A2(n5610), .A3(n5611), .ZN(n5601) );
  NAND2_X1 U4045 ( .A1(n4687), .A2(n4559), .ZN(n5611) );
  NAND3_X1 U4046 ( .A1(n4688), .A2(n5612), .A3(KEYINPUT6), .ZN(n5610) );
  NAND2_X1 U4047 ( .A1(n4558), .A2(n5613), .ZN(n5609) );
  OR2_X1 U4048 ( .A1(n5612), .A2(n4688), .ZN(n5613) );
  NAND2_X1 U4049 ( .A1(n5614), .A2(n5615), .ZN(n4688) );
  OR2_X1 U4050 ( .A1(n4527), .A2(G2239), .ZN(n5615) );
  NAND2_X1 U4051 ( .A1(G63), .A2(n4527), .ZN(n5614) );
  NAND3_X1 U4052 ( .A1(n5616), .A2(n5617), .A3(n5618), .ZN(n5612) );
  NAND2_X1 U4053 ( .A1(n4701), .A2(n4571), .ZN(n5618) );
  NAND2_X1 U4054 ( .A1(n5619), .A2(n5620), .ZN(n5617) );
  XOR2_X1 U4055 ( .A(n5621), .B(KEYINPUT57), .Z(n5619) );
  NAND4_X1 U4056 ( .A1(n5622), .A2(n5623), .A3(n5624), .A4(n5625), .ZN(n5621) );
  NOR2_X1 U4057 ( .A1(n4550), .A2(n4694), .ZN(n5625) );
  INV_X1 U4058 ( .A(n5626), .ZN(n4550) );
  NAND2_X1 U4059 ( .A1(n4703), .A2(n4566), .ZN(n5624) );
  OR2_X1 U4060 ( .A1(n4700), .A2(n4555), .ZN(n5622) );
  NAND2_X1 U4061 ( .A1(n5627), .A2(n5623), .ZN(n5616) );
  OR2_X1 U4062 ( .A1(n4701), .A2(n4571), .ZN(n5623) );
  NAND2_X1 U4063 ( .A1(n4541), .A2(n5628), .ZN(n4571) );
  NAND2_X1 U4064 ( .A1(G177), .A2(n4543), .ZN(n5628) );
  NAND2_X1 U4065 ( .A1(n5629), .A2(n5630), .ZN(n4701) );
  NAND2_X1 U4066 ( .A1(G64), .A2(n4527), .ZN(n5630) );
  NAND2_X1 U4067 ( .A1(n5631), .A2(G18), .ZN(n5629) );
  XOR2_X1 U4068 ( .A(KEYINPUT16), .B(G2236), .Z(n5631) );
  NAND2_X1 U4069 ( .A1(n5632), .A2(n5633), .ZN(n5627) );
  NAND2_X1 U4070 ( .A1(n4555), .A2(n5634), .ZN(n5633) );
  OR2_X1 U4071 ( .A1(n5635), .A2(n4700), .ZN(n5634) );
  NAND2_X1 U4072 ( .A1(n5636), .A2(n5637), .ZN(n4555) );
  NAND2_X1 U4073 ( .A1(G178), .A2(G18), .ZN(n5636) );
  NAND2_X1 U4074 ( .A1(n4700), .A2(n5635), .ZN(n5632) );
  NAND2_X1 U4075 ( .A1(n5638), .A2(n5639), .ZN(n5635) );
  NAND2_X1 U4076 ( .A1(n5640), .A2(n5641), .ZN(n5639) );
  OR2_X1 U4077 ( .A1(n5642), .A2(n5643), .ZN(n5641) );
  INV_X1 U4078 ( .A(n4703), .ZN(n5640) );
  NAND2_X1 U4079 ( .A1(n5644), .A2(n5645), .ZN(n4703) );
  NAND2_X1 U4080 ( .A1(G2224), .A2(G18), .ZN(n5645) );
  OR2_X1 U4081 ( .A1(G84), .A2(G18), .ZN(n5644) );
  NAND2_X1 U4082 ( .A1(n5643), .A2(n5642), .ZN(n5638) );
  NAND2_X1 U4083 ( .A1(n5646), .A2(n5647), .ZN(n5642) );
  NAND2_X1 U4084 ( .A1(n4702), .A2(n4567), .ZN(n5647) );
  NAND3_X1 U4085 ( .A1(n5620), .A2(n5539), .A3(n5648), .ZN(n5646) );
  XNOR2_X1 U4086 ( .A(n4694), .B(n5626), .ZN(n5648) );
  NAND2_X1 U4087 ( .A1(n5649), .A2(n5650), .ZN(n5626) );
  NAND2_X1 U4088 ( .A1(G147), .A2(n4527), .ZN(n5650) );
  NAND2_X1 U4089 ( .A1(G171), .A2(G18), .ZN(n5649) );
  NAND2_X1 U4090 ( .A1(n5651), .A2(n5652), .ZN(n4694) );
  NAND2_X1 U4091 ( .A1(G2211), .A2(G18), .ZN(n5652) );
  OR2_X1 U4092 ( .A1(G65), .A2(G18), .ZN(n5651) );
  NAND2_X1 U4093 ( .A1(n5535), .A2(n5653), .ZN(n5539) );
  NAND2_X1 U4094 ( .A1(n5537), .A2(n5538), .ZN(n5653) );
  NAND3_X1 U4095 ( .A1(n5654), .A2(n5655), .A3(n5656), .ZN(n5538) );
  NAND2_X1 U4096 ( .A1(n4590), .A2(n4717), .ZN(n5656) );
  NAND4_X1 U4097 ( .A1(n5657), .A2(n5658), .A3(n5659), .A4(n5660), .ZN(n5655) );
  NOR3_X1 U4098 ( .A1(n5661), .A2(n5662), .A3(n5663), .ZN(n5660) );
  NOR2_X1 U4099 ( .A1(n4584), .A2(n4724), .ZN(n5663) );
  NOR2_X1 U4100 ( .A1(n4651), .A2(n5664), .ZN(n5662) );
  NAND2_X1 U4101 ( .A1(n4598), .A2(n5665), .ZN(n5659) );
  NAND2_X1 U4102 ( .A1(n5666), .A2(n5664), .ZN(n5665) );
  NAND2_X1 U4103 ( .A1(n5667), .A2(n5668), .ZN(n5664) );
  NAND2_X1 U4104 ( .A1(n5669), .A2(n5670), .ZN(n5668) );
  NAND2_X1 U4105 ( .A1(n5671), .A2(n5672), .ZN(n5670) );
  NAND3_X1 U4106 ( .A1(n5673), .A2(n5674), .A3(n5675), .ZN(n5672) );
  NAND2_X1 U4107 ( .A1(n4619), .A2(n4644), .ZN(n5675) );
  NAND4_X1 U4108 ( .A1(n5676), .A2(n5677), .A3(n5678), .A4(n5679), .ZN(n5674) );
  NOR2_X1 U4109 ( .A1(n5680), .A2(n5681), .ZN(n5679) );
  NOR2_X1 U4110 ( .A1(n4619), .A2(n4644), .ZN(n5681) );
  NAND2_X1 U4111 ( .A1(n5682), .A2(n5683), .ZN(n4644) );
  OR2_X1 U4112 ( .A1(G53), .A2(G18), .ZN(n5683) );
  NAND2_X1 U4113 ( .A1(G18), .A2(n5684), .ZN(n5682) );
  AND2_X1 U4114 ( .A1(n5685), .A2(n5686), .ZN(n4619) );
  NAND2_X1 U4115 ( .A1(G130), .A2(n4583), .ZN(n5686) );
  NAND2_X1 U4116 ( .A1(G203), .A2(n4586), .ZN(n5685) );
  NOR2_X1 U4117 ( .A1(n4608), .A2(n4647), .ZN(n5680) );
  NAND2_X1 U4118 ( .A1(n5687), .A2(n5688), .ZN(n5678) );
  NAND2_X1 U4119 ( .A1(n5689), .A2(n5690), .ZN(n5687) );
  NAND2_X1 U4120 ( .A1(n5691), .A2(n5692), .ZN(n5690) );
  NAND2_X1 U4121 ( .A1(n5693), .A2(n5694), .ZN(n5691) );
  NAND3_X1 U4122 ( .A1(n4620), .A2(n5695), .A3(n4639), .ZN(n5694) );
  NAND2_X1 U4123 ( .A1(n4646), .A2(n4621), .ZN(n5693) );
  NAND2_X1 U4124 ( .A1(n4645), .A2(n4609), .ZN(n5689) );
  NAND3_X1 U4125 ( .A1(G89), .A2(n5696), .A3(n5697), .ZN(n5677) );
  XOR2_X1 U4126 ( .A(n5698), .B(n4616), .Z(n5697) );
  XOR2_X1 U4127 ( .A(KEYINPUT51), .B(n5699), .Z(n5696) );
  NAND3_X1 U4128 ( .A1(n4616), .A2(n5698), .A3(n5699), .ZN(n5676) );
  AND4_X1 U4129 ( .A1(n5695), .A2(n5700), .A3(n5692), .A4(n5688), .ZN(n5699) );
  NAND2_X1 U4130 ( .A1(n4647), .A2(n4608), .ZN(n5688) );
  AND2_X1 U4131 ( .A1(n5701), .A2(n5702), .ZN(n4608) );
  NAND2_X1 U4132 ( .A1(n5703), .A2(G103), .ZN(n5702) );
  XNOR2_X1 U4133 ( .A(n4586), .B(KEYINPUT108), .ZN(n5703) );
  NAND2_X1 U4134 ( .A1(G204), .A2(n4586), .ZN(n5701) );
  AND2_X1 U4135 ( .A1(n5704), .A2(n5705), .ZN(n4647) );
  NAND2_X1 U4136 ( .A1(G18), .A2(n5706), .ZN(n5705) );
  NAND2_X1 U4137 ( .A1(G73), .A2(n4527), .ZN(n5704) );
  OR2_X1 U4138 ( .A1(n4645), .A2(n4609), .ZN(n5692) );
  NAND2_X1 U4139 ( .A1(n5707), .A2(n5708), .ZN(n4609) );
  NAND2_X1 U4140 ( .A1(G205), .A2(G18), .ZN(n5707) );
  NAND2_X1 U4141 ( .A1(n5709), .A2(n5710), .ZN(n4645) );
  NAND2_X1 U4142 ( .A1(G18), .A2(n5711), .ZN(n5710) );
  NAND2_X1 U4143 ( .A1(G75), .A2(n4527), .ZN(n5709) );
  OR2_X1 U4144 ( .A1(n4639), .A2(n4620), .ZN(n5700) );
  NAND2_X1 U4145 ( .A1(n5712), .A2(n5713), .ZN(n4620) );
  NAND2_X1 U4146 ( .A1(G207), .A2(G18), .ZN(n5712) );
  NAND2_X1 U4147 ( .A1(n5714), .A2(n5715), .ZN(n4639) );
  NAND2_X1 U4148 ( .A1(G18), .A2(n5454), .ZN(n5715) );
  INV_X1 U4149 ( .A(G3705), .ZN(n5454) );
  NAND2_X1 U4150 ( .A1(G74), .A2(n4527), .ZN(n5714) );
  OR2_X1 U4151 ( .A1(n4646), .A2(n4621), .ZN(n5695) );
  NAND2_X1 U4152 ( .A1(n5716), .A2(n5717), .ZN(n4621) );
  NAND2_X1 U4153 ( .A1(G26), .A2(n4527), .ZN(n5717) );
  NAND2_X1 U4154 ( .A1(G206), .A2(G18), .ZN(n5716) );
  NAND2_X1 U4155 ( .A1(n5718), .A2(n5719), .ZN(n4646) );
  NAND2_X1 U4156 ( .A1(G76), .A2(n4527), .ZN(n5719) );
  OR2_X1 U4157 ( .A1(n5720), .A2(n4527), .ZN(n5718) );
  NAND2_X1 U4158 ( .A1(n4527), .A2(n5721), .ZN(n5698) );
  NAND2_X1 U4159 ( .A1(KEYINPUT70), .A2(G70), .ZN(n5721) );
  AND2_X1 U4160 ( .A1(n4615), .A2(n4527), .ZN(n4616) );
  NAND2_X1 U4161 ( .A1(n5722), .A2(n5723), .ZN(n4615) );
  NAND2_X1 U4162 ( .A1(G198), .A2(G18), .ZN(n5722) );
  OR2_X1 U4163 ( .A1(n4650), .A2(n4622), .ZN(n5673) );
  NAND2_X1 U4164 ( .A1(n4650), .A2(n4622), .ZN(n5671) );
  NAND2_X1 U4165 ( .A1(n5724), .A2(n5725), .ZN(n4622) );
  NAND2_X1 U4166 ( .A1(n4583), .A2(G127), .ZN(n5725) );
  NAND2_X1 U4167 ( .A1(G202), .A2(n4586), .ZN(n5724) );
  NAND2_X1 U4168 ( .A1(n5726), .A2(n5727), .ZN(n4650) );
  NAND2_X1 U4169 ( .A1(G18), .A2(n5728), .ZN(n5727) );
  NAND2_X1 U4170 ( .A1(G54), .A2(n4527), .ZN(n5726) );
  XOR2_X1 U4171 ( .A(n4652), .B(n5729), .Z(n5669) );
  XNOR2_X1 U4172 ( .A(KEYINPUT79), .B(n4603), .ZN(n5729) );
  NAND2_X1 U4173 ( .A1(n4652), .A2(n4603), .ZN(n5667) );
  NAND2_X1 U4174 ( .A1(n5730), .A2(n5731), .ZN(n4603) );
  NAND2_X1 U4175 ( .A1(n4583), .A2(G124), .ZN(n5731) );
  NAND2_X1 U4176 ( .A1(G201), .A2(n4586), .ZN(n5730) );
  NAND2_X1 U4177 ( .A1(n5732), .A2(n5733), .ZN(n4652) );
  NAND2_X1 U4178 ( .A1(G18), .A2(n5734), .ZN(n5733) );
  NAND2_X1 U4179 ( .A1(G55), .A2(n4527), .ZN(n5732) );
  XNOR2_X1 U4180 ( .A(KEYINPUT60), .B(n4651), .ZN(n5666) );
  NAND2_X1 U4181 ( .A1(n5735), .A2(n5736), .ZN(n4651) );
  NAND2_X1 U4182 ( .A1(G18), .A2(n5737), .ZN(n5736) );
  NAND2_X1 U4183 ( .A1(G56), .A2(n4527), .ZN(n5735) );
  NAND2_X1 U4184 ( .A1(n5738), .A2(n5739), .ZN(n4598) );
  OR2_X1 U4185 ( .A1(G200), .A2(n4583), .ZN(n5739) );
  OR2_X1 U4186 ( .A1(n4586), .A2(G100), .ZN(n5738) );
  NAND2_X1 U4187 ( .A1(n5740), .A2(n5657), .ZN(n5654) );
  OR2_X1 U4188 ( .A1(n4717), .A2(n4590), .ZN(n5657) );
  NAND2_X1 U4189 ( .A1(n5741), .A2(n5742), .ZN(n4590) );
  NAND2_X1 U4190 ( .A1(G193), .A2(G18), .ZN(n5741) );
  NAND2_X1 U4191 ( .A1(n5743), .A2(n5744), .ZN(n4717) );
  NAND2_X1 U4192 ( .A1(G18), .A2(n5745), .ZN(n5744) );
  XOR2_X1 U4193 ( .A(n5746), .B(KEYINPUT65), .Z(n5743) );
  NAND2_X1 U4194 ( .A1(G80), .A2(n4527), .ZN(n5746) );
  NAND2_X1 U4195 ( .A1(n5747), .A2(n5748), .ZN(n5740) );
  NAND2_X1 U4196 ( .A1(n5749), .A2(n5750), .ZN(n5748) );
  NAND3_X1 U4197 ( .A1(n5751), .A2(n5752), .A3(n5753), .ZN(n5750) );
  NAND2_X1 U4198 ( .A1(n4720), .A2(n4588), .ZN(n5753) );
  NAND3_X1 U4199 ( .A1(n4584), .A2(n5658), .A3(n4724), .ZN(n5752) );
  NAND2_X1 U4200 ( .A1(n5754), .A2(n5755), .ZN(n4724) );
  OR2_X1 U4201 ( .A1(n4527), .A2(G4394), .ZN(n5755) );
  NAND2_X1 U4202 ( .A1(G77), .A2(n4527), .ZN(n5754) );
  OR2_X1 U4203 ( .A1(n4719), .A2(n4579), .ZN(n5658) );
  NAND2_X1 U4204 ( .A1(n5756), .A2(n5757), .ZN(n4584) );
  NAND2_X1 U4205 ( .A1(G118), .A2(n4583), .ZN(n5757) );
  NAND2_X1 U4206 ( .A1(G187), .A2(n4586), .ZN(n5756) );
  NAND2_X1 U4207 ( .A1(n4719), .A2(n4579), .ZN(n5751) );
  NAND2_X1 U4208 ( .A1(n5758), .A2(n5759), .ZN(n4579) );
  NAND2_X1 U4209 ( .A1(n4583), .A2(G97), .ZN(n5759) );
  NAND2_X1 U4210 ( .A1(G196), .A2(n4586), .ZN(n5758) );
  NAND2_X1 U4211 ( .A1(n5760), .A2(n5761), .ZN(n4719) );
  OR2_X1 U4212 ( .A1(n4527), .A2(G4400), .ZN(n5761) );
  NAND2_X1 U4213 ( .A1(G78), .A2(n4527), .ZN(n5760) );
  INV_X1 U4214 ( .A(n5661), .ZN(n5749) );
  NAND2_X1 U4215 ( .A1(n5762), .A2(n5763), .ZN(n5661) );
  OR2_X1 U4216 ( .A1(n4720), .A2(n4588), .ZN(n5763) );
  NAND2_X1 U4217 ( .A1(n5764), .A2(n5765), .ZN(n4588) );
  NAND2_X1 U4218 ( .A1(G94), .A2(n4583), .ZN(n5765) );
  NAND2_X1 U4219 ( .A1(G195), .A2(n4586), .ZN(n5764) );
  NAND2_X1 U4220 ( .A1(n5766), .A2(n5767), .ZN(n4720) );
  NAND2_X1 U4221 ( .A1(G18), .A2(n5768), .ZN(n5767) );
  NAND2_X1 U4222 ( .A1(G59), .A2(n4527), .ZN(n5766) );
  OR2_X1 U4223 ( .A1(n4718), .A2(n4593), .ZN(n5762) );
  NAND2_X1 U4224 ( .A1(n4718), .A2(n4593), .ZN(n5747) );
  NAND2_X1 U4225 ( .A1(n5769), .A2(n5770), .ZN(n4593) );
  NAND2_X1 U4226 ( .A1(G121), .A2(n4583), .ZN(n5770) );
  INV_X1 U4227 ( .A(n4586), .ZN(n4583) );
  NAND2_X1 U4228 ( .A1(G194), .A2(n4586), .ZN(n5769) );
  XOR2_X1 U4229 ( .A(G18), .B(KEYINPUT88), .Z(n4586) );
  NAND2_X1 U4230 ( .A1(n5771), .A2(n5772), .ZN(n4718) );
  NAND2_X1 U4231 ( .A1(G18), .A2(n5773), .ZN(n5772) );
  NAND2_X1 U4232 ( .A1(G81), .A2(n4527), .ZN(n5771) );
  AND3_X1 U4233 ( .A1(n5774), .A2(n5775), .A3(n5776), .ZN(n5537) );
  XOR2_X1 U4234 ( .A(n4732), .B(n5777), .Z(n5776) );
  XNOR2_X1 U4235 ( .A(KEYINPUT15), .B(n4594), .ZN(n5777) );
  AND2_X1 U4236 ( .A1(n5778), .A2(n5779), .ZN(n5535) );
  NAND2_X1 U4237 ( .A1(n5780), .A2(n5775), .ZN(n5779) );
  OR2_X1 U4238 ( .A1(n4729), .A2(n4572), .ZN(n5775) );
  NAND2_X1 U4239 ( .A1(n5781), .A2(n5782), .ZN(n5780) );
  NAND2_X1 U4240 ( .A1(n5774), .A2(n5783), .ZN(n5782) );
  NAND2_X1 U4241 ( .A1(n5784), .A2(n5785), .ZN(n5783) );
  NAND2_X1 U4242 ( .A1(n4732), .A2(n4594), .ZN(n5785) );
  NAND2_X1 U4243 ( .A1(n5786), .A2(n5787), .ZN(n4594) );
  NAND2_X1 U4244 ( .A1(G192), .A2(G18), .ZN(n5786) );
  NAND2_X1 U4245 ( .A1(n5788), .A2(n5789), .ZN(n4732) );
  NAND2_X1 U4246 ( .A1(G18), .A2(n5472), .ZN(n5789) );
  NAND2_X1 U4247 ( .A1(G79), .A2(n4527), .ZN(n5788) );
  NAND2_X1 U4248 ( .A1(n4731), .A2(n4596), .ZN(n5784) );
  AND2_X1 U4249 ( .A1(n5790), .A2(n5791), .ZN(n5774) );
  OR2_X1 U4250 ( .A1(n4731), .A2(n4596), .ZN(n5791) );
  NAND2_X1 U4251 ( .A1(n5792), .A2(n5793), .ZN(n4596) );
  NAND2_X1 U4252 ( .A1(G191), .A2(G18), .ZN(n5792) );
  NAND2_X1 U4253 ( .A1(n5794), .A2(n5795), .ZN(n4731) );
  NAND2_X1 U4254 ( .A1(G18), .A2(n4510), .ZN(n5795) );
  NAND2_X1 U4255 ( .A1(G60), .A2(n4527), .ZN(n5794) );
  OR2_X1 U4256 ( .A1(n4730), .A2(n4595), .ZN(n5790) );
  NAND2_X1 U4257 ( .A1(n4730), .A2(n4595), .ZN(n5781) );
  NAND2_X1 U4258 ( .A1(n5796), .A2(n5797), .ZN(n4595) );
  NAND2_X1 U4259 ( .A1(G190), .A2(G18), .ZN(n5796) );
  NAND2_X1 U4260 ( .A1(n5798), .A2(n5799), .ZN(n4730) );
  NAND2_X1 U4261 ( .A1(G61), .A2(n4527), .ZN(n5799) );
  NAND2_X1 U4262 ( .A1(G18), .A2(n5494), .ZN(n5798) );
  NAND2_X1 U4263 ( .A1(n4729), .A2(n4572), .ZN(n5778) );
  NAND2_X1 U4264 ( .A1(n5800), .A2(n5801), .ZN(n4572) );
  NAND2_X1 U4265 ( .A1(G189), .A2(G18), .ZN(n5800) );
  NAND2_X1 U4266 ( .A1(n5802), .A2(n5803), .ZN(n4729) );
  NAND2_X1 U4267 ( .A1(G18), .A2(n5804), .ZN(n5803) );
  NAND2_X1 U4268 ( .A1(G62), .A2(n4527), .ZN(n5802) );
  XOR2_X1 U4269 ( .A(n4702), .B(n4567), .Z(n5620) );
  NAND2_X1 U4270 ( .A1(n5805), .A2(n5806), .ZN(n4567) );
  NAND2_X1 U4271 ( .A1(G138), .A2(n4527), .ZN(n5806) );
  NAND2_X1 U4272 ( .A1(G180), .A2(G18), .ZN(n5805) );
  NAND2_X1 U4273 ( .A1(n5807), .A2(n5808), .ZN(n4702) );
  OR2_X1 U4274 ( .A1(n4527), .A2(G2218), .ZN(n5808) );
  NAND2_X1 U4275 ( .A1(G83), .A2(n4527), .ZN(n5807) );
  INV_X1 U4276 ( .A(n4566), .ZN(n5643) );
  NAND2_X1 U4277 ( .A1(n5809), .A2(n5810), .ZN(n4566) );
  OR2_X1 U4278 ( .A1(G179), .A2(n4527), .ZN(n5810) );
  NAND2_X1 U4279 ( .A1(n5811), .A2(n5812), .ZN(n4700) );
  NAND2_X1 U4280 ( .A1(G18), .A2(n5513), .ZN(n5812) );
  NAND2_X1 U4281 ( .A1(G85), .A2(n4527), .ZN(n5811) );
  AND2_X1 U4282 ( .A1(n4543), .A2(n5813), .ZN(n4558) );
  OR2_X1 U4283 ( .A1(G176), .A2(n4545), .ZN(n5813) );
  OR2_X1 U4284 ( .A1(n4687), .A2(n4559), .ZN(n5600) );
  NAND2_X1 U4285 ( .A1(n4541), .A2(n5814), .ZN(n4559) );
  NAND2_X1 U4286 ( .A1(G175), .A2(n4543), .ZN(n5814) );
  NAND2_X1 U4287 ( .A1(n5815), .A2(n5816), .ZN(n4687) );
  OR2_X1 U4288 ( .A1(n4527), .A2(G2247), .ZN(n5816) );
  NAND2_X1 U4289 ( .A1(G86), .A2(n4527), .ZN(n5815) );
  NAND2_X1 U4290 ( .A1(n4704), .A2(n4563), .ZN(n5597) );
  NAND2_X1 U4291 ( .A1(n5817), .A2(n5818), .ZN(n4563) );
  OR2_X1 U4292 ( .A1(n5819), .A2(n4536), .ZN(n5818) );
  NAND2_X1 U4293 ( .A1(G18), .A2(n4543), .ZN(n4536) );
  NOR2_X1 U4294 ( .A1(G173), .A2(KEYINPUT33), .ZN(n5819) );
  OR2_X1 U4295 ( .A1(n4541), .A2(KEYINPUT33), .ZN(n5817) );
  NAND2_X1 U4296 ( .A1(n5820), .A2(n5821), .ZN(n4704) );
  NAND2_X1 U4297 ( .A1(G18), .A2(n5822), .ZN(n5821) );
  NAND2_X1 U4298 ( .A1(G110), .A2(n4527), .ZN(n5820) );
  NAND2_X1 U4299 ( .A1(G38), .A2(n5823), .ZN(n5557) );
  OR4_X1 U4300 ( .A1(n5593), .A2(G1455), .A3(G2204), .A4(KEYINPUT46), .ZN(n5823) );
  INV_X1 U4301 ( .A(G4528), .ZN(n5593) );
  NAND2_X1 U4302 ( .A1(n5414), .A2(n5824), .ZN(G246) );
  NAND2_X1 U4303 ( .A1(n5231), .A2(n5825), .ZN(n5824) );
  NAND2_X1 U4304 ( .A1(n5416), .A2(n5826), .ZN(n5825) );
  NAND2_X1 U4305 ( .A1(n5418), .A2(n5827), .ZN(n5826) );
  NAND2_X1 U4306 ( .A1(n5419), .A2(n5828), .ZN(n5827) );
  NAND2_X1 U4307 ( .A1(n5424), .A2(n5355), .ZN(n5828) );
  OR2_X1 U4308 ( .A1(n5425), .A2(n5423), .ZN(n5355) );
  AND4_X1 U4309 ( .A1(n5079), .A2(n5136), .A3(n5139), .A4(n5829), .ZN(n5423) );
  NAND2_X1 U4310 ( .A1(n5144), .A2(n5830), .ZN(n5829) );
  NAND2_X1 U4311 ( .A1(n5146), .A2(n5147), .ZN(n5830) );
  NAND3_X1 U4312 ( .A1(n5831), .A2(n5450), .A3(n5447), .ZN(n5147) );
  AND2_X1 U4313 ( .A1(n5832), .A2(n5833), .ZN(n5447) );
  NAND2_X1 U4314 ( .A1(n4881), .A2(n4899), .ZN(n5833) );
  NAND2_X1 U4315 ( .A1(n4959), .A2(n5834), .ZN(n4899) );
  NAND2_X1 U4316 ( .A1(n4854), .A2(n4960), .ZN(n5834) );
  INV_X1 U4317 ( .A(n4889), .ZN(n4960) );
  NAND2_X1 U4318 ( .A1(n4809), .A2(n5711), .ZN(n4959) );
  INV_X1 U4319 ( .A(G3717), .ZN(n5711) );
  NAND2_X1 U4320 ( .A1(n4808), .A2(n5706), .ZN(n5832) );
  INV_X1 U4321 ( .A(G3723), .ZN(n5706) );
  NAND2_X1 U4322 ( .A1(n4870), .A2(n5443), .ZN(n5450) );
  INV_X1 U4323 ( .A(n5835), .ZN(n5443) );
  NAND2_X1 U4324 ( .A1(n5451), .A2(n4948), .ZN(n5831) );
  NOR2_X1 U4325 ( .A1(n4851), .A2(n5835), .ZN(n5451) );
  AND2_X1 U4326 ( .A1(n5061), .A2(n5836), .ZN(n5144) );
  NAND2_X1 U4327 ( .A1(n4947), .A2(n4984), .ZN(n5836) );
  NAND2_X1 U4328 ( .A1(n5455), .A2(n5837), .ZN(n4984) );
  NAND2_X1 U4329 ( .A1(n5457), .A2(n4976), .ZN(n5837) );
  NAND2_X1 U4330 ( .A1(n5458), .A2(n5838), .ZN(n4976) );
  NAND2_X1 U4331 ( .A1(n4916), .A2(n4968), .ZN(n5838) );
  NAND2_X1 U4332 ( .A1(n4790), .A2(n5728), .ZN(n5458) );
  NAND2_X1 U4333 ( .A1(n4788), .A2(n5734), .ZN(n5455) );
  NAND2_X1 U4334 ( .A1(n5463), .A2(n5839), .ZN(n5425) );
  NAND2_X1 U4335 ( .A1(n5079), .A2(n5840), .ZN(n5839) );
  NAND2_X1 U4336 ( .A1(n5132), .A2(n5841), .ZN(n5840) );
  NAND2_X1 U4337 ( .A1(n5136), .A2(n5842), .ZN(n5841) );
  NAND2_X1 U4338 ( .A1(n5137), .A2(n5843), .ZN(n5842) );
  NAND3_X1 U4339 ( .A1(n5148), .A2(n5139), .A3(n5146), .ZN(n5843) );
  AND2_X1 U4340 ( .A1(n4947), .A2(n4983), .ZN(n5146) );
  NOR3_X1 U4341 ( .A1(n4925), .A2(n5460), .A3(n4923), .ZN(n4983) );
  NAND2_X1 U4342 ( .A1(n4918), .A2(n4939), .ZN(n4923) );
  NAND2_X1 U4343 ( .A1(n4786), .A2(n5684), .ZN(n4939) );
  INV_X1 U4344 ( .A(n4916), .ZN(n4918) );
  NOR2_X1 U4345 ( .A1(n5684), .A2(n4786), .ZN(n4916) );
  AND2_X1 U4346 ( .A1(n5844), .A2(n5845), .ZN(n4786) );
  NAND2_X1 U4347 ( .A1(G130), .A2(n4527), .ZN(n5845) );
  NAND2_X1 U4348 ( .A1(G234), .A2(G18), .ZN(n5844) );
  XOR2_X1 U4349 ( .A(KEYINPUT36), .B(G3729), .Z(n5684) );
  INV_X1 U4350 ( .A(n4968), .ZN(n5460) );
  XOR2_X1 U4351 ( .A(n4790), .B(n5728), .Z(n4968) );
  INV_X1 U4352 ( .A(G3737), .ZN(n5728) );
  AND2_X1 U4353 ( .A1(n5846), .A2(n5847), .ZN(n4790) );
  OR2_X1 U4354 ( .A1(G233), .A2(n4527), .ZN(n5847) );
  OR2_X1 U4355 ( .A1(G127), .A2(G18), .ZN(n5846) );
  INV_X1 U4356 ( .A(n5457), .ZN(n4925) );
  XOR2_X1 U4357 ( .A(n4788), .B(n5734), .Z(n5457) );
  INV_X1 U4358 ( .A(G3743), .ZN(n5734) );
  AND2_X1 U4359 ( .A1(n5848), .A2(n5849), .ZN(n4788) );
  OR2_X1 U4360 ( .A1(G232), .A2(n4527), .ZN(n5849) );
  OR2_X1 U4361 ( .A1(G124), .A2(G18), .ZN(n5848) );
  INV_X1 U4362 ( .A(n4915), .ZN(n4947) );
  NAND2_X1 U4363 ( .A1(n5061), .A2(n5850), .ZN(n4915) );
  OR2_X1 U4364 ( .A1(n5737), .A2(n4787), .ZN(n5850) );
  NAND2_X1 U4365 ( .A1(n4787), .A2(n5737), .ZN(n5061) );
  INV_X1 U4366 ( .A(G3749), .ZN(n5737) );
  NAND2_X1 U4367 ( .A1(n5851), .A2(n5852), .ZN(n4787) );
  NAND2_X1 U4368 ( .A1(G100), .A2(n4527), .ZN(n5852) );
  NAND2_X1 U4369 ( .A1(G231), .A2(G18), .ZN(n5851) );
  AND4_X1 U4370 ( .A1(n5096), .A2(n5436), .A3(n5093), .A4(n5095), .ZN(n5139) );
  AND2_X1 U4371 ( .A1(n5086), .A2(n5011), .ZN(n5096) );
  NAND2_X1 U4372 ( .A1(G4394), .A2(n4764), .ZN(n5011) );
  INV_X1 U4373 ( .A(n5019), .ZN(n5086) );
  NOR2_X1 U4374 ( .A1(n4962), .A2(n5835), .ZN(n5148) );
  NAND2_X1 U4375 ( .A1(n4892), .A2(n4881), .ZN(n5835) );
  INV_X1 U4376 ( .A(n4880), .ZN(n4881) );
  XOR2_X1 U4377 ( .A(G3723), .B(n4808), .Z(n4880) );
  NAND2_X1 U4378 ( .A1(n5853), .A2(n5854), .ZN(n4808) );
  NAND2_X1 U4379 ( .A1(G103), .A2(n4527), .ZN(n5854) );
  NAND2_X1 U4380 ( .A1(G235), .A2(G18), .ZN(n5853) );
  NOR2_X1 U4381 ( .A1(n4866), .A2(n4889), .ZN(n4892) );
  XOR2_X1 U4382 ( .A(G3717), .B(n4809), .Z(n4889) );
  NAND2_X1 U4383 ( .A1(n5855), .A2(n5708), .ZN(n4809) );
  NAND2_X1 U4384 ( .A1(G23), .A2(n4527), .ZN(n5708) );
  NAND2_X1 U4385 ( .A1(G236), .A2(G18), .ZN(n5855) );
  NAND2_X1 U4386 ( .A1(n4954), .A2(n5856), .ZN(n4866) );
  NAND2_X1 U4387 ( .A1(n4804), .A2(n5720), .ZN(n5856) );
  INV_X1 U4388 ( .A(n4854), .ZN(n4954) );
  NOR2_X1 U4389 ( .A1(n5720), .A2(n4804), .ZN(n4854) );
  NAND2_X1 U4390 ( .A1(n5857), .A2(n5858), .ZN(n4804) );
  OR2_X1 U4391 ( .A1(G237), .A2(n4527), .ZN(n5858) );
  OR2_X1 U4392 ( .A1(G18), .A2(G26), .ZN(n5857) );
  XOR2_X1 U4393 ( .A(KEYINPUT59), .B(G3711), .Z(n5720) );
  NAND3_X1 U4394 ( .A1(n4882), .A2(n4948), .A3(G4526), .ZN(n4962) );
  AND2_X1 U4395 ( .A1(n5859), .A2(n4869), .ZN(n4948) );
  INV_X1 U4396 ( .A(n4870), .ZN(n4869) );
  NOR2_X1 U4397 ( .A1(n4807), .A2(G3705), .ZN(n4870) );
  NAND2_X1 U4398 ( .A1(G3705), .A2(n4807), .ZN(n5859) );
  INV_X1 U4399 ( .A(n4805), .ZN(n4807) );
  NAND2_X1 U4400 ( .A1(n5860), .A2(n5713), .ZN(n4805) );
  NAND2_X1 U4401 ( .A1(G29), .A2(n4527), .ZN(n5713) );
  NAND2_X1 U4402 ( .A1(G238), .A2(G18), .ZN(n5860) );
  NOR2_X1 U4403 ( .A1(n4861), .A2(n4902), .ZN(n4882) );
  INV_X1 U4404 ( .A(n4851), .ZN(n4902) );
  NAND3_X1 U4405 ( .A1(n4527), .A2(n4630), .A3(n4798), .ZN(n4851) );
  NOR3_X1 U4406 ( .A1(n4798), .A2(G18), .A3(n4630), .ZN(n4861) );
  INV_X1 U4407 ( .A(G3701), .ZN(n4630) );
  NAND2_X1 U4408 ( .A1(n5861), .A2(n5723), .ZN(n4798) );
  NAND2_X1 U4409 ( .A1(G41), .A2(n4527), .ZN(n5723) );
  NAND2_X1 U4410 ( .A1(G229), .A2(G18), .ZN(n5861) );
  AND2_X1 U4411 ( .A1(n5470), .A2(n5469), .ZN(n5137) );
  NAND2_X1 U4412 ( .A1(n5436), .A2(n5014), .ZN(n5469) );
  NAND2_X1 U4413 ( .A1(n5097), .A2(n5862), .ZN(n5014) );
  NAND2_X1 U4414 ( .A1(n5093), .A2(n5024), .ZN(n5862) );
  NAND3_X1 U4415 ( .A1(n5863), .A2(n5864), .A3(n5865), .ZN(n5024) );
  NAND2_X1 U4416 ( .A1(n4771), .A2(n5768), .ZN(n5865) );
  INV_X1 U4417 ( .A(G4405), .ZN(n5768) );
  NAND2_X1 U4418 ( .A1(n5019), .A2(n5095), .ZN(n5864) );
  NOR2_X1 U4419 ( .A1(n5081), .A2(n5034), .ZN(n5095) );
  NAND2_X1 U4420 ( .A1(n5026), .A2(n5866), .ZN(n5081) );
  NAND2_X1 U4421 ( .A1(G4400), .A2(n4768), .ZN(n5866) );
  INV_X1 U4422 ( .A(n5867), .ZN(n5026) );
  NOR2_X1 U4423 ( .A1(n4764), .A2(G4394), .ZN(n5019) );
  AND2_X1 U4424 ( .A1(n5868), .A2(n5869), .ZN(n4764) );
  NAND2_X1 U4425 ( .A1(G118), .A2(n4527), .ZN(n5869) );
  NAND2_X1 U4426 ( .A1(G217), .A2(G18), .ZN(n5868) );
  NAND2_X1 U4427 ( .A1(n5867), .A2(n4998), .ZN(n5863) );
  INV_X1 U4428 ( .A(n5034), .ZN(n4998) );
  XOR2_X1 U4429 ( .A(G4405), .B(n4771), .Z(n5034) );
  NAND2_X1 U4430 ( .A1(n5870), .A2(n5871), .ZN(n4771) );
  NAND2_X1 U4431 ( .A1(G94), .A2(n4527), .ZN(n5871) );
  NAND2_X1 U4432 ( .A1(G225), .A2(G18), .ZN(n5870) );
  NOR2_X1 U4433 ( .A1(n4768), .A2(G4400), .ZN(n5867) );
  NAND2_X1 U4434 ( .A1(n5872), .A2(n5873), .ZN(n4768) );
  OR2_X1 U4435 ( .A1(G226), .A2(n4527), .ZN(n5873) );
  OR2_X1 U4436 ( .A1(G18), .A2(G97), .ZN(n5872) );
  INV_X1 U4437 ( .A(n5032), .ZN(n5093) );
  NAND2_X1 U4438 ( .A1(n5874), .A2(n5097), .ZN(n5032) );
  OR2_X1 U4439 ( .A1(n5773), .A2(n4769), .ZN(n5874) );
  NAND2_X1 U4440 ( .A1(n4769), .A2(n5773), .ZN(n5097) );
  INV_X1 U4441 ( .A(G4410), .ZN(n5773) );
  NAND2_X1 U4442 ( .A1(n5875), .A2(n5876), .ZN(n4769) );
  NAND2_X1 U4443 ( .A1(G121), .A2(n4527), .ZN(n5876) );
  NAND2_X1 U4444 ( .A1(G224), .A2(G18), .ZN(n5875) );
  INV_X1 U4445 ( .A(n5008), .ZN(n5436) );
  NAND2_X1 U4446 ( .A1(n5470), .A2(n5877), .ZN(n5008) );
  OR2_X1 U4447 ( .A1(n5745), .A2(n4757), .ZN(n5877) );
  NAND2_X1 U4448 ( .A1(n4757), .A2(n5745), .ZN(n5470) );
  INV_X1 U4449 ( .A(G4415), .ZN(n5745) );
  NAND2_X1 U4450 ( .A1(n5878), .A2(n5742), .ZN(n4757) );
  NAND2_X1 U4451 ( .A1(G47), .A2(n4527), .ZN(n5742) );
  NAND2_X1 U4452 ( .A1(G223), .A2(G18), .ZN(n5878) );
  NOR2_X1 U4453 ( .A1(n5122), .A2(n5117), .ZN(n5136) );
  OR2_X1 U4454 ( .A1(n5100), .A2(n5106), .ZN(n5122) );
  XOR2_X1 U4455 ( .A(n5879), .B(n5472), .Z(n5100) );
  INV_X1 U4456 ( .A(G4420), .ZN(n5472) );
  NAND2_X1 U4457 ( .A1(KEYINPUT97), .A2(n5880), .ZN(n5879) );
  XNOR2_X1 U4458 ( .A(n4776), .B(KEYINPUT58), .ZN(n5880) );
  INV_X1 U4459 ( .A(n5133), .ZN(n5132) );
  NAND2_X1 U4460 ( .A1(n5495), .A2(n5881), .ZN(n5133) );
  OR2_X1 U4461 ( .A1(n5117), .A2(n5118), .ZN(n5881) );
  AND2_X1 U4462 ( .A1(n5112), .A2(n5476), .ZN(n5118) );
  OR2_X1 U4463 ( .A1(n5106), .A2(n5077), .ZN(n5112) );
  INV_X1 U4464 ( .A(n5072), .ZN(n5077) );
  NOR2_X1 U4465 ( .A1(n4776), .A2(G4420), .ZN(n5072) );
  INV_X1 U4466 ( .A(n4780), .ZN(n4776) );
  NAND2_X1 U4467 ( .A1(n5882), .A2(n5787), .ZN(n4780) );
  NAND2_X1 U4468 ( .A1(G35), .A2(n4527), .ZN(n5787) );
  NAND2_X1 U4469 ( .A1(G222), .A2(G18), .ZN(n5882) );
  NAND2_X1 U4470 ( .A1(n5476), .A2(n5883), .ZN(n5106) );
  NAND2_X1 U4471 ( .A1(n4782), .A2(G4427), .ZN(n5883) );
  INV_X1 U4472 ( .A(n4779), .ZN(n4782) );
  NAND2_X1 U4473 ( .A1(n4779), .A2(n4510), .ZN(n5476) );
  INV_X1 U4474 ( .A(G4427), .ZN(n4510) );
  NAND2_X1 U4475 ( .A1(n5884), .A2(n5793), .ZN(n4779) );
  NAND2_X1 U4476 ( .A1(G32), .A2(n4527), .ZN(n5793) );
  NAND2_X1 U4477 ( .A1(G221), .A2(G18), .ZN(n5884) );
  NAND2_X1 U4478 ( .A1(n5495), .A2(n5885), .ZN(n5117) );
  OR2_X1 U4479 ( .A1(n4765), .A2(n5494), .ZN(n5885) );
  NAND2_X1 U4480 ( .A1(n5494), .A2(n4765), .ZN(n5495) );
  NAND2_X1 U4481 ( .A1(n5886), .A2(n5797), .ZN(n4765) );
  NAND2_X1 U4482 ( .A1(G50), .A2(n4527), .ZN(n5797) );
  NAND2_X1 U4483 ( .A1(G220), .A2(G18), .ZN(n5886) );
  XOR2_X1 U4484 ( .A(KEYINPUT37), .B(G4432), .Z(n5494) );
  INV_X1 U4485 ( .A(n5126), .ZN(n5079) );
  NAND2_X1 U4486 ( .A1(n5463), .A2(n5887), .ZN(n5126) );
  OR2_X1 U4487 ( .A1(n5804), .A2(n4758), .ZN(n5887) );
  NAND2_X1 U4488 ( .A1(n4758), .A2(n5804), .ZN(n5463) );
  INV_X1 U4489 ( .A(G4437), .ZN(n5804) );
  NAND2_X1 U4490 ( .A1(n5888), .A2(n5801), .ZN(n4758) );
  NAND2_X1 U4491 ( .A1(G66), .A2(n4527), .ZN(n5801) );
  NAND2_X1 U4492 ( .A1(G219), .A2(G18), .ZN(n5888) );
  AND4_X1 U4493 ( .A1(n5297), .A2(n5889), .A3(n5362), .A4(n5287), .ZN(n5424) );
  AND2_X1 U4494 ( .A1(n5292), .A2(n5281), .ZN(n5297) );
  AND2_X1 U4495 ( .A1(n5271), .A2(n5286), .ZN(n5292) );
  AND2_X1 U4496 ( .A1(n5890), .A2(n5353), .ZN(n5271) );
  INV_X1 U4497 ( .A(n5270), .ZN(n5353) );
  NAND2_X1 U4498 ( .A1(G2211), .A2(n4821), .ZN(n5890) );
  AND3_X1 U4499 ( .A1(n5891), .A2(n5892), .A3(n5496), .ZN(n5419) );
  NAND2_X1 U4500 ( .A1(n4832), .A2(n5822), .ZN(n5496) );
  INV_X1 U4501 ( .A(G2256), .ZN(n5822) );
  NAND2_X1 U4502 ( .A1(n5889), .A2(n5399), .ZN(n5892) );
  NAND3_X1 U4503 ( .A1(n5893), .A2(n5894), .A3(n5506), .ZN(n5399) );
  NAND2_X1 U4504 ( .A1(n5287), .A2(n5895), .ZN(n5894) );
  NAND2_X1 U4505 ( .A1(n5896), .A2(n5897), .ZN(n5895) );
  OR2_X1 U4506 ( .A1(n5366), .A2(KEYINPUT10), .ZN(n5897) );
  NAND2_X1 U4507 ( .A1(n5362), .A2(n5275), .ZN(n5896) );
  NAND2_X1 U4508 ( .A1(n5898), .A2(n5899), .ZN(n5275) );
  NAND2_X1 U4509 ( .A1(n5281), .A2(n5360), .ZN(n5899) );
  NAND2_X1 U4510 ( .A1(n5293), .A2(n5900), .ZN(n5360) );
  NAND2_X1 U4511 ( .A1(n5270), .A2(n5286), .ZN(n5900) );
  INV_X1 U4512 ( .A(n5352), .ZN(n5286) );
  NAND2_X1 U4513 ( .A1(n5293), .A2(n5901), .ZN(n5352) );
  NAND2_X1 U4514 ( .A1(G2218), .A2(n4829), .ZN(n5901) );
  NOR2_X1 U4515 ( .A1(n4821), .A2(G2211), .ZN(n5270) );
  NAND2_X1 U4516 ( .A1(n5902), .A2(n5903), .ZN(n4821) );
  OR2_X1 U4517 ( .A1(G151), .A2(n4527), .ZN(n5903) );
  OR2_X1 U4518 ( .A1(G147), .A2(G18), .ZN(n5902) );
  OR2_X1 U4519 ( .A1(n4829), .A2(G2218), .ZN(n5293) );
  NAND2_X1 U4520 ( .A1(n5904), .A2(n5905), .ZN(n4829) );
  OR2_X1 U4521 ( .A1(G160), .A2(n4527), .ZN(n5905) );
  OR2_X1 U4522 ( .A1(G138), .A2(G18), .ZN(n5904) );
  XOR2_X1 U4523 ( .A(n4830), .B(G2224), .Z(n5281) );
  OR2_X1 U4524 ( .A1(n4830), .A2(G2224), .ZN(n5898) );
  NAND2_X1 U4525 ( .A1(n5809), .A2(n5906), .ZN(n4830) );
  OR2_X1 U4526 ( .A1(G159), .A2(n4527), .ZN(n5906) );
  NAND2_X1 U4527 ( .A1(n5907), .A2(n4527), .ZN(n5809) );
  INV_X1 U4528 ( .A(G144), .ZN(n5907) );
  XNOR2_X1 U4529 ( .A(n5513), .B(n5512), .ZN(n5362) );
  INV_X1 U4530 ( .A(n5364), .ZN(n5287) );
  NAND3_X1 U4531 ( .A1(KEYINPUT10), .A2(n5908), .A3(n5364), .ZN(n5893) );
  NAND2_X1 U4532 ( .A1(n5506), .A2(n5909), .ZN(n5364) );
  NAND2_X1 U4533 ( .A1(G2236), .A2(n4831), .ZN(n5909) );
  OR2_X1 U4534 ( .A1(n4831), .A2(G2236), .ZN(n5506) );
  NAND2_X1 U4535 ( .A1(n5910), .A2(n4543), .ZN(n4831) );
  OR2_X1 U4536 ( .A1(G157), .A2(n4545), .ZN(n5910) );
  INV_X1 U4537 ( .A(n5366), .ZN(n5908) );
  NAND2_X1 U4538 ( .A1(n5911), .A2(n5513), .ZN(n5366) );
  INV_X1 U4539 ( .A(G2230), .ZN(n5513) );
  XNOR2_X1 U4540 ( .A(n5512), .B(KEYINPUT96), .ZN(n5911) );
  INV_X1 U4541 ( .A(n4822), .ZN(n5512) );
  NAND2_X1 U4542 ( .A1(n5912), .A2(n5637), .ZN(n4822) );
  NAND2_X1 U4543 ( .A1(G135), .A2(n4527), .ZN(n5637) );
  NAND2_X1 U4544 ( .A1(G158), .A2(G18), .ZN(n5912) );
  NOR4_X1 U4545 ( .A1(n5329), .A2(n5395), .A3(n5326), .A4(n5393), .ZN(n5889) );
  INV_X1 U4546 ( .A(n5391), .ZN(n5393) );
  INV_X1 U4547 ( .A(n5327), .ZN(n5329) );
  NOR2_X1 U4548 ( .A1(n5309), .A2(n5350), .ZN(n5327) );
  INV_X1 U4549 ( .A(n5312), .ZN(n5309) );
  NAND2_X1 U4550 ( .A1(G2239), .A2(n4814), .ZN(n5312) );
  NAND2_X1 U4551 ( .A1(n5391), .A2(n5398), .ZN(n5891) );
  NAND2_X1 U4552 ( .A1(n5347), .A2(n5913), .ZN(n5398) );
  NAND2_X1 U4553 ( .A1(n5381), .A2(n5310), .ZN(n5913) );
  NAND2_X1 U4554 ( .A1(n5504), .A2(n5377), .ZN(n5310) );
  NAND2_X1 U4555 ( .A1(n5350), .A2(n5330), .ZN(n5377) );
  INV_X1 U4556 ( .A(n5326), .ZN(n5330) );
  NAND2_X1 U4557 ( .A1(n5504), .A2(n5914), .ZN(n5326) );
  NAND2_X1 U4558 ( .A1(G2247), .A2(n4825), .ZN(n5914) );
  NOR2_X1 U4559 ( .A1(n4814), .A2(G2239), .ZN(n5350) );
  NAND2_X1 U4560 ( .A1(n5915), .A2(n4543), .ZN(n4814) );
  OR2_X1 U4561 ( .A1(G156), .A2(n4545), .ZN(n5915) );
  INV_X1 U4562 ( .A(n5505), .ZN(n5504) );
  NOR2_X1 U4563 ( .A1(n4825), .A2(G2247), .ZN(n5505) );
  NAND2_X1 U4564 ( .A1(n5916), .A2(n4543), .ZN(n4825) );
  OR2_X1 U4565 ( .A1(n4545), .A2(G155), .ZN(n5916) );
  INV_X1 U4566 ( .A(n5395), .ZN(n5381) );
  NAND2_X1 U4567 ( .A1(n5917), .A2(n5918), .ZN(n5395) );
  NAND2_X1 U4568 ( .A1(G2253), .A2(n5919), .ZN(n5918) );
  NAND2_X1 U4569 ( .A1(KEYINPUT90), .A2(n4815), .ZN(n5919) );
  NAND2_X1 U4570 ( .A1(n5920), .A2(KEYINPUT90), .ZN(n5917) );
  INV_X1 U4571 ( .A(n5920), .ZN(n5347) );
  NOR2_X1 U4572 ( .A1(n5516), .A2(G2253), .ZN(n5920) );
  INV_X1 U4573 ( .A(n4815), .ZN(n5516) );
  NAND2_X1 U4574 ( .A1(n4541), .A2(n5921), .ZN(n4815) );
  NAND2_X1 U4575 ( .A1(G154), .A2(n4543), .ZN(n5921) );
  XOR2_X1 U4576 ( .A(n5305), .B(KEYINPUT119), .Z(n5391) );
  XNOR2_X1 U4577 ( .A(G2256), .B(n4832), .ZN(n5305) );
  NAND2_X1 U4578 ( .A1(n4541), .A2(n5922), .ZN(n4832) );
  NAND2_X1 U4579 ( .A1(G153), .A2(n4543), .ZN(n5922) );
  AND3_X1 U4580 ( .A1(n5517), .A2(n5923), .A3(n5192), .ZN(n5418) );
  INV_X1 U4581 ( .A(n5189), .ZN(n5192) );
  NAND2_X1 U4582 ( .A1(n5197), .A2(n5170), .ZN(n5189) );
  NAND2_X1 U4583 ( .A1(G1462), .A2(n5924), .ZN(n5170) );
  INV_X1 U4584 ( .A(n5215), .ZN(n5197) );
  AND2_X1 U4585 ( .A1(n5925), .A2(n5926), .ZN(n5416) );
  NAND2_X1 U4586 ( .A1(n5517), .A2(n5927), .ZN(n5926) );
  NAND3_X1 U4587 ( .A1(n5928), .A2(n5929), .A3(n5930), .ZN(n5927) );
  XNOR2_X1 U4588 ( .A(KEYINPUT21), .B(n5248), .ZN(n5930) );
  NAND2_X1 U4589 ( .A1(n5215), .A2(n5923), .ZN(n5929) );
  NOR3_X1 U4590 ( .A1(n5173), .A2(n5250), .A3(n5252), .ZN(n5923) );
  NAND2_X1 U4591 ( .A1(n5931), .A2(n5195), .ZN(n5252) );
  INV_X1 U4592 ( .A(n5523), .ZN(n5195) );
  NAND2_X1 U4593 ( .A1(G1469), .A2(n4745), .ZN(n5931) );
  INV_X1 U4594 ( .A(n5244), .ZN(n5250) );
  NOR2_X1 U4595 ( .A1(n5924), .A2(G1462), .ZN(n5215) );
  AND2_X1 U4596 ( .A1(n4541), .A2(n5932), .ZN(n5924) );
  NAND2_X1 U4597 ( .A1(G209), .A2(n4543), .ZN(n5932) );
  NAND2_X1 U4598 ( .A1(n5213), .A2(n5244), .ZN(n5928) );
  NAND2_X1 U4599 ( .A1(n5933), .A2(n5934), .ZN(n5244) );
  NAND3_X1 U4600 ( .A1(n5248), .A2(n5567), .A3(KEYINPUT54), .ZN(n5934) );
  NAND2_X1 U4601 ( .A1(n5935), .A2(n4744), .ZN(n5933) );
  NAND2_X1 U4602 ( .A1(n5201), .A2(KEYINPUT54), .ZN(n5935) );
  INV_X1 U4603 ( .A(n5248), .ZN(n5201) );
  NAND2_X1 U4604 ( .A1(n5567), .A2(n4744), .ZN(n5248) );
  NAND2_X1 U4605 ( .A1(n4541), .A2(n5936), .ZN(n4744) );
  NAND2_X1 U4606 ( .A1(G214), .A2(n4543), .ZN(n5936) );
  INV_X1 U4607 ( .A(G1480), .ZN(n5567) );
  NAND2_X1 U4608 ( .A1(n5205), .A2(n5937), .ZN(n5213) );
  NAND2_X1 U4609 ( .A1(n5523), .A2(n5166), .ZN(n5937) );
  INV_X1 U4610 ( .A(n5173), .ZN(n5166) );
  NAND2_X1 U4611 ( .A1(n5205), .A2(n5938), .ZN(n5173) );
  NAND2_X1 U4612 ( .A1(G106), .A2(n4749), .ZN(n5938) );
  NOR2_X1 U4613 ( .A1(G1469), .A2(n4745), .ZN(n5523) );
  AND2_X1 U4614 ( .A1(n4541), .A2(n5939), .ZN(n4745) );
  NAND2_X1 U4615 ( .A1(G216), .A2(n4543), .ZN(n5939) );
  INV_X1 U4616 ( .A(n4545), .ZN(n4541) );
  OR2_X1 U4617 ( .A1(n4749), .A2(G106), .ZN(n5205) );
  NAND2_X1 U4618 ( .A1(n5940), .A2(n4543), .ZN(n4749) );
  OR2_X1 U4619 ( .A1(n4545), .A2(G215), .ZN(n5940) );
  INV_X1 U4620 ( .A(n5255), .ZN(n5517) );
  NAND2_X1 U4621 ( .A1(n5429), .A2(n5941), .ZN(n5255) );
  NAND2_X1 U4622 ( .A1(G1486), .A2(n4748), .ZN(n5941) );
  XNOR2_X1 U4623 ( .A(KEYINPUT50), .B(n5429), .ZN(n5925) );
  OR2_X1 U4624 ( .A1(n4748), .A2(G1486), .ZN(n5429) );
  NAND2_X1 U4625 ( .A1(n4543), .A2(n5942), .ZN(n4748) );
  OR2_X1 U4626 ( .A1(G213), .A2(n4545), .ZN(n5942) );
  NOR2_X1 U4627 ( .A1(G18), .A2(n4746), .ZN(n4545) );
  INV_X1 U4628 ( .A(n4543), .ZN(n4746) );
  NAND2_X1 U4629 ( .A1(G9), .A2(G12), .ZN(n4543) );
  NOR2_X1 U4630 ( .A1(n4514), .A2(n4511), .ZN(n5231) );
  NAND2_X1 U4631 ( .A1(n5233), .A2(n4515), .ZN(n4511) );
  NAND2_X1 U4632 ( .A1(n5943), .A2(n5590), .ZN(n5233) );
  XNOR2_X1 U4633 ( .A(KEYINPUT18), .B(n5944), .ZN(n5943) );
  XOR2_X1 U4634 ( .A(n5945), .B(n5590), .Z(n4514) );
  INV_X1 U4635 ( .A(G38), .ZN(n5590) );
  INV_X1 U4636 ( .A(n5234), .ZN(n5414) );
  NAND2_X1 U4637 ( .A1(n4515), .A2(n5946), .ZN(n5234) );
  NAND2_X1 U4638 ( .A1(G38), .A2(n5945), .ZN(n5946) );
  NAND2_X1 U4639 ( .A1(G1496), .A2(G4528), .ZN(n5945) );
  NAND2_X1 U4640 ( .A1(n5947), .A2(G38), .ZN(n4515) );
  XOR2_X1 U4641 ( .A(n5944), .B(KEYINPUT18), .Z(n5947) );
  NAND2_X1 U4642 ( .A1(G4528), .A2(G1492), .ZN(n5944) );
endmodule

