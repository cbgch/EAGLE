//Key = 0001000001110001101010111111010111010111001110101011001000011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315;

XOR2_X1 U726 ( .A(G107), .B(n1001), .Z(G9) );
NOR2_X1 U727 ( .A1(KEYINPUT5), .A2(n1002), .ZN(n1001) );
NOR2_X1 U728 ( .A1(n1003), .A2(n1004), .ZN(G75) );
XOR2_X1 U729 ( .A(KEYINPUT30), .B(n1005), .Z(n1004) );
NOR3_X1 U730 ( .A1(n1006), .A2(G953), .A3(G952), .ZN(n1005) );
NOR4_X1 U731 ( .A1(n1007), .A2(n1008), .A3(n1006), .A4(n1009), .ZN(n1003) );
NOR2_X1 U732 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR2_X1 U733 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U734 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
INV_X1 U735 ( .A(n1016), .ZN(n1015) );
NOR2_X1 U736 ( .A1(n1017), .A2(n1018), .ZN(n1014) );
NOR2_X1 U737 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U738 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U739 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U741 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U742 ( .A1(n1029), .A2(n1030), .ZN(n1021) );
NOR2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR3_X1 U745 ( .A1(n1030), .A2(n1035), .A3(n1024), .ZN(n1017) );
NOR2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR4_X1 U747 ( .A1(n1038), .A2(n1024), .A3(n1020), .A4(n1030), .ZN(n1012) );
INV_X1 U748 ( .A(n1039), .ZN(n1030) );
NOR2_X1 U749 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
XOR2_X1 U750 ( .A(KEYINPUT53), .B(n1042), .Z(n1041) );
NOR2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
AND4_X1 U752 ( .A1(n1016), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1006) );
NOR4_X1 U753 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
XNOR2_X1 U755 ( .A(G475), .B(KEYINPUT55), .ZN(n1053) );
INV_X1 U756 ( .A(n1054), .ZN(n1052) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1046) );
XNOR2_X1 U758 ( .A(n1057), .B(n1058), .ZN(n1056) );
XOR2_X1 U759 ( .A(KEYINPUT44), .B(G478), .Z(n1058) );
INV_X1 U760 ( .A(G952), .ZN(n1008) );
NAND2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1007) );
XNOR2_X1 U762 ( .A(G953), .B(KEYINPUT40), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1061), .A2(n1062), .ZN(G72) );
NAND3_X1 U764 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
INV_X1 U765 ( .A(n1066), .ZN(n1065) );
XOR2_X1 U766 ( .A(n1067), .B(KEYINPUT63), .Z(n1061) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1068), .ZN(n1067) );
NAND2_X1 U768 ( .A1(n1063), .A2(n1064), .ZN(n1068) );
NAND2_X1 U769 ( .A1(G900), .A2(G227), .ZN(n1064) );
XNOR2_X1 U770 ( .A(KEYINPUT0), .B(n1069), .ZN(n1063) );
NAND2_X1 U771 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
NAND2_X1 U772 ( .A1(n1072), .A2(n1069), .ZN(n1071) );
XOR2_X1 U773 ( .A(n1073), .B(n1074), .Z(n1072) );
NAND2_X1 U774 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
INV_X1 U775 ( .A(n1077), .ZN(n1076) );
XOR2_X1 U776 ( .A(n1078), .B(KEYINPUT24), .Z(n1075) );
NAND3_X1 U777 ( .A1(G900), .A2(n1074), .A3(G953), .ZN(n1070) );
XNOR2_X1 U778 ( .A(n1079), .B(n1080), .ZN(n1074) );
XNOR2_X1 U779 ( .A(n1081), .B(n1082), .ZN(n1080) );
XNOR2_X1 U780 ( .A(n1083), .B(n1084), .ZN(n1079) );
XOR2_X1 U781 ( .A(KEYINPUT43), .B(n1085), .Z(n1084) );
XOR2_X1 U782 ( .A(n1086), .B(n1087), .Z(G69) );
NAND2_X1 U783 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1088) );
NAND2_X1 U785 ( .A1(KEYINPUT9), .A2(n1089), .ZN(n1086) );
XOR2_X1 U786 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U788 ( .A(KEYINPUT29), .B(n1069), .ZN(n1092) );
NAND2_X1 U789 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
NAND2_X1 U790 ( .A1(G953), .A2(n1096), .ZN(n1095) );
XOR2_X1 U791 ( .A(n1097), .B(n1098), .Z(n1094) );
XOR2_X1 U792 ( .A(KEYINPUT49), .B(n1099), .Z(n1098) );
NOR2_X1 U793 ( .A1(n1100), .A2(n1101), .ZN(G66) );
XOR2_X1 U794 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR2_X1 U796 ( .A1(n1100), .A2(n1106), .ZN(G63) );
XOR2_X1 U797 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U798 ( .A1(KEYINPUT46), .A2(n1109), .ZN(n1108) );
NAND2_X1 U799 ( .A1(n1104), .A2(G478), .ZN(n1107) );
NOR2_X1 U800 ( .A1(n1100), .A2(n1110), .ZN(G60) );
XOR2_X1 U801 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND2_X1 U802 ( .A1(n1104), .A2(G475), .ZN(n1111) );
XNOR2_X1 U803 ( .A(G104), .B(n1113), .ZN(G6) );
NAND4_X1 U804 ( .A1(n1114), .A2(n1037), .A3(n1115), .A4(n1045), .ZN(n1113) );
XNOR2_X1 U805 ( .A(n1040), .B(KEYINPUT42), .ZN(n1114) );
NOR2_X1 U806 ( .A1(n1100), .A2(n1116), .ZN(G57) );
XOR2_X1 U807 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U808 ( .A(n1119), .B(n1120), .Z(n1118) );
AND2_X1 U809 ( .A1(G472), .A2(n1104), .ZN(n1119) );
NOR3_X1 U810 ( .A1(n1121), .A2(n1100), .A3(n1122), .ZN(G54) );
NOR4_X1 U811 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1122) );
NOR2_X1 U812 ( .A1(KEYINPUT27), .A2(n1127), .ZN(n1124) );
NOR2_X1 U813 ( .A1(n1128), .A2(n1129), .ZN(n1123) );
INV_X1 U814 ( .A(KEYINPUT27), .ZN(n1129) );
NOR2_X1 U815 ( .A1(n1128), .A2(n1130), .ZN(n1121) );
NOR2_X1 U816 ( .A1(n1125), .A2(n1126), .ZN(n1130) );
INV_X1 U817 ( .A(n1104), .ZN(n1126) );
NOR2_X1 U818 ( .A1(n1127), .A2(n1131), .ZN(n1128) );
INV_X1 U819 ( .A(KEYINPUT51), .ZN(n1131) );
XNOR2_X1 U820 ( .A(n1132), .B(n1133), .ZN(n1127) );
XNOR2_X1 U821 ( .A(n1134), .B(n1135), .ZN(n1132) );
NAND2_X1 U822 ( .A1(KEYINPUT31), .A2(n1136), .ZN(n1135) );
XOR2_X1 U823 ( .A(KEYINPUT28), .B(n1137), .Z(n1136) );
NAND2_X1 U824 ( .A1(n1138), .A2(KEYINPUT33), .ZN(n1134) );
XOR2_X1 U825 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U826 ( .A1(KEYINPUT35), .A2(n1141), .ZN(n1139) );
NOR2_X1 U827 ( .A1(n1100), .A2(n1142), .ZN(G51) );
XOR2_X1 U828 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U829 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U830 ( .A1(KEYINPUT32), .A2(n1147), .ZN(n1145) );
XOR2_X1 U831 ( .A(n1148), .B(KEYINPUT54), .Z(n1143) );
NAND2_X1 U832 ( .A1(n1104), .A2(n1149), .ZN(n1148) );
NOR2_X1 U833 ( .A1(n1150), .A2(n1060), .ZN(n1104) );
NOR3_X1 U834 ( .A1(n1077), .A2(n1078), .A3(n1093), .ZN(n1060) );
NAND4_X1 U835 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1093) );
NOR4_X1 U836 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
INV_X1 U837 ( .A(n1002), .ZN(n1155) );
NAND4_X1 U838 ( .A1(n1040), .A2(n1115), .A3(n1036), .A4(n1045), .ZN(n1002) );
OR2_X1 U839 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
NAND3_X1 U840 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1152) );
XNOR2_X1 U841 ( .A(n1026), .B(KEYINPUT60), .ZN(n1163) );
XNOR2_X1 U842 ( .A(KEYINPUT23), .B(n1164), .ZN(n1162) );
INV_X1 U843 ( .A(n1165), .ZN(n1161) );
NAND3_X1 U844 ( .A1(n1045), .A2(n1166), .A3(n1115), .ZN(n1151) );
NAND2_X1 U845 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND3_X1 U846 ( .A1(n1169), .A2(n1170), .A3(n1016), .ZN(n1168) );
NAND2_X1 U847 ( .A1(n1037), .A2(n1040), .ZN(n1167) );
NAND4_X1 U848 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1078) );
NAND3_X1 U849 ( .A1(n1016), .A2(n1026), .A3(n1175), .ZN(n1171) );
NAND4_X1 U850 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1077) );
NOR2_X1 U851 ( .A1(n1069), .A2(G952), .ZN(n1100) );
NAND2_X1 U852 ( .A1(n1180), .A2(n1181), .ZN(G48) );
NAND2_X1 U853 ( .A1(G146), .A2(n1176), .ZN(n1181) );
XOR2_X1 U854 ( .A(KEYINPUT25), .B(n1182), .Z(n1180) );
NOR2_X1 U855 ( .A1(G146), .A2(n1176), .ZN(n1182) );
NAND3_X1 U856 ( .A1(n1037), .A2(n1026), .A3(n1183), .ZN(n1176) );
XNOR2_X1 U857 ( .A(G143), .B(n1177), .ZN(G45) );
NAND4_X1 U858 ( .A1(n1169), .A2(n1184), .A3(n1026), .A4(n1170), .ZN(n1177) );
XNOR2_X1 U859 ( .A(G140), .B(n1178), .ZN(G42) );
NAND3_X1 U860 ( .A1(n1039), .A2(n1040), .A3(n1175), .ZN(n1178) );
XNOR2_X1 U861 ( .A(G137), .B(n1179), .ZN(G39) );
NAND3_X1 U862 ( .A1(n1039), .A2(n1185), .A3(n1183), .ZN(n1179) );
XNOR2_X1 U863 ( .A(G134), .B(n1172), .ZN(G36) );
NAND3_X1 U864 ( .A1(n1039), .A2(n1036), .A3(n1184), .ZN(n1172) );
XNOR2_X1 U865 ( .A(G131), .B(n1173), .ZN(G33) );
NAND3_X1 U866 ( .A1(n1039), .A2(n1037), .A3(n1184), .ZN(n1173) );
AND3_X1 U867 ( .A1(n1040), .A2(n1186), .A3(n1032), .ZN(n1184) );
NOR2_X1 U868 ( .A1(n1027), .A2(n1055), .ZN(n1039) );
INV_X1 U869 ( .A(n1028), .ZN(n1055) );
XNOR2_X1 U870 ( .A(G128), .B(n1174), .ZN(G30) );
NAND3_X1 U871 ( .A1(n1036), .A2(n1026), .A3(n1183), .ZN(n1174) );
AND4_X1 U872 ( .A1(n1040), .A2(n1187), .A3(n1034), .A4(n1186), .ZN(n1183) );
XNOR2_X1 U873 ( .A(n1188), .B(n1189), .ZN(G3) );
NOR2_X1 U874 ( .A1(n1190), .A2(n1160), .ZN(n1189) );
XOR2_X1 U875 ( .A(n1159), .B(KEYINPUT57), .Z(n1190) );
NAND4_X1 U876 ( .A1(n1032), .A2(n1185), .A3(n1040), .A4(n1164), .ZN(n1159) );
XNOR2_X1 U877 ( .A(G125), .B(n1191), .ZN(G27) );
NAND4_X1 U878 ( .A1(KEYINPUT3), .A2(n1175), .A3(n1016), .A4(n1026), .ZN(n1191) );
AND4_X1 U879 ( .A1(n1192), .A2(n1037), .A3(n1187), .A4(n1186), .ZN(n1175) );
NAND2_X1 U880 ( .A1(n1011), .A2(n1193), .ZN(n1186) );
NAND4_X1 U881 ( .A1(G953), .A2(G902), .A3(n1194), .A4(n1195), .ZN(n1193) );
INV_X1 U882 ( .A(G900), .ZN(n1195) );
XNOR2_X1 U883 ( .A(G122), .B(n1196), .ZN(G24) );
NAND4_X1 U884 ( .A1(n1197), .A2(n1198), .A3(n1016), .A4(n1199), .ZN(n1196) );
NOR3_X1 U885 ( .A1(n1024), .A2(n1200), .A3(n1201), .ZN(n1199) );
INV_X1 U886 ( .A(n1045), .ZN(n1024) );
NOR2_X1 U887 ( .A1(n1034), .A2(n1187), .ZN(n1045) );
NAND2_X1 U888 ( .A1(KEYINPUT18), .A2(n1202), .ZN(n1198) );
NAND2_X1 U889 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
INV_X1 U890 ( .A(KEYINPUT18), .ZN(n1204) );
NAND2_X1 U891 ( .A1(n1160), .A2(n1164), .ZN(n1203) );
XNOR2_X1 U892 ( .A(n1205), .B(n1158), .ZN(G21) );
AND3_X1 U893 ( .A1(n1016), .A2(n1034), .A3(n1206), .ZN(n1158) );
XOR2_X1 U894 ( .A(G116), .B(n1157), .Z(G18) );
AND4_X1 U895 ( .A1(n1032), .A2(n1016), .A3(n1115), .A4(n1036), .ZN(n1157) );
NOR2_X1 U896 ( .A1(n1170), .A2(n1201), .ZN(n1036) );
INV_X1 U897 ( .A(n1202), .ZN(n1115) );
XOR2_X1 U898 ( .A(n1207), .B(n1208), .Z(G15) );
NOR2_X1 U899 ( .A1(n1202), .A2(n1165), .ZN(n1208) );
NAND3_X1 U900 ( .A1(n1032), .A2(n1016), .A3(n1037), .ZN(n1165) );
AND2_X1 U901 ( .A1(n1209), .A2(n1170), .ZN(n1037) );
XNOR2_X1 U902 ( .A(KEYINPUT13), .B(n1169), .ZN(n1209) );
NOR2_X1 U903 ( .A1(n1043), .A2(n1210), .ZN(n1016) );
INV_X1 U904 ( .A(n1044), .ZN(n1210) );
NOR2_X1 U905 ( .A1(n1187), .A2(n1192), .ZN(n1032) );
NOR2_X1 U906 ( .A1(KEYINPUT19), .A2(n1211), .ZN(n1207) );
INV_X1 U907 ( .A(G113), .ZN(n1211) );
XOR2_X1 U908 ( .A(n1156), .B(n1212), .Z(G12) );
XNOR2_X1 U909 ( .A(KEYINPUT1), .B(n1213), .ZN(n1212) );
AND3_X1 U910 ( .A1(n1192), .A2(n1040), .A3(n1206), .ZN(n1156) );
NOR3_X1 U911 ( .A1(n1202), .A2(n1033), .A3(n1020), .ZN(n1206) );
INV_X1 U912 ( .A(n1185), .ZN(n1020) );
NOR2_X1 U913 ( .A1(n1170), .A2(n1169), .ZN(n1185) );
INV_X1 U914 ( .A(n1201), .ZN(n1169) );
XOR2_X1 U915 ( .A(G478), .B(n1214), .Z(n1201) );
NOR2_X1 U916 ( .A1(n1057), .A2(KEYINPUT45), .ZN(n1214) );
NOR2_X1 U917 ( .A1(n1109), .A2(G902), .ZN(n1057) );
AND2_X1 U918 ( .A1(n1215), .A2(n1216), .ZN(n1109) );
NAND4_X1 U919 ( .A1(G234), .A2(n1069), .A3(G217), .A4(n1217), .ZN(n1216) );
INV_X1 U920 ( .A(n1218), .ZN(n1217) );
NAND2_X1 U921 ( .A1(n1218), .A2(n1219), .ZN(n1215) );
NAND3_X1 U922 ( .A1(G234), .A2(n1069), .A3(G217), .ZN(n1219) );
XNOR2_X1 U923 ( .A(n1220), .B(n1221), .ZN(n1218) );
NOR2_X1 U924 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR2_X1 U925 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XNOR2_X1 U926 ( .A(KEYINPUT59), .B(n1226), .ZN(n1224) );
NOR2_X1 U927 ( .A1(G143), .A2(n1227), .ZN(n1222) );
XNOR2_X1 U928 ( .A(G128), .B(n1228), .ZN(n1227) );
XNOR2_X1 U929 ( .A(KEYINPUT8), .B(KEYINPUT58), .ZN(n1228) );
XNOR2_X1 U930 ( .A(n1229), .B(n1230), .ZN(n1220) );
INV_X1 U931 ( .A(G134), .ZN(n1230) );
NAND2_X1 U932 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
NAND2_X1 U933 ( .A1(G107), .A2(n1233), .ZN(n1232) );
XOR2_X1 U934 ( .A(KEYINPUT37), .B(n1234), .Z(n1231) );
NOR2_X1 U935 ( .A1(G107), .A2(n1233), .ZN(n1234) );
XNOR2_X1 U936 ( .A(n1235), .B(n1236), .ZN(n1233) );
NOR2_X1 U937 ( .A1(KEYINPUT36), .A2(n1237), .ZN(n1236) );
INV_X1 U938 ( .A(n1200), .ZN(n1170) );
NOR2_X1 U939 ( .A1(n1048), .A2(n1238), .ZN(n1200) );
AND2_X1 U940 ( .A1(G475), .A2(n1054), .ZN(n1238) );
NOR2_X1 U941 ( .A1(n1054), .A2(G475), .ZN(n1048) );
NAND2_X1 U942 ( .A1(n1112), .A2(n1150), .ZN(n1054) );
XNOR2_X1 U943 ( .A(n1239), .B(n1240), .ZN(n1112) );
XOR2_X1 U944 ( .A(n1241), .B(n1242), .Z(n1240) );
XNOR2_X1 U945 ( .A(n1237), .B(G113), .ZN(n1242) );
INV_X1 U946 ( .A(G122), .ZN(n1237) );
XNOR2_X1 U947 ( .A(KEYINPUT26), .B(n1225), .ZN(n1241) );
XOR2_X1 U948 ( .A(n1243), .B(n1244), .Z(n1239) );
XNOR2_X1 U949 ( .A(G104), .B(n1245), .ZN(n1244) );
NAND2_X1 U950 ( .A1(KEYINPUT38), .A2(n1081), .ZN(n1245) );
XOR2_X1 U951 ( .A(n1246), .B(n1247), .Z(n1243) );
NAND4_X1 U952 ( .A1(KEYINPUT16), .A2(G214), .A3(n1248), .A4(n1069), .ZN(n1246) );
INV_X1 U953 ( .A(n1187), .ZN(n1033) );
XNOR2_X1 U954 ( .A(n1249), .B(n1105), .ZN(n1187) );
AND2_X1 U955 ( .A1(G217), .A2(n1250), .ZN(n1105) );
NAND2_X1 U956 ( .A1(n1103), .A2(n1150), .ZN(n1249) );
XNOR2_X1 U957 ( .A(n1251), .B(n1252), .ZN(n1103) );
XOR2_X1 U958 ( .A(n1253), .B(n1247), .Z(n1252) );
XNOR2_X1 U959 ( .A(n1254), .B(n1085), .ZN(n1247) );
XOR2_X1 U960 ( .A(G140), .B(G125), .Z(n1085) );
NOR2_X1 U961 ( .A1(KEYINPUT2), .A2(n1255), .ZN(n1253) );
XNOR2_X1 U962 ( .A(G137), .B(n1256), .ZN(n1255) );
AND3_X1 U963 ( .A1(G221), .A2(n1069), .A3(G234), .ZN(n1256) );
XOR2_X1 U964 ( .A(n1257), .B(n1258), .Z(n1251) );
NOR2_X1 U965 ( .A1(KEYINPUT6), .A2(n1259), .ZN(n1258) );
XNOR2_X1 U966 ( .A(n1226), .B(G119), .ZN(n1259) );
INV_X1 U967 ( .A(G128), .ZN(n1226) );
XNOR2_X1 U968 ( .A(G110), .B(KEYINPUT20), .ZN(n1257) );
NAND2_X1 U969 ( .A1(n1026), .A2(n1164), .ZN(n1202) );
NAND2_X1 U970 ( .A1(n1011), .A2(n1260), .ZN(n1164) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1194), .A4(n1096), .ZN(n1260) );
INV_X1 U972 ( .A(G898), .ZN(n1096) );
NAND3_X1 U973 ( .A1(n1194), .A2(n1069), .A3(G952), .ZN(n1011) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1194) );
INV_X1 U975 ( .A(n1160), .ZN(n1026) );
NAND2_X1 U976 ( .A1(n1261), .A2(n1028), .ZN(n1160) );
NAND2_X1 U977 ( .A1(n1262), .A2(n1263), .ZN(n1028) );
XOR2_X1 U978 ( .A(KEYINPUT41), .B(G214), .Z(n1262) );
XOR2_X1 U979 ( .A(n1027), .B(KEYINPUT21), .Z(n1261) );
NAND3_X1 U980 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1027) );
INV_X1 U981 ( .A(n1049), .ZN(n1266) );
NOR2_X1 U982 ( .A1(n1267), .A2(n1149), .ZN(n1049) );
NAND2_X1 U983 ( .A1(KEYINPUT12), .A2(n1268), .ZN(n1265) );
NAND2_X1 U984 ( .A1(n1051), .A2(n1269), .ZN(n1264) );
INV_X1 U985 ( .A(KEYINPUT12), .ZN(n1269) );
AND2_X1 U986 ( .A1(n1149), .A2(n1267), .ZN(n1051) );
NAND2_X1 U987 ( .A1(n1270), .A2(n1150), .ZN(n1267) );
XOR2_X1 U988 ( .A(n1146), .B(n1271), .Z(n1270) );
XNOR2_X1 U989 ( .A(KEYINPUT10), .B(n1147), .ZN(n1271) );
INV_X1 U990 ( .A(G125), .ZN(n1147) );
XOR2_X1 U991 ( .A(n1272), .B(n1273), .Z(n1146) );
XOR2_X1 U992 ( .A(n1274), .B(n1275), .Z(n1273) );
NAND2_X1 U993 ( .A1(KEYINPUT39), .A2(n1099), .ZN(n1275) );
XNOR2_X1 U994 ( .A(n1213), .B(G122), .ZN(n1099) );
XOR2_X1 U995 ( .A(n1097), .B(n1276), .Z(n1272) );
NOR2_X1 U996 ( .A1(G953), .A2(n1277), .ZN(n1276) );
XOR2_X1 U997 ( .A(KEYINPUT48), .B(G224), .Z(n1277) );
XOR2_X1 U998 ( .A(n1278), .B(n1279), .Z(n1097) );
XOR2_X1 U999 ( .A(n1280), .B(n1281), .Z(n1279) );
NOR2_X1 U1000 ( .A1(G101), .A2(KEYINPUT34), .ZN(n1280) );
XOR2_X1 U1001 ( .A(n1282), .B(n1283), .Z(n1278) );
XNOR2_X1 U1002 ( .A(n1205), .B(n1284), .ZN(n1283) );
NOR2_X1 U1003 ( .A1(G113), .A2(KEYINPUT17), .ZN(n1284) );
NAND2_X1 U1004 ( .A1(KEYINPUT11), .A2(n1285), .ZN(n1282) );
INV_X1 U1005 ( .A(n1268), .ZN(n1149) );
NAND2_X1 U1006 ( .A1(G210), .A2(n1263), .ZN(n1268) );
NAND2_X1 U1007 ( .A1(n1248), .A2(n1150), .ZN(n1263) );
AND2_X1 U1008 ( .A1(n1043), .A2(n1044), .ZN(n1040) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1250), .ZN(n1044) );
NAND2_X1 U1010 ( .A1(n1286), .A2(n1150), .ZN(n1250) );
XOR2_X1 U1011 ( .A(KEYINPUT47), .B(G234), .Z(n1286) );
XOR2_X1 U1012 ( .A(n1287), .B(n1125), .Z(n1043) );
INV_X1 U1013 ( .A(G469), .ZN(n1125) );
NAND2_X1 U1014 ( .A1(n1288), .A2(n1150), .ZN(n1287) );
XOR2_X1 U1015 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U1016 ( .A(n1141), .B(n1140), .ZN(n1290) );
XNOR2_X1 U1017 ( .A(n1188), .B(n1281), .ZN(n1140) );
XOR2_X1 U1018 ( .A(G104), .B(G107), .Z(n1281) );
INV_X1 U1019 ( .A(n1082), .ZN(n1141) );
XNOR2_X1 U1020 ( .A(n1291), .B(n1292), .ZN(n1082) );
NOR2_X1 U1021 ( .A1(KEYINPUT14), .A2(n1254), .ZN(n1292) );
INV_X1 U1022 ( .A(G146), .ZN(n1254) );
XNOR2_X1 U1023 ( .A(G128), .B(G143), .ZN(n1291) );
XNOR2_X1 U1024 ( .A(n1133), .B(n1293), .ZN(n1289) );
XNOR2_X1 U1025 ( .A(n1137), .B(KEYINPUT22), .ZN(n1293) );
XNOR2_X1 U1026 ( .A(G140), .B(n1213), .ZN(n1137) );
INV_X1 U1027 ( .A(G110), .ZN(n1213) );
XNOR2_X1 U1028 ( .A(n1294), .B(n1295), .ZN(n1133) );
AND2_X1 U1029 ( .A1(n1069), .A2(G227), .ZN(n1295) );
INV_X1 U1030 ( .A(n1034), .ZN(n1192) );
XNOR2_X1 U1031 ( .A(n1296), .B(G472), .ZN(n1034) );
NAND2_X1 U1032 ( .A1(n1297), .A2(n1150), .ZN(n1296) );
INV_X1 U1033 ( .A(G902), .ZN(n1150) );
XOR2_X1 U1034 ( .A(n1298), .B(n1120), .Z(n1297) );
XNOR2_X1 U1035 ( .A(n1299), .B(n1300), .ZN(n1120) );
XNOR2_X1 U1036 ( .A(G113), .B(n1274), .ZN(n1300) );
NAND2_X1 U1037 ( .A1(n1301), .A2(n1302), .ZN(n1274) );
OR2_X1 U1038 ( .A1(n1303), .A2(G128), .ZN(n1302) );
XOR2_X1 U1039 ( .A(n1304), .B(KEYINPUT62), .Z(n1301) );
NAND2_X1 U1040 ( .A1(G128), .A2(n1303), .ZN(n1304) );
XNOR2_X1 U1041 ( .A(G146), .B(n1225), .ZN(n1303) );
INV_X1 U1042 ( .A(G143), .ZN(n1225) );
XOR2_X1 U1043 ( .A(n1294), .B(n1305), .Z(n1299) );
NOR2_X1 U1044 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NOR2_X1 U1045 ( .A1(n1235), .A2(n1205), .ZN(n1307) );
INV_X1 U1046 ( .A(G119), .ZN(n1205) );
NOR2_X1 U1047 ( .A1(G119), .A2(n1308), .ZN(n1306) );
XNOR2_X1 U1048 ( .A(n1309), .B(n1235), .ZN(n1308) );
INV_X1 U1049 ( .A(n1285), .ZN(n1235) );
XOR2_X1 U1050 ( .A(G116), .B(KEYINPUT56), .Z(n1285) );
XNOR2_X1 U1051 ( .A(KEYINPUT61), .B(KEYINPUT4), .ZN(n1309) );
XNOR2_X1 U1052 ( .A(n1310), .B(n1311), .ZN(n1294) );
INV_X1 U1053 ( .A(n1083), .ZN(n1311) );
XOR2_X1 U1054 ( .A(G134), .B(n1312), .Z(n1083) );
XOR2_X1 U1055 ( .A(KEYINPUT52), .B(G137), .Z(n1312) );
NAND2_X1 U1056 ( .A1(KEYINPUT50), .A2(n1081), .ZN(n1310) );
XNOR2_X1 U1057 ( .A(G131), .B(KEYINPUT7), .ZN(n1081) );
NAND2_X1 U1058 ( .A1(KEYINPUT15), .A2(n1117), .ZN(n1298) );
AND2_X1 U1059 ( .A1(n1313), .A2(n1314), .ZN(n1117) );
NAND2_X1 U1060 ( .A1(n1315), .A2(n1188), .ZN(n1314) );
INV_X1 U1061 ( .A(G101), .ZN(n1188) );
NAND3_X1 U1062 ( .A1(n1248), .A2(n1069), .A3(G210), .ZN(n1315) );
NAND4_X1 U1063 ( .A1(n1248), .A2(n1069), .A3(G210), .A4(G101), .ZN(n1313) );
INV_X1 U1064 ( .A(G953), .ZN(n1069) );
INV_X1 U1065 ( .A(G237), .ZN(n1248) );
endmodule


