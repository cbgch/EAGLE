//Key = 1111110000001111011001010010000100001111100011101101110101010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;

XNOR2_X1 U754 ( .A(G107), .B(n1038), .ZN(G9) );
NOR2_X1 U755 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR2_X1 U756 ( .A1(G952), .A2(n1041), .ZN(n1040) );
NOR4_X1 U757 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1039) );
NOR2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR3_X1 U759 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1046) );
NOR2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR3_X1 U762 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1049) );
NOR2_X1 U763 ( .A1(KEYINPUT56), .A2(n1058), .ZN(n1048) );
NOR4_X1 U764 ( .A1(n1059), .A2(n1052), .A3(n1055), .A4(n1060), .ZN(n1044) );
NOR2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U766 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR3_X1 U767 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1063) );
AND2_X1 U768 ( .A1(n1068), .A2(KEYINPUT16), .ZN(n1067) );
NOR3_X1 U769 ( .A1(KEYINPUT16), .A2(n1069), .A3(n1070), .ZN(n1066) );
NOR2_X1 U770 ( .A1(n1071), .A2(n1072), .ZN(n1061) );
NOR2_X1 U771 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1043) );
INV_X1 U773 ( .A(KEYINPUT56), .ZN(n1076) );
NOR2_X1 U774 ( .A1(n1058), .A2(n1047), .ZN(n1075) );
OR3_X1 U775 ( .A1(n1064), .A2(n1072), .A3(n1060), .ZN(n1047) );
OR2_X1 U776 ( .A1(n1077), .A2(n1041), .ZN(n1042) );
NAND2_X1 U777 ( .A1(n1078), .A2(n1079), .ZN(n1041) );
NAND4_X1 U778 ( .A1(n1080), .A2(n1056), .A3(n1081), .A4(n1082), .ZN(n1079) );
NOR4_X1 U779 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
XNOR2_X1 U780 ( .A(n1087), .B(n1088), .ZN(n1086) );
XNOR2_X1 U781 ( .A(KEYINPUT62), .B(KEYINPUT20), .ZN(n1087) );
AND2_X1 U782 ( .A1(n1089), .A2(G469), .ZN(n1085) );
NOR3_X1 U783 ( .A1(n1057), .A2(n1090), .A3(n1091), .ZN(n1081) );
NOR2_X1 U784 ( .A1(KEYINPUT26), .A2(n1053), .ZN(n1091) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1053) );
AND2_X1 U786 ( .A1(n1055), .A2(KEYINPUT26), .ZN(n1090) );
XOR2_X1 U787 ( .A(n1094), .B(n1095), .Z(G72) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1097) );
NAND2_X1 U790 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
NAND2_X1 U791 ( .A1(n1100), .A2(G953), .ZN(n1099) );
XNOR2_X1 U792 ( .A(G900), .B(KEYINPUT47), .ZN(n1100) );
XOR2_X1 U793 ( .A(n1101), .B(n1102), .Z(n1098) );
NOR2_X1 U794 ( .A1(KEYINPUT8), .A2(n1103), .ZN(n1102) );
XOR2_X1 U795 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U797 ( .A1(KEYINPUT9), .A2(n1108), .ZN(n1106) );
XOR2_X1 U798 ( .A(n1109), .B(n1110), .Z(n1104) );
NOR2_X1 U799 ( .A1(n1111), .A2(G953), .ZN(n1101) );
NOR2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(G69) );
XOR2_X1 U802 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U803 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U804 ( .A1(G953), .A2(n1120), .ZN(n1119) );
XOR2_X1 U805 ( .A(KEYINPUT15), .B(n1121), .Z(n1118) );
NAND2_X1 U806 ( .A1(n1096), .A2(n1122), .ZN(n1116) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1122) );
XNOR2_X1 U808 ( .A(n1078), .B(KEYINPUT33), .ZN(n1096) );
NOR2_X1 U809 ( .A1(n1123), .A2(G953), .ZN(n1114) );
NOR2_X1 U810 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XNOR2_X1 U811 ( .A(n1126), .B(n1127), .ZN(n1125) );
NAND2_X1 U812 ( .A1(n1128), .A2(G217), .ZN(n1126) );
NOR2_X1 U813 ( .A1(n1124), .A2(n1129), .ZN(G63) );
XOR2_X1 U814 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U815 ( .A1(n1128), .A2(G478), .ZN(n1130) );
NOR2_X1 U816 ( .A1(n1124), .A2(n1132), .ZN(G60) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U818 ( .A1(n1128), .A2(G475), .ZN(n1133) );
NAND2_X1 U819 ( .A1(n1135), .A2(n1136), .ZN(G6) );
OR2_X1 U820 ( .A1(n1137), .A2(G104), .ZN(n1136) );
XOR2_X1 U821 ( .A(n1138), .B(KEYINPUT11), .Z(n1135) );
NAND2_X1 U822 ( .A1(G104), .A2(n1137), .ZN(n1138) );
NOR3_X1 U823 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(G57) );
AND2_X1 U824 ( .A1(KEYINPUT1), .A2(n1124), .ZN(n1141) );
NOR3_X1 U825 ( .A1(KEYINPUT1), .A2(n1078), .A3(n1142), .ZN(n1140) );
XOR2_X1 U826 ( .A(n1143), .B(n1144), .Z(n1139) );
XNOR2_X1 U827 ( .A(n1145), .B(n1146), .ZN(n1144) );
XOR2_X1 U828 ( .A(n1147), .B(n1148), .Z(n1143) );
XNOR2_X1 U829 ( .A(G101), .B(n1149), .ZN(n1148) );
NAND2_X1 U830 ( .A1(KEYINPUT40), .A2(n1150), .ZN(n1149) );
NAND2_X1 U831 ( .A1(n1128), .A2(G472), .ZN(n1147) );
NOR3_X1 U832 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(G54) );
AND2_X1 U833 ( .A1(n1124), .A2(KEYINPUT21), .ZN(n1153) );
NOR2_X1 U834 ( .A1(n1078), .A2(G952), .ZN(n1124) );
NOR3_X1 U835 ( .A1(KEYINPUT21), .A2(G953), .A3(G952), .ZN(n1152) );
NOR3_X1 U836 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1151) );
AND2_X1 U837 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR3_X1 U838 ( .A1(n1158), .A2(n1159), .A3(n1157), .ZN(n1155) );
NOR2_X1 U839 ( .A1(n1160), .A2(n1161), .ZN(n1154) );
INV_X1 U840 ( .A(n1159), .ZN(n1161) );
XNOR2_X1 U841 ( .A(n1162), .B(n1163), .ZN(n1159) );
XOR2_X1 U842 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U843 ( .A1(n1166), .A2(KEYINPUT12), .ZN(n1164) );
XNOR2_X1 U844 ( .A(n1167), .B(G101), .ZN(n1166) );
XNOR2_X1 U845 ( .A(n1168), .B(n1169), .ZN(n1162) );
XOR2_X1 U846 ( .A(KEYINPUT50), .B(G110), .Z(n1169) );
NOR2_X1 U847 ( .A1(n1157), .A2(n1170), .ZN(n1160) );
XNOR2_X1 U848 ( .A(KEYINPUT53), .B(n1158), .ZN(n1170) );
NAND2_X1 U849 ( .A1(n1128), .A2(G469), .ZN(n1158) );
INV_X1 U850 ( .A(KEYINPUT37), .ZN(n1157) );
NOR2_X1 U851 ( .A1(n1171), .A2(n1172), .ZN(G51) );
XOR2_X1 U852 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U853 ( .A(n1175), .B(KEYINPUT18), .Z(n1174) );
NAND2_X1 U854 ( .A1(n1176), .A2(KEYINPUT49), .ZN(n1175) );
XOR2_X1 U855 ( .A(n1177), .B(n1121), .Z(n1176) );
NAND3_X1 U856 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
NAND2_X1 U857 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U858 ( .A(n1183), .B(n1184), .ZN(n1181) );
NAND3_X1 U859 ( .A1(G125), .A2(n1184), .A3(n1185), .ZN(n1179) );
NAND2_X1 U860 ( .A1(n1186), .A2(n1183), .ZN(n1178) );
NAND2_X1 U861 ( .A1(n1128), .A2(n1187), .ZN(n1173) );
AND2_X1 U862 ( .A1(G902), .A2(n1077), .ZN(n1128) );
NAND3_X1 U863 ( .A1(n1123), .A2(n1188), .A3(n1189), .ZN(n1077) );
XNOR2_X1 U864 ( .A(n1112), .B(KEYINPUT63), .ZN(n1189) );
AND4_X1 U865 ( .A1(n1190), .A2(n1068), .A3(n1054), .A4(n1191), .ZN(n1112) );
XNOR2_X1 U866 ( .A(KEYINPUT4), .B(n1192), .ZN(n1191) );
INV_X1 U867 ( .A(n1113), .ZN(n1188) );
NAND4_X1 U868 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1113) );
NOR4_X1 U869 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196) );
NOR3_X1 U870 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
XNOR2_X1 U871 ( .A(n1054), .B(KEYINPUT32), .ZN(n1202) );
NAND2_X1 U872 ( .A1(n1204), .A2(n1205), .ZN(n1195) );
NAND3_X1 U873 ( .A1(n1206), .A2(n1074), .A3(n1207), .ZN(n1194) );
NAND2_X1 U874 ( .A1(n1208), .A2(n1054), .ZN(n1193) );
XNOR2_X1 U875 ( .A(n1209), .B(KEYINPUT3), .ZN(n1208) );
AND4_X1 U876 ( .A1(n1137), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1123) );
NOR4_X1 U877 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1212) );
AND2_X1 U878 ( .A1(n1038), .A2(n1217), .ZN(n1211) );
NAND3_X1 U879 ( .A1(n1073), .A2(n1218), .A3(n1065), .ZN(n1038) );
NAND3_X1 U880 ( .A1(n1065), .A2(n1218), .A3(n1074), .ZN(n1137) );
NOR2_X1 U881 ( .A1(n1078), .A2(n1219), .ZN(n1171) );
XNOR2_X1 U882 ( .A(KEYINPUT24), .B(n1142), .ZN(n1219) );
INV_X1 U883 ( .A(G952), .ZN(n1142) );
XOR2_X1 U884 ( .A(n1220), .B(G146), .Z(G48) );
NAND2_X1 U885 ( .A1(KEYINPUT13), .A2(n1221), .ZN(n1220) );
NAND4_X1 U886 ( .A1(n1222), .A2(n1223), .A3(n1074), .A4(n1224), .ZN(n1221) );
NOR3_X1 U887 ( .A1(n1225), .A2(n1056), .A3(n1226), .ZN(n1224) );
OR2_X1 U888 ( .A1(n1227), .A2(n1206), .ZN(n1223) );
NAND2_X1 U889 ( .A1(n1228), .A2(n1227), .ZN(n1222) );
INV_X1 U890 ( .A(KEYINPUT17), .ZN(n1227) );
NAND2_X1 U891 ( .A1(n1229), .A2(n1065), .ZN(n1228) );
XOR2_X1 U892 ( .A(G143), .B(n1199), .Z(G45) );
AND3_X1 U893 ( .A1(n1206), .A2(n1230), .A3(n1231), .ZN(n1199) );
NOR3_X1 U894 ( .A1(n1225), .A2(n1080), .A3(n1088), .ZN(n1231) );
XNOR2_X1 U895 ( .A(n1232), .B(n1198), .ZN(G42) );
AND3_X1 U896 ( .A1(n1206), .A2(n1205), .A3(n1190), .ZN(n1198) );
XNOR2_X1 U897 ( .A(n1233), .B(n1197), .ZN(G39) );
NOR3_X1 U898 ( .A1(n1055), .A2(n1064), .A3(n1201), .ZN(n1197) );
XNOR2_X1 U899 ( .A(G134), .B(n1234), .ZN(G36) );
NAND3_X1 U900 ( .A1(n1205), .A2(n1235), .A3(KEYINPUT39), .ZN(n1234) );
XOR2_X1 U901 ( .A(KEYINPUT6), .B(n1204), .Z(n1235) );
AND3_X1 U902 ( .A1(n1230), .A2(n1073), .A3(n1206), .ZN(n1204) );
XOR2_X1 U903 ( .A(n1236), .B(n1237), .Z(G33) );
NAND2_X1 U904 ( .A1(KEYINPUT48), .A2(G131), .ZN(n1237) );
NAND4_X1 U905 ( .A1(n1238), .A2(n1207), .A3(n1074), .A4(n1192), .ZN(n1236) );
INV_X1 U906 ( .A(n1058), .ZN(n1207) );
NAND2_X1 U907 ( .A1(n1230), .A2(n1205), .ZN(n1058) );
INV_X1 U908 ( .A(n1055), .ZN(n1205) );
NAND2_X1 U909 ( .A1(n1239), .A2(n1093), .ZN(n1055) );
INV_X1 U910 ( .A(n1092), .ZN(n1239) );
XNOR2_X1 U911 ( .A(n1065), .B(KEYINPUT38), .ZN(n1238) );
XNOR2_X1 U912 ( .A(G128), .B(n1240), .ZN(G30) );
NAND2_X1 U913 ( .A1(n1209), .A2(n1054), .ZN(n1240) );
NOR2_X1 U914 ( .A1(n1201), .A2(n1241), .ZN(n1209) );
NAND3_X1 U915 ( .A1(n1057), .A2(n1242), .A3(n1206), .ZN(n1201) );
NOR2_X1 U916 ( .A1(n1243), .A2(n1229), .ZN(n1206) );
NAND2_X1 U917 ( .A1(n1244), .A2(n1245), .ZN(G3) );
OR2_X1 U918 ( .A1(n1246), .A2(G101), .ZN(n1245) );
NAND2_X1 U919 ( .A1(n1247), .A2(G101), .ZN(n1244) );
NAND2_X1 U920 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U921 ( .A1(n1216), .A2(n1250), .ZN(n1249) );
INV_X1 U922 ( .A(KEYINPUT36), .ZN(n1250) );
NAND2_X1 U923 ( .A1(KEYINPUT36), .A2(n1246), .ZN(n1248) );
NAND2_X1 U924 ( .A1(KEYINPUT52), .A2(n1216), .ZN(n1246) );
AND2_X1 U925 ( .A1(n1230), .A2(n1251), .ZN(n1216) );
XNOR2_X1 U926 ( .A(G125), .B(n1252), .ZN(G27) );
NAND3_X1 U927 ( .A1(KEYINPUT51), .A2(n1190), .A3(n1253), .ZN(n1252) );
NOR3_X1 U928 ( .A1(n1072), .A2(n1229), .A3(n1225), .ZN(n1253) );
INV_X1 U929 ( .A(n1192), .ZN(n1229) );
NAND2_X1 U930 ( .A1(n1060), .A2(n1254), .ZN(n1192) );
NAND4_X1 U931 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1256), .ZN(n1254) );
INV_X1 U932 ( .A(G900), .ZN(n1256) );
NOR3_X1 U933 ( .A1(n1057), .A2(n1056), .A3(n1203), .ZN(n1190) );
INV_X1 U934 ( .A(n1074), .ZN(n1203) );
INV_X1 U935 ( .A(n1242), .ZN(n1056) );
XNOR2_X1 U936 ( .A(G122), .B(n1210), .ZN(G24) );
NAND4_X1 U937 ( .A1(n1068), .A2(n1218), .A3(n1257), .A4(n1258), .ZN(n1210) );
NOR2_X1 U938 ( .A1(n1259), .A2(n1052), .ZN(n1218) );
NAND2_X1 U939 ( .A1(n1226), .A2(n1260), .ZN(n1052) );
XNOR2_X1 U940 ( .A(KEYINPUT27), .B(n1242), .ZN(n1260) );
XNOR2_X1 U941 ( .A(n1215), .B(n1261), .ZN(G21) );
NOR2_X1 U942 ( .A1(G119), .A2(KEYINPUT42), .ZN(n1261) );
AND4_X1 U943 ( .A1(n1057), .A2(n1242), .A3(n1262), .A4(n1263), .ZN(n1215) );
NOR2_X1 U944 ( .A1(n1072), .A2(n1064), .ZN(n1263) );
INV_X1 U945 ( .A(n1068), .ZN(n1072) );
XNOR2_X1 U946 ( .A(G116), .B(n1264), .ZN(G18) );
NAND2_X1 U947 ( .A1(KEYINPUT55), .A2(n1214), .ZN(n1264) );
AND4_X1 U948 ( .A1(n1230), .A2(n1068), .A3(n1073), .A4(n1262), .ZN(n1214) );
INV_X1 U949 ( .A(n1241), .ZN(n1073) );
NAND2_X1 U950 ( .A1(n1080), .A2(n1257), .ZN(n1241) );
XNOR2_X1 U951 ( .A(G113), .B(n1217), .ZN(G15) );
NAND4_X1 U952 ( .A1(n1074), .A2(n1230), .A3(n1068), .A4(n1262), .ZN(n1217) );
INV_X1 U953 ( .A(n1259), .ZN(n1262) );
NOR2_X1 U954 ( .A1(n1069), .A2(n1084), .ZN(n1068) );
INV_X1 U955 ( .A(n1265), .ZN(n1069) );
NOR2_X1 U956 ( .A1(n1242), .A2(n1226), .ZN(n1230) );
NOR2_X1 U957 ( .A1(n1257), .A2(n1080), .ZN(n1074) );
XOR2_X1 U958 ( .A(G110), .B(n1213), .Z(G12) );
AND3_X1 U959 ( .A1(n1226), .A2(n1242), .A3(n1251), .ZN(n1213) );
NOR3_X1 U960 ( .A1(n1243), .A2(n1259), .A3(n1064), .ZN(n1251) );
NAND2_X1 U961 ( .A1(n1088), .A2(n1080), .ZN(n1064) );
INV_X1 U962 ( .A(n1258), .ZN(n1080) );
XNOR2_X1 U963 ( .A(n1266), .B(G475), .ZN(n1258) );
NAND2_X1 U964 ( .A1(n1134), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U965 ( .A(n1268), .B(n1269), .ZN(n1134) );
XOR2_X1 U966 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U967 ( .A(n1272), .B(n1273), .ZN(n1271) );
XNOR2_X1 U968 ( .A(n1274), .B(n1275), .ZN(n1270) );
NOR2_X1 U969 ( .A1(KEYINPUT60), .A2(n1232), .ZN(n1275) );
NOR2_X1 U970 ( .A1(G104), .A2(KEYINPUT54), .ZN(n1274) );
XOR2_X1 U971 ( .A(n1276), .B(n1277), .Z(n1268) );
XNOR2_X1 U972 ( .A(G143), .B(n1182), .ZN(n1277) );
XOR2_X1 U973 ( .A(n1278), .B(n1279), .Z(n1276) );
AND3_X1 U974 ( .A1(G214), .A2(n1078), .A3(n1280), .ZN(n1279) );
NAND2_X1 U975 ( .A1(KEYINPUT14), .A2(n1281), .ZN(n1278) );
INV_X1 U976 ( .A(n1257), .ZN(n1088) );
XNOR2_X1 U977 ( .A(n1282), .B(G478), .ZN(n1257) );
NAND2_X1 U978 ( .A1(n1131), .A2(n1267), .ZN(n1282) );
XOR2_X1 U979 ( .A(n1283), .B(n1284), .Z(n1131) );
NOR2_X1 U980 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U981 ( .A1(n1287), .A2(KEYINPUT0), .ZN(n1283) );
XOR2_X1 U982 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U983 ( .A(n1290), .B(n1291), .ZN(n1289) );
NOR2_X1 U984 ( .A1(KEYINPUT22), .A2(n1292), .ZN(n1291) );
XOR2_X1 U985 ( .A(n1293), .B(n1108), .Z(n1292) );
NAND2_X1 U986 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NAND2_X1 U987 ( .A1(KEYINPUT10), .A2(n1296), .ZN(n1295) );
INV_X1 U988 ( .A(n1297), .ZN(n1296) );
NAND2_X1 U989 ( .A1(KEYINPUT44), .A2(n1297), .ZN(n1294) );
XOR2_X1 U990 ( .A(G128), .B(G143), .Z(n1297) );
NAND2_X1 U991 ( .A1(KEYINPUT57), .A2(n1298), .ZN(n1290) );
XNOR2_X1 U992 ( .A(G116), .B(G107), .ZN(n1288) );
NAND2_X1 U993 ( .A1(n1054), .A2(n1299), .ZN(n1259) );
NAND2_X1 U994 ( .A1(n1060), .A2(n1300), .ZN(n1299) );
NAND4_X1 U995 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1120), .ZN(n1300) );
INV_X1 U996 ( .A(G898), .ZN(n1120) );
NAND3_X1 U997 ( .A1(n1255), .A2(n1078), .A3(G952), .ZN(n1060) );
NAND2_X1 U998 ( .A1(G237), .A2(G234), .ZN(n1255) );
INV_X1 U999 ( .A(n1225), .ZN(n1054) );
NAND2_X1 U1000 ( .A1(n1092), .A2(n1093), .ZN(n1225) );
NAND2_X1 U1001 ( .A1(G214), .A2(n1301), .ZN(n1093) );
XNOR2_X1 U1002 ( .A(n1302), .B(n1187), .ZN(n1092) );
AND2_X1 U1003 ( .A1(G210), .A2(n1301), .ZN(n1187) );
NAND2_X1 U1004 ( .A1(n1280), .A2(n1267), .ZN(n1301) );
NAND2_X1 U1005 ( .A1(n1303), .A2(n1267), .ZN(n1302) );
XOR2_X1 U1006 ( .A(n1304), .B(n1121), .Z(n1303) );
XNOR2_X1 U1007 ( .A(n1305), .B(n1306), .ZN(n1121) );
XOR2_X1 U1008 ( .A(n1272), .B(n1307), .Z(n1306) );
XNOR2_X1 U1009 ( .A(G113), .B(n1298), .ZN(n1272) );
INV_X1 U1010 ( .A(G122), .ZN(n1298) );
XOR2_X1 U1011 ( .A(n1308), .B(n1309), .Z(n1305) );
XNOR2_X1 U1012 ( .A(G104), .B(G107), .ZN(n1308) );
NAND2_X1 U1013 ( .A1(n1310), .A2(n1311), .ZN(n1304) );
NAND3_X1 U1014 ( .A1(n1312), .A2(n1313), .A3(n1185), .ZN(n1311) );
INV_X1 U1015 ( .A(n1183), .ZN(n1185) );
XOR2_X1 U1016 ( .A(n1314), .B(KEYINPUT29), .Z(n1310) );
NAND2_X1 U1017 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1018 ( .A1(n1312), .A2(n1313), .ZN(n1316) );
INV_X1 U1019 ( .A(n1186), .ZN(n1313) );
NOR2_X1 U1020 ( .A1(n1184), .A2(n1182), .ZN(n1186) );
XOR2_X1 U1021 ( .A(n1317), .B(KEYINPUT28), .Z(n1312) );
NAND2_X1 U1022 ( .A1(n1184), .A2(n1182), .ZN(n1317) );
INV_X1 U1023 ( .A(G125), .ZN(n1182) );
XNOR2_X1 U1024 ( .A(n1318), .B(n1183), .ZN(n1315) );
NAND2_X1 U1025 ( .A1(G224), .A2(n1078), .ZN(n1183) );
XNOR2_X1 U1026 ( .A(KEYINPUT34), .B(KEYINPUT25), .ZN(n1318) );
INV_X1 U1027 ( .A(n1065), .ZN(n1243) );
NOR2_X1 U1028 ( .A1(n1084), .A2(n1265), .ZN(n1065) );
NOR2_X1 U1029 ( .A1(n1319), .A2(n1083), .ZN(n1265) );
NOR2_X1 U1030 ( .A1(n1089), .A2(G469), .ZN(n1083) );
AND2_X1 U1031 ( .A1(n1320), .A2(n1089), .ZN(n1319) );
NAND2_X1 U1032 ( .A1(n1321), .A2(n1267), .ZN(n1089) );
XOR2_X1 U1033 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1034 ( .A(n1324), .B(n1307), .ZN(n1323) );
XOR2_X1 U1035 ( .A(G110), .B(G101), .Z(n1307) );
NAND2_X1 U1036 ( .A1(KEYINPUT31), .A2(n1168), .ZN(n1324) );
AND2_X1 U1037 ( .A1(G227), .A2(n1078), .ZN(n1168) );
XNOR2_X1 U1038 ( .A(n1165), .B(n1325), .ZN(n1322) );
INV_X1 U1039 ( .A(n1167), .ZN(n1325) );
XNOR2_X1 U1040 ( .A(n1326), .B(n1110), .ZN(n1167) );
XNOR2_X1 U1041 ( .A(n1327), .B(n1328), .ZN(n1110) );
NOR2_X1 U1042 ( .A1(KEYINPUT7), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1043 ( .A(G107), .B(n1330), .ZN(n1326) );
NOR2_X1 U1044 ( .A1(KEYINPUT41), .A2(n1331), .ZN(n1330) );
INV_X1 U1045 ( .A(G104), .ZN(n1331) );
XNOR2_X1 U1046 ( .A(n1332), .B(n1232), .ZN(n1165) );
XNOR2_X1 U1047 ( .A(G469), .B(KEYINPUT5), .ZN(n1320) );
INV_X1 U1048 ( .A(n1070), .ZN(n1084) );
NAND2_X1 U1049 ( .A1(G221), .A2(n1333), .ZN(n1070) );
NAND2_X1 U1050 ( .A1(G234), .A2(n1267), .ZN(n1333) );
NAND3_X1 U1051 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1242) );
NAND2_X1 U1052 ( .A1(n1337), .A2(n1127), .ZN(n1336) );
OR3_X1 U1053 ( .A1(n1127), .A2(n1337), .A3(G902), .ZN(n1335) );
NOR2_X1 U1054 ( .A1(n1286), .A2(G234), .ZN(n1337) );
INV_X1 U1055 ( .A(G217), .ZN(n1286) );
XOR2_X1 U1056 ( .A(n1338), .B(n1339), .Z(n1127) );
NOR2_X1 U1057 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1058 ( .A(KEYINPUT35), .B(n1342), .Z(n1341) );
NOR3_X1 U1059 ( .A1(n1285), .A2(n1233), .A3(n1343), .ZN(n1342) );
INV_X1 U1060 ( .A(G137), .ZN(n1233) );
NOR2_X1 U1061 ( .A1(n1344), .A2(G137), .ZN(n1340) );
NOR2_X1 U1062 ( .A1(n1343), .A2(n1285), .ZN(n1344) );
NAND2_X1 U1063 ( .A1(G234), .A2(n1078), .ZN(n1285) );
INV_X1 U1064 ( .A(G221), .ZN(n1343) );
NAND4_X1 U1065 ( .A1(n1345), .A2(n1346), .A3(n1347), .A4(n1348), .ZN(n1338) );
NAND3_X1 U1066 ( .A1(KEYINPUT2), .A2(n1349), .A3(n1350), .ZN(n1348) );
XNOR2_X1 U1067 ( .A(n1351), .B(KEYINPUT58), .ZN(n1349) );
OR2_X1 U1068 ( .A1(n1350), .A2(KEYINPUT2), .ZN(n1347) );
NAND3_X1 U1069 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1346) );
INV_X1 U1070 ( .A(KEYINPUT59), .ZN(n1354) );
NAND2_X1 U1071 ( .A1(n1350), .A2(KEYINPUT58), .ZN(n1353) );
INV_X1 U1072 ( .A(n1351), .ZN(n1352) );
NAND3_X1 U1073 ( .A1(n1351), .A2(n1355), .A3(KEYINPUT59), .ZN(n1345) );
NAND2_X1 U1074 ( .A1(n1350), .A2(n1356), .ZN(n1355) );
INV_X1 U1075 ( .A(KEYINPUT58), .ZN(n1356) );
XNOR2_X1 U1076 ( .A(n1357), .B(n1281), .ZN(n1350) );
XNOR2_X1 U1077 ( .A(G146), .B(KEYINPUT30), .ZN(n1281) );
NAND2_X1 U1078 ( .A1(KEYINPUT46), .A2(n1107), .ZN(n1357) );
XNOR2_X1 U1079 ( .A(n1232), .B(G125), .ZN(n1107) );
INV_X1 U1080 ( .A(G140), .ZN(n1232) );
XOR2_X1 U1081 ( .A(G110), .B(n1358), .Z(n1351) );
XNOR2_X1 U1082 ( .A(n1329), .B(G119), .ZN(n1358) );
INV_X1 U1083 ( .A(G128), .ZN(n1329) );
NAND2_X1 U1084 ( .A1(G902), .A2(G217), .ZN(n1334) );
INV_X1 U1085 ( .A(n1057), .ZN(n1226) );
XNOR2_X1 U1086 ( .A(n1359), .B(G472), .ZN(n1057) );
NAND2_X1 U1087 ( .A1(n1360), .A2(n1267), .ZN(n1359) );
INV_X1 U1088 ( .A(G902), .ZN(n1267) );
XOR2_X1 U1089 ( .A(n1361), .B(n1362), .Z(n1360) );
XNOR2_X1 U1090 ( .A(n1150), .B(n1146), .ZN(n1362) );
XOR2_X1 U1091 ( .A(G113), .B(n1309), .Z(n1146) );
XNOR2_X1 U1092 ( .A(n1363), .B(G119), .ZN(n1309) );
INV_X1 U1093 ( .A(G116), .ZN(n1363) );
NAND3_X1 U1094 ( .A1(n1280), .A2(n1078), .A3(G210), .ZN(n1150) );
INV_X1 U1095 ( .A(G953), .ZN(n1078) );
INV_X1 U1096 ( .A(G237), .ZN(n1280) );
XOR2_X1 U1097 ( .A(n1364), .B(n1365), .Z(n1361) );
XNOR2_X1 U1098 ( .A(KEYINPUT45), .B(n1366), .ZN(n1365) );
NOR2_X1 U1099 ( .A1(KEYINPUT19), .A2(n1145), .ZN(n1366) );
XOR2_X1 U1100 ( .A(n1332), .B(n1184), .Z(n1145) );
XNOR2_X1 U1101 ( .A(G128), .B(n1327), .ZN(n1184) );
XNOR2_X1 U1102 ( .A(G146), .B(G143), .ZN(n1327) );
XNOR2_X1 U1103 ( .A(n1109), .B(n1108), .ZN(n1332) );
XNOR2_X1 U1104 ( .A(G134), .B(KEYINPUT23), .ZN(n1108) );
XNOR2_X1 U1105 ( .A(G137), .B(n1273), .ZN(n1109) );
XOR2_X1 U1106 ( .A(G131), .B(KEYINPUT43), .Z(n1273) );
NAND2_X1 U1107 ( .A1(KEYINPUT61), .A2(G101), .ZN(n1364) );
endmodule


