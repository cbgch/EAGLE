//Key = 0100111100000110000010011111000100111000101011001010000100110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;

XOR2_X1 U710 ( .A(G107), .B(n973), .Z(G9) );
NOR2_X1 U711 ( .A1(n974), .A2(n975), .ZN(G75) );
NOR4_X1 U712 ( .A1(G953), .A2(n976), .A3(n977), .A4(n978), .ZN(n975) );
NOR2_X1 U713 ( .A1(n979), .A2(n980), .ZN(n977) );
NOR2_X1 U714 ( .A1(n981), .A2(n982), .ZN(n979) );
NOR3_X1 U715 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n982) );
NOR2_X1 U716 ( .A1(n986), .A2(n987), .ZN(n984) );
AND2_X1 U717 ( .A1(n988), .A2(n989), .ZN(n987) );
NOR3_X1 U718 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n986) );
NOR3_X1 U719 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NOR2_X1 U720 ( .A1(n989), .A2(n996), .ZN(n991) );
NOR3_X1 U721 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n981) );
INV_X1 U722 ( .A(n989), .ZN(n999) );
NOR2_X1 U723 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR2_X1 U724 ( .A1(n1002), .A2(n985), .ZN(n1001) );
INV_X1 U725 ( .A(n1003), .ZN(n985) );
NOR2_X1 U726 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NOR2_X1 U727 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U728 ( .A1(n1008), .A2(n983), .ZN(n1000) );
NOR2_X1 U729 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
AND2_X1 U730 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR3_X1 U731 ( .A1(n976), .A2(G953), .A3(G952), .ZN(n974) );
AND4_X1 U732 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n976) );
NOR4_X1 U733 ( .A1(n1017), .A2(n993), .A3(n1018), .A4(n1019), .ZN(n1016) );
NOR2_X1 U734 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
INV_X1 U735 ( .A(G478), .ZN(n1021) );
NOR2_X1 U736 ( .A1(G902), .A2(n1022), .ZN(n1020) );
NOR2_X1 U737 ( .A1(n983), .A2(n1023), .ZN(n1015) );
XOR2_X1 U738 ( .A(n1024), .B(n1025), .Z(n1014) );
NAND2_X1 U739 ( .A1(KEYINPUT36), .A2(n1026), .ZN(n1024) );
XOR2_X1 U740 ( .A(n1027), .B(n1028), .Z(n1013) );
XOR2_X1 U741 ( .A(n1029), .B(n1030), .Z(G72) );
XOR2_X1 U742 ( .A(n1031), .B(n1032), .Z(n1030) );
NAND2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U744 ( .A1(G953), .A2(n1035), .ZN(n1034) );
XOR2_X1 U745 ( .A(n1036), .B(n1037), .Z(n1033) );
XOR2_X1 U746 ( .A(n1038), .B(n1039), .Z(n1037) );
NAND2_X1 U747 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND3_X1 U748 ( .A1(G131), .A2(n1042), .A3(n1043), .ZN(n1041) );
OR2_X1 U749 ( .A1(n1044), .A2(n1043), .ZN(n1040) );
INV_X1 U750 ( .A(KEYINPUT7), .ZN(n1043) );
XOR2_X1 U751 ( .A(n1045), .B(KEYINPUT43), .Z(n1036) );
NAND2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1031) );
NAND2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U754 ( .A(KEYINPUT8), .B(n1050), .Z(n1049) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U756 ( .A(KEYINPUT41), .B(n1053), .ZN(n1052) );
INV_X1 U757 ( .A(n1054), .ZN(n1048) );
XOR2_X1 U758 ( .A(KEYINPUT55), .B(G953), .Z(n1046) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1029) );
AND2_X1 U760 ( .A1(G227), .A2(G900), .ZN(n1055) );
XOR2_X1 U761 ( .A(n1057), .B(n1058), .Z(G69) );
NOR2_X1 U762 ( .A1(n1059), .A2(n1056), .ZN(n1058) );
AND2_X1 U763 ( .A1(G224), .A2(G898), .ZN(n1059) );
NOR3_X1 U764 ( .A1(KEYINPUT61), .A2(n1060), .A3(n1061), .ZN(n1057) );
NOR2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
INV_X1 U766 ( .A(n1064), .ZN(n1063) );
NOR2_X1 U767 ( .A1(n1065), .A2(n1064), .ZN(n1060) );
XOR2_X1 U768 ( .A(n1066), .B(n1067), .Z(n1064) );
XOR2_X1 U769 ( .A(KEYINPUT51), .B(n1068), .Z(n1067) );
XOR2_X1 U770 ( .A(n1069), .B(n1070), .Z(n1066) );
NOR2_X1 U771 ( .A1(n1062), .A2(n1071), .ZN(n1065) );
NOR2_X1 U772 ( .A1(n1056), .A2(n1072), .ZN(n1071) );
XOR2_X1 U773 ( .A(KEYINPUT3), .B(G898), .Z(n1072) );
AND2_X1 U774 ( .A1(n1056), .A2(n1073), .ZN(n1062) );
NOR2_X1 U775 ( .A1(n1074), .A2(n1075), .ZN(G66) );
XNOR2_X1 U776 ( .A(n1076), .B(n1077), .ZN(n1075) );
XNOR2_X1 U777 ( .A(KEYINPUT50), .B(n1078), .ZN(n1077) );
NOR3_X1 U778 ( .A1(n1079), .A2(KEYINPUT49), .A3(n1080), .ZN(n1078) );
NOR2_X1 U779 ( .A1(n1074), .A2(n1081), .ZN(G63) );
XOR2_X1 U780 ( .A(n1082), .B(n1083), .Z(n1081) );
NAND3_X1 U781 ( .A1(n1084), .A2(n1085), .A3(G478), .ZN(n1082) );
NAND2_X1 U782 ( .A1(KEYINPUT48), .A2(n1079), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
INV_X1 U784 ( .A(KEYINPUT48), .ZN(n1087) );
NAND2_X1 U785 ( .A1(n1088), .A2(G902), .ZN(n1086) );
NOR2_X1 U786 ( .A1(n1074), .A2(n1089), .ZN(G60) );
XNOR2_X1 U787 ( .A(n1090), .B(n1091), .ZN(n1089) );
AND2_X1 U788 ( .A1(G475), .A2(n1092), .ZN(n1091) );
XNOR2_X1 U789 ( .A(G104), .B(n1093), .ZN(G6) );
NAND2_X1 U790 ( .A1(KEYINPUT58), .A2(n1094), .ZN(n1093) );
NOR2_X1 U791 ( .A1(n1074), .A2(n1095), .ZN(G57) );
XOR2_X1 U792 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U793 ( .A(n1045), .B(n1098), .Z(n1096) );
AND2_X1 U794 ( .A1(G472), .A2(n1092), .ZN(n1098) );
NOR2_X1 U795 ( .A1(n1074), .A2(n1099), .ZN(G54) );
XOR2_X1 U796 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U797 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U798 ( .A(n1104), .B(n1105), .Z(n1103) );
XNOR2_X1 U799 ( .A(n1106), .B(n1107), .ZN(n1102) );
NAND2_X1 U800 ( .A1(KEYINPUT42), .A2(n1044), .ZN(n1107) );
NAND2_X1 U801 ( .A1(KEYINPUT26), .A2(n1108), .ZN(n1106) );
XOR2_X1 U802 ( .A(n1109), .B(n1110), .Z(n1100) );
XOR2_X1 U803 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR3_X1 U804 ( .A1(n1079), .A2(KEYINPUT56), .A3(n1028), .ZN(n1112) );
XOR2_X1 U805 ( .A(KEYINPUT31), .B(G101), .Z(n1109) );
NOR2_X1 U806 ( .A1(n1074), .A2(n1113), .ZN(G51) );
XOR2_X1 U807 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U808 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND3_X1 U809 ( .A1(n1092), .A2(G210), .A3(KEYINPUT44), .ZN(n1116) );
INV_X1 U810 ( .A(n1079), .ZN(n1092) );
NAND2_X1 U811 ( .A1(G902), .A2(n978), .ZN(n1079) );
INV_X1 U812 ( .A(n1088), .ZN(n978) );
NOR4_X1 U813 ( .A1(n1118), .A2(n1073), .A3(n1051), .A4(n1054), .ZN(n1088) );
NAND4_X1 U814 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1054) );
NAND3_X1 U815 ( .A1(n1123), .A2(n989), .A3(n1124), .ZN(n1119) );
XOR2_X1 U816 ( .A(n983), .B(KEYINPUT27), .Z(n1124) );
INV_X1 U817 ( .A(n1125), .ZN(n983) );
NAND3_X1 U818 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1051) );
NAND3_X1 U819 ( .A1(n1125), .A2(n995), .A3(n1129), .ZN(n1128) );
NAND2_X1 U820 ( .A1(n1130), .A2(n1131), .ZN(n1073) );
NOR4_X1 U821 ( .A1(n1132), .A2(n973), .A3(n1133), .A4(n1134), .ZN(n1131) );
AND3_X1 U822 ( .A1(n995), .A2(n1135), .A3(n1003), .ZN(n973) );
NOR4_X1 U823 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1094), .ZN(n1130) );
AND3_X1 U824 ( .A1(n1003), .A2(n1135), .A3(n994), .ZN(n1094) );
INV_X1 U825 ( .A(n1139), .ZN(n1138) );
NOR2_X1 U826 ( .A1(n1140), .A2(n1141), .ZN(n1136) );
XNOR2_X1 U827 ( .A(n1053), .B(KEYINPUT60), .ZN(n1118) );
XOR2_X1 U828 ( .A(n1142), .B(n1143), .Z(n1114) );
NOR2_X1 U829 ( .A1(KEYINPUT33), .A2(n1144), .ZN(n1143) );
XOR2_X1 U830 ( .A(n1145), .B(KEYINPUT6), .Z(n1144) );
NOR2_X1 U831 ( .A1(n1056), .A2(G952), .ZN(n1074) );
NAND2_X1 U832 ( .A1(n1146), .A2(n1147), .ZN(G48) );
NAND2_X1 U833 ( .A1(G146), .A2(n1121), .ZN(n1147) );
XOR2_X1 U834 ( .A(KEYINPUT40), .B(n1148), .Z(n1146) );
NOR2_X1 U835 ( .A1(G146), .A2(n1121), .ZN(n1148) );
NAND3_X1 U836 ( .A1(n994), .A2(n1005), .A3(n1123), .ZN(n1121) );
NAND2_X1 U837 ( .A1(n1149), .A2(n1150), .ZN(G45) );
NAND2_X1 U838 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U839 ( .A(n1153), .B(KEYINPUT47), .Z(n1149) );
OR2_X1 U840 ( .A1(n1151), .A2(n1152), .ZN(n1153) );
NAND2_X1 U841 ( .A1(n1154), .A2(n1155), .ZN(n1151) );
OR2_X1 U842 ( .A1(n1120), .A2(KEYINPUT32), .ZN(n1155) );
NAND4_X1 U843 ( .A1(n1129), .A2(n1005), .A3(n1023), .A4(n1156), .ZN(n1120) );
NAND4_X1 U844 ( .A1(n1157), .A2(n1156), .A3(n1158), .A4(KEYINPUT32), .ZN(n1154) );
NOR2_X1 U845 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U846 ( .A(G140), .B(n1122), .ZN(G42) );
NAND3_X1 U847 ( .A1(n1125), .A2(n990), .A3(n1161), .ZN(n1122) );
NAND2_X1 U848 ( .A1(n1162), .A2(n1163), .ZN(G39) );
NAND3_X1 U849 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1163) );
INV_X1 U850 ( .A(KEYINPUT9), .ZN(n1165) );
NAND2_X1 U851 ( .A1(n1167), .A2(n1168), .ZN(n1162) );
NAND2_X1 U852 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND2_X1 U853 ( .A1(n1164), .A2(n1171), .ZN(n1170) );
OR2_X1 U854 ( .A1(KEYINPUT29), .A2(KEYINPUT9), .ZN(n1171) );
OR2_X1 U855 ( .A1(n1164), .A2(KEYINPUT29), .ZN(n1169) );
XOR2_X1 U856 ( .A(G137), .B(KEYINPUT2), .Z(n1164) );
INV_X1 U857 ( .A(n1166), .ZN(n1167) );
NAND3_X1 U858 ( .A1(n989), .A2(n1125), .A3(n1123), .ZN(n1166) );
XNOR2_X1 U859 ( .A(G134), .B(n1172), .ZN(G36) );
NAND2_X1 U860 ( .A1(n1125), .A2(n1173), .ZN(n1172) );
XOR2_X1 U861 ( .A(KEYINPUT11), .B(n1174), .Z(n1173) );
NOR2_X1 U862 ( .A1(n1175), .A2(n1160), .ZN(n1174) );
XNOR2_X1 U863 ( .A(n1126), .B(n1176), .ZN(G33) );
XOR2_X1 U864 ( .A(KEYINPUT39), .B(G131), .Z(n1176) );
NAND3_X1 U865 ( .A1(n994), .A2(n1125), .A3(n1129), .ZN(n1126) );
INV_X1 U866 ( .A(n1160), .ZN(n1129) );
NAND3_X1 U867 ( .A1(n988), .A2(n1177), .A3(n1010), .ZN(n1160) );
NOR2_X1 U868 ( .A1(n1006), .A2(n1178), .ZN(n1125) );
XNOR2_X1 U869 ( .A(G128), .B(n1053), .ZN(G30) );
NAND3_X1 U870 ( .A1(n995), .A2(n1005), .A3(n1123), .ZN(n1053) );
AND4_X1 U871 ( .A1(n1012), .A2(n1179), .A3(n988), .A4(n1177), .ZN(n1123) );
XOR2_X1 U872 ( .A(n1132), .B(n1180), .Z(G3) );
NOR2_X1 U873 ( .A1(KEYINPUT15), .A2(n1181), .ZN(n1180) );
AND3_X1 U874 ( .A1(n1010), .A2(n1135), .A3(n989), .ZN(n1132) );
NOR2_X1 U875 ( .A1(n1140), .A2(n1182), .ZN(n1135) );
XOR2_X1 U876 ( .A(G125), .B(n1183), .Z(G27) );
NOR2_X1 U877 ( .A1(KEYINPUT62), .A2(n1127), .ZN(n1183) );
NAND3_X1 U878 ( .A1(n1184), .A2(n1005), .A3(n1161), .ZN(n1127) );
AND3_X1 U879 ( .A1(n1012), .A2(n994), .A3(n1185), .ZN(n1161) );
AND3_X1 U880 ( .A1(n1011), .A2(n1177), .A3(n996), .ZN(n1185) );
NAND2_X1 U881 ( .A1(n1186), .A2(n980), .ZN(n1177) );
NAND2_X1 U882 ( .A1(n1187), .A2(n1035), .ZN(n1186) );
INV_X1 U883 ( .A(G900), .ZN(n1035) );
INV_X1 U884 ( .A(n1157), .ZN(n1005) );
XOR2_X1 U885 ( .A(n1188), .B(n1139), .Z(G24) );
NAND4_X1 U886 ( .A1(n1189), .A2(n1003), .A3(n1023), .A4(n1156), .ZN(n1139) );
NOR2_X1 U887 ( .A1(n1019), .A2(n1179), .ZN(n1003) );
XOR2_X1 U888 ( .A(G119), .B(n1137), .Z(G21) );
AND4_X1 U889 ( .A1(n1012), .A2(n1189), .A3(n1179), .A4(n989), .ZN(n1137) );
XOR2_X1 U890 ( .A(n1190), .B(G116), .Z(G18) );
NAND2_X1 U891 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND2_X1 U892 ( .A1(n1133), .A2(n1193), .ZN(n1192) );
INV_X1 U893 ( .A(KEYINPUT17), .ZN(n1193) );
AND3_X1 U894 ( .A1(n1010), .A2(n995), .A3(n1189), .ZN(n1133) );
NAND4_X1 U895 ( .A1(n995), .A2(n1194), .A3(n1189), .A4(KEYINPUT17), .ZN(n1191) );
NOR3_X1 U896 ( .A1(n1157), .A2(n1195), .A3(n997), .ZN(n1189) );
XOR2_X1 U897 ( .A(n1140), .B(KEYINPUT22), .Z(n1157) );
INV_X1 U898 ( .A(n1175), .ZN(n995) );
NAND2_X1 U899 ( .A1(n1196), .A2(n1156), .ZN(n1175) );
XOR2_X1 U900 ( .A(KEYINPUT35), .B(n1023), .Z(n1196) );
XOR2_X1 U901 ( .A(G113), .B(n1197), .Z(G15) );
NOR3_X1 U902 ( .A1(KEYINPUT18), .A2(n1198), .A3(n1199), .ZN(n1197) );
NOR2_X1 U903 ( .A1(KEYINPUT45), .A2(n1200), .ZN(n1199) );
NOR3_X1 U904 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
NOR2_X1 U905 ( .A1(n1134), .A2(n1204), .ZN(n1198) );
INV_X1 U906 ( .A(KEYINPUT45), .ZN(n1204) );
NOR3_X1 U907 ( .A1(n1202), .A2(n1195), .A3(n1203), .ZN(n1134) );
INV_X1 U908 ( .A(n994), .ZN(n1203) );
NOR2_X1 U909 ( .A1(n1156), .A2(n1159), .ZN(n994) );
INV_X1 U910 ( .A(n1201), .ZN(n1195) );
OR3_X1 U911 ( .A1(n1194), .A2(n1140), .A3(n997), .ZN(n1202) );
NAND2_X1 U912 ( .A1(n1184), .A2(n996), .ZN(n997) );
INV_X1 U913 ( .A(n1010), .ZN(n1194) );
NOR2_X1 U914 ( .A1(n1011), .A2(n1019), .ZN(n1010) );
XOR2_X1 U915 ( .A(G110), .B(n1205), .Z(G12) );
NOR2_X1 U916 ( .A1(n1140), .A2(n1206), .ZN(n1205) );
XNOR2_X1 U917 ( .A(KEYINPUT59), .B(n1141), .ZN(n1206) );
NAND4_X1 U918 ( .A1(n1012), .A2(n989), .A3(n1207), .A4(n1011), .ZN(n1141) );
INV_X1 U919 ( .A(n1179), .ZN(n1011) );
XOR2_X1 U920 ( .A(n1026), .B(n1025), .Z(n1179) );
XOR2_X1 U921 ( .A(G472), .B(KEYINPUT4), .Z(n1025) );
NAND2_X1 U922 ( .A1(n1208), .A2(n1209), .ZN(n1026) );
XOR2_X1 U923 ( .A(n1210), .B(n1211), .Z(n1208) );
XNOR2_X1 U924 ( .A(n1097), .B(n1212), .ZN(n1211) );
NOR2_X1 U925 ( .A1(KEYINPUT21), .A2(n1213), .ZN(n1212) );
XOR2_X1 U926 ( .A(KEYINPUT37), .B(n1105), .Z(n1213) );
XNOR2_X1 U927 ( .A(n1214), .B(n1215), .ZN(n1097) );
XNOR2_X1 U928 ( .A(G113), .B(n1216), .ZN(n1215) );
NAND2_X1 U929 ( .A1(G210), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U930 ( .A(n1218), .B(n1219), .ZN(n1214) );
XNOR2_X1 U931 ( .A(KEYINPUT54), .B(KEYINPUT20), .ZN(n1210) );
INV_X1 U932 ( .A(n1182), .ZN(n1207) );
NAND2_X1 U933 ( .A1(n988), .A2(n1201), .ZN(n1182) );
NAND2_X1 U934 ( .A1(n1220), .A2(n980), .ZN(n1201) );
NAND3_X1 U935 ( .A1(n1221), .A2(n1056), .A3(G952), .ZN(n980) );
NAND2_X1 U936 ( .A1(n1187), .A2(n1222), .ZN(n1220) );
INV_X1 U937 ( .A(G898), .ZN(n1222) );
AND3_X1 U938 ( .A1(G902), .A2(n1221), .A3(G953), .ZN(n1187) );
NAND2_X1 U939 ( .A1(G237), .A2(G234), .ZN(n1221) );
NOR2_X1 U940 ( .A1(n993), .A2(n1184), .ZN(n988) );
INV_X1 U941 ( .A(n990), .ZN(n1184) );
NAND2_X1 U942 ( .A1(n1223), .A2(n1224), .ZN(n990) );
NAND2_X1 U943 ( .A1(n1225), .A2(n1027), .ZN(n1224) );
XOR2_X1 U944 ( .A(KEYINPUT34), .B(n1226), .Z(n1223) );
NOR2_X1 U945 ( .A1(n1027), .A2(n1225), .ZN(n1226) );
XOR2_X1 U946 ( .A(KEYINPUT46), .B(n1028), .Z(n1225) );
INV_X1 U947 ( .A(G469), .ZN(n1028) );
AND4_X1 U948 ( .A1(n1227), .A2(n1209), .A3(n1228), .A4(n1229), .ZN(n1027) );
NAND2_X1 U949 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U950 ( .A(n1232), .B(n1108), .Z(n1230) );
OR3_X1 U951 ( .A1(n1108), .A2(n1232), .A3(n1231), .ZN(n1228) );
NAND3_X1 U952 ( .A1(n1111), .A2(n1108), .A3(n1232), .ZN(n1227) );
NOR2_X1 U953 ( .A1(KEYINPUT16), .A2(n1233), .ZN(n1232) );
XOR2_X1 U954 ( .A(n1234), .B(n1235), .Z(n1233) );
INV_X1 U955 ( .A(n1104), .ZN(n1235) );
XOR2_X1 U956 ( .A(n1236), .B(n1237), .Z(n1104) );
NOR2_X1 U957 ( .A1(KEYINPUT19), .A2(G107), .ZN(n1237) );
XNOR2_X1 U958 ( .A(G104), .B(KEYINPUT53), .ZN(n1236) );
XOR2_X1 U959 ( .A(n1238), .B(n1218), .Z(n1234) );
XNOR2_X1 U960 ( .A(n1044), .B(G101), .ZN(n1218) );
XOR2_X1 U961 ( .A(n1239), .B(n1042), .Z(n1044) );
XOR2_X1 U962 ( .A(G134), .B(G137), .Z(n1042) );
INV_X1 U963 ( .A(G131), .ZN(n1239) );
NAND2_X1 U964 ( .A1(KEYINPUT13), .A2(n1105), .ZN(n1238) );
INV_X1 U965 ( .A(n1045), .ZN(n1105) );
XOR2_X1 U966 ( .A(G140), .B(G110), .Z(n1108) );
INV_X1 U967 ( .A(n1231), .ZN(n1111) );
NAND2_X1 U968 ( .A1(G227), .A2(n1056), .ZN(n1231) );
INV_X1 U969 ( .A(n996), .ZN(n993) );
NAND2_X1 U970 ( .A1(G221), .A2(n1240), .ZN(n996) );
NOR2_X1 U971 ( .A1(n1156), .A2(n1023), .ZN(n989) );
INV_X1 U972 ( .A(n1159), .ZN(n1023) );
XOR2_X1 U973 ( .A(n1241), .B(G475), .Z(n1159) );
NAND2_X1 U974 ( .A1(n1090), .A2(n1209), .ZN(n1241) );
XNOR2_X1 U975 ( .A(n1242), .B(n1243), .ZN(n1090) );
XNOR2_X1 U976 ( .A(n1244), .B(n1245), .ZN(n1243) );
XOR2_X1 U977 ( .A(n1246), .B(G131), .Z(n1245) );
NAND2_X1 U978 ( .A1(G214), .A2(n1217), .ZN(n1246) );
NOR2_X1 U979 ( .A1(G953), .A2(G237), .ZN(n1217) );
XNOR2_X1 U980 ( .A(n1070), .B(n1039), .ZN(n1242) );
XNOR2_X1 U981 ( .A(n1188), .B(n1247), .ZN(n1070) );
INV_X1 U982 ( .A(G122), .ZN(n1188) );
OR2_X1 U983 ( .A1(n1248), .A2(n1017), .ZN(n1156) );
NOR3_X1 U984 ( .A1(G478), .A2(G902), .A3(n1022), .ZN(n1017) );
INV_X1 U985 ( .A(n1083), .ZN(n1022) );
AND2_X1 U986 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NAND2_X1 U987 ( .A1(n1083), .A2(n1209), .ZN(n1250) );
XOR2_X1 U988 ( .A(n1251), .B(n1252), .Z(n1083) );
XNOR2_X1 U989 ( .A(n1253), .B(n1254), .ZN(n1252) );
NAND2_X1 U990 ( .A1(n1255), .A2(KEYINPUT23), .ZN(n1253) );
XNOR2_X1 U991 ( .A(G107), .B(n1256), .ZN(n1255) );
XOR2_X1 U992 ( .A(G122), .B(G116), .Z(n1256) );
XOR2_X1 U993 ( .A(n1257), .B(n1258), .Z(n1251) );
XOR2_X1 U994 ( .A(G143), .B(G134), .Z(n1258) );
NAND3_X1 U995 ( .A1(G234), .A2(n1056), .A3(G217), .ZN(n1257) );
XOR2_X1 U996 ( .A(KEYINPUT30), .B(G478), .Z(n1249) );
XNOR2_X1 U997 ( .A(n1019), .B(KEYINPUT1), .ZN(n1012) );
XOR2_X1 U998 ( .A(n1259), .B(n1080), .Z(n1019) );
NAND2_X1 U999 ( .A1(G217), .A2(n1240), .ZN(n1080) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1209), .ZN(n1240) );
NAND2_X1 U1001 ( .A1(n1076), .A2(n1209), .ZN(n1259) );
XNOR2_X1 U1002 ( .A(n1260), .B(n1261), .ZN(n1076) );
XNOR2_X1 U1003 ( .A(n1262), .B(n1039), .ZN(n1261) );
XOR2_X1 U1004 ( .A(G140), .B(G125), .Z(n1039) );
NAND2_X1 U1005 ( .A1(KEYINPUT24), .A2(n1263), .ZN(n1262) );
XOR2_X1 U1006 ( .A(G137), .B(n1264), .Z(n1263) );
AND3_X1 U1007 ( .A1(G221), .A2(n1056), .A3(G234), .ZN(n1264) );
XOR2_X1 U1008 ( .A(n1265), .B(G146), .Z(n1260) );
NAND3_X1 U1009 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1265) );
NAND2_X1 U1010 ( .A1(G110), .A2(n1269), .ZN(n1268) );
NAND2_X1 U1011 ( .A1(n1270), .A2(n1271), .ZN(n1267) );
INV_X1 U1012 ( .A(KEYINPUT25), .ZN(n1271) );
NAND2_X1 U1013 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
INV_X1 U1014 ( .A(G110), .ZN(n1273) );
XNOR2_X1 U1015 ( .A(KEYINPUT28), .B(n1269), .ZN(n1272) );
NAND2_X1 U1016 ( .A1(KEYINPUT25), .A2(n1274), .ZN(n1266) );
NAND2_X1 U1017 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
OR3_X1 U1018 ( .A1(n1269), .A2(G110), .A3(KEYINPUT28), .ZN(n1276) );
NAND2_X1 U1019 ( .A1(KEYINPUT28), .A2(n1269), .ZN(n1275) );
XOR2_X1 U1020 ( .A(n1277), .B(n1278), .Z(n1269) );
NOR2_X1 U1021 ( .A1(KEYINPUT63), .A2(n1254), .ZN(n1278) );
NAND2_X1 U1022 ( .A1(n1006), .A2(n1007), .ZN(n1140) );
INV_X1 U1023 ( .A(n1178), .ZN(n1007) );
NOR2_X1 U1024 ( .A1(n1279), .A2(n1280), .ZN(n1178) );
INV_X1 U1025 ( .A(G214), .ZN(n1279) );
XNOR2_X1 U1026 ( .A(n1281), .B(n1282), .ZN(n1006) );
NOR2_X1 U1027 ( .A1(n1280), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U1028 ( .A(G210), .B(KEYINPUT38), .ZN(n1283) );
NOR2_X1 U1029 ( .A1(G902), .A2(G237), .ZN(n1280) );
NAND2_X1 U1030 ( .A1(n1284), .A2(n1209), .ZN(n1281) );
INV_X1 U1031 ( .A(G902), .ZN(n1209) );
XOR2_X1 U1032 ( .A(n1117), .B(n1285), .Z(n1284) );
XNOR2_X1 U1033 ( .A(n1145), .B(n1286), .ZN(n1285) );
NOR2_X1 U1034 ( .A1(KEYINPUT52), .A2(n1142), .ZN(n1286) );
INV_X1 U1035 ( .A(G125), .ZN(n1142) );
NAND2_X1 U1036 ( .A1(G224), .A2(n1056), .ZN(n1145) );
INV_X1 U1037 ( .A(G953), .ZN(n1056) );
XOR2_X1 U1038 ( .A(n1287), .B(n1288), .Z(n1117) );
XOR2_X1 U1039 ( .A(n1045), .B(n1289), .Z(n1288) );
XNOR2_X1 U1040 ( .A(KEYINPUT5), .B(n1290), .ZN(n1289) );
NOR2_X1 U1041 ( .A1(KEYINPUT10), .A2(n1291), .ZN(n1290) );
XOR2_X1 U1042 ( .A(G122), .B(n1068), .Z(n1291) );
XOR2_X1 U1043 ( .A(G110), .B(KEYINPUT0), .Z(n1068) );
XNOR2_X1 U1044 ( .A(n1254), .B(n1244), .ZN(n1045) );
XNOR2_X1 U1045 ( .A(n1152), .B(G146), .ZN(n1244) );
INV_X1 U1046 ( .A(G143), .ZN(n1152) );
XOR2_X1 U1047 ( .A(G128), .B(KEYINPUT12), .Z(n1254) );
XOR2_X1 U1048 ( .A(n1069), .B(n1247), .Z(n1287) );
XOR2_X1 U1049 ( .A(G104), .B(G113), .Z(n1247) );
XNOR2_X1 U1050 ( .A(n1219), .B(n1292), .ZN(n1069) );
XNOR2_X1 U1051 ( .A(G107), .B(n1293), .ZN(n1292) );
NAND2_X1 U1052 ( .A1(KEYINPUT14), .A2(n1181), .ZN(n1293) );
INV_X1 U1053 ( .A(G101), .ZN(n1181) );
XOR2_X1 U1054 ( .A(G116), .B(n1294), .Z(n1219) );
INV_X1 U1055 ( .A(n1277), .ZN(n1294) );
XNOR2_X1 U1056 ( .A(G119), .B(KEYINPUT57), .ZN(n1277) );
endmodule


