//Key = 0100110000100100000111001100111000100010011110010001110000001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353;

XNOR2_X1 U739 ( .A(G107), .B(n1026), .ZN(G9) );
NAND2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U741 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1031), .A2(n1032), .A3(G953), .A4(n1033), .ZN(n1030) );
NOR2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U744 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR3_X1 U745 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NOR2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U747 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U748 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U750 ( .A1(n1049), .A2(n1050), .ZN(n1041) );
NOR2_X1 U751 ( .A1(n1051), .A2(n1027), .ZN(n1049) );
NOR3_X1 U752 ( .A1(n1050), .A2(n1052), .A3(n1044), .ZN(n1036) );
INV_X1 U753 ( .A(n1053), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1056), .A2(n1040), .ZN(n1055) );
NOR2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U758 ( .A1(n1061), .A2(n1038), .ZN(n1054) );
NOR2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR3_X1 U761 ( .A1(n1033), .A2(G953), .A3(G952), .ZN(n1029) );
AND4_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1033) );
NOR4_X1 U763 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
XOR2_X1 U764 ( .A(n1074), .B(n1075), .Z(n1073) );
XNOR2_X1 U765 ( .A(KEYINPUT58), .B(n1076), .ZN(n1072) );
NOR3_X1 U766 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1068) );
INV_X1 U767 ( .A(n1060), .ZN(n1079) );
INV_X1 U768 ( .A(n1048), .ZN(n1078) );
NOR2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1077) );
XOR2_X1 U770 ( .A(n1082), .B(KEYINPUT31), .Z(n1081) );
XOR2_X1 U771 ( .A(n1083), .B(n1084), .Z(n1066) );
XOR2_X1 U772 ( .A(KEYINPUT15), .B(n1085), .Z(n1084) );
NOR2_X1 U773 ( .A1(G472), .A2(KEYINPUT45), .ZN(n1083) );
XOR2_X1 U774 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
AND2_X1 U776 ( .A1(G227), .A2(G900), .ZN(n1088) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1086) );
NAND3_X1 U778 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NAND2_X1 U779 ( .A1(n1095), .A2(n1089), .ZN(n1092) );
NAND2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1090) );
NAND2_X1 U781 ( .A1(n1094), .A2(n1093), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
XOR2_X1 U783 ( .A(KEYINPUT26), .B(n1100), .Z(n1098) );
XOR2_X1 U784 ( .A(n1101), .B(n1102), .Z(n1094) );
XNOR2_X1 U785 ( .A(n1103), .B(n1104), .ZN(n1102) );
NOR2_X1 U786 ( .A1(KEYINPUT57), .A2(n1105), .ZN(n1104) );
NAND2_X1 U787 ( .A1(KEYINPUT4), .A2(n1106), .ZN(n1103) );
XOR2_X1 U788 ( .A(KEYINPUT6), .B(n1107), .Z(n1096) );
NOR2_X1 U789 ( .A1(n1108), .A2(G953), .ZN(n1107) );
XOR2_X1 U790 ( .A(n1109), .B(n1110), .Z(G69) );
XOR2_X1 U791 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U792 ( .A1(KEYINPUT40), .A2(n1113), .ZN(n1112) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XNOR2_X1 U794 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
OR2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U797 ( .A(n1122), .B(KEYINPUT49), .Z(n1118) );
NAND2_X1 U798 ( .A1(n1121), .A2(n1120), .ZN(n1122) );
NOR2_X1 U799 ( .A1(G898), .A2(n1123), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1124), .A2(n1125), .ZN(n1111) );
XOR2_X1 U801 ( .A(n1089), .B(KEYINPUT10), .Z(n1125) );
NAND2_X1 U802 ( .A1(n1126), .A2(n1127), .ZN(n1109) );
NAND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1127) );
XOR2_X1 U804 ( .A(n1089), .B(KEYINPUT43), .Z(n1126) );
NOR2_X1 U805 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XNOR2_X1 U806 ( .A(n1130), .B(n1131), .ZN(n1129) );
NOR2_X1 U807 ( .A1(n1082), .A2(n1132), .ZN(n1131) );
NOR2_X1 U808 ( .A1(n1128), .A2(n1133), .ZN(G63) );
XOR2_X1 U809 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U810 ( .A1(KEYINPUT32), .A2(n1136), .ZN(n1135) );
XOR2_X1 U811 ( .A(KEYINPUT14), .B(n1137), .Z(n1136) );
NAND2_X1 U812 ( .A1(n1138), .A2(G478), .ZN(n1134) );
NOR2_X1 U813 ( .A1(n1128), .A2(n1139), .ZN(G60) );
XNOR2_X1 U814 ( .A(n1140), .B(n1141), .ZN(n1139) );
AND2_X1 U815 ( .A1(G475), .A2(n1138), .ZN(n1140) );
XNOR2_X1 U816 ( .A(G104), .B(n1142), .ZN(G6) );
NOR3_X1 U817 ( .A1(n1128), .A2(n1143), .A3(n1144), .ZN(G57) );
NOR2_X1 U818 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U819 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND2_X1 U820 ( .A1(KEYINPUT63), .A2(n1149), .ZN(n1147) );
NOR2_X1 U821 ( .A1(G101), .A2(n1150), .ZN(n1143) );
XOR2_X1 U822 ( .A(n1151), .B(n1148), .Z(n1150) );
XOR2_X1 U823 ( .A(n1121), .B(n1152), .Z(n1148) );
XOR2_X1 U824 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U825 ( .A1(KEYINPUT16), .A2(n1155), .ZN(n1154) );
AND2_X1 U826 ( .A1(G472), .A2(n1138), .ZN(n1153) );
NAND2_X1 U827 ( .A1(KEYINPUT63), .A2(n1156), .ZN(n1151) );
NOR3_X1 U828 ( .A1(n1128), .A2(n1157), .A3(n1158), .ZN(G54) );
NOR2_X1 U829 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U830 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U831 ( .A1(KEYINPUT50), .A2(n1163), .ZN(n1161) );
NOR2_X1 U832 ( .A1(n1164), .A2(n1165), .ZN(n1157) );
XOR2_X1 U833 ( .A(n1166), .B(n1162), .Z(n1165) );
XNOR2_X1 U834 ( .A(n1167), .B(n1168), .ZN(n1162) );
NOR2_X1 U835 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR3_X1 U836 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
INV_X1 U837 ( .A(KEYINPUT0), .ZN(n1171) );
NOR2_X1 U838 ( .A1(KEYINPUT0), .A2(n1174), .ZN(n1169) );
XOR2_X1 U839 ( .A(n1172), .B(n1105), .Z(n1174) );
INV_X1 U840 ( .A(n1173), .ZN(n1105) );
XOR2_X1 U841 ( .A(n1175), .B(n1176), .Z(n1167) );
AND2_X1 U842 ( .A1(G469), .A2(n1138), .ZN(n1176) );
NOR2_X1 U843 ( .A1(KEYINPUT50), .A2(n1177), .ZN(n1166) );
INV_X1 U844 ( .A(n1159), .ZN(n1164) );
NOR3_X1 U845 ( .A1(n1128), .A2(n1178), .A3(n1179), .ZN(G51) );
NOR2_X1 U846 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U847 ( .A(n1182), .B(KEYINPUT61), .Z(n1181) );
INV_X1 U848 ( .A(n1183), .ZN(n1180) );
NOR2_X1 U849 ( .A1(n1183), .A2(n1184), .ZN(n1178) );
XOR2_X1 U850 ( .A(n1182), .B(KEYINPUT37), .Z(n1184) );
NAND3_X1 U851 ( .A1(n1138), .A2(G210), .A3(KEYINPUT51), .ZN(n1182) );
INV_X1 U852 ( .A(n1132), .ZN(n1138) );
NAND2_X1 U853 ( .A1(G902), .A2(n1031), .ZN(n1132) );
NAND2_X1 U854 ( .A1(n1124), .A2(n1108), .ZN(n1031) );
INV_X1 U855 ( .A(n1095), .ZN(n1108) );
NAND4_X1 U856 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1095) );
AND4_X1 U857 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
NOR2_X1 U858 ( .A1(n1193), .A2(n1194), .ZN(n1187) );
INV_X1 U859 ( .A(n1195), .ZN(n1193) );
NAND3_X1 U860 ( .A1(n1051), .A2(n1058), .A3(n1196), .ZN(n1186) );
NAND2_X1 U861 ( .A1(n1197), .A2(n1198), .ZN(n1185) );
XOR2_X1 U862 ( .A(KEYINPUT22), .B(n1199), .Z(n1198) );
AND2_X1 U863 ( .A1(n1027), .A2(n1200), .ZN(n1199) );
AND4_X1 U864 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1124) );
AND4_X1 U865 ( .A1(n1205), .A2(n1206), .A3(n1142), .A4(n1207), .ZN(n1204) );
OR4_X1 U866 ( .A1(n1208), .A2(n1209), .A3(n1040), .A4(n1210), .ZN(n1207) );
INV_X1 U867 ( .A(n1027), .ZN(n1210) );
NOR2_X1 U868 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
INV_X1 U869 ( .A(KEYINPUT59), .ZN(n1212) );
NOR3_X1 U870 ( .A1(n1213), .A2(n1058), .A3(n1214), .ZN(n1211) );
NOR2_X1 U871 ( .A1(KEYINPUT59), .A2(n1215), .ZN(n1208) );
NAND2_X1 U872 ( .A1(n1051), .A2(n1028), .ZN(n1142) );
AND2_X1 U873 ( .A1(n1215), .A2(n1216), .ZN(n1028) );
NOR2_X1 U874 ( .A1(n1217), .A2(n1218), .ZN(n1203) );
INV_X1 U875 ( .A(n1219), .ZN(n1217) );
NAND2_X1 U876 ( .A1(n1220), .A2(n1221), .ZN(n1183) );
NAND3_X1 U877 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1221) );
INV_X1 U878 ( .A(KEYINPUT34), .ZN(n1224) );
NAND2_X1 U879 ( .A1(n1225), .A2(KEYINPUT34), .ZN(n1220) );
NOR2_X1 U880 ( .A1(n1089), .A2(G952), .ZN(n1128) );
XOR2_X1 U881 ( .A(n1226), .B(n1227), .Z(G48) );
XOR2_X1 U882 ( .A(KEYINPUT13), .B(G146), .Z(n1227) );
NAND4_X1 U883 ( .A1(KEYINPUT42), .A2(n1196), .A3(n1051), .A4(n1058), .ZN(n1226) );
XNOR2_X1 U884 ( .A(G143), .B(n1228), .ZN(G45) );
NAND2_X1 U885 ( .A1(n1194), .A2(n1229), .ZN(n1228) );
XOR2_X1 U886 ( .A(KEYINPUT60), .B(KEYINPUT2), .Z(n1229) );
AND3_X1 U887 ( .A1(n1230), .A2(n1058), .A3(n1200), .ZN(n1194) );
XNOR2_X1 U888 ( .A(G140), .B(n1192), .ZN(G42) );
NAND4_X1 U889 ( .A1(n1197), .A2(n1231), .A3(n1232), .A4(n1051), .ZN(n1192) );
XNOR2_X1 U890 ( .A(G137), .B(n1191), .ZN(G39) );
NAND3_X1 U891 ( .A1(n1196), .A2(n1053), .A3(n1197), .ZN(n1191) );
XNOR2_X1 U892 ( .A(G134), .B(n1233), .ZN(G36) );
NAND4_X1 U893 ( .A1(n1234), .A2(n1235), .A3(n1027), .A4(n1236), .ZN(n1233) );
NOR2_X1 U894 ( .A1(n1237), .A2(n1038), .ZN(n1236) );
XOR2_X1 U895 ( .A(KEYINPUT54), .B(n1046), .Z(n1234) );
INV_X1 U896 ( .A(n1213), .ZN(n1046) );
XNOR2_X1 U897 ( .A(G131), .B(n1190), .ZN(G33) );
NAND3_X1 U898 ( .A1(n1200), .A2(n1051), .A3(n1197), .ZN(n1190) );
INV_X1 U899 ( .A(n1038), .ZN(n1197) );
NAND2_X1 U900 ( .A1(n1238), .A2(n1060), .ZN(n1038) );
NOR3_X1 U901 ( .A1(n1213), .A2(n1239), .A3(n1237), .ZN(n1200) );
XOR2_X1 U902 ( .A(n1240), .B(n1189), .Z(G30) );
NAND3_X1 U903 ( .A1(n1027), .A2(n1058), .A3(n1196), .ZN(n1189) );
AND2_X1 U904 ( .A1(n1231), .A2(n1065), .ZN(n1196) );
NOR3_X1 U905 ( .A1(n1239), .A2(n1064), .A3(n1213), .ZN(n1231) );
INV_X1 U906 ( .A(n1241), .ZN(n1058) );
XOR2_X1 U907 ( .A(G101), .B(n1242), .Z(G3) );
NOR2_X1 U908 ( .A1(KEYINPUT35), .A2(n1206), .ZN(n1242) );
NAND3_X1 U909 ( .A1(n1215), .A2(n1053), .A3(n1063), .ZN(n1206) );
XOR2_X1 U910 ( .A(G125), .B(n1243), .Z(G27) );
NOR2_X1 U911 ( .A1(KEYINPUT27), .A2(n1195), .ZN(n1243) );
NAND4_X1 U912 ( .A1(n1232), .A2(n1244), .A3(n1051), .A4(n1245), .ZN(n1195) );
NOR3_X1 U913 ( .A1(n1241), .A2(n1064), .A3(n1239), .ZN(n1245) );
INV_X1 U914 ( .A(n1235), .ZN(n1239) );
NAND2_X1 U915 ( .A1(n1035), .A2(n1246), .ZN(n1235) );
NAND4_X1 U916 ( .A1(G902), .A2(n1100), .A3(n1247), .A4(n1099), .ZN(n1246) );
INV_X1 U917 ( .A(G900), .ZN(n1099) );
INV_X1 U918 ( .A(n1050), .ZN(n1244) );
XNOR2_X1 U919 ( .A(G122), .B(n1205), .ZN(G24) );
NAND3_X1 U920 ( .A1(n1248), .A2(n1216), .A3(n1230), .ZN(n1205) );
AND2_X1 U921 ( .A1(n1249), .A2(n1071), .ZN(n1230) );
XOR2_X1 U922 ( .A(n1250), .B(KEYINPUT20), .Z(n1249) );
INV_X1 U923 ( .A(n1040), .ZN(n1216) );
NAND2_X1 U924 ( .A1(n1064), .A2(n1232), .ZN(n1040) );
XNOR2_X1 U925 ( .A(G119), .B(n1201), .ZN(G21) );
NAND4_X1 U926 ( .A1(n1248), .A2(n1053), .A3(n1065), .A4(n1251), .ZN(n1201) );
XNOR2_X1 U927 ( .A(n1252), .B(n1202), .ZN(G18) );
NAND3_X1 U928 ( .A1(n1063), .A2(n1027), .A3(n1248), .ZN(n1202) );
NAND2_X1 U929 ( .A1(KEYINPUT1), .A2(n1253), .ZN(n1252) );
XOR2_X1 U930 ( .A(G113), .B(n1218), .Z(G15) );
AND3_X1 U931 ( .A1(n1051), .A2(n1063), .A3(n1248), .ZN(n1218) );
NOR3_X1 U932 ( .A1(n1241), .A2(n1214), .A3(n1050), .ZN(n1248) );
NAND2_X1 U933 ( .A1(n1254), .A2(n1048), .ZN(n1050) );
XOR2_X1 U934 ( .A(KEYINPUT12), .B(n1067), .Z(n1254) );
INV_X1 U935 ( .A(n1047), .ZN(n1067) );
INV_X1 U936 ( .A(n1237), .ZN(n1063) );
NAND2_X1 U937 ( .A1(n1064), .A2(n1065), .ZN(n1237) );
INV_X1 U938 ( .A(n1232), .ZN(n1065) );
INV_X1 U939 ( .A(n1251), .ZN(n1064) );
AND2_X1 U940 ( .A1(n1255), .A2(n1071), .ZN(n1051) );
XOR2_X1 U941 ( .A(n1250), .B(KEYINPUT7), .Z(n1255) );
XOR2_X1 U942 ( .A(G110), .B(n1256), .Z(G12) );
NOR2_X1 U943 ( .A1(KEYINPUT46), .A2(n1219), .ZN(n1256) );
NAND4_X1 U944 ( .A1(n1232), .A2(n1215), .A3(n1053), .A4(n1251), .ZN(n1219) );
NAND2_X1 U945 ( .A1(n1257), .A2(n1076), .ZN(n1251) );
NAND2_X1 U946 ( .A1(n1080), .A2(n1082), .ZN(n1076) );
OR2_X1 U947 ( .A1(n1082), .A2(n1080), .ZN(n1257) );
AND2_X1 U948 ( .A1(n1258), .A2(n1130), .ZN(n1080) );
NAND2_X1 U949 ( .A1(n1259), .A2(n1260), .ZN(n1130) );
NAND2_X1 U950 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U951 ( .A(KEYINPUT38), .B(n1263), .Z(n1259) );
NOR2_X1 U952 ( .A1(n1261), .A2(n1262), .ZN(n1263) );
XOR2_X1 U953 ( .A(n1264), .B(G137), .Z(n1262) );
NAND2_X1 U954 ( .A1(G221), .A2(n1265), .ZN(n1264) );
AND2_X1 U955 ( .A1(n1266), .A2(n1267), .ZN(n1261) );
NAND2_X1 U956 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U957 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U958 ( .A1(n1272), .A2(n1273), .ZN(n1268) );
NAND2_X1 U959 ( .A1(KEYINPUT41), .A2(n1274), .ZN(n1272) );
XNOR2_X1 U960 ( .A(n1275), .B(n1276), .ZN(n1274) );
NAND2_X1 U961 ( .A1(n1277), .A2(n1278), .ZN(n1266) );
NAND2_X1 U962 ( .A1(KEYINPUT41), .A2(n1279), .ZN(n1278) );
NAND3_X1 U963 ( .A1(n1271), .A2(n1273), .A3(n1270), .ZN(n1279) );
XOR2_X1 U964 ( .A(n1280), .B(KEYINPUT8), .Z(n1270) );
OR2_X1 U965 ( .A1(n1281), .A2(G146), .ZN(n1280) );
INV_X1 U966 ( .A(KEYINPUT9), .ZN(n1273) );
NAND2_X1 U967 ( .A1(G146), .A2(n1281), .ZN(n1271) );
XOR2_X1 U968 ( .A(n1275), .B(n1276), .Z(n1277) );
XOR2_X1 U969 ( .A(G119), .B(G110), .Z(n1276) );
NAND2_X1 U970 ( .A1(KEYINPUT29), .A2(n1240), .ZN(n1275) );
NAND2_X1 U971 ( .A1(G217), .A2(n1282), .ZN(n1082) );
NAND2_X1 U972 ( .A1(n1283), .A2(n1284), .ZN(n1053) );
OR3_X1 U973 ( .A1(n1071), .A2(n1070), .A3(KEYINPUT7), .ZN(n1284) );
INV_X1 U974 ( .A(n1250), .ZN(n1070) );
NAND2_X1 U975 ( .A1(KEYINPUT7), .A2(n1027), .ZN(n1283) );
NOR2_X1 U976 ( .A1(n1071), .A2(n1250), .ZN(n1027) );
XOR2_X1 U977 ( .A(n1285), .B(G478), .Z(n1250) );
OR2_X1 U978 ( .A1(n1137), .A2(G902), .ZN(n1285) );
XNOR2_X1 U979 ( .A(n1286), .B(n1287), .ZN(n1137) );
XOR2_X1 U980 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U981 ( .A(G107), .B(n1290), .Z(n1289) );
NOR2_X1 U982 ( .A1(KEYINPUT11), .A2(n1291), .ZN(n1290) );
XOR2_X1 U983 ( .A(G143), .B(G128), .Z(n1291) );
AND2_X1 U984 ( .A1(n1265), .A2(G217), .ZN(n1288) );
AND2_X1 U985 ( .A1(G234), .A2(n1089), .ZN(n1265) );
XOR2_X1 U986 ( .A(n1253), .B(n1292), .Z(n1286) );
XOR2_X1 U987 ( .A(G134), .B(G122), .Z(n1292) );
INV_X1 U988 ( .A(G116), .ZN(n1253) );
XNOR2_X1 U989 ( .A(n1293), .B(G475), .ZN(n1071) );
NAND2_X1 U990 ( .A1(n1294), .A2(n1141), .ZN(n1293) );
XOR2_X1 U991 ( .A(n1295), .B(n1296), .Z(n1141) );
XOR2_X1 U992 ( .A(G113), .B(n1297), .Z(n1296) );
XOR2_X1 U993 ( .A(KEYINPUT39), .B(G122), .Z(n1297) );
XOR2_X1 U994 ( .A(n1298), .B(G104), .Z(n1295) );
NAND3_X1 U995 ( .A1(n1299), .A2(n1300), .A3(KEYINPUT53), .ZN(n1298) );
NAND3_X1 U996 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1300) );
INV_X1 U997 ( .A(KEYINPUT25), .ZN(n1303) );
NAND2_X1 U998 ( .A1(n1304), .A2(KEYINPUT25), .ZN(n1299) );
XOR2_X1 U999 ( .A(n1302), .B(n1301), .Z(n1304) );
XNOR2_X1 U1000 ( .A(n1305), .B(G131), .ZN(n1301) );
NAND2_X1 U1001 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND4_X1 U1002 ( .A1(G214), .A2(G143), .A3(n1308), .A4(n1089), .ZN(n1307) );
NAND2_X1 U1003 ( .A1(n1309), .A2(n1310), .ZN(n1306) );
NAND3_X1 U1004 ( .A1(n1308), .A2(n1089), .A3(G214), .ZN(n1310) );
XOR2_X1 U1005 ( .A(KEYINPUT47), .B(G143), .Z(n1309) );
XOR2_X1 U1006 ( .A(G146), .B(n1281), .Z(n1302) );
XNOR2_X1 U1007 ( .A(n1106), .B(KEYINPUT56), .ZN(n1281) );
XNOR2_X1 U1008 ( .A(G125), .B(G140), .ZN(n1106) );
XOR2_X1 U1009 ( .A(n1258), .B(KEYINPUT55), .Z(n1294) );
NOR3_X1 U1010 ( .A1(n1213), .A2(n1214), .A3(n1241), .ZN(n1215) );
NAND2_X1 U1011 ( .A1(n1059), .A2(n1060), .ZN(n1241) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1311), .ZN(n1060) );
INV_X1 U1013 ( .A(n1238), .ZN(n1059) );
XOR2_X1 U1014 ( .A(n1074), .B(n1312), .Z(n1238) );
NOR2_X1 U1015 ( .A1(KEYINPUT48), .A2(n1075), .ZN(n1312) );
OR2_X1 U1016 ( .A1(n1225), .A2(G902), .ZN(n1075) );
XOR2_X1 U1017 ( .A(n1222), .B(n1223), .Z(n1225) );
XNOR2_X1 U1018 ( .A(n1313), .B(n1314), .ZN(n1223) );
XOR2_X1 U1019 ( .A(G125), .B(n1315), .Z(n1314) );
AND2_X1 U1020 ( .A1(n1089), .A2(G224), .ZN(n1315) );
XNOR2_X1 U1021 ( .A(n1316), .B(n1117), .ZN(n1222) );
XNOR2_X1 U1022 ( .A(n1317), .B(G122), .ZN(n1117) );
INV_X1 U1023 ( .A(G110), .ZN(n1317) );
XOR2_X1 U1024 ( .A(n1120), .B(n1121), .Z(n1316) );
NAND2_X1 U1025 ( .A1(n1318), .A2(n1319), .ZN(n1120) );
OR2_X1 U1026 ( .A1(n1320), .A2(G101), .ZN(n1319) );
XOR2_X1 U1027 ( .A(n1321), .B(KEYINPUT36), .Z(n1318) );
NAND2_X1 U1028 ( .A1(n1322), .A2(n1320), .ZN(n1321) );
XNOR2_X1 U1029 ( .A(n1323), .B(n1324), .ZN(n1320) );
NOR2_X1 U1030 ( .A1(KEYINPUT17), .A2(G107), .ZN(n1324) );
XNOR2_X1 U1031 ( .A(G104), .B(KEYINPUT24), .ZN(n1323) );
XOR2_X1 U1032 ( .A(n1145), .B(KEYINPUT28), .Z(n1322) );
NAND2_X1 U1033 ( .A1(G210), .A2(n1311), .ZN(n1074) );
NAND2_X1 U1034 ( .A1(n1308), .A2(n1258), .ZN(n1311) );
AND2_X1 U1035 ( .A1(n1035), .A2(n1325), .ZN(n1214) );
NAND4_X1 U1036 ( .A1(G902), .A2(n1100), .A3(n1247), .A4(n1326), .ZN(n1325) );
INV_X1 U1037 ( .A(G898), .ZN(n1326) );
INV_X1 U1038 ( .A(n1123), .ZN(n1100) );
XOR2_X1 U1039 ( .A(n1089), .B(KEYINPUT18), .Z(n1123) );
NAND3_X1 U1040 ( .A1(n1247), .A2(n1089), .A3(G952), .ZN(n1035) );
NAND2_X1 U1041 ( .A1(G237), .A2(G234), .ZN(n1247) );
NAND2_X1 U1042 ( .A1(n1047), .A2(n1048), .ZN(n1213) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1282), .ZN(n1048) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1258), .ZN(n1282) );
XOR2_X1 U1045 ( .A(n1327), .B(n1328), .Z(n1047) );
XOR2_X1 U1046 ( .A(KEYINPUT19), .B(G469), .Z(n1328) );
NAND2_X1 U1047 ( .A1(n1329), .A2(n1258), .ZN(n1327) );
XOR2_X1 U1048 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1049 ( .A(n1332), .B(n1159), .Z(n1331) );
NAND2_X1 U1050 ( .A1(G227), .A2(n1089), .ZN(n1159) );
NAND2_X1 U1051 ( .A1(n1333), .A2(KEYINPUT21), .ZN(n1332) );
XOR2_X1 U1052 ( .A(n1175), .B(n1334), .Z(n1333) );
NOR2_X1 U1053 ( .A1(KEYINPUT33), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1054 ( .A(n1172), .B(n1173), .Z(n1335) );
XNOR2_X1 U1055 ( .A(n1336), .B(n1337), .ZN(n1173) );
NOR2_X1 U1056 ( .A1(G128), .A2(KEYINPUT23), .ZN(n1337) );
XNOR2_X1 U1057 ( .A(n1145), .B(n1338), .ZN(n1172) );
XOR2_X1 U1058 ( .A(G107), .B(G104), .Z(n1338) );
INV_X1 U1059 ( .A(G101), .ZN(n1145) );
NAND2_X1 U1060 ( .A1(KEYINPUT52), .A2(n1163), .ZN(n1330) );
INV_X1 U1061 ( .A(n1177), .ZN(n1163) );
XOR2_X1 U1062 ( .A(G140), .B(G110), .Z(n1177) );
XOR2_X1 U1063 ( .A(n1339), .B(G472), .Z(n1232) );
NAND2_X1 U1064 ( .A1(KEYINPUT30), .A2(n1085), .ZN(n1339) );
AND2_X1 U1065 ( .A1(n1340), .A2(n1258), .ZN(n1085) );
INV_X1 U1066 ( .A(G902), .ZN(n1258) );
NAND2_X1 U1067 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1068 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XOR2_X1 U1069 ( .A(KEYINPUT62), .B(n1345), .Z(n1344) );
XOR2_X1 U1070 ( .A(n1155), .B(n1121), .Z(n1343) );
INV_X1 U1071 ( .A(n1346), .ZN(n1121) );
NAND2_X1 U1072 ( .A1(n1347), .A2(n1348), .ZN(n1341) );
XOR2_X1 U1073 ( .A(n1346), .B(n1155), .Z(n1348) );
XOR2_X1 U1074 ( .A(n1313), .B(n1101), .Z(n1155) );
INV_X1 U1075 ( .A(n1175), .ZN(n1101) );
XNOR2_X1 U1076 ( .A(G131), .B(n1349), .ZN(n1175) );
XOR2_X1 U1077 ( .A(G137), .B(G134), .Z(n1349) );
XOR2_X1 U1078 ( .A(n1240), .B(n1336), .Z(n1313) );
XOR2_X1 U1079 ( .A(G143), .B(G146), .Z(n1336) );
INV_X1 U1080 ( .A(G128), .ZN(n1240) );
XOR2_X1 U1081 ( .A(n1350), .B(n1351), .Z(n1346) );
XOR2_X1 U1082 ( .A(KEYINPUT44), .B(G119), .Z(n1351) );
XOR2_X1 U1083 ( .A(n1352), .B(G116), .Z(n1350) );
INV_X1 U1084 ( .A(G113), .ZN(n1352) );
XOR2_X1 U1085 ( .A(KEYINPUT5), .B(n1345), .Z(n1347) );
XOR2_X1 U1086 ( .A(n1156), .B(n1353), .Z(n1345) );
NOR2_X1 U1087 ( .A1(G101), .A2(KEYINPUT3), .ZN(n1353) );
INV_X1 U1088 ( .A(n1149), .ZN(n1156) );
NAND3_X1 U1089 ( .A1(n1308), .A2(n1089), .A3(G210), .ZN(n1149) );
INV_X1 U1090 ( .A(G953), .ZN(n1089) );
INV_X1 U1091 ( .A(G237), .ZN(n1308) );
endmodule


