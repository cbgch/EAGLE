//Key = 1101100001101101111010001110111101011110001111110000111101111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334;

XOR2_X1 U733 ( .A(n1013), .B(n1014), .Z(G9) );
NAND2_X1 U734 ( .A1(KEYINPUT35), .A2(G107), .ZN(n1014) );
NOR2_X1 U735 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR3_X1 U736 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
INV_X1 U737 ( .A(n1020), .ZN(n1019) );
NOR3_X1 U738 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1018) );
NOR2_X1 U739 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR3_X1 U740 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NOR2_X1 U741 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR2_X1 U742 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1029) );
NOR2_X1 U745 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
AND2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1024) );
NAND3_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1017) );
NAND4_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
NOR3_X1 U750 ( .A1(n1032), .A2(n1036), .A3(n1026), .ZN(n1049) );
INV_X1 U751 ( .A(n1041), .ZN(n1036) );
INV_X1 U752 ( .A(n1021), .ZN(n1048) );
NAND2_X1 U753 ( .A1(n1027), .A2(n1023), .ZN(n1047) );
OR3_X1 U754 ( .A1(n1050), .A2(n1051), .A3(n1027), .ZN(n1046) );
NOR3_X1 U755 ( .A1(n1052), .A2(G953), .A3(G952), .ZN(n1015) );
INV_X1 U756 ( .A(n1043), .ZN(n1052) );
NAND4_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1043) );
NOR4_X1 U758 ( .A1(n1027), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1056) );
NOR3_X1 U759 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1055) );
NOR2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U761 ( .A1(G472), .A2(n1065), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
AND2_X1 U763 ( .A1(n1063), .A2(KEYINPUT43), .ZN(n1067) );
NAND2_X1 U764 ( .A1(KEYINPUT17), .A2(n1068), .ZN(n1063) );
NOR2_X1 U765 ( .A1(KEYINPUT43), .A2(n1069), .ZN(n1066) );
XNOR2_X1 U766 ( .A(n1070), .B(n1071), .ZN(n1060) );
XNOR2_X1 U767 ( .A(n1072), .B(G475), .ZN(n1054) );
XOR2_X1 U768 ( .A(n1073), .B(G469), .Z(n1053) );
XOR2_X1 U769 ( .A(n1074), .B(n1075), .Z(G72) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
AND2_X1 U771 ( .A1(G227), .A2(G900), .ZN(n1076) );
NAND2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
NAND2_X1 U773 ( .A1(n1080), .A2(n1044), .ZN(n1079) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND3_X1 U775 ( .A1(G900), .A2(n1082), .A3(G953), .ZN(n1078) );
XOR2_X1 U776 ( .A(n1083), .B(n1084), .Z(n1082) );
XNOR2_X1 U777 ( .A(n1085), .B(n1086), .ZN(n1083) );
NOR2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U779 ( .A1(KEYINPUT9), .A2(n1089), .ZN(n1088) );
AND2_X1 U780 ( .A1(KEYINPUT18), .A2(n1089), .ZN(n1087) );
XOR2_X1 U781 ( .A(n1090), .B(n1091), .Z(G69) );
XOR2_X1 U782 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1095) );
INV_X1 U785 ( .A(n1077), .ZN(n1094) );
XOR2_X1 U786 ( .A(G953), .B(KEYINPUT42), .Z(n1077) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
NAND2_X1 U788 ( .A1(G953), .A2(n1098), .ZN(n1097) );
XNOR2_X1 U789 ( .A(n1099), .B(n1100), .ZN(n1096) );
XNOR2_X1 U790 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR3_X1 U791 ( .A1(n1103), .A2(KEYINPUT56), .A3(G953), .ZN(n1090) );
NOR2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U793 ( .A1(n1106), .A2(n1107), .ZN(G66) );
XOR2_X1 U794 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U795 ( .A1(n1110), .A2(n1071), .ZN(n1109) );
INV_X1 U796 ( .A(n1111), .ZN(n1071) );
NAND2_X1 U797 ( .A1(KEYINPUT26), .A2(n1112), .ZN(n1108) );
INV_X1 U798 ( .A(n1113), .ZN(n1112) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1115), .ZN(G63) );
XOR2_X1 U800 ( .A(KEYINPUT11), .B(n1106), .Z(n1115) );
XOR2_X1 U801 ( .A(n1116), .B(n1117), .Z(n1114) );
NAND2_X1 U802 ( .A1(n1110), .A2(G478), .ZN(n1116) );
NOR2_X1 U803 ( .A1(n1106), .A2(n1118), .ZN(G60) );
NOR3_X1 U804 ( .A1(n1072), .A2(n1119), .A3(n1120), .ZN(n1118) );
AND3_X1 U805 ( .A1(n1121), .A2(G475), .A3(n1110), .ZN(n1120) );
NOR2_X1 U806 ( .A1(n1122), .A2(n1121), .ZN(n1119) );
NOR2_X1 U807 ( .A1(n1020), .A2(n1123), .ZN(n1122) );
XOR2_X1 U808 ( .A(G104), .B(n1124), .Z(G6) );
NOR2_X1 U809 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U810 ( .A1(n1106), .A2(n1127), .ZN(G57) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
XNOR2_X1 U812 ( .A(n1130), .B(n1131), .ZN(n1129) );
NAND3_X1 U813 ( .A1(n1132), .A2(n1133), .A3(KEYINPUT12), .ZN(n1130) );
NAND2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
INV_X1 U815 ( .A(G101), .ZN(n1135) );
XOR2_X1 U816 ( .A(n1136), .B(n1137), .Z(n1128) );
NAND4_X1 U817 ( .A1(KEYINPUT58), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1137) );
NAND3_X1 U818 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
INV_X1 U819 ( .A(KEYINPUT48), .ZN(n1142) );
OR2_X1 U820 ( .A1(n1143), .A2(n1141), .ZN(n1139) );
NOR2_X1 U821 ( .A1(KEYINPUT32), .A2(n1085), .ZN(n1141) );
NAND2_X1 U822 ( .A1(KEYINPUT48), .A2(n1085), .ZN(n1138) );
NAND2_X1 U823 ( .A1(n1144), .A2(n1110), .ZN(n1136) );
XNOR2_X1 U824 ( .A(G472), .B(KEYINPUT55), .ZN(n1144) );
NOR2_X1 U825 ( .A1(n1106), .A2(n1145), .ZN(G54) );
XOR2_X1 U826 ( .A(n1146), .B(n1147), .Z(n1145) );
AND2_X1 U827 ( .A1(G469), .A2(n1110), .ZN(n1147) );
NOR2_X1 U828 ( .A1(KEYINPUT7), .A2(n1148), .ZN(n1146) );
XOR2_X1 U829 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U831 ( .A(KEYINPUT15), .B(G110), .Z(n1152) );
XOR2_X1 U832 ( .A(n1153), .B(n1154), .Z(n1149) );
NOR2_X1 U833 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
AND2_X1 U834 ( .A1(KEYINPUT45), .A2(n1157), .ZN(n1156) );
NOR2_X1 U835 ( .A1(KEYINPUT31), .A2(n1157), .ZN(n1155) );
XNOR2_X1 U836 ( .A(n1158), .B(n1159), .ZN(n1153) );
NAND2_X1 U837 ( .A1(n1160), .A2(KEYINPUT13), .ZN(n1158) );
XNOR2_X1 U838 ( .A(n1161), .B(n1143), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1106), .A2(n1162), .ZN(G51) );
XOR2_X1 U840 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U841 ( .A(n1165), .B(n1166), .Z(n1163) );
NOR2_X1 U842 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U843 ( .A(KEYINPUT23), .B(n1169), .Z(n1168) );
NOR2_X1 U844 ( .A1(n1084), .A2(n1170), .ZN(n1169) );
AND2_X1 U845 ( .A1(n1084), .A2(n1170), .ZN(n1167) );
XOR2_X1 U846 ( .A(n1171), .B(KEYINPUT33), .Z(n1170) );
NAND2_X1 U847 ( .A1(n1110), .A2(n1172), .ZN(n1165) );
NOR2_X1 U848 ( .A1(n1173), .A2(n1020), .ZN(n1110) );
NOR3_X1 U849 ( .A1(n1081), .A2(n1105), .A3(n1174), .ZN(n1020) );
XOR2_X1 U850 ( .A(n1104), .B(KEYINPUT6), .Z(n1174) );
NAND4_X1 U851 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1105) );
AND4_X1 U852 ( .A1(n1013), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1178) );
NAND3_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1034), .ZN(n1013) );
NOR2_X1 U854 ( .A1(n1184), .A2(n1185), .ZN(n1177) );
NOR2_X1 U855 ( .A1(KEYINPUT22), .A2(n1186), .ZN(n1185) );
INV_X1 U856 ( .A(n1187), .ZN(n1184) );
NAND4_X1 U857 ( .A1(KEYINPUT22), .A2(n1188), .A3(n1189), .A4(n1125), .ZN(n1176) );
AND3_X1 U858 ( .A1(n1033), .A2(n1190), .A3(n1051), .ZN(n1189) );
NAND2_X1 U859 ( .A1(n1191), .A2(n1192), .ZN(n1175) );
XOR2_X1 U860 ( .A(n1126), .B(KEYINPUT16), .Z(n1191) );
NAND4_X1 U861 ( .A1(n1033), .A2(n1182), .A3(n1038), .A4(n1190), .ZN(n1126) );
NAND4_X1 U862 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1081) );
NOR4_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196) );
INV_X1 U864 ( .A(n1201), .ZN(n1200) );
NOR2_X1 U865 ( .A1(n1202), .A2(n1203), .ZN(n1195) );
NOR2_X1 U866 ( .A1(n1204), .A2(n1125), .ZN(n1203) );
XOR2_X1 U867 ( .A(n1205), .B(KEYINPUT62), .Z(n1204) );
NAND3_X1 U868 ( .A1(n1206), .A2(n1034), .A3(n1207), .ZN(n1194) );
NOR2_X1 U869 ( .A1(n1044), .A2(G952), .ZN(n1106) );
XNOR2_X1 U870 ( .A(G146), .B(n1201), .ZN(G48) );
NAND3_X1 U871 ( .A1(n1033), .A2(n1206), .A3(n1207), .ZN(n1201) );
XOR2_X1 U872 ( .A(G143), .B(n1208), .Z(G45) );
NOR2_X1 U873 ( .A1(n1125), .A2(n1205), .ZN(n1208) );
NAND4_X1 U874 ( .A1(n1051), .A2(n1206), .A3(n1209), .A4(n1059), .ZN(n1205) );
INV_X1 U875 ( .A(n1210), .ZN(n1206) );
XOR2_X1 U876 ( .A(G140), .B(n1199), .Z(G42) );
AND3_X1 U877 ( .A1(n1033), .A2(n1211), .A3(n1050), .ZN(n1199) );
XOR2_X1 U878 ( .A(G137), .B(n1198), .Z(G39) );
AND4_X1 U879 ( .A1(n1212), .A2(n1041), .A3(n1211), .A4(n1213), .ZN(n1198) );
NAND2_X1 U880 ( .A1(n1214), .A2(n1215), .ZN(G36) );
NAND2_X1 U881 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XNOR2_X1 U882 ( .A(n1202), .B(KEYINPUT44), .ZN(n1216) );
INV_X1 U883 ( .A(n1218), .ZN(n1202) );
NAND2_X1 U884 ( .A1(n1219), .A2(G134), .ZN(n1214) );
XNOR2_X1 U885 ( .A(KEYINPUT25), .B(n1218), .ZN(n1219) );
NAND3_X1 U886 ( .A1(n1211), .A2(n1034), .A3(n1051), .ZN(n1218) );
XOR2_X1 U887 ( .A(G131), .B(n1197), .Z(G33) );
AND3_X1 U888 ( .A1(n1051), .A2(n1211), .A3(n1033), .ZN(n1197) );
NOR3_X1 U889 ( .A1(n1026), .A2(n1027), .A3(n1210), .ZN(n1211) );
NAND2_X1 U890 ( .A1(n1038), .A2(n1220), .ZN(n1210) );
XOR2_X1 U891 ( .A(n1058), .B(KEYINPUT27), .Z(n1026) );
XNOR2_X1 U892 ( .A(G128), .B(n1221), .ZN(G30) );
NAND4_X1 U893 ( .A1(n1222), .A2(n1207), .A3(n1034), .A4(n1220), .ZN(n1221) );
XNOR2_X1 U894 ( .A(n1038), .B(KEYINPUT4), .ZN(n1222) );
INV_X1 U895 ( .A(n1223), .ZN(n1038) );
XNOR2_X1 U896 ( .A(G101), .B(n1187), .ZN(G3) );
NAND3_X1 U897 ( .A1(n1051), .A2(n1183), .A3(n1041), .ZN(n1187) );
XNOR2_X1 U898 ( .A(G125), .B(n1193), .ZN(G27) );
NAND4_X1 U899 ( .A1(n1042), .A2(n1050), .A3(n1033), .A4(n1220), .ZN(n1193) );
NAND2_X1 U900 ( .A1(n1021), .A2(n1224), .ZN(n1220) );
NAND2_X1 U901 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
INV_X1 U902 ( .A(G900), .ZN(n1226) );
XOR2_X1 U903 ( .A(G122), .B(n1104), .Z(G24) );
AND3_X1 U904 ( .A1(n1209), .A2(n1042), .A3(n1227), .ZN(n1104) );
NOR3_X1 U905 ( .A1(n1023), .A2(n1228), .A3(n1229), .ZN(n1227) );
INV_X1 U906 ( .A(n1182), .ZN(n1023) );
NOR2_X1 U907 ( .A1(n1213), .A2(n1212), .ZN(n1182) );
XOR2_X1 U908 ( .A(n1230), .B(G119), .Z(G21) );
NAND2_X1 U909 ( .A1(KEYINPUT28), .A2(n1181), .ZN(n1230) );
NAND4_X1 U910 ( .A1(n1188), .A2(n1207), .A3(n1041), .A4(n1190), .ZN(n1181) );
AND3_X1 U911 ( .A1(n1192), .A2(n1213), .A3(n1212), .ZN(n1207) );
INV_X1 U912 ( .A(n1231), .ZN(n1212) );
XNOR2_X1 U913 ( .A(G116), .B(n1180), .ZN(G18) );
NAND4_X1 U914 ( .A1(n1042), .A2(n1051), .A3(n1034), .A4(n1190), .ZN(n1180) );
NOR2_X1 U915 ( .A1(n1229), .A2(n1209), .ZN(n1034) );
INV_X1 U916 ( .A(n1059), .ZN(n1229) );
XNOR2_X1 U917 ( .A(n1186), .B(n1232), .ZN(G15) );
NOR2_X1 U918 ( .A1(KEYINPUT34), .A2(n1233), .ZN(n1232) );
NAND4_X1 U919 ( .A1(n1042), .A2(n1033), .A3(n1051), .A4(n1190), .ZN(n1186) );
AND2_X1 U920 ( .A1(n1231), .A2(n1213), .ZN(n1051) );
NOR2_X1 U921 ( .A1(n1234), .A2(n1059), .ZN(n1033) );
NOR2_X1 U922 ( .A1(n1032), .A2(n1125), .ZN(n1042) );
INV_X1 U923 ( .A(n1188), .ZN(n1032) );
NOR2_X1 U924 ( .A1(n1039), .A2(n1057), .ZN(n1188) );
INV_X1 U925 ( .A(n1040), .ZN(n1057) );
XOR2_X1 U926 ( .A(n1179), .B(n1235), .Z(G12) );
NAND2_X1 U927 ( .A1(n1236), .A2(G110), .ZN(n1235) );
XNOR2_X1 U928 ( .A(KEYINPUT59), .B(KEYINPUT53), .ZN(n1236) );
NAND3_X1 U929 ( .A1(n1041), .A2(n1183), .A3(n1050), .ZN(n1179) );
NOR2_X1 U930 ( .A1(n1231), .A2(n1213), .ZN(n1050) );
XNOR2_X1 U931 ( .A(n1069), .B(n1064), .ZN(n1213) );
INV_X1 U932 ( .A(G472), .ZN(n1064) );
INV_X1 U933 ( .A(n1068), .ZN(n1069) );
NAND2_X1 U934 ( .A1(n1237), .A2(n1173), .ZN(n1068) );
XOR2_X1 U935 ( .A(n1238), .B(n1239), .Z(n1237) );
XNOR2_X1 U936 ( .A(n1240), .B(n1241), .ZN(n1239) );
INV_X1 U937 ( .A(n1131), .ZN(n1241) );
XNOR2_X1 U938 ( .A(n1242), .B(KEYINPUT10), .ZN(n1131) );
NAND2_X1 U939 ( .A1(n1243), .A2(n1244), .ZN(n1240) );
NAND2_X1 U940 ( .A1(n1143), .A2(n1085), .ZN(n1244) );
XOR2_X1 U941 ( .A(n1245), .B(KEYINPUT63), .Z(n1243) );
NAND2_X1 U942 ( .A1(n1159), .A2(n1246), .ZN(n1245) );
INV_X1 U943 ( .A(n1085), .ZN(n1159) );
XOR2_X1 U944 ( .A(n1247), .B(KEYINPUT41), .Z(n1238) );
NAND2_X1 U945 ( .A1(n1133), .A2(n1248), .ZN(n1247) );
NAND2_X1 U946 ( .A1(n1249), .A2(n1134), .ZN(n1248) );
INV_X1 U947 ( .A(n1250), .ZN(n1134) );
XNOR2_X1 U948 ( .A(G101), .B(KEYINPUT21), .ZN(n1249) );
NAND2_X1 U949 ( .A1(G101), .A2(n1250), .ZN(n1133) );
NAND3_X1 U950 ( .A1(n1251), .A2(n1044), .A3(G210), .ZN(n1250) );
XOR2_X1 U951 ( .A(n1252), .B(n1111), .Z(n1231) );
NAND2_X1 U952 ( .A1(G217), .A2(n1253), .ZN(n1111) );
NAND2_X1 U953 ( .A1(KEYINPUT20), .A2(n1070), .ZN(n1252) );
NAND2_X1 U954 ( .A1(n1113), .A2(n1173), .ZN(n1070) );
NAND2_X1 U955 ( .A1(n1254), .A2(n1255), .ZN(n1113) );
NAND2_X1 U956 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XNOR2_X1 U957 ( .A(G137), .B(n1258), .ZN(n1257) );
XOR2_X1 U958 ( .A(n1259), .B(n1260), .Z(n1256) );
XOR2_X1 U959 ( .A(n1261), .B(KEYINPUT14), .Z(n1254) );
NAND2_X1 U960 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U961 ( .A(n1260), .B(n1259), .ZN(n1263) );
XNOR2_X1 U962 ( .A(n1264), .B(n1265), .ZN(n1259) );
XOR2_X1 U963 ( .A(G119), .B(n1266), .Z(n1265) );
XOR2_X1 U964 ( .A(n1267), .B(n1268), .Z(n1260) );
XNOR2_X1 U965 ( .A(KEYINPUT40), .B(KEYINPUT38), .ZN(n1267) );
XOR2_X1 U966 ( .A(n1258), .B(G137), .Z(n1262) );
NAND3_X1 U967 ( .A1(G221), .A2(n1269), .A3(KEYINPUT52), .ZN(n1258) );
INV_X1 U968 ( .A(n1270), .ZN(n1269) );
NOR3_X1 U969 ( .A1(n1223), .A2(n1228), .A3(n1125), .ZN(n1183) );
INV_X1 U970 ( .A(n1192), .ZN(n1125) );
NOR2_X1 U971 ( .A1(n1271), .A2(n1027), .ZN(n1192) );
AND2_X1 U972 ( .A1(G214), .A2(n1272), .ZN(n1027) );
INV_X1 U973 ( .A(n1058), .ZN(n1271) );
XNOR2_X1 U974 ( .A(n1273), .B(n1172), .ZN(n1058) );
AND2_X1 U975 ( .A1(G210), .A2(n1272), .ZN(n1172) );
NAND2_X1 U976 ( .A1(n1173), .A2(n1251), .ZN(n1272) );
NAND2_X1 U977 ( .A1(n1274), .A2(n1173), .ZN(n1273) );
XNOR2_X1 U978 ( .A(n1164), .B(n1275), .ZN(n1274) );
XNOR2_X1 U979 ( .A(n1276), .B(n1084), .ZN(n1275) );
XNOR2_X1 U980 ( .A(G125), .B(n1246), .ZN(n1084) );
NAND2_X1 U981 ( .A1(KEYINPUT24), .A2(n1171), .ZN(n1276) );
AND2_X1 U982 ( .A1(G224), .A2(n1044), .ZN(n1171) );
XNOR2_X1 U983 ( .A(n1277), .B(n1102), .ZN(n1164) );
XOR2_X1 U984 ( .A(G110), .B(G122), .Z(n1102) );
NAND2_X1 U985 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NAND2_X1 U986 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U987 ( .A1(KEYINPUT3), .A2(n1282), .ZN(n1281) );
NAND2_X1 U988 ( .A1(KEYINPUT54), .A2(n1161), .ZN(n1282) );
NAND2_X1 U989 ( .A1(n1101), .A2(n1283), .ZN(n1278) );
NAND2_X1 U990 ( .A1(KEYINPUT54), .A2(n1284), .ZN(n1283) );
NAND2_X1 U991 ( .A1(n1099), .A2(KEYINPUT3), .ZN(n1284) );
INV_X1 U992 ( .A(n1280), .ZN(n1099) );
XNOR2_X1 U993 ( .A(n1242), .B(KEYINPUT57), .ZN(n1280) );
XNOR2_X1 U994 ( .A(G113), .B(n1285), .ZN(n1242) );
XOR2_X1 U995 ( .A(G119), .B(G116), .Z(n1285) );
INV_X1 U996 ( .A(n1161), .ZN(n1101) );
INV_X1 U997 ( .A(n1190), .ZN(n1228) );
NAND2_X1 U998 ( .A1(n1021), .A2(n1286), .ZN(n1190) );
NAND2_X1 U999 ( .A1(n1225), .A2(n1098), .ZN(n1286) );
INV_X1 U1000 ( .A(G898), .ZN(n1098) );
AND3_X1 U1001 ( .A1(G953), .A2(n1287), .A3(n1288), .ZN(n1225) );
XNOR2_X1 U1002 ( .A(G902), .B(KEYINPUT0), .ZN(n1288) );
NAND3_X1 U1003 ( .A1(n1287), .A2(n1044), .A3(G952), .ZN(n1021) );
NAND2_X1 U1004 ( .A1(G234), .A2(G237), .ZN(n1287) );
NAND2_X1 U1005 ( .A1(n1039), .A2(n1040), .ZN(n1223) );
NAND2_X1 U1006 ( .A1(G221), .A2(n1253), .ZN(n1040) );
NAND2_X1 U1007 ( .A1(G234), .A2(n1173), .ZN(n1253) );
NAND2_X1 U1008 ( .A1(n1289), .A2(n1290), .ZN(n1039) );
OR2_X1 U1009 ( .A1(n1073), .A2(G469), .ZN(n1290) );
NAND2_X1 U1010 ( .A1(n1291), .A2(G469), .ZN(n1289) );
XNOR2_X1 U1011 ( .A(KEYINPUT29), .B(n1073), .ZN(n1291) );
NAND2_X1 U1012 ( .A1(n1292), .A2(n1173), .ZN(n1073) );
XOR2_X1 U1013 ( .A(n1293), .B(n1266), .Z(n1292) );
XNOR2_X1 U1014 ( .A(G110), .B(n1157), .ZN(n1266) );
XOR2_X1 U1015 ( .A(n1294), .B(n1151), .Z(n1293) );
AND2_X1 U1016 ( .A1(n1295), .A2(G227), .ZN(n1151) );
XNOR2_X1 U1017 ( .A(G953), .B(KEYINPUT5), .ZN(n1295) );
NAND2_X1 U1018 ( .A1(n1296), .A2(n1297), .ZN(n1294) );
XOR2_X1 U1019 ( .A(KEYINPUT51), .B(KEYINPUT47), .Z(n1297) );
XOR2_X1 U1020 ( .A(n1298), .B(n1299), .Z(n1296) );
XNOR2_X1 U1021 ( .A(n1300), .B(KEYINPUT46), .ZN(n1299) );
NAND2_X1 U1022 ( .A1(KEYINPUT37), .A2(n1143), .ZN(n1300) );
INV_X1 U1023 ( .A(n1246), .ZN(n1143) );
XNOR2_X1 U1024 ( .A(G143), .B(n1264), .ZN(n1246) );
XOR2_X1 U1025 ( .A(G146), .B(G128), .Z(n1264) );
XNOR2_X1 U1026 ( .A(n1085), .B(n1161), .ZN(n1298) );
XOR2_X1 U1027 ( .A(G101), .B(n1301), .Z(n1161) );
XOR2_X1 U1028 ( .A(G107), .B(G104), .Z(n1301) );
XOR2_X1 U1029 ( .A(G131), .B(n1302), .Z(n1085) );
XNOR2_X1 U1030 ( .A(G137), .B(n1217), .ZN(n1302) );
NOR2_X1 U1031 ( .A1(n1059), .A2(n1209), .ZN(n1041) );
INV_X1 U1032 ( .A(n1234), .ZN(n1209) );
XNOR2_X1 U1033 ( .A(n1303), .B(n1304), .ZN(n1234) );
XOR2_X1 U1034 ( .A(KEYINPUT50), .B(n1072), .Z(n1304) );
NOR2_X1 U1035 ( .A1(n1121), .A2(G902), .ZN(n1072) );
XNOR2_X1 U1036 ( .A(n1305), .B(n1306), .ZN(n1121) );
XOR2_X1 U1037 ( .A(G131), .B(n1307), .Z(n1306) );
XNOR2_X1 U1038 ( .A(n1308), .B(G143), .ZN(n1307) );
INV_X1 U1039 ( .A(G146), .ZN(n1308) );
XOR2_X1 U1040 ( .A(n1309), .B(n1310), .Z(n1305) );
NOR3_X1 U1041 ( .A1(n1311), .A2(G953), .A3(n1312), .ZN(n1310) );
INV_X1 U1042 ( .A(G214), .ZN(n1312) );
XNOR2_X1 U1043 ( .A(KEYINPUT39), .B(n1251), .ZN(n1311) );
INV_X1 U1044 ( .A(G237), .ZN(n1251) );
XNOR2_X1 U1045 ( .A(n1313), .B(n1314), .ZN(n1309) );
NOR2_X1 U1046 ( .A1(KEYINPUT2), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1047 ( .A(G104), .B(n1316), .Z(n1315) );
XNOR2_X1 U1048 ( .A(G122), .B(n1233), .ZN(n1316) );
INV_X1 U1049 ( .A(G113), .ZN(n1233) );
NOR2_X1 U1050 ( .A1(KEYINPUT19), .A2(n1317), .ZN(n1313) );
NOR2_X1 U1051 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XOR2_X1 U1052 ( .A(KEYINPUT61), .B(n1320), .Z(n1319) );
NOR2_X1 U1053 ( .A1(n1321), .A2(n1089), .ZN(n1320) );
XNOR2_X1 U1054 ( .A(G125), .B(KEYINPUT30), .ZN(n1321) );
NOR2_X1 U1055 ( .A1(n1157), .A2(n1268), .ZN(n1318) );
INV_X1 U1056 ( .A(G125), .ZN(n1268) );
INV_X1 U1057 ( .A(n1089), .ZN(n1157) );
XOR2_X1 U1058 ( .A(G140), .B(KEYINPUT60), .Z(n1089) );
NAND2_X1 U1059 ( .A1(KEYINPUT1), .A2(n1123), .ZN(n1303) );
INV_X1 U1060 ( .A(G475), .ZN(n1123) );
XNOR2_X1 U1061 ( .A(n1322), .B(G478), .ZN(n1059) );
NAND2_X1 U1062 ( .A1(n1117), .A2(n1173), .ZN(n1322) );
INV_X1 U1063 ( .A(G902), .ZN(n1173) );
XOR2_X1 U1064 ( .A(n1323), .B(n1324), .Z(n1117) );
XOR2_X1 U1065 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1066 ( .A(G107), .B(n1327), .Z(n1326) );
NOR2_X1 U1067 ( .A1(n1328), .A2(n1270), .ZN(n1327) );
NAND2_X1 U1068 ( .A1(n1329), .A2(n1044), .ZN(n1270) );
INV_X1 U1069 ( .A(G953), .ZN(n1044) );
XNOR2_X1 U1070 ( .A(G234), .B(KEYINPUT36), .ZN(n1329) );
XNOR2_X1 U1071 ( .A(G217), .B(KEYINPUT49), .ZN(n1328) );
NOR2_X1 U1072 ( .A1(n1330), .A2(n1331), .ZN(n1325) );
XOR2_X1 U1073 ( .A(KEYINPUT8), .B(n1332), .Z(n1331) );
NOR2_X1 U1074 ( .A1(G143), .A2(n1333), .ZN(n1332) );
AND2_X1 U1075 ( .A1(n1333), .A2(G143), .ZN(n1330) );
INV_X1 U1076 ( .A(G128), .ZN(n1333) );
XNOR2_X1 U1077 ( .A(G116), .B(n1334), .ZN(n1323) );
XNOR2_X1 U1078 ( .A(n1217), .B(G122), .ZN(n1334) );
INV_X1 U1079 ( .A(G134), .ZN(n1217) );
endmodule


