//Key = 0010010010000100010001011111101100110010010100010111100000001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360;

XNOR2_X1 U743 ( .A(n1028), .B(n1029), .ZN(G9) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U745 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
XOR2_X1 U746 ( .A(n1036), .B(KEYINPUT2), .Z(n1034) );
NAND2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND3_X1 U749 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NAND2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1039) );
NAND3_X1 U751 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NAND2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND3_X1 U753 ( .A1(n1051), .A2(n1052), .A3(n1043), .ZN(n1047) );
NAND3_X1 U754 ( .A1(n1053), .A2(n1042), .A3(n1054), .ZN(n1046) );
NAND4_X1 U755 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1032) );
NAND4_X1 U756 ( .A1(n1043), .A2(n1059), .A3(n1060), .A4(n1044), .ZN(n1056) );
NOR2_X1 U757 ( .A1(n1061), .A2(n1051), .ZN(n1060) );
XNOR2_X1 U758 ( .A(n1037), .B(KEYINPUT56), .ZN(n1061) );
NAND3_X1 U759 ( .A1(n1042), .A2(n1062), .A3(n1037), .ZN(n1055) );
INV_X1 U760 ( .A(n1063), .ZN(n1037) );
NAND2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1044), .A2(n1066), .ZN(n1065) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U764 ( .A1(n1069), .A2(n1050), .A3(n1070), .ZN(n1068) );
NAND2_X1 U765 ( .A1(n1053), .A2(n1071), .ZN(n1067) );
NAND2_X1 U766 ( .A1(n1043), .A2(n1072), .ZN(n1064) );
AND2_X1 U767 ( .A1(n1053), .A2(n1050), .ZN(n1043) );
NOR3_X1 U768 ( .A1(n1073), .A2(G953), .A3(G952), .ZN(n1030) );
INV_X1 U769 ( .A(n1057), .ZN(n1073) );
NAND4_X1 U770 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1057) );
NOR4_X1 U771 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
XOR2_X1 U772 ( .A(n1082), .B(n1083), .Z(n1079) );
XNOR2_X1 U773 ( .A(G469), .B(KEYINPUT36), .ZN(n1083) );
NAND3_X1 U774 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1078) );
XOR2_X1 U775 ( .A(n1087), .B(KEYINPUT48), .Z(n1086) );
NAND2_X1 U776 ( .A1(KEYINPUT1), .A2(n1088), .ZN(n1085) );
OR3_X1 U777 ( .A1(n1089), .A2(KEYINPUT1), .A3(n1088), .ZN(n1084) );
NOR3_X1 U778 ( .A1(n1059), .A2(n1090), .A3(n1070), .ZN(n1076) );
XNOR2_X1 U779 ( .A(n1091), .B(n1092), .ZN(n1074) );
NOR2_X1 U780 ( .A1(n1093), .A2(KEYINPUT53), .ZN(n1092) );
INV_X1 U781 ( .A(n1094), .ZN(n1093) );
XOR2_X1 U782 ( .A(n1095), .B(n1096), .Z(G72) );
NOR2_X1 U783 ( .A1(n1058), .A2(n1097), .ZN(n1096) );
XOR2_X1 U784 ( .A(KEYINPUT29), .B(n1098), .Z(n1097) );
NOR2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1095) );
NAND2_X1 U787 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U788 ( .A(n1105), .B(n1106), .Z(n1101) );
NOR2_X1 U789 ( .A1(n1107), .A2(G953), .ZN(n1106) );
OR2_X1 U790 ( .A1(n1104), .A2(n1103), .ZN(n1105) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1103) );
NAND2_X1 U792 ( .A1(G953), .A2(n1100), .ZN(n1109) );
XOR2_X1 U793 ( .A(n1110), .B(n1111), .Z(n1108) );
XNOR2_X1 U794 ( .A(KEYINPUT39), .B(n1112), .ZN(n1111) );
XNOR2_X1 U795 ( .A(n1113), .B(n1114), .ZN(n1110) );
NOR2_X1 U796 ( .A1(G140), .A2(KEYINPUT44), .ZN(n1114) );
NOR2_X1 U797 ( .A1(KEYINPUT33), .A2(n1115), .ZN(n1113) );
XOR2_X1 U798 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND3_X1 U799 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1116) );
OR2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND3_X1 U801 ( .A1(n1122), .A2(n1121), .A3(G131), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1123), .A2(n1124), .ZN(n1118) );
NAND2_X1 U803 ( .A1(n1125), .A2(n1121), .ZN(n1123) );
INV_X1 U804 ( .A(KEYINPUT4), .ZN(n1121) );
XOR2_X1 U805 ( .A(KEYINPUT14), .B(n1122), .Z(n1125) );
INV_X1 U806 ( .A(KEYINPUT17), .ZN(n1104) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(G69) );
AND2_X1 U808 ( .A1(n1035), .A2(n1058), .ZN(n1127) );
NAND2_X1 U809 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NAND2_X1 U810 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
INV_X1 U811 ( .A(n1132), .ZN(n1130) );
NAND2_X1 U812 ( .A1(n1133), .A2(n1132), .ZN(n1128) );
NAND2_X1 U813 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
XOR2_X1 U814 ( .A(n1136), .B(KEYINPUT62), .Z(n1134) );
NAND2_X1 U815 ( .A1(n1135), .A2(n1131), .ZN(n1133) );
NAND2_X1 U816 ( .A1(G953), .A2(n1137), .ZN(n1131) );
INV_X1 U817 ( .A(n1138), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XNOR2_X1 U819 ( .A(n1141), .B(n1142), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U821 ( .A1(n1139), .A2(n1145), .ZN(G63) );
XOR2_X1 U822 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U823 ( .A(n1148), .B(KEYINPUT57), .Z(n1147) );
NAND3_X1 U824 ( .A1(G478), .A2(n1149), .A3(n1150), .ZN(n1146) );
XNOR2_X1 U825 ( .A(G902), .B(KEYINPUT13), .ZN(n1150) );
NOR2_X1 U826 ( .A1(n1139), .A2(n1151), .ZN(G60) );
XOR2_X1 U827 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND3_X1 U828 ( .A1(n1154), .A2(G475), .A3(KEYINPUT5), .ZN(n1152) );
XOR2_X1 U829 ( .A(G104), .B(n1155), .Z(G6) );
NOR2_X1 U830 ( .A1(n1139), .A2(n1156), .ZN(G57) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U832 ( .A1(n1088), .A2(n1144), .ZN(n1157) );
NOR2_X1 U833 ( .A1(n1139), .A2(n1159), .ZN(G54) );
XOR2_X1 U834 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U836 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
OR2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U838 ( .A(n1168), .B(KEYINPUT55), .Z(n1164) );
NAND2_X1 U839 ( .A1(n1167), .A2(n1166), .ZN(n1168) );
XOR2_X1 U840 ( .A(n1169), .B(n1117), .Z(n1166) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1160) );
NOR2_X1 U842 ( .A1(n1172), .A2(KEYINPUT22), .ZN(n1171) );
AND2_X1 U843 ( .A1(G469), .A2(n1154), .ZN(n1172) );
INV_X1 U844 ( .A(n1144), .ZN(n1154) );
NOR2_X1 U845 ( .A1(n1139), .A2(n1173), .ZN(G51) );
XOR2_X1 U846 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U847 ( .A(n1176), .B(n1136), .ZN(n1175) );
XOR2_X1 U848 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U849 ( .A1(KEYINPUT49), .A2(n1179), .ZN(n1177) );
XOR2_X1 U850 ( .A(n1180), .B(n1181), .Z(n1174) );
NOR2_X1 U851 ( .A1(n1094), .A2(n1144), .ZN(n1181) );
NAND2_X1 U852 ( .A1(G902), .A2(n1149), .ZN(n1144) );
NAND2_X1 U853 ( .A1(n1107), .A2(n1182), .ZN(n1149) );
XNOR2_X1 U854 ( .A(KEYINPUT3), .B(n1035), .ZN(n1182) );
NAND2_X1 U855 ( .A1(n1183), .A2(n1184), .ZN(n1035) );
NOR4_X1 U856 ( .A1(n1185), .A2(n1155), .A3(n1029), .A4(n1186), .ZN(n1184) );
NOR4_X1 U857 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1186) );
NOR2_X1 U858 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
INV_X1 U859 ( .A(KEYINPUT15), .ZN(n1192) );
NOR2_X1 U860 ( .A1(KEYINPUT15), .A2(n1193), .ZN(n1187) );
AND3_X1 U861 ( .A1(n1072), .A2(n1194), .A3(n1050), .ZN(n1029) );
AND3_X1 U862 ( .A1(n1050), .A2(n1194), .A3(n1041), .ZN(n1155) );
NOR4_X1 U863 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1183) );
AND3_X1 U864 ( .A1(n1044), .A2(n1194), .A3(n1071), .ZN(n1198) );
INV_X1 U865 ( .A(n1199), .ZN(n1194) );
INV_X1 U866 ( .A(n1200), .ZN(n1196) );
NOR3_X1 U867 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1195) );
NOR2_X1 U868 ( .A1(n1191), .A2(n1204), .ZN(n1203) );
INV_X1 U869 ( .A(KEYINPUT7), .ZN(n1204) );
NOR3_X1 U870 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1191) );
INV_X1 U871 ( .A(n1208), .ZN(n1207) );
INV_X1 U872 ( .A(n1042), .ZN(n1205) );
NOR2_X1 U873 ( .A1(KEYINPUT7), .A2(n1193), .ZN(n1202) );
INV_X1 U874 ( .A(n1033), .ZN(n1107) );
NAND2_X1 U875 ( .A1(n1209), .A2(n1210), .ZN(n1033) );
NOR4_X1 U876 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
AND4_X1 U877 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1209) );
OR3_X1 U878 ( .A1(n1201), .A2(n1219), .A3(n1220), .ZN(n1218) );
XNOR2_X1 U879 ( .A(n1053), .B(KEYINPUT9), .ZN(n1219) );
XNOR2_X1 U880 ( .A(G125), .B(KEYINPUT63), .ZN(n1180) );
NOR2_X1 U881 ( .A1(n1058), .A2(G952), .ZN(n1139) );
XNOR2_X1 U882 ( .A(G146), .B(n1217), .ZN(G48) );
NAND3_X1 U883 ( .A1(n1041), .A2(n1206), .A3(n1221), .ZN(n1217) );
XNOR2_X1 U884 ( .A(G143), .B(n1216), .ZN(G45) );
NAND4_X1 U885 ( .A1(n1080), .A2(n1222), .A3(n1206), .A4(n1223), .ZN(n1216) );
NOR2_X1 U886 ( .A1(n1220), .A2(n1190), .ZN(n1223) );
XNOR2_X1 U887 ( .A(G140), .B(n1215), .ZN(G42) );
NAND4_X1 U888 ( .A1(n1053), .A2(n1224), .A3(n1071), .A4(n1041), .ZN(n1215) );
XOR2_X1 U889 ( .A(G137), .B(n1214), .Z(G39) );
AND3_X1 U890 ( .A1(n1053), .A2(n1221), .A3(n1044), .ZN(n1214) );
XNOR2_X1 U891 ( .A(G134), .B(n1225), .ZN(G36) );
NAND4_X1 U892 ( .A1(KEYINPUT23), .A2(n1226), .A3(n1053), .A4(n1224), .ZN(n1225) );
NAND2_X1 U893 ( .A1(n1227), .A2(n1228), .ZN(G33) );
NAND2_X1 U894 ( .A1(n1213), .A2(n1124), .ZN(n1228) );
XOR2_X1 U895 ( .A(KEYINPUT8), .B(n1229), .Z(n1227) );
NOR2_X1 U896 ( .A1(n1213), .A2(n1124), .ZN(n1229) );
INV_X1 U897 ( .A(G131), .ZN(n1124) );
AND4_X1 U898 ( .A1(n1054), .A2(n1053), .A3(n1224), .A4(n1041), .ZN(n1213) );
NOR2_X1 U899 ( .A1(n1230), .A2(n1070), .ZN(n1053) );
XNOR2_X1 U900 ( .A(n1212), .B(n1231), .ZN(G30) );
XOR2_X1 U901 ( .A(KEYINPUT26), .B(G128), .Z(n1231) );
AND3_X1 U902 ( .A1(n1072), .A2(n1206), .A3(n1221), .ZN(n1212) );
AND3_X1 U903 ( .A1(n1232), .A2(n1233), .A3(n1224), .ZN(n1221) );
INV_X1 U904 ( .A(n1220), .ZN(n1224) );
NAND3_X1 U905 ( .A1(n1051), .A2(n1052), .A3(n1234), .ZN(n1220) );
NAND2_X1 U906 ( .A1(KEYINPUT40), .A2(n1190), .ZN(n1233) );
NAND2_X1 U907 ( .A1(n1235), .A2(n1236), .ZN(n1232) );
INV_X1 U908 ( .A(KEYINPUT40), .ZN(n1236) );
NAND2_X1 U909 ( .A1(n1081), .A2(n1237), .ZN(n1235) );
XOR2_X1 U910 ( .A(G101), .B(n1185), .Z(G3) );
NOR3_X1 U911 ( .A1(n1190), .A2(n1199), .A3(n1238), .ZN(n1185) );
XOR2_X1 U912 ( .A(n1239), .B(n1211), .Z(G27) );
AND4_X1 U913 ( .A1(n1071), .A2(n1049), .A3(n1041), .A4(n1234), .ZN(n1211) );
NAND2_X1 U914 ( .A1(n1063), .A2(n1240), .ZN(n1234) );
NAND4_X1 U915 ( .A1(G902), .A2(G953), .A3(n1241), .A4(n1100), .ZN(n1240) );
INV_X1 U916 ( .A(G900), .ZN(n1100) );
INV_X1 U917 ( .A(n1189), .ZN(n1041) );
NAND2_X1 U918 ( .A1(KEYINPUT24), .A2(n1112), .ZN(n1239) );
XOR2_X1 U919 ( .A(G122), .B(n1197), .Z(G24) );
AND4_X1 U920 ( .A1(n1193), .A2(n1050), .A3(n1080), .A4(n1222), .ZN(n1197) );
NOR2_X1 U921 ( .A1(n1237), .A2(n1081), .ZN(n1050) );
XNOR2_X1 U922 ( .A(G119), .B(n1200), .ZN(G21) );
NAND4_X1 U923 ( .A1(n1193), .A2(n1044), .A3(n1242), .A4(n1237), .ZN(n1200) );
XNOR2_X1 U924 ( .A(KEYINPUT40), .B(n1243), .ZN(n1242) );
XOR2_X1 U925 ( .A(n1244), .B(n1245), .Z(G18) );
XNOR2_X1 U926 ( .A(G116), .B(KEYINPUT45), .ZN(n1245) );
NAND2_X1 U927 ( .A1(n1193), .A2(n1226), .ZN(n1244) );
INV_X1 U928 ( .A(n1201), .ZN(n1226) );
NAND2_X1 U929 ( .A1(n1054), .A2(n1072), .ZN(n1201) );
NOR2_X1 U930 ( .A1(n1222), .A2(n1246), .ZN(n1072) );
INV_X1 U931 ( .A(n1190), .ZN(n1054) );
INV_X1 U932 ( .A(n1247), .ZN(n1193) );
XNOR2_X1 U933 ( .A(n1248), .B(n1249), .ZN(G15) );
NOR4_X1 U934 ( .A1(KEYINPUT11), .A2(n1189), .A3(n1190), .A4(n1247), .ZN(n1249) );
NAND2_X1 U935 ( .A1(n1049), .A2(n1208), .ZN(n1247) );
AND2_X1 U936 ( .A1(n1042), .A2(n1206), .ZN(n1049) );
NOR2_X1 U937 ( .A1(n1051), .A2(n1059), .ZN(n1042) );
INV_X1 U938 ( .A(n1052), .ZN(n1059) );
NAND2_X1 U939 ( .A1(n1243), .A2(n1237), .ZN(n1190) );
NAND2_X1 U940 ( .A1(n1246), .A2(n1222), .ZN(n1189) );
INV_X1 U941 ( .A(n1080), .ZN(n1246) );
XNOR2_X1 U942 ( .A(n1250), .B(n1251), .ZN(G12) );
NOR3_X1 U943 ( .A1(n1252), .A2(n1199), .A3(n1238), .ZN(n1251) );
INV_X1 U944 ( .A(n1044), .ZN(n1238) );
NOR2_X1 U945 ( .A1(n1080), .A2(n1222), .ZN(n1044) );
NAND2_X1 U946 ( .A1(n1087), .A2(n1075), .ZN(n1222) );
NAND2_X1 U947 ( .A1(G475), .A2(n1253), .ZN(n1075) );
OR2_X1 U948 ( .A1(n1253), .A2(G475), .ZN(n1087) );
NAND2_X1 U949 ( .A1(n1153), .A2(n1254), .ZN(n1253) );
XOR2_X1 U950 ( .A(n1255), .B(n1256), .Z(n1153) );
XOR2_X1 U951 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U952 ( .A(n1259), .B(n1260), .Z(n1258) );
NAND2_X1 U953 ( .A1(KEYINPUT25), .A2(n1261), .ZN(n1259) );
XNOR2_X1 U954 ( .A(n1262), .B(n1263), .ZN(n1257) );
NOR2_X1 U955 ( .A1(KEYINPUT37), .A2(n1248), .ZN(n1263) );
INV_X1 U956 ( .A(G113), .ZN(n1248) );
NOR4_X1 U957 ( .A1(KEYINPUT10), .A2(G953), .A3(G237), .A4(n1264), .ZN(n1262) );
INV_X1 U958 ( .A(G214), .ZN(n1264) );
XOR2_X1 U959 ( .A(n1265), .B(n1266), .Z(n1255) );
XOR2_X1 U960 ( .A(G122), .B(G104), .Z(n1266) );
XNOR2_X1 U961 ( .A(G143), .B(G131), .ZN(n1265) );
XOR2_X1 U962 ( .A(G478), .B(n1267), .Z(n1080) );
NOR2_X1 U963 ( .A1(G902), .A2(n1268), .ZN(n1267) );
XOR2_X1 U964 ( .A(n1148), .B(KEYINPUT51), .Z(n1268) );
NAND3_X1 U965 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1148) );
NAND2_X1 U966 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND3_X1 U967 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
NAND2_X1 U968 ( .A1(KEYINPUT38), .A2(n1277), .ZN(n1276) );
NAND2_X1 U969 ( .A1(KEYINPUT35), .A2(n1278), .ZN(n1275) );
NAND2_X1 U970 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U971 ( .A1(KEYINPUT30), .A2(n1281), .ZN(n1280) );
NAND2_X1 U972 ( .A1(n1279), .A2(n1282), .ZN(n1274) );
INV_X1 U973 ( .A(KEYINPUT35), .ZN(n1282) );
INV_X1 U974 ( .A(n1283), .ZN(n1272) );
NAND4_X1 U975 ( .A1(n1279), .A2(n1283), .A3(KEYINPUT38), .A4(KEYINPUT30), .ZN(n1270) );
NAND2_X1 U976 ( .A1(n1284), .A2(n1277), .ZN(n1269) );
INV_X1 U977 ( .A(KEYINPUT30), .ZN(n1277) );
NAND2_X1 U978 ( .A1(n1279), .A2(n1285), .ZN(n1284) );
NAND2_X1 U979 ( .A1(n1283), .A2(n1281), .ZN(n1285) );
INV_X1 U980 ( .A(KEYINPUT38), .ZN(n1281) );
NAND3_X1 U981 ( .A1(G234), .A2(n1058), .A3(G217), .ZN(n1283) );
XNOR2_X1 U982 ( .A(n1286), .B(n1287), .ZN(n1279) );
XOR2_X1 U983 ( .A(KEYINPUT21), .B(G134), .Z(n1287) );
XNOR2_X1 U984 ( .A(n1288), .B(n1289), .ZN(n1286) );
NOR2_X1 U985 ( .A1(KEYINPUT12), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U986 ( .A(n1028), .B(n1291), .ZN(n1290) );
XOR2_X1 U987 ( .A(G122), .B(G116), .Z(n1291) );
INV_X1 U988 ( .A(G107), .ZN(n1028) );
NAND4_X1 U989 ( .A1(n1206), .A2(n1051), .A3(n1208), .A4(n1052), .ZN(n1199) );
NAND2_X1 U990 ( .A1(G221), .A2(n1292), .ZN(n1052) );
NAND2_X1 U991 ( .A1(n1063), .A2(n1293), .ZN(n1208) );
NAND3_X1 U992 ( .A1(n1138), .A2(n1241), .A3(G902), .ZN(n1293) );
NOR2_X1 U993 ( .A1(G898), .A2(n1058), .ZN(n1138) );
NAND3_X1 U994 ( .A1(n1241), .A2(n1058), .A3(n1294), .ZN(n1063) );
XNOR2_X1 U995 ( .A(G952), .B(KEYINPUT41), .ZN(n1294) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1241) );
NAND2_X1 U997 ( .A1(n1295), .A2(n1296), .ZN(n1051) );
NAND2_X1 U998 ( .A1(G469), .A2(n1082), .ZN(n1296) );
XOR2_X1 U999 ( .A(KEYINPUT61), .B(n1297), .Z(n1295) );
NOR2_X1 U1000 ( .A1(G469), .A2(n1082), .ZN(n1297) );
NAND2_X1 U1001 ( .A1(n1298), .A2(n1254), .ZN(n1082) );
XOR2_X1 U1002 ( .A(n1299), .B(n1300), .Z(n1298) );
XOR2_X1 U1003 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1004 ( .A(n1117), .B(n1167), .Z(n1302) );
XOR2_X1 U1005 ( .A(n1178), .B(KEYINPUT60), .Z(n1117) );
NAND2_X1 U1006 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
NAND2_X1 U1007 ( .A1(KEYINPUT43), .A2(n1163), .ZN(n1304) );
XNOR2_X1 U1008 ( .A(G140), .B(G110), .ZN(n1163) );
NAND3_X1 U1009 ( .A1(G140), .A2(n1250), .A3(n1305), .ZN(n1303) );
INV_X1 U1010 ( .A(KEYINPUT43), .ZN(n1305) );
XNOR2_X1 U1011 ( .A(n1170), .B(n1306), .ZN(n1299) );
XNOR2_X1 U1012 ( .A(KEYINPUT54), .B(n1307), .ZN(n1306) );
NOR2_X1 U1013 ( .A1(KEYINPUT6), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U1014 ( .A(KEYINPUT59), .B(n1309), .ZN(n1308) );
INV_X1 U1015 ( .A(n1169), .ZN(n1309) );
XNOR2_X1 U1016 ( .A(n1310), .B(n1311), .ZN(n1169) );
XOR2_X1 U1017 ( .A(G101), .B(n1312), .Z(n1311) );
NOR2_X1 U1018 ( .A1(G104), .A2(KEYINPUT19), .ZN(n1312) );
XNOR2_X1 U1019 ( .A(G107), .B(KEYINPUT31), .ZN(n1310) );
NOR2_X1 U1020 ( .A1(n1099), .A2(G953), .ZN(n1170) );
INV_X1 U1021 ( .A(G227), .ZN(n1099) );
NOR2_X1 U1022 ( .A1(n1069), .A2(n1070), .ZN(n1206) );
AND2_X1 U1023 ( .A1(G214), .A2(n1313), .ZN(n1070) );
INV_X1 U1024 ( .A(n1230), .ZN(n1069) );
XOR2_X1 U1025 ( .A(n1091), .B(n1094), .Z(n1230) );
NAND2_X1 U1026 ( .A1(G210), .A2(n1313), .ZN(n1094) );
NAND2_X1 U1027 ( .A1(n1314), .A2(n1254), .ZN(n1313) );
XNOR2_X1 U1028 ( .A(G237), .B(KEYINPUT0), .ZN(n1314) );
NAND3_X1 U1029 ( .A1(n1315), .A2(n1316), .A3(n1254), .ZN(n1091) );
NAND2_X1 U1030 ( .A1(n1317), .A2(n1136), .ZN(n1316) );
NAND2_X1 U1031 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND2_X1 U1032 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
INV_X1 U1033 ( .A(KEYINPUT46), .ZN(n1321) );
NAND2_X1 U1034 ( .A1(KEYINPUT46), .A2(n1322), .ZN(n1318) );
OR2_X1 U1035 ( .A1(n1136), .A2(n1320), .ZN(n1315) );
NAND2_X1 U1036 ( .A1(KEYINPUT34), .A2(n1322), .ZN(n1320) );
XOR2_X1 U1037 ( .A(n1323), .B(n1324), .Z(n1322) );
XNOR2_X1 U1038 ( .A(G125), .B(n1325), .ZN(n1324) );
NAND2_X1 U1039 ( .A1(KEYINPUT47), .A2(n1178), .ZN(n1325) );
NAND2_X1 U1040 ( .A1(KEYINPUT50), .A2(n1179), .ZN(n1323) );
NOR2_X1 U1041 ( .A1(n1137), .A2(G953), .ZN(n1179) );
INV_X1 U1042 ( .A(G224), .ZN(n1137) );
XOR2_X1 U1043 ( .A(n1326), .B(n1327), .Z(n1136) );
XOR2_X1 U1044 ( .A(n1328), .B(n1329), .Z(n1327) );
NAND2_X1 U1045 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1046 ( .A1(G122), .A2(n1250), .ZN(n1331) );
XOR2_X1 U1047 ( .A(n1332), .B(KEYINPUT18), .Z(n1330) );
OR2_X1 U1048 ( .A1(n1250), .A2(G122), .ZN(n1332) );
NAND2_X1 U1049 ( .A1(n1333), .A2(n1334), .ZN(n1328) );
NAND2_X1 U1050 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
XOR2_X1 U1051 ( .A(n1337), .B(KEYINPUT58), .Z(n1333) );
OR2_X1 U1052 ( .A1(n1336), .A2(n1335), .ZN(n1337) );
XOR2_X1 U1053 ( .A(n1338), .B(KEYINPUT16), .Z(n1336) );
XNOR2_X1 U1054 ( .A(G101), .B(n1339), .ZN(n1326) );
NOR2_X1 U1055 ( .A1(KEYINPUT32), .A2(n1340), .ZN(n1339) );
XNOR2_X1 U1056 ( .A(G104), .B(G107), .ZN(n1340) );
XOR2_X1 U1057 ( .A(KEYINPUT27), .B(n1071), .Z(n1252) );
NOR2_X1 U1058 ( .A1(n1237), .A2(n1243), .ZN(n1071) );
INV_X1 U1059 ( .A(n1081), .ZN(n1243) );
XOR2_X1 U1060 ( .A(n1341), .B(n1143), .Z(n1081) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1292), .ZN(n1143) );
NAND2_X1 U1062 ( .A1(G234), .A2(n1254), .ZN(n1292) );
NAND2_X1 U1063 ( .A1(n1141), .A2(n1254), .ZN(n1341) );
INV_X1 U1064 ( .A(G902), .ZN(n1254) );
XNOR2_X1 U1065 ( .A(n1342), .B(n1343), .ZN(n1141) );
XOR2_X1 U1066 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1067 ( .A(n1261), .B(G110), .ZN(n1345) );
INV_X1 U1068 ( .A(G146), .ZN(n1261) );
NOR3_X1 U1069 ( .A1(n1346), .A2(KEYINPUT42), .A3(n1347), .ZN(n1344) );
NOR2_X1 U1070 ( .A1(n1348), .A2(G137), .ZN(n1347) );
AND3_X1 U1071 ( .A1(G221), .A2(n1058), .A3(G234), .ZN(n1348) );
XOR2_X1 U1072 ( .A(KEYINPUT20), .B(n1349), .Z(n1346) );
AND4_X1 U1073 ( .A1(n1058), .A2(G137), .A3(G234), .A4(G221), .ZN(n1349) );
INV_X1 U1074 ( .A(G953), .ZN(n1058) );
XOR2_X1 U1075 ( .A(n1350), .B(n1260), .Z(n1342) );
XNOR2_X1 U1076 ( .A(n1112), .B(G140), .ZN(n1260) );
INV_X1 U1077 ( .A(G125), .ZN(n1112) );
NAND2_X1 U1078 ( .A1(KEYINPUT52), .A2(n1351), .ZN(n1350) );
XNOR2_X1 U1079 ( .A(G128), .B(n1352), .ZN(n1351) );
INV_X1 U1080 ( .A(G119), .ZN(n1352) );
OR2_X1 U1081 ( .A1(n1353), .A2(n1090), .ZN(n1237) );
AND2_X1 U1082 ( .A1(n1089), .A2(n1088), .ZN(n1090) );
NOR2_X1 U1083 ( .A1(n1088), .A2(n1089), .ZN(n1353) );
NOR2_X1 U1084 ( .A1(n1158), .A2(G902), .ZN(n1089) );
XNOR2_X1 U1085 ( .A(n1354), .B(n1355), .ZN(n1158) );
XNOR2_X1 U1086 ( .A(n1167), .B(n1356), .ZN(n1355) );
XOR2_X1 U1087 ( .A(G101), .B(n1357), .Z(n1356) );
NOR3_X1 U1088 ( .A1(n1358), .A2(G953), .A3(G237), .ZN(n1357) );
INV_X1 U1089 ( .A(G210), .ZN(n1358) );
XNOR2_X1 U1090 ( .A(G131), .B(n1122), .ZN(n1167) );
XOR2_X1 U1091 ( .A(G134), .B(G137), .Z(n1122) );
XNOR2_X1 U1092 ( .A(n1359), .B(n1335), .ZN(n1354) );
XNOR2_X1 U1093 ( .A(G116), .B(G119), .ZN(n1335) );
XNOR2_X1 U1094 ( .A(n1178), .B(n1338), .ZN(n1359) );
XOR2_X1 U1095 ( .A(G113), .B(KEYINPUT28), .Z(n1338) );
XOR2_X1 U1096 ( .A(G146), .B(n1288), .Z(n1178) );
XNOR2_X1 U1097 ( .A(G128), .B(n1360), .ZN(n1288) );
INV_X1 U1098 ( .A(G143), .ZN(n1360) );
INV_X1 U1099 ( .A(G472), .ZN(n1088) );
INV_X1 U1100 ( .A(G110), .ZN(n1250) );
endmodule


