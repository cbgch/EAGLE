//Key = 1010100011111101100101011010110000111110010001011000001010011111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366;

XNOR2_X1 U756 ( .A(n1054), .B(n1055), .ZN(G9) );
NAND2_X1 U757 ( .A1(KEYINPUT54), .A2(n1056), .ZN(n1054) );
NOR2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(G75) );
NOR3_X1 U759 ( .A1(n1059), .A2(G953), .A3(G952), .ZN(n1058) );
NOR4_X1 U760 ( .A1(G953), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1057) );
NOR2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U764 ( .A(n1068), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U769 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(n1073) );
NOR2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR3_X1 U773 ( .A1(n1082), .A2(n1085), .A3(n1076), .ZN(n1069) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR4_X1 U776 ( .A1(n1090), .A2(n1076), .A3(n1072), .A4(n1082), .ZN(n1064) );
NOR2_X1 U777 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
AND4_X1 U778 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1059) );
NOR4_X1 U779 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XOR2_X1 U780 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U781 ( .A1(G475), .A2(KEYINPUT31), .ZN(n1102) );
XOR2_X1 U782 ( .A(n1103), .B(KEYINPUT17), .Z(n1101) );
XOR2_X1 U783 ( .A(n1104), .B(KEYINPUT26), .Z(n1099) );
INV_X1 U784 ( .A(n1105), .ZN(n1098) );
NOR2_X1 U785 ( .A1(n1072), .A2(n1106), .ZN(n1095) );
XNOR2_X1 U786 ( .A(KEYINPUT3), .B(n1107), .ZN(n1106) );
XNOR2_X1 U787 ( .A(G472), .B(n1108), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U789 ( .A(KEYINPUT41), .B(KEYINPUT16), .ZN(n1109) );
XOR2_X1 U790 ( .A(n1111), .B(n1112), .Z(G72) );
NOR2_X1 U791 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR3_X1 U792 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NOR2_X1 U793 ( .A1(G953), .A2(n1118), .ZN(n1113) );
XNOR2_X1 U794 ( .A(n1119), .B(n1116), .ZN(n1118) );
XNOR2_X1 U795 ( .A(n1120), .B(n1121), .ZN(n1116) );
XOR2_X1 U796 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U797 ( .A(G131), .B(G140), .ZN(n1123) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NAND2_X1 U799 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U800 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NAND2_X1 U801 ( .A1(KEYINPUT51), .A2(KEYINPUT4), .ZN(n1129) );
NAND3_X1 U802 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1124) );
INV_X1 U803 ( .A(KEYINPUT51), .ZN(n1132) );
OR2_X1 U804 ( .A1(G137), .A2(KEYINPUT4), .ZN(n1131) );
NAND2_X1 U805 ( .A1(KEYINPUT4), .A2(n1133), .ZN(n1130) );
NAND2_X1 U806 ( .A1(G134), .A2(n1128), .ZN(n1133) );
XNOR2_X1 U807 ( .A(n1134), .B(n1135), .ZN(n1120) );
NOR2_X1 U808 ( .A1(G125), .A2(KEYINPUT57), .ZN(n1135) );
NOR2_X1 U809 ( .A1(KEYINPUT50), .A2(n1136), .ZN(n1134) );
NAND3_X1 U810 ( .A1(G953), .A2(n1137), .A3(KEYINPUT35), .ZN(n1111) );
NAND2_X1 U811 ( .A1(G900), .A2(G227), .ZN(n1137) );
XOR2_X1 U812 ( .A(n1138), .B(n1139), .Z(G69) );
NOR2_X1 U813 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U814 ( .A(n1142), .B(KEYINPUT24), .Z(n1141) );
NAND3_X1 U815 ( .A1(n1143), .A2(n1115), .A3(n1144), .ZN(n1142) );
NOR3_X1 U816 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1140) );
AND2_X1 U817 ( .A1(n1115), .A2(n1143), .ZN(n1146) );
NAND2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
XOR2_X1 U819 ( .A(n1055), .B(KEYINPUT25), .Z(n1147) );
NOR2_X1 U820 ( .A1(G898), .A2(n1115), .ZN(n1145) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(n1144) );
XNOR2_X1 U822 ( .A(n1151), .B(n1152), .ZN(n1149) );
NAND2_X1 U823 ( .A1(G953), .A2(n1153), .ZN(n1138) );
NAND2_X1 U824 ( .A1(G898), .A2(G224), .ZN(n1153) );
NOR2_X1 U825 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U826 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U828 ( .A1(n1154), .A2(n1160), .ZN(G63) );
XOR2_X1 U829 ( .A(n1161), .B(n1162), .Z(n1160) );
AND2_X1 U830 ( .A1(G478), .A2(n1158), .ZN(n1162) );
NAND2_X1 U831 ( .A1(KEYINPUT61), .A2(n1163), .ZN(n1161) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1164), .ZN(G60) );
XOR2_X1 U833 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U834 ( .A(n1167), .B(KEYINPUT46), .Z(n1165) );
NAND2_X1 U835 ( .A1(n1158), .A2(G475), .ZN(n1167) );
XNOR2_X1 U836 ( .A(G104), .B(n1168), .ZN(G6) );
NOR2_X1 U837 ( .A1(n1154), .A2(n1169), .ZN(G57) );
XOR2_X1 U838 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U839 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U840 ( .A1(G101), .A2(KEYINPUT20), .ZN(n1172) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1170) );
XOR2_X1 U842 ( .A(n1176), .B(KEYINPUT55), .Z(n1175) );
NAND2_X1 U843 ( .A1(n1158), .A2(G472), .ZN(n1174) );
NOR2_X1 U844 ( .A1(n1154), .A2(n1177), .ZN(G54) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U847 ( .A1(n1182), .A2(KEYINPUT6), .ZN(n1181) );
AND2_X1 U848 ( .A1(G469), .A2(n1158), .ZN(n1182) );
XOR2_X1 U849 ( .A(n1183), .B(n1184), .Z(n1178) );
NOR2_X1 U850 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U851 ( .A(n1187), .B(KEYINPUT19), .Z(n1186) );
NAND2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XNOR2_X1 U853 ( .A(n1190), .B(KEYINPUT43), .ZN(n1188) );
NOR2_X1 U854 ( .A1(n1191), .A2(n1189), .ZN(n1185) );
XOR2_X1 U855 ( .A(n1136), .B(n1192), .Z(n1189) );
NAND2_X1 U856 ( .A1(KEYINPUT9), .A2(n1193), .ZN(n1192) );
NAND2_X1 U857 ( .A1(n1194), .A2(n1195), .ZN(n1183) );
NAND2_X1 U858 ( .A1(G110), .A2(n1196), .ZN(n1195) );
XOR2_X1 U859 ( .A(n1197), .B(KEYINPUT58), .Z(n1194) );
OR2_X1 U860 ( .A1(n1196), .A2(G110), .ZN(n1197) );
XOR2_X1 U861 ( .A(G140), .B(KEYINPUT38), .Z(n1196) );
NOR2_X1 U862 ( .A1(n1154), .A2(n1198), .ZN(G51) );
XOR2_X1 U863 ( .A(n1199), .B(n1200), .Z(n1198) );
XNOR2_X1 U864 ( .A(n1201), .B(n1202), .ZN(n1200) );
XOR2_X1 U865 ( .A(n1203), .B(KEYINPUT28), .Z(n1199) );
NAND2_X1 U866 ( .A1(n1158), .A2(n1204), .ZN(n1203) );
AND2_X1 U867 ( .A1(n1205), .A2(n1061), .ZN(n1158) );
NAND3_X1 U868 ( .A1(n1148), .A2(n1055), .A3(n1119), .ZN(n1061) );
AND4_X1 U869 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1119) );
AND4_X1 U870 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
NAND2_X1 U871 ( .A1(n1078), .A2(n1214), .ZN(n1208) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND4_X1 U873 ( .A1(n1084), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1216) );
XNOR2_X1 U874 ( .A(KEYINPUT21), .B(n1220), .ZN(n1215) );
NAND3_X1 U875 ( .A1(n1091), .A2(n1221), .A3(n1222), .ZN(n1055) );
AND4_X1 U876 ( .A1(n1168), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1148) );
AND4_X1 U877 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
NAND2_X1 U878 ( .A1(n1230), .A2(n1231), .ZN(n1224) );
NAND3_X1 U879 ( .A1(n1222), .A2(n1221), .A3(n1092), .ZN(n1168) );
XNOR2_X1 U880 ( .A(G902), .B(KEYINPUT47), .ZN(n1205) );
AND2_X1 U881 ( .A1(n1232), .A2(G953), .ZN(n1154) );
XNOR2_X1 U882 ( .A(G952), .B(KEYINPUT18), .ZN(n1232) );
XNOR2_X1 U883 ( .A(G146), .B(n1207), .ZN(G48) );
NAND2_X1 U884 ( .A1(n1233), .A2(n1234), .ZN(n1207) );
NAND2_X1 U885 ( .A1(n1235), .A2(n1236), .ZN(G45) );
NAND2_X1 U886 ( .A1(G143), .A2(n1237), .ZN(n1236) );
XOR2_X1 U887 ( .A(KEYINPUT36), .B(n1238), .Z(n1235) );
NOR2_X1 U888 ( .A1(G143), .A2(n1237), .ZN(n1238) );
NAND4_X1 U889 ( .A1(n1084), .A2(n1078), .A3(n1239), .A4(n1240), .ZN(n1237) );
NOR3_X1 U890 ( .A1(n1241), .A2(n1242), .A3(n1093), .ZN(n1240) );
XNOR2_X1 U891 ( .A(n1087), .B(KEYINPUT0), .ZN(n1239) );
XNOR2_X1 U892 ( .A(G140), .B(n1213), .ZN(G42) );
NAND3_X1 U893 ( .A1(n1233), .A2(n1243), .A3(n1083), .ZN(n1213) );
XOR2_X1 U894 ( .A(n1212), .B(n1244), .Z(G39) );
NAND2_X1 U895 ( .A1(KEYINPUT63), .A2(G137), .ZN(n1244) );
NAND3_X1 U896 ( .A1(n1217), .A2(n1068), .A3(n1245), .ZN(n1212) );
NOR3_X1 U897 ( .A1(n1082), .A2(n1246), .A3(n1247), .ZN(n1245) );
XNOR2_X1 U898 ( .A(n1127), .B(n1248), .ZN(G36) );
NOR3_X1 U899 ( .A1(KEYINPUT27), .A2(n1249), .A3(n1250), .ZN(n1248) );
NOR2_X1 U900 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NOR2_X1 U901 ( .A1(n1253), .A2(n1082), .ZN(n1251) );
INV_X1 U902 ( .A(n1243), .ZN(n1082) );
AND2_X1 U903 ( .A1(n1252), .A2(n1206), .ZN(n1249) );
NAND2_X1 U904 ( .A1(n1253), .A2(n1243), .ZN(n1206) );
AND3_X1 U905 ( .A1(n1217), .A2(n1091), .A3(n1084), .ZN(n1253) );
INV_X1 U906 ( .A(KEYINPUT5), .ZN(n1252) );
XNOR2_X1 U907 ( .A(G131), .B(n1211), .ZN(G33) );
NAND3_X1 U908 ( .A1(n1233), .A2(n1243), .A3(n1084), .ZN(n1211) );
NOR2_X1 U909 ( .A1(n1079), .A2(n1097), .ZN(n1243) );
INV_X1 U910 ( .A(n1080), .ZN(n1097) );
AND2_X1 U911 ( .A1(n1092), .A2(n1217), .ZN(n1233) );
NOR2_X1 U912 ( .A1(n1254), .A2(n1242), .ZN(n1217) );
INV_X1 U913 ( .A(n1255), .ZN(n1242) );
INV_X1 U914 ( .A(n1087), .ZN(n1254) );
XOR2_X1 U915 ( .A(n1256), .B(KEYINPUT30), .Z(n1087) );
XNOR2_X1 U916 ( .A(G128), .B(n1210), .ZN(G30) );
NAND4_X1 U917 ( .A1(n1234), .A2(n1091), .A3(n1256), .A4(n1255), .ZN(n1210) );
XNOR2_X1 U918 ( .A(G101), .B(n1223), .ZN(G3) );
NAND3_X1 U919 ( .A1(n1068), .A2(n1222), .A3(n1084), .ZN(n1223) );
XOR2_X1 U920 ( .A(G125), .B(n1257), .Z(G27) );
NOR2_X1 U921 ( .A1(n1258), .A2(n1220), .ZN(n1257) );
NAND4_X1 U922 ( .A1(n1083), .A2(n1092), .A3(n1259), .A4(n1255), .ZN(n1220) );
NAND2_X1 U923 ( .A1(n1063), .A2(n1260), .ZN(n1255) );
NAND4_X1 U924 ( .A1(G953), .A2(G902), .A3(n1261), .A4(n1117), .ZN(n1260) );
INV_X1 U925 ( .A(G900), .ZN(n1117) );
XNOR2_X1 U926 ( .A(G122), .B(n1229), .ZN(G24) );
NAND4_X1 U927 ( .A1(n1262), .A2(n1221), .A3(n1218), .A4(n1219), .ZN(n1229) );
INV_X1 U928 ( .A(n1076), .ZN(n1221) );
NAND2_X1 U929 ( .A1(n1246), .A2(n1247), .ZN(n1076) );
XNOR2_X1 U930 ( .A(G119), .B(n1228), .ZN(G21) );
NAND4_X1 U931 ( .A1(n1234), .A2(n1068), .A3(n1259), .A4(n1263), .ZN(n1228) );
NOR3_X1 U932 ( .A1(n1247), .A2(n1246), .A3(n1258), .ZN(n1234) );
INV_X1 U933 ( .A(n1264), .ZN(n1246) );
XNOR2_X1 U934 ( .A(G116), .B(n1227), .ZN(G18) );
NAND3_X1 U935 ( .A1(n1084), .A2(n1091), .A3(n1262), .ZN(n1227) );
AND3_X1 U936 ( .A1(n1078), .A2(n1263), .A3(n1259), .ZN(n1262) );
NOR2_X1 U937 ( .A1(n1218), .A2(n1093), .ZN(n1091) );
INV_X1 U938 ( .A(n1219), .ZN(n1093) );
XNOR2_X1 U939 ( .A(G113), .B(n1265), .ZN(G15) );
NAND2_X1 U940 ( .A1(n1266), .A2(n1231), .ZN(n1265) );
XNOR2_X1 U941 ( .A(n1230), .B(KEYINPUT8), .ZN(n1266) );
AND4_X1 U942 ( .A1(n1084), .A2(n1092), .A3(n1259), .A4(n1263), .ZN(n1230) );
INV_X1 U943 ( .A(n1072), .ZN(n1259) );
NAND2_X1 U944 ( .A1(n1267), .A2(n1089), .ZN(n1072) );
INV_X1 U945 ( .A(n1088), .ZN(n1267) );
NOR2_X1 U946 ( .A1(n1219), .A2(n1241), .ZN(n1092) );
INV_X1 U947 ( .A(n1218), .ZN(n1241) );
NOR2_X1 U948 ( .A1(n1264), .A2(n1247), .ZN(n1084) );
XNOR2_X1 U949 ( .A(G110), .B(n1226), .ZN(G12) );
NAND3_X1 U950 ( .A1(n1068), .A2(n1222), .A3(n1083), .ZN(n1226) );
AND2_X1 U951 ( .A1(n1247), .A2(n1264), .ZN(n1083) );
NAND2_X1 U952 ( .A1(n1107), .A2(n1105), .ZN(n1264) );
NAND3_X1 U953 ( .A1(n1156), .A2(n1268), .A3(n1269), .ZN(n1105) );
NAND2_X1 U954 ( .A1(n1159), .A2(n1270), .ZN(n1107) );
NAND2_X1 U955 ( .A1(n1269), .A2(n1156), .ZN(n1270) );
NAND2_X1 U956 ( .A1(n1271), .A2(n1272), .ZN(n1156) );
NAND2_X1 U957 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U958 ( .A(KEYINPUT12), .B(n1275), .Z(n1271) );
NOR2_X1 U959 ( .A1(n1273), .A2(n1274), .ZN(n1275) );
XNOR2_X1 U960 ( .A(n1276), .B(n1277), .ZN(n1274) );
NOR2_X1 U961 ( .A1(KEYINPUT14), .A2(G137), .ZN(n1277) );
NAND2_X1 U962 ( .A1(n1278), .A2(G221), .ZN(n1276) );
NAND2_X1 U963 ( .A1(n1279), .A2(n1280), .ZN(n1273) );
NAND2_X1 U964 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XNOR2_X1 U965 ( .A(n1283), .B(KEYINPUT29), .ZN(n1281) );
NAND2_X1 U966 ( .A1(n1284), .A2(G140), .ZN(n1279) );
XNOR2_X1 U967 ( .A(KEYINPUT11), .B(n1285), .ZN(n1284) );
INV_X1 U968 ( .A(n1283), .ZN(n1285) );
XNOR2_X1 U969 ( .A(n1286), .B(n1287), .ZN(n1283) );
XNOR2_X1 U970 ( .A(n1288), .B(G125), .ZN(n1287) );
NAND2_X1 U971 ( .A1(n1289), .A2(KEYINPUT48), .ZN(n1286) );
XOR2_X1 U972 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U973 ( .A(KEYINPUT13), .B(n1292), .ZN(n1291) );
XNOR2_X1 U974 ( .A(G119), .B(G110), .ZN(n1290) );
XNOR2_X1 U975 ( .A(KEYINPUT15), .B(n1293), .ZN(n1269) );
INV_X1 U976 ( .A(n1268), .ZN(n1159) );
NAND2_X1 U977 ( .A1(G217), .A2(n1294), .ZN(n1268) );
XOR2_X1 U978 ( .A(n1110), .B(G472), .Z(n1247) );
NAND2_X1 U979 ( .A1(n1295), .A2(n1293), .ZN(n1110) );
XOR2_X1 U980 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U981 ( .A(n1173), .B(n1176), .Z(n1297) );
NAND3_X1 U982 ( .A1(n1298), .A2(n1115), .A3(G210), .ZN(n1176) );
XNOR2_X1 U983 ( .A(n1299), .B(n1300), .ZN(n1173) );
XNOR2_X1 U984 ( .A(n1301), .B(n1302), .ZN(n1300) );
XNOR2_X1 U985 ( .A(KEYINPUT49), .B(n1303), .ZN(n1302) );
INV_X1 U986 ( .A(n1304), .ZN(n1301) );
XNOR2_X1 U987 ( .A(n1190), .B(n1305), .ZN(n1299) );
XNOR2_X1 U988 ( .A(G101), .B(KEYINPUT53), .ZN(n1296) );
AND3_X1 U989 ( .A1(n1231), .A2(n1263), .A3(n1256), .ZN(n1222) );
AND2_X1 U990 ( .A1(n1088), .A2(n1089), .ZN(n1256) );
NAND2_X1 U991 ( .A1(G221), .A2(n1294), .ZN(n1089) );
NAND2_X1 U992 ( .A1(G234), .A2(n1293), .ZN(n1294) );
XNOR2_X1 U993 ( .A(n1306), .B(G469), .ZN(n1088) );
NAND2_X1 U994 ( .A1(n1307), .A2(n1293), .ZN(n1306) );
XOR2_X1 U995 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U996 ( .A(n1310), .B(n1180), .Z(n1309) );
AND2_X1 U997 ( .A1(G227), .A2(n1115), .ZN(n1180) );
NAND2_X1 U998 ( .A1(n1311), .A2(KEYINPUT10), .ZN(n1310) );
XOR2_X1 U999 ( .A(n1312), .B(n1193), .Z(n1311) );
XNOR2_X1 U1000 ( .A(n1313), .B(n1314), .ZN(n1193) );
NOR2_X1 U1001 ( .A1(KEYINPUT44), .A2(n1315), .ZN(n1314) );
XOR2_X1 U1002 ( .A(n1316), .B(n1317), .Z(n1315) );
XOR2_X1 U1003 ( .A(KEYINPUT1), .B(G104), .Z(n1317) );
NAND2_X1 U1004 ( .A1(KEYINPUT37), .A2(n1056), .ZN(n1316) );
XNOR2_X1 U1005 ( .A(n1318), .B(n1191), .ZN(n1312) );
INV_X1 U1006 ( .A(n1190), .ZN(n1191) );
XOR2_X1 U1007 ( .A(G131), .B(n1319), .Z(n1190) );
XNOR2_X1 U1008 ( .A(n1128), .B(G134), .ZN(n1319) );
INV_X1 U1009 ( .A(G137), .ZN(n1128) );
NAND2_X1 U1010 ( .A1(KEYINPUT60), .A2(n1320), .ZN(n1318) );
XNOR2_X1 U1011 ( .A(KEYINPUT7), .B(n1136), .ZN(n1320) );
NAND2_X1 U1012 ( .A1(n1321), .A2(n1322), .ZN(n1136) );
OR2_X1 U1013 ( .A1(n1292), .A2(n1323), .ZN(n1322) );
XOR2_X1 U1014 ( .A(n1324), .B(KEYINPUT42), .Z(n1321) );
NAND2_X1 U1015 ( .A1(n1323), .A2(n1292), .ZN(n1324) );
XNOR2_X1 U1016 ( .A(n1325), .B(G143), .ZN(n1323) );
NAND2_X1 U1017 ( .A1(KEYINPUT62), .A2(n1288), .ZN(n1325) );
INV_X1 U1018 ( .A(G146), .ZN(n1288) );
XNOR2_X1 U1019 ( .A(G110), .B(G140), .ZN(n1308) );
NAND2_X1 U1020 ( .A1(n1326), .A2(n1063), .ZN(n1263) );
NAND3_X1 U1021 ( .A1(n1261), .A2(n1115), .A3(G952), .ZN(n1063) );
XOR2_X1 U1022 ( .A(KEYINPUT45), .B(n1327), .Z(n1326) );
NOR4_X1 U1023 ( .A1(G898), .A2(n1328), .A3(n1293), .A4(n1115), .ZN(n1327) );
INV_X1 U1024 ( .A(n1261), .ZN(n1328) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1261) );
XNOR2_X1 U1026 ( .A(n1078), .B(KEYINPUT59), .ZN(n1231) );
INV_X1 U1027 ( .A(n1258), .ZN(n1078) );
NAND2_X1 U1028 ( .A1(n1329), .A2(n1080), .ZN(n1258) );
NAND2_X1 U1029 ( .A1(G214), .A2(n1330), .ZN(n1080) );
XOR2_X1 U1030 ( .A(n1079), .B(KEYINPUT32), .Z(n1329) );
XOR2_X1 U1031 ( .A(n1104), .B(KEYINPUT23), .Z(n1079) );
XOR2_X1 U1032 ( .A(n1331), .B(n1204), .Z(n1104) );
AND2_X1 U1033 ( .A1(G210), .A2(n1330), .ZN(n1204) );
NAND2_X1 U1034 ( .A1(n1298), .A2(n1293), .ZN(n1330) );
NAND2_X1 U1035 ( .A1(n1332), .A2(n1293), .ZN(n1331) );
XNOR2_X1 U1036 ( .A(n1333), .B(n1334), .ZN(n1332) );
INV_X1 U1037 ( .A(n1201), .ZN(n1334) );
XNOR2_X1 U1038 ( .A(n1335), .B(n1336), .ZN(n1201) );
XOR2_X1 U1039 ( .A(n1152), .B(n1337), .Z(n1336) );
NAND2_X1 U1040 ( .A1(KEYINPUT56), .A2(n1150), .ZN(n1337) );
XNOR2_X1 U1041 ( .A(n1313), .B(n1338), .ZN(n1150) );
XNOR2_X1 U1042 ( .A(n1056), .B(G104), .ZN(n1338) );
INV_X1 U1043 ( .A(G101), .ZN(n1313) );
NAND2_X1 U1044 ( .A1(n1339), .A2(n1340), .ZN(n1152) );
NAND2_X1 U1045 ( .A1(G122), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1046 ( .A(KEYINPUT2), .B(n1342), .Z(n1339) );
NOR2_X1 U1047 ( .A1(G122), .A2(n1341), .ZN(n1342) );
INV_X1 U1048 ( .A(G110), .ZN(n1341) );
XOR2_X1 U1049 ( .A(n1151), .B(n1343), .Z(n1335) );
AND2_X1 U1050 ( .A1(n1115), .A2(G224), .ZN(n1343) );
NAND2_X1 U1051 ( .A1(n1344), .A2(n1345), .ZN(n1151) );
OR2_X1 U1052 ( .A1(n1305), .A2(G113), .ZN(n1345) );
XOR2_X1 U1053 ( .A(n1346), .B(KEYINPUT40), .Z(n1344) );
NAND2_X1 U1054 ( .A1(n1347), .A2(n1305), .ZN(n1346) );
XNOR2_X1 U1055 ( .A(G116), .B(n1348), .ZN(n1305) );
INV_X1 U1056 ( .A(G119), .ZN(n1348) );
XNOR2_X1 U1057 ( .A(KEYINPUT52), .B(n1303), .ZN(n1347) );
INV_X1 U1058 ( .A(G113), .ZN(n1303) );
NOR2_X1 U1059 ( .A1(KEYINPUT33), .A2(n1349), .ZN(n1333) );
XOR2_X1 U1060 ( .A(n1202), .B(KEYINPUT34), .Z(n1349) );
XNOR2_X1 U1061 ( .A(n1304), .B(G125), .ZN(n1202) );
XOR2_X1 U1062 ( .A(G128), .B(n1350), .Z(n1304) );
NOR2_X1 U1063 ( .A1(n1219), .A2(n1218), .ZN(n1068) );
XNOR2_X1 U1064 ( .A(n1103), .B(G475), .ZN(n1218) );
NAND2_X1 U1065 ( .A1(n1166), .A2(n1293), .ZN(n1103) );
XNOR2_X1 U1066 ( .A(n1351), .B(n1352), .ZN(n1166) );
XOR2_X1 U1067 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1068 ( .A(G125), .B(G122), .Z(n1354) );
XNOR2_X1 U1069 ( .A(n1282), .B(G131), .ZN(n1353) );
INV_X1 U1070 ( .A(G140), .ZN(n1282) );
XOR2_X1 U1071 ( .A(n1355), .B(n1356), .Z(n1351) );
XOR2_X1 U1072 ( .A(n1357), .B(n1350), .Z(n1356) );
XOR2_X1 U1073 ( .A(G143), .B(G146), .Z(n1350) );
AND3_X1 U1074 ( .A1(G214), .A2(n1115), .A3(n1298), .ZN(n1357) );
INV_X1 U1075 ( .A(G237), .ZN(n1298) );
XNOR2_X1 U1076 ( .A(G104), .B(G113), .ZN(n1355) );
XNOR2_X1 U1077 ( .A(n1358), .B(G478), .ZN(n1219) );
NAND2_X1 U1078 ( .A1(n1163), .A2(n1293), .ZN(n1358) );
INV_X1 U1079 ( .A(G902), .ZN(n1293) );
XOR2_X1 U1080 ( .A(n1359), .B(n1360), .Z(n1163) );
XOR2_X1 U1081 ( .A(n1361), .B(n1362), .Z(n1360) );
XNOR2_X1 U1082 ( .A(n1292), .B(G122), .ZN(n1362) );
INV_X1 U1083 ( .A(G128), .ZN(n1292) );
XNOR2_X1 U1084 ( .A(KEYINPUT39), .B(n1127), .ZN(n1361) );
INV_X1 U1085 ( .A(G134), .ZN(n1127) );
XOR2_X1 U1086 ( .A(n1363), .B(n1364), .Z(n1359) );
XNOR2_X1 U1087 ( .A(G116), .B(n1056), .ZN(n1364) );
INV_X1 U1088 ( .A(G107), .ZN(n1056) );
XOR2_X1 U1089 ( .A(n1365), .B(n1366), .Z(n1363) );
NOR2_X1 U1090 ( .A1(G143), .A2(KEYINPUT22), .ZN(n1366) );
NAND2_X1 U1091 ( .A1(G217), .A2(n1278), .ZN(n1365) );
AND2_X1 U1092 ( .A1(G234), .A2(n1115), .ZN(n1278) );
INV_X1 U1093 ( .A(G953), .ZN(n1115) );
endmodule


