//Key = 1001100100000110100101001101001010000100111101011001011000011101


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274;

XNOR2_X1 U1267 ( .A(n1923), .B(KEYINPUT30), .ZN(n1705) );
INV_X2 U1268 ( .A(n1705), .ZN(n1706) );
NAND2_X2 U1269 ( .A1(n1707), .A2(n2274), .ZN(n1854) );
XOR2_X1 U1270 ( .A(n1707), .B(KEYINPUT19), .Z(U375) );
NAND2_X1 U1271 ( .A1(n1708), .A2(n1709), .ZN(U344) );
NAND2_X1 U1272 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1710), .ZN(n1709) );
NAND2_X1 U1273 ( .A1(n1711), .A2(DATA_IN_7_), .ZN(n1708) );
NAND2_X1 U1274 ( .A1(n1712), .A2(n1713), .ZN(U343) );
NAND2_X1 U1275 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1710), .ZN(n1713) );
NAND2_X1 U1276 ( .A1(n1711), .A2(DATA_IN_6_), .ZN(n1712) );
NAND2_X1 U1277 ( .A1(n1714), .A2(n1715), .ZN(U342) );
NAND2_X1 U1278 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1710), .ZN(n1715) );
XOR2_X1 U1279 ( .A(n1716), .B(KEYINPUT35), .Z(n1714) );
NAND2_X1 U1280 ( .A1(n1711), .A2(DATA_IN_5_), .ZN(n1716) );
NAND2_X1 U1281 ( .A1(n1717), .A2(n1718), .ZN(U341) );
NAND2_X1 U1282 ( .A1(n1719), .A2(DATA_IN_4_), .ZN(n1718) );
XOR2_X1 U1283 ( .A(n1710), .B(KEYINPUT54), .Z(n1719) );
XOR2_X1 U1284 ( .A(KEYINPUT59), .B(n1720), .Z(n1717) );
NOR2_X1 U1285 ( .A1(n1711), .A2(n1721), .ZN(n1720) );
XNOR2_X1 U1286 ( .A(RMAX_REG_4__SCAN_IN), .B(KEYINPUT9), .ZN(n1721) );
NAND2_X1 U1287 ( .A1(n1722), .A2(n1723), .ZN(U340) );
NAND2_X1 U1288 ( .A1(n1724), .A2(DATA_IN_3_), .ZN(n1723) );
XOR2_X1 U1289 ( .A(n1710), .B(KEYINPUT43), .Z(n1724) );
NAND2_X1 U1290 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1710), .ZN(n1722) );
NAND2_X1 U1291 ( .A1(n1725), .A2(n1726), .ZN(U339) );
NAND2_X1 U1292 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1710), .ZN(n1726) );
NAND2_X1 U1293 ( .A1(n1711), .A2(DATA_IN_2_), .ZN(n1725) );
NAND2_X1 U1294 ( .A1(n1727), .A2(n1728), .ZN(U338) );
NAND2_X1 U1295 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1710), .ZN(n1728) );
NAND2_X1 U1296 ( .A1(n1711), .A2(DATA_IN_1_), .ZN(n1727) );
NAND2_X1 U1297 ( .A1(n1729), .A2(n1730), .ZN(U337) );
NAND2_X1 U1298 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1710), .ZN(n1730) );
NAND2_X1 U1299 ( .A1(n1731), .A2(n1711), .ZN(n1729) );
INV_X1 U1300 ( .A(n1710), .ZN(n1711) );
NAND2_X1 U1301 ( .A1(n1707), .A2(n1732), .ZN(n1710) );
NAND3_X1 U1302 ( .A1(n1733), .A2(n1734), .A3(n1735), .ZN(n1732) );
XOR2_X1 U1303 ( .A(KEYINPUT46), .B(DATA_IN_0_), .Z(n1731) );
NAND2_X1 U1304 ( .A1(n1736), .A2(n1737), .ZN(U336) );
NAND2_X1 U1305 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1738), .ZN(n1737) );
NAND2_X1 U1306 ( .A1(n1739), .A2(DATA_IN_7_), .ZN(n1736) );
NAND2_X1 U1307 ( .A1(n1740), .A2(n1741), .ZN(U335) );
NAND2_X1 U1308 ( .A1(n1739), .A2(DATA_IN_6_), .ZN(n1741) );
XOR2_X1 U1309 ( .A(KEYINPUT32), .B(n1742), .Z(n1740) );
NOR2_X1 U1310 ( .A1(n1739), .A2(n1743), .ZN(n1742) );
NAND2_X1 U1311 ( .A1(n1744), .A2(n1745), .ZN(U334) );
NAND2_X1 U1312 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1738), .ZN(n1745) );
NAND2_X1 U1313 ( .A1(n1739), .A2(DATA_IN_5_), .ZN(n1744) );
NAND2_X1 U1314 ( .A1(n1746), .A2(n1747), .ZN(U333) );
NAND2_X1 U1315 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1738), .ZN(n1747) );
NAND2_X1 U1316 ( .A1(n1739), .A2(DATA_IN_4_), .ZN(n1746) );
NAND2_X1 U1317 ( .A1(n1748), .A2(n1749), .ZN(U332) );
NAND2_X1 U1318 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1738), .ZN(n1749) );
NAND2_X1 U1319 ( .A1(n1739), .A2(DATA_IN_3_), .ZN(n1748) );
NAND2_X1 U1320 ( .A1(n1750), .A2(n1751), .ZN(U331) );
NAND2_X1 U1321 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1738), .ZN(n1751) );
NAND2_X1 U1322 ( .A1(n1739), .A2(DATA_IN_2_), .ZN(n1750) );
NAND2_X1 U1323 ( .A1(n1752), .A2(n1753), .ZN(U330) );
NAND2_X1 U1324 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1738), .ZN(n1753) );
NAND2_X1 U1325 ( .A1(n1739), .A2(DATA_IN_1_), .ZN(n1752) );
NAND2_X1 U1326 ( .A1(n1754), .A2(n1755), .ZN(U329) );
NAND2_X1 U1327 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1738), .ZN(n1755) );
NAND2_X1 U1328 ( .A1(n1739), .A2(DATA_IN_0_), .ZN(n1754) );
INV_X1 U1329 ( .A(n1738), .ZN(n1739) );
NAND2_X1 U1330 ( .A1(n1707), .A2(n1756), .ZN(n1738) );
NAND2_X1 U1331 ( .A1(n1734), .A2(n1757), .ZN(n1756) );
NAND3_X1 U1332 ( .A1(n1758), .A2(n1733), .A3(n1735), .ZN(n1757) );
XNOR2_X1 U1333 ( .A(n1759), .B(KEYINPUT0), .ZN(n1735) );
NAND2_X1 U1334 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1760), .ZN(n1759) );
NAND3_X1 U1335 ( .A1(n1761), .A2(n1762), .A3(n1763), .ZN(n1733) );
OR2_X1 U1336 ( .A1(n1760), .A2(RMAX_REG_7__SCAN_IN), .ZN(n1763) );
NAND3_X1 U1337 ( .A1(n1764), .A2(n1765), .A3(n1766), .ZN(n1762) );
OR2_X1 U1338 ( .A1(n1767), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1766) );
NAND3_X1 U1339 ( .A1(n1768), .A2(n1769), .A3(n1770), .ZN(n1765) );
NAND2_X1 U1340 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1771), .ZN(n1770) );
NAND3_X1 U1341 ( .A1(n1772), .A2(n1773), .A3(n1774), .ZN(n1769) );
OR2_X1 U1342 ( .A1(n1775), .A2(RMAX_REG_4__SCAN_IN), .ZN(n1774) );
NAND3_X1 U1343 ( .A1(n1776), .A2(n1777), .A3(n1778), .ZN(n1773) );
XOR2_X1 U1344 ( .A(KEYINPUT51), .B(n1779), .Z(n1778) );
NOR3_X1 U1345 ( .A1(n1780), .A2(n1781), .A3(n1782), .ZN(n1779) );
NOR2_X1 U1346 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1783), .ZN(n1782) );
NOR3_X1 U1347 ( .A1(n1784), .A2(RMAX_REG_0__SCAN_IN), .A3(n1785), .ZN(n1781));
NOR2_X1 U1348 ( .A1(DATA_IN_1_), .A2(n1786), .ZN(n1785) );
NOR2_X1 U1349 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1787), .ZN(n1780) );
NAND2_X1 U1350 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1788), .ZN(n1777) );
XOR2_X1 U1351 ( .A(KEYINPUT4), .B(DATA_IN_2_), .Z(n1788) );
NAND2_X1 U1352 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1789), .ZN(n1776) );
NAND2_X1 U1353 ( .A1(DATA_IN_3_), .A2(n1790), .ZN(n1772) );
XOR2_X1 U1354 ( .A(RMAX_REG_3__SCAN_IN), .B(KEYINPUT63), .Z(n1790) );
NAND2_X1 U1355 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1775), .ZN(n1768) );
NAND2_X1 U1356 ( .A1(n1791), .A2(DATA_IN_5_), .ZN(n1764) );
XOR2_X1 U1357 ( .A(n1792), .B(KEYINPUT17), .Z(n1791) );
NAND2_X1 U1358 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1767), .ZN(n1761) );
NAND2_X1 U1359 ( .A1(n1793), .A2(n1794), .ZN(n1758) );
NAND2_X1 U1360 ( .A1(DATA_IN_7_), .A2(n1795), .ZN(n1794) );
XOR2_X1 U1361 ( .A(KEYINPUT60), .B(n1796), .Z(n1793) );
NOR3_X1 U1362 ( .A1(n1797), .A2(n1798), .A3(n1799), .ZN(n1796) );
NOR2_X1 U1363 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1767), .ZN(n1799) );
INV_X1 U1364 ( .A(DATA_IN_6_), .ZN(n1767) );
NOR2_X1 U1365 ( .A1(DATA_IN_7_), .A2(n1795), .ZN(n1798) );
NOR3_X1 U1366 ( .A1(n1800), .A2(n1801), .A3(n1802), .ZN(n1797) );
AND2_X1 U1367 ( .A1(n1771), .A2(n1803), .ZN(n1802) );
NOR2_X1 U1368 ( .A1(n1804), .A2(n1805), .ZN(n1801) );
NOR2_X1 U1369 ( .A1(n1771), .A2(n1803), .ZN(n1804) );
NAND2_X1 U1370 ( .A1(n1806), .A2(n1807), .ZN(n1803) );
NAND2_X1 U1371 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1808), .ZN(n1807) );
NAND2_X1 U1372 ( .A1(DATA_IN_4_), .A2(n1809), .ZN(n1808) );
OR2_X1 U1373 ( .A1(n1809), .A2(DATA_IN_4_), .ZN(n1806) );
NAND2_X1 U1374 ( .A1(n1810), .A2(n1811), .ZN(n1809) );
NAND2_X1 U1375 ( .A1(n1812), .A2(n1813), .ZN(n1811) );
NAND2_X1 U1376 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1789), .ZN(n1813) );
NAND2_X1 U1377 ( .A1(n1814), .A2(n1815), .ZN(n1812) );
NAND2_X1 U1378 ( .A1(DATA_IN_2_), .A2(n1816), .ZN(n1815) );
NAND4_X1 U1379 ( .A1(n1817), .A2(n1818), .A3(n1819), .A4(n1820), .ZN(n1814));
NAND3_X1 U1380 ( .A1(n1784), .A2(n1787), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1820) );
NAND2_X1 U1381 ( .A1(n1821), .A2(RMIN_REG_2__SCAN_IN), .ZN(n1819) );
XOR2_X1 U1382 ( .A(n1783), .B(KEYINPUT56), .Z(n1821) );
NAND2_X1 U1383 ( .A1(KEYINPUT10), .A2(n1822), .ZN(n1818) );
NAND2_X1 U1384 ( .A1(n1823), .A2(RMIN_REG_1__SCAN_IN), .ZN(n1822) );
NAND2_X1 U1385 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1824), .ZN(n1817) );
NAND2_X1 U1386 ( .A1(n1825), .A2(n1826), .ZN(n1824) );
NAND2_X1 U1387 ( .A1(n1823), .A2(n1827), .ZN(n1826) );
INV_X1 U1388 ( .A(KEYINPUT10), .ZN(n1827) );
XOR2_X1 U1389 ( .A(KEYINPUT2), .B(n1787), .Z(n1823) );
NAND2_X1 U1390 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1784), .ZN(n1825) );
NAND2_X1 U1391 ( .A1(DATA_IN_3_), .A2(n1828), .ZN(n1810) );
NOR2_X1 U1392 ( .A1(DATA_IN_6_), .A2(n1743), .ZN(n1800) );
NAND2_X1 U1393 ( .A1(n1829), .A2(n1830), .ZN(U328) );
NAND2_X1 U1394 ( .A1(n1831), .A2(DATA_IN_7_), .ZN(n1830) );
NAND2_X1 U1395 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1832), .ZN(n1829) );
NAND2_X1 U1396 ( .A1(n1833), .A2(n1834), .ZN(U327) );
NAND2_X1 U1397 ( .A1(DATA_IN_6_), .A2(n1835), .ZN(n1834) );
XOR2_X1 U1398 ( .A(KEYINPUT20), .B(n1831), .Z(n1835) );
NAND2_X1 U1399 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1832), .ZN(n1833) );
NAND2_X1 U1400 ( .A1(n1836), .A2(n1837), .ZN(U326) );
NAND2_X1 U1401 ( .A1(n1831), .A2(DATA_IN_5_), .ZN(n1837) );
NAND2_X1 U1402 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1832), .ZN(n1836) );
NAND2_X1 U1403 ( .A1(n1838), .A2(n1839), .ZN(U325) );
NAND2_X1 U1404 ( .A1(n1831), .A2(DATA_IN_4_), .ZN(n1839) );
NAND2_X1 U1405 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1832), .ZN(n1838) );
NAND2_X1 U1406 ( .A1(n1840), .A2(n1841), .ZN(U324) );
NAND2_X1 U1407 ( .A1(n1831), .A2(DATA_IN_3_), .ZN(n1841) );
NAND2_X1 U1408 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1832), .ZN(n1840) );
NAND2_X1 U1409 ( .A1(n1842), .A2(n1843), .ZN(U323) );
NAND2_X1 U1410 ( .A1(n1831), .A2(DATA_IN_2_), .ZN(n1843) );
NAND2_X1 U1411 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1832), .ZN(n1842) );
NAND2_X1 U1412 ( .A1(n1844), .A2(n1845), .ZN(U322) );
NAND2_X1 U1413 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1832), .ZN(n1845) );
XOR2_X1 U1414 ( .A(KEYINPUT41), .B(n1846), .Z(n1844) );
NOR2_X1 U1415 ( .A1(n1787), .A2(n1847), .ZN(n1846) );
NAND2_X1 U1416 ( .A1(n1848), .A2(n1849), .ZN(U321) );
NAND2_X1 U1417 ( .A1(n1831), .A2(DATA_IN_0_), .ZN(n1849) );
INV_X1 U1418 ( .A(n1847), .ZN(n1831) );
NAND2_X1 U1419 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1850), .ZN(n1847) );
NAND2_X1 U1420 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1832), .ZN(n1848) );
NAND2_X1 U1421 ( .A1(n1707), .A2(n1850), .ZN(n1832) );
NAND2_X1 U1422 ( .A1(n1851), .A2(n1734), .ZN(n1850) );
NAND2_X1 U1423 ( .A1(n1852), .A2(n1853), .ZN(U320) );
NAND2_X1 U1424 ( .A1(n1706), .A2(DATA_IN_7_), .ZN(n1853) );
NAND2_X1 U1425 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1854), .ZN(n1852) );
NAND2_X1 U1426 ( .A1(n1855), .A2(n1856), .ZN(U319) );
NAND2_X1 U1427 ( .A1(n1706), .A2(DATA_IN_6_), .ZN(n1856) );
NAND2_X1 U1428 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1854), .ZN(n1855) );
NAND2_X1 U1429 ( .A1(n1857), .A2(n1858), .ZN(U318) );
NAND2_X1 U1430 ( .A1(n1859), .A2(n1854), .ZN(n1858) );
XOR2_X1 U1431 ( .A(REG1_REG_5__SCAN_IN), .B(KEYINPUT36), .Z(n1859) );
NAND2_X1 U1432 ( .A1(n1860), .A2(DATA_IN_5_), .ZN(n1857) );
XOR2_X1 U1433 ( .A(n1706), .B(KEYINPUT55), .Z(n1860) );
NAND2_X1 U1434 ( .A1(n1861), .A2(n1862), .ZN(U317) );
NAND2_X1 U1435 ( .A1(n1706), .A2(DATA_IN_4_), .ZN(n1862) );
NAND2_X1 U1436 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1854), .ZN(n1861) );
NAND2_X1 U1437 ( .A1(n1863), .A2(n1864), .ZN(U316) );
NAND2_X1 U1438 ( .A1(n1706), .A2(DATA_IN_3_), .ZN(n1864) );
NAND2_X1 U1439 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1854), .ZN(n1863) );
NAND2_X1 U1440 ( .A1(n1865), .A2(n1866), .ZN(U315) );
NAND2_X1 U1441 ( .A1(n1706), .A2(DATA_IN_2_), .ZN(n1866) );
NAND2_X1 U1442 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1854), .ZN(n1865) );
NAND2_X1 U1443 ( .A1(n1867), .A2(n1868), .ZN(U314) );
NAND2_X1 U1444 ( .A1(n1706), .A2(DATA_IN_1_), .ZN(n1868) );
NAND2_X1 U1445 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1854), .ZN(n1867) );
NAND2_X1 U1446 ( .A1(n1869), .A2(n1870), .ZN(U313) );
NAND2_X1 U1447 ( .A1(n1706), .A2(DATA_IN_0_), .ZN(n1870) );
NAND2_X1 U1448 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1854), .ZN(n1869) );
NAND2_X1 U1449 ( .A1(n1871), .A2(n1872), .ZN(U312) );
NAND2_X1 U1450 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1706), .ZN(n1872) );
NAND2_X1 U1451 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1854), .ZN(n1871) );
NAND2_X1 U1452 ( .A1(n1873), .A2(n1874), .ZN(U311) );
NAND2_X1 U1453 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1706), .ZN(n1874) );
NAND2_X1 U1454 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1854), .ZN(n1873) );
NAND2_X1 U1455 ( .A1(n1875), .A2(n1876), .ZN(U310) );
NAND2_X1 U1456 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1706), .ZN(n1876) );
NAND2_X1 U1457 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1854), .ZN(n1875) );
NAND2_X1 U1458 ( .A1(n1877), .A2(n1878), .ZN(U309) );
NAND2_X1 U1459 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1706), .ZN(n1878) );
NAND2_X1 U1460 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1854), .ZN(n1877) );
NAND2_X1 U1461 ( .A1(n1879), .A2(n1880), .ZN(U308) );
NAND2_X1 U1462 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1881), .ZN(n1880) );
XNOR2_X1 U1463 ( .A(KEYINPUT27), .B(n1706), .ZN(n1881) );
NAND2_X1 U1464 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1854), .ZN(n1879) );
NAND2_X1 U1465 ( .A1(n1882), .A2(n1883), .ZN(U307) );
NAND2_X1 U1466 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1706), .ZN(n1883) );
NAND2_X1 U1467 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1854), .ZN(n1882) );
NAND2_X1 U1468 ( .A1(n1884), .A2(n1885), .ZN(U306) );
NAND2_X1 U1469 ( .A1(n1706), .A2(n1886), .ZN(n1885) );
XOR2_X1 U1470 ( .A(REG1_REG_1__SCAN_IN), .B(KEYINPUT57), .Z(n1886) );
NAND2_X1 U1471 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1854), .ZN(n1884) );
NAND2_X1 U1472 ( .A1(n1887), .A2(n1888), .ZN(U305) );
NAND2_X1 U1473 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1706), .ZN(n1888) );
NAND2_X1 U1474 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1854), .ZN(n1887) );
NAND2_X1 U1475 ( .A1(n1889), .A2(n1890), .ZN(U304) );
NAND2_X1 U1476 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1706), .ZN(n1890) );
NAND2_X1 U1477 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1854), .ZN(n1889) );
NAND2_X1 U1478 ( .A1(n1891), .A2(n1892), .ZN(U303) );
NAND2_X1 U1479 ( .A1(n1706), .A2(n1893), .ZN(n1892) );
XOR2_X1 U1480 ( .A(REG2_REG_6__SCAN_IN), .B(KEYINPUT23), .Z(n1893) );
NAND2_X1 U1481 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1854), .ZN(n1891) );
NAND2_X1 U1482 ( .A1(n1894), .A2(n1895), .ZN(U302) );
NAND2_X1 U1483 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1706), .ZN(n1895) );
NAND2_X1 U1484 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1854), .ZN(n1894) );
NAND2_X1 U1485 ( .A1(n1896), .A2(n1897), .ZN(U301) );
NAND2_X1 U1486 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1706), .ZN(n1897) );
NAND2_X1 U1487 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1854), .ZN(n1896) );
NAND2_X1 U1488 ( .A1(n1898), .A2(n1899), .ZN(U300) );
NAND2_X1 U1489 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1854), .ZN(n1899) );
XOR2_X1 U1490 ( .A(n1900), .B(KEYINPUT44), .Z(n1898) );
NAND2_X1 U1491 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1706), .ZN(n1900) );
NAND2_X1 U1492 ( .A1(n1901), .A2(n1902), .ZN(U299) );
NAND2_X1 U1493 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1706), .ZN(n1902) );
NAND2_X1 U1494 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1854), .ZN(n1901) );
NAND2_X1 U1495 ( .A1(n1903), .A2(n1904), .ZN(U298) );
NAND2_X1 U1496 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1706), .ZN(n1904) );
NAND2_X1 U1497 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1854), .ZN(n1903) );
NAND2_X1 U1498 ( .A1(n1905), .A2(n1906), .ZN(U297) );
NAND2_X1 U1499 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1706), .ZN(n1906) );
NAND2_X1 U1500 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1854), .ZN(n1905) );
NAND2_X1 U1501 ( .A1(n1907), .A2(n1908), .ZN(U296) );
NAND2_X1 U1502 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1706), .ZN(n1908) );
NAND2_X1 U1503 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1854), .ZN(n1907) );
NAND2_X1 U1504 ( .A1(n1909), .A2(n1910), .ZN(U295) );
NAND2_X1 U1505 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1706), .ZN(n1910) );
NAND2_X1 U1506 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1854), .ZN(n1909) );
NAND2_X1 U1507 ( .A1(n1911), .A2(n1912), .ZN(U294) );
NAND2_X1 U1508 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1706), .ZN(n1912) );
NAND2_X1 U1509 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1854), .ZN(n1911) );
NAND2_X1 U1510 ( .A1(n1913), .A2(n1914), .ZN(U293) );
NAND2_X1 U1511 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1706), .ZN(n1914) );
NAND2_X1 U1512 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1854), .ZN(n1913) );
NAND2_X1 U1513 ( .A1(n1915), .A2(n1916), .ZN(U292) );
NAND2_X1 U1514 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1706), .ZN(n1916) );
NAND2_X1 U1515 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1854), .ZN(n1915) );
NAND2_X1 U1516 ( .A1(n1917), .A2(n1918), .ZN(U291) );
NAND2_X1 U1517 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1706), .ZN(n1918) );
NAND2_X1 U1518 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1854), .ZN(n1917) );
NAND2_X1 U1519 ( .A1(n1919), .A2(n1920), .ZN(U290) );
NAND2_X1 U1520 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1706), .ZN(n1920) );
NAND2_X1 U1521 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1854), .ZN(n1919) );
NAND2_X1 U1522 ( .A1(n1921), .A2(n1922), .ZN(U289) );
NAND2_X1 U1523 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1706), .ZN(n1922) );
NAND2_X1 U1524 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1734), .ZN(n1923) );
INV_X1 U1525 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1734) );
NAND2_X1 U1526 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1854), .ZN(n1921) );
NAND4_X1 U1527 ( .A1(n1924), .A2(n1925), .A3(n1926), .A4(n1927), .ZN(U288));
NAND2_X1 U1528 ( .A1(n1928), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1927) );
NAND2_X1 U1529 ( .A1(n1929), .A2(REG4_REG_7__SCAN_IN), .ZN(n1926) );
NAND2_X1 U1530 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1854), .ZN(n1925) );
NAND4_X1 U1531 ( .A1(n1930), .A2(n1931), .A3(n1924), .A4(n1932), .ZN(U287));
NOR3_X1 U1532 ( .A1(n1933), .A2(n1934), .A3(n1935), .ZN(n1932) );
NOR3_X1 U1533 ( .A1(n1936), .A2(n1937), .A3(n1938), .ZN(n1935) );
NOR4_X1 U1534 ( .A1(n1939), .A2(n1940), .A3(n1941), .A4(n1942), .ZN(n1934));
AND2_X1 U1535 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1928), .ZN(n1933) );
AND2_X1 U1536 ( .A1(n1943), .A2(n1944), .ZN(n1924) );
NAND3_X1 U1537 ( .A1(n1937), .A2(n1936), .A3(n1945), .ZN(n1944) );
NAND2_X1 U1538 ( .A1(n1946), .A2(n1947), .ZN(n1936) );
XOR2_X1 U1539 ( .A(n1948), .B(KEYINPUT61), .Z(n1946) );
INV_X1 U1540 ( .A(n1949), .ZN(n1937) );
NAND3_X1 U1541 ( .A1(n1950), .A2(n1939), .A3(n1940), .ZN(n1943) );
NAND2_X1 U1542 ( .A1(n1929), .A2(REG4_REG_6__SCAN_IN), .ZN(n1931) );
NAND2_X1 U1543 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1854), .ZN(n1930) );
NAND4_X1 U1544 ( .A1(n1951), .A2(n1952), .A3(n1953), .A4(n1954), .ZN(U286));
NOR3_X1 U1545 ( .A1(n1955), .A2(n1956), .A3(n1957), .ZN(n1954) );
NOR2_X1 U1546 ( .A1(n1958), .A2(n1938), .ZN(n1957) );
XOR2_X1 U1547 ( .A(n1959), .B(n1960), .Z(n1958) );
NAND2_X1 U1548 ( .A1(KEYINPUT61), .A2(n1947), .ZN(n1959) );
NAND2_X1 U1549 ( .A1(n1961), .A2(n1949), .ZN(n1947) );
NAND3_X1 U1550 ( .A1(n1962), .A2(n1963), .A3(n1964), .ZN(n1949) );
NAND2_X1 U1551 ( .A1(n1965), .A2(n1966), .ZN(n1961) );
NAND2_X1 U1552 ( .A1(n1964), .A2(n1962), .ZN(n1966) );
NOR2_X1 U1553 ( .A1(n1941), .A2(n1967), .ZN(n1956) );
XOR2_X1 U1554 ( .A(n1940), .B(n1968), .Z(n1967) );
AND3_X1 U1555 ( .A1(n1969), .A2(n1970), .A3(n1971), .ZN(n1940) );
NAND2_X1 U1556 ( .A1(n1972), .A2(n1973), .ZN(n1971) );
XOR2_X1 U1557 ( .A(KEYINPUT18), .B(n1965), .Z(n1972) );
NAND3_X1 U1558 ( .A1(n1974), .A2(n1965), .A3(KEYINPUT15), .ZN(n1970) );
NAND2_X1 U1559 ( .A1(n1939), .A2(n1975), .ZN(n1969) );
INV_X1 U1560 ( .A(KEYINPUT15), .ZN(n1975) );
NOR2_X1 U1561 ( .A1(n1973), .A2(n1965), .ZN(n1939) );
INV_X1 U1562 ( .A(n1963), .ZN(n1965) );
NOR2_X1 U1563 ( .A1(n1963), .A2(n1976), .ZN(n1955) );
NAND2_X1 U1564 ( .A1(n1977), .A2(n1978), .ZN(n1963) );
NAND4_X1 U1565 ( .A1(n1979), .A2(n1980), .A3(n1981), .A4(n1982), .ZN(n1978));
XOR2_X1 U1566 ( .A(KEYINPUT7), .B(n1983), .Z(n1979) );
AND2_X1 U1567 ( .A1(n1984), .A2(n1985), .ZN(n1983) );
NAND3_X1 U1568 ( .A1(n1986), .A2(n1984), .A3(n1987), .ZN(n1977) );
NAND2_X1 U1569 ( .A1(n1981), .A2(n1982), .ZN(n1987) );
NAND3_X1 U1570 ( .A1(n1988), .A2(n1989), .A3(n1990), .ZN(n1982) );
XOR2_X1 U1571 ( .A(n1991), .B(KEYINPUT48), .Z(n1990) );
NAND2_X1 U1572 ( .A1(RESTART), .A2(n1743), .ZN(n1989) );
NAND2_X1 U1573 ( .A1(n1992), .A2(n1993), .ZN(n1988) );
NAND3_X1 U1574 ( .A1(n1994), .A2(n1995), .A3(n1991), .ZN(n1981) );
NAND2_X1 U1575 ( .A1(n1996), .A2(n1997), .ZN(n1991) );
NAND2_X1 U1576 ( .A1(DATA_IN_6_), .A2(n1993), .ZN(n1997) );
NAND2_X1 U1577 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1996) );
NAND2_X1 U1578 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1993), .ZN(n1995) );
NAND2_X1 U1579 ( .A1(RESTART), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1994) );
NAND2_X1 U1580 ( .A1(n1998), .A2(n1999), .ZN(n1984) );
NAND2_X1 U1581 ( .A1(n2000), .A2(n2001), .ZN(n1986) );
XNOR2_X1 U1582 ( .A(KEYINPUT3), .B(n1980), .ZN(n2001) );
OR2_X1 U1583 ( .A1(n1999), .A2(n1998), .ZN(n1980) );
NAND2_X1 U1584 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1854), .ZN(n1953) );
NAND2_X1 U1585 ( .A1(n1928), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1952) );
NAND2_X1 U1586 ( .A1(n1929), .A2(REG4_REG_5__SCAN_IN), .ZN(n1951) );
NAND4_X1 U1587 ( .A1(n2002), .A2(n2003), .A3(n2004), .A4(n2005), .ZN(U285));
NOR3_X1 U1588 ( .A1(n2006), .A2(n2007), .A3(n2008), .ZN(n2005) );
NOR3_X1 U1589 ( .A1(n1938), .A2(n1960), .A3(n2009), .ZN(n2008) );
NOR2_X1 U1590 ( .A1(n2010), .A2(n2011), .ZN(n2009) );
XOR2_X1 U1591 ( .A(KEYINPUT28), .B(n2012), .Z(n2011) );
INV_X1 U1592 ( .A(n1948), .ZN(n1960) );
NAND2_X1 U1593 ( .A1(n2012), .A2(n2010), .ZN(n1948) );
XOR2_X1 U1594 ( .A(n2013), .B(n1964), .Z(n2010) );
NOR3_X1 U1595 ( .A1(n1941), .A2(n1968), .A3(n2014), .ZN(n2007) );
NOR2_X1 U1596 ( .A1(n2015), .A2(n2013), .ZN(n2014) );
INV_X1 U1597 ( .A(n1942), .ZN(n1968) );
NAND2_X1 U1598 ( .A1(n2015), .A2(n2016), .ZN(n1942) );
NAND2_X1 U1599 ( .A1(n2017), .A2(n1973), .ZN(n2016) );
INV_X1 U1600 ( .A(n1974), .ZN(n1973) );
NOR2_X1 U1601 ( .A1(n2018), .A2(n2013), .ZN(n1974) );
NAND2_X1 U1602 ( .A1(n2013), .A2(n2018), .ZN(n2017) );
NOR2_X1 U1603 ( .A1(n1962), .A2(n1976), .ZN(n2006) );
INV_X1 U1604 ( .A(n2013), .ZN(n1962) );
NAND2_X1 U1605 ( .A1(n2019), .A2(n2020), .ZN(n2013) );
NAND2_X1 U1606 ( .A1(n2000), .A2(n2021), .ZN(n2020) );
XOR2_X1 U1607 ( .A(n2022), .B(KEYINPUT49), .Z(n2019) );
OR2_X1 U1608 ( .A1(n2021), .A2(n2000), .ZN(n2022) );
INV_X1 U1609 ( .A(n1985), .ZN(n2000) );
NAND2_X1 U1610 ( .A1(n2023), .A2(n2024), .ZN(n1985) );
NAND2_X1 U1611 ( .A1(n2025), .A2(n2026), .ZN(n2024) );
XOR2_X1 U1612 ( .A(n2027), .B(KEYINPUT22), .Z(n2025) );
XOR2_X1 U1613 ( .A(n1998), .B(n1999), .Z(n2021) );
NAND2_X1 U1614 ( .A1(n2028), .A2(n2029), .ZN(n1999) );
NAND2_X1 U1615 ( .A1(RESTART), .A2(n1805), .ZN(n2029) );
INV_X1 U1616 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1805) );
NAND2_X1 U1617 ( .A1(n2030), .A2(n1993), .ZN(n2028) );
NAND2_X1 U1618 ( .A1(n2031), .A2(n2032), .ZN(n1998) );
NAND2_X1 U1619 ( .A1(RESTART), .A2(n1792), .ZN(n2032) );
INV_X1 U1620 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1792) );
NAND2_X1 U1621 ( .A1(n1771), .A2(n1993), .ZN(n2031) );
INV_X1 U1622 ( .A(DATA_IN_5_), .ZN(n1771) );
NAND2_X1 U1623 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1854), .ZN(n2004) );
NAND2_X1 U1624 ( .A1(n1928), .A2(RLAST_REG_4__SCAN_IN), .ZN(n2003) );
NAND2_X1 U1625 ( .A1(n1929), .A2(REG4_REG_4__SCAN_IN), .ZN(n2002) );
NAND4_X1 U1626 ( .A1(n2033), .A2(n2034), .A3(n2035), .A4(n2036), .ZN(U284));
NOR3_X1 U1627 ( .A1(n2037), .A2(n2038), .A3(n2039), .ZN(n2036) );
NOR2_X1 U1628 ( .A1(n2040), .A2(n2041), .ZN(n2039) );
INV_X1 U1629 ( .A(RLAST_REG_3__SCAN_IN), .ZN(n2041) );
XNOR2_X1 U1630 ( .A(n1928), .B(KEYINPUT11), .ZN(n2040) );
NOR3_X1 U1631 ( .A1(n2042), .A2(n2043), .A3(n1941), .ZN(n2038) );
NOR2_X1 U1632 ( .A1(n2044), .A2(n2045), .ZN(n2043) );
XOR2_X1 U1633 ( .A(KEYINPUT1), .B(n2015), .Z(n2042) );
AND2_X1 U1634 ( .A1(n2044), .A2(n2045), .ZN(n2015) );
NAND2_X1 U1635 ( .A1(n2018), .A2(n2046), .ZN(n2045) );
NAND2_X1 U1636 ( .A1(n2047), .A2(n2048), .ZN(n2046) );
NAND2_X1 U1637 ( .A1(n2049), .A2(n2050), .ZN(n2048) );
OR3_X1 U1638 ( .A1(n2051), .A2(n2052), .A3(n2047), .ZN(n2018) );
NOR3_X1 U1639 ( .A1(n1938), .A2(n2053), .A3(n2054), .ZN(n2037) );
NOR2_X1 U1640 ( .A1(n2055), .A2(n2056), .ZN(n2054) );
XOR2_X1 U1641 ( .A(n2057), .B(n2058), .Z(n2056) );
INV_X1 U1642 ( .A(KEYINPUT40), .ZN(n2055) );
NOR3_X1 U1643 ( .A1(KEYINPUT40), .A2(n2012), .A3(n2059), .ZN(n2053) );
AND2_X1 U1644 ( .A1(n2057), .A2(n2058), .ZN(n2059) );
NOR2_X1 U1645 ( .A1(n2057), .A2(n2058), .ZN(n2012) );
NOR2_X1 U1646 ( .A1(n2060), .A2(n1964), .ZN(n2058) );
NOR3_X1 U1647 ( .A1(n2051), .A2(n2061), .A3(n2047), .ZN(n1964) );
AND2_X1 U1648 ( .A1(n2047), .A2(n2062), .ZN(n2060) );
NAND2_X1 U1649 ( .A1(n2050), .A2(n2063), .ZN(n2062) );
NAND2_X1 U1650 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1854), .ZN(n2035) );
NAND2_X1 U1651 ( .A1(n2064), .A2(n2047), .ZN(n2034) );
NAND2_X1 U1652 ( .A1(n2065), .A2(n2066), .ZN(n2047) );
NAND2_X1 U1653 ( .A1(n2067), .A2(n2026), .ZN(n2066) );
NAND2_X1 U1654 ( .A1(n2027), .A2(n2023), .ZN(n2067) );
NAND2_X1 U1655 ( .A1(n2068), .A2(n2069), .ZN(n2023) );
OR2_X1 U1656 ( .A1(n2069), .A2(n2068), .ZN(n2027) );
NAND2_X1 U1657 ( .A1(n2070), .A2(n2071), .ZN(n2065) );
XOR2_X1 U1658 ( .A(n2069), .B(n2068), .Z(n2071) );
NAND2_X1 U1659 ( .A1(n2072), .A2(n2073), .ZN(n2068) );
NAND2_X1 U1660 ( .A1(DATA_IN_4_), .A2(n1993), .ZN(n2073) );
NAND2_X1 U1661 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2072) );
NAND3_X1 U1662 ( .A1(n2074), .A2(n2075), .A3(n2076), .ZN(n2069) );
OR2_X1 U1663 ( .A1(KEYINPUT25), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2076) );
NAND3_X1 U1664 ( .A1(KEYINPUT25), .A2(RMIN_REG_4__SCAN_IN), .A3(RESTART),
.ZN(n2075) );
NAND2_X1 U1665 ( .A1(n2077), .A2(n1993), .ZN(n2074) );
NAND2_X1 U1666 ( .A1(KEYINPUT25), .A2(n2078), .ZN(n2077) );
INV_X1 U1667 ( .A(n2026), .ZN(n2070) );
NAND2_X1 U1668 ( .A1(n2079), .A2(n2080), .ZN(n2026) );
NAND2_X1 U1669 ( .A1(n2081), .A2(n2082), .ZN(n2080) );
XOR2_X1 U1670 ( .A(KEYINPUT24), .B(n2083), .Z(n2081) );
NOR2_X1 U1671 ( .A1(n2084), .A2(n2085), .ZN(n2083) );
NAND2_X1 U1672 ( .A1(n2084), .A2(n2085), .ZN(n2079) );
INV_X1 U1673 ( .A(n2086), .ZN(n2084) );
INV_X1 U1674 ( .A(n1976), .ZN(n2064) );
NAND2_X1 U1675 ( .A1(n1929), .A2(REG4_REG_3__SCAN_IN), .ZN(n2033) );
NAND4_X1 U1676 ( .A1(n2087), .A2(n2088), .A3(n2089), .A4(n2090), .ZN(U283));
NOR3_X1 U1677 ( .A1(n2091), .A2(n2092), .A3(n2093), .ZN(n2090) );
NOR3_X1 U1678 ( .A1(n1938), .A2(n2094), .A3(n2095), .ZN(n2093) );
NOR3_X1 U1679 ( .A1(n2096), .A2(n2097), .A3(n2098), .ZN(n2095) );
NOR2_X1 U1680 ( .A1(n2099), .A2(n2051), .ZN(n2098) );
NOR2_X1 U1681 ( .A1(n2100), .A2(n2101), .ZN(n2099) );
NOR2_X1 U1682 ( .A1(n2101), .A2(n2050), .ZN(n2097) );
NOR2_X1 U1683 ( .A1(n2102), .A2(n2103), .ZN(n2096) );
INV_X1 U1684 ( .A(n2057), .ZN(n2094) );
NAND4_X1 U1685 ( .A1(n2104), .A2(n2105), .A3(n2106), .A4(n2107), .ZN(n2057));
NAND2_X1 U1686 ( .A1(n2049), .A2(n2108), .ZN(n2106) );
NAND2_X1 U1687 ( .A1(n2100), .A2(n2050), .ZN(n2108) );
XOR2_X1 U1688 ( .A(KEYINPUT14), .B(n2103), .Z(n2105) );
NOR2_X1 U1689 ( .A1(n2109), .A2(n2110), .ZN(n2104) );
NOR3_X1 U1690 ( .A1(n2101), .A2(n2051), .A3(n2100), .ZN(n2110) );
XOR2_X1 U1691 ( .A(n2063), .B(KEYINPUT5), .Z(n2100) );
INV_X1 U1692 ( .A(n2061), .ZN(n2063) );
XOR2_X1 U1693 ( .A(n2052), .B(KEYINPUT50), .Z(n2061) );
INV_X1 U1694 ( .A(KEYINPUT47), .ZN(n2101) );
NOR2_X1 U1695 ( .A1(KEYINPUT47), .A2(n2050), .ZN(n2109) );
NOR3_X1 U1696 ( .A1(n1941), .A2(n2044), .A3(n2111), .ZN(n2092) );
NOR2_X1 U1697 ( .A1(n2112), .A2(n2113), .ZN(n2111) );
INV_X1 U1698 ( .A(n2114), .ZN(n2113) );
NOR2_X1 U1699 ( .A1(n2102), .A2(n2115), .ZN(n2112) );
NOR3_X1 U1700 ( .A1(n2115), .A2(n2102), .A3(n2114), .ZN(n2044) );
XNOR2_X1 U1701 ( .A(n2051), .B(n2049), .ZN(n2114) );
INV_X1 U1702 ( .A(n2052), .ZN(n2049) );
INV_X1 U1703 ( .A(n2050), .ZN(n2051) );
INV_X1 U1704 ( .A(n2107), .ZN(n2102) );
NOR2_X1 U1705 ( .A1(n2050), .A2(n1976), .ZN(n2091) );
XNOR2_X1 U1706 ( .A(n2116), .B(n2085), .ZN(n2050) );
NAND2_X1 U1707 ( .A1(n2117), .A2(n2118), .ZN(n2085) );
NAND2_X1 U1708 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1993), .ZN(n2118) );
NAND2_X1 U1709 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2117) );
XOR2_X1 U1710 ( .A(n2082), .B(n2119), .Z(n2116) );
NOR2_X1 U1711 ( .A1(KEYINPUT29), .A2(n2086), .ZN(n2119) );
NAND2_X1 U1712 ( .A1(n2120), .A2(n2121), .ZN(n2086) );
NAND2_X1 U1713 ( .A1(RESTART), .A2(n2122), .ZN(n2121) );
NAND2_X1 U1714 ( .A1(n1789), .A2(n1993), .ZN(n2120) );
INV_X1 U1715 ( .A(DATA_IN_3_), .ZN(n1789) );
NAND2_X1 U1716 ( .A1(n2123), .A2(n2124), .ZN(n2082) );
NAND2_X1 U1717 ( .A1(n2125), .A2(n2126), .ZN(n2124) );
NAND2_X1 U1718 ( .A1(n2127), .A2(n2128), .ZN(n2126) );
OR2_X1 U1719 ( .A1(n2128), .A2(n2127), .ZN(n2123) );
NAND2_X1 U1720 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1854), .ZN(n2089) );
NAND2_X1 U1721 ( .A1(n1928), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2088) );
NAND2_X1 U1722 ( .A1(n1929), .A2(REG4_REG_2__SCAN_IN), .ZN(n2087) );
NAND4_X1 U1723 ( .A1(n2129), .A2(n2130), .A3(n2131), .A4(n2132), .ZN(U282));
NOR3_X1 U1724 ( .A1(n2133), .A2(n2134), .A3(n2135), .ZN(n2132) );
NOR2_X1 U1725 ( .A1(n1938), .A2(n2136), .ZN(n2135) );
XOR2_X1 U1726 ( .A(n2137), .B(n2138), .Z(n2136) );
NAND2_X1 U1727 ( .A1(KEYINPUT45), .A2(n2107), .ZN(n2137) );
INV_X1 U1728 ( .A(n1945), .ZN(n1938) );
NOR2_X1 U1729 ( .A1(n1941), .A2(n2139), .ZN(n2134) );
XOR2_X1 U1730 ( .A(n2107), .B(n2115), .Z(n2139) );
NAND2_X1 U1731 ( .A1(n2052), .A2(n2140), .ZN(n2107) );
NAND2_X1 U1732 ( .A1(n2141), .A2(n2142), .ZN(n2140) );
NAND2_X1 U1733 ( .A1(n2143), .A2(n2144), .ZN(n2142) );
NAND3_X1 U1734 ( .A1(n2145), .A2(n2144), .A3(n2143), .ZN(n2052) );
NOR2_X1 U1735 ( .A1(n2145), .A2(n1976), .ZN(n2133) );
INV_X1 U1736 ( .A(n2141), .ZN(n2145) );
NAND2_X1 U1737 ( .A1(n2146), .A2(n2147), .ZN(n2141) );
NAND2_X1 U1738 ( .A1(n2148), .A2(n2149), .ZN(n2147) );
NAND2_X1 U1739 ( .A1(n2150), .A2(n2151), .ZN(n2148) );
NAND2_X1 U1740 ( .A1(KEYINPUT31), .A2(n2152), .ZN(n2151) );
NAND2_X1 U1741 ( .A1(n2125), .A2(n2153), .ZN(n2152) );
INV_X1 U1742 ( .A(KEYINPUT13), .ZN(n2153) );
XNOR2_X1 U1743 ( .A(n2125), .B(n2128), .ZN(n2150) );
NAND3_X1 U1744 ( .A1(n2154), .A2(n2155), .A3(n2127), .ZN(n2146) );
INV_X1 U1745 ( .A(n2149), .ZN(n2127) );
NAND2_X1 U1746 ( .A1(n2156), .A2(n2157), .ZN(n2149) );
NAND2_X1 U1747 ( .A1(n2158), .A2(n2159), .ZN(n2157) );
NAND2_X1 U1748 ( .A1(n2160), .A2(n2161), .ZN(n2159) );
XOR2_X1 U1749 ( .A(n2162), .B(KEYINPUT33), .Z(n2160) );
XOR2_X1 U1750 ( .A(KEYINPUT26), .B(n2163), .Z(n2158) );
XOR2_X1 U1751 ( .A(n2164), .B(KEYINPUT6), .Z(n2156) );
INV_X1 U1752 ( .A(KEYINPUT31), .ZN(n2155) );
XOR2_X1 U1753 ( .A(n2165), .B(n2125), .Z(n2154) );
NAND2_X1 U1754 ( .A1(n2166), .A2(n2167), .ZN(n2125) );
NAND2_X1 U1755 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1993), .ZN(n2167) );
NAND2_X1 U1756 ( .A1(RESTART), .A2(RMIN_REG_2__SCAN_IN), .ZN(n2166) );
NAND2_X1 U1757 ( .A1(KEYINPUT13), .A2(n2128), .ZN(n2165) );
NAND2_X1 U1758 ( .A1(n2168), .A2(n2169), .ZN(n2128) );
NAND2_X1 U1759 ( .A1(RESTART), .A2(n2170), .ZN(n2169) );
NAND2_X1 U1760 ( .A1(n1783), .A2(n1993), .ZN(n2168) );
INV_X1 U1761 ( .A(DATA_IN_2_), .ZN(n1783) );
NAND2_X1 U1762 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1854), .ZN(n2131) );
NAND2_X1 U1763 ( .A1(n1928), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2130) );
NAND2_X1 U1764 ( .A1(n1929), .A2(REG4_REG_1__SCAN_IN), .ZN(n2129) );
NAND4_X1 U1765 ( .A1(n2171), .A2(n2172), .A3(n2173), .A4(n2174), .ZN(U281));
NOR3_X1 U1766 ( .A1(n2175), .A2(n2176), .A3(n2177), .ZN(n2174) );
NOR2_X1 U1767 ( .A1(n2143), .A2(n1976), .ZN(n2177) );
NAND4_X1 U1768 ( .A1(U280), .A2(STATO_REG_1__SCAN_IN), .A3(n2178), .A4(n2179), .ZN(n1976) );
NAND2_X1 U1769 ( .A1(n2180), .A2(n1993), .ZN(n2179) );
NAND4_X1 U1770 ( .A1(ENABLE), .A2(n2181), .A3(n2182), .A4(n2183), .ZN(n2180));
NAND2_X1 U1771 ( .A1(KEYINPUT34), .A2(n2184), .ZN(n2181) );
NAND3_X1 U1772 ( .A1(n2184), .A2(n2185), .A3(RESTART), .ZN(n2178) );
INV_X1 U1773 ( .A(KEYINPUT34), .ZN(n2185) );
AND2_X1 U1774 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1928), .ZN(n2176) );
NOR2_X1 U1775 ( .A1(n2186), .A2(ENABLE), .ZN(n1928) );
AND2_X1 U1776 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1929), .ZN(n2175) );
NOR3_X1 U1777 ( .A1(n1851), .A2(n2186), .A3(n2183), .ZN(n1929) );
INV_X1 U1778 ( .A(AVERAGE), .ZN(n2183) );
NAND2_X1 U1779 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1854), .ZN(n2173) );
NAND2_X1 U1780 ( .A1(n2115), .A2(n1950), .ZN(n2172) );
INV_X1 U1781 ( .A(n1941), .ZN(n1950) );
NAND4_X1 U1782 ( .A1(RESTART), .A2(U280), .A3(STATO_REG_1__SCAN_IN), .A4(
n2184), .ZN(n1941) );
NAND2_X1 U1783 ( .A1(n2187), .A2(n2188), .ZN(n2184) );
NAND2_X1 U1784 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2188) );
NAND2_X1 U1785 ( .A1(n2189), .A2(n2190), .ZN(n2187) );
NAND2_X1 U1786 ( .A1(n2191), .A2(n2192), .ZN(n2190) );
NAND3_X1 U1787 ( .A1(n2193), .A2(n2194), .A3(n2195), .ZN(n2192) );
NAND2_X1 U1788 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n2196), .ZN(n2195) );
NAND2_X1 U1789 ( .A1(n2197), .A2(n2198), .ZN(n2194) );
NAND2_X1 U1790 ( .A1(n2199), .A2(n2200), .ZN(n2198) );
NAND3_X1 U1791 ( .A1(n2201), .A2(n2202), .A3(n2203), .ZN(n2200) );
OR2_X1 U1792 ( .A1(RMAX_REG_4__SCAN_IN), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2203) );
NAND3_X1 U1793 ( .A1(n2204), .A2(n2205), .A3(n2206), .ZN(n2202) );
NAND2_X1 U1794 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2206) );
NAND3_X1 U1795 ( .A1(n2207), .A2(n2208), .A3(n2209), .ZN(n2205) );
NAND2_X1 U1796 ( .A1(n2170), .A2(n1816), .ZN(n2209) );
INV_X1 U1797 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1816) );
INV_X1 U1798 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n2170) );
NAND2_X1 U1799 ( .A1(n2210), .A2(n2211), .ZN(n2208) );
NAND2_X1 U1800 ( .A1(n2212), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2210) );
OR2_X1 U1801 ( .A1(n2212), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2207) );
NOR2_X1 U1802 ( .A1(n2213), .A2(n2214), .ZN(n2212) );
NAND2_X1 U1803 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2204) );
NAND2_X1 U1804 ( .A1(n2122), .A2(n1828), .ZN(n2201) );
INV_X1 U1805 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1828) );
INV_X1 U1806 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n2122) );
NAND2_X1 U1807 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2199) );
XOR2_X1 U1808 ( .A(KEYINPUT53), .B(n2215), .Z(n2197) );
NOR2_X1 U1809 ( .A1(RMAX_REG_5__SCAN_IN), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2215) );
NAND2_X1 U1810 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n2216), .ZN(n2193) );
XOR2_X1 U1811 ( .A(RMAX_REG_5__SCAN_IN), .B(KEYINPUT12), .Z(n2216) );
OR2_X1 U1812 ( .A1(n2196), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2191) );
XNOR2_X1 U1813 ( .A(n1743), .B(KEYINPUT52), .ZN(n2196) );
INV_X1 U1814 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1743) );
NAND2_X1 U1815 ( .A1(n2217), .A2(n1795), .ZN(n2189) );
INV_X1 U1816 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1795) );
XNOR2_X1 U1817 ( .A(RMAX_REG_7__SCAN_IN), .B(KEYINPUT39), .ZN(n2217) );
XNOR2_X1 U1818 ( .A(n2143), .B(n2218), .ZN(n2115) );
NOR2_X1 U1819 ( .A1(KEYINPUT8), .A2(n2144), .ZN(n2218) );
NAND2_X1 U1820 ( .A1(n1945), .A2(n2103), .ZN(n2171) );
INV_X1 U1821 ( .A(n2138), .ZN(n2103) );
XNOR2_X1 U1822 ( .A(n2143), .B(n2144), .ZN(n2138) );
XNOR2_X1 U1823 ( .A(n2219), .B(n2220), .ZN(n2144) );
NOR2_X1 U1824 ( .A1(KEYINPUT62), .A2(n2221), .ZN(n2220) );
AND3_X1 U1825 ( .A1(n2222), .A2(n2223), .A3(n2224), .ZN(n2143) );
NAND3_X1 U1826 ( .A1(n2225), .A2(n2226), .A3(n2161), .ZN(n2224) );
NAND2_X1 U1827 ( .A1(n2227), .A2(n2228), .ZN(n2226) );
INV_X1 U1828 ( .A(KEYINPUT38), .ZN(n2228) );
XOR2_X1 U1829 ( .A(n2162), .B(n2163), .Z(n2227) );
NAND3_X1 U1830 ( .A1(n2163), .A2(n2162), .A3(KEYINPUT38), .ZN(n2225) );
NAND3_X1 U1831 ( .A1(n2229), .A2(n2162), .A3(n2230), .ZN(n2223) );
NAND2_X1 U1832 ( .A1(n2163), .A2(n2231), .ZN(n2222) );
XOR2_X1 U1833 ( .A(n2164), .B(KEYINPUT16), .Z(n2231) );
OR2_X1 U1834 ( .A1(n2162), .A2(n2161), .ZN(n2164) );
INV_X1 U1835 ( .A(n2229), .ZN(n2161) );
NAND3_X1 U1836 ( .A1(n2232), .A2(n2233), .A3(n2234), .ZN(n2229) );
OR2_X1 U1837 ( .A1(DATA_IN_1_), .A2(KEYINPUT37), .ZN(n2234) );
NAND3_X1 U1838 ( .A1(KEYINPUT37), .A2(DATA_IN_1_), .A3(n1993), .ZN(n2233) );
NAND2_X1 U1839 ( .A1(RESTART), .A2(n2235), .ZN(n2232) );
NAND2_X1 U1840 ( .A1(KEYINPUT37), .A2(n1786), .ZN(n2235) );
INV_X1 U1841 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1786) );
NAND2_X1 U1842 ( .A1(n2236), .A2(n2219), .ZN(n2162) );
NAND3_X1 U1843 ( .A1(n2237), .A2(n2238), .A3(n2239), .ZN(n2219) );
NAND2_X1 U1844 ( .A1(KEYINPUT58), .A2(n2214), .ZN(n2239) );
INV_X1 U1845 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n2214) );
NAND3_X1 U1846 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n2240), .A3(RESTART), .ZN(n2238) );
NAND2_X1 U1847 ( .A1(n2241), .A2(n1993), .ZN(n2237) );
NAND2_X1 U1848 ( .A1(n2240), .A2(n1784), .ZN(n2241) );
INV_X1 U1849 ( .A(DATA_IN_0_), .ZN(n1784) );
INV_X1 U1850 ( .A(KEYINPUT58), .ZN(n2240) );
XOR2_X1 U1851 ( .A(n2221), .B(KEYINPUT42), .Z(n2236) );
NAND2_X1 U1852 ( .A1(n2242), .A2(n2243), .ZN(n2221) );
NAND2_X1 U1853 ( .A1(RESTART), .A2(n2213), .ZN(n2243) );
INV_X1 U1854 ( .A(RMIN_REG_0__SCAN_IN), .ZN(n2213) );
OR2_X1 U1855 ( .A1(REG4_REG_0__SCAN_IN), .A2(RESTART), .ZN(n2242) );
INV_X1 U1856 ( .A(n2230), .ZN(n2163) );
NAND2_X1 U1857 ( .A1(n2244), .A2(n2245), .ZN(n2230) );
NAND2_X1 U1858 ( .A1(RESTART), .A2(n2211), .ZN(n2245) );
INV_X1 U1859 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n2211) );
NAND2_X1 U1860 ( .A1(n2246), .A2(n1993), .ZN(n2244) );
NOR4_X1 U1861 ( .A1(n1851), .A2(n2186), .A3(n2182), .A4(AVERAGE), .ZN(n1945));
NAND2_X1 U1862 ( .A1(n2247), .A2(n2248), .ZN(n2182) );
NAND2_X1 U1863 ( .A1(n2249), .A2(n2250), .ZN(n2248) );
INV_X1 U1864 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2250) );
OR2_X1 U1865 ( .A1(n2251), .A2(n1760), .ZN(n2249) );
NAND2_X1 U1866 ( .A1(n2251), .A2(n1760), .ZN(n2247) );
INV_X1 U1867 ( .A(DATA_IN_7_), .ZN(n1760) );
NAND2_X1 U1868 ( .A1(n2252), .A2(n2253), .ZN(n2251) );
NAND2_X1 U1869 ( .A1(DATA_IN_6_), .A2(n2254), .ZN(n2253) );
NAND2_X1 U1870 ( .A1(n2255), .A2(n1992), .ZN(n2254) );
INV_X1 U1871 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1992) );
XOR2_X1 U1872 ( .A(KEYINPUT21), .B(n2256), .Z(n2255) );
NAND2_X1 U1873 ( .A1(n2256), .A2(REG4_REG_6__SCAN_IN), .ZN(n2252) );
AND2_X1 U1874 ( .A1(n2257), .A2(n2258), .ZN(n2256) );
NAND2_X1 U1875 ( .A1(n2030), .A2(n2259), .ZN(n2258) );
NAND2_X1 U1876 ( .A1(DATA_IN_5_), .A2(n2260), .ZN(n2259) );
INV_X1 U1877 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2030) );
OR2_X1 U1878 ( .A1(n2260), .A2(DATA_IN_5_), .ZN(n2257) );
NAND2_X1 U1879 ( .A1(n2261), .A2(n2262), .ZN(n2260) );
NAND2_X1 U1880 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2262) );
NAND3_X1 U1881 ( .A1(n2263), .A2(n2264), .A3(n2265), .ZN(n2261) );
NAND2_X1 U1882 ( .A1(n1775), .A2(n2078), .ZN(n2265) );
INV_X1 U1883 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2078) );
INV_X1 U1884 ( .A(DATA_IN_4_), .ZN(n1775) );
NAND3_X1 U1885 ( .A1(n2266), .A2(n2267), .A3(n2268), .ZN(n2264) );
NAND2_X1 U1886 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2268) );
NAND3_X1 U1887 ( .A1(n2269), .A2(n2270), .A3(n2271), .ZN(n2267) );
OR2_X1 U1888 ( .A1(DATA_IN_2_), .A2(REG4_REG_2__SCAN_IN), .ZN(n2271) );
NAND2_X1 U1889 ( .A1(n2272), .A2(n2273), .ZN(n2270) );
NAND2_X1 U1890 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2273) );
NAND2_X1 U1891 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2272) );
NAND2_X1 U1892 ( .A1(n1787), .A2(n2246), .ZN(n2269) );
INV_X1 U1893 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2246) );
INV_X1 U1894 ( .A(DATA_IN_1_), .ZN(n1787) );
NAND2_X1 U1895 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2266) );
OR2_X1 U1896 ( .A1(DATA_IN_3_), .A2(REG4_REG_3__SCAN_IN), .ZN(n2263) );
NAND3_X1 U1897 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1993), .A3(U280), .ZN(n2186) );
INV_X1 U1898 ( .A(RESTART), .ZN(n1993) );
INV_X1 U1899 ( .A(ENABLE), .ZN(n1851) );
INV_X1 U1900 ( .A(n1854), .ZN(U280) );
NAND2_X1 U1901 ( .A1(STATO_REG_0__SCAN_IN), .A2(STATO_REG_1__SCAN_IN), .ZN(n2274) );
OR2_X1 U1902 ( .A1(STATO_REG_1__SCAN_IN), .A2(STATO_REG_0__SCAN_IN), .ZN(n1707) );
endmodule


