//Key = 0011100010100100011100101000111110011101001000001000101011000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;

XNOR2_X1 U698 ( .A(G107), .B(n946), .ZN(G9) );
NAND3_X1 U699 ( .A1(n947), .A2(n948), .A3(n949), .ZN(G75) );
NAND2_X1 U700 ( .A1(G952), .A2(n950), .ZN(n949) );
NAND2_X1 U701 ( .A1(n951), .A2(n952), .ZN(n950) );
NAND2_X1 U702 ( .A1(n953), .A2(n954), .ZN(n952) );
NAND2_X1 U703 ( .A1(n955), .A2(n956), .ZN(n953) );
NAND3_X1 U704 ( .A1(n957), .A2(n958), .A3(n959), .ZN(n956) );
NAND3_X1 U705 ( .A1(n960), .A2(n961), .A3(n962), .ZN(n958) );
NAND2_X1 U706 ( .A1(n963), .A2(n964), .ZN(n962) );
NAND2_X1 U707 ( .A1(n965), .A2(n966), .ZN(n964) );
NAND2_X1 U708 ( .A1(n967), .A2(n968), .ZN(n961) );
NAND2_X1 U709 ( .A1(n969), .A2(n970), .ZN(n968) );
NAND2_X1 U710 ( .A1(KEYINPUT42), .A2(n971), .ZN(n970) );
NAND2_X1 U711 ( .A1(n972), .A2(n973), .ZN(n969) );
OR3_X1 U712 ( .A1(n974), .A2(KEYINPUT42), .A3(n967), .ZN(n960) );
NAND4_X1 U713 ( .A1(n967), .A2(n963), .A3(n975), .A4(n976), .ZN(n955) );
NAND2_X1 U714 ( .A1(n959), .A2(n977), .ZN(n976) );
NAND2_X1 U715 ( .A1(n978), .A2(n979), .ZN(n977) );
NAND2_X1 U716 ( .A1(n980), .A2(n981), .ZN(n979) );
INV_X1 U717 ( .A(n957), .ZN(n978) );
NAND2_X1 U718 ( .A1(n982), .A2(n983), .ZN(n975) );
NAND2_X1 U719 ( .A1(n957), .A2(n984), .ZN(n982) );
NAND2_X1 U720 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND4_X1 U721 ( .A1(n987), .A2(n963), .A3(n988), .A4(n989), .ZN(n947) );
NOR4_X1 U722 ( .A1(n985), .A2(n990), .A3(n991), .A4(n992), .ZN(n989) );
XNOR2_X1 U723 ( .A(G478), .B(n993), .ZN(n991) );
NOR2_X1 U724 ( .A1(n994), .A2(KEYINPUT43), .ZN(n993) );
XNOR2_X1 U725 ( .A(n995), .B(n996), .ZN(n990) );
NOR2_X1 U726 ( .A1(KEYINPUT53), .A2(n997), .ZN(n996) );
XNOR2_X1 U727 ( .A(G469), .B(n998), .ZN(n988) );
NOR2_X1 U728 ( .A1(KEYINPUT1), .A2(n999), .ZN(n998) );
XOR2_X1 U729 ( .A(n1000), .B(n1001), .Z(G72) );
NOR2_X1 U730 ( .A1(n1002), .A2(n948), .ZN(n1001) );
NOR2_X1 U731 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NOR3_X1 U732 ( .A1(KEYINPUT33), .A2(n1005), .A3(n1006), .ZN(n1000) );
NOR2_X1 U733 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
XOR2_X1 U734 ( .A(KEYINPUT38), .B(n1009), .Z(n1008) );
AND2_X1 U735 ( .A1(n1007), .A2(n1009), .ZN(n1005) );
NOR2_X1 U736 ( .A1(G953), .A2(n1010), .ZN(n1009) );
AND2_X1 U737 ( .A1(n1011), .A2(n1012), .ZN(n1007) );
NAND2_X1 U738 ( .A1(G953), .A2(n1004), .ZN(n1012) );
XOR2_X1 U739 ( .A(n1013), .B(n1014), .Z(n1011) );
NOR2_X1 U740 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
XOR2_X1 U741 ( .A(n1017), .B(KEYINPUT10), .Z(n1016) );
NAND2_X1 U742 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
XNOR2_X1 U743 ( .A(G140), .B(KEYINPUT56), .ZN(n1018) );
NAND2_X1 U744 ( .A1(n1020), .A2(n1021), .ZN(G69) );
NAND2_X1 U745 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U746 ( .A1(G953), .A2(n1024), .ZN(n1023) );
NAND3_X1 U747 ( .A1(G953), .A2(n1025), .A3(n1026), .ZN(n1020) );
INV_X1 U748 ( .A(n1022), .ZN(n1026) );
XNOR2_X1 U749 ( .A(n1027), .B(n1028), .ZN(n1022) );
NOR3_X1 U750 ( .A1(n1029), .A2(KEYINPUT5), .A3(G953), .ZN(n1028) );
AND3_X1 U751 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
XNOR2_X1 U752 ( .A(n946), .B(KEYINPUT37), .ZN(n1032) );
NAND2_X1 U753 ( .A1(n1033), .A2(n1034), .ZN(n1027) );
NAND2_X1 U754 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U755 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
XNOR2_X1 U756 ( .A(KEYINPUT28), .B(n1039), .ZN(n1038) );
XNOR2_X1 U757 ( .A(n1040), .B(KEYINPUT50), .ZN(n1037) );
NAND2_X1 U758 ( .A1(n1041), .A2(n1040), .ZN(n1035) );
XOR2_X1 U759 ( .A(n1042), .B(n1043), .Z(n1040) );
XOR2_X1 U760 ( .A(KEYINPUT7), .B(n1044), .Z(n1043) );
XNOR2_X1 U761 ( .A(n1045), .B(KEYINPUT28), .ZN(n1041) );
NAND2_X1 U762 ( .A1(G953), .A2(n1046), .ZN(n1033) );
NAND2_X1 U763 ( .A1(G898), .A2(G224), .ZN(n1025) );
NOR2_X1 U764 ( .A1(n1047), .A2(n1048), .ZN(G66) );
XNOR2_X1 U765 ( .A(n1049), .B(n1050), .ZN(n1048) );
XOR2_X1 U766 ( .A(KEYINPUT0), .B(n1051), .Z(n1050) );
NOR2_X1 U767 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U768 ( .A1(n1047), .A2(n1054), .ZN(G63) );
XNOR2_X1 U769 ( .A(n1055), .B(n1056), .ZN(n1054) );
NOR2_X1 U770 ( .A1(n1057), .A2(n1053), .ZN(n1056) );
NOR2_X1 U771 ( .A1(n1047), .A2(n1058), .ZN(G60) );
XOR2_X1 U772 ( .A(n1059), .B(n1060), .Z(n1058) );
AND2_X1 U773 ( .A1(G475), .A2(n1061), .ZN(n1060) );
XOR2_X1 U774 ( .A(G104), .B(n1062), .Z(G6) );
NOR2_X1 U775 ( .A1(n1047), .A2(n1063), .ZN(G57) );
XOR2_X1 U776 ( .A(n1064), .B(n1065), .Z(n1063) );
XOR2_X1 U777 ( .A(n1066), .B(n1067), .Z(n1065) );
XNOR2_X1 U778 ( .A(G101), .B(n1068), .ZN(n1064) );
AND2_X1 U779 ( .A1(G472), .A2(n1061), .ZN(n1068) );
NOR2_X1 U780 ( .A1(n1047), .A2(n1069), .ZN(G54) );
NOR2_X1 U781 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U782 ( .A(KEYINPUT9), .B(n1072), .Z(n1071) );
NOR2_X1 U783 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
AND2_X1 U784 ( .A1(n1074), .A2(n1073), .ZN(n1070) );
XNOR2_X1 U785 ( .A(n1075), .B(n1076), .ZN(n1073) );
XOR2_X1 U786 ( .A(n1077), .B(n1078), .Z(n1075) );
NAND2_X1 U787 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NAND2_X1 U788 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U789 ( .A(KEYINPUT13), .B(n1083), .Z(n1079) );
NOR2_X1 U790 ( .A1(n1081), .A2(n1082), .ZN(n1083) );
NAND2_X1 U791 ( .A1(n1061), .A2(G469), .ZN(n1074) );
NOR2_X1 U792 ( .A1(n1047), .A2(n1084), .ZN(G51) );
XOR2_X1 U793 ( .A(n1085), .B(n1086), .Z(n1084) );
XOR2_X1 U794 ( .A(KEYINPUT3), .B(n1087), .Z(n1086) );
NOR2_X1 U795 ( .A1(n1088), .A2(n1053), .ZN(n1087) );
INV_X1 U796 ( .A(n1061), .ZN(n1053) );
NOR2_X1 U797 ( .A1(n1089), .A2(n951), .ZN(n1061) );
AND4_X1 U798 ( .A1(n1010), .A2(n1030), .A3(n1090), .A4(n946), .ZN(n951) );
NAND3_X1 U799 ( .A1(n1091), .A2(n957), .A3(n1092), .ZN(n946) );
XNOR2_X1 U800 ( .A(KEYINPUT22), .B(n1031), .ZN(n1090) );
NOR4_X1 U801 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1030) );
OR3_X1 U802 ( .A1(n1097), .A2(n1098), .A3(n1062), .ZN(n1096) );
AND3_X1 U803 ( .A1(n1092), .A2(n957), .A3(n1099), .ZN(n1062) );
INV_X1 U804 ( .A(n1100), .ZN(n1098) );
NOR4_X1 U805 ( .A1(n1101), .A2(n1102), .A3(n965), .A4(n980), .ZN(n1097) );
NOR2_X1 U806 ( .A1(KEYINPUT17), .A2(n1103), .ZN(n1102) );
NOR4_X1 U807 ( .A1(n1104), .A2(n974), .A3(n983), .A4(n1105), .ZN(n1103) );
INV_X1 U808 ( .A(n959), .ZN(n983) );
AND2_X1 U809 ( .A1(n1106), .A2(KEYINPUT17), .ZN(n1101) );
AND4_X1 U810 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1010) );
NOR4_X1 U811 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1110) );
NOR2_X1 U812 ( .A1(n974), .A2(n1115), .ZN(n1114) );
NOR3_X1 U813 ( .A1(n1116), .A2(n966), .A3(n1117), .ZN(n1113) );
AND2_X1 U814 ( .A1(n1118), .A2(n1119), .ZN(n1109) );
XNOR2_X1 U815 ( .A(n1120), .B(n1121), .ZN(n1085) );
NOR2_X1 U816 ( .A1(n948), .A2(G952), .ZN(n1047) );
XNOR2_X1 U817 ( .A(G146), .B(n1107), .ZN(G48) );
NAND3_X1 U818 ( .A1(n1099), .A2(n971), .A3(n1122), .ZN(n1107) );
XNOR2_X1 U819 ( .A(G143), .B(n1123), .ZN(G45) );
NAND2_X1 U820 ( .A1(n1124), .A2(n971), .ZN(n1123) );
XOR2_X1 U821 ( .A(n1115), .B(KEYINPUT18), .Z(n1124) );
OR3_X1 U822 ( .A1(n1125), .A2(n1126), .A3(n1116), .ZN(n1115) );
NAND2_X1 U823 ( .A1(n1127), .A2(n1128), .ZN(G42) );
NAND3_X1 U824 ( .A1(n1112), .A2(n1129), .A3(n1130), .ZN(n1128) );
INV_X1 U825 ( .A(n1131), .ZN(n1130) );
NAND2_X1 U826 ( .A1(n1131), .A2(n1132), .ZN(n1127) );
NAND2_X1 U827 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U828 ( .A1(n1112), .A2(n1135), .ZN(n1134) );
INV_X1 U829 ( .A(KEYINPUT8), .ZN(n1135) );
NAND2_X1 U830 ( .A1(KEYINPUT8), .A2(n1136), .ZN(n1133) );
NAND2_X1 U831 ( .A1(n1112), .A2(n1129), .ZN(n1136) );
INV_X1 U832 ( .A(KEYINPUT47), .ZN(n1129) );
AND3_X1 U833 ( .A1(n1137), .A2(n1099), .A3(n1138), .ZN(n1112) );
NOR3_X1 U834 ( .A1(n1117), .A2(n987), .A3(n981), .ZN(n1138) );
XOR2_X1 U835 ( .A(G140), .B(KEYINPUT16), .Z(n1131) );
XOR2_X1 U836 ( .A(n1111), .B(n1139), .Z(G39) );
NOR2_X1 U837 ( .A1(KEYINPUT61), .A2(n1140), .ZN(n1139) );
AND3_X1 U838 ( .A1(n1122), .A2(n963), .A3(n967), .ZN(n1111) );
XOR2_X1 U839 ( .A(G134), .B(n1141), .Z(G36) );
NOR3_X1 U840 ( .A1(n1116), .A2(n1142), .A3(n966), .ZN(n1141) );
XNOR2_X1 U841 ( .A(n963), .B(KEYINPUT34), .ZN(n1142) );
INV_X1 U842 ( .A(n1117), .ZN(n963) );
XNOR2_X1 U843 ( .A(G131), .B(n1119), .ZN(G33) );
OR3_X1 U844 ( .A1(n965), .A2(n1117), .A3(n1116), .ZN(n1119) );
NAND3_X1 U845 ( .A1(n987), .A2(n981), .A3(n1137), .ZN(n1116) );
NAND2_X1 U846 ( .A1(n973), .A2(n1143), .ZN(n1117) );
XNOR2_X1 U847 ( .A(G128), .B(n1118), .ZN(G30) );
NAND3_X1 U848 ( .A1(n1091), .A2(n971), .A3(n1122), .ZN(n1118) );
AND3_X1 U849 ( .A1(n980), .A2(n981), .A3(n1137), .ZN(n1122) );
NOR3_X1 U850 ( .A1(n1144), .A2(n985), .A3(n1145), .ZN(n1137) );
XNOR2_X1 U851 ( .A(n1146), .B(n1147), .ZN(G3) );
NOR2_X1 U852 ( .A1(KEYINPUT46), .A2(n1031), .ZN(n1147) );
NAND4_X1 U853 ( .A1(n967), .A2(n1092), .A3(n987), .A4(n981), .ZN(n1031) );
XOR2_X1 U854 ( .A(n1108), .B(n1148), .Z(G27) );
NAND2_X1 U855 ( .A1(KEYINPUT63), .A2(G125), .ZN(n1148) );
NAND4_X1 U856 ( .A1(n1104), .A2(n1099), .A3(n959), .A4(n1149), .ZN(n1108) );
NOR3_X1 U857 ( .A1(n974), .A2(n1144), .A3(n987), .ZN(n1149) );
AND2_X1 U858 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
NAND2_X1 U859 ( .A1(n1152), .A2(n1004), .ZN(n1151) );
INV_X1 U860 ( .A(G900), .ZN(n1004) );
INV_X1 U861 ( .A(n971), .ZN(n974) );
XNOR2_X1 U862 ( .A(G122), .B(n1100), .ZN(G24) );
NAND4_X1 U863 ( .A1(n1153), .A2(n1154), .A3(n957), .A4(n1155), .ZN(n1100) );
NOR2_X1 U864 ( .A1(n981), .A2(n980), .ZN(n957) );
XOR2_X1 U865 ( .A(G119), .B(n1095), .Z(G21) );
NOR3_X1 U866 ( .A1(n1156), .A2(n987), .A3(n1106), .ZN(n1095) );
INV_X1 U867 ( .A(n980), .ZN(n987) );
INV_X1 U868 ( .A(n967), .ZN(n1156) );
XNOR2_X1 U869 ( .A(G116), .B(n1157), .ZN(G18) );
NAND2_X1 U870 ( .A1(KEYINPUT52), .A2(n1093), .ZN(n1157) );
NOR3_X1 U871 ( .A1(n980), .A2(n966), .A3(n1106), .ZN(n1093) );
INV_X1 U872 ( .A(n1091), .ZN(n966) );
NOR2_X1 U873 ( .A1(n1153), .A2(n1126), .ZN(n1091) );
INV_X1 U874 ( .A(n1155), .ZN(n1126) );
XNOR2_X1 U875 ( .A(n1158), .B(n1159), .ZN(G15) );
NOR3_X1 U876 ( .A1(n1106), .A2(n965), .A3(n980), .ZN(n1159) );
INV_X1 U877 ( .A(n1099), .ZN(n965) );
NOR2_X1 U878 ( .A1(n1155), .A2(n1125), .ZN(n1099) );
NAND2_X1 U879 ( .A1(n1154), .A2(n981), .ZN(n1106) );
AND3_X1 U880 ( .A1(n971), .A2(n1105), .A3(n959), .ZN(n1154) );
NOR2_X1 U881 ( .A1(n986), .A2(n985), .ZN(n959) );
INV_X1 U882 ( .A(n1160), .ZN(n985) );
XOR2_X1 U883 ( .A(G110), .B(n1094), .Z(G12) );
AND4_X1 U884 ( .A1(n967), .A2(n1092), .A3(n1104), .A4(n980), .ZN(n1094) );
XOR2_X1 U885 ( .A(n1161), .B(n1052), .Z(n980) );
NAND2_X1 U886 ( .A1(G217), .A2(n1162), .ZN(n1052) );
NAND2_X1 U887 ( .A1(n1049), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U888 ( .A(n1164), .B(n1165), .ZN(n1049) );
XOR2_X1 U889 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U890 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U891 ( .A1(KEYINPUT59), .A2(n1170), .ZN(n1168) );
XOR2_X1 U892 ( .A(n1078), .B(n1171), .Z(n1170) );
XNOR2_X1 U893 ( .A(n1172), .B(G119), .ZN(n1171) );
INV_X1 U894 ( .A(G128), .ZN(n1172) );
NOR3_X1 U895 ( .A1(n1173), .A2(KEYINPUT40), .A3(n1174), .ZN(n1166) );
INV_X1 U896 ( .A(G221), .ZN(n1174) );
XNOR2_X1 U897 ( .A(G137), .B(n1175), .ZN(n1164) );
XOR2_X1 U898 ( .A(KEYINPUT62), .B(G146), .Z(n1175) );
INV_X1 U899 ( .A(n981), .ZN(n1104) );
XOR2_X1 U900 ( .A(n992), .B(KEYINPUT51), .Z(n981) );
XNOR2_X1 U901 ( .A(n1176), .B(G472), .ZN(n992) );
NAND2_X1 U902 ( .A1(n1177), .A2(n1163), .ZN(n1176) );
XOR2_X1 U903 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U904 ( .A(n1067), .B(n1180), .Z(n1179) );
NOR2_X1 U905 ( .A1(G101), .A2(KEYINPUT27), .ZN(n1180) );
XOR2_X1 U906 ( .A(n1181), .B(n1014), .Z(n1067) );
XNOR2_X1 U907 ( .A(n1182), .B(n1183), .ZN(n1014) );
INV_X1 U908 ( .A(n1082), .ZN(n1182) );
NAND2_X1 U909 ( .A1(n1184), .A2(G210), .ZN(n1181) );
XOR2_X1 U910 ( .A(n1185), .B(n1186), .Z(n1178) );
NOR2_X1 U911 ( .A1(KEYINPUT55), .A2(n1066), .ZN(n1186) );
XNOR2_X1 U912 ( .A(KEYINPUT57), .B(KEYINPUT14), .ZN(n1185) );
AND4_X1 U913 ( .A1(n986), .A2(n971), .A3(n1105), .A4(n1160), .ZN(n1092) );
NAND2_X1 U914 ( .A1(G221), .A2(n1162), .ZN(n1160) );
NAND2_X1 U915 ( .A1(G234), .A2(n1089), .ZN(n1162) );
NAND2_X1 U916 ( .A1(n1150), .A2(n1187), .ZN(n1105) );
NAND2_X1 U917 ( .A1(n1152), .A2(n1046), .ZN(n1187) );
INV_X1 U918 ( .A(G898), .ZN(n1046) );
AND3_X1 U919 ( .A1(G902), .A2(n954), .A3(G953), .ZN(n1152) );
NAND3_X1 U920 ( .A1(G952), .A2(n948), .A3(n1188), .ZN(n1150) );
XOR2_X1 U921 ( .A(n954), .B(KEYINPUT49), .Z(n1188) );
NAND2_X1 U922 ( .A1(G237), .A2(G234), .ZN(n954) );
NOR2_X1 U923 ( .A1(n973), .A2(n972), .ZN(n971) );
INV_X1 U924 ( .A(n1143), .ZN(n972) );
NAND2_X1 U925 ( .A1(G214), .A2(n1189), .ZN(n1143) );
XNOR2_X1 U926 ( .A(n1190), .B(n1088), .ZN(n973) );
NAND2_X1 U927 ( .A1(G210), .A2(n1189), .ZN(n1088) );
NAND2_X1 U928 ( .A1(n1191), .A2(n1089), .ZN(n1189) );
INV_X1 U929 ( .A(G237), .ZN(n1191) );
NAND2_X1 U930 ( .A1(n1192), .A2(n1163), .ZN(n1190) );
XOR2_X1 U931 ( .A(n1193), .B(n1121), .Z(n1192) );
XNOR2_X1 U932 ( .A(n1194), .B(n1195), .ZN(n1121) );
XOR2_X1 U933 ( .A(n1044), .B(n1196), .Z(n1195) );
NOR2_X1 U934 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U935 ( .A1(KEYINPUT39), .A2(n1042), .ZN(n1198) );
AND2_X1 U936 ( .A1(KEYINPUT32), .A2(n1042), .ZN(n1197) );
XNOR2_X1 U937 ( .A(n1066), .B(KEYINPUT45), .ZN(n1042) );
XNOR2_X1 U938 ( .A(G113), .B(n1199), .ZN(n1066) );
XNOR2_X1 U939 ( .A(G119), .B(n1200), .ZN(n1199) );
INV_X1 U940 ( .A(G116), .ZN(n1200) );
XNOR2_X1 U941 ( .A(n1146), .B(n1201), .ZN(n1044) );
NOR2_X1 U942 ( .A1(KEYINPUT25), .A2(n1202), .ZN(n1201) );
XOR2_X1 U943 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U944 ( .A(KEYINPUT24), .B(KEYINPUT11), .Z(n1204) );
XNOR2_X1 U945 ( .A(n1205), .B(n1039), .ZN(n1194) );
INV_X1 U946 ( .A(n1045), .ZN(n1039) );
XOR2_X1 U947 ( .A(G122), .B(n1078), .Z(n1045) );
XNOR2_X1 U948 ( .A(n1183), .B(n1206), .ZN(n1205) );
NOR2_X1 U949 ( .A1(n1024), .A2(n1207), .ZN(n1206) );
XNOR2_X1 U950 ( .A(KEYINPUT15), .B(n948), .ZN(n1207) );
INV_X1 U951 ( .A(G224), .ZN(n1024) );
NOR2_X1 U952 ( .A1(KEYINPUT20), .A2(n1120), .ZN(n1193) );
INV_X1 U953 ( .A(n1145), .ZN(n986) );
XOR2_X1 U954 ( .A(G469), .B(n1208), .Z(n1145) );
NOR2_X1 U955 ( .A1(n1209), .A2(KEYINPUT44), .ZN(n1208) );
INV_X1 U956 ( .A(n999), .ZN(n1209) );
NAND2_X1 U957 ( .A1(n1210), .A2(n1163), .ZN(n999) );
XOR2_X1 U958 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U959 ( .A(n1213), .B(n1076), .Z(n1212) );
XNOR2_X1 U960 ( .A(n1214), .B(n1215), .ZN(n1076) );
NOR2_X1 U961 ( .A1(G953), .A2(n1003), .ZN(n1215) );
INV_X1 U962 ( .A(G227), .ZN(n1003) );
NAND2_X1 U963 ( .A1(n1216), .A2(n1217), .ZN(n1213) );
NAND2_X1 U964 ( .A1(KEYINPUT36), .A2(n1081), .ZN(n1217) );
XOR2_X1 U965 ( .A(n1218), .B(n1183), .Z(n1081) );
OR3_X1 U966 ( .A1(n1218), .A2(n1183), .A3(KEYINPUT36), .ZN(n1216) );
XOR2_X1 U967 ( .A(G128), .B(n1219), .Z(n1183) );
XNOR2_X1 U968 ( .A(n1203), .B(n1146), .ZN(n1218) );
INV_X1 U969 ( .A(G101), .ZN(n1146) );
XNOR2_X1 U970 ( .A(G107), .B(n1220), .ZN(n1203) );
XNOR2_X1 U971 ( .A(n1082), .B(n1221), .ZN(n1211) );
XNOR2_X1 U972 ( .A(n1222), .B(KEYINPUT54), .ZN(n1221) );
NAND2_X1 U973 ( .A1(KEYINPUT31), .A2(n1078), .ZN(n1222) );
XOR2_X1 U974 ( .A(G110), .B(KEYINPUT60), .Z(n1078) );
XOR2_X1 U975 ( .A(G131), .B(n1223), .Z(n1082) );
XNOR2_X1 U976 ( .A(n1140), .B(G134), .ZN(n1223) );
INV_X1 U977 ( .A(G137), .ZN(n1140) );
NOR2_X1 U978 ( .A1(n1155), .A2(n1153), .ZN(n967) );
INV_X1 U979 ( .A(n1125), .ZN(n1153) );
XOR2_X1 U980 ( .A(n1224), .B(n997), .Z(n1125) );
XNOR2_X1 U981 ( .A(G475), .B(KEYINPUT35), .ZN(n997) );
XNOR2_X1 U982 ( .A(KEYINPUT2), .B(n1225), .ZN(n1224) );
NOR2_X1 U983 ( .A1(n995), .A2(KEYINPUT26), .ZN(n1225) );
AND2_X1 U984 ( .A1(n1226), .A2(n1163), .ZN(n995) );
XOR2_X1 U985 ( .A(n1059), .B(KEYINPUT4), .Z(n1226) );
XOR2_X1 U986 ( .A(n1227), .B(n1228), .Z(n1059) );
XNOR2_X1 U987 ( .A(n1158), .B(n1229), .ZN(n1228) );
XNOR2_X1 U988 ( .A(KEYINPUT30), .B(n1230), .ZN(n1229) );
INV_X1 U989 ( .A(G113), .ZN(n1158) );
XNOR2_X1 U990 ( .A(n1220), .B(n1231), .ZN(n1227) );
NOR2_X1 U991 ( .A1(KEYINPUT6), .A2(n1232), .ZN(n1231) );
XOR2_X1 U992 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U993 ( .A(n1169), .B(n1219), .ZN(n1234) );
XOR2_X1 U994 ( .A(G143), .B(G146), .Z(n1219) );
NOR2_X1 U995 ( .A1(n1015), .A2(n1235), .ZN(n1169) );
NOR2_X1 U996 ( .A1(n1214), .A2(n1120), .ZN(n1235) );
INV_X1 U997 ( .A(G140), .ZN(n1214) );
NOR2_X1 U998 ( .A1(n1019), .A2(G140), .ZN(n1015) );
INV_X1 U999 ( .A(n1120), .ZN(n1019) );
XOR2_X1 U1000 ( .A(G125), .B(KEYINPUT41), .Z(n1120) );
XOR2_X1 U1001 ( .A(n1236), .B(G131), .Z(n1233) );
NAND2_X1 U1002 ( .A1(n1184), .A2(G214), .ZN(n1236) );
NOR2_X1 U1003 ( .A1(G953), .A2(G237), .ZN(n1184) );
XOR2_X1 U1004 ( .A(G104), .B(KEYINPUT48), .Z(n1220) );
XOR2_X1 U1005 ( .A(n994), .B(n1237), .Z(n1155) );
XNOR2_X1 U1006 ( .A(KEYINPUT58), .B(n1057), .ZN(n1237) );
INV_X1 U1007 ( .A(G478), .ZN(n1057) );
AND2_X1 U1008 ( .A1(n1055), .A2(n1163), .ZN(n994) );
XNOR2_X1 U1009 ( .A(n1089), .B(KEYINPUT29), .ZN(n1163) );
INV_X1 U1010 ( .A(G902), .ZN(n1089) );
XNOR2_X1 U1011 ( .A(n1238), .B(n1239), .ZN(n1055) );
XOR2_X1 U1012 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U1013 ( .A(n1242), .B(n1243), .ZN(n1241) );
NOR2_X1 U1014 ( .A1(KEYINPUT23), .A2(n1244), .ZN(n1243) );
XOR2_X1 U1015 ( .A(KEYINPUT12), .B(G107), .Z(n1244) );
NAND2_X1 U1016 ( .A1(KEYINPUT19), .A2(n1230), .ZN(n1242) );
INV_X1 U1017 ( .A(G122), .ZN(n1230) );
NOR2_X1 U1018 ( .A1(n1173), .A2(n1245), .ZN(n1240) );
INV_X1 U1019 ( .A(G217), .ZN(n1245) );
NAND2_X1 U1020 ( .A1(G234), .A2(n948), .ZN(n1173) );
INV_X1 U1021 ( .A(G953), .ZN(n948) );
XOR2_X1 U1022 ( .A(n1246), .B(n1247), .Z(n1238) );
NOR2_X1 U1023 ( .A1(KEYINPUT21), .A2(n1248), .ZN(n1247) );
XNOR2_X1 U1024 ( .A(G143), .B(G128), .ZN(n1248) );
XNOR2_X1 U1025 ( .A(G116), .B(G134), .ZN(n1246) );
endmodule


