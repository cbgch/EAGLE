//Key = 1010001110001000110111001101101101010101011100111110101101011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338;

XNOR2_X1 U746 ( .A(G107), .B(n1025), .ZN(G9) );
NAND2_X1 U747 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U748 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U749 ( .A1(G953), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
NOR2_X1 U750 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U751 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U752 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U753 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U754 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR3_X1 U755 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1041) );
NOR3_X1 U756 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
XNOR2_X1 U757 ( .A(KEYINPUT24), .B(n1049), .ZN(n1048) );
INV_X1 U758 ( .A(n1050), .ZN(n1047) );
NOR3_X1 U759 ( .A1(n1051), .A2(n1049), .A3(n1050), .ZN(n1044) );
NOR2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1043) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR3_X1 U763 ( .A1(n1049), .A2(n1058), .A3(n1053), .ZN(n1039) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR4_X1 U765 ( .A1(n1061), .A2(n1042), .A3(n1053), .A4(n1049), .ZN(n1035) );
NOR2_X1 U766 ( .A1(n1026), .A2(n1062), .ZN(n1061) );
NOR3_X1 U767 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n1028) );
AND4_X1 U768 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1030) );
NOR4_X1 U769 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
XOR2_X1 U770 ( .A(n1071), .B(n1072), .Z(n1069) );
NOR2_X1 U771 ( .A1(KEYINPUT38), .A2(n1073), .ZN(n1072) );
INV_X1 U772 ( .A(G475), .ZN(n1073) );
XNOR2_X1 U773 ( .A(n1074), .B(KEYINPUT12), .ZN(n1071) );
XOR2_X1 U774 ( .A(n1075), .B(n1076), .Z(n1068) );
XOR2_X1 U775 ( .A(KEYINPUT27), .B(G472), .Z(n1076) );
XOR2_X1 U776 ( .A(n1077), .B(n1078), .Z(n1065) );
XOR2_X1 U777 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n1078) );
XOR2_X1 U778 ( .A(n1079), .B(n1080), .Z(n1077) );
XOR2_X1 U779 ( .A(n1081), .B(n1082), .Z(G72) );
NOR3_X1 U780 ( .A1(n1083), .A2(KEYINPUT62), .A3(n1084), .ZN(n1082) );
AND2_X1 U781 ( .A1(G227), .A2(G900), .ZN(n1084) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
NAND2_X1 U783 ( .A1(n1087), .A2(n1083), .ZN(n1086) );
XOR2_X1 U784 ( .A(n1088), .B(n1089), .Z(n1087) );
OR3_X1 U785 ( .A1(n1090), .A2(n1089), .A3(n1083), .ZN(n1085) );
XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(n1089) );
NOR2_X1 U787 ( .A1(KEYINPUT26), .A2(n1093), .ZN(n1092) );
XOR2_X1 U788 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U789 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U790 ( .A1(KEYINPUT6), .A2(n1098), .ZN(n1096) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(n1094) );
NAND2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(G69) );
NAND2_X1 U793 ( .A1(n1103), .A2(n1083), .ZN(n1102) );
XNOR2_X1 U794 ( .A(n1104), .B(n1105), .ZN(n1103) );
NAND2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
XNOR2_X1 U796 ( .A(n1108), .B(KEYINPUT49), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1109), .A2(G953), .ZN(n1101) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1105), .A2(n1112), .ZN(n1111) );
INV_X1 U800 ( .A(G224), .ZN(n1112) );
NAND2_X1 U801 ( .A1(G224), .A2(n1113), .ZN(n1110) );
NAND2_X1 U802 ( .A1(G898), .A2(n1105), .ZN(n1113) );
NAND2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(n1105) );
NAND2_X1 U804 ( .A1(G953), .A2(n1116), .ZN(n1115) );
XOR2_X1 U805 ( .A(n1117), .B(n1118), .Z(n1114) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XOR2_X1 U808 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U809 ( .A1(KEYINPUT22), .A2(n1125), .ZN(n1124) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1123) );
NOR2_X1 U811 ( .A1(n1121), .A2(n1128), .ZN(G63) );
XOR2_X1 U812 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U813 ( .A1(n1131), .A2(G478), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1121), .A2(n1132), .ZN(G60) );
NOR3_X1 U815 ( .A1(n1074), .A2(n1133), .A3(n1134), .ZN(n1132) );
AND3_X1 U816 ( .A1(n1135), .A2(G475), .A3(n1131), .ZN(n1134) );
NOR2_X1 U817 ( .A1(n1136), .A2(n1135), .ZN(n1133) );
AND2_X1 U818 ( .A1(n1032), .A2(G475), .ZN(n1136) );
XNOR2_X1 U819 ( .A(G104), .B(n1137), .ZN(G6) );
NOR2_X1 U820 ( .A1(n1138), .A2(n1139), .ZN(G57) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U822 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U823 ( .A(n1144), .B(n1145), .Z(n1142) );
NAND3_X1 U824 ( .A1(n1131), .A2(G472), .A3(KEYINPUT54), .ZN(n1144) );
XOR2_X1 U825 ( .A(n1146), .B(n1147), .Z(n1140) );
XOR2_X1 U826 ( .A(KEYINPUT3), .B(G101), .Z(n1147) );
NOR2_X1 U827 ( .A1(n1148), .A2(n1083), .ZN(n1138) );
XNOR2_X1 U828 ( .A(G952), .B(KEYINPUT57), .ZN(n1148) );
NOR2_X1 U829 ( .A1(n1121), .A2(n1149), .ZN(G54) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1149) );
XNOR2_X1 U831 ( .A(n1152), .B(n1153), .ZN(n1151) );
NAND2_X1 U832 ( .A1(n1154), .A2(KEYINPUT50), .ZN(n1152) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1150) );
NOR2_X1 U835 ( .A1(KEYINPUT34), .A2(n1159), .ZN(n1158) );
NAND2_X1 U836 ( .A1(n1131), .A2(G469), .ZN(n1157) );
NOR2_X1 U837 ( .A1(n1121), .A2(n1160), .ZN(G51) );
XOR2_X1 U838 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U839 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND3_X1 U840 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1164) );
NAND2_X1 U841 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U842 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
INV_X1 U843 ( .A(KEYINPUT8), .ZN(n1171) );
NAND2_X1 U844 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
XOR2_X1 U845 ( .A(KEYINPUT37), .B(n1169), .Z(n1172) );
NAND2_X1 U846 ( .A1(KEYINPUT8), .A2(n1174), .ZN(n1165) );
NAND2_X1 U847 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
OR2_X1 U848 ( .A1(G125), .A2(KEYINPUT37), .ZN(n1176) );
NAND3_X1 U849 ( .A1(G125), .A2(n1173), .A3(KEYINPUT37), .ZN(n1175) );
XOR2_X1 U850 ( .A(n1177), .B(n1178), .Z(n1161) );
NOR2_X1 U851 ( .A1(KEYINPUT29), .A2(n1179), .ZN(n1178) );
NAND2_X1 U852 ( .A1(n1131), .A2(n1080), .ZN(n1177) );
INV_X1 U853 ( .A(n1127), .ZN(n1131) );
NAND2_X1 U854 ( .A1(G902), .A2(n1032), .ZN(n1127) );
NAND3_X1 U855 ( .A1(n1107), .A2(n1088), .A3(n1108), .ZN(n1032) );
AND3_X1 U856 ( .A1(n1137), .A2(n1180), .A3(n1181), .ZN(n1108) );
NAND2_X1 U857 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U858 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U859 ( .A1(n1186), .A2(n1026), .ZN(n1185) );
XOR2_X1 U860 ( .A(n1042), .B(KEYINPUT31), .Z(n1186) );
NAND2_X1 U861 ( .A1(n1059), .A2(n1187), .ZN(n1184) );
NAND2_X1 U862 ( .A1(n1062), .A2(n1027), .ZN(n1137) );
NOR2_X1 U863 ( .A1(n1188), .A2(n1042), .ZN(n1027) );
AND4_X1 U864 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1088) );
AND4_X1 U865 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
AND2_X1 U866 ( .A1(n1197), .A2(n1198), .ZN(n1191) );
NAND3_X1 U867 ( .A1(n1199), .A2(n1060), .A3(n1200), .ZN(n1190) );
XNOR2_X1 U868 ( .A(n1062), .B(KEYINPUT42), .ZN(n1200) );
NAND2_X1 U869 ( .A1(n1201), .A2(n1055), .ZN(n1189) );
XOR2_X1 U870 ( .A(n1202), .B(KEYINPUT43), .Z(n1201) );
AND4_X1 U871 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1107) );
NAND3_X1 U872 ( .A1(n1207), .A2(n1062), .A3(n1208), .ZN(n1203) );
XOR2_X1 U873 ( .A(n1209), .B(KEYINPUT16), .Z(n1208) );
NOR2_X1 U874 ( .A1(n1083), .A2(G952), .ZN(n1121) );
XOR2_X1 U875 ( .A(G146), .B(n1210), .Z(G48) );
NOR2_X1 U876 ( .A1(n1211), .A2(n1202), .ZN(n1210) );
NAND3_X1 U877 ( .A1(n1212), .A2(n1062), .A3(n1213), .ZN(n1202) );
XOR2_X1 U878 ( .A(n1214), .B(n1197), .Z(G45) );
NAND4_X1 U879 ( .A1(n1215), .A2(n1216), .A3(n1055), .A4(n1217), .ZN(n1197) );
NOR2_X1 U880 ( .A1(n1209), .A2(n1218), .ZN(n1217) );
XOR2_X1 U881 ( .A(G140), .B(n1219), .Z(G42) );
NOR2_X1 U882 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
AND2_X1 U883 ( .A1(KEYINPUT21), .A2(n1222), .ZN(n1221) );
NAND2_X1 U884 ( .A1(n1199), .A2(n1223), .ZN(n1222) );
NOR3_X1 U885 ( .A1(n1224), .A2(KEYINPUT59), .A3(n1225), .ZN(n1220) );
INV_X1 U886 ( .A(n1199), .ZN(n1224) );
XNOR2_X1 U887 ( .A(G137), .B(n1196), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1212), .A2(n1187), .A3(n1199), .ZN(n1196) );
XNOR2_X1 U889 ( .A(G134), .B(n1195), .ZN(G36) );
NAND3_X1 U890 ( .A1(n1059), .A2(n1026), .A3(n1199), .ZN(n1195) );
XOR2_X1 U891 ( .A(n1098), .B(n1194), .Z(G33) );
NAND3_X1 U892 ( .A1(n1059), .A2(n1062), .A3(n1199), .ZN(n1194) );
NOR2_X1 U893 ( .A1(n1218), .A2(n1049), .ZN(n1199) );
OR2_X1 U894 ( .A1(n1056), .A2(n1067), .ZN(n1049) );
INV_X1 U895 ( .A(n1057), .ZN(n1067) );
XOR2_X1 U896 ( .A(n1099), .B(n1198), .Z(G30) );
NAND4_X1 U897 ( .A1(n1213), .A2(n1212), .A3(n1026), .A4(n1055), .ZN(n1198) );
INV_X1 U898 ( .A(n1218), .ZN(n1213) );
NAND3_X1 U899 ( .A1(n1050), .A2(n1226), .A3(n1051), .ZN(n1218) );
XOR2_X1 U900 ( .A(G101), .B(n1227), .Z(G3) );
NOR4_X1 U901 ( .A1(KEYINPUT51), .A2(n1188), .A3(n1038), .A4(n1209), .ZN(n1227) );
XOR2_X1 U902 ( .A(n1169), .B(n1193), .Z(G27) );
NAND4_X1 U903 ( .A1(n1223), .A2(n1064), .A3(n1055), .A4(n1226), .ZN(n1193) );
NAND2_X1 U904 ( .A1(n1228), .A2(n1034), .ZN(n1226) );
NAND2_X1 U905 ( .A1(n1090), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U906 ( .A(G900), .B(KEYINPUT1), .ZN(n1090) );
INV_X1 U907 ( .A(n1225), .ZN(n1223) );
NAND2_X1 U908 ( .A1(n1062), .A2(n1060), .ZN(n1225) );
INV_X1 U909 ( .A(G125), .ZN(n1169) );
XNOR2_X1 U910 ( .A(G122), .B(n1204), .ZN(G24) );
NAND4_X1 U911 ( .A1(n1207), .A2(n1230), .A3(n1215), .A4(n1216), .ZN(n1204) );
INV_X1 U912 ( .A(n1042), .ZN(n1230) );
NAND2_X1 U913 ( .A1(n1063), .A2(n1231), .ZN(n1042) );
XNOR2_X1 U914 ( .A(G119), .B(n1205), .ZN(G21) );
NAND3_X1 U915 ( .A1(n1207), .A2(n1187), .A3(n1212), .ZN(n1205) );
NOR2_X1 U916 ( .A1(n1231), .A2(n1063), .ZN(n1212) );
NAND2_X1 U917 ( .A1(n1232), .A2(n1233), .ZN(G18) );
OR2_X1 U918 ( .A1(n1206), .A2(G116), .ZN(n1233) );
XOR2_X1 U919 ( .A(n1234), .B(KEYINPUT23), .Z(n1232) );
NAND2_X1 U920 ( .A1(G116), .A2(n1206), .ZN(n1234) );
NAND3_X1 U921 ( .A1(n1059), .A2(n1026), .A3(n1207), .ZN(n1206) );
AND2_X1 U922 ( .A1(n1235), .A2(n1215), .ZN(n1026) );
XOR2_X1 U923 ( .A(n1070), .B(KEYINPUT10), .Z(n1215) );
XOR2_X1 U924 ( .A(n1236), .B(n1237), .Z(G15) );
AND3_X1 U925 ( .A1(n1207), .A2(n1062), .A3(n1059), .ZN(n1237) );
INV_X1 U926 ( .A(n1209), .ZN(n1059) );
NAND2_X1 U927 ( .A1(n1063), .A2(n1238), .ZN(n1209) );
NOR2_X1 U928 ( .A1(n1070), .A2(n1235), .ZN(n1062) );
INV_X1 U929 ( .A(n1239), .ZN(n1070) );
AND2_X1 U930 ( .A1(n1064), .A2(n1240), .ZN(n1207) );
INV_X1 U931 ( .A(n1053), .ZN(n1064) );
NAND2_X1 U932 ( .A1(n1046), .A2(n1050), .ZN(n1053) );
NOR2_X1 U933 ( .A1(KEYINPUT56), .A2(n1241), .ZN(n1236) );
XOR2_X1 U934 ( .A(KEYINPUT46), .B(G113), .Z(n1241) );
XOR2_X1 U935 ( .A(n1156), .B(n1180), .Z(G12) );
NAND3_X1 U936 ( .A1(n1060), .A2(n1182), .A3(n1187), .ZN(n1180) );
INV_X1 U937 ( .A(n1038), .ZN(n1187) );
NAND2_X1 U938 ( .A1(n1235), .A2(n1239), .ZN(n1038) );
XOR2_X1 U939 ( .A(n1242), .B(G478), .Z(n1239) );
NAND2_X1 U940 ( .A1(n1130), .A2(n1243), .ZN(n1242) );
XOR2_X1 U941 ( .A(n1244), .B(n1245), .Z(n1130) );
XOR2_X1 U942 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U943 ( .A(n1248), .B(n1249), .Z(n1244) );
XOR2_X1 U944 ( .A(n1250), .B(G116), .Z(n1248) );
NAND2_X1 U945 ( .A1(G217), .A2(n1251), .ZN(n1250) );
INV_X1 U946 ( .A(n1216), .ZN(n1235) );
XOR2_X1 U947 ( .A(n1074), .B(G475), .Z(n1216) );
NOR2_X1 U948 ( .A1(n1135), .A2(G902), .ZN(n1074) );
XNOR2_X1 U949 ( .A(n1252), .B(KEYINPUT25), .ZN(n1135) );
XOR2_X1 U950 ( .A(n1253), .B(n1254), .Z(n1252) );
XOR2_X1 U951 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U952 ( .A(G131), .B(G113), .Z(n1256) );
XOR2_X1 U953 ( .A(KEYINPUT20), .B(G146), .Z(n1255) );
XOR2_X1 U954 ( .A(n1257), .B(n1258), .Z(n1253) );
XOR2_X1 U955 ( .A(n1259), .B(n1247), .Z(n1258) );
XOR2_X1 U956 ( .A(G122), .B(G143), .Z(n1247) );
XOR2_X1 U957 ( .A(n1260), .B(n1091), .Z(n1257) );
NAND3_X1 U958 ( .A1(n1261), .A2(n1083), .A3(G214), .ZN(n1260) );
INV_X1 U959 ( .A(n1188), .ZN(n1182) );
NAND3_X1 U960 ( .A1(n1051), .A2(n1050), .A3(n1240), .ZN(n1188) );
AND2_X1 U961 ( .A1(n1055), .A2(n1262), .ZN(n1240) );
NAND2_X1 U962 ( .A1(n1034), .A2(n1263), .ZN(n1262) );
NAND2_X1 U963 ( .A1(n1229), .A2(n1116), .ZN(n1263) );
INV_X1 U964 ( .A(G898), .ZN(n1116) );
AND3_X1 U965 ( .A1(G902), .A2(n1264), .A3(G953), .ZN(n1229) );
NAND3_X1 U966 ( .A1(n1264), .A2(n1083), .A3(G952), .ZN(n1034) );
NAND2_X1 U967 ( .A1(G237), .A2(G234), .ZN(n1264) );
INV_X1 U968 ( .A(n1211), .ZN(n1055) );
NAND2_X1 U969 ( .A1(n1056), .A2(n1057), .ZN(n1211) );
NAND2_X1 U970 ( .A1(G214), .A2(n1265), .ZN(n1057) );
XOR2_X1 U971 ( .A(n1266), .B(n1267), .Z(n1056) );
XOR2_X1 U972 ( .A(KEYINPUT9), .B(n1080), .Z(n1267) );
AND2_X1 U973 ( .A1(G210), .A2(n1265), .ZN(n1080) );
NAND2_X1 U974 ( .A1(n1261), .A2(n1243), .ZN(n1265) );
NAND2_X1 U975 ( .A1(n1268), .A2(n1079), .ZN(n1266) );
NAND2_X1 U976 ( .A1(n1269), .A2(n1243), .ZN(n1079) );
XOR2_X1 U977 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U978 ( .A(n1272), .B(n1179), .Z(n1271) );
NAND2_X1 U979 ( .A1(G224), .A2(n1083), .ZN(n1179) );
NAND2_X1 U980 ( .A1(KEYINPUT30), .A2(n1273), .ZN(n1272) );
XOR2_X1 U981 ( .A(G125), .B(n1168), .Z(n1273) );
INV_X1 U982 ( .A(n1173), .ZN(n1168) );
XOR2_X1 U983 ( .A(n1163), .B(KEYINPUT14), .Z(n1270) );
NAND2_X1 U984 ( .A1(n1274), .A2(n1275), .ZN(n1163) );
NAND2_X1 U985 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U986 ( .A(n1278), .B(n1120), .Z(n1277) );
XOR2_X1 U987 ( .A(KEYINPUT61), .B(n1279), .Z(n1276) );
XOR2_X1 U988 ( .A(n1280), .B(KEYINPUT11), .Z(n1274) );
NAND2_X1 U989 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XNOR2_X1 U990 ( .A(n1120), .B(n1278), .ZN(n1282) );
NOR2_X1 U991 ( .A1(KEYINPUT32), .A2(n1119), .ZN(n1278) );
XOR2_X1 U992 ( .A(n1283), .B(n1284), .Z(n1119) );
XOR2_X1 U993 ( .A(KEYINPUT39), .B(n1285), .Z(n1284) );
XNOR2_X1 U994 ( .A(n1286), .B(n1287), .ZN(n1120) );
XOR2_X1 U995 ( .A(KEYINPUT61), .B(n1117), .Z(n1281) );
INV_X1 U996 ( .A(n1279), .ZN(n1117) );
XOR2_X1 U997 ( .A(G122), .B(G110), .Z(n1279) );
XNOR2_X1 U998 ( .A(KEYINPUT40), .B(KEYINPUT4), .ZN(n1268) );
NAND2_X1 U999 ( .A1(G221), .A2(n1288), .ZN(n1050) );
INV_X1 U1000 ( .A(n1046), .ZN(n1051) );
XOR2_X1 U1001 ( .A(n1289), .B(G469), .Z(n1046) );
NAND2_X1 U1002 ( .A1(n1290), .A2(n1243), .ZN(n1289) );
XOR2_X1 U1003 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U1004 ( .A(n1159), .B(n1293), .Z(n1292) );
NAND2_X1 U1005 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NAND2_X1 U1006 ( .A1(n1155), .A2(G110), .ZN(n1295) );
NAND2_X1 U1007 ( .A1(n1296), .A2(n1156), .ZN(n1294) );
XNOR2_X1 U1008 ( .A(n1155), .B(KEYINPUT15), .ZN(n1296) );
XNOR2_X1 U1009 ( .A(n1297), .B(n1298), .ZN(n1155) );
XOR2_X1 U1010 ( .A(KEYINPUT7), .B(G140), .Z(n1298) );
NAND2_X1 U1011 ( .A1(G227), .A2(n1083), .ZN(n1297) );
XOR2_X1 U1012 ( .A(n1299), .B(n1300), .Z(n1159) );
INV_X1 U1013 ( .A(n1283), .ZN(n1300) );
XNOR2_X1 U1014 ( .A(G101), .B(n1259), .ZN(n1283) );
XOR2_X1 U1015 ( .A(G104), .B(KEYINPUT60), .Z(n1259) );
XOR2_X1 U1016 ( .A(n1100), .B(n1246), .Z(n1299) );
XOR2_X1 U1017 ( .A(G128), .B(n1285), .Z(n1246) );
XOR2_X1 U1018 ( .A(G107), .B(KEYINPUT44), .Z(n1285) );
NAND2_X1 U1019 ( .A1(n1301), .A2(n1302), .ZN(n1100) );
NAND2_X1 U1020 ( .A1(G146), .A2(n1214), .ZN(n1302) );
XOR2_X1 U1021 ( .A(KEYINPUT2), .B(n1303), .Z(n1301) );
NOR2_X1 U1022 ( .A1(G146), .A2(n1214), .ZN(n1303) );
XNOR2_X1 U1023 ( .A(KEYINPUT58), .B(n1153), .ZN(n1291) );
NOR2_X1 U1024 ( .A1(n1238), .A2(n1063), .ZN(n1060) );
XNOR2_X1 U1025 ( .A(n1304), .B(n1126), .ZN(n1063) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1288), .ZN(n1126) );
NAND2_X1 U1027 ( .A1(G234), .A2(n1243), .ZN(n1288) );
NAND2_X1 U1028 ( .A1(n1125), .A2(n1243), .ZN(n1304) );
XNOR2_X1 U1029 ( .A(n1305), .B(n1306), .ZN(n1125) );
XOR2_X1 U1030 ( .A(n1307), .B(n1308), .Z(n1306) );
AND2_X1 U1031 ( .A1(n1251), .A2(G221), .ZN(n1308) );
AND2_X1 U1032 ( .A1(G234), .A2(n1083), .ZN(n1251) );
NOR2_X1 U1033 ( .A1(KEYINPUT53), .A2(n1309), .ZN(n1307) );
XOR2_X1 U1034 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1035 ( .A(n1286), .B(n1312), .Z(n1311) );
NOR2_X1 U1036 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1037 ( .A(n1315), .B(KEYINPUT55), .Z(n1314) );
NAND2_X1 U1038 ( .A1(n1316), .A2(G146), .ZN(n1315) );
NOR2_X1 U1039 ( .A1(G146), .A2(n1316), .ZN(n1313) );
XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n1091), .ZN(n1316) );
XOR2_X1 U1041 ( .A(G140), .B(G125), .Z(n1091) );
XOR2_X1 U1042 ( .A(n1156), .B(G128), .Z(n1310) );
NAND2_X1 U1043 ( .A1(KEYINPUT48), .A2(G137), .ZN(n1305) );
INV_X1 U1044 ( .A(n1231), .ZN(n1238) );
XNOR2_X1 U1045 ( .A(G472), .B(n1317), .ZN(n1231) );
NOR2_X1 U1046 ( .A1(KEYINPUT13), .A2(n1075), .ZN(n1317) );
NAND2_X1 U1047 ( .A1(n1318), .A2(n1243), .ZN(n1075) );
INV_X1 U1048 ( .A(G902), .ZN(n1243) );
XOR2_X1 U1049 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1050 ( .A(n1321), .B(n1145), .ZN(n1320) );
XNOR2_X1 U1051 ( .A(n1322), .B(n1287), .ZN(n1145) );
XOR2_X1 U1052 ( .A(G113), .B(G116), .Z(n1287) );
NAND2_X1 U1053 ( .A1(KEYINPUT33), .A2(n1286), .ZN(n1322) );
XNOR2_X1 U1054 ( .A(G119), .B(KEYINPUT28), .ZN(n1286) );
NAND2_X1 U1055 ( .A1(KEYINPUT35), .A2(n1143), .ZN(n1321) );
XOR2_X1 U1056 ( .A(n1153), .B(n1173), .Z(n1143) );
NAND2_X1 U1057 ( .A1(n1323), .A2(n1324), .ZN(n1173) );
NAND2_X1 U1058 ( .A1(n1325), .A2(n1099), .ZN(n1324) );
XOR2_X1 U1059 ( .A(n1326), .B(KEYINPUT36), .Z(n1323) );
OR2_X1 U1060 ( .A1(n1325), .A2(n1099), .ZN(n1326) );
INV_X1 U1061 ( .A(G128), .ZN(n1099) );
NAND4_X1 U1062 ( .A1(n1327), .A2(n1328), .A3(n1329), .A4(n1330), .ZN(n1325) );
OR2_X1 U1063 ( .A1(n1214), .A2(KEYINPUT41), .ZN(n1330) );
NAND3_X1 U1064 ( .A1(n1331), .A2(n1214), .A3(KEYINPUT41), .ZN(n1329) );
XOR2_X1 U1065 ( .A(KEYINPUT18), .B(n1332), .Z(n1331) );
NAND3_X1 U1066 ( .A1(KEYINPUT5), .A2(n1333), .A3(n1332), .ZN(n1328) );
INV_X1 U1067 ( .A(G146), .ZN(n1332) );
NAND2_X1 U1068 ( .A1(KEYINPUT18), .A2(n1214), .ZN(n1333) );
INV_X1 U1069 ( .A(G143), .ZN(n1214) );
NAND3_X1 U1070 ( .A1(n1334), .A2(n1335), .A3(G146), .ZN(n1327) );
INV_X1 U1071 ( .A(KEYINPUT5), .ZN(n1335) );
OR2_X1 U1072 ( .A1(KEYINPUT18), .A2(G143), .ZN(n1334) );
XNOR2_X1 U1073 ( .A(n1097), .B(n1098), .ZN(n1153) );
INV_X1 U1074 ( .A(G131), .ZN(n1098) );
XNOR2_X1 U1075 ( .A(G137), .B(n1249), .ZN(n1097) );
XOR2_X1 U1076 ( .A(G134), .B(KEYINPUT63), .Z(n1249) );
XOR2_X1 U1077 ( .A(n1336), .B(n1337), .Z(n1319) );
XNOR2_X1 U1078 ( .A(KEYINPUT45), .B(n1146), .ZN(n1337) );
NAND3_X1 U1079 ( .A1(n1261), .A2(n1083), .A3(G210), .ZN(n1146) );
INV_X1 U1080 ( .A(G953), .ZN(n1083) );
INV_X1 U1081 ( .A(G237), .ZN(n1261) );
NOR2_X1 U1082 ( .A1(G101), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1083 ( .A(KEYINPUT47), .B(KEYINPUT0), .Z(n1338) );
INV_X1 U1084 ( .A(G110), .ZN(n1156) );
endmodule


