//Key = 1000110000001111000101010001111110110100010111110100000001001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384;

XNOR2_X1 U756 ( .A(G107), .B(n1049), .ZN(G9) );
NOR2_X1 U757 ( .A1(n1050), .A2(n1051), .ZN(G75) );
NOR4_X1 U758 ( .A1(G953), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1051) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U762 ( .A(n1061), .ZN(n1060) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1062) );
NOR2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR3_X1 U770 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1074) );
AND2_X1 U771 ( .A1(n1079), .A2(KEYINPUT50), .ZN(n1078) );
NOR3_X1 U772 ( .A1(KEYINPUT50), .A2(n1080), .A3(n1081), .ZN(n1077) );
NOR2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(n1072) );
NOR2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR3_X1 U775 ( .A1(n1065), .A2(n1086), .A3(n1071), .ZN(n1057) );
INV_X1 U776 ( .A(n1087), .ZN(n1071) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
INV_X1 U778 ( .A(n1090), .ZN(n1065) );
NOR3_X1 U779 ( .A1(n1052), .A2(G953), .A3(G952), .ZN(n1050) );
AND4_X1 U780 ( .A1(n1087), .A2(n1061), .A3(n1091), .A4(n1092), .ZN(n1052) );
NOR3_X1 U781 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U783 ( .A1(G475), .A2(KEYINPUT17), .ZN(n1097) );
XOR2_X1 U784 ( .A(n1098), .B(n1099), .Z(n1091) );
XOR2_X1 U785 ( .A(n1100), .B(n1101), .Z(G72) );
NOR2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
AND2_X1 U787 ( .A1(G227), .A2(G900), .ZN(n1102) );
NAND2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1103), .ZN(n1105) );
XNOR2_X1 U790 ( .A(n1107), .B(n1108), .ZN(n1106) );
NAND3_X1 U791 ( .A1(G900), .A2(n1107), .A3(G953), .ZN(n1104) );
XNOR2_X1 U792 ( .A(n1109), .B(n1110), .ZN(n1107) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1110) );
XNOR2_X1 U794 ( .A(n1113), .B(G131), .ZN(n1112) );
NOR2_X1 U795 ( .A1(G137), .A2(KEYINPUT42), .ZN(n1111) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(n1109) );
NOR3_X1 U797 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
AND2_X1 U798 ( .A1(n1119), .A2(KEYINPUT11), .ZN(n1118) );
NOR2_X1 U799 ( .A1(KEYINPUT11), .A2(n1120), .ZN(n1117) );
NAND2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(G69) );
NAND2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U802 ( .A1(G953), .A2(n1125), .ZN(n1124) );
NAND3_X1 U803 ( .A1(G953), .A2(n1126), .A3(n1127), .ZN(n1121) );
XNOR2_X1 U804 ( .A(n1123), .B(KEYINPUT2), .ZN(n1127) );
XNOR2_X1 U805 ( .A(n1128), .B(n1129), .ZN(n1123) );
NOR2_X1 U806 ( .A1(n1130), .A2(G953), .ZN(n1129) );
AND2_X1 U807 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1128) );
NAND2_X1 U809 ( .A1(G953), .A2(n1135), .ZN(n1134) );
XOR2_X1 U810 ( .A(KEYINPUT38), .B(n1136), .Z(n1133) );
NOR2_X1 U811 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U812 ( .A(KEYINPUT53), .B(n1139), .Z(n1138) );
NOR2_X1 U813 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U814 ( .A(KEYINPUT16), .B(n1142), .Z(n1141) );
AND2_X1 U815 ( .A1(n1142), .A2(n1140), .ZN(n1137) );
XOR2_X1 U816 ( .A(n1143), .B(n1144), .Z(n1140) );
XOR2_X1 U817 ( .A(KEYINPUT26), .B(G113), .Z(n1144) );
XOR2_X1 U818 ( .A(G122), .B(G110), .Z(n1142) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1126) );
NOR2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XNOR2_X1 U821 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U822 ( .A(KEYINPUT52), .B(n1149), .Z(n1148) );
NOR2_X1 U823 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1145), .A2(n1152), .ZN(G63) );
XOR2_X1 U825 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U826 ( .A1(n1155), .A2(KEYINPUT63), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1156), .A2(n1151), .ZN(n1155) );
NOR2_X1 U828 ( .A1(n1145), .A2(n1157), .ZN(G60) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND3_X1 U830 ( .A1(G475), .A2(n1054), .A3(n1160), .ZN(n1158) );
XNOR2_X1 U831 ( .A(G902), .B(KEYINPUT31), .ZN(n1160) );
XOR2_X1 U832 ( .A(n1161), .B(n1162), .Z(G6) );
NOR2_X1 U833 ( .A1(KEYINPUT36), .A2(n1163), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1145), .A2(n1164), .ZN(G57) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND2_X1 U837 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
NAND2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
OR2_X1 U839 ( .A1(n1151), .A2(n1173), .ZN(n1172) );
XOR2_X1 U840 ( .A(KEYINPUT57), .B(n1174), .Z(n1169) );
NOR3_X1 U841 ( .A1(n1151), .A2(n1173), .A3(n1171), .ZN(n1174) );
NOR2_X1 U842 ( .A1(G101), .A2(KEYINPUT1), .ZN(n1165) );
NOR2_X1 U843 ( .A1(n1145), .A2(n1175), .ZN(G54) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U846 ( .A1(n1180), .A2(n1151), .ZN(n1178) );
XOR2_X1 U847 ( .A(n1181), .B(n1182), .Z(n1176) );
NOR2_X1 U848 ( .A1(KEYINPUT61), .A2(n1183), .ZN(n1182) );
NOR2_X1 U849 ( .A1(n1184), .A2(n1185), .ZN(n1181) );
NOR2_X1 U850 ( .A1(n1186), .A2(n1114), .ZN(n1185) );
NOR2_X1 U851 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
INV_X1 U852 ( .A(KEYINPUT27), .ZN(n1188) );
NOR2_X1 U853 ( .A1(KEYINPUT8), .A2(n1189), .ZN(n1187) );
NOR2_X1 U854 ( .A1(n1190), .A2(n1191), .ZN(n1184) );
NOR2_X1 U855 ( .A1(n1192), .A2(KEYINPUT8), .ZN(n1190) );
AND2_X1 U856 ( .A1(n1114), .A2(KEYINPUT27), .ZN(n1192) );
NOR3_X1 U857 ( .A1(n1145), .A2(n1193), .A3(n1194), .ZN(G51) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U859 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U860 ( .A1(KEYINPUT22), .A2(n1199), .ZN(n1198) );
INV_X1 U861 ( .A(KEYINPUT62), .ZN(n1195) );
NOR2_X1 U862 ( .A1(KEYINPUT62), .A2(n1200), .ZN(n1193) );
XOR2_X1 U863 ( .A(n1197), .B(n1201), .Z(n1200) );
NOR2_X1 U864 ( .A1(KEYINPUT22), .A2(n1202), .ZN(n1201) );
INV_X1 U865 ( .A(n1199), .ZN(n1202) );
XOR2_X1 U866 ( .A(n1203), .B(n1204), .Z(n1197) );
XOR2_X1 U867 ( .A(n1205), .B(n1206), .Z(n1203) );
NOR3_X1 U868 ( .A1(n1151), .A2(n1207), .A3(n1208), .ZN(n1206) );
INV_X1 U869 ( .A(G210), .ZN(n1208) );
NAND2_X1 U870 ( .A1(G902), .A2(n1054), .ZN(n1151) );
NAND3_X1 U871 ( .A1(n1132), .A2(n1209), .A3(n1108), .ZN(n1054) );
AND4_X1 U872 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1108) );
NOR4_X1 U873 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
INV_X1 U874 ( .A(n1218), .ZN(n1217) );
NOR3_X1 U875 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1216) );
NOR2_X1 U876 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
AND2_X1 U877 ( .A1(n1084), .A2(n1079), .ZN(n1222) );
INV_X1 U878 ( .A(n1224), .ZN(n1212) );
NAND2_X1 U879 ( .A1(n1225), .A2(n1079), .ZN(n1210) );
XNOR2_X1 U880 ( .A(n1226), .B(KEYINPUT21), .ZN(n1225) );
XNOR2_X1 U881 ( .A(KEYINPUT34), .B(n1131), .ZN(n1209) );
AND4_X1 U882 ( .A1(n1227), .A2(n1228), .A3(n1049), .A4(n1229), .ZN(n1132) );
NOR3_X1 U883 ( .A1(n1230), .A2(n1231), .A3(n1161), .ZN(n1229) );
AND3_X1 U884 ( .A1(n1061), .A2(n1232), .A3(n1085), .ZN(n1161) );
NOR2_X1 U885 ( .A1(n1233), .A2(n1234), .ZN(n1230) );
NOR2_X1 U886 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
XNOR2_X1 U887 ( .A(KEYINPUT48), .B(n1237), .ZN(n1236) );
XOR2_X1 U888 ( .A(n1238), .B(KEYINPUT15), .Z(n1235) );
NAND3_X1 U889 ( .A1(n1061), .A2(n1232), .A3(n1084), .ZN(n1049) );
NAND3_X1 U890 ( .A1(n1089), .A2(n1232), .A3(n1239), .ZN(n1227) );
XNOR2_X1 U891 ( .A(n1240), .B(KEYINPUT12), .ZN(n1239) );
NAND2_X1 U892 ( .A1(KEYINPUT45), .A2(n1241), .ZN(n1205) );
NOR2_X1 U893 ( .A1(n1103), .A2(G952), .ZN(n1145) );
XNOR2_X1 U894 ( .A(G146), .B(n1242), .ZN(G48) );
NAND2_X1 U895 ( .A1(KEYINPUT46), .A2(n1215), .ZN(n1242) );
AND3_X1 U896 ( .A1(n1085), .A2(n1076), .A3(n1243), .ZN(n1215) );
XOR2_X1 U897 ( .A(G143), .B(n1244), .Z(G45) );
NOR4_X1 U898 ( .A1(KEYINPUT39), .A2(n1221), .A3(n1219), .A4(n1245), .ZN(n1244) );
INV_X1 U899 ( .A(n1223), .ZN(n1245) );
XNOR2_X1 U900 ( .A(G140), .B(n1218), .ZN(G42) );
NAND4_X1 U901 ( .A1(n1079), .A2(n1246), .A3(n1085), .A4(n1088), .ZN(n1218) );
XOR2_X1 U902 ( .A(n1247), .B(n1248), .Z(G39) );
NOR2_X1 U903 ( .A1(KEYINPUT40), .A2(n1249), .ZN(n1248) );
NAND2_X1 U904 ( .A1(n1250), .A2(n1251), .ZN(n1247) );
NAND4_X1 U905 ( .A1(n1243), .A2(n1083), .A3(n1240), .A4(n1252), .ZN(n1251) );
OR2_X1 U906 ( .A1(n1211), .A2(n1252), .ZN(n1250) );
INV_X1 U907 ( .A(KEYINPUT47), .ZN(n1252) );
NAND2_X1 U908 ( .A1(n1090), .A2(n1243), .ZN(n1211) );
NOR2_X1 U909 ( .A1(n1075), .A2(n1083), .ZN(n1090) );
INV_X1 U910 ( .A(n1079), .ZN(n1083) );
INV_X1 U911 ( .A(n1240), .ZN(n1075) );
XOR2_X1 U912 ( .A(n1253), .B(n1254), .Z(G36) );
XNOR2_X1 U913 ( .A(KEYINPUT32), .B(n1113), .ZN(n1254) );
NAND4_X1 U914 ( .A1(n1255), .A2(n1079), .A3(n1246), .A4(n1084), .ZN(n1253) );
XNOR2_X1 U915 ( .A(n1089), .B(KEYINPUT35), .ZN(n1255) );
XOR2_X1 U916 ( .A(n1256), .B(n1257), .Z(G33) );
XNOR2_X1 U917 ( .A(G131), .B(KEYINPUT24), .ZN(n1257) );
NAND2_X1 U918 ( .A1(n1226), .A2(n1079), .ZN(n1256) );
NOR2_X1 U919 ( .A1(n1080), .A2(n1094), .ZN(n1079) );
INV_X1 U920 ( .A(n1081), .ZN(n1094) );
XOR2_X1 U921 ( .A(n1258), .B(KEYINPUT9), .Z(n1080) );
AND3_X1 U922 ( .A1(n1246), .A2(n1085), .A3(n1089), .ZN(n1226) );
XOR2_X1 U923 ( .A(n1259), .B(G128), .Z(G30) );
NAND2_X1 U924 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND3_X1 U925 ( .A1(n1076), .A2(n1262), .A3(n1263), .ZN(n1261) );
INV_X1 U926 ( .A(KEYINPUT29), .ZN(n1263) );
NAND2_X1 U927 ( .A1(n1224), .A2(KEYINPUT29), .ZN(n1260) );
NOR2_X1 U928 ( .A1(n1262), .A2(n1234), .ZN(n1224) );
NAND2_X1 U929 ( .A1(n1243), .A2(n1084), .ZN(n1262) );
AND3_X1 U930 ( .A1(n1264), .A2(n1265), .A3(n1246), .ZN(n1243) );
INV_X1 U931 ( .A(n1221), .ZN(n1246) );
NAND2_X1 U932 ( .A1(n1067), .A2(n1266), .ZN(n1221) );
XNOR2_X1 U933 ( .A(G101), .B(n1267), .ZN(G3) );
NAND3_X1 U934 ( .A1(n1089), .A2(n1232), .A3(n1240), .ZN(n1267) );
XOR2_X1 U935 ( .A(G125), .B(n1214), .Z(G27) );
AND4_X1 U936 ( .A1(n1085), .A2(n1088), .A3(n1268), .A4(n1087), .ZN(n1214) );
AND2_X1 U937 ( .A1(n1266), .A2(n1076), .ZN(n1268) );
NAND2_X1 U938 ( .A1(n1056), .A2(n1269), .ZN(n1266) );
NAND4_X1 U939 ( .A1(G953), .A2(G902), .A3(n1270), .A4(n1271), .ZN(n1269) );
INV_X1 U940 ( .A(G900), .ZN(n1271) );
XOR2_X1 U941 ( .A(n1231), .B(n1272), .Z(G24) );
NOR2_X1 U942 ( .A1(KEYINPUT3), .A2(n1273), .ZN(n1272) );
AND3_X1 U943 ( .A1(n1274), .A2(n1061), .A3(n1223), .ZN(n1231) );
NOR3_X1 U944 ( .A1(n1275), .A2(n1234), .A3(n1276), .ZN(n1223) );
NOR2_X1 U945 ( .A1(n1265), .A2(n1264), .ZN(n1061) );
XNOR2_X1 U946 ( .A(n1277), .B(n1278), .ZN(G21) );
NOR2_X1 U947 ( .A1(n1234), .A2(n1238), .ZN(n1278) );
NAND4_X1 U948 ( .A1(n1274), .A2(n1240), .A3(n1264), .A4(n1265), .ZN(n1238) );
XNOR2_X1 U949 ( .A(n1279), .B(n1280), .ZN(G18) );
NOR2_X1 U950 ( .A1(KEYINPUT10), .A2(n1131), .ZN(n1280) );
NAND4_X1 U951 ( .A1(n1274), .A2(n1089), .A3(n1084), .A4(n1076), .ZN(n1131) );
NOR2_X1 U952 ( .A1(n1275), .A2(n1281), .ZN(n1084) );
XOR2_X1 U953 ( .A(G113), .B(n1282), .Z(G15) );
NOR2_X1 U954 ( .A1(n1234), .A2(n1237), .ZN(n1282) );
NAND3_X1 U955 ( .A1(n1089), .A2(n1085), .A3(n1274), .ZN(n1237) );
AND2_X1 U956 ( .A1(n1087), .A2(n1283), .ZN(n1274) );
NOR2_X1 U957 ( .A1(n1068), .A2(n1284), .ZN(n1087) );
INV_X1 U958 ( .A(n1069), .ZN(n1284) );
NOR2_X1 U959 ( .A1(n1276), .A2(n1285), .ZN(n1085) );
INV_X1 U960 ( .A(n1219), .ZN(n1089) );
NAND2_X1 U961 ( .A1(n1286), .A2(n1265), .ZN(n1219) );
NAND2_X1 U962 ( .A1(n1287), .A2(n1288), .ZN(G12) );
NAND2_X1 U963 ( .A1(G110), .A2(n1228), .ZN(n1288) );
XOR2_X1 U964 ( .A(KEYINPUT19), .B(n1289), .Z(n1287) );
NOR2_X1 U965 ( .A1(G110), .A2(n1228), .ZN(n1289) );
NAND3_X1 U966 ( .A1(n1088), .A2(n1232), .A3(n1240), .ZN(n1228) );
NOR2_X1 U967 ( .A1(n1281), .A2(n1285), .ZN(n1240) );
INV_X1 U968 ( .A(n1275), .ZN(n1285) );
XOR2_X1 U969 ( .A(n1093), .B(KEYINPUT37), .Z(n1275) );
XOR2_X1 U970 ( .A(n1290), .B(n1156), .Z(n1093) );
INV_X1 U971 ( .A(G478), .ZN(n1156) );
NAND2_X1 U972 ( .A1(n1153), .A2(n1291), .ZN(n1290) );
XOR2_X1 U973 ( .A(n1292), .B(n1293), .Z(n1153) );
XNOR2_X1 U974 ( .A(n1294), .B(n1295), .ZN(n1293) );
XNOR2_X1 U975 ( .A(n1113), .B(G122), .ZN(n1295) );
XOR2_X1 U976 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U977 ( .A(n1298), .B(n1299), .Z(n1296) );
NOR2_X1 U978 ( .A1(KEYINPUT25), .A2(G116), .ZN(n1299) );
NAND2_X1 U979 ( .A1(G217), .A2(n1300), .ZN(n1298) );
INV_X1 U980 ( .A(n1276), .ZN(n1281) );
XNOR2_X1 U981 ( .A(n1096), .B(n1301), .ZN(n1276) );
XOR2_X1 U982 ( .A(KEYINPUT5), .B(G475), .Z(n1301) );
NAND2_X1 U983 ( .A1(n1159), .A2(n1291), .ZN(n1096) );
XNOR2_X1 U984 ( .A(n1302), .B(n1303), .ZN(n1159) );
XNOR2_X1 U985 ( .A(n1163), .B(n1304), .ZN(n1303) );
NOR2_X1 U986 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U987 ( .A(n1307), .B(KEYINPUT0), .Z(n1306) );
NAND2_X1 U988 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NOR2_X1 U989 ( .A1(n1309), .A2(n1308), .ZN(n1305) );
XNOR2_X1 U990 ( .A(KEYINPUT43), .B(n1310), .ZN(n1308) );
XNOR2_X1 U991 ( .A(n1311), .B(G143), .ZN(n1309) );
NAND2_X1 U992 ( .A1(G214), .A2(n1312), .ZN(n1311) );
INV_X1 U993 ( .A(G104), .ZN(n1163) );
XOR2_X1 U994 ( .A(n1313), .B(n1314), .Z(n1302) );
NOR2_X1 U995 ( .A1(KEYINPUT55), .A2(n1315), .ZN(n1314) );
INV_X1 U996 ( .A(G146), .ZN(n1315) );
NAND2_X1 U997 ( .A1(n1316), .A2(n1317), .ZN(n1313) );
NAND2_X1 U998 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND2_X1 U999 ( .A1(n1320), .A2(n1120), .ZN(n1319) );
INV_X1 U1000 ( .A(n1321), .ZN(n1120) );
INV_X1 U1001 ( .A(n1322), .ZN(n1318) );
NAND2_X1 U1002 ( .A1(n1323), .A2(n1322), .ZN(n1316) );
XNOR2_X1 U1003 ( .A(n1324), .B(n1119), .ZN(n1323) );
AND3_X1 U1004 ( .A1(n1067), .A2(n1283), .A3(n1076), .ZN(n1232) );
INV_X1 U1005 ( .A(n1234), .ZN(n1076) );
NAND2_X1 U1006 ( .A1(n1258), .A2(n1081), .ZN(n1234) );
NAND2_X1 U1007 ( .A1(G214), .A2(n1325), .ZN(n1081) );
XOR2_X1 U1008 ( .A(n1098), .B(n1326), .Z(n1258) );
NOR2_X1 U1009 ( .A1(n1099), .A2(KEYINPUT18), .ZN(n1326) );
AND2_X1 U1010 ( .A1(G210), .A2(n1327), .ZN(n1099) );
XNOR2_X1 U1011 ( .A(KEYINPUT13), .B(n1325), .ZN(n1327) );
INV_X1 U1012 ( .A(n1207), .ZN(n1325) );
NOR2_X1 U1013 ( .A1(n1328), .A2(G237), .ZN(n1207) );
INV_X1 U1014 ( .A(n1329), .ZN(n1328) );
NAND2_X1 U1015 ( .A1(n1330), .A2(n1291), .ZN(n1098) );
XNOR2_X1 U1016 ( .A(n1199), .B(n1331), .ZN(n1330) );
XNOR2_X1 U1017 ( .A(n1204), .B(n1119), .ZN(n1331) );
XNOR2_X1 U1018 ( .A(n1332), .B(n1333), .ZN(n1204) );
NOR2_X1 U1019 ( .A1(G953), .A2(n1125), .ZN(n1333) );
INV_X1 U1020 ( .A(G224), .ZN(n1125) );
XNOR2_X1 U1021 ( .A(n1334), .B(n1335), .ZN(n1199) );
XOR2_X1 U1022 ( .A(KEYINPUT59), .B(G110), .Z(n1335) );
XNOR2_X1 U1023 ( .A(n1143), .B(n1322), .ZN(n1334) );
XOR2_X1 U1024 ( .A(G113), .B(n1273), .Z(n1322) );
INV_X1 U1025 ( .A(G122), .ZN(n1273) );
XOR2_X1 U1026 ( .A(n1336), .B(n1337), .Z(n1143) );
XOR2_X1 U1027 ( .A(n1338), .B(n1339), .Z(n1337) );
NOR2_X1 U1028 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
AND2_X1 U1029 ( .A1(KEYINPUT54), .A2(n1342), .ZN(n1341) );
NOR2_X1 U1030 ( .A1(KEYINPUT7), .A2(n1342), .ZN(n1340) );
XNOR2_X1 U1031 ( .A(G116), .B(G119), .ZN(n1336) );
NAND2_X1 U1032 ( .A1(n1056), .A2(n1343), .ZN(n1283) );
NAND4_X1 U1033 ( .A1(G953), .A2(G902), .A3(n1270), .A4(n1135), .ZN(n1343) );
INV_X1 U1034 ( .A(G898), .ZN(n1135) );
NAND3_X1 U1035 ( .A1(n1270), .A2(n1103), .A3(G952), .ZN(n1056) );
NAND2_X1 U1036 ( .A1(G237), .A2(G234), .ZN(n1270) );
AND2_X1 U1037 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1344), .ZN(n1069) );
XOR2_X1 U1039 ( .A(n1345), .B(n1180), .Z(n1068) );
INV_X1 U1040 ( .A(G469), .ZN(n1180) );
NAND2_X1 U1041 ( .A1(n1346), .A2(n1291), .ZN(n1345) );
XOR2_X1 U1042 ( .A(n1347), .B(n1348), .Z(n1346) );
XNOR2_X1 U1043 ( .A(n1191), .B(n1179), .ZN(n1348) );
XNOR2_X1 U1044 ( .A(n1349), .B(n1350), .ZN(n1179) );
XNOR2_X1 U1045 ( .A(n1324), .B(G110), .ZN(n1350) );
NAND2_X1 U1046 ( .A1(G227), .A2(n1103), .ZN(n1349) );
INV_X1 U1047 ( .A(n1189), .ZN(n1191) );
XNOR2_X1 U1048 ( .A(n1342), .B(n1351), .ZN(n1189) );
NOR2_X1 U1049 ( .A1(KEYINPUT33), .A2(n1352), .ZN(n1351) );
XNOR2_X1 U1050 ( .A(n1338), .B(KEYINPUT44), .ZN(n1352) );
XNOR2_X1 U1051 ( .A(G104), .B(n1294), .ZN(n1338) );
INV_X1 U1052 ( .A(G107), .ZN(n1294) );
XNOR2_X1 U1053 ( .A(G101), .B(KEYINPUT49), .ZN(n1342) );
XOR2_X1 U1054 ( .A(n1114), .B(n1353), .Z(n1347) );
XOR2_X1 U1055 ( .A(n1183), .B(KEYINPUT6), .Z(n1353) );
XNOR2_X1 U1056 ( .A(G146), .B(n1354), .ZN(n1114) );
NOR2_X1 U1057 ( .A1(n1265), .A2(n1286), .ZN(n1088) );
INV_X1 U1058 ( .A(n1264), .ZN(n1286) );
XOR2_X1 U1059 ( .A(n1355), .B(n1150), .Z(n1264) );
NAND2_X1 U1060 ( .A1(G217), .A2(n1344), .ZN(n1150) );
NAND2_X1 U1061 ( .A1(G234), .A2(n1329), .ZN(n1344) );
XNOR2_X1 U1062 ( .A(n1291), .B(KEYINPUT30), .ZN(n1329) );
NAND2_X1 U1063 ( .A1(n1147), .A2(n1291), .ZN(n1355) );
XNOR2_X1 U1064 ( .A(n1356), .B(n1357), .ZN(n1147) );
XOR2_X1 U1065 ( .A(n1358), .B(n1359), .Z(n1357) );
XNOR2_X1 U1066 ( .A(G137), .B(G146), .ZN(n1359) );
NAND3_X1 U1067 ( .A1(n1360), .A2(n1361), .A3(n1320), .ZN(n1358) );
INV_X1 U1068 ( .A(n1116), .ZN(n1320) );
NOR2_X1 U1069 ( .A1(n1324), .A2(n1241), .ZN(n1116) );
INV_X1 U1070 ( .A(n1119), .ZN(n1241) );
OR2_X1 U1071 ( .A1(n1324), .A2(KEYINPUT23), .ZN(n1361) );
INV_X1 U1072 ( .A(G140), .ZN(n1324) );
NAND2_X1 U1073 ( .A1(n1321), .A2(KEYINPUT23), .ZN(n1360) );
NOR2_X1 U1074 ( .A1(n1119), .A2(G140), .ZN(n1321) );
XOR2_X1 U1075 ( .A(G125), .B(KEYINPUT20), .Z(n1119) );
XOR2_X1 U1076 ( .A(n1362), .B(n1363), .Z(n1356) );
AND2_X1 U1077 ( .A1(n1300), .A2(G221), .ZN(n1363) );
AND2_X1 U1078 ( .A1(G234), .A2(n1103), .ZN(n1300) );
INV_X1 U1079 ( .A(G953), .ZN(n1103) );
NAND2_X1 U1080 ( .A1(KEYINPUT14), .A2(n1364), .ZN(n1362) );
XOR2_X1 U1081 ( .A(G110), .B(n1365), .Z(n1364) );
XNOR2_X1 U1082 ( .A(G128), .B(n1277), .ZN(n1365) );
XOR2_X1 U1083 ( .A(n1366), .B(n1173), .Z(n1265) );
INV_X1 U1084 ( .A(G472), .ZN(n1173) );
NAND2_X1 U1085 ( .A1(n1367), .A2(n1291), .ZN(n1366) );
INV_X1 U1086 ( .A(G902), .ZN(n1291) );
XNOR2_X1 U1087 ( .A(n1171), .B(n1368), .ZN(n1367) );
XNOR2_X1 U1088 ( .A(G101), .B(n1168), .ZN(n1368) );
NAND2_X1 U1089 ( .A1(G210), .A2(n1312), .ZN(n1168) );
NOR2_X1 U1090 ( .A1(G953), .A2(G237), .ZN(n1312) );
XNOR2_X1 U1091 ( .A(n1369), .B(n1370), .ZN(n1171) );
XNOR2_X1 U1092 ( .A(G113), .B(n1183), .ZN(n1370) );
NAND2_X1 U1093 ( .A1(n1371), .A2(n1372), .ZN(n1183) );
NAND3_X1 U1094 ( .A1(n1373), .A2(n1113), .A3(KEYINPUT28), .ZN(n1372) );
XNOR2_X1 U1095 ( .A(n1310), .B(n1374), .ZN(n1373) );
AND2_X1 U1096 ( .A1(n1249), .A2(KEYINPUT60), .ZN(n1374) );
INV_X1 U1097 ( .A(G137), .ZN(n1249) );
INV_X1 U1098 ( .A(G131), .ZN(n1310) );
NAND2_X1 U1099 ( .A1(n1375), .A2(n1376), .ZN(n1371) );
NAND2_X1 U1100 ( .A1(KEYINPUT28), .A2(n1113), .ZN(n1376) );
INV_X1 U1101 ( .A(G134), .ZN(n1113) );
XNOR2_X1 U1102 ( .A(G131), .B(n1377), .ZN(n1375) );
NAND2_X1 U1103 ( .A1(G137), .A2(KEYINPUT60), .ZN(n1377) );
XOR2_X1 U1104 ( .A(n1332), .B(n1378), .Z(n1369) );
NOR2_X1 U1105 ( .A1(n1379), .A2(n1380), .ZN(n1378) );
NOR2_X1 U1106 ( .A1(n1381), .A2(n1277), .ZN(n1380) );
INV_X1 U1107 ( .A(G119), .ZN(n1277) );
XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1279), .ZN(n1381) );
INV_X1 U1109 ( .A(G116), .ZN(n1279) );
NOR2_X1 U1110 ( .A1(G119), .A2(n1382), .ZN(n1379) );
XNOR2_X1 U1111 ( .A(G116), .B(KEYINPUT51), .ZN(n1382) );
XOR2_X1 U1112 ( .A(n1383), .B(n1354), .Z(n1332) );
XOR2_X1 U1113 ( .A(n1297), .B(KEYINPUT56), .Z(n1354) );
XOR2_X1 U1114 ( .A(G128), .B(G143), .Z(n1297) );
NAND2_X1 U1115 ( .A1(n1384), .A2(KEYINPUT41), .ZN(n1383) );
XNOR2_X1 U1116 ( .A(G146), .B(KEYINPUT4), .ZN(n1384) );
endmodule


