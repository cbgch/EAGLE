//Key = 0111000101111000110001011100110000101001001011110010000010010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392;

XNOR2_X1 U758 ( .A(G107), .B(n1056), .ZN(G9) );
NOR2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(G75) );
NOR4_X1 U760 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U763 ( .A1(KEYINPUT29), .A2(n1067), .ZN(n1066) );
NOR4_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1068), .A2(n1072), .ZN(n1065) );
NOR2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U769 ( .A1(n1079), .A2(n1071), .ZN(n1078) );
NOR3_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U771 ( .A1(n1069), .A2(n1083), .ZN(n1082) );
NOR2_X1 U772 ( .A1(KEYINPUT18), .A2(n1084), .ZN(n1080) );
NOR2_X1 U773 ( .A1(n1085), .A2(n1069), .ZN(n1077) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR3_X1 U776 ( .A1(n1071), .A2(n1090), .A3(n1069), .ZN(n1073) );
INV_X1 U777 ( .A(n1091), .ZN(n1069) );
NOR2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
AND2_X1 U779 ( .A1(n1094), .A2(KEYINPUT29), .ZN(n1092) );
NAND3_X1 U780 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1059) );
NAND4_X1 U781 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND3_X1 U783 ( .A1(n1104), .A2(n1064), .A3(KEYINPUT18), .ZN(n1103) );
INV_X1 U784 ( .A(n1105), .ZN(n1064) );
NAND2_X1 U785 ( .A1(n1091), .A2(n1106), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND3_X1 U787 ( .A1(n1109), .A2(n1083), .A3(n1110), .ZN(n1108) );
INV_X1 U788 ( .A(KEYINPUT4), .ZN(n1083) );
NOR3_X1 U789 ( .A1(n1111), .A2(G953), .A3(G952), .ZN(n1057) );
INV_X1 U790 ( .A(n1095), .ZN(n1111) );
NAND4_X1 U791 ( .A1(n1112), .A2(n1099), .A3(n1113), .A4(n1114), .ZN(n1095) );
NOR4_X1 U792 ( .A1(n1110), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1114) );
XOR2_X1 U793 ( .A(n1118), .B(n1119), .Z(n1115) );
XOR2_X1 U794 ( .A(KEYINPUT50), .B(G472), .Z(n1119) );
XOR2_X1 U795 ( .A(n1120), .B(n1121), .Z(n1113) );
XOR2_X1 U796 ( .A(n1122), .B(G478), .Z(n1112) );
NAND2_X1 U797 ( .A1(n1123), .A2(n1124), .ZN(G72) );
NAND3_X1 U798 ( .A1(n1125), .A2(n1126), .A3(KEYINPUT9), .ZN(n1124) );
NAND2_X1 U799 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U800 ( .A1(n1062), .A2(n1096), .ZN(n1127) );
NAND2_X1 U801 ( .A1(n1129), .A2(n1130), .ZN(n1125) );
NAND2_X1 U802 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND3_X1 U803 ( .A1(G953), .A2(n1133), .A3(KEYINPUT59), .ZN(n1132) );
NAND4_X1 U804 ( .A1(G953), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1123) );
NAND2_X1 U805 ( .A1(n1129), .A2(KEYINPUT9), .ZN(n1136) );
OR2_X1 U806 ( .A1(n1129), .A2(KEYINPUT59), .ZN(n1135) );
INV_X1 U807 ( .A(n1128), .ZN(n1129) );
NAND2_X1 U808 ( .A1(n1137), .A2(n1138), .ZN(n1128) );
NAND2_X1 U809 ( .A1(G953), .A2(n1139), .ZN(n1138) );
XOR2_X1 U810 ( .A(n1140), .B(n1141), .Z(n1137) );
XNOR2_X1 U811 ( .A(KEYINPUT17), .B(n1142), .ZN(n1140) );
NOR2_X1 U812 ( .A1(KEYINPUT40), .A2(n1143), .ZN(n1142) );
XNOR2_X1 U813 ( .A(n1144), .B(n1145), .ZN(n1143) );
NAND2_X1 U814 ( .A1(KEYINPUT44), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U815 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U816 ( .A(KEYINPUT11), .B(n1149), .Z(n1148) );
NAND2_X1 U817 ( .A1(G900), .A2(G227), .ZN(n1134) );
XOR2_X1 U818 ( .A(n1150), .B(n1151), .Z(G69) );
XOR2_X1 U819 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U820 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U821 ( .A1(G953), .A2(n1156), .ZN(n1155) );
XOR2_X1 U822 ( .A(n1157), .B(n1158), .Z(n1154) );
NAND2_X1 U823 ( .A1(KEYINPUT61), .A2(n1159), .ZN(n1157) );
NAND2_X1 U824 ( .A1(n1160), .A2(n1161), .ZN(n1152) );
NAND2_X1 U825 ( .A1(G898), .A2(G224), .ZN(n1161) );
XNOR2_X1 U826 ( .A(KEYINPUT20), .B(n1096), .ZN(n1160) );
NOR2_X1 U827 ( .A1(n1162), .A2(G953), .ZN(n1150) );
NOR2_X1 U828 ( .A1(n1163), .A2(n1164), .ZN(G66) );
XOR2_X1 U829 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U830 ( .A1(KEYINPUT51), .A2(n1167), .ZN(n1166) );
NOR2_X1 U831 ( .A1(n1168), .A2(n1169), .ZN(n1165) );
NOR2_X1 U832 ( .A1(n1163), .A2(n1170), .ZN(G63) );
XOR2_X1 U833 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U834 ( .A1(KEYINPUT14), .A2(n1173), .ZN(n1172) );
NAND2_X1 U835 ( .A1(n1174), .A2(G478), .ZN(n1171) );
NOR2_X1 U836 ( .A1(n1163), .A2(n1175), .ZN(G60) );
XOR2_X1 U837 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U838 ( .A(n1178), .B(KEYINPUT38), .Z(n1177) );
NAND2_X1 U839 ( .A1(n1174), .A2(G475), .ZN(n1176) );
XNOR2_X1 U840 ( .A(G104), .B(n1179), .ZN(G6) );
NOR2_X1 U841 ( .A1(n1163), .A2(n1180), .ZN(G57) );
NOR2_X1 U842 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U843 ( .A(n1183), .B(KEYINPUT21), .Z(n1182) );
NAND2_X1 U844 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U845 ( .A1(n1184), .A2(n1185), .ZN(n1181) );
NAND2_X1 U846 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XOR2_X1 U847 ( .A(n1188), .B(n1189), .Z(n1184) );
XOR2_X1 U848 ( .A(n1190), .B(n1191), .Z(n1188) );
NAND2_X1 U849 ( .A1(n1174), .A2(G472), .ZN(n1190) );
NOR2_X1 U850 ( .A1(n1163), .A2(n1192), .ZN(G54) );
XOR2_X1 U851 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U852 ( .A(n1195), .B(n1196), .Z(n1194) );
NAND2_X1 U853 ( .A1(n1174), .A2(G469), .ZN(n1195) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(n1193) );
NOR2_X1 U855 ( .A1(KEYINPUT43), .A2(n1199), .ZN(n1198) );
NOR2_X1 U856 ( .A1(KEYINPUT57), .A2(n1200), .ZN(n1197) );
XOR2_X1 U857 ( .A(n1201), .B(n1202), .Z(n1200) );
NAND3_X1 U858 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1201) );
NAND2_X1 U859 ( .A1(KEYINPUT52), .A2(n1206), .ZN(n1205) );
NAND3_X1 U860 ( .A1(n1207), .A2(n1208), .A3(n1145), .ZN(n1204) );
NAND2_X1 U861 ( .A1(n1209), .A2(n1210), .ZN(n1203) );
NAND2_X1 U862 ( .A1(n1211), .A2(n1208), .ZN(n1210) );
INV_X1 U863 ( .A(KEYINPUT52), .ZN(n1208) );
XNOR2_X1 U864 ( .A(n1206), .B(KEYINPUT54), .ZN(n1211) );
NOR2_X1 U865 ( .A1(n1163), .A2(n1212), .ZN(G51) );
XOR2_X1 U866 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U867 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR2_X1 U868 ( .A1(KEYINPUT62), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U869 ( .A(n1218), .B(n1219), .ZN(n1217) );
NOR2_X1 U870 ( .A1(n1220), .A2(KEYINPUT33), .ZN(n1219) );
XOR2_X1 U871 ( .A(n1221), .B(n1222), .Z(n1213) );
NAND2_X1 U872 ( .A1(n1174), .A2(G210), .ZN(n1221) );
INV_X1 U873 ( .A(n1169), .ZN(n1174) );
NAND2_X1 U874 ( .A1(G902), .A2(n1223), .ZN(n1169) );
NAND2_X1 U875 ( .A1(n1162), .A2(n1131), .ZN(n1223) );
INV_X1 U876 ( .A(n1062), .ZN(n1131) );
NAND4_X1 U877 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1062) );
AND3_X1 U878 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1227) );
NAND2_X1 U879 ( .A1(n1231), .A2(n1232), .ZN(n1226) );
NAND2_X1 U880 ( .A1(n1233), .A2(n1084), .ZN(n1232) );
XOR2_X1 U881 ( .A(KEYINPUT24), .B(n1081), .Z(n1233) );
NAND3_X1 U882 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1224) );
NAND2_X1 U883 ( .A1(n1237), .A2(n1238), .ZN(n1235) );
NAND2_X1 U884 ( .A1(n1105), .A2(n1098), .ZN(n1238) );
NAND2_X1 U885 ( .A1(n1094), .A2(n1239), .ZN(n1237) );
INV_X1 U886 ( .A(n1060), .ZN(n1162) );
NAND4_X1 U887 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1060) );
AND4_X1 U888 ( .A1(n1244), .A2(n1245), .A3(n1056), .A4(n1246), .ZN(n1243) );
NAND3_X1 U889 ( .A1(n1091), .A2(n1247), .A3(n1094), .ZN(n1056) );
NOR2_X1 U890 ( .A1(n1248), .A2(n1249), .ZN(n1242) );
NOR2_X1 U891 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NOR2_X1 U892 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
NOR2_X1 U893 ( .A1(n1076), .A2(n1254), .ZN(n1253) );
INV_X1 U894 ( .A(n1098), .ZN(n1076) );
NOR2_X1 U895 ( .A1(n1255), .A2(n1256), .ZN(n1252) );
NAND3_X1 U896 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1241) );
NAND2_X1 U897 ( .A1(n1260), .A2(n1107), .ZN(n1258) );
NAND4_X1 U898 ( .A1(KEYINPUT30), .A2(n1093), .A3(n1091), .A4(n1087), .ZN(n1260) );
NAND2_X1 U899 ( .A1(n1239), .A2(n1261), .ZN(n1257) );
NAND3_X1 U900 ( .A1(n1071), .A2(n1256), .A3(n1262), .ZN(n1261) );
INV_X1 U901 ( .A(KEYINPUT46), .ZN(n1256) );
OR2_X1 U902 ( .A1(n1179), .A2(KEYINPUT30), .ZN(n1240) );
NAND3_X1 U903 ( .A1(n1091), .A2(n1247), .A3(n1093), .ZN(n1179) );
NOR2_X1 U904 ( .A1(n1096), .A2(G952), .ZN(n1163) );
XNOR2_X1 U905 ( .A(G146), .B(n1225), .ZN(G48) );
NAND4_X1 U906 ( .A1(n1236), .A2(n1234), .A3(n1093), .A4(n1239), .ZN(n1225) );
XNOR2_X1 U907 ( .A(G143), .B(n1228), .ZN(G45) );
NAND4_X1 U908 ( .A1(n1236), .A2(n1104), .A3(n1263), .A4(n1239), .ZN(n1228) );
NOR2_X1 U909 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U910 ( .A(n1266), .B(n1267), .Z(G42) );
NOR2_X1 U911 ( .A1(G140), .A2(KEYINPUT5), .ZN(n1267) );
NAND2_X1 U912 ( .A1(n1231), .A2(n1081), .ZN(n1266) );
INV_X1 U913 ( .A(n1268), .ZN(n1231) );
XNOR2_X1 U914 ( .A(G137), .B(n1269), .ZN(G39) );
NAND4_X1 U915 ( .A1(n1105), .A2(n1234), .A3(n1270), .A4(n1098), .ZN(n1269) );
NOR2_X1 U916 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XNOR2_X1 U917 ( .A(n1087), .B(KEYINPUT27), .ZN(n1272) );
NAND2_X1 U918 ( .A1(n1273), .A2(n1274), .ZN(G36) );
NAND2_X1 U919 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XOR2_X1 U920 ( .A(KEYINPUT3), .B(n1277), .Z(n1273) );
NOR2_X1 U921 ( .A1(n1275), .A2(n1276), .ZN(n1277) );
INV_X1 U922 ( .A(G134), .ZN(n1276) );
INV_X1 U923 ( .A(n1230), .ZN(n1275) );
NAND3_X1 U924 ( .A1(n1236), .A2(n1262), .A3(n1105), .ZN(n1230) );
XOR2_X1 U925 ( .A(G131), .B(n1278), .Z(G33) );
NOR2_X1 U926 ( .A1(n1084), .A2(n1268), .ZN(n1278) );
NAND3_X1 U927 ( .A1(n1236), .A2(n1093), .A3(n1105), .ZN(n1268) );
NOR2_X1 U928 ( .A1(n1279), .A2(n1110), .ZN(n1105) );
XNOR2_X1 U929 ( .A(G128), .B(n1280), .ZN(G30) );
NAND4_X1 U930 ( .A1(n1281), .A2(n1236), .A3(n1234), .A4(n1094), .ZN(n1280) );
INV_X1 U931 ( .A(n1254), .ZN(n1234) );
NOR2_X1 U932 ( .A1(n1282), .A2(n1271), .ZN(n1236) );
XNOR2_X1 U933 ( .A(n1239), .B(KEYINPUT23), .ZN(n1281) );
XOR2_X1 U934 ( .A(G101), .B(n1248), .Z(G3) );
AND3_X1 U935 ( .A1(n1098), .A2(n1247), .A3(n1104), .ZN(n1248) );
XNOR2_X1 U936 ( .A(G125), .B(n1229), .ZN(G27) );
NAND3_X1 U937 ( .A1(n1093), .A2(n1081), .A3(n1283), .ZN(n1229) );
NOR3_X1 U938 ( .A1(n1071), .A2(n1271), .A3(n1107), .ZN(n1283) );
INV_X1 U939 ( .A(n1239), .ZN(n1107) );
AND2_X1 U940 ( .A1(n1284), .A2(n1285), .ZN(n1271) );
NAND2_X1 U941 ( .A1(n1286), .A2(n1139), .ZN(n1285) );
INV_X1 U942 ( .A(G900), .ZN(n1139) );
XNOR2_X1 U943 ( .A(G122), .B(n1246), .ZN(G24) );
NAND4_X1 U944 ( .A1(n1287), .A2(n1091), .A3(n1288), .A4(n1117), .ZN(n1246) );
NOR2_X1 U945 ( .A1(n1289), .A2(n1116), .ZN(n1091) );
XNOR2_X1 U946 ( .A(G119), .B(n1290), .ZN(G21) );
NAND3_X1 U947 ( .A1(n1098), .A2(n1291), .A3(n1287), .ZN(n1290) );
XNOR2_X1 U948 ( .A(KEYINPUT0), .B(n1254), .ZN(n1291) );
NAND2_X1 U949 ( .A1(n1116), .A2(n1289), .ZN(n1254) );
XNOR2_X1 U950 ( .A(n1292), .B(n1293), .ZN(G18) );
NOR2_X1 U951 ( .A1(n1251), .A2(n1255), .ZN(n1293) );
INV_X1 U952 ( .A(n1262), .ZN(n1255) );
NOR2_X1 U953 ( .A1(n1084), .A2(n1070), .ZN(n1262) );
INV_X1 U954 ( .A(n1094), .ZN(n1070) );
NOR2_X1 U955 ( .A1(n1117), .A2(n1265), .ZN(n1094) );
INV_X1 U956 ( .A(n1104), .ZN(n1084) );
XNOR2_X1 U957 ( .A(G113), .B(n1245), .ZN(G15) );
NAND3_X1 U958 ( .A1(n1287), .A2(n1104), .A3(n1093), .ZN(n1245) );
NOR2_X1 U959 ( .A1(n1288), .A2(n1264), .ZN(n1093) );
INV_X1 U960 ( .A(n1117), .ZN(n1264) );
NOR2_X1 U961 ( .A1(n1116), .A2(n1294), .ZN(n1104) );
INV_X1 U962 ( .A(n1251), .ZN(n1287) );
NAND3_X1 U963 ( .A1(n1239), .A2(n1259), .A3(n1099), .ZN(n1251) );
INV_X1 U964 ( .A(n1071), .ZN(n1099) );
NAND2_X1 U965 ( .A1(n1295), .A2(n1089), .ZN(n1071) );
INV_X1 U966 ( .A(n1088), .ZN(n1295) );
XNOR2_X1 U967 ( .A(G110), .B(n1244), .ZN(G12) );
NAND3_X1 U968 ( .A1(n1098), .A2(n1247), .A3(n1081), .ZN(n1244) );
AND2_X1 U969 ( .A1(n1294), .A2(n1116), .ZN(n1081) );
XOR2_X1 U970 ( .A(n1296), .B(n1168), .Z(n1116) );
OR2_X1 U971 ( .A1(n1297), .A2(n1298), .ZN(n1168) );
NAND2_X1 U972 ( .A1(n1167), .A2(n1299), .ZN(n1296) );
XOR2_X1 U973 ( .A(n1300), .B(KEYINPUT32), .Z(n1167) );
XOR2_X1 U974 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U975 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U976 ( .A(G137), .B(n1305), .ZN(n1304) );
XOR2_X1 U977 ( .A(KEYINPUT28), .B(G146), .Z(n1303) );
XOR2_X1 U978 ( .A(n1306), .B(n1307), .Z(n1301) );
XOR2_X1 U979 ( .A(n1308), .B(n1141), .Z(n1307) );
XNOR2_X1 U980 ( .A(n1309), .B(G125), .ZN(n1141) );
NOR2_X1 U981 ( .A1(KEYINPUT6), .A2(n1199), .ZN(n1308) );
XNOR2_X1 U982 ( .A(G119), .B(n1310), .ZN(n1306) );
AND3_X1 U983 ( .A1(G221), .A2(n1096), .A3(G234), .ZN(n1310) );
INV_X1 U984 ( .A(n1289), .ZN(n1294) );
XOR2_X1 U985 ( .A(G472), .B(n1311), .Z(n1289) );
NOR2_X1 U986 ( .A1(KEYINPUT49), .A2(n1118), .ZN(n1311) );
NAND2_X1 U987 ( .A1(n1312), .A2(n1299), .ZN(n1118) );
XOR2_X1 U988 ( .A(n1313), .B(n1191), .Z(n1312) );
XOR2_X1 U989 ( .A(n1314), .B(n1315), .Z(n1313) );
NOR2_X1 U990 ( .A1(KEYINPUT22), .A2(n1316), .ZN(n1315) );
XOR2_X1 U991 ( .A(KEYINPUT42), .B(n1189), .Z(n1316) );
XOR2_X1 U992 ( .A(n1202), .B(n1220), .Z(n1189) );
NAND2_X1 U993 ( .A1(n1317), .A2(n1187), .ZN(n1314) );
NAND2_X1 U994 ( .A1(G101), .A2(n1318), .ZN(n1187) );
XNOR2_X1 U995 ( .A(KEYINPUT7), .B(n1186), .ZN(n1317) );
OR2_X1 U996 ( .A1(G101), .A2(n1318), .ZN(n1186) );
NOR3_X1 U997 ( .A1(G237), .A2(G953), .A3(n1319), .ZN(n1318) );
INV_X1 U998 ( .A(G210), .ZN(n1319) );
AND3_X1 U999 ( .A1(n1087), .A2(n1259), .A3(n1239), .ZN(n1247) );
NOR2_X1 U1000 ( .A1(n1109), .A2(n1110), .ZN(n1239) );
NOR2_X1 U1001 ( .A1(n1320), .A2(n1321), .ZN(n1110) );
INV_X1 U1002 ( .A(n1279), .ZN(n1109) );
XOR2_X1 U1003 ( .A(n1120), .B(n1322), .Z(n1279) );
NOR2_X1 U1004 ( .A1(n1121), .A2(KEYINPUT58), .ZN(n1322) );
AND2_X1 U1005 ( .A1(G210), .A2(n1323), .ZN(n1121) );
XOR2_X1 U1006 ( .A(KEYINPUT1), .B(n1321), .Z(n1323) );
NOR2_X1 U1007 ( .A1(G902), .A2(G237), .ZN(n1321) );
NAND2_X1 U1008 ( .A1(n1324), .A2(n1299), .ZN(n1120) );
XOR2_X1 U1009 ( .A(n1325), .B(n1326), .Z(n1324) );
XNOR2_X1 U1010 ( .A(n1220), .B(n1327), .ZN(n1326) );
XNOR2_X1 U1011 ( .A(G125), .B(KEYINPUT16), .ZN(n1327) );
AND2_X1 U1012 ( .A1(n1328), .A2(n1329), .ZN(n1220) );
NAND2_X1 U1013 ( .A1(n1330), .A2(n1305), .ZN(n1329) );
XNOR2_X1 U1014 ( .A(n1331), .B(n1332), .ZN(n1330) );
NAND2_X1 U1015 ( .A1(n1333), .A2(n1334), .ZN(n1328) );
XNOR2_X1 U1016 ( .A(KEYINPUT13), .B(n1305), .ZN(n1334) );
INV_X1 U1017 ( .A(G128), .ZN(n1305) );
XNOR2_X1 U1018 ( .A(G143), .B(n1332), .ZN(n1333) );
NOR2_X1 U1019 ( .A1(G146), .A2(KEYINPUT19), .ZN(n1332) );
XNOR2_X1 U1020 ( .A(n1222), .B(n1215), .ZN(n1325) );
AND2_X1 U1021 ( .A1(G224), .A2(n1096), .ZN(n1215) );
XOR2_X1 U1022 ( .A(n1158), .B(n1159), .Z(n1222) );
XNOR2_X1 U1023 ( .A(n1199), .B(n1335), .ZN(n1159) );
INV_X1 U1024 ( .A(G110), .ZN(n1199) );
XOR2_X1 U1025 ( .A(n1336), .B(n1191), .Z(n1158) );
XOR2_X1 U1026 ( .A(G113), .B(n1337), .Z(n1191) );
XNOR2_X1 U1027 ( .A(G119), .B(n1292), .ZN(n1337) );
XNOR2_X1 U1028 ( .A(G104), .B(n1338), .ZN(n1336) );
NAND2_X1 U1029 ( .A1(n1284), .A2(n1339), .ZN(n1259) );
NAND2_X1 U1030 ( .A1(n1286), .A2(n1156), .ZN(n1339) );
INV_X1 U1031 ( .A(G898), .ZN(n1156) );
NOR3_X1 U1032 ( .A1(n1299), .A2(n1068), .A3(n1096), .ZN(n1286) );
INV_X1 U1033 ( .A(n1101), .ZN(n1068) );
NAND3_X1 U1034 ( .A1(n1101), .A2(n1096), .A3(n1340), .ZN(n1284) );
XOR2_X1 U1035 ( .A(KEYINPUT31), .B(G952), .Z(n1340) );
INV_X1 U1036 ( .A(G953), .ZN(n1096) );
NAND2_X1 U1037 ( .A1(G237), .A2(n1341), .ZN(n1101) );
XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(n1342), .ZN(n1341) );
INV_X1 U1039 ( .A(n1282), .ZN(n1087) );
NAND2_X1 U1040 ( .A1(n1088), .A2(n1089), .ZN(n1282) );
NAND2_X1 U1041 ( .A1(G221), .A2(n1343), .ZN(n1089) );
XOR2_X1 U1042 ( .A(KEYINPUT2), .B(n1298), .Z(n1343) );
NOR2_X1 U1043 ( .A1(n1342), .A2(G902), .ZN(n1298) );
XNOR2_X1 U1044 ( .A(n1344), .B(G469), .ZN(n1088) );
NAND2_X1 U1045 ( .A1(n1345), .A2(n1299), .ZN(n1344) );
XOR2_X1 U1046 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1047 ( .A(n1348), .B(n1349), .Z(n1347) );
XNOR2_X1 U1048 ( .A(G110), .B(KEYINPUT48), .ZN(n1349) );
NAND2_X1 U1049 ( .A1(n1350), .A2(n1351), .ZN(n1348) );
NAND2_X1 U1050 ( .A1(n1207), .A2(n1145), .ZN(n1351) );
INV_X1 U1051 ( .A(n1206), .ZN(n1207) );
XOR2_X1 U1052 ( .A(n1352), .B(KEYINPUT53), .Z(n1350) );
NAND2_X1 U1053 ( .A1(n1209), .A2(n1206), .ZN(n1352) );
XNOR2_X1 U1054 ( .A(n1353), .B(n1338), .ZN(n1206) );
XOR2_X1 U1055 ( .A(G107), .B(G101), .Z(n1338) );
NAND2_X1 U1056 ( .A1(KEYINPUT10), .A2(n1354), .ZN(n1353) );
INV_X1 U1057 ( .A(G104), .ZN(n1354) );
INV_X1 U1058 ( .A(n1145), .ZN(n1209) );
XOR2_X1 U1059 ( .A(G128), .B(n1355), .Z(n1145) );
XOR2_X1 U1060 ( .A(n1196), .B(n1202), .Z(n1346) );
XOR2_X1 U1061 ( .A(n1149), .B(n1356), .Z(n1202) );
NOR2_X1 U1062 ( .A1(KEYINPUT8), .A2(n1147), .ZN(n1356) );
INV_X1 U1063 ( .A(n1357), .ZN(n1147) );
XOR2_X1 U1064 ( .A(G131), .B(G137), .Z(n1149) );
XNOR2_X1 U1065 ( .A(G140), .B(n1358), .ZN(n1196) );
NOR2_X1 U1066 ( .A1(G953), .A2(n1133), .ZN(n1358) );
INV_X1 U1067 ( .A(G227), .ZN(n1133) );
NOR2_X1 U1068 ( .A1(n1117), .A2(n1288), .ZN(n1098) );
INV_X1 U1069 ( .A(n1265), .ZN(n1288) );
XNOR2_X1 U1070 ( .A(n1122), .B(n1359), .ZN(n1265) );
NOR2_X1 U1071 ( .A1(G478), .A2(KEYINPUT60), .ZN(n1359) );
NAND2_X1 U1072 ( .A1(n1360), .A2(n1299), .ZN(n1122) );
XNOR2_X1 U1073 ( .A(KEYINPUT63), .B(n1173), .ZN(n1360) );
XOR2_X1 U1074 ( .A(n1361), .B(n1362), .Z(n1173) );
NOR3_X1 U1075 ( .A1(n1342), .A2(G953), .A3(n1297), .ZN(n1362) );
INV_X1 U1076 ( .A(G217), .ZN(n1297) );
INV_X1 U1077 ( .A(G234), .ZN(n1342) );
NAND2_X1 U1078 ( .A1(n1363), .A2(KEYINPUT25), .ZN(n1361) );
XOR2_X1 U1079 ( .A(n1364), .B(n1365), .Z(n1363) );
XOR2_X1 U1080 ( .A(n1366), .B(n1367), .Z(n1365) );
NAND2_X1 U1081 ( .A1(KEYINPUT47), .A2(n1292), .ZN(n1367) );
INV_X1 U1082 ( .A(G116), .ZN(n1292) );
NAND2_X1 U1083 ( .A1(n1368), .A2(n1369), .ZN(n1366) );
NAND2_X1 U1084 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XNOR2_X1 U1085 ( .A(n1372), .B(KEYINPUT35), .ZN(n1371) );
XNOR2_X1 U1086 ( .A(n1357), .B(KEYINPUT26), .ZN(n1370) );
XOR2_X1 U1087 ( .A(n1373), .B(KEYINPUT15), .Z(n1368) );
NAND2_X1 U1088 ( .A1(n1357), .A2(n1372), .ZN(n1373) );
XOR2_X1 U1089 ( .A(G128), .B(n1374), .Z(n1372) );
XNOR2_X1 U1090 ( .A(KEYINPUT34), .B(n1331), .ZN(n1374) );
INV_X1 U1091 ( .A(G143), .ZN(n1331) );
XOR2_X1 U1092 ( .A(G134), .B(KEYINPUT39), .Z(n1357) );
XNOR2_X1 U1093 ( .A(G107), .B(G122), .ZN(n1364) );
XOR2_X1 U1094 ( .A(G475), .B(n1375), .Z(n1117) );
AND2_X1 U1095 ( .A1(n1178), .A2(n1299), .ZN(n1375) );
INV_X1 U1096 ( .A(G902), .ZN(n1299) );
NAND2_X1 U1097 ( .A1(n1376), .A2(n1377), .ZN(n1178) );
NAND2_X1 U1098 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
XOR2_X1 U1099 ( .A(KEYINPUT12), .B(n1380), .Z(n1376) );
NOR2_X1 U1100 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
XNOR2_X1 U1101 ( .A(KEYINPUT56), .B(n1379), .ZN(n1382) );
XOR2_X1 U1102 ( .A(n1383), .B(n1384), .Z(n1379) );
XNOR2_X1 U1103 ( .A(n1355), .B(n1385), .ZN(n1384) );
NAND2_X1 U1104 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
NAND2_X1 U1105 ( .A1(n1388), .A2(n1309), .ZN(n1387) );
INV_X1 U1106 ( .A(G140), .ZN(n1309) );
XNOR2_X1 U1107 ( .A(KEYINPUT36), .B(n1218), .ZN(n1388) );
INV_X1 U1108 ( .A(G125), .ZN(n1218) );
NAND2_X1 U1109 ( .A1(G140), .A2(n1389), .ZN(n1386) );
XNOR2_X1 U1110 ( .A(G125), .B(KEYINPUT45), .ZN(n1389) );
XOR2_X1 U1111 ( .A(G143), .B(G146), .Z(n1355) );
XNOR2_X1 U1112 ( .A(G131), .B(n1390), .ZN(n1383) );
NOR3_X1 U1113 ( .A1(n1320), .A2(G953), .A3(G237), .ZN(n1390) );
INV_X1 U1114 ( .A(G214), .ZN(n1320) );
XOR2_X1 U1115 ( .A(n1378), .B(KEYINPUT37), .Z(n1381) );
XNOR2_X1 U1116 ( .A(G104), .B(n1391), .ZN(n1378) );
NOR2_X1 U1117 ( .A1(KEYINPUT41), .A2(n1392), .ZN(n1391) );
XNOR2_X1 U1118 ( .A(n1335), .B(G113), .ZN(n1392) );
INV_X1 U1119 ( .A(G122), .ZN(n1335) );
endmodule


