//Key = 0100000100101110110101110110001010110010101100010011000010111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448;

XOR2_X1 U797 ( .A(n1100), .B(n1101), .Z(G9) );
NOR2_X1 U798 ( .A1(n1102), .A2(n1103), .ZN(G75) );
XOR2_X1 U799 ( .A(n1104), .B(KEYINPUT7), .Z(n1103) );
NAND4_X1 U800 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1104) );
NAND4_X1 U801 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1107) );
NAND2_X1 U802 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U803 ( .A1(n1115), .A2(n1116), .A3(KEYINPUT41), .ZN(n1114) );
NAND2_X1 U804 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
NAND2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1106) );
NAND3_X1 U808 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
NAND2_X1 U809 ( .A1(KEYINPUT20), .A2(n1128), .ZN(n1127) );
NAND4_X1 U810 ( .A1(n1109), .A2(n1110), .A3(n1117), .A4(n1129), .ZN(n1128) );
NAND3_X1 U811 ( .A1(n1117), .A2(n1130), .A3(n1109), .ZN(n1126) );
NAND2_X1 U812 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND3_X1 U813 ( .A1(n1111), .A2(n1133), .A3(n1134), .ZN(n1132) );
INV_X1 U814 ( .A(n1135), .ZN(n1134) );
NAND2_X1 U815 ( .A1(n1110), .A2(n1136), .ZN(n1131) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
OR2_X1 U817 ( .A1(n1139), .A2(KEYINPUT20), .ZN(n1138) );
NAND2_X1 U818 ( .A1(n1111), .A2(n1140), .ZN(n1125) );
NAND3_X1 U819 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
NAND2_X1 U820 ( .A1(n1109), .A2(n1144), .ZN(n1142) );
NAND3_X1 U821 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
OR2_X1 U822 ( .A1(n1148), .A2(KEYINPUT3), .ZN(n1147) );
NAND3_X1 U823 ( .A1(n1110), .A2(n1149), .A3(n1115), .ZN(n1146) );
INV_X1 U824 ( .A(KEYINPUT41), .ZN(n1149) );
NAND2_X1 U825 ( .A1(n1117), .A2(n1150), .ZN(n1145) );
INV_X1 U826 ( .A(n1151), .ZN(n1109) );
NAND3_X1 U827 ( .A1(KEYINPUT3), .A2(n1152), .A3(n1151), .ZN(n1141) );
NOR3_X1 U828 ( .A1(n1153), .A2(G953), .A3(G952), .ZN(n1102) );
NOR3_X1 U829 ( .A1(n1143), .A2(n1116), .A3(n1154), .ZN(n1153) );
NAND3_X1 U830 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1143) );
AND2_X1 U831 ( .A1(n1158), .A2(n1135), .ZN(n1157) );
XOR2_X1 U832 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U833 ( .A1(n1161), .A2(KEYINPUT15), .ZN(n1160) );
XOR2_X1 U834 ( .A(n1162), .B(n1163), .Z(G72) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR3_X1 U836 ( .A1(n1166), .A2(KEYINPUT53), .A3(G953), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U838 ( .A(n1169), .B(KEYINPUT26), .Z(n1167) );
NAND2_X1 U839 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
NAND2_X1 U840 ( .A1(G900), .A2(G227), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1172), .A2(n1173), .ZN(n1162) );
NAND2_X1 U842 ( .A1(G953), .A2(n1174), .ZN(n1173) );
XOR2_X1 U843 ( .A(n1175), .B(n1176), .Z(n1172) );
XNOR2_X1 U844 ( .A(n1177), .B(n1178), .ZN(n1176) );
NAND2_X1 U845 ( .A1(n1179), .A2(n1180), .ZN(n1177) );
NAND2_X1 U846 ( .A1(G125), .A2(n1181), .ZN(n1180) );
XOR2_X1 U847 ( .A(KEYINPUT43), .B(n1182), .Z(n1179) );
NOR2_X1 U848 ( .A1(G125), .A2(n1181), .ZN(n1182) );
XOR2_X1 U849 ( .A(n1183), .B(G131), .Z(n1175) );
NAND2_X1 U850 ( .A1(KEYINPUT30), .A2(n1184), .ZN(n1183) );
XOR2_X1 U851 ( .A(n1185), .B(n1186), .Z(G69) );
XOR2_X1 U852 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND3_X1 U853 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1188) );
INV_X1 U854 ( .A(n1192), .ZN(n1190) );
NAND2_X1 U855 ( .A1(n1193), .A2(n1194), .ZN(n1189) );
NAND2_X1 U856 ( .A1(n1170), .A2(n1195), .ZN(n1187) );
NAND2_X1 U857 ( .A1(G898), .A2(G224), .ZN(n1195) );
XOR2_X1 U858 ( .A(G953), .B(KEYINPUT6), .Z(n1170) );
NOR2_X1 U859 ( .A1(n1196), .A2(G953), .ZN(n1185) );
NOR2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U861 ( .A1(n1199), .A2(n1200), .ZN(G66) );
NOR3_X1 U862 ( .A1(n1159), .A2(n1201), .A3(n1202), .ZN(n1200) );
NOR3_X1 U863 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
NOR2_X1 U864 ( .A1(n1206), .A2(n1207), .ZN(n1201) );
NOR2_X1 U865 ( .A1(n1105), .A2(n1204), .ZN(n1206) );
INV_X1 U866 ( .A(G217), .ZN(n1204) );
NOR2_X1 U867 ( .A1(n1199), .A2(n1208), .ZN(G63) );
XOR2_X1 U868 ( .A(n1209), .B(n1210), .Z(n1208) );
NOR2_X1 U869 ( .A1(n1211), .A2(n1205), .ZN(n1210) );
INV_X1 U870 ( .A(G478), .ZN(n1211) );
NOR2_X1 U871 ( .A1(n1199), .A2(n1212), .ZN(G60) );
XNOR2_X1 U872 ( .A(n1213), .B(n1214), .ZN(n1212) );
NOR2_X1 U873 ( .A1(n1215), .A2(n1205), .ZN(n1214) );
INV_X1 U874 ( .A(G475), .ZN(n1215) );
XNOR2_X1 U875 ( .A(G104), .B(n1216), .ZN(G6) );
NOR2_X1 U876 ( .A1(n1199), .A2(n1217), .ZN(G57) );
XOR2_X1 U877 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U878 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U879 ( .A(n1222), .B(n1223), .Z(n1218) );
XOR2_X1 U880 ( .A(n1224), .B(n1225), .Z(n1223) );
NOR2_X1 U881 ( .A1(n1226), .A2(n1205), .ZN(n1225) );
INV_X1 U882 ( .A(G472), .ZN(n1226) );
NOR2_X1 U883 ( .A1(KEYINPUT33), .A2(n1227), .ZN(n1224) );
XOR2_X1 U884 ( .A(n1228), .B(n1229), .Z(n1227) );
NAND4_X1 U885 ( .A1(KEYINPUT16), .A2(G210), .A3(n1230), .A4(n1108), .ZN(n1229) );
NAND2_X1 U886 ( .A1(KEYINPUT58), .A2(n1231), .ZN(n1222) );
INV_X1 U887 ( .A(n1232), .ZN(n1231) );
NOR2_X1 U888 ( .A1(n1199), .A2(n1233), .ZN(G54) );
XOR2_X1 U889 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U890 ( .A(n1236), .B(n1237), .Z(n1235) );
NOR2_X1 U891 ( .A1(n1238), .A2(n1205), .ZN(n1237) );
INV_X1 U892 ( .A(G469), .ZN(n1238) );
NAND2_X1 U893 ( .A1(n1239), .A2(n1240), .ZN(n1236) );
NAND2_X1 U894 ( .A1(n1241), .A2(G140), .ZN(n1239) );
XNOR2_X1 U895 ( .A(n1242), .B(KEYINPUT29), .ZN(n1241) );
NOR2_X1 U896 ( .A1(n1199), .A2(n1243), .ZN(G51) );
XNOR2_X1 U897 ( .A(n1244), .B(n1245), .ZN(n1243) );
NOR2_X1 U898 ( .A1(n1246), .A2(n1205), .ZN(n1245) );
OR2_X1 U899 ( .A1(n1247), .A2(n1105), .ZN(n1205) );
NOR4_X1 U900 ( .A1(n1198), .A2(n1168), .A3(n1248), .A4(n1249), .ZN(n1105) );
INV_X1 U901 ( .A(n1169), .ZN(n1249) );
XOR2_X1 U902 ( .A(KEYINPUT39), .B(n1197), .Z(n1248) );
NAND4_X1 U903 ( .A1(n1250), .A2(n1216), .A3(n1251), .A4(n1101), .ZN(n1197) );
NAND3_X1 U904 ( .A1(n1117), .A2(n1252), .A3(n1253), .ZN(n1101) );
NAND4_X1 U905 ( .A1(n1254), .A2(n1253), .A3(n1117), .A4(n1255), .ZN(n1216) );
NAND2_X1 U906 ( .A1(n1256), .A2(n1255), .ZN(n1250) );
INV_X1 U907 ( .A(n1257), .ZN(n1256) );
NAND4_X1 U908 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1168) );
NOR4_X1 U909 ( .A1(n1262), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(n1261) );
NOR3_X1 U910 ( .A1(n1266), .A2(n1119), .A3(n1267), .ZN(n1265) );
INV_X1 U911 ( .A(n1268), .ZN(n1264) );
AND2_X1 U912 ( .A1(KEYINPUT47), .A2(n1269), .ZN(n1263) );
NOR3_X1 U913 ( .A1(KEYINPUT47), .A2(n1270), .A3(n1271), .ZN(n1262) );
NOR2_X1 U914 ( .A1(n1272), .A2(n1273), .ZN(n1260) );
NAND4_X1 U915 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1198) );
NAND2_X1 U916 ( .A1(n1152), .A2(n1278), .ZN(n1275) );
NAND3_X1 U917 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1278) );
NAND4_X1 U918 ( .A1(KEYINPUT28), .A2(n1254), .A3(n1282), .A4(n1119), .ZN(n1281) );
OR4_X1 U919 ( .A1(n1139), .A2(n1119), .A3(n1282), .A4(KEYINPUT1), .ZN(n1280) );
NAND2_X1 U920 ( .A1(KEYINPUT1), .A2(n1252), .ZN(n1279) );
INV_X1 U921 ( .A(n1283), .ZN(n1252) );
NAND2_X1 U922 ( .A1(n1284), .A2(n1285), .ZN(n1274) );
INV_X1 U923 ( .A(KEYINPUT28), .ZN(n1285) );
NOR2_X1 U924 ( .A1(n1108), .A2(G952), .ZN(n1199) );
XOR2_X1 U925 ( .A(n1286), .B(n1287), .Z(G48) );
NOR2_X1 U926 ( .A1(KEYINPUT48), .A2(n1169), .ZN(n1287) );
NAND3_X1 U927 ( .A1(n1288), .A2(n1289), .A3(n1254), .ZN(n1169) );
XNOR2_X1 U928 ( .A(G146), .B(KEYINPUT56), .ZN(n1286) );
NAND2_X1 U929 ( .A1(n1290), .A2(n1291), .ZN(G45) );
OR2_X1 U930 ( .A1(n1292), .A2(G143), .ZN(n1291) );
NAND2_X1 U931 ( .A1(n1293), .A2(G143), .ZN(n1290) );
NAND2_X1 U932 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
OR2_X1 U933 ( .A1(n1258), .A2(KEYINPUT60), .ZN(n1295) );
INV_X1 U934 ( .A(n1296), .ZN(n1258) );
NAND2_X1 U935 ( .A1(KEYINPUT60), .A2(n1292), .ZN(n1294) );
NAND2_X1 U936 ( .A1(KEYINPUT42), .A2(n1296), .ZN(n1292) );
NOR4_X1 U937 ( .A1(n1297), .A2(n1119), .A3(n1298), .A4(n1299), .ZN(n1296) );
XOR2_X1 U938 ( .A(n1181), .B(n1259), .Z(G42) );
NAND3_X1 U939 ( .A1(n1123), .A2(n1150), .A3(n1300), .ZN(n1259) );
NAND2_X1 U940 ( .A1(n1301), .A2(n1302), .ZN(G39) );
NAND2_X1 U941 ( .A1(G137), .A2(n1268), .ZN(n1302) );
XOR2_X1 U942 ( .A(KEYINPUT22), .B(n1303), .Z(n1301) );
NOR2_X1 U943 ( .A1(G137), .A2(n1268), .ZN(n1303) );
NAND3_X1 U944 ( .A1(n1111), .A2(n1123), .A3(n1288), .ZN(n1268) );
AND3_X1 U945 ( .A1(n1150), .A2(n1304), .A3(n1270), .ZN(n1288) );
INV_X1 U946 ( .A(n1116), .ZN(n1123) );
NAND2_X1 U947 ( .A1(n1305), .A2(n1306), .ZN(G36) );
NAND2_X1 U948 ( .A1(n1273), .A2(n1307), .ZN(n1306) );
NAND2_X1 U949 ( .A1(G134), .A2(n1308), .ZN(n1307) );
OR2_X1 U950 ( .A1(n1309), .A2(KEYINPUT38), .ZN(n1308) );
NAND3_X1 U951 ( .A1(n1310), .A2(n1311), .A3(KEYINPUT38), .ZN(n1305) );
NAND2_X1 U952 ( .A1(G134), .A2(n1309), .ZN(n1311) );
INV_X1 U953 ( .A(KEYINPUT19), .ZN(n1309) );
NAND2_X1 U954 ( .A1(KEYINPUT19), .A2(n1312), .ZN(n1310) );
NAND2_X1 U955 ( .A1(G134), .A2(n1313), .ZN(n1312) );
INV_X1 U956 ( .A(n1273), .ZN(n1313) );
NOR3_X1 U957 ( .A1(n1116), .A2(n1139), .A3(n1297), .ZN(n1273) );
INV_X1 U958 ( .A(n1129), .ZN(n1139) );
XOR2_X1 U959 ( .A(n1314), .B(n1272), .Z(G33) );
NOR3_X1 U960 ( .A1(n1137), .A2(n1116), .A3(n1297), .ZN(n1272) );
NAND4_X1 U961 ( .A1(n1315), .A2(n1150), .A3(n1316), .A4(n1304), .ZN(n1297) );
XOR2_X1 U962 ( .A(n1253), .B(KEYINPUT36), .Z(n1150) );
NAND2_X1 U963 ( .A1(n1122), .A2(n1317), .ZN(n1116) );
XOR2_X1 U964 ( .A(n1318), .B(KEYINPUT10), .Z(n1314) );
XOR2_X1 U965 ( .A(G128), .B(n1269), .Z(G30) );
NOR2_X1 U966 ( .A1(n1271), .A2(n1319), .ZN(n1269) );
NAND4_X1 U967 ( .A1(n1253), .A2(n1129), .A3(n1289), .A4(n1304), .ZN(n1271) );
XOR2_X1 U968 ( .A(n1320), .B(n1321), .Z(G3) );
NOR2_X1 U969 ( .A1(KEYINPUT57), .A2(n1228), .ZN(n1321) );
INV_X1 U970 ( .A(G101), .ZN(n1228) );
NOR3_X1 U971 ( .A1(n1257), .A2(n1322), .A3(n1323), .ZN(n1320) );
NOR2_X1 U972 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
INV_X1 U973 ( .A(KEYINPUT0), .ZN(n1325) );
NOR2_X1 U974 ( .A1(n1119), .A2(n1282), .ZN(n1324) );
NOR2_X1 U975 ( .A1(KEYINPUT0), .A2(n1255), .ZN(n1322) );
NAND4_X1 U976 ( .A1(n1111), .A2(n1253), .A3(n1315), .A4(n1316), .ZN(n1257) );
XOR2_X1 U977 ( .A(n1326), .B(n1327), .Z(G27) );
XOR2_X1 U978 ( .A(n1328), .B(KEYINPUT27), .Z(n1327) );
NAND3_X1 U979 ( .A1(n1300), .A2(n1110), .A3(n1329), .ZN(n1326) );
XOR2_X1 U980 ( .A(n1119), .B(KEYINPUT17), .Z(n1329) );
INV_X1 U981 ( .A(n1289), .ZN(n1119) );
INV_X1 U982 ( .A(n1266), .ZN(n1300) );
NAND3_X1 U983 ( .A1(n1254), .A2(n1304), .A3(n1115), .ZN(n1266) );
NAND2_X1 U984 ( .A1(n1151), .A2(n1330), .ZN(n1304) );
NAND4_X1 U985 ( .A1(G902), .A2(G953), .A3(n1331), .A4(n1174), .ZN(n1330) );
INV_X1 U986 ( .A(G900), .ZN(n1174) );
XNOR2_X1 U987 ( .A(n1276), .B(n1332), .ZN(G24) );
NOR2_X1 U988 ( .A1(KEYINPUT11), .A2(n1333), .ZN(n1332) );
NAND4_X1 U989 ( .A1(n1110), .A2(n1117), .A3(n1334), .A4(n1255), .ZN(n1276) );
NOR2_X1 U990 ( .A1(n1299), .A2(n1298), .ZN(n1334) );
NOR2_X1 U991 ( .A1(n1316), .A2(n1335), .ZN(n1117) );
XOR2_X1 U992 ( .A(n1336), .B(n1277), .Z(G21) );
NAND4_X1 U993 ( .A1(n1110), .A2(n1270), .A3(n1111), .A4(n1255), .ZN(n1277) );
INV_X1 U994 ( .A(n1319), .ZN(n1270) );
NAND2_X1 U995 ( .A1(n1335), .A2(n1316), .ZN(n1319) );
INV_X1 U996 ( .A(n1315), .ZN(n1335) );
XOR2_X1 U997 ( .A(G116), .B(n1337), .Z(G18) );
NOR2_X1 U998 ( .A1(n1283), .A2(n1148), .ZN(n1337) );
NAND2_X1 U999 ( .A1(n1129), .A2(n1255), .ZN(n1283) );
NOR2_X1 U1000 ( .A1(n1298), .A2(n1338), .ZN(n1129) );
XNOR2_X1 U1001 ( .A(n1339), .B(KEYINPUT13), .ZN(n1298) );
XOR2_X1 U1002 ( .A(n1284), .B(n1340), .Z(G15) );
NOR2_X1 U1003 ( .A1(KEYINPUT52), .A2(n1341), .ZN(n1340) );
AND3_X1 U1004 ( .A1(n1254), .A2(n1255), .A3(n1152), .ZN(n1284) );
INV_X1 U1005 ( .A(n1148), .ZN(n1152) );
NAND3_X1 U1006 ( .A1(n1315), .A2(n1316), .A3(n1110), .ZN(n1148) );
INV_X1 U1007 ( .A(n1267), .ZN(n1110) );
NAND2_X1 U1008 ( .A1(n1133), .A2(n1135), .ZN(n1267) );
XNOR2_X1 U1009 ( .A(n1155), .B(KEYINPUT59), .ZN(n1133) );
INV_X1 U1010 ( .A(n1137), .ZN(n1254) );
NAND2_X1 U1011 ( .A1(n1339), .A2(n1338), .ZN(n1137) );
INV_X1 U1012 ( .A(n1299), .ZN(n1338) );
XOR2_X1 U1013 ( .A(n1342), .B(n1251), .Z(G12) );
NAND4_X1 U1014 ( .A1(n1115), .A2(n1111), .A3(n1253), .A4(n1255), .ZN(n1251) );
AND2_X1 U1015 ( .A1(n1289), .A2(n1282), .ZN(n1255) );
NAND2_X1 U1016 ( .A1(n1151), .A2(n1343), .ZN(n1282) );
NAND3_X1 U1017 ( .A1(n1192), .A2(n1331), .A3(G902), .ZN(n1343) );
NOR2_X1 U1018 ( .A1(n1108), .A2(G898), .ZN(n1192) );
NAND3_X1 U1019 ( .A1(n1331), .A2(n1108), .A3(G952), .ZN(n1151) );
NAND2_X1 U1020 ( .A1(G237), .A2(G234), .ZN(n1331) );
NOR2_X1 U1021 ( .A1(n1122), .A2(n1121), .ZN(n1289) );
INV_X1 U1022 ( .A(n1317), .ZN(n1121) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1344), .ZN(n1317) );
XNOR2_X1 U1024 ( .A(n1345), .B(n1246), .ZN(n1122) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1344), .ZN(n1246) );
NAND2_X1 U1026 ( .A1(n1230), .A2(n1247), .ZN(n1344) );
NAND2_X1 U1027 ( .A1(n1244), .A2(n1247), .ZN(n1345) );
XNOR2_X1 U1028 ( .A(n1346), .B(n1347), .ZN(n1244) );
XOR2_X1 U1029 ( .A(n1348), .B(n1349), .Z(n1347) );
NAND3_X1 U1030 ( .A1(n1350), .A2(n1351), .A3(n1352), .ZN(n1348) );
OR2_X1 U1031 ( .A1(n1191), .A2(KEYINPUT2), .ZN(n1352) );
OR2_X1 U1032 ( .A1(n1194), .A2(n1193), .ZN(n1191) );
NAND2_X1 U1033 ( .A1(n1353), .A2(n1354), .ZN(n1194) );
INV_X1 U1034 ( .A(n1355), .ZN(n1353) );
NAND3_X1 U1035 ( .A1(n1355), .A2(KEYINPUT2), .A3(n1356), .ZN(n1351) );
NAND2_X1 U1036 ( .A1(n1193), .A2(n1357), .ZN(n1350) );
NAND2_X1 U1037 ( .A1(n1358), .A2(n1354), .ZN(n1357) );
NAND2_X1 U1038 ( .A1(n1359), .A2(n1360), .ZN(n1354) );
XNOR2_X1 U1039 ( .A(n1355), .B(KEYINPUT2), .ZN(n1358) );
NOR2_X1 U1040 ( .A1(n1360), .A2(n1359), .ZN(n1355) );
XNOR2_X1 U1041 ( .A(n1361), .B(G101), .ZN(n1359) );
NAND2_X1 U1042 ( .A1(n1362), .A2(KEYINPUT62), .ZN(n1361) );
XOR2_X1 U1043 ( .A(n1100), .B(n1363), .Z(n1362) );
XNOR2_X1 U1044 ( .A(n1364), .B(G113), .ZN(n1360) );
NAND2_X1 U1045 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NAND2_X1 U1046 ( .A1(G116), .A2(n1336), .ZN(n1366) );
XOR2_X1 U1047 ( .A(KEYINPUT32), .B(n1367), .Z(n1365) );
NOR2_X1 U1048 ( .A1(G116), .A2(n1336), .ZN(n1367) );
INV_X1 U1049 ( .A(n1356), .ZN(n1193) );
XOR2_X1 U1050 ( .A(n1368), .B(n1369), .Z(n1356) );
NOR2_X1 U1051 ( .A1(KEYINPUT45), .A2(G122), .ZN(n1369) );
XOR2_X1 U1052 ( .A(n1342), .B(KEYINPUT23), .Z(n1368) );
XOR2_X1 U1053 ( .A(n1328), .B(n1370), .Z(n1346) );
NOR2_X1 U1054 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
XOR2_X1 U1055 ( .A(KEYINPUT9), .B(G953), .Z(n1372) );
INV_X1 U1056 ( .A(G224), .ZN(n1371) );
AND2_X1 U1057 ( .A1(n1373), .A2(n1135), .ZN(n1253) );
NAND2_X1 U1058 ( .A1(G221), .A2(n1374), .ZN(n1135) );
XOR2_X1 U1059 ( .A(n1155), .B(KEYINPUT40), .Z(n1373) );
XOR2_X1 U1060 ( .A(n1375), .B(G469), .Z(n1155) );
NAND2_X1 U1061 ( .A1(n1376), .A2(n1247), .ZN(n1375) );
XOR2_X1 U1062 ( .A(n1234), .B(n1377), .Z(n1376) );
NOR2_X1 U1063 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
NOR2_X1 U1064 ( .A1(n1242), .A2(n1181), .ZN(n1379) );
XNOR2_X1 U1065 ( .A(n1342), .B(n1380), .ZN(n1242) );
INV_X1 U1066 ( .A(n1240), .ZN(n1378) );
NAND2_X1 U1067 ( .A1(n1381), .A2(n1181), .ZN(n1240) );
XOR2_X1 U1068 ( .A(G110), .B(n1380), .Z(n1381) );
AND2_X1 U1069 ( .A1(G227), .A2(n1108), .ZN(n1380) );
XOR2_X1 U1070 ( .A(n1382), .B(n1383), .Z(n1234) );
XOR2_X1 U1071 ( .A(n1100), .B(n1384), .Z(n1383) );
NAND2_X1 U1072 ( .A1(KEYINPUT35), .A2(n1385), .ZN(n1384) );
XNOR2_X1 U1073 ( .A(n1386), .B(n1178), .ZN(n1382) );
XNOR2_X1 U1074 ( .A(n1387), .B(n1388), .ZN(n1178) );
NOR2_X1 U1075 ( .A1(KEYINPUT4), .A2(n1389), .ZN(n1388) );
XNOR2_X1 U1076 ( .A(KEYINPUT50), .B(G143), .ZN(n1389) );
XOR2_X1 U1077 ( .A(G146), .B(n1390), .Z(n1387) );
INV_X1 U1078 ( .A(n1154), .ZN(n1111) );
NAND2_X1 U1079 ( .A1(n1299), .A2(n1339), .ZN(n1154) );
XOR2_X1 U1080 ( .A(n1391), .B(G478), .Z(n1339) );
NAND2_X1 U1081 ( .A1(n1392), .A2(n1247), .ZN(n1391) );
XOR2_X1 U1082 ( .A(n1209), .B(KEYINPUT21), .Z(n1392) );
XOR2_X1 U1083 ( .A(n1393), .B(n1394), .Z(n1209) );
XOR2_X1 U1084 ( .A(n1395), .B(n1396), .Z(n1394) );
XOR2_X1 U1085 ( .A(n1397), .B(n1398), .Z(n1396) );
NOR2_X1 U1086 ( .A1(KEYINPUT61), .A2(n1100), .ZN(n1398) );
INV_X1 U1087 ( .A(G107), .ZN(n1100) );
NAND2_X1 U1088 ( .A1(n1399), .A2(n1400), .ZN(n1397) );
NAND2_X1 U1089 ( .A1(G143), .A2(n1390), .ZN(n1400) );
XOR2_X1 U1090 ( .A(n1401), .B(KEYINPUT54), .Z(n1399) );
OR2_X1 U1091 ( .A1(n1390), .A2(G143), .ZN(n1401) );
NAND2_X1 U1092 ( .A1(G217), .A2(n1402), .ZN(n1395) );
XOR2_X1 U1093 ( .A(n1403), .B(n1404), .Z(n1393) );
XOR2_X1 U1094 ( .A(KEYINPUT25), .B(G134), .Z(n1404) );
XOR2_X1 U1095 ( .A(G116), .B(n1333), .Z(n1403) );
INV_X1 U1096 ( .A(G122), .ZN(n1333) );
XOR2_X1 U1097 ( .A(n1405), .B(G475), .Z(n1299) );
NAND2_X1 U1098 ( .A1(n1213), .A2(n1247), .ZN(n1405) );
XNOR2_X1 U1099 ( .A(n1406), .B(n1407), .ZN(n1213) );
XOR2_X1 U1100 ( .A(n1408), .B(n1409), .Z(n1407) );
XOR2_X1 U1101 ( .A(n1410), .B(n1411), .Z(n1409) );
NAND2_X1 U1102 ( .A1(KEYINPUT14), .A2(n1181), .ZN(n1410) );
XOR2_X1 U1103 ( .A(n1412), .B(n1413), .Z(n1408) );
NOR2_X1 U1104 ( .A1(KEYINPUT8), .A2(n1363), .ZN(n1413) );
INV_X1 U1105 ( .A(n1385), .ZN(n1363) );
XNOR2_X1 U1106 ( .A(G104), .B(KEYINPUT44), .ZN(n1385) );
NAND3_X1 U1107 ( .A1(n1230), .A2(n1108), .A3(G214), .ZN(n1412) );
INV_X1 U1108 ( .A(G237), .ZN(n1230) );
XOR2_X1 U1109 ( .A(n1414), .B(n1415), .Z(n1406) );
XOR2_X1 U1110 ( .A(G131), .B(G125), .Z(n1415) );
XOR2_X1 U1111 ( .A(n1341), .B(G122), .Z(n1414) );
NOR2_X1 U1112 ( .A1(n1316), .A2(n1315), .ZN(n1115) );
XNOR2_X1 U1113 ( .A(n1159), .B(n1161), .ZN(n1315) );
AND2_X1 U1114 ( .A1(n1416), .A2(n1374), .ZN(n1161) );
NAND2_X1 U1115 ( .A1(G234), .A2(n1247), .ZN(n1374) );
XOR2_X1 U1116 ( .A(KEYINPUT31), .B(G217), .Z(n1416) );
NOR2_X1 U1117 ( .A1(n1207), .A2(G902), .ZN(n1159) );
INV_X1 U1118 ( .A(n1203), .ZN(n1207) );
XOR2_X1 U1119 ( .A(n1417), .B(n1418), .Z(n1203) );
XOR2_X1 U1120 ( .A(KEYINPUT5), .B(G137), .Z(n1418) );
XOR2_X1 U1121 ( .A(n1419), .B(n1420), .Z(n1417) );
NOR2_X1 U1122 ( .A1(n1421), .A2(n1422), .ZN(n1420) );
XOR2_X1 U1123 ( .A(n1423), .B(KEYINPUT12), .Z(n1422) );
NAND3_X1 U1124 ( .A1(n1424), .A2(n1425), .A3(n1426), .ZN(n1423) );
XOR2_X1 U1125 ( .A(KEYINPUT55), .B(n1427), .Z(n1424) );
NOR2_X1 U1126 ( .A1(n1428), .A2(n1427), .ZN(n1421) );
XNOR2_X1 U1127 ( .A(n1429), .B(n1430), .ZN(n1427) );
XOR2_X1 U1128 ( .A(n1181), .B(n1431), .Z(n1430) );
NAND2_X1 U1129 ( .A1(KEYINPUT34), .A2(n1328), .ZN(n1431) );
INV_X1 U1130 ( .A(G125), .ZN(n1328) );
INV_X1 U1131 ( .A(G140), .ZN(n1181) );
NAND2_X1 U1132 ( .A1(KEYINPUT51), .A2(G146), .ZN(n1429) );
AND2_X1 U1133 ( .A1(n1425), .A2(n1426), .ZN(n1428) );
XOR2_X1 U1134 ( .A(n1432), .B(KEYINPUT24), .Z(n1426) );
NAND2_X1 U1135 ( .A1(G110), .A2(n1433), .ZN(n1432) );
XOR2_X1 U1136 ( .A(G128), .B(G119), .Z(n1433) );
NAND2_X1 U1137 ( .A1(n1434), .A2(n1342), .ZN(n1425) );
XOR2_X1 U1138 ( .A(n1336), .B(G128), .Z(n1434) );
NAND2_X1 U1139 ( .A1(n1402), .A2(G221), .ZN(n1419) );
AND2_X1 U1140 ( .A1(G234), .A2(n1108), .ZN(n1402) );
INV_X1 U1141 ( .A(G953), .ZN(n1108) );
INV_X1 U1142 ( .A(n1156), .ZN(n1316) );
XOR2_X1 U1143 ( .A(n1435), .B(G472), .Z(n1156) );
NAND2_X1 U1144 ( .A1(n1436), .A2(n1247), .ZN(n1435) );
INV_X1 U1145 ( .A(G902), .ZN(n1247) );
XOR2_X1 U1146 ( .A(n1437), .B(n1438), .Z(n1436) );
XOR2_X1 U1147 ( .A(n1220), .B(n1386), .Z(n1438) );
XOR2_X1 U1148 ( .A(n1221), .B(G101), .Z(n1386) );
XNOR2_X1 U1149 ( .A(n1318), .B(n1184), .ZN(n1221) );
XOR2_X1 U1150 ( .A(G134), .B(G137), .Z(n1184) );
INV_X1 U1151 ( .A(G131), .ZN(n1318) );
INV_X1 U1152 ( .A(n1349), .ZN(n1220) );
XOR2_X1 U1153 ( .A(n1390), .B(n1439), .Z(n1349) );
NOR2_X1 U1154 ( .A1(KEYINPUT18), .A2(n1440), .ZN(n1439) );
XNOR2_X1 U1155 ( .A(KEYINPUT50), .B(n1411), .ZN(n1440) );
XOR2_X1 U1156 ( .A(G146), .B(G143), .Z(n1411) );
INV_X1 U1157 ( .A(G128), .ZN(n1390) );
XNOR2_X1 U1158 ( .A(n1441), .B(n1442), .ZN(n1437) );
NOR2_X1 U1159 ( .A1(KEYINPUT46), .A2(n1232), .ZN(n1442) );
NAND2_X1 U1160 ( .A1(n1443), .A2(n1444), .ZN(n1232) );
OR2_X1 U1161 ( .A1(n1341), .A2(n1445), .ZN(n1444) );
XOR2_X1 U1162 ( .A(n1446), .B(KEYINPUT37), .Z(n1443) );
NAND2_X1 U1163 ( .A1(n1445), .A2(n1341), .ZN(n1446) );
INV_X1 U1164 ( .A(G113), .ZN(n1341) );
XNOR2_X1 U1165 ( .A(n1336), .B(n1447), .ZN(n1445) );
NOR2_X1 U1166 ( .A1(G116), .A2(KEYINPUT49), .ZN(n1447) );
INV_X1 U1167 ( .A(G119), .ZN(n1336) );
NOR4_X1 U1168 ( .A1(KEYINPUT63), .A2(G953), .A3(G237), .A4(n1448), .ZN(n1441) );
INV_X1 U1169 ( .A(G210), .ZN(n1448) );
INV_X1 U1170 ( .A(G110), .ZN(n1342) );
endmodule


