//Key = 0011110010101100010001101111000001001101010111110001001101010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379;

XNOR2_X1 U755 ( .A(G107), .B(n1048), .ZN(G9) );
NAND4_X1 U756 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(G75) );
NAND3_X1 U757 ( .A1(KEYINPUT32), .A2(n1053), .A3(n1054), .ZN(n1052) );
NAND2_X1 U758 ( .A1(G952), .A2(n1055), .ZN(n1051) );
NAND3_X1 U759 ( .A1(n1056), .A2(n1053), .A3(n1057), .ZN(n1055) );
XOR2_X1 U760 ( .A(KEYINPUT26), .B(n1058), .Z(n1056) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NOR2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR3_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1066) );
NOR3_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1071) );
NOR4_X1 U770 ( .A1(n1073), .A2(n1080), .A3(n1069), .A4(n1070), .ZN(n1061) );
NOR3_X1 U771 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U773 ( .A(KEYINPUT12), .B(n1086), .Z(n1085) );
NOR2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1082) );
XOR2_X1 U775 ( .A(KEYINPUT8), .B(n1086), .Z(n1088) );
NOR2_X1 U776 ( .A1(n1089), .A2(n1063), .ZN(n1081) );
NOR2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
OR2_X1 U779 ( .A1(n1053), .A2(KEYINPUT32), .ZN(n1049) );
NAND4_X1 U780 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1053) );
NOR4_X1 U781 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1070), .ZN(n1097) );
XOR2_X1 U782 ( .A(n1101), .B(n1102), .Z(n1098) );
XOR2_X1 U783 ( .A(KEYINPUT10), .B(G472), .Z(n1102) );
NOR2_X1 U784 ( .A1(n1073), .A2(n1103), .ZN(n1096) );
XOR2_X1 U785 ( .A(n1104), .B(n1105), .Z(n1095) );
XOR2_X1 U786 ( .A(KEYINPUT31), .B(G469), .Z(n1105) );
NOR2_X1 U787 ( .A1(n1106), .A2(KEYINPUT48), .ZN(n1104) );
XNOR2_X1 U788 ( .A(n1107), .B(n1108), .ZN(n1094) );
NAND2_X1 U789 ( .A1(KEYINPUT21), .A2(n1109), .ZN(n1108) );
XOR2_X1 U790 ( .A(n1110), .B(n1111), .Z(G72) );
XOR2_X1 U791 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U792 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1114) );
NAND2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1112) );
NAND2_X1 U795 ( .A1(n1117), .A2(G953), .ZN(n1116) );
XOR2_X1 U796 ( .A(n1118), .B(KEYINPUT49), .Z(n1117) );
XOR2_X1 U797 ( .A(n1119), .B(n1120), .Z(n1115) );
XOR2_X1 U798 ( .A(G125), .B(n1121), .Z(n1120) );
XOR2_X1 U799 ( .A(G140), .B(G131), .Z(n1121) );
XOR2_X1 U800 ( .A(n1122), .B(n1123), .Z(n1119) );
NOR2_X1 U801 ( .A1(n1124), .A2(G953), .ZN(n1110) );
XOR2_X1 U802 ( .A(n1125), .B(n1126), .Z(G69) );
NOR2_X1 U803 ( .A1(n1127), .A2(n1050), .ZN(n1126) );
AND2_X1 U804 ( .A1(G224), .A2(G898), .ZN(n1127) );
NAND2_X1 U805 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
NAND2_X1 U806 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
OR3_X1 U807 ( .A1(n1130), .A2(n1132), .A3(n1131), .ZN(n1128) );
AND2_X1 U808 ( .A1(n1050), .A2(n1133), .ZN(n1130) );
NAND3_X1 U809 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR3_X1 U810 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(G66) );
AND2_X1 U811 ( .A1(KEYINPUT51), .A2(n1140), .ZN(n1139) );
NOR3_X1 U812 ( .A1(KEYINPUT51), .A2(n1050), .A3(n1054), .ZN(n1138) );
INV_X1 U813 ( .A(G952), .ZN(n1054) );
XNOR2_X1 U814 ( .A(n1141), .B(n1142), .ZN(n1137) );
NOR2_X1 U815 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1145), .ZN(G63) );
NOR3_X1 U817 ( .A1(n1107), .A2(n1146), .A3(n1147), .ZN(n1145) );
AND4_X1 U818 ( .A1(n1148), .A2(KEYINPUT59), .A3(G478), .A4(n1149), .ZN(n1147) );
NOR2_X1 U819 ( .A1(n1150), .A2(n1148), .ZN(n1146) );
NOR3_X1 U820 ( .A1(n1151), .A2(n1057), .A3(n1109), .ZN(n1150) );
INV_X1 U821 ( .A(KEYINPUT59), .ZN(n1151) );
NOR2_X1 U822 ( .A1(n1140), .A2(n1152), .ZN(G60) );
NOR2_X1 U823 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U824 ( .A(KEYINPUT50), .B(n1155), .Z(n1154) );
NOR2_X1 U825 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
INV_X1 U826 ( .A(n1158), .ZN(n1157) );
XOR2_X1 U827 ( .A(n1159), .B(KEYINPUT37), .Z(n1156) );
NOR2_X1 U828 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
NAND2_X1 U829 ( .A1(n1149), .A2(G475), .ZN(n1159) );
XNOR2_X1 U830 ( .A(n1160), .B(n1161), .ZN(G6) );
NOR2_X1 U831 ( .A1(KEYINPUT61), .A2(n1162), .ZN(n1161) );
NOR2_X1 U832 ( .A1(n1140), .A2(n1163), .ZN(G57) );
XOR2_X1 U833 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U834 ( .A(n1166), .B(n1167), .Z(n1165) );
AND2_X1 U835 ( .A1(G472), .A2(n1149), .ZN(n1167) );
NOR2_X1 U836 ( .A1(KEYINPUT6), .A2(n1168), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U838 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U839 ( .A1(KEYINPUT9), .A2(n1173), .ZN(n1172) );
XOR2_X1 U840 ( .A(n1174), .B(KEYINPUT17), .Z(n1169) );
NOR2_X1 U841 ( .A1(n1140), .A2(n1175), .ZN(G54) );
XOR2_X1 U842 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U843 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U844 ( .A(n1180), .B(n1174), .Z(n1179) );
XOR2_X1 U845 ( .A(KEYINPUT13), .B(n1181), .Z(n1178) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1176) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U848 ( .A1(n1186), .A2(n1144), .ZN(n1185) );
NOR2_X1 U849 ( .A1(n1187), .A2(n1188), .ZN(n1184) );
XOR2_X1 U850 ( .A(KEYINPUT30), .B(n1189), .Z(n1188) );
AND2_X1 U851 ( .A1(n1190), .A2(G140), .ZN(n1189) );
NOR2_X1 U852 ( .A1(G140), .A2(n1190), .ZN(n1187) );
NAND2_X1 U853 ( .A1(KEYINPUT27), .A2(n1191), .ZN(n1182) );
NOR2_X1 U854 ( .A1(n1140), .A2(n1192), .ZN(G51) );
XOR2_X1 U855 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U856 ( .A1(n1195), .A2(n1144), .ZN(n1194) );
INV_X1 U857 ( .A(n1149), .ZN(n1144) );
NOR2_X1 U858 ( .A1(n1196), .A2(n1057), .ZN(n1149) );
AND4_X1 U859 ( .A1(n1124), .A2(n1136), .A3(n1197), .A4(n1135), .ZN(n1057) );
XOR2_X1 U860 ( .A(KEYINPUT56), .B(n1134), .Z(n1197) );
AND4_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1134) );
NAND3_X1 U862 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1199) );
XOR2_X1 U863 ( .A(n1063), .B(KEYINPUT57), .Z(n1204) );
NAND4_X1 U864 ( .A1(n1205), .A2(n1091), .A3(n1206), .A4(n1207), .ZN(n1198) );
OR2_X1 U865 ( .A1(n1202), .A2(KEYINPUT15), .ZN(n1207) );
NAND2_X1 U866 ( .A1(KEYINPUT15), .A2(n1208), .ZN(n1206) );
NAND3_X1 U867 ( .A1(n1209), .A2(n1069), .A3(n1210), .ZN(n1208) );
INV_X1 U868 ( .A(n1078), .ZN(n1069) );
AND3_X1 U869 ( .A1(n1211), .A2(n1048), .A3(n1160), .ZN(n1136) );
NAND3_X1 U870 ( .A1(n1212), .A2(n1086), .A3(n1205), .ZN(n1160) );
NAND3_X1 U871 ( .A1(n1086), .A2(n1213), .A3(n1212), .ZN(n1048) );
INV_X1 U872 ( .A(n1065), .ZN(n1086) );
AND4_X1 U873 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1124) );
NOR4_X1 U874 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
NOR2_X1 U875 ( .A1(n1222), .A2(n1223), .ZN(n1216) );
NOR2_X1 U876 ( .A1(KEYINPUT0), .A2(n1224), .ZN(n1193) );
XOR2_X1 U877 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U878 ( .A(n1227), .B(n1171), .Z(n1226) );
XNOR2_X1 U879 ( .A(n1228), .B(n1229), .ZN(n1225) );
NOR2_X1 U880 ( .A1(G125), .A2(KEYINPUT14), .ZN(n1229) );
NOR3_X1 U881 ( .A1(n1230), .A2(KEYINPUT20), .A3(G953), .ZN(n1228) );
NOR2_X1 U882 ( .A1(n1050), .A2(G952), .ZN(n1140) );
XOR2_X1 U883 ( .A(G146), .B(n1223), .Z(G48) );
AND3_X1 U884 ( .A1(n1074), .A2(n1093), .A3(n1231), .ZN(n1223) );
XOR2_X1 U885 ( .A(G143), .B(n1222), .Z(G45) );
AND4_X1 U886 ( .A1(n1100), .A2(n1232), .A3(n1091), .A4(n1233), .ZN(n1222) );
NOR3_X1 U887 ( .A1(n1234), .A2(n1235), .A3(n1068), .ZN(n1233) );
INV_X1 U888 ( .A(n1236), .ZN(n1100) );
XNOR2_X1 U889 ( .A(G140), .B(n1214), .ZN(G42) );
NAND4_X1 U890 ( .A1(n1237), .A2(n1205), .A3(n1238), .A4(n1099), .ZN(n1214) );
XOR2_X1 U891 ( .A(G137), .B(n1221), .Z(G39) );
AND3_X1 U892 ( .A1(n1203), .A2(n1237), .A3(n1239), .ZN(n1221) );
XOR2_X1 U893 ( .A(G134), .B(n1220), .Z(G36) );
AND3_X1 U894 ( .A1(n1213), .A2(n1091), .A3(n1237), .ZN(n1220) );
XNOR2_X1 U895 ( .A(n1219), .B(n1240), .ZN(G33) );
XOR2_X1 U896 ( .A(KEYINPUT2), .B(G131), .Z(n1240) );
AND3_X1 U897 ( .A1(n1205), .A2(n1091), .A3(n1237), .ZN(n1219) );
NOR4_X1 U898 ( .A1(n1070), .A2(n1235), .A3(n1241), .A4(n1073), .ZN(n1237) );
INV_X1 U899 ( .A(n1079), .ZN(n1073) );
XOR2_X1 U900 ( .A(n1242), .B(n1215), .Z(G30) );
NAND4_X1 U901 ( .A1(n1203), .A2(n1213), .A3(n1243), .A4(n1210), .ZN(n1215) );
NOR2_X1 U902 ( .A1(n1241), .A2(n1235), .ZN(n1243) );
INV_X1 U903 ( .A(n1087), .ZN(n1213) );
XNOR2_X1 U904 ( .A(G101), .B(n1211), .ZN(G3) );
NAND3_X1 U905 ( .A1(n1212), .A2(n1091), .A3(n1239), .ZN(n1211) );
XOR2_X1 U906 ( .A(G125), .B(n1218), .Z(G27) );
AND3_X1 U907 ( .A1(n1231), .A2(n1238), .A3(n1078), .ZN(n1218) );
NOR4_X1 U908 ( .A1(n1084), .A2(n1068), .A3(n1092), .A4(n1241), .ZN(n1231) );
INV_X1 U909 ( .A(n1232), .ZN(n1241) );
NAND2_X1 U910 ( .A1(n1060), .A2(n1244), .ZN(n1232) );
NAND4_X1 U911 ( .A1(G902), .A2(G953), .A3(n1245), .A4(n1118), .ZN(n1244) );
INV_X1 U912 ( .A(G900), .ZN(n1118) );
NAND2_X1 U913 ( .A1(n1246), .A2(n1247), .ZN(G24) );
NAND2_X1 U914 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U915 ( .A1(G122), .A2(n1250), .ZN(n1246) );
NAND2_X1 U916 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U917 ( .A1(KEYINPUT16), .A2(n1253), .ZN(n1252) );
OR2_X1 U918 ( .A1(n1248), .A2(KEYINPUT16), .ZN(n1251) );
NOR2_X1 U919 ( .A1(KEYINPUT62), .A2(n1201), .ZN(n1248) );
INV_X1 U920 ( .A(n1253), .ZN(n1201) );
NOR4_X1 U921 ( .A1(n1234), .A2(n1254), .A3(n1065), .A4(n1236), .ZN(n1253) );
XOR2_X1 U922 ( .A(n1255), .B(KEYINPUT36), .Z(n1234) );
XOR2_X1 U923 ( .A(G119), .B(n1256), .Z(G21) );
NOR2_X1 U924 ( .A1(n1257), .A2(n1068), .ZN(n1256) );
XOR2_X1 U925 ( .A(n1258), .B(KEYINPUT60), .Z(n1257) );
NAND4_X1 U926 ( .A1(n1239), .A2(n1203), .A3(n1078), .A4(n1209), .ZN(n1258) );
NOR2_X1 U927 ( .A1(n1092), .A2(n1238), .ZN(n1203) );
XNOR2_X1 U928 ( .A(G116), .B(n1200), .ZN(G18) );
OR2_X1 U929 ( .A1(n1259), .A2(n1087), .ZN(n1200) );
NAND2_X1 U930 ( .A1(n1236), .A2(n1255), .ZN(n1087) );
XOR2_X1 U931 ( .A(n1260), .B(KEYINPUT7), .Z(n1255) );
XOR2_X1 U932 ( .A(G113), .B(n1261), .Z(G15) );
NOR2_X1 U933 ( .A1(n1084), .A2(n1259), .ZN(n1261) );
NAND2_X1 U934 ( .A1(n1202), .A2(n1091), .ZN(n1259) );
NAND2_X1 U935 ( .A1(n1262), .A2(n1263), .ZN(n1091) );
OR2_X1 U936 ( .A1(n1065), .A2(KEYINPUT24), .ZN(n1263) );
NAND2_X1 U937 ( .A1(n1238), .A2(n1092), .ZN(n1065) );
NAND3_X1 U938 ( .A1(n1092), .A2(n1093), .A3(KEYINPUT24), .ZN(n1262) );
INV_X1 U939 ( .A(n1254), .ZN(n1202) );
NAND3_X1 U940 ( .A1(n1210), .A2(n1209), .A3(n1078), .ZN(n1254) );
NOR2_X1 U941 ( .A1(n1076), .A2(n1103), .ZN(n1078) );
INV_X1 U942 ( .A(n1077), .ZN(n1103) );
INV_X1 U943 ( .A(n1205), .ZN(n1084) );
NOR2_X1 U944 ( .A1(n1260), .A2(n1236), .ZN(n1205) );
INV_X1 U945 ( .A(n1264), .ZN(n1260) );
NAND2_X1 U946 ( .A1(n1265), .A2(n1266), .ZN(G12) );
OR2_X1 U947 ( .A1(n1267), .A2(G110), .ZN(n1266) );
NAND2_X1 U948 ( .A1(n1268), .A2(G110), .ZN(n1265) );
NAND2_X1 U949 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
OR2_X1 U950 ( .A1(n1135), .A2(KEYINPUT41), .ZN(n1270) );
NAND2_X1 U951 ( .A1(KEYINPUT41), .A2(n1267), .ZN(n1269) );
NAND2_X1 U952 ( .A1(KEYINPUT25), .A2(n1271), .ZN(n1267) );
INV_X1 U953 ( .A(n1135), .ZN(n1271) );
NAND4_X1 U954 ( .A1(n1239), .A2(n1212), .A3(n1238), .A4(n1099), .ZN(n1135) );
INV_X1 U955 ( .A(n1092), .ZN(n1099) );
XNOR2_X1 U956 ( .A(n1272), .B(n1143), .ZN(n1092) );
NAND2_X1 U957 ( .A1(G217), .A2(n1273), .ZN(n1143) );
NAND2_X1 U958 ( .A1(n1141), .A2(n1196), .ZN(n1272) );
XNOR2_X1 U959 ( .A(n1274), .B(n1275), .ZN(n1141) );
XOR2_X1 U960 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U961 ( .A(n1278), .B(G125), .Z(n1277) );
INV_X1 U962 ( .A(G119), .ZN(n1278) );
NAND2_X1 U963 ( .A1(n1279), .A2(n1280), .ZN(n1276) );
NAND3_X1 U964 ( .A1(G137), .A2(G221), .A3(n1281), .ZN(n1280) );
XOR2_X1 U965 ( .A(n1282), .B(KEYINPUT40), .Z(n1279) );
NAND2_X1 U966 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
INV_X1 U967 ( .A(G137), .ZN(n1284) );
XOR2_X1 U968 ( .A(KEYINPUT22), .B(n1285), .Z(n1283) );
AND2_X1 U969 ( .A1(G221), .A2(n1281), .ZN(n1285) );
INV_X1 U970 ( .A(n1286), .ZN(n1281) );
XNOR2_X1 U971 ( .A(n1287), .B(n1288), .ZN(n1274) );
INV_X1 U972 ( .A(n1093), .ZN(n1238) );
NAND2_X1 U973 ( .A1(n1289), .A2(n1290), .ZN(n1093) );
NAND2_X1 U974 ( .A1(G472), .A2(n1101), .ZN(n1290) );
XOR2_X1 U975 ( .A(KEYINPUT54), .B(n1291), .Z(n1289) );
NOR2_X1 U976 ( .A1(G472), .A2(n1101), .ZN(n1291) );
NAND2_X1 U977 ( .A1(n1292), .A2(n1196), .ZN(n1101) );
XNOR2_X1 U978 ( .A(n1293), .B(n1164), .ZN(n1292) );
XNOR2_X1 U979 ( .A(n1294), .B(G101), .ZN(n1164) );
NAND2_X1 U980 ( .A1(n1295), .A2(G210), .ZN(n1294) );
NAND2_X1 U981 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
NAND2_X1 U982 ( .A1(n1173), .A2(n1298), .ZN(n1297) );
XOR2_X1 U983 ( .A(n1299), .B(KEYINPUT34), .Z(n1296) );
OR2_X1 U984 ( .A1(n1298), .A2(n1173), .ZN(n1299) );
NAND2_X1 U985 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
NAND2_X1 U986 ( .A1(n1302), .A2(n1171), .ZN(n1301) );
XOR2_X1 U987 ( .A(KEYINPUT44), .B(n1303), .Z(n1300) );
NOR2_X1 U988 ( .A1(n1302), .A2(n1171), .ZN(n1303) );
INV_X1 U989 ( .A(n1174), .ZN(n1302) );
AND3_X1 U990 ( .A1(n1074), .A2(n1209), .A3(n1210), .ZN(n1212) );
INV_X1 U991 ( .A(n1068), .ZN(n1210) );
NAND2_X1 U992 ( .A1(n1070), .A2(n1079), .ZN(n1068) );
NAND2_X1 U993 ( .A1(G214), .A2(n1304), .ZN(n1079) );
XOR2_X1 U994 ( .A(n1305), .B(n1195), .Z(n1070) );
NAND2_X1 U995 ( .A1(G210), .A2(n1304), .ZN(n1195) );
NAND2_X1 U996 ( .A1(n1306), .A2(n1196), .ZN(n1304) );
INV_X1 U997 ( .A(G237), .ZN(n1306) );
NAND3_X1 U998 ( .A1(n1307), .A2(n1308), .A3(n1196), .ZN(n1305) );
OR2_X1 U999 ( .A1(n1227), .A2(n1309), .ZN(n1308) );
NAND2_X1 U1000 ( .A1(n1227), .A2(n1310), .ZN(n1307) );
NAND2_X1 U1001 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND2_X1 U1002 ( .A1(KEYINPUT45), .A2(n1309), .ZN(n1312) );
OR2_X1 U1003 ( .A1(KEYINPUT28), .A2(n1313), .ZN(n1309) );
OR2_X1 U1004 ( .A1(n1313), .A2(KEYINPUT45), .ZN(n1311) );
XNOR2_X1 U1005 ( .A(n1314), .B(n1171), .ZN(n1313) );
XNOR2_X1 U1006 ( .A(n1287), .B(n1315), .ZN(n1171) );
NOR2_X1 U1007 ( .A1(G143), .A2(KEYINPUT29), .ZN(n1315) );
XOR2_X1 U1008 ( .A(n1316), .B(n1317), .Z(n1314) );
NOR2_X1 U1009 ( .A1(G953), .A2(n1230), .ZN(n1317) );
INV_X1 U1010 ( .A(G224), .ZN(n1230) );
XNOR2_X1 U1011 ( .A(n1131), .B(KEYINPUT55), .ZN(n1227) );
XOR2_X1 U1012 ( .A(n1318), .B(n1319), .Z(n1131) );
XOR2_X1 U1013 ( .A(n1320), .B(n1173), .Z(n1319) );
XNOR2_X1 U1014 ( .A(G113), .B(n1321), .ZN(n1173) );
XOR2_X1 U1015 ( .A(G119), .B(G116), .Z(n1321) );
NAND2_X1 U1016 ( .A1(KEYINPUT3), .A2(n1190), .ZN(n1320) );
INV_X1 U1017 ( .A(G110), .ZN(n1190) );
XOR2_X1 U1018 ( .A(n1322), .B(n1323), .Z(n1318) );
XOR2_X1 U1019 ( .A(G122), .B(G101), .Z(n1323) );
NAND3_X1 U1020 ( .A1(n1324), .A2(n1325), .A3(n1326), .ZN(n1322) );
NAND2_X1 U1021 ( .A1(KEYINPUT23), .A2(n1327), .ZN(n1326) );
NAND3_X1 U1022 ( .A1(n1328), .A2(n1329), .A3(n1162), .ZN(n1325) );
INV_X1 U1023 ( .A(KEYINPUT23), .ZN(n1329) );
OR2_X1 U1024 ( .A1(n1162), .A2(n1328), .ZN(n1324) );
NOR2_X1 U1025 ( .A1(KEYINPUT52), .A2(n1327), .ZN(n1328) );
NAND2_X1 U1026 ( .A1(n1060), .A2(n1330), .ZN(n1209) );
NAND3_X1 U1027 ( .A1(n1132), .A2(n1245), .A3(G902), .ZN(n1330) );
NOR2_X1 U1028 ( .A1(n1050), .A2(G898), .ZN(n1132) );
NAND3_X1 U1029 ( .A1(n1245), .A2(n1050), .A3(G952), .ZN(n1060) );
NAND2_X1 U1030 ( .A1(G237), .A2(G234), .ZN(n1245) );
INV_X1 U1031 ( .A(n1235), .ZN(n1074) );
NAND2_X1 U1032 ( .A1(n1076), .A2(n1077), .ZN(n1235) );
NAND2_X1 U1033 ( .A1(G221), .A2(n1273), .ZN(n1077) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1196), .ZN(n1273) );
XOR2_X1 U1035 ( .A(n1186), .B(n1331), .Z(n1076) );
NOR2_X1 U1036 ( .A1(n1106), .A2(KEYINPUT18), .ZN(n1331) );
AND3_X1 U1037 ( .A1(n1332), .A2(n1196), .A3(n1333), .ZN(n1106) );
NAND2_X1 U1038 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XNOR2_X1 U1039 ( .A(KEYINPUT19), .B(n1288), .ZN(n1335) );
XOR2_X1 U1040 ( .A(n1336), .B(KEYINPUT42), .Z(n1334) );
NAND2_X1 U1041 ( .A1(n1337), .A2(n1338), .ZN(n1332) );
XOR2_X1 U1042 ( .A(KEYINPUT19), .B(n1288), .Z(n1338) );
XOR2_X1 U1043 ( .A(G110), .B(G140), .Z(n1288) );
XOR2_X1 U1044 ( .A(n1336), .B(KEYINPUT5), .Z(n1337) );
XOR2_X1 U1045 ( .A(n1339), .B(n1340), .Z(n1336) );
XOR2_X1 U1046 ( .A(n1341), .B(n1191), .Z(n1340) );
INV_X1 U1047 ( .A(n1122), .ZN(n1191) );
XNOR2_X1 U1048 ( .A(G143), .B(n1287), .ZN(n1122) );
XNOR2_X1 U1049 ( .A(n1242), .B(G146), .ZN(n1287) );
INV_X1 U1050 ( .A(G128), .ZN(n1242) );
NOR2_X1 U1051 ( .A1(KEYINPUT35), .A2(n1174), .ZN(n1341) );
NAND2_X1 U1052 ( .A1(n1342), .A2(n1343), .ZN(n1174) );
NAND2_X1 U1053 ( .A1(G131), .A2(n1123), .ZN(n1343) );
XOR2_X1 U1054 ( .A(n1344), .B(KEYINPUT1), .Z(n1342) );
OR2_X1 U1055 ( .A1(n1123), .A2(G131), .ZN(n1344) );
XOR2_X1 U1056 ( .A(G134), .B(G137), .Z(n1123) );
XOR2_X1 U1057 ( .A(n1180), .B(n1181), .Z(n1339) );
AND2_X1 U1058 ( .A1(n1345), .A2(G227), .ZN(n1181) );
XOR2_X1 U1059 ( .A(n1050), .B(KEYINPUT58), .Z(n1345) );
NAND2_X1 U1060 ( .A1(n1346), .A2(n1347), .ZN(n1180) );
NAND2_X1 U1061 ( .A1(n1348), .A2(G101), .ZN(n1347) );
XOR2_X1 U1062 ( .A(KEYINPUT63), .B(n1349), .Z(n1346) );
NOR2_X1 U1063 ( .A1(G101), .A2(n1348), .ZN(n1349) );
XOR2_X1 U1064 ( .A(n1162), .B(n1350), .Z(n1348) );
INV_X1 U1065 ( .A(G104), .ZN(n1162) );
INV_X1 U1066 ( .A(G469), .ZN(n1186) );
INV_X1 U1067 ( .A(n1063), .ZN(n1239) );
NAND2_X1 U1068 ( .A1(n1236), .A2(n1264), .ZN(n1063) );
XOR2_X1 U1069 ( .A(n1107), .B(n1109), .Z(n1264) );
INV_X1 U1070 ( .A(G478), .ZN(n1109) );
NOR2_X1 U1071 ( .A1(n1148), .A2(G902), .ZN(n1107) );
XNOR2_X1 U1072 ( .A(n1351), .B(n1352), .ZN(n1148) );
NOR3_X1 U1073 ( .A1(n1286), .A2(KEYINPUT38), .A3(n1353), .ZN(n1352) );
INV_X1 U1074 ( .A(G217), .ZN(n1353) );
NAND2_X1 U1075 ( .A1(n1354), .A2(n1050), .ZN(n1286) );
INV_X1 U1076 ( .A(G953), .ZN(n1050) );
XOR2_X1 U1077 ( .A(KEYINPUT53), .B(G234), .Z(n1354) );
NAND2_X1 U1078 ( .A1(n1355), .A2(n1356), .ZN(n1351) );
NAND2_X1 U1079 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
XOR2_X1 U1080 ( .A(KEYINPUT46), .B(n1359), .Z(n1355) );
NOR2_X1 U1081 ( .A1(n1358), .A2(n1357), .ZN(n1359) );
XOR2_X1 U1082 ( .A(n1350), .B(n1360), .Z(n1357) );
XOR2_X1 U1083 ( .A(n1361), .B(n1249), .Z(n1360) );
INV_X1 U1084 ( .A(G122), .ZN(n1249) );
NAND2_X1 U1085 ( .A1(KEYINPUT33), .A2(G116), .ZN(n1361) );
INV_X1 U1086 ( .A(n1327), .ZN(n1350) );
XNOR2_X1 U1087 ( .A(G107), .B(KEYINPUT4), .ZN(n1327) );
XOR2_X1 U1088 ( .A(G128), .B(n1362), .Z(n1358) );
XOR2_X1 U1089 ( .A(G143), .B(G134), .Z(n1362) );
XOR2_X1 U1090 ( .A(n1363), .B(G475), .Z(n1236) );
NAND2_X1 U1091 ( .A1(n1158), .A2(n1196), .ZN(n1363) );
INV_X1 U1092 ( .A(G902), .ZN(n1196) );
XOR2_X1 U1093 ( .A(n1364), .B(n1365), .Z(n1158) );
XOR2_X1 U1094 ( .A(G113), .B(n1366), .Z(n1365) );
XOR2_X1 U1095 ( .A(KEYINPUT43), .B(G122), .Z(n1366) );
XOR2_X1 U1096 ( .A(n1367), .B(G104), .Z(n1364) );
NAND2_X1 U1097 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
NAND2_X1 U1098 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1099 ( .A(KEYINPUT39), .B(n1372), .Z(n1368) );
NOR2_X1 U1100 ( .A1(n1370), .A2(n1371), .ZN(n1372) );
XOR2_X1 U1101 ( .A(n1373), .B(n1374), .Z(n1371) );
XOR2_X1 U1102 ( .A(G143), .B(G131), .Z(n1374) );
NAND2_X1 U1103 ( .A1(n1295), .A2(G214), .ZN(n1373) );
NOR2_X1 U1104 ( .A1(G953), .A2(G237), .ZN(n1295) );
XOR2_X1 U1105 ( .A(n1375), .B(n1376), .Z(n1370) );
NOR2_X1 U1106 ( .A1(G146), .A2(KEYINPUT11), .ZN(n1376) );
NAND2_X1 U1107 ( .A1(n1377), .A2(n1378), .ZN(n1375) );
NAND2_X1 U1108 ( .A1(G140), .A2(n1316), .ZN(n1378) );
XOR2_X1 U1109 ( .A(KEYINPUT47), .B(n1379), .Z(n1377) );
NOR2_X1 U1110 ( .A1(G140), .A2(n1316), .ZN(n1379) );
INV_X1 U1111 ( .A(G125), .ZN(n1316) );
endmodule


