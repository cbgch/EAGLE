//Key = 0111001010010111100101100110000010010101100011110010011101111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356;

XNOR2_X1 U756 ( .A(n1034), .B(n1035), .ZN(G9) );
NOR2_X1 U757 ( .A1(n1036), .A2(n1037), .ZN(G75) );
NOR4_X1 U758 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1037) );
NAND3_X1 U759 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1038) );
NAND2_X1 U760 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U761 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND4_X1 U762 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
NAND2_X1 U763 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
NAND2_X1 U764 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U765 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1053) );
NAND2_X1 U768 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U769 ( .A1(G214), .A2(n1065), .A3(n1066), .ZN(n1064) );
NAND3_X1 U770 ( .A1(n1061), .A2(n1067), .A3(n1055), .ZN(n1047) );
NAND2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U772 ( .A1(n1070), .A2(n1071), .A3(n1052), .ZN(n1069) );
OR2_X1 U773 ( .A1(n1051), .A2(n1049), .ZN(n1071) );
NAND3_X1 U774 ( .A1(n1072), .A2(n1073), .A3(n1051), .ZN(n1070) );
NAND2_X1 U775 ( .A1(n1074), .A2(n1049), .ZN(n1068) );
INV_X1 U776 ( .A(n1075), .ZN(n1045) );
NOR3_X1 U777 ( .A1(n1076), .A2(G953), .A3(n1077), .ZN(n1036) );
INV_X1 U778 ( .A(n1042), .ZN(n1077) );
NAND4_X1 U779 ( .A1(n1078), .A2(n1079), .A3(n1055), .A4(n1080), .ZN(n1042) );
NOR4_X1 U780 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1080) );
XOR2_X1 U781 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U782 ( .A1(G469), .A2(KEYINPUT36), .ZN(n1086) );
XOR2_X1 U783 ( .A(n1087), .B(n1088), .Z(n1083) );
NOR3_X1 U784 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1082) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
AND3_X1 U786 ( .A1(n1093), .A2(n1092), .A3(KEYINPUT61), .ZN(n1090) );
AND2_X1 U787 ( .A1(KEYINPUT63), .A2(n1094), .ZN(n1092) );
NOR2_X1 U788 ( .A1(KEYINPUT61), .A2(n1094), .ZN(n1089) );
XNOR2_X1 U789 ( .A(G478), .B(KEYINPUT24), .ZN(n1094) );
XOR2_X1 U790 ( .A(n1095), .B(n1096), .Z(n1079) );
NOR2_X1 U791 ( .A1(n1097), .A2(KEYINPUT5), .ZN(n1096) );
INV_X1 U792 ( .A(n1098), .ZN(n1097) );
XNOR2_X1 U793 ( .A(KEYINPUT18), .B(n1040), .ZN(n1076) );
XOR2_X1 U794 ( .A(n1099), .B(n1100), .Z(G72) );
NOR2_X1 U795 ( .A1(n1101), .A2(G953), .ZN(n1100) );
NAND2_X1 U796 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
NAND2_X1 U797 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
OR2_X1 U798 ( .A1(n1043), .A2(G227), .ZN(n1105) );
NAND2_X1 U799 ( .A1(G953), .A2(n1106), .ZN(n1102) );
NAND2_X1 U800 ( .A1(G900), .A2(n1107), .ZN(n1106) );
OR2_X1 U801 ( .A1(n1104), .A2(G227), .ZN(n1107) );
XNOR2_X1 U802 ( .A(n1108), .B(n1109), .ZN(n1104) );
XNOR2_X1 U803 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U804 ( .A1(G131), .A2(KEYINPUT4), .ZN(n1111) );
NAND2_X1 U805 ( .A1(KEYINPUT21), .A2(n1112), .ZN(n1110) );
XNOR2_X1 U806 ( .A(n1113), .B(n1114), .ZN(n1108) );
XOR2_X1 U807 ( .A(n1115), .B(n1116), .Z(G69) );
NOR2_X1 U808 ( .A1(n1117), .A2(n1043), .ZN(n1116) );
NOR2_X1 U809 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U810 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NAND3_X1 U811 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
NAND2_X1 U812 ( .A1(G953), .A2(n1119), .ZN(n1123) );
XOR2_X1 U813 ( .A(KEYINPUT37), .B(n1125), .Z(n1120) );
NOR3_X1 U814 ( .A1(n1122), .A2(G953), .A3(n1124), .ZN(n1125) );
XNOR2_X1 U815 ( .A(n1126), .B(n1127), .ZN(n1122) );
NAND2_X1 U816 ( .A1(KEYINPUT54), .A2(n1128), .ZN(n1126) );
NOR3_X1 U817 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(G66) );
AND3_X1 U818 ( .A1(KEYINPUT30), .A2(G953), .A3(G952), .ZN(n1131) );
NOR2_X1 U819 ( .A1(KEYINPUT30), .A2(n1132), .ZN(n1130) );
INV_X1 U820 ( .A(n1133), .ZN(n1132) );
XOR2_X1 U821 ( .A(n1134), .B(n1135), .Z(n1129) );
NOR2_X1 U822 ( .A1(n1098), .A2(n1136), .ZN(n1134) );
NOR2_X1 U823 ( .A1(n1133), .A2(n1137), .ZN(G63) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U825 ( .A1(n1140), .A2(n1136), .ZN(n1139) );
NAND2_X1 U826 ( .A1(KEYINPUT11), .A2(n1141), .ZN(n1138) );
NOR2_X1 U827 ( .A1(n1133), .A2(n1142), .ZN(G60) );
XNOR2_X1 U828 ( .A(n1143), .B(n1144), .ZN(n1142) );
NOR2_X1 U829 ( .A1(n1145), .A2(n1136), .ZN(n1144) );
XNOR2_X1 U830 ( .A(G104), .B(n1146), .ZN(G6) );
NAND4_X1 U831 ( .A1(n1147), .A2(n1148), .A3(n1061), .A4(n1149), .ZN(n1146) );
XNOR2_X1 U832 ( .A(KEYINPUT49), .B(n1150), .ZN(n1149) );
NOR2_X1 U833 ( .A1(n1133), .A2(n1151), .ZN(G57) );
XOR2_X1 U834 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U835 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U836 ( .A(n1156), .B(n1157), .Z(n1152) );
NOR2_X1 U837 ( .A1(KEYINPUT31), .A2(n1158), .ZN(n1157) );
XOR2_X1 U838 ( .A(n1159), .B(G101), .Z(n1158) );
NAND3_X1 U839 ( .A1(G472), .A2(n1160), .A3(n1161), .ZN(n1156) );
XNOR2_X1 U840 ( .A(G902), .B(KEYINPUT16), .ZN(n1161) );
NOR3_X1 U841 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(G54) );
AND2_X1 U842 ( .A1(n1133), .A2(KEYINPUT26), .ZN(n1164) );
NOR3_X1 U843 ( .A1(KEYINPUT26), .A2(n1043), .A3(n1040), .ZN(n1163) );
INV_X1 U844 ( .A(G952), .ZN(n1040) );
XOR2_X1 U845 ( .A(n1165), .B(n1166), .Z(n1162) );
XOR2_X1 U846 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U847 ( .A(n1169), .B(n1170), .Z(n1165) );
NOR2_X1 U848 ( .A1(KEYINPUT27), .A2(n1171), .ZN(n1170) );
NOR2_X1 U849 ( .A1(n1172), .A2(n1136), .ZN(n1169) );
NOR2_X1 U850 ( .A1(n1133), .A2(n1173), .ZN(G51) );
XOR2_X1 U851 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U852 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U853 ( .A1(KEYINPUT44), .A2(n1178), .ZN(n1176) );
XNOR2_X1 U854 ( .A(n1179), .B(n1180), .ZN(n1174) );
NOR2_X1 U855 ( .A1(n1181), .A2(n1136), .ZN(n1180) );
NAND2_X1 U856 ( .A1(G902), .A2(n1160), .ZN(n1136) );
NAND2_X1 U857 ( .A1(n1101), .A2(n1124), .ZN(n1160) );
INV_X1 U858 ( .A(n1041), .ZN(n1124) );
NAND4_X1 U859 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1041) );
NOR4_X1 U860 ( .A1(n1186), .A2(n1187), .A3(n1035), .A4(n1188), .ZN(n1185) );
NOR4_X1 U861 ( .A1(n1150), .A2(n1189), .A3(n1072), .A4(n1190), .ZN(n1035) );
NOR2_X1 U862 ( .A1(n1191), .A2(n1192), .ZN(n1184) );
NOR4_X1 U863 ( .A1(n1190), .A2(n1189), .A3(n1150), .A4(n1193), .ZN(n1192) );
XNOR2_X1 U864 ( .A(KEYINPUT57), .B(n1073), .ZN(n1193) );
INV_X1 U865 ( .A(n1061), .ZN(n1190) );
INV_X1 U866 ( .A(n1039), .ZN(n1101) );
NAND4_X1 U867 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1039) );
NOR4_X1 U868 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
INV_X1 U869 ( .A(n1202), .ZN(n1199) );
NOR4_X1 U870 ( .A1(n1203), .A2(n1204), .A3(n1057), .A4(n1073), .ZN(n1198) );
XNOR2_X1 U871 ( .A(n1055), .B(KEYINPUT38), .ZN(n1203) );
NOR3_X1 U872 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1196) );
NOR2_X1 U873 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
AND4_X1 U874 ( .A1(n1208), .A2(n1210), .A3(n1150), .A4(n1211), .ZN(n1206) );
INV_X1 U875 ( .A(KEYINPUT35), .ZN(n1208) );
AND3_X1 U876 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1205) );
INV_X1 U877 ( .A(n1215), .ZN(n1194) );
NOR2_X1 U878 ( .A1(n1043), .A2(G952), .ZN(n1133) );
XNOR2_X1 U879 ( .A(G146), .B(n1216), .ZN(G48) );
NAND4_X1 U880 ( .A1(KEYINPUT59), .A2(n1212), .A3(n1217), .A4(n1213), .ZN(n1216) );
NOR2_X1 U881 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XNOR2_X1 U882 ( .A(n1074), .B(KEYINPUT52), .ZN(n1219) );
XNOR2_X1 U883 ( .A(G143), .B(n1209), .ZN(G45) );
NAND2_X1 U884 ( .A1(n1210), .A2(n1214), .ZN(n1209) );
NOR4_X1 U885 ( .A1(n1057), .A2(n1063), .A3(n1078), .A4(n1220), .ZN(n1210) );
XNOR2_X1 U886 ( .A(n1221), .B(n1215), .ZN(G42) );
NOR3_X1 U887 ( .A1(n1222), .A2(n1213), .A3(n1223), .ZN(n1215) );
XNOR2_X1 U888 ( .A(G137), .B(n1195), .ZN(G39) );
NAND3_X1 U889 ( .A1(n1055), .A2(n1049), .A3(n1224), .ZN(n1195) );
NAND3_X1 U890 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(G36) );
NAND2_X1 U891 ( .A1(KEYINPUT12), .A2(G134), .ZN(n1227) );
NAND3_X1 U892 ( .A1(n1228), .A2(n1229), .A3(n1201), .ZN(n1226) );
NAND2_X1 U893 ( .A1(n1230), .A2(n1231), .ZN(n1225) );
INV_X1 U894 ( .A(n1201), .ZN(n1231) );
NOR4_X1 U895 ( .A1(n1057), .A2(n1204), .A3(n1232), .A4(n1072), .ZN(n1201) );
NAND2_X1 U896 ( .A1(n1233), .A2(n1229), .ZN(n1230) );
INV_X1 U897 ( .A(KEYINPUT12), .ZN(n1229) );
XNOR2_X1 U898 ( .A(KEYINPUT46), .B(n1228), .ZN(n1233) );
XOR2_X1 U899 ( .A(G131), .B(n1234), .Z(G33) );
NOR2_X1 U900 ( .A1(n1057), .A2(n1223), .ZN(n1234) );
NAND3_X1 U901 ( .A1(n1214), .A2(n1055), .A3(n1147), .ZN(n1223) );
INV_X1 U902 ( .A(n1232), .ZN(n1055) );
NAND2_X1 U903 ( .A1(n1066), .A2(n1235), .ZN(n1232) );
NAND2_X1 U904 ( .A1(G214), .A2(n1065), .ZN(n1235) );
INV_X1 U905 ( .A(n1236), .ZN(n1057) );
XNOR2_X1 U906 ( .A(G128), .B(n1237), .ZN(G30) );
NAND2_X1 U907 ( .A1(KEYINPUT1), .A2(n1200), .ZN(n1237) );
AND3_X1 U908 ( .A1(n1238), .A2(n1239), .A3(n1224), .ZN(n1200) );
NOR3_X1 U909 ( .A1(n1204), .A2(n1060), .A3(n1222), .ZN(n1224) );
INV_X1 U910 ( .A(n1214), .ZN(n1204) );
NOR2_X1 U911 ( .A1(n1150), .A2(n1218), .ZN(n1214) );
INV_X1 U912 ( .A(n1211), .ZN(n1218) );
INV_X1 U913 ( .A(n1074), .ZN(n1150) );
XNOR2_X1 U914 ( .A(n1191), .B(n1240), .ZN(G3) );
NAND2_X1 U915 ( .A1(KEYINPUT8), .A2(G101), .ZN(n1240) );
AND2_X1 U916 ( .A1(n1241), .A2(n1236), .ZN(n1191) );
XNOR2_X1 U917 ( .A(G125), .B(n1202), .ZN(G27) );
NAND3_X1 U918 ( .A1(n1212), .A2(n1211), .A3(n1242), .ZN(n1202) );
AND3_X1 U919 ( .A1(n1060), .A2(n1052), .A3(n1051), .ZN(n1242) );
NAND2_X1 U920 ( .A1(n1075), .A2(n1243), .ZN(n1211) );
NAND4_X1 U921 ( .A1(G953), .A2(G902), .A3(n1244), .A4(n1245), .ZN(n1243) );
INV_X1 U922 ( .A(G900), .ZN(n1245) );
NOR3_X1 U923 ( .A1(n1073), .A2(n1063), .A3(n1222), .ZN(n1212) );
INV_X1 U924 ( .A(n1239), .ZN(n1063) );
XNOR2_X1 U925 ( .A(n1246), .B(n1182), .ZN(G24) );
NAND4_X1 U926 ( .A1(n1247), .A2(n1061), .A3(n1248), .A4(n1249), .ZN(n1182) );
NOR2_X1 U927 ( .A1(n1059), .A2(n1213), .ZN(n1061) );
NAND2_X1 U928 ( .A1(KEYINPUT25), .A2(n1250), .ZN(n1246) );
XNOR2_X1 U929 ( .A(G119), .B(n1183), .ZN(G21) );
NAND4_X1 U930 ( .A1(n1059), .A2(n1247), .A3(n1213), .A4(n1049), .ZN(n1183) );
INV_X1 U931 ( .A(n1060), .ZN(n1213) );
XNOR2_X1 U932 ( .A(n1251), .B(n1187), .ZN(G18) );
AND3_X1 U933 ( .A1(n1236), .A2(n1238), .A3(n1247), .ZN(n1187) );
INV_X1 U934 ( .A(n1072), .ZN(n1238) );
NAND2_X1 U935 ( .A1(n1252), .A2(n1249), .ZN(n1072) );
XNOR2_X1 U936 ( .A(KEYINPUT13), .B(n1078), .ZN(n1252) );
XOR2_X1 U937 ( .A(G113), .B(n1186), .Z(G15) );
AND3_X1 U938 ( .A1(n1147), .A2(n1236), .A3(n1247), .ZN(n1186) );
AND3_X1 U939 ( .A1(n1051), .A2(n1052), .A3(n1148), .ZN(n1247) );
NOR2_X1 U940 ( .A1(n1060), .A2(n1059), .ZN(n1236) );
XOR2_X1 U941 ( .A(G110), .B(n1188), .Z(G12) );
AND3_X1 U942 ( .A1(n1059), .A2(n1060), .A3(n1241), .ZN(n1188) );
AND3_X1 U943 ( .A1(n1148), .A2(n1049), .A3(n1074), .ZN(n1241) );
NOR2_X1 U944 ( .A1(n1052), .A2(n1081), .ZN(n1074) );
INV_X1 U945 ( .A(n1051), .ZN(n1081) );
NAND2_X1 U946 ( .A1(G221), .A2(n1253), .ZN(n1051) );
NAND2_X1 U947 ( .A1(n1254), .A2(n1255), .ZN(n1052) );
NAND2_X1 U948 ( .A1(n1256), .A2(n1085), .ZN(n1255) );
NAND2_X1 U949 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U950 ( .A1(n1172), .A2(n1259), .ZN(n1258) );
INV_X1 U951 ( .A(G469), .ZN(n1172) );
INV_X1 U952 ( .A(KEYINPUT10), .ZN(n1257) );
NAND2_X1 U953 ( .A1(G469), .A2(n1260), .ZN(n1254) );
NAND2_X1 U954 ( .A1(n1259), .A2(n1261), .ZN(n1260) );
OR2_X1 U955 ( .A1(n1085), .A2(KEYINPUT10), .ZN(n1261) );
NAND4_X1 U956 ( .A1(n1262), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(n1085) );
NAND3_X1 U957 ( .A1(n1266), .A2(n1267), .A3(n1168), .ZN(n1265) );
INV_X1 U958 ( .A(KEYINPUT51), .ZN(n1267) );
OR2_X1 U959 ( .A1(n1168), .A2(n1266), .ZN(n1264) );
NOR2_X1 U960 ( .A1(KEYINPUT20), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U961 ( .A(n1269), .B(n1270), .ZN(n1168) );
XNOR2_X1 U962 ( .A(n1221), .B(G110), .ZN(n1270) );
INV_X1 U963 ( .A(G140), .ZN(n1221) );
NAND2_X1 U964 ( .A1(G227), .A2(n1043), .ZN(n1269) );
NAND2_X1 U965 ( .A1(KEYINPUT51), .A2(n1268), .ZN(n1262) );
XNOR2_X1 U966 ( .A(n1171), .B(n1167), .ZN(n1268) );
XNOR2_X1 U967 ( .A(n1271), .B(n1112), .ZN(n1171) );
XNOR2_X1 U968 ( .A(n1272), .B(n1273), .ZN(n1112) );
NOR2_X1 U969 ( .A1(G128), .A2(KEYINPUT42), .ZN(n1273) );
XNOR2_X1 U970 ( .A(G101), .B(n1274), .ZN(n1271) );
NOR2_X1 U971 ( .A1(KEYINPUT41), .A2(n1275), .ZN(n1274) );
NOR2_X1 U972 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XOR2_X1 U973 ( .A(KEYINPUT62), .B(n1278), .Z(n1277) );
NOR2_X1 U974 ( .A1(G107), .A2(n1279), .ZN(n1278) );
NOR2_X1 U975 ( .A1(G104), .A2(n1034), .ZN(n1276) );
INV_X1 U976 ( .A(KEYINPUT9), .ZN(n1259) );
NAND2_X1 U977 ( .A1(n1280), .A2(n1281), .ZN(n1049) );
OR2_X1 U978 ( .A1(n1073), .A2(KEYINPUT13), .ZN(n1281) );
INV_X1 U979 ( .A(n1147), .ZN(n1073) );
NOR2_X1 U980 ( .A1(n1249), .A2(n1078), .ZN(n1147) );
NAND3_X1 U981 ( .A1(n1078), .A2(n1220), .A3(KEYINPUT13), .ZN(n1280) );
INV_X1 U982 ( .A(n1249), .ZN(n1220) );
XOR2_X1 U983 ( .A(n1093), .B(n1140), .Z(n1249) );
INV_X1 U984 ( .A(G478), .ZN(n1140) );
NAND2_X1 U985 ( .A1(n1282), .A2(n1263), .ZN(n1093) );
XNOR2_X1 U986 ( .A(KEYINPUT14), .B(n1141), .ZN(n1282) );
XOR2_X1 U987 ( .A(n1283), .B(n1284), .Z(n1141) );
XNOR2_X1 U988 ( .A(n1251), .B(n1285), .ZN(n1284) );
XNOR2_X1 U989 ( .A(KEYINPUT60), .B(n1250), .ZN(n1285) );
INV_X1 U990 ( .A(G122), .ZN(n1250) );
XOR2_X1 U991 ( .A(n1286), .B(n1287), .Z(n1283) );
XNOR2_X1 U992 ( .A(n1288), .B(n1289), .ZN(n1287) );
NOR2_X1 U993 ( .A1(KEYINPUT56), .A2(n1290), .ZN(n1289) );
NOR3_X1 U994 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1290) );
NOR2_X1 U995 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NOR2_X1 U996 ( .A1(n1296), .A2(n1297), .ZN(n1294) );
INV_X1 U997 ( .A(KEYINPUT55), .ZN(n1297) );
XNOR2_X1 U998 ( .A(G134), .B(KEYINPUT22), .ZN(n1296) );
AND3_X1 U999 ( .A1(n1295), .A2(n1228), .A3(KEYINPUT55), .ZN(n1292) );
XOR2_X1 U1000 ( .A(n1298), .B(G128), .Z(n1295) );
NAND2_X1 U1001 ( .A1(KEYINPUT3), .A2(G143), .ZN(n1298) );
NOR2_X1 U1002 ( .A1(KEYINPUT55), .A2(n1228), .ZN(n1291) );
NAND2_X1 U1003 ( .A1(KEYINPUT15), .A2(n1034), .ZN(n1288) );
INV_X1 U1004 ( .A(G107), .ZN(n1034) );
NAND2_X1 U1005 ( .A1(G217), .A2(n1299), .ZN(n1286) );
INV_X1 U1006 ( .A(n1248), .ZN(n1078) );
XNOR2_X1 U1007 ( .A(n1300), .B(n1301), .ZN(n1248) );
XNOR2_X1 U1008 ( .A(KEYINPUT0), .B(n1145), .ZN(n1301) );
INV_X1 U1009 ( .A(G475), .ZN(n1145) );
NAND2_X1 U1010 ( .A1(n1143), .A2(n1263), .ZN(n1300) );
XNOR2_X1 U1011 ( .A(n1302), .B(n1303), .ZN(n1143) );
XOR2_X1 U1012 ( .A(n1304), .B(n1305), .Z(n1303) );
NAND2_X1 U1013 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1014 ( .A1(n1308), .A2(n1279), .ZN(n1307) );
XOR2_X1 U1015 ( .A(KEYINPUT39), .B(n1309), .Z(n1306) );
NOR2_X1 U1016 ( .A1(n1279), .A2(n1308), .ZN(n1309) );
XOR2_X1 U1017 ( .A(G113), .B(n1310), .Z(n1308) );
NOR2_X1 U1018 ( .A1(G122), .A2(KEYINPUT17), .ZN(n1310) );
NAND2_X1 U1019 ( .A1(n1311), .A2(n1312), .ZN(n1304) );
NAND2_X1 U1020 ( .A1(n1313), .A2(n1114), .ZN(n1312) );
XOR2_X1 U1021 ( .A(n1314), .B(KEYINPUT7), .Z(n1311) );
OR2_X1 U1022 ( .A1(n1114), .A2(n1313), .ZN(n1314) );
XNOR2_X1 U1023 ( .A(G146), .B(KEYINPUT32), .ZN(n1313) );
XOR2_X1 U1024 ( .A(n1315), .B(n1316), .Z(n1302) );
AND3_X1 U1025 ( .A1(G214), .A2(n1043), .A3(n1317), .ZN(n1316) );
XNOR2_X1 U1026 ( .A(G131), .B(G143), .ZN(n1315) );
INV_X1 U1027 ( .A(n1189), .ZN(n1148) );
NAND2_X1 U1028 ( .A1(n1239), .A2(n1318), .ZN(n1189) );
NAND2_X1 U1029 ( .A1(n1075), .A2(n1319), .ZN(n1318) );
NAND4_X1 U1030 ( .A1(G953), .A2(G902), .A3(n1244), .A4(n1119), .ZN(n1319) );
INV_X1 U1031 ( .A(G898), .ZN(n1119) );
NAND3_X1 U1032 ( .A1(n1244), .A2(n1043), .A3(G952), .ZN(n1075) );
NAND2_X1 U1033 ( .A1(G237), .A2(G234), .ZN(n1244) );
NOR2_X1 U1034 ( .A1(n1066), .A2(n1320), .ZN(n1239) );
AND2_X1 U1035 ( .A1(G214), .A2(n1065), .ZN(n1320) );
XNOR2_X1 U1036 ( .A(n1321), .B(n1181), .ZN(n1066) );
NAND2_X1 U1037 ( .A1(G210), .A2(n1065), .ZN(n1181) );
NAND2_X1 U1038 ( .A1(n1322), .A2(n1317), .ZN(n1065) );
NAND2_X1 U1039 ( .A1(n1323), .A2(n1263), .ZN(n1321) );
XOR2_X1 U1040 ( .A(n1177), .B(n1324), .Z(n1323) );
XOR2_X1 U1041 ( .A(n1325), .B(n1178), .Z(n1324) );
NOR2_X1 U1042 ( .A1(n1118), .A2(G953), .ZN(n1178) );
INV_X1 U1043 ( .A(G224), .ZN(n1118) );
NAND2_X1 U1044 ( .A1(KEYINPUT6), .A2(n1179), .ZN(n1325) );
XOR2_X1 U1045 ( .A(n1326), .B(n1327), .Z(n1177) );
XOR2_X1 U1046 ( .A(KEYINPUT19), .B(n1328), .Z(n1327) );
XOR2_X1 U1047 ( .A(n1127), .B(n1128), .Z(n1326) );
XNOR2_X1 U1048 ( .A(G110), .B(G122), .ZN(n1128) );
XNOR2_X1 U1049 ( .A(n1329), .B(n1330), .ZN(n1127) );
XNOR2_X1 U1050 ( .A(G107), .B(n1331), .ZN(n1330) );
NAND2_X1 U1051 ( .A1(KEYINPUT47), .A2(n1279), .ZN(n1331) );
INV_X1 U1052 ( .A(G104), .ZN(n1279) );
XOR2_X1 U1053 ( .A(n1332), .B(n1333), .Z(n1329) );
NAND2_X1 U1054 ( .A1(KEYINPUT2), .A2(n1251), .ZN(n1332) );
INV_X1 U1055 ( .A(G116), .ZN(n1251) );
NAND3_X1 U1056 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1060) );
OR2_X1 U1057 ( .A1(n1337), .A2(n1087), .ZN(n1336) );
NAND3_X1 U1058 ( .A1(n1338), .A2(n1337), .A3(n1088), .ZN(n1335) );
INV_X1 U1059 ( .A(KEYINPUT29), .ZN(n1337) );
OR2_X1 U1060 ( .A1(n1088), .A2(n1338), .ZN(n1334) );
AND2_X1 U1061 ( .A1(n1339), .A2(n1087), .ZN(n1338) );
NAND2_X1 U1062 ( .A1(n1340), .A2(n1263), .ZN(n1087) );
INV_X1 U1063 ( .A(G902), .ZN(n1263) );
XOR2_X1 U1064 ( .A(n1341), .B(n1342), .Z(n1340) );
XNOR2_X1 U1065 ( .A(KEYINPUT23), .B(n1159), .ZN(n1342) );
NAND3_X1 U1066 ( .A1(n1317), .A2(n1043), .A3(G210), .ZN(n1159) );
INV_X1 U1067 ( .A(G237), .ZN(n1317) );
XOR2_X1 U1068 ( .A(n1154), .B(n1333), .Z(n1341) );
XOR2_X1 U1069 ( .A(G101), .B(n1155), .Z(n1333) );
XOR2_X1 U1070 ( .A(G113), .B(G119), .Z(n1155) );
XOR2_X1 U1071 ( .A(n1343), .B(n1344), .Z(n1154) );
XOR2_X1 U1072 ( .A(KEYINPUT34), .B(n1345), .Z(n1344) );
NOR2_X1 U1073 ( .A1(G116), .A2(KEYINPUT43), .ZN(n1345) );
XNOR2_X1 U1074 ( .A(n1167), .B(n1328), .ZN(n1343) );
XOR2_X1 U1075 ( .A(G128), .B(n1272), .Z(n1328) );
XOR2_X1 U1076 ( .A(G143), .B(G146), .Z(n1272) );
XOR2_X1 U1077 ( .A(G131), .B(n1113), .Z(n1167) );
XNOR2_X1 U1078 ( .A(G137), .B(n1228), .ZN(n1113) );
INV_X1 U1079 ( .A(G134), .ZN(n1228) );
XNOR2_X1 U1080 ( .A(KEYINPUT48), .B(KEYINPUT28), .ZN(n1339) );
XOR2_X1 U1081 ( .A(G472), .B(KEYINPUT45), .Z(n1088) );
INV_X1 U1082 ( .A(n1222), .ZN(n1059) );
XOR2_X1 U1083 ( .A(n1346), .B(n1098), .Z(n1222) );
NAND2_X1 U1084 ( .A1(G217), .A2(n1253), .ZN(n1098) );
NAND2_X1 U1085 ( .A1(G234), .A2(n1322), .ZN(n1253) );
XNOR2_X1 U1086 ( .A(G902), .B(KEYINPUT33), .ZN(n1322) );
XNOR2_X1 U1087 ( .A(n1095), .B(KEYINPUT50), .ZN(n1346) );
NOR2_X1 U1088 ( .A1(n1135), .A2(G902), .ZN(n1095) );
XNOR2_X1 U1089 ( .A(n1347), .B(n1348), .ZN(n1135) );
XOR2_X1 U1090 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1091 ( .A(n1351), .B(G110), .Z(n1350) );
NAND2_X1 U1092 ( .A1(KEYINPUT58), .A2(G137), .ZN(n1351) );
XNOR2_X1 U1093 ( .A(G128), .B(G146), .ZN(n1349) );
XOR2_X1 U1094 ( .A(n1352), .B(n1353), .Z(n1347) );
NOR2_X1 U1095 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NOR2_X1 U1096 ( .A1(KEYINPUT40), .A2(G119), .ZN(n1355) );
AND2_X1 U1097 ( .A1(KEYINPUT53), .A2(G119), .ZN(n1354) );
XOR2_X1 U1098 ( .A(n1356), .B(n1114), .Z(n1352) );
XNOR2_X1 U1099 ( .A(G140), .B(n1179), .ZN(n1114) );
INV_X1 U1100 ( .A(G125), .ZN(n1179) );
NAND2_X1 U1101 ( .A1(n1299), .A2(G221), .ZN(n1356) );
AND2_X1 U1102 ( .A1(G234), .A2(n1043), .ZN(n1299) );
INV_X1 U1103 ( .A(G953), .ZN(n1043) );
endmodule


