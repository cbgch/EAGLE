//Key = 0000110001000111011000100011101000101111011110000101100110111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;

XOR2_X1 U731 ( .A(n1019), .B(n1020), .Z(G9) );
XOR2_X1 U732 ( .A(KEYINPUT48), .B(G107), .Z(n1020) );
NOR2_X1 U733 ( .A1(KEYINPUT12), .A2(n1021), .ZN(n1019) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
NAND2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1025) );
OR3_X1 U737 ( .A1(n1030), .A2(n1031), .A3(KEYINPUT41), .ZN(n1029) );
AND3_X1 U738 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND2_X1 U739 ( .A1(KEYINPUT41), .A2(n1030), .ZN(n1028) );
NAND2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1030) );
NAND4_X1 U741 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
NAND2_X1 U742 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U743 ( .A1(KEYINPUT51), .A2(n1043), .ZN(n1042) );
NAND3_X1 U744 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1039) );
OR3_X1 U745 ( .A1(n1047), .A2(KEYINPUT31), .A3(n1048), .ZN(n1045) );
NAND2_X1 U746 ( .A1(n1043), .A2(n1049), .ZN(n1044) );
INV_X1 U747 ( .A(KEYINPUT51), .ZN(n1049) );
XOR2_X1 U748 ( .A(n1050), .B(KEYINPUT54), .Z(n1043) );
NAND3_X1 U749 ( .A1(n1051), .A2(n1052), .A3(n1034), .ZN(n1035) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U751 ( .A1(KEYINPUT31), .A2(n1033), .ZN(n1054) );
NAND4_X1 U752 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1024) );
NAND2_X1 U753 ( .A1(n1037), .A2(n1059), .ZN(n1056) );
NAND2_X1 U754 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U755 ( .A1(n1038), .A2(n1046), .A3(n1062), .ZN(n1061) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1063), .ZN(n1060) );
AND3_X1 U757 ( .A1(n1051), .A2(n1033), .A3(n1064), .ZN(n1037) );
NAND2_X1 U758 ( .A1(n1034), .A2(n1065), .ZN(n1055) );
NAND2_X1 U759 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U760 ( .A1(n1033), .A2(n1068), .ZN(n1067) );
NAND2_X1 U761 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U762 ( .A1(KEYINPUT41), .A2(n1032), .ZN(n1070) );
NAND2_X1 U763 ( .A1(n1071), .A2(n1051), .ZN(n1066) );
AND4_X1 U764 ( .A1(n1064), .A2(n1050), .A3(n1038), .A4(n1046), .ZN(n1034) );
INV_X1 U765 ( .A(n1072), .ZN(n1064) );
NOR3_X1 U766 ( .A1(n1073), .A2(G953), .A3(G952), .ZN(n1022) );
INV_X1 U767 ( .A(n1057), .ZN(n1073) );
NAND4_X1 U768 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1057) );
NOR4_X1 U769 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
NOR2_X1 U770 ( .A1(G469), .A2(n1082), .ZN(n1079) );
XNOR2_X1 U771 ( .A(KEYINPUT36), .B(n1083), .ZN(n1082) );
AND2_X1 U772 ( .A1(n1083), .A2(G469), .ZN(n1078) );
NOR2_X1 U773 ( .A1(n1041), .A2(n1084), .ZN(n1076) );
INV_X1 U774 ( .A(n1048), .ZN(n1084) );
XOR2_X1 U775 ( .A(n1085), .B(n1086), .Z(n1075) );
NAND2_X1 U776 ( .A1(KEYINPUT17), .A2(n1087), .ZN(n1086) );
NAND2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(G72) );
NAND2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U779 ( .A(n1092), .B(KEYINPUT21), .Z(n1088) );
NAND2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U781 ( .A(KEYINPUT14), .B(n1090), .Z(n1094) );
XNOR2_X1 U782 ( .A(n1095), .B(n1096), .ZN(n1090) );
NOR2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U784 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U785 ( .A1(G900), .A2(n1058), .ZN(n1097) );
NAND2_X1 U786 ( .A1(n1058), .A2(n1027), .ZN(n1095) );
INV_X1 U787 ( .A(n1091), .ZN(n1093) );
NAND2_X1 U788 ( .A1(G953), .A2(n1101), .ZN(n1091) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1101) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(G69) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1026), .ZN(n1103) );
NOR2_X1 U792 ( .A1(n1105), .A2(n1058), .ZN(n1104) );
NOR2_X1 U793 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U794 ( .A(G224), .B(KEYINPUT11), .ZN(n1106) );
NAND3_X1 U795 ( .A1(n1108), .A2(n1109), .A3(KEYINPUT28), .ZN(n1102) );
XOR2_X1 U796 ( .A(KEYINPUT58), .B(n1110), .Z(n1109) );
NOR2_X1 U797 ( .A1(n1111), .A2(n1058), .ZN(n1110) );
XOR2_X1 U798 ( .A(n1107), .B(KEYINPUT44), .Z(n1111) );
XOR2_X1 U799 ( .A(n1112), .B(n1113), .Z(n1108) );
NOR2_X1 U800 ( .A1(KEYINPUT53), .A2(n1114), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XOR2_X1 U802 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND3_X1 U803 ( .A1(n1119), .A2(G217), .A3(KEYINPUT43), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1120), .ZN(G63) );
XNOR2_X1 U805 ( .A(n1121), .B(n1122), .ZN(n1120) );
AND2_X1 U806 ( .A1(G478), .A2(n1119), .ZN(n1122) );
NOR2_X1 U807 ( .A1(n1115), .A2(n1123), .ZN(G60) );
XOR2_X1 U808 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U809 ( .A1(n1119), .A2(G475), .ZN(n1124) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(G6) );
NAND3_X1 U811 ( .A1(n1128), .A2(n1033), .A3(n1129), .ZN(n1127) );
NOR2_X1 U812 ( .A1(n1115), .A2(n1130), .ZN(G57) );
XOR2_X1 U813 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U814 ( .A(n1133), .B(n1134), .Z(n1132) );
AND2_X1 U815 ( .A1(G472), .A2(n1119), .ZN(n1134) );
XNOR2_X1 U816 ( .A(G101), .B(n1135), .ZN(n1131) );
NOR2_X1 U817 ( .A1(KEYINPUT7), .A2(n1136), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1115), .A2(n1137), .ZN(G54) );
XOR2_X1 U819 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U821 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U822 ( .A(n1144), .B(n1145), .Z(n1140) );
AND2_X1 U823 ( .A1(G469), .A2(n1119), .ZN(n1145) );
INV_X1 U824 ( .A(n1146), .ZN(n1119) );
NAND2_X1 U825 ( .A1(KEYINPUT27), .A2(n1147), .ZN(n1144) );
XOR2_X1 U826 ( .A(n1148), .B(n1149), .Z(n1138) );
XOR2_X1 U827 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR3_X1 U828 ( .A1(n1152), .A2(KEYINPUT3), .A3(G953), .ZN(n1151) );
INV_X1 U829 ( .A(G227), .ZN(n1152) );
NAND2_X1 U830 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
XOR2_X1 U831 ( .A(G128), .B(n1155), .Z(n1154) );
XNOR2_X1 U832 ( .A(KEYINPUT62), .B(KEYINPUT42), .ZN(n1153) );
XNOR2_X1 U833 ( .A(G134), .B(G140), .ZN(n1148) );
NOR2_X1 U834 ( .A1(n1156), .A2(G952), .ZN(n1115) );
NOR2_X1 U835 ( .A1(n1157), .A2(n1158), .ZN(G51) );
XOR2_X1 U836 ( .A(n1159), .B(n1160), .Z(n1158) );
XNOR2_X1 U837 ( .A(n1161), .B(n1162), .ZN(n1160) );
XOR2_X1 U838 ( .A(n1163), .B(n1164), .Z(n1159) );
NOR2_X1 U839 ( .A1(n1085), .A2(n1146), .ZN(n1164) );
NAND2_X1 U840 ( .A1(G902), .A2(n1165), .ZN(n1146) );
OR2_X1 U841 ( .A1(n1027), .A2(n1026), .ZN(n1165) );
NAND4_X1 U842 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1026) );
AND4_X1 U843 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1021), .ZN(n1169) );
NAND3_X1 U844 ( .A1(n1032), .A2(n1033), .A3(n1128), .ZN(n1021) );
NOR2_X1 U845 ( .A1(n1173), .A2(n1174), .ZN(n1168) );
NOR3_X1 U846 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
XOR2_X1 U847 ( .A(KEYINPUT9), .B(n1051), .Z(n1175) );
NOR3_X1 U848 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1173) );
XOR2_X1 U849 ( .A(KEYINPUT56), .B(n1062), .Z(n1180) );
XOR2_X1 U850 ( .A(KEYINPUT15), .B(n1063), .Z(n1179) );
NAND3_X1 U851 ( .A1(n1033), .A2(n1181), .A3(n1129), .ZN(n1178) );
NAND4_X1 U852 ( .A1(n1182), .A2(n1051), .A3(n1183), .A4(n1184), .ZN(n1167) );
OR2_X1 U853 ( .A1(n1185), .A2(n1128), .ZN(n1184) );
NAND2_X1 U854 ( .A1(n1186), .A2(n1185), .ZN(n1183) );
INV_X1 U855 ( .A(KEYINPUT37), .ZN(n1185) );
NAND3_X1 U856 ( .A1(n1181), .A2(n1187), .A3(n1062), .ZN(n1186) );
NAND2_X1 U857 ( .A1(n1188), .A2(n1063), .ZN(n1166) );
NAND4_X1 U858 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1027) );
NOR4_X1 U859 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
INV_X1 U860 ( .A(n1197), .ZN(n1196) );
NOR3_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1191) );
NOR4_X1 U862 ( .A1(n1201), .A2(n1202), .A3(n1053), .A4(n1203), .ZN(n1200) );
NAND3_X1 U863 ( .A1(n1204), .A2(n1187), .A3(n1129), .ZN(n1202) );
INV_X1 U864 ( .A(KEYINPUT50), .ZN(n1201) );
NOR2_X1 U865 ( .A1(KEYINPUT50), .A2(n1205), .ZN(n1199) );
XNOR2_X1 U866 ( .A(n1206), .B(n1207), .ZN(n1163) );
NOR2_X1 U867 ( .A1(KEYINPUT10), .A2(n1208), .ZN(n1207) );
NOR2_X1 U868 ( .A1(G952), .A2(n1209), .ZN(n1157) );
XOR2_X1 U869 ( .A(n1156), .B(KEYINPUT8), .Z(n1209) );
XOR2_X1 U870 ( .A(n1058), .B(KEYINPUT57), .Z(n1156) );
XOR2_X1 U871 ( .A(G146), .B(n1198), .Z(G48) );
AND2_X1 U872 ( .A1(n1129), .A2(n1210), .ZN(n1198) );
XNOR2_X1 U873 ( .A(G143), .B(n1189), .ZN(G45) );
NAND4_X1 U874 ( .A1(n1211), .A2(n1071), .A3(n1212), .A4(n1213), .ZN(n1189) );
NOR2_X1 U875 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
XNOR2_X1 U876 ( .A(G140), .B(n1190), .ZN(G42) );
NAND3_X1 U877 ( .A1(n1129), .A2(n1216), .A3(n1182), .ZN(n1190) );
XOR2_X1 U878 ( .A(G137), .B(n1193), .Z(G39) );
AND3_X1 U879 ( .A1(n1216), .A2(n1217), .A3(n1051), .ZN(n1193) );
NAND2_X1 U880 ( .A1(n1218), .A2(n1219), .ZN(G36) );
NAND2_X1 U881 ( .A1(G134), .A2(n1197), .ZN(n1219) );
XOR2_X1 U882 ( .A(n1220), .B(KEYINPUT19), .Z(n1218) );
OR2_X1 U883 ( .A1(n1197), .A2(G134), .ZN(n1220) );
NAND3_X1 U884 ( .A1(n1216), .A2(n1032), .A3(n1071), .ZN(n1197) );
NAND3_X1 U885 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(G33) );
NAND2_X1 U886 ( .A1(n1195), .A2(n1224), .ZN(n1223) );
NAND2_X1 U887 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
INV_X1 U888 ( .A(KEYINPUT30), .ZN(n1226) );
NAND2_X1 U889 ( .A1(n1227), .A2(G131), .ZN(n1225) );
XNOR2_X1 U890 ( .A(KEYINPUT2), .B(n1195), .ZN(n1227) );
NAND2_X1 U891 ( .A1(KEYINPUT30), .A2(n1228), .ZN(n1221) );
NAND2_X1 U892 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
OR3_X1 U893 ( .A1(n1224), .A2(n1195), .A3(KEYINPUT2), .ZN(n1230) );
NAND2_X1 U894 ( .A1(KEYINPUT2), .A2(n1195), .ZN(n1229) );
AND3_X1 U895 ( .A1(n1129), .A2(n1216), .A3(n1071), .ZN(n1195) );
AND4_X1 U896 ( .A1(n1062), .A2(n1038), .A3(n1204), .A4(n1046), .ZN(n1216) );
XNOR2_X1 U897 ( .A(n1194), .B(n1231), .ZN(G30) );
NAND2_X1 U898 ( .A1(KEYINPUT34), .A2(G128), .ZN(n1231) );
AND2_X1 U899 ( .A1(n1210), .A2(n1032), .ZN(n1194) );
AND3_X1 U900 ( .A1(n1217), .A2(n1062), .A3(n1213), .ZN(n1210) );
INV_X1 U901 ( .A(n1215), .ZN(n1062) );
XNOR2_X1 U902 ( .A(G101), .B(n1172), .ZN(G3) );
NAND3_X1 U903 ( .A1(n1051), .A2(n1128), .A3(n1071), .ZN(n1172) );
XOR2_X1 U904 ( .A(n1205), .B(n1232), .Z(G27) );
XOR2_X1 U905 ( .A(n1208), .B(KEYINPUT45), .Z(n1232) );
NAND4_X1 U906 ( .A1(n1050), .A2(n1182), .A3(n1129), .A4(n1213), .ZN(n1205) );
AND2_X1 U907 ( .A1(n1063), .A2(n1204), .ZN(n1213) );
NAND2_X1 U908 ( .A1(n1072), .A2(n1233), .ZN(n1204) );
NAND4_X1 U909 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1235), .ZN(n1233) );
INV_X1 U910 ( .A(G900), .ZN(n1235) );
XOR2_X1 U911 ( .A(n1236), .B(n1237), .Z(G24) );
NOR2_X1 U912 ( .A1(G122), .A2(KEYINPUT6), .ZN(n1237) );
NAND2_X1 U913 ( .A1(n1063), .A2(n1238), .ZN(n1236) );
XOR2_X1 U914 ( .A(KEYINPUT46), .B(n1188), .Z(n1238) );
AND3_X1 U915 ( .A1(n1211), .A2(n1050), .A3(n1239), .ZN(n1188) );
NOR3_X1 U916 ( .A1(n1080), .A2(n1240), .A3(n1214), .ZN(n1239) );
INV_X1 U917 ( .A(n1033), .ZN(n1080) );
NOR2_X1 U918 ( .A1(n1241), .A2(n1242), .ZN(n1033) );
XNOR2_X1 U919 ( .A(G119), .B(n1243), .ZN(G21) );
NAND3_X1 U920 ( .A1(n1051), .A2(n1217), .A3(n1244), .ZN(n1243) );
INV_X1 U921 ( .A(n1176), .ZN(n1217) );
NAND2_X1 U922 ( .A1(n1242), .A2(n1241), .ZN(n1176) );
INV_X1 U923 ( .A(n1245), .ZN(n1242) );
XNOR2_X1 U924 ( .A(G116), .B(n1171), .ZN(G18) );
NAND3_X1 U925 ( .A1(n1071), .A2(n1032), .A3(n1244), .ZN(n1171) );
NOR2_X1 U926 ( .A1(n1211), .A2(n1214), .ZN(n1032) );
XNOR2_X1 U927 ( .A(G113), .B(n1170), .ZN(G15) );
NAND3_X1 U928 ( .A1(n1071), .A2(n1129), .A3(n1244), .ZN(n1170) );
INV_X1 U929 ( .A(n1177), .ZN(n1244) );
NAND3_X1 U930 ( .A1(n1063), .A2(n1181), .A3(n1050), .ZN(n1177) );
INV_X1 U931 ( .A(n1203), .ZN(n1050) );
NAND2_X1 U932 ( .A1(n1246), .A2(n1048), .ZN(n1203) );
INV_X1 U933 ( .A(n1069), .ZN(n1129) );
NAND2_X1 U934 ( .A1(n1211), .A2(n1214), .ZN(n1069) );
NOR2_X1 U935 ( .A1(n1241), .A2(n1245), .ZN(n1071) );
XOR2_X1 U936 ( .A(n1147), .B(n1247), .Z(G12) );
NAND3_X1 U937 ( .A1(n1051), .A2(n1128), .A3(n1182), .ZN(n1247) );
INV_X1 U938 ( .A(n1053), .ZN(n1182) );
NAND2_X1 U939 ( .A1(n1245), .A2(n1241), .ZN(n1053) );
NAND3_X1 U940 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1241) );
OR2_X1 U941 ( .A1(n1251), .A2(n1118), .ZN(n1250) );
NAND3_X1 U942 ( .A1(n1118), .A2(n1251), .A3(n1252), .ZN(n1249) );
NAND2_X1 U943 ( .A1(G217), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U944 ( .A(n1254), .B(n1255), .ZN(n1118) );
XOR2_X1 U945 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U946 ( .A(G110), .B(n1258), .Z(n1257) );
NOR2_X1 U947 ( .A1(KEYINPUT40), .A2(n1259), .ZN(n1258) );
XOR2_X1 U948 ( .A(KEYINPUT32), .B(G146), .Z(n1259) );
XOR2_X1 U949 ( .A(G137), .B(G125), .Z(n1256) );
XOR2_X1 U950 ( .A(n1260), .B(n1261), .Z(n1254) );
XNOR2_X1 U951 ( .A(n1262), .B(n1263), .ZN(n1261) );
NOR2_X1 U952 ( .A1(KEYINPUT23), .A2(n1264), .ZN(n1263) );
XOR2_X1 U953 ( .A(G128), .B(G119), .Z(n1264) );
NAND2_X1 U954 ( .A1(KEYINPUT5), .A2(G140), .ZN(n1262) );
NAND2_X1 U955 ( .A1(n1265), .A2(G221), .ZN(n1260) );
NAND2_X1 U956 ( .A1(G217), .A2(G902), .ZN(n1248) );
XOR2_X1 U957 ( .A(n1266), .B(G472), .Z(n1245) );
NAND2_X1 U958 ( .A1(n1267), .A2(n1252), .ZN(n1266) );
XOR2_X1 U959 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U960 ( .A(n1133), .B(n1136), .Z(n1269) );
XNOR2_X1 U961 ( .A(n1270), .B(n1271), .ZN(n1136) );
XOR2_X1 U962 ( .A(n1272), .B(n1273), .Z(n1133) );
AND2_X1 U963 ( .A1(G210), .A2(n1274), .ZN(n1273) );
XOR2_X1 U964 ( .A(n1275), .B(n1276), .Z(n1268) );
XOR2_X1 U965 ( .A(KEYINPUT22), .B(KEYINPUT1), .Z(n1276) );
NAND2_X1 U966 ( .A1(n1277), .A2(KEYINPUT13), .ZN(n1275) );
XNOR2_X1 U967 ( .A(G101), .B(KEYINPUT24), .ZN(n1277) );
NOR3_X1 U968 ( .A1(n1187), .A2(n1240), .A3(n1215), .ZN(n1128) );
NAND2_X1 U969 ( .A1(n1047), .A2(n1048), .ZN(n1215) );
NAND2_X1 U970 ( .A1(G221), .A2(n1278), .ZN(n1048) );
NAND2_X1 U971 ( .A1(G234), .A2(n1252), .ZN(n1278) );
INV_X1 U972 ( .A(n1246), .ZN(n1047) );
XNOR2_X1 U973 ( .A(G469), .B(n1279), .ZN(n1246) );
NOR2_X1 U974 ( .A1(KEYINPUT29), .A2(n1083), .ZN(n1279) );
NAND2_X1 U975 ( .A1(n1280), .A2(n1252), .ZN(n1083) );
XOR2_X1 U976 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U977 ( .A(G110), .B(n1283), .Z(n1282) );
XOR2_X1 U978 ( .A(KEYINPUT33), .B(G227), .Z(n1283) );
XOR2_X1 U979 ( .A(n1284), .B(n1100), .Z(n1281) );
XOR2_X1 U980 ( .A(n1155), .B(n1270), .Z(n1100) );
XOR2_X1 U981 ( .A(n1143), .B(n1285), .Z(n1270) );
XOR2_X1 U982 ( .A(n1286), .B(n1224), .Z(n1143) );
INV_X1 U983 ( .A(G131), .ZN(n1224) );
INV_X1 U984 ( .A(G137), .ZN(n1286) );
XOR2_X1 U985 ( .A(n1142), .B(n1287), .Z(n1284) );
NOR2_X1 U986 ( .A1(G140), .A2(KEYINPUT20), .ZN(n1287) );
XOR2_X1 U987 ( .A(n1288), .B(KEYINPUT61), .Z(n1142) );
INV_X1 U988 ( .A(n1181), .ZN(n1240) );
NAND2_X1 U989 ( .A1(n1072), .A2(n1289), .ZN(n1181) );
NAND4_X1 U990 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1107), .ZN(n1289) );
INV_X1 U991 ( .A(G898), .ZN(n1107) );
NAND3_X1 U992 ( .A1(n1234), .A2(n1058), .A3(G952), .ZN(n1072) );
NAND2_X1 U993 ( .A1(G237), .A2(G234), .ZN(n1234) );
INV_X1 U994 ( .A(n1063), .ZN(n1187) );
NOR2_X1 U995 ( .A1(n1038), .A2(n1041), .ZN(n1063) );
INV_X1 U996 ( .A(n1046), .ZN(n1041) );
NAND2_X1 U997 ( .A1(G214), .A2(n1290), .ZN(n1046) );
XOR2_X1 U998 ( .A(n1291), .B(n1085), .Z(n1038) );
NAND2_X1 U999 ( .A1(G210), .A2(n1290), .ZN(n1085) );
NAND2_X1 U1000 ( .A1(n1292), .A2(n1252), .ZN(n1290) );
INV_X1 U1001 ( .A(G237), .ZN(n1292) );
XOR2_X1 U1002 ( .A(n1087), .B(KEYINPUT59), .Z(n1291) );
NAND2_X1 U1003 ( .A1(n1293), .A2(n1252), .ZN(n1087) );
XOR2_X1 U1004 ( .A(n1161), .B(n1294), .Z(n1293) );
NOR2_X1 U1005 ( .A1(KEYINPUT25), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1006 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U1007 ( .A(n1298), .B(n1299), .ZN(n1297) );
NAND2_X1 U1008 ( .A1(KEYINPUT18), .A2(n1162), .ZN(n1299) );
XNOR2_X1 U1009 ( .A(G128), .B(n1271), .ZN(n1162) );
NOR2_X1 U1010 ( .A1(KEYINPUT63), .A2(n1300), .ZN(n1271) );
XNOR2_X1 U1011 ( .A(n1155), .B(KEYINPUT39), .ZN(n1300) );
XOR2_X1 U1012 ( .A(G143), .B(G146), .Z(n1155) );
NAND2_X1 U1013 ( .A1(KEYINPUT55), .A2(n1206), .ZN(n1298) );
AND2_X1 U1014 ( .A1(G224), .A2(n1058), .ZN(n1206) );
INV_X1 U1015 ( .A(G953), .ZN(n1058) );
XOR2_X1 U1016 ( .A(n1208), .B(KEYINPUT47), .Z(n1296) );
INV_X1 U1017 ( .A(G125), .ZN(n1208) );
XNOR2_X1 U1018 ( .A(n1114), .B(n1112), .ZN(n1161) );
AND2_X1 U1019 ( .A1(n1301), .A2(n1302), .ZN(n1112) );
NAND2_X1 U1020 ( .A1(G122), .A2(n1147), .ZN(n1302) );
XOR2_X1 U1021 ( .A(n1303), .B(KEYINPUT16), .Z(n1301) );
NAND2_X1 U1022 ( .A1(G110), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U1023 ( .A(n1305), .B(n1306), .ZN(n1114) );
INV_X1 U1024 ( .A(n1288), .ZN(n1306) );
XNOR2_X1 U1025 ( .A(G101), .B(n1307), .ZN(n1288) );
XOR2_X1 U1026 ( .A(G107), .B(G104), .Z(n1307) );
XOR2_X1 U1027 ( .A(n1272), .B(KEYINPUT38), .Z(n1305) );
XNOR2_X1 U1028 ( .A(G113), .B(n1308), .ZN(n1272) );
XOR2_X1 U1029 ( .A(G119), .B(G116), .Z(n1308) );
NOR2_X1 U1030 ( .A1(n1081), .A2(n1211), .ZN(n1051) );
XOR2_X1 U1031 ( .A(n1074), .B(KEYINPUT49), .Z(n1211) );
XOR2_X1 U1032 ( .A(n1309), .B(G475), .Z(n1074) );
NAND2_X1 U1033 ( .A1(n1125), .A2(n1252), .ZN(n1309) );
XOR2_X1 U1034 ( .A(n1310), .B(n1311), .Z(n1125) );
XOR2_X1 U1035 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1036 ( .A(n1126), .B(n1314), .Z(n1313) );
NOR2_X1 U1037 ( .A1(G143), .A2(KEYINPUT0), .ZN(n1314) );
INV_X1 U1038 ( .A(G104), .ZN(n1126) );
XOR2_X1 U1039 ( .A(G113), .B(n1304), .Z(n1312) );
XOR2_X1 U1040 ( .A(n1315), .B(n1316), .Z(n1310) );
XNOR2_X1 U1041 ( .A(n1317), .B(n1318), .ZN(n1316) );
NOR2_X1 U1042 ( .A1(G131), .A2(KEYINPUT35), .ZN(n1318) );
NAND2_X1 U1043 ( .A1(KEYINPUT60), .A2(n1319), .ZN(n1317) );
INV_X1 U1044 ( .A(G146), .ZN(n1319) );
XOR2_X1 U1045 ( .A(n1320), .B(n1099), .Z(n1315) );
XOR2_X1 U1046 ( .A(G125), .B(G140), .Z(n1099) );
NAND2_X1 U1047 ( .A1(n1274), .A2(G214), .ZN(n1320) );
NOR2_X1 U1048 ( .A1(G953), .A2(G237), .ZN(n1274) );
INV_X1 U1049 ( .A(n1214), .ZN(n1081) );
XOR2_X1 U1050 ( .A(n1321), .B(G478), .Z(n1214) );
NAND2_X1 U1051 ( .A1(n1121), .A2(n1252), .ZN(n1321) );
INV_X1 U1052 ( .A(G902), .ZN(n1252) );
XNOR2_X1 U1053 ( .A(n1322), .B(n1323), .ZN(n1121) );
XOR2_X1 U1054 ( .A(n1324), .B(n1325), .Z(n1323) );
XNOR2_X1 U1055 ( .A(G107), .B(G116), .ZN(n1325) );
NAND2_X1 U1056 ( .A1(n1326), .A2(KEYINPUT52), .ZN(n1324) );
XNOR2_X1 U1057 ( .A(G143), .B(n1285), .ZN(n1326) );
XOR2_X1 U1058 ( .A(G128), .B(G134), .Z(n1285) );
XNOR2_X1 U1059 ( .A(n1327), .B(n1328), .ZN(n1322) );
NAND2_X1 U1060 ( .A1(KEYINPUT4), .A2(n1304), .ZN(n1328) );
INV_X1 U1061 ( .A(G122), .ZN(n1304) );
NAND3_X1 U1062 ( .A1(G217), .A2(n1265), .A3(KEYINPUT26), .ZN(n1327) );
NOR2_X1 U1063 ( .A1(n1253), .A2(G953), .ZN(n1265) );
INV_X1 U1064 ( .A(G234), .ZN(n1253) );
INV_X1 U1065 ( .A(G110), .ZN(n1147) );
endmodule


