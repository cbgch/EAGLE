//Key = 0111000010111000000111010001001110100111101110110001100110111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301;

XOR2_X1 U719 ( .A(n996), .B(n997), .Z(G9) );
XNOR2_X1 U720 ( .A(KEYINPUT56), .B(n998), .ZN(n997) );
NOR2_X1 U721 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U722 ( .A1(n1001), .A2(n1002), .A3(G953), .A4(n1003), .ZN(n1000) );
NOR3_X1 U723 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1002) );
NOR4_X1 U724 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1005) );
NAND3_X1 U725 ( .A1(G952), .A2(n1011), .A3(n1012), .ZN(n1001) );
NAND2_X1 U726 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NAND2_X1 U727 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND3_X1 U728 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NAND2_X1 U729 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NAND2_X1 U730 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U731 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U732 ( .A1(n1026), .A2(n1004), .ZN(n1025) );
INV_X1 U733 ( .A(KEYINPUT13), .ZN(n1004) );
INV_X1 U734 ( .A(n1027), .ZN(n1024) );
NAND2_X1 U735 ( .A1(n1028), .A2(n1029), .ZN(n1020) );
NAND2_X1 U736 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U737 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
INV_X1 U738 ( .A(n1034), .ZN(n1030) );
NAND3_X1 U739 ( .A1(n1035), .A2(n1036), .A3(n1028), .ZN(n1015) );
NAND2_X1 U740 ( .A1(n1037), .A2(n1007), .ZN(n1036) );
NAND4_X1 U741 ( .A1(n1038), .A2(n1017), .A3(n1039), .A4(n1040), .ZN(n1037) );
INV_X1 U742 ( .A(KEYINPUT51), .ZN(n1040) );
NAND4_X1 U743 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1022), .ZN(n1035) );
NAND2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
XNOR2_X1 U745 ( .A(n1017), .B(KEYINPUT19), .ZN(n1044) );
NAND4_X1 U746 ( .A1(KEYINPUT51), .A2(n1038), .A3(n1039), .A4(n1017), .ZN(n1042) );
NAND2_X1 U747 ( .A1(n1019), .A2(n1046), .ZN(n1041) );
NAND2_X1 U748 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U749 ( .A1(G214), .A2(n1049), .A3(n1050), .ZN(n1048) );
INV_X1 U750 ( .A(n1010), .ZN(n1013) );
NOR3_X1 U751 ( .A1(n1051), .A2(G953), .A3(n1003), .ZN(n999) );
AND4_X1 U752 ( .A1(n1032), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1003) );
NOR4_X1 U753 ( .A1(n1055), .A2(n1056), .A3(n1006), .A4(n1057), .ZN(n1054) );
XOR2_X1 U754 ( .A(n1058), .B(n1059), .Z(n1057) );
NAND2_X1 U755 ( .A1(KEYINPUT47), .A2(n1060), .ZN(n1059) );
AND2_X1 U756 ( .A1(n1008), .A2(KEYINPUT11), .ZN(n1056) );
NOR2_X1 U757 ( .A1(KEYINPUT11), .A2(n1045), .ZN(n1055) );
XNOR2_X1 U758 ( .A(KEYINPUT38), .B(n1061), .ZN(n1052) );
XOR2_X1 U759 ( .A(KEYINPUT14), .B(G952), .Z(n1051) );
XOR2_X1 U760 ( .A(n1062), .B(n1063), .Z(G72) );
NOR2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND2_X1 U762 ( .A1(G227), .A2(G900), .ZN(n1064) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U766 ( .A(KEYINPUT43), .B(n1072), .Z(n1066) );
NOR4_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
XOR2_X1 U768 ( .A(KEYINPUT25), .B(n1068), .Z(n1076) );
AND2_X1 U769 ( .A1(n1077), .A2(n1065), .ZN(n1068) );
NAND2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
INV_X1 U771 ( .A(n1071), .ZN(n1075) );
NAND3_X1 U772 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1071) );
INV_X1 U773 ( .A(n1070), .ZN(n1074) );
NAND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1070) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1084) );
NAND2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
XNOR2_X1 U777 ( .A(KEYINPUT60), .B(n1087), .ZN(n1080) );
NAND2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U779 ( .A(KEYINPUT53), .B(n1085), .ZN(n1089) );
INV_X1 U780 ( .A(n1086), .ZN(n1088) );
XOR2_X1 U781 ( .A(G131), .B(n1090), .Z(n1086) );
XNOR2_X1 U782 ( .A(n1091), .B(G134), .ZN(n1090) );
XOR2_X1 U783 ( .A(n1092), .B(n1093), .Z(G69) );
XOR2_X1 U784 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U785 ( .A1(n1096), .A2(G953), .ZN(n1095) );
NOR2_X1 U786 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
XNOR2_X1 U787 ( .A(n1099), .B(KEYINPUT40), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1100), .A2(n1065), .ZN(n1092) );
AND2_X1 U789 ( .A1(G224), .A2(G898), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(G66) );
XOR2_X1 U791 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U792 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
INV_X1 U793 ( .A(n1107), .ZN(n1106) );
NOR2_X1 U794 ( .A1(n1101), .A2(n1108), .ZN(G63) );
XOR2_X1 U795 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U796 ( .A1(KEYINPUT17), .A2(n1111), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1107), .A2(G478), .ZN(n1109) );
NOR2_X1 U798 ( .A1(n1101), .A2(n1112), .ZN(G60) );
XOR2_X1 U799 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND3_X1 U800 ( .A1(n1107), .A2(G475), .A3(KEYINPUT27), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(G6) );
NAND2_X1 U802 ( .A1(KEYINPUT59), .A2(G104), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
XOR2_X1 U804 ( .A(n1119), .B(KEYINPUT31), .Z(n1117) );
NOR2_X1 U805 ( .A1(n1101), .A2(n1120), .ZN(G57) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U807 ( .A(n1123), .B(n1124), .Z(n1122) );
AND2_X1 U808 ( .A1(G472), .A2(n1107), .ZN(n1123) );
XOR2_X1 U809 ( .A(KEYINPUT54), .B(n1125), .Z(n1121) );
NOR2_X1 U810 ( .A1(KEYINPUT9), .A2(n1126), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1101), .A2(n1127), .ZN(G54) );
XOR2_X1 U812 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U813 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U814 ( .A(n1132), .B(n1133), .ZN(n1131) );
AND2_X1 U815 ( .A1(G469), .A2(n1107), .ZN(n1132) );
XOR2_X1 U816 ( .A(n1134), .B(n1135), .Z(n1128) );
XNOR2_X1 U817 ( .A(KEYINPUT20), .B(n1136), .ZN(n1134) );
NOR2_X1 U818 ( .A1(KEYINPUT24), .A2(n1137), .ZN(n1136) );
XOR2_X1 U819 ( .A(KEYINPUT10), .B(n1138), .Z(n1137) );
NOR2_X1 U820 ( .A1(n1101), .A2(n1139), .ZN(G51) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U822 ( .A(n1142), .B(n1143), .ZN(n1141) );
XOR2_X1 U823 ( .A(n1144), .B(n1145), .Z(n1140) );
NOR2_X1 U824 ( .A1(KEYINPUT6), .A2(n1146), .ZN(n1145) );
NAND4_X1 U825 ( .A1(G210), .A2(n1049), .A3(n1147), .A4(n1148), .ZN(n1144) );
OR2_X1 U826 ( .A1(n1107), .A2(KEYINPUT48), .ZN(n1148) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1012), .ZN(n1107) );
NAND2_X1 U828 ( .A1(KEYINPUT48), .A2(n1150), .ZN(n1147) );
NAND2_X1 U829 ( .A1(n1012), .A2(G902), .ZN(n1150) );
AND3_X1 U830 ( .A1(n1078), .A2(n1151), .A3(n1096), .ZN(n1012) );
AND4_X1 U831 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1096) );
NOR4_X1 U832 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NOR2_X1 U833 ( .A1(n1047), .A2(n1119), .ZN(n1159) );
NAND3_X1 U834 ( .A1(n1160), .A2(n1045), .A3(n1026), .ZN(n1119) );
NOR3_X1 U835 ( .A1(n1161), .A2(n1047), .A3(n1162), .ZN(n1158) );
XNOR2_X1 U836 ( .A(KEYINPUT46), .B(n1008), .ZN(n1161) );
INV_X1 U837 ( .A(n1163), .ZN(n1156) );
AND2_X1 U838 ( .A1(n1164), .A2(n996), .ZN(n1154) );
NAND3_X1 U839 ( .A1(n1160), .A2(n1165), .A3(n1027), .ZN(n996) );
XOR2_X1 U840 ( .A(KEYINPUT28), .B(n1079), .Z(n1151) );
AND4_X1 U841 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1079) );
AND4_X1 U842 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1078) );
NAND2_X1 U843 ( .A1(n1174), .A2(n1175), .ZN(n1170) );
XNOR2_X1 U844 ( .A(n1017), .B(KEYINPUT52), .ZN(n1174) );
AND2_X1 U845 ( .A1(n1176), .A2(G953), .ZN(n1101) );
XNOR2_X1 U846 ( .A(G952), .B(KEYINPUT41), .ZN(n1176) );
XNOR2_X1 U847 ( .A(G146), .B(n1171), .ZN(G48) );
NAND3_X1 U848 ( .A1(n1026), .A2(n1118), .A3(n1177), .ZN(n1171) );
XNOR2_X1 U849 ( .A(G143), .B(n1172), .ZN(G45) );
NAND4_X1 U850 ( .A1(n1178), .A2(n1034), .A3(n1179), .A4(n1165), .ZN(n1172) );
AND2_X1 U851 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XNOR2_X1 U852 ( .A(G140), .B(n1173), .ZN(G42) );
NAND2_X1 U853 ( .A1(n1182), .A2(n1183), .ZN(n1173) );
XNOR2_X1 U854 ( .A(G137), .B(n1184), .ZN(G39) );
NAND2_X1 U855 ( .A1(n1175), .A2(n1017), .ZN(n1184) );
AND2_X1 U856 ( .A1(n1177), .A2(n1028), .ZN(n1175) );
XNOR2_X1 U857 ( .A(G134), .B(n1166), .ZN(G36) );
NAND3_X1 U858 ( .A1(n1034), .A2(n1027), .A3(n1183), .ZN(n1166) );
XNOR2_X1 U859 ( .A(G131), .B(n1167), .ZN(G33) );
NAND3_X1 U860 ( .A1(n1034), .A2(n1026), .A3(n1183), .ZN(n1167) );
AND3_X1 U861 ( .A1(n1045), .A2(n1180), .A3(n1017), .ZN(n1183) );
INV_X1 U862 ( .A(n1006), .ZN(n1017) );
NAND2_X1 U863 ( .A1(n1050), .A2(n1185), .ZN(n1006) );
NAND2_X1 U864 ( .A1(G214), .A2(n1049), .ZN(n1185) );
XNOR2_X1 U865 ( .A(G128), .B(n1168), .ZN(G30) );
NAND3_X1 U866 ( .A1(n1027), .A2(n1118), .A3(n1177), .ZN(n1168) );
AND4_X1 U867 ( .A1(n1045), .A2(n1033), .A3(n1186), .A4(n1180), .ZN(n1177) );
XNOR2_X1 U868 ( .A(G101), .B(n1164), .ZN(G3) );
NAND4_X1 U869 ( .A1(n1028), .A2(n1034), .A3(n1165), .A4(n1187), .ZN(n1164) );
XOR2_X1 U870 ( .A(n1169), .B(n1188), .Z(G27) );
NAND2_X1 U871 ( .A1(KEYINPUT44), .A2(G125), .ZN(n1188) );
NAND4_X1 U872 ( .A1(n1182), .A2(n1019), .A3(n1118), .A4(n1180), .ZN(n1169) );
NAND2_X1 U873 ( .A1(n1010), .A2(n1189), .ZN(n1180) );
NAND3_X1 U874 ( .A1(G902), .A2(n1190), .A3(n1073), .ZN(n1189) );
NOR2_X1 U875 ( .A1(n1065), .A2(G900), .ZN(n1073) );
NOR3_X1 U876 ( .A1(n1186), .A2(n1061), .A3(n1009), .ZN(n1182) );
INV_X1 U877 ( .A(n1026), .ZN(n1009) );
XOR2_X1 U878 ( .A(G122), .B(n1157), .Z(G24) );
AND4_X1 U879 ( .A1(n1178), .A2(n1019), .A3(n1191), .A4(n1160), .ZN(n1157) );
NOR2_X1 U880 ( .A1(n1007), .A2(n1192), .ZN(n1160) );
INV_X1 U881 ( .A(n1022), .ZN(n1007) );
NOR2_X1 U882 ( .A1(n1186), .A2(n1033), .ZN(n1022) );
NOR2_X1 U883 ( .A1(n1053), .A2(n1047), .ZN(n1191) );
INV_X1 U884 ( .A(n1008), .ZN(n1019) );
XNOR2_X1 U885 ( .A(G119), .B(n1152), .ZN(G21) );
NAND4_X1 U886 ( .A1(n1028), .A2(n1193), .A3(n1033), .A4(n1186), .ZN(n1152) );
XOR2_X1 U887 ( .A(G116), .B(n1194), .Z(G18) );
NOR3_X1 U888 ( .A1(n1162), .A2(n1195), .A3(n1008), .ZN(n1194) );
XNOR2_X1 U889 ( .A(n1118), .B(KEYINPUT15), .ZN(n1195) );
NAND3_X1 U890 ( .A1(n1027), .A2(n1187), .A3(n1034), .ZN(n1162) );
NOR2_X1 U891 ( .A1(n1053), .A2(n1178), .ZN(n1027) );
INV_X1 U892 ( .A(n1181), .ZN(n1053) );
XNOR2_X1 U893 ( .A(G113), .B(n1153), .ZN(G15) );
NAND3_X1 U894 ( .A1(n1026), .A2(n1193), .A3(n1034), .ZN(n1153) );
NOR2_X1 U895 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
INV_X1 U896 ( .A(n1186), .ZN(n1032) );
NOR3_X1 U897 ( .A1(n1047), .A2(n1192), .A3(n1008), .ZN(n1193) );
NAND2_X1 U898 ( .A1(n1039), .A2(n1196), .ZN(n1008) );
INV_X1 U899 ( .A(n1118), .ZN(n1047) );
NOR2_X1 U900 ( .A1(n1197), .A2(n1181), .ZN(n1026) );
NAND2_X1 U901 ( .A1(n1198), .A2(n1199), .ZN(G12) );
OR2_X1 U902 ( .A1(n1163), .A2(G110), .ZN(n1199) );
XOR2_X1 U903 ( .A(n1200), .B(KEYINPUT22), .Z(n1198) );
NAND2_X1 U904 ( .A1(G110), .A2(n1163), .ZN(n1200) );
NAND3_X1 U905 ( .A1(n1028), .A2(n1165), .A3(n1201), .ZN(n1163) );
NOR3_X1 U906 ( .A1(n1186), .A2(n1192), .A3(n1061), .ZN(n1201) );
INV_X1 U907 ( .A(n1033), .ZN(n1061) );
XOR2_X1 U908 ( .A(n1202), .B(n1105), .Z(n1033) );
NAND2_X1 U909 ( .A1(G217), .A2(n1203), .ZN(n1105) );
OR2_X1 U910 ( .A1(n1104), .A2(G902), .ZN(n1202) );
XNOR2_X1 U911 ( .A(n1204), .B(n1205), .ZN(n1104) );
XOR2_X1 U912 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U913 ( .A(G119), .B(G128), .ZN(n1207) );
NAND2_X1 U914 ( .A1(KEYINPUT8), .A2(n1208), .ZN(n1206) );
XNOR2_X1 U915 ( .A(G137), .B(n1209), .ZN(n1208) );
NAND2_X1 U916 ( .A1(G221), .A2(n1210), .ZN(n1209) );
XOR2_X1 U917 ( .A(n1211), .B(n1212), .Z(n1204) );
NOR2_X1 U918 ( .A1(G110), .A2(KEYINPUT49), .ZN(n1212) );
NAND2_X1 U919 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
NAND2_X1 U920 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U921 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XNOR2_X1 U922 ( .A(KEYINPUT3), .B(n1219), .ZN(n1217) );
INV_X1 U923 ( .A(n1220), .ZN(n1215) );
NAND2_X1 U924 ( .A1(n1221), .A2(n1220), .ZN(n1213) );
NAND2_X1 U925 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
OR2_X1 U926 ( .A1(n1219), .A2(KEYINPUT3), .ZN(n1223) );
NAND2_X1 U927 ( .A1(KEYINPUT3), .A2(n1082), .ZN(n1222) );
INV_X1 U928 ( .A(n1187), .ZN(n1192) );
NAND2_X1 U929 ( .A1(n1010), .A2(n1224), .ZN(n1187) );
NAND3_X1 U930 ( .A1(G902), .A2(n1190), .A3(n1099), .ZN(n1224) );
NOR2_X1 U931 ( .A1(n1065), .A2(G898), .ZN(n1099) );
NAND3_X1 U932 ( .A1(n1190), .A2(n1065), .A3(G952), .ZN(n1010) );
NAND2_X1 U933 ( .A1(G237), .A2(G234), .ZN(n1190) );
XNOR2_X1 U934 ( .A(n1225), .B(G472), .ZN(n1186) );
NAND2_X1 U935 ( .A1(n1226), .A2(n1149), .ZN(n1225) );
XNOR2_X1 U936 ( .A(n1143), .B(n1124), .ZN(n1226) );
XNOR2_X1 U937 ( .A(n1227), .B(n1228), .ZN(n1124) );
XNOR2_X1 U938 ( .A(n1229), .B(n1230), .ZN(n1228) );
XNOR2_X1 U939 ( .A(n1231), .B(n1232), .ZN(n1230) );
NOR2_X1 U940 ( .A1(G113), .A2(KEYINPUT57), .ZN(n1232) );
XOR2_X1 U941 ( .A(n1233), .B(n1234), .Z(n1227) );
XNOR2_X1 U942 ( .A(n1235), .B(G101), .ZN(n1234) );
NAND2_X1 U943 ( .A1(G210), .A2(n1236), .ZN(n1233) );
AND2_X1 U944 ( .A1(n1045), .A2(n1118), .ZN(n1165) );
NOR2_X1 U945 ( .A1(n1050), .A2(n1237), .ZN(n1118) );
AND2_X1 U946 ( .A1(G214), .A2(n1049), .ZN(n1237) );
XOR2_X1 U947 ( .A(n1238), .B(n1239), .Z(n1050) );
AND2_X1 U948 ( .A1(n1049), .A2(G210), .ZN(n1239) );
NAND2_X1 U949 ( .A1(n1240), .A2(n1241), .ZN(n1049) );
INV_X1 U950 ( .A(G237), .ZN(n1241) );
NAND2_X1 U951 ( .A1(n1242), .A2(n1149), .ZN(n1238) );
XNOR2_X1 U952 ( .A(n1142), .B(n1243), .ZN(n1242) );
NOR2_X1 U953 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U954 ( .A(KEYINPUT50), .B(n1246), .Z(n1245) );
NOR2_X1 U955 ( .A1(n1146), .A2(n1126), .ZN(n1246) );
NOR2_X1 U956 ( .A1(G125), .A2(n1143), .ZN(n1244) );
INV_X1 U957 ( .A(n1126), .ZN(n1143) );
XNOR2_X1 U958 ( .A(n1247), .B(n1248), .ZN(n1126) );
XOR2_X1 U959 ( .A(n1249), .B(G143), .Z(n1247) );
NAND2_X1 U960 ( .A1(KEYINPUT42), .A2(n1220), .ZN(n1249) );
XNOR2_X1 U961 ( .A(n1250), .B(n1098), .ZN(n1142) );
XNOR2_X1 U962 ( .A(n1251), .B(n1252), .ZN(n1098) );
XOR2_X1 U963 ( .A(n1133), .B(n1253), .Z(n1252) );
XNOR2_X1 U964 ( .A(n1254), .B(n1255), .ZN(n1253) );
NOR2_X1 U965 ( .A1(KEYINPUT5), .A2(n1231), .ZN(n1255) );
XOR2_X1 U966 ( .A(n1256), .B(n1257), .Z(n1251) );
XNOR2_X1 U967 ( .A(KEYINPUT1), .B(n1235), .ZN(n1257) );
INV_X1 U968 ( .A(G119), .ZN(n1235) );
XOR2_X1 U969 ( .A(n1258), .B(G113), .Z(n1256) );
NAND2_X1 U970 ( .A1(KEYINPUT12), .A2(G110), .ZN(n1258) );
NAND2_X1 U971 ( .A1(G224), .A2(n1065), .ZN(n1250) );
NOR2_X1 U972 ( .A1(n1039), .A2(n1038), .ZN(n1045) );
INV_X1 U973 ( .A(n1196), .ZN(n1038) );
NAND2_X1 U974 ( .A1(G221), .A2(n1203), .ZN(n1196) );
NAND2_X1 U975 ( .A1(n1240), .A2(G234), .ZN(n1203) );
XNOR2_X1 U976 ( .A(G902), .B(KEYINPUT4), .ZN(n1240) );
XOR2_X1 U977 ( .A(n1259), .B(G469), .Z(n1039) );
NAND2_X1 U978 ( .A1(n1260), .A2(n1149), .ZN(n1259) );
XOR2_X1 U979 ( .A(n1130), .B(n1261), .Z(n1260) );
XOR2_X1 U980 ( .A(n1262), .B(n1263), .Z(n1261) );
NOR2_X1 U981 ( .A1(KEYINPUT36), .A2(n1133), .ZN(n1263) );
XNOR2_X1 U982 ( .A(G101), .B(n1264), .ZN(n1133) );
XNOR2_X1 U983 ( .A(n998), .B(G104), .ZN(n1264) );
NAND2_X1 U984 ( .A1(KEYINPUT32), .A2(n1265), .ZN(n1262) );
XOR2_X1 U985 ( .A(n1138), .B(n1266), .Z(n1265) );
XNOR2_X1 U986 ( .A(n1267), .B(KEYINPUT7), .ZN(n1266) );
NAND2_X1 U987 ( .A1(KEYINPUT23), .A2(n1135), .ZN(n1267) );
AND2_X1 U988 ( .A1(G227), .A2(n1065), .ZN(n1135) );
XOR2_X1 U989 ( .A(G110), .B(n1268), .Z(n1138) );
XNOR2_X1 U990 ( .A(KEYINPUT63), .B(n1269), .ZN(n1268) );
XOR2_X1 U991 ( .A(n1085), .B(n1229), .Z(n1130) );
AND2_X1 U992 ( .A1(n1270), .A2(n1271), .ZN(n1229) );
NAND2_X1 U993 ( .A1(n1272), .A2(n1091), .ZN(n1271) );
INV_X1 U994 ( .A(G137), .ZN(n1091) );
XOR2_X1 U995 ( .A(KEYINPUT45), .B(n1273), .Z(n1272) );
NAND2_X1 U996 ( .A1(n1274), .A2(G137), .ZN(n1270) );
XOR2_X1 U997 ( .A(KEYINPUT62), .B(n1273), .Z(n1274) );
XNOR2_X1 U998 ( .A(n1275), .B(G134), .ZN(n1273) );
NAND2_X1 U999 ( .A1(KEYINPUT34), .A2(G131), .ZN(n1275) );
XNOR2_X1 U1000 ( .A(n1220), .B(n1276), .ZN(n1085) );
XOR2_X1 U1001 ( .A(n1277), .B(n1248), .Z(n1276) );
XOR2_X1 U1002 ( .A(G128), .B(KEYINPUT55), .Z(n1248) );
NOR2_X1 U1003 ( .A1(G143), .A2(KEYINPUT35), .ZN(n1277) );
NOR2_X1 U1004 ( .A1(n1181), .A2(n1178), .ZN(n1028) );
INV_X1 U1005 ( .A(n1197), .ZN(n1178) );
XOR2_X1 U1006 ( .A(n1058), .B(n1060), .Z(n1197) );
XNOR2_X1 U1007 ( .A(G475), .B(KEYINPUT37), .ZN(n1060) );
NAND2_X1 U1008 ( .A1(n1114), .A2(n1149), .ZN(n1058) );
INV_X1 U1009 ( .A(G902), .ZN(n1149) );
XNOR2_X1 U1010 ( .A(n1278), .B(n1279), .ZN(n1114) );
XNOR2_X1 U1011 ( .A(n1280), .B(n1220), .ZN(n1279) );
XOR2_X1 U1012 ( .A(G146), .B(KEYINPUT30), .Z(n1220) );
NAND2_X1 U1013 ( .A1(KEYINPUT21), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1014 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U1015 ( .A(n1284), .B(n1254), .Z(n1283) );
NOR2_X1 U1016 ( .A1(G113), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U1017 ( .A(KEYINPUT58), .B(KEYINPUT16), .ZN(n1285) );
XOR2_X1 U1018 ( .A(KEYINPUT0), .B(G104), .Z(n1282) );
XNOR2_X1 U1019 ( .A(n1082), .B(n1286), .ZN(n1278) );
NOR2_X1 U1020 ( .A1(KEYINPUT26), .A2(n1287), .ZN(n1286) );
XOR2_X1 U1021 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U1022 ( .A(G131), .B(n1290), .Z(n1289) );
NOR2_X1 U1023 ( .A1(G143), .A2(KEYINPUT29), .ZN(n1290) );
NAND2_X1 U1024 ( .A1(G214), .A2(n1236), .ZN(n1288) );
NOR2_X1 U1025 ( .A1(G953), .A2(G237), .ZN(n1236) );
INV_X1 U1026 ( .A(n1083), .ZN(n1082) );
NAND2_X1 U1027 ( .A1(n1219), .A2(n1218), .ZN(n1083) );
NAND2_X1 U1028 ( .A1(G140), .A2(n1146), .ZN(n1218) );
INV_X1 U1029 ( .A(G125), .ZN(n1146) );
NAND2_X1 U1030 ( .A1(G125), .A2(n1269), .ZN(n1219) );
INV_X1 U1031 ( .A(G140), .ZN(n1269) );
XNOR2_X1 U1032 ( .A(n1291), .B(G478), .ZN(n1181) );
OR2_X1 U1033 ( .A1(n1111), .A2(G902), .ZN(n1291) );
XOR2_X1 U1034 ( .A(n1292), .B(n1293), .Z(n1111) );
XOR2_X1 U1035 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U1036 ( .A(n1296), .B(G128), .Z(n1295) );
NAND2_X1 U1037 ( .A1(G217), .A2(n1210), .ZN(n1296) );
AND2_X1 U1038 ( .A1(G234), .A2(n1065), .ZN(n1210) );
INV_X1 U1039 ( .A(G953), .ZN(n1065) );
XNOR2_X1 U1040 ( .A(G134), .B(G143), .ZN(n1294) );
XOR2_X1 U1041 ( .A(n1297), .B(n1298), .Z(n1292) );
NOR2_X1 U1042 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NOR2_X1 U1043 ( .A1(KEYINPUT2), .A2(n1254), .ZN(n1300) );
AND2_X1 U1044 ( .A1(KEYINPUT39), .A2(n1254), .ZN(n1299) );
XOR2_X1 U1045 ( .A(G122), .B(KEYINPUT18), .Z(n1254) );
XOR2_X1 U1046 ( .A(n1301), .B(n1231), .Z(n1297) );
XOR2_X1 U1047 ( .A(G116), .B(KEYINPUT33), .Z(n1231) );
NAND2_X1 U1048 ( .A1(KEYINPUT61), .A2(n998), .ZN(n1301) );
INV_X1 U1049 ( .A(G107), .ZN(n998) );
endmodule


