//Key = 1110011000111110100100001101100001110000100010000111010001011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360;

XOR2_X1 U740 ( .A(n1033), .B(n1034), .Z(G9) );
NAND2_X1 U741 ( .A1(KEYINPUT12), .A2(G107), .ZN(n1034) );
NOR2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U743 ( .A1(G953), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1036) );
NOR2_X1 U744 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U745 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR3_X1 U746 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NOR2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U748 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U751 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U753 ( .A1(n1059), .A2(n1060), .ZN(n1051) );
NOR2_X1 U754 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U755 ( .A1(n1060), .A2(n1063), .A3(n1054), .ZN(n1047) );
NOR2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR4_X1 U757 ( .A1(n1066), .A2(n1054), .A3(n1060), .A4(n1050), .ZN(n1042) );
NOR2_X1 U758 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U759 ( .A1(n1069), .A2(n1044), .ZN(n1067) );
NOR3_X1 U760 ( .A1(n1037), .A2(G953), .A3(G952), .ZN(n1035) );
AND4_X1 U761 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1037) );
NOR4_X1 U762 ( .A1(n1074), .A2(n1044), .A3(n1075), .A4(n1076), .ZN(n1073) );
XOR2_X1 U763 ( .A(KEYINPUT23), .B(n1058), .Z(n1076) );
XNOR2_X1 U764 ( .A(KEYINPUT47), .B(n1057), .ZN(n1075) );
NOR3_X1 U765 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1072) );
INV_X1 U766 ( .A(n1069), .ZN(n1079) );
NOR2_X1 U767 ( .A1(n1080), .A2(n1081), .ZN(n1077) );
XOR2_X1 U768 ( .A(KEYINPUT2), .B(n1082), .Z(n1081) );
XNOR2_X1 U769 ( .A(n1083), .B(n1084), .ZN(n1071) );
NOR2_X1 U770 ( .A1(G472), .A2(KEYINPUT63), .ZN(n1084) );
XOR2_X1 U771 ( .A(n1085), .B(n1086), .Z(G72) );
XOR2_X1 U772 ( .A(n1087), .B(n1088), .Z(n1086) );
NOR2_X1 U773 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U774 ( .A(KEYINPUT18), .B(n1091), .Z(n1090) );
NOR2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U776 ( .A(KEYINPUT41), .B(G900), .Z(n1093) );
XOR2_X1 U777 ( .A(n1094), .B(n1095), .Z(n1089) );
NAND2_X1 U778 ( .A1(n1096), .A2(KEYINPUT57), .ZN(n1094) );
XOR2_X1 U779 ( .A(n1097), .B(n1098), .Z(n1096) );
XOR2_X1 U780 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U781 ( .A1(n1101), .A2(n1102), .ZN(n1087) );
NOR2_X1 U782 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR2_X1 U783 ( .A1(n1105), .A2(n1106), .ZN(n1085) );
XOR2_X1 U784 ( .A(KEYINPUT29), .B(G953), .Z(n1106) );
XOR2_X1 U785 ( .A(n1107), .B(n1108), .Z(G69) );
NAND2_X1 U786 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1110) );
INV_X1 U788 ( .A(n1102), .ZN(n1109) );
XOR2_X1 U789 ( .A(n1092), .B(KEYINPUT9), .Z(n1102) );
NAND2_X1 U790 ( .A1(KEYINPUT6), .A2(n1111), .ZN(n1107) );
XOR2_X1 U791 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U792 ( .A1(n1114), .A2(G953), .ZN(n1113) );
NOR2_X1 U793 ( .A1(n1115), .A2(n1116), .ZN(n1112) );
XOR2_X1 U794 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U795 ( .A1(G898), .A2(n1092), .ZN(n1115) );
NOR2_X1 U796 ( .A1(n1119), .A2(n1120), .ZN(G66) );
NOR3_X1 U797 ( .A1(n1082), .A2(n1121), .A3(n1122), .ZN(n1120) );
AND3_X1 U798 ( .A1(n1123), .A2(n1080), .A3(n1124), .ZN(n1122) );
NOR2_X1 U799 ( .A1(n1125), .A2(n1123), .ZN(n1121) );
AND2_X1 U800 ( .A1(n1039), .A2(n1080), .ZN(n1125) );
INV_X1 U801 ( .A(n1126), .ZN(n1080) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1128), .ZN(G63) );
XOR2_X1 U803 ( .A(n1129), .B(n1130), .Z(n1128) );
AND2_X1 U804 ( .A1(G478), .A2(n1124), .ZN(n1130) );
NOR2_X1 U805 ( .A1(G952), .A2(n1131), .ZN(n1127) );
XOR2_X1 U806 ( .A(KEYINPUT25), .B(G953), .Z(n1131) );
NOR2_X1 U807 ( .A1(n1119), .A2(n1132), .ZN(G60) );
NOR2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U809 ( .A(KEYINPUT26), .B(n1135), .Z(n1134) );
NOR2_X1 U810 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
AND2_X1 U811 ( .A1(n1137), .A2(n1136), .ZN(n1133) );
NAND2_X1 U812 ( .A1(n1124), .A2(G475), .ZN(n1137) );
XOR2_X1 U813 ( .A(n1138), .B(n1139), .Z(G6) );
NOR2_X1 U814 ( .A1(n1119), .A2(n1140), .ZN(G57) );
XOR2_X1 U815 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U816 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND3_X1 U817 ( .A1(n1124), .A2(G472), .A3(KEYINPUT51), .ZN(n1143) );
XNOR2_X1 U818 ( .A(G101), .B(n1145), .ZN(n1141) );
NOR2_X1 U819 ( .A1(n1119), .A2(n1146), .ZN(G54) );
XOR2_X1 U820 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U822 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U823 ( .A1(G469), .A2(n1124), .ZN(n1152) );
INV_X1 U824 ( .A(n1153), .ZN(n1124) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1147) );
XOR2_X1 U826 ( .A(KEYINPUT39), .B(G110), .Z(n1155) );
NAND2_X1 U827 ( .A1(KEYINPUT34), .A2(n1156), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1119), .A2(n1157), .ZN(G51) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U830 ( .A1(n1160), .A2(n1153), .ZN(n1159) );
NAND2_X1 U831 ( .A1(G902), .A2(n1039), .ZN(n1153) );
NAND2_X1 U832 ( .A1(n1105), .A2(n1114), .ZN(n1039) );
AND4_X1 U833 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1114) );
AND4_X1 U834 ( .A1(n1165), .A2(n1166), .A3(n1139), .A4(n1033), .ZN(n1164) );
NAND3_X1 U835 ( .A1(n1064), .A2(n1167), .A3(n1168), .ZN(n1033) );
NAND3_X1 U836 ( .A1(n1168), .A2(n1167), .A3(n1065), .ZN(n1139) );
NOR2_X1 U837 ( .A1(n1169), .A2(n1170), .ZN(n1163) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
AND3_X1 U839 ( .A1(n1173), .A2(n1168), .A3(n1062), .ZN(n1169) );
AND4_X1 U840 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1105) );
NOR4_X1 U841 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR2_X1 U842 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U843 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
NOR2_X1 U844 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U845 ( .A1(n1188), .A2(n1189), .ZN(n1184) );
XNOR2_X1 U846 ( .A(n1062), .B(KEYINPUT52), .ZN(n1188) );
INV_X1 U847 ( .A(n1190), .ZN(n1180) );
NOR4_X1 U848 ( .A1(n1191), .A2(n1192), .A3(n1060), .A4(n1186), .ZN(n1179) );
NAND2_X1 U849 ( .A1(n1068), .A2(n1187), .ZN(n1192) );
INV_X1 U850 ( .A(KEYINPUT16), .ZN(n1187) );
NOR3_X1 U851 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1178) );
NOR2_X1 U852 ( .A1(n1196), .A2(n1197), .ZN(n1176) );
NAND3_X1 U853 ( .A1(n1198), .A2(n1199), .A3(KEYINPUT19), .ZN(n1158) );
NAND2_X1 U854 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
INV_X1 U855 ( .A(KEYINPUT17), .ZN(n1201) );
XOR2_X1 U856 ( .A(n1202), .B(n1203), .Z(n1200) );
NAND3_X1 U857 ( .A1(n1202), .A2(n1203), .A3(KEYINPUT17), .ZN(n1198) );
XOR2_X1 U858 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U859 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U860 ( .A1(G125), .A2(KEYINPUT46), .ZN(n1207) );
NOR2_X1 U861 ( .A1(n1092), .A2(G952), .ZN(n1119) );
XOR2_X1 U862 ( .A(n1208), .B(n1190), .Z(G48) );
NAND2_X1 U863 ( .A1(n1209), .A2(n1065), .ZN(n1190) );
XOR2_X1 U864 ( .A(G143), .B(n1210), .Z(G45) );
NOR3_X1 U865 ( .A1(n1195), .A2(n1193), .A3(n1211), .ZN(n1210) );
XOR2_X1 U866 ( .A(n1194), .B(KEYINPUT3), .Z(n1211) );
NAND4_X1 U867 ( .A1(n1062), .A2(n1068), .A3(n1074), .A4(n1212), .ZN(n1195) );
XOR2_X1 U868 ( .A(n1156), .B(n1213), .Z(G42) );
NAND2_X1 U869 ( .A1(KEYINPUT27), .A2(n1197), .ZN(n1213) );
AND3_X1 U870 ( .A1(n1065), .A2(n1214), .A3(n1061), .ZN(n1197) );
INV_X1 U871 ( .A(G140), .ZN(n1156) );
XOR2_X1 U872 ( .A(G137), .B(n1215), .Z(G39) );
NOR2_X1 U873 ( .A1(n1183), .A2(n1186), .ZN(n1215) );
INV_X1 U874 ( .A(n1216), .ZN(n1186) );
XOR2_X1 U875 ( .A(G134), .B(n1217), .Z(G36) );
NOR2_X1 U876 ( .A1(n1183), .A2(n1172), .ZN(n1217) );
INV_X1 U877 ( .A(n1214), .ZN(n1183) );
NAND3_X1 U878 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(G33) );
OR2_X1 U879 ( .A1(G131), .A2(KEYINPUT60), .ZN(n1220) );
NAND3_X1 U880 ( .A1(KEYINPUT60), .A2(G131), .A3(n1221), .ZN(n1219) );
NAND2_X1 U881 ( .A1(n1196), .A2(n1222), .ZN(n1218) );
NAND2_X1 U882 ( .A1(KEYINPUT60), .A2(n1223), .ZN(n1222) );
XOR2_X1 U883 ( .A(KEYINPUT7), .B(G131), .Z(n1223) );
INV_X1 U884 ( .A(n1221), .ZN(n1196) );
NAND3_X1 U885 ( .A1(n1065), .A2(n1214), .A3(n1062), .ZN(n1221) );
NOR3_X1 U886 ( .A1(n1224), .A2(n1193), .A3(n1060), .ZN(n1214) );
NAND2_X1 U887 ( .A1(n1225), .A2(n1057), .ZN(n1060) );
INV_X1 U888 ( .A(n1068), .ZN(n1224) );
XNOR2_X1 U889 ( .A(G128), .B(n1174), .ZN(G30) );
NAND2_X1 U890 ( .A1(n1209), .A2(n1064), .ZN(n1174) );
AND3_X1 U891 ( .A1(n1056), .A2(n1068), .A3(n1226), .ZN(n1209) );
NOR3_X1 U892 ( .A1(n1227), .A2(n1228), .A3(n1193), .ZN(n1226) );
INV_X1 U893 ( .A(n1191), .ZN(n1193) );
XNOR2_X1 U894 ( .A(G101), .B(n1229), .ZN(G3) );
NAND3_X1 U895 ( .A1(n1168), .A2(n1230), .A3(n1062), .ZN(n1229) );
XOR2_X1 U896 ( .A(KEYINPUT58), .B(n1173), .Z(n1230) );
XOR2_X1 U897 ( .A(n1175), .B(n1231), .Z(G27) );
XOR2_X1 U898 ( .A(n1232), .B(KEYINPUT54), .Z(n1231) );
NAND4_X1 U899 ( .A1(n1233), .A2(n1061), .A3(n1065), .A4(n1191), .ZN(n1175) );
NAND2_X1 U900 ( .A1(n1234), .A2(n1235), .ZN(n1191) );
NAND2_X1 U901 ( .A1(n1236), .A2(n1104), .ZN(n1235) );
INV_X1 U902 ( .A(G900), .ZN(n1104) );
XOR2_X1 U903 ( .A(n1237), .B(n1161), .Z(G24) );
NAND4_X1 U904 ( .A1(n1238), .A2(n1167), .A3(n1074), .A4(n1212), .ZN(n1161) );
INV_X1 U905 ( .A(n1054), .ZN(n1167) );
NAND2_X1 U906 ( .A1(n1228), .A2(n1227), .ZN(n1054) );
XOR2_X1 U907 ( .A(n1162), .B(n1239), .Z(G21) );
XOR2_X1 U908 ( .A(n1240), .B(KEYINPUT30), .Z(n1239) );
NAND2_X1 U909 ( .A1(n1238), .A2(n1216), .ZN(n1162) );
NOR3_X1 U910 ( .A1(n1227), .A2(n1228), .A3(n1050), .ZN(n1216) );
XOR2_X1 U911 ( .A(G116), .B(n1241), .Z(G18) );
NOR3_X1 U912 ( .A1(n1172), .A2(KEYINPUT20), .A3(n1171), .ZN(n1241) );
NAND2_X1 U913 ( .A1(n1062), .A2(n1064), .ZN(n1172) );
INV_X1 U914 ( .A(n1189), .ZN(n1064) );
NAND2_X1 U915 ( .A1(n1070), .A2(n1074), .ZN(n1189) );
INV_X1 U916 ( .A(n1242), .ZN(n1074) );
XOR2_X1 U917 ( .A(n1166), .B(n1243), .Z(G15) );
NAND2_X1 U918 ( .A1(KEYINPUT44), .A2(G113), .ZN(n1243) );
NAND3_X1 U919 ( .A1(n1062), .A2(n1065), .A3(n1238), .ZN(n1166) );
INV_X1 U920 ( .A(n1171), .ZN(n1238) );
NAND2_X1 U921 ( .A1(n1233), .A2(n1244), .ZN(n1171) );
NOR3_X1 U922 ( .A1(n1046), .A2(n1194), .A3(n1044), .ZN(n1233) );
INV_X1 U923 ( .A(n1245), .ZN(n1044) );
AND2_X1 U924 ( .A1(n1246), .A2(n1212), .ZN(n1065) );
INV_X1 U925 ( .A(n1070), .ZN(n1212) );
NOR2_X1 U926 ( .A1(n1247), .A2(n1227), .ZN(n1062) );
XOR2_X1 U927 ( .A(n1248), .B(n1165), .Z(G12) );
NAND3_X1 U928 ( .A1(n1061), .A2(n1168), .A3(n1173), .ZN(n1165) );
INV_X1 U929 ( .A(n1050), .ZN(n1173) );
NAND2_X1 U930 ( .A1(n1246), .A2(n1070), .ZN(n1050) );
XOR2_X1 U931 ( .A(n1249), .B(G475), .Z(n1070) );
NAND2_X1 U932 ( .A1(n1136), .A2(n1250), .ZN(n1249) );
XNOR2_X1 U933 ( .A(n1251), .B(n1252), .ZN(n1136) );
XOR2_X1 U934 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U935 ( .A(n1255), .B(n1256), .ZN(n1254) );
NOR2_X1 U936 ( .A1(KEYINPUT43), .A2(n1257), .ZN(n1256) );
XOR2_X1 U937 ( .A(G146), .B(n1095), .Z(n1257) );
NOR2_X1 U938 ( .A1(KEYINPUT55), .A2(G131), .ZN(n1255) );
NAND2_X1 U939 ( .A1(n1258), .A2(G214), .ZN(n1253) );
XOR2_X1 U940 ( .A(n1259), .B(n1260), .Z(n1251) );
XOR2_X1 U941 ( .A(G113), .B(G104), .Z(n1260) );
XOR2_X1 U942 ( .A(G143), .B(n1237), .Z(n1259) );
INV_X1 U943 ( .A(G122), .ZN(n1237) );
XOR2_X1 U944 ( .A(n1242), .B(KEYINPUT37), .Z(n1246) );
XNOR2_X1 U945 ( .A(G478), .B(n1261), .ZN(n1242) );
NOR2_X1 U946 ( .A1(G902), .A2(n1129), .ZN(n1261) );
XOR2_X1 U947 ( .A(n1262), .B(n1263), .Z(n1129) );
NOR2_X1 U948 ( .A1(KEYINPUT36), .A2(n1264), .ZN(n1263) );
XOR2_X1 U949 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U950 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U951 ( .A(n1269), .B(G107), .Z(n1265) );
NAND2_X1 U952 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U953 ( .A1(G122), .A2(n1272), .ZN(n1271) );
XOR2_X1 U954 ( .A(KEYINPUT14), .B(n1273), .Z(n1270) );
NOR2_X1 U955 ( .A1(G122), .A2(n1272), .ZN(n1273) );
NAND2_X1 U956 ( .A1(G217), .A2(n1274), .ZN(n1262) );
AND3_X1 U957 ( .A1(n1068), .A2(n1244), .A3(n1056), .ZN(n1168) );
INV_X1 U958 ( .A(n1194), .ZN(n1056) );
NAND2_X1 U959 ( .A1(n1058), .A2(n1057), .ZN(n1194) );
NAND2_X1 U960 ( .A1(G214), .A2(n1275), .ZN(n1057) );
INV_X1 U961 ( .A(n1225), .ZN(n1058) );
XNOR2_X1 U962 ( .A(n1276), .B(n1160), .ZN(n1225) );
NAND2_X1 U963 ( .A1(G210), .A2(n1275), .ZN(n1160) );
NAND2_X1 U964 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
INV_X1 U965 ( .A(G237), .ZN(n1278) );
NAND2_X1 U966 ( .A1(n1279), .A2(n1250), .ZN(n1276) );
XOR2_X1 U967 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U968 ( .A(n1204), .B(n1202), .Z(n1281) );
NAND2_X1 U969 ( .A1(n1282), .A2(n1283), .ZN(n1202) );
NAND2_X1 U970 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
INV_X1 U971 ( .A(KEYINPUT15), .ZN(n1285) );
XNOR2_X1 U972 ( .A(n1117), .B(n1118), .ZN(n1284) );
NAND2_X1 U973 ( .A1(n1286), .A2(n1287), .ZN(n1117) );
NAND2_X1 U974 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U975 ( .A1(n1290), .A2(KEYINPUT15), .ZN(n1282) );
XNOR2_X1 U976 ( .A(n1286), .B(n1118), .ZN(n1290) );
XNOR2_X1 U977 ( .A(n1291), .B(n1292), .ZN(n1118) );
XOR2_X1 U978 ( .A(KEYINPUT21), .B(G122), .Z(n1292) );
NAND2_X1 U979 ( .A1(KEYINPUT5), .A2(n1248), .ZN(n1291) );
OR2_X1 U980 ( .A1(n1289), .A2(n1288), .ZN(n1286) );
NAND2_X1 U981 ( .A1(n1293), .A2(n1294), .ZN(n1288) );
NAND2_X1 U982 ( .A1(n1295), .A2(KEYINPUT28), .ZN(n1294) );
NAND2_X1 U983 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
INV_X1 U984 ( .A(KEYINPUT28), .ZN(n1297) );
NAND2_X1 U985 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
NAND2_X1 U986 ( .A1(G113), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U987 ( .A(n1301), .B(n1302), .ZN(n1289) );
XOR2_X1 U988 ( .A(G107), .B(G101), .Z(n1302) );
NAND2_X1 U989 ( .A1(KEYINPUT0), .A2(n1138), .ZN(n1301) );
INV_X1 U990 ( .A(G104), .ZN(n1138) );
XOR2_X1 U991 ( .A(n1206), .B(n1303), .Z(n1280) );
NOR2_X1 U992 ( .A1(KEYINPUT48), .A2(n1232), .ZN(n1303) );
INV_X1 U993 ( .A(G125), .ZN(n1232) );
AND2_X1 U994 ( .A1(G224), .A2(n1092), .ZN(n1206) );
NAND2_X1 U995 ( .A1(n1234), .A2(n1304), .ZN(n1244) );
NAND2_X1 U996 ( .A1(n1236), .A2(n1305), .ZN(n1304) );
INV_X1 U997 ( .A(G898), .ZN(n1305) );
NOR3_X1 U998 ( .A1(n1250), .A2(n1040), .A3(n1092), .ZN(n1236) );
INV_X1 U999 ( .A(n1306), .ZN(n1040) );
NAND3_X1 U1000 ( .A1(n1306), .A2(n1092), .A3(G952), .ZN(n1234) );
NAND2_X1 U1001 ( .A1(G237), .A2(n1307), .ZN(n1306) );
NOR2_X1 U1002 ( .A1(n1046), .A2(n1245), .ZN(n1068) );
XOR2_X1 U1003 ( .A(n1308), .B(G469), .Z(n1245) );
NAND2_X1 U1004 ( .A1(n1309), .A2(n1250), .ZN(n1308) );
XOR2_X1 U1005 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1006 ( .A(n1312), .B(n1151), .Z(n1311) );
XNOR2_X1 U1007 ( .A(n1313), .B(n1314), .ZN(n1151) );
NOR2_X1 U1008 ( .A1(G953), .A2(n1103), .ZN(n1314) );
INV_X1 U1009 ( .A(G227), .ZN(n1103) );
NAND2_X1 U1010 ( .A1(KEYINPUT10), .A2(n1149), .ZN(n1312) );
XOR2_X1 U1011 ( .A(n1315), .B(n1316), .Z(n1149) );
XOR2_X1 U1012 ( .A(n1317), .B(n1097), .Z(n1316) );
NAND2_X1 U1013 ( .A1(n1318), .A2(n1319), .ZN(n1097) );
NAND2_X1 U1014 ( .A1(n1320), .A2(n1208), .ZN(n1319) );
XOR2_X1 U1015 ( .A(KEYINPUT50), .B(n1267), .Z(n1320) );
NAND2_X1 U1016 ( .A1(n1321), .A2(n1322), .ZN(n1317) );
NAND2_X1 U1017 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1018 ( .A(KEYINPUT11), .B(G104), .Z(n1324) );
XNOR2_X1 U1019 ( .A(n1325), .B(KEYINPUT56), .ZN(n1323) );
XOR2_X1 U1020 ( .A(n1326), .B(KEYINPUT32), .Z(n1321) );
NAND2_X1 U1021 ( .A1(G104), .A2(n1325), .ZN(n1326) );
XNOR2_X1 U1022 ( .A(n1327), .B(KEYINPUT49), .ZN(n1325) );
INV_X1 U1023 ( .A(G107), .ZN(n1327) );
XNOR2_X1 U1024 ( .A(G101), .B(KEYINPUT62), .ZN(n1315) );
XOR2_X1 U1025 ( .A(G140), .B(G110), .Z(n1310) );
XNOR2_X1 U1026 ( .A(n1069), .B(KEYINPUT45), .ZN(n1046) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1328), .ZN(n1069) );
AND2_X1 U1028 ( .A1(n1227), .A2(n1247), .ZN(n1061) );
INV_X1 U1029 ( .A(n1228), .ZN(n1247) );
NOR2_X1 U1030 ( .A1(n1329), .A2(n1078), .ZN(n1228) );
NOR2_X1 U1031 ( .A1(n1126), .A2(n1082), .ZN(n1078) );
AND2_X1 U1032 ( .A1(n1082), .A2(n1126), .ZN(n1329) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1328), .ZN(n1126) );
NAND2_X1 U1034 ( .A1(n1307), .A2(n1277), .ZN(n1328) );
XOR2_X1 U1035 ( .A(G902), .B(KEYINPUT33), .Z(n1277) );
XNOR2_X1 U1036 ( .A(G234), .B(KEYINPUT13), .ZN(n1307) );
NOR2_X1 U1037 ( .A1(n1123), .A2(G902), .ZN(n1082) );
XOR2_X1 U1038 ( .A(n1330), .B(n1331), .Z(n1123) );
XOR2_X1 U1039 ( .A(n1332), .B(n1333), .Z(n1331) );
NAND2_X1 U1040 ( .A1(KEYINPUT59), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1041 ( .A(G137), .B(n1335), .ZN(n1334) );
NAND2_X1 U1042 ( .A1(n1274), .A2(G221), .ZN(n1335) );
AND2_X1 U1043 ( .A1(G234), .A2(n1092), .ZN(n1274) );
INV_X1 U1044 ( .A(G953), .ZN(n1092) );
NAND2_X1 U1045 ( .A1(n1336), .A2(KEYINPUT40), .ZN(n1332) );
XOR2_X1 U1046 ( .A(n1208), .B(n1095), .Z(n1336) );
XOR2_X1 U1047 ( .A(G125), .B(G140), .Z(n1095) );
NAND2_X1 U1048 ( .A1(n1337), .A2(n1338), .ZN(n1330) );
NAND2_X1 U1049 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NAND2_X1 U1050 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1051 ( .A1(G110), .A2(n1343), .ZN(n1342) );
INV_X1 U1052 ( .A(KEYINPUT31), .ZN(n1341) );
NAND2_X1 U1053 ( .A1(n1344), .A2(n1248), .ZN(n1337) );
NAND2_X1 U1054 ( .A1(n1343), .A2(n1345), .ZN(n1344) );
OR2_X1 U1055 ( .A1(n1339), .A2(KEYINPUT31), .ZN(n1345) );
XOR2_X1 U1056 ( .A(n1240), .B(n1346), .Z(n1339) );
XOR2_X1 U1057 ( .A(KEYINPUT22), .B(G128), .Z(n1346) );
INV_X1 U1058 ( .A(KEYINPUT42), .ZN(n1343) );
XOR2_X1 U1059 ( .A(n1083), .B(G472), .Z(n1227) );
NAND2_X1 U1060 ( .A1(n1347), .A2(n1250), .ZN(n1083) );
INV_X1 U1061 ( .A(G902), .ZN(n1250) );
XOR2_X1 U1062 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1063 ( .A(KEYINPUT8), .B(G101), .Z(n1349) );
XOR2_X1 U1064 ( .A(n1350), .B(n1351), .Z(n1348) );
INV_X1 U1065 ( .A(n1144), .ZN(n1351) );
XNOR2_X1 U1066 ( .A(n1352), .B(n1204), .ZN(n1144) );
NAND2_X1 U1067 ( .A1(n1318), .A2(n1353), .ZN(n1204) );
NAND2_X1 U1068 ( .A1(n1354), .A2(n1208), .ZN(n1353) );
INV_X1 U1069 ( .A(G146), .ZN(n1208) );
XOR2_X1 U1070 ( .A(KEYINPUT24), .B(n1267), .Z(n1354) );
NAND2_X1 U1071 ( .A1(n1267), .A2(G146), .ZN(n1318) );
XOR2_X1 U1072 ( .A(G128), .B(G143), .Z(n1267) );
XNOR2_X1 U1073 ( .A(n1295), .B(n1313), .ZN(n1352) );
XNOR2_X1 U1074 ( .A(n1099), .B(n1355), .ZN(n1313) );
NOR2_X1 U1075 ( .A1(KEYINPUT38), .A2(n1100), .ZN(n1355) );
XOR2_X1 U1076 ( .A(G131), .B(KEYINPUT4), .Z(n1100) );
XNOR2_X1 U1077 ( .A(G137), .B(n1268), .ZN(n1099) );
XOR2_X1 U1078 ( .A(G134), .B(KEYINPUT53), .Z(n1268) );
AND3_X1 U1079 ( .A1(n1356), .A2(n1357), .A3(n1298), .ZN(n1295) );
OR2_X1 U1080 ( .A1(n1300), .A2(G113), .ZN(n1298) );
OR2_X1 U1081 ( .A1(n1358), .A2(G119), .ZN(n1300) );
NAND2_X1 U1082 ( .A1(G119), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1083 ( .A(G113), .B(n1358), .Z(n1359) );
NAND3_X1 U1084 ( .A1(G113), .A2(n1358), .A3(n1240), .ZN(n1356) );
INV_X1 U1085 ( .A(G119), .ZN(n1240) );
XOR2_X1 U1086 ( .A(n1272), .B(KEYINPUT61), .Z(n1358) );
INV_X1 U1087 ( .A(G116), .ZN(n1272) );
NAND2_X1 U1088 ( .A1(n1360), .A2(KEYINPUT1), .ZN(n1350) );
XOR2_X1 U1089 ( .A(n1145), .B(KEYINPUT35), .Z(n1360) );
NAND2_X1 U1090 ( .A1(n1258), .A2(G210), .ZN(n1145) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1258) );
INV_X1 U1092 ( .A(G110), .ZN(n1248) );
endmodule


