//Key = 1110100111000111111010011011010010010000110000000101010110111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340;

XNOR2_X1 U732 ( .A(n1010), .B(n1011), .ZN(G9) );
XNOR2_X1 U733 ( .A(G107), .B(KEYINPUT47), .ZN(n1011) );
NOR2_X1 U734 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
NAND3_X1 U736 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1014) );
NAND2_X1 U737 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U738 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND3_X1 U739 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
OR2_X1 U740 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND2_X1 U741 ( .A1(n1030), .A2(n1029), .ZN(n1025) );
OR4_X1 U742 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(KEYINPUT17), .ZN(n1030) );
NAND2_X1 U743 ( .A1(KEYINPUT6), .A2(n1034), .ZN(n1023) );
NAND4_X1 U744 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
NAND3_X1 U745 ( .A1(n1037), .A2(n1039), .A3(n1035), .ZN(n1018) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U747 ( .A1(n1027), .A2(n1042), .ZN(n1041) );
NAND2_X1 U748 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND4_X1 U749 ( .A1(KEYINPUT17), .A2(n1021), .A3(n1045), .A4(n1046), .ZN(n1044) );
NAND3_X1 U750 ( .A1(n1028), .A2(n1047), .A3(n1048), .ZN(n1043) );
INV_X1 U751 ( .A(KEYINPUT55), .ZN(n1047) );
NAND4_X1 U752 ( .A1(n1021), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1028) );
NAND2_X1 U753 ( .A1(n1036), .A2(n1052), .ZN(n1051) );
NAND2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
OR2_X1 U755 ( .A1(n1055), .A2(KEYINPUT31), .ZN(n1054) );
NAND3_X1 U756 ( .A1(KEYINPUT31), .A2(n1056), .A3(n1057), .ZN(n1050) );
NAND3_X1 U757 ( .A1(n1037), .A2(n1048), .A3(KEYINPUT55), .ZN(n1049) );
NAND2_X1 U758 ( .A1(n1036), .A2(n1058), .ZN(n1040) );
NAND2_X1 U759 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U760 ( .A1(n1021), .A2(n1061), .ZN(n1060) );
NAND2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
OR2_X1 U762 ( .A1(n1064), .A2(KEYINPUT6), .ZN(n1063) );
NAND2_X1 U763 ( .A1(n1027), .A2(n1065), .ZN(n1059) );
NAND2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR3_X1 U766 ( .A1(n1017), .A2(G952), .A3(n1070), .ZN(n1012) );
INV_X1 U767 ( .A(n1019), .ZN(n1070) );
NAND4_X1 U768 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1019) );
NOR4_X1 U769 ( .A1(n1046), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1074) );
XOR2_X1 U770 ( .A(n1078), .B(n1079), .Z(n1076) );
NOR2_X1 U771 ( .A1(n1080), .A2(KEYINPUT39), .ZN(n1079) );
NOR2_X1 U772 ( .A1(n1081), .A2(n1082), .ZN(n1075) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1031), .ZN(n1073) );
XOR2_X1 U774 ( .A(n1084), .B(KEYINPUT56), .Z(n1072) );
NAND2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U776 ( .A(n1087), .B(KEYINPUT57), .Z(n1085) );
XOR2_X1 U777 ( .A(n1088), .B(KEYINPUT61), .Z(n1071) );
XOR2_X1 U778 ( .A(n1089), .B(n1090), .Z(G72) );
NOR2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(n1089) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1092), .ZN(n1094) );
XOR2_X1 U783 ( .A(n1096), .B(n1015), .Z(n1095) );
NAND3_X1 U784 ( .A1(n1096), .A2(G900), .A3(G953), .ZN(n1093) );
NOR2_X1 U785 ( .A1(KEYINPUT28), .A2(n1097), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(n1097) );
XNOR2_X1 U787 ( .A(n1100), .B(n1101), .ZN(n1099) );
XOR2_X1 U788 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U789 ( .A(n1104), .B(n1105), .Z(n1098) );
XNOR2_X1 U790 ( .A(KEYINPUT40), .B(KEYINPUT16), .ZN(n1105) );
NAND2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(G69) );
NAND2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U793 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND3_X1 U794 ( .A1(G953), .A2(n1111), .A3(n1112), .ZN(n1106) );
XNOR2_X1 U795 ( .A(n1108), .B(KEYINPUT54), .ZN(n1112) );
XNOR2_X1 U796 ( .A(n1113), .B(n1114), .ZN(n1108) );
NOR2_X1 U797 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U798 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U799 ( .A1(KEYINPUT50), .A2(n1119), .ZN(n1118) );
NOR2_X1 U800 ( .A1(G898), .A2(n1092), .ZN(n1115) );
NAND2_X1 U801 ( .A1(n1092), .A2(n1016), .ZN(n1113) );
NAND2_X1 U802 ( .A1(G898), .A2(G224), .ZN(n1111) );
NOR3_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(G66) );
AND2_X1 U804 ( .A1(KEYINPUT0), .A2(n1123), .ZN(n1122) );
NOR3_X1 U805 ( .A1(KEYINPUT0), .A2(G952), .A3(n1124), .ZN(n1121) );
XOR2_X1 U806 ( .A(n1125), .B(n1126), .Z(n1120) );
NOR2_X1 U807 ( .A1(n1078), .A2(n1127), .ZN(n1126) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1128), .ZN(G63) );
XOR2_X1 U809 ( .A(n1129), .B(n1130), .Z(n1128) );
AND2_X1 U810 ( .A1(G478), .A2(n1131), .ZN(n1129) );
NOR2_X1 U811 ( .A1(n1123), .A2(n1132), .ZN(G60) );
XOR2_X1 U812 ( .A(n1133), .B(n1134), .Z(n1132) );
AND2_X1 U813 ( .A1(G475), .A2(n1131), .ZN(n1133) );
XNOR2_X1 U814 ( .A(G104), .B(n1135), .ZN(G6) );
NAND4_X1 U815 ( .A1(KEYINPUT24), .A2(n1056), .A3(n1136), .A4(n1027), .ZN(n1135) );
NOR2_X1 U816 ( .A1(n1123), .A2(n1137), .ZN(G57) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U818 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NAND2_X1 U819 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XOR2_X1 U820 ( .A(n1144), .B(KEYINPUT34), .Z(n1142) );
NAND2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(n1140) );
XOR2_X1 U822 ( .A(n1144), .B(KEYINPUT9), .Z(n1146) );
NAND2_X1 U823 ( .A1(n1131), .A2(G472), .ZN(n1144) );
INV_X1 U824 ( .A(n1143), .ZN(n1145) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1143) );
NOR2_X1 U826 ( .A1(KEYINPUT48), .A2(n1149), .ZN(n1148) );
NOR2_X1 U827 ( .A1(n1123), .A2(n1150), .ZN(G54) );
XOR2_X1 U828 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U829 ( .A1(G469), .A2(n1131), .ZN(n1152) );
INV_X1 U830 ( .A(n1127), .ZN(n1131) );
NAND2_X1 U831 ( .A1(n1153), .A2(KEYINPUT20), .ZN(n1151) );
XOR2_X1 U832 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U833 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U834 ( .A(n1158), .B(n1159), .Z(n1156) );
XOR2_X1 U835 ( .A(n1160), .B(n1161), .Z(n1154) );
XNOR2_X1 U836 ( .A(n1162), .B(n1163), .ZN(n1161) );
NOR2_X1 U837 ( .A1(KEYINPUT38), .A2(n1164), .ZN(n1163) );
XOR2_X1 U838 ( .A(KEYINPUT62), .B(n1165), .Z(n1164) );
NAND2_X1 U839 ( .A1(KEYINPUT32), .A2(n1166), .ZN(n1162) );
XNOR2_X1 U840 ( .A(KEYINPUT8), .B(KEYINPUT5), .ZN(n1160) );
NOR2_X1 U841 ( .A1(n1123), .A2(n1167), .ZN(G51) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U844 ( .A(n1172), .B(n1173), .Z(n1168) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1127), .ZN(n1173) );
NAND2_X1 U846 ( .A1(G902), .A2(n1175), .ZN(n1127) );
OR2_X1 U847 ( .A1(n1015), .A2(n1016), .ZN(n1175) );
NAND4_X1 U848 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1016) );
NOR4_X1 U849 ( .A1(n1010), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1179) );
AND3_X1 U850 ( .A1(n1183), .A2(n1027), .A3(n1136), .ZN(n1010) );
NAND2_X1 U851 ( .A1(n1056), .A2(n1184), .ZN(n1178) );
NAND3_X1 U852 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NAND3_X1 U853 ( .A1(n1188), .A2(n1189), .A3(n1027), .ZN(n1187) );
NAND2_X1 U854 ( .A1(KEYINPUT60), .A2(n1190), .ZN(n1189) );
NAND2_X1 U855 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
INV_X1 U856 ( .A(KEYINPUT60), .ZN(n1192) );
NAND3_X1 U857 ( .A1(n1048), .A2(n1193), .A3(n1194), .ZN(n1191) );
NAND4_X1 U858 ( .A1(n1195), .A2(n1066), .A3(n1196), .A4(n1197), .ZN(n1186) );
INV_X1 U859 ( .A(KEYINPUT26), .ZN(n1197) );
NOR2_X1 U860 ( .A1(n1064), .A2(n1057), .ZN(n1196) );
NAND2_X1 U861 ( .A1(KEYINPUT26), .A2(n1198), .ZN(n1185) );
NAND3_X1 U862 ( .A1(n1199), .A2(n1027), .A3(n1200), .ZN(n1177) );
NAND3_X1 U863 ( .A1(n1038), .A2(n1136), .A3(n1037), .ZN(n1176) );
INV_X1 U864 ( .A(n1190), .ZN(n1136) );
NAND4_X1 U865 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1015) );
NOR4_X1 U866 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1204) );
NOR3_X1 U867 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1203) );
NOR4_X1 U868 ( .A1(n1212), .A2(n1213), .A3(n1062), .A4(n1057), .ZN(n1211) );
NAND3_X1 U869 ( .A1(n1214), .A2(n1055), .A3(n1193), .ZN(n1213) );
INV_X1 U870 ( .A(KEYINPUT36), .ZN(n1212) );
NOR2_X1 U871 ( .A1(KEYINPUT36), .A2(n1215), .ZN(n1210) );
NOR3_X1 U872 ( .A1(n1216), .A2(n1217), .A3(n1053), .ZN(n1209) );
INV_X1 U873 ( .A(n1183), .ZN(n1053) );
XOR2_X1 U874 ( .A(n1083), .B(KEYINPUT42), .Z(n1217) );
NAND2_X1 U875 ( .A1(KEYINPUT51), .A2(n1218), .ZN(n1172) );
AND2_X1 U876 ( .A1(n1124), .A2(n1219), .ZN(n1123) );
XOR2_X1 U877 ( .A(G953), .B(KEYINPUT37), .Z(n1124) );
XOR2_X1 U878 ( .A(n1202), .B(n1220), .Z(G48) );
NAND2_X1 U879 ( .A1(KEYINPUT29), .A2(G146), .ZN(n1220) );
NAND3_X1 U880 ( .A1(n1221), .A2(n1193), .A3(n1056), .ZN(n1202) );
XOR2_X1 U881 ( .A(G143), .B(n1208), .Z(G45) );
AND3_X1 U882 ( .A1(n1222), .A2(n1193), .A3(n1199), .ZN(n1208) );
XOR2_X1 U883 ( .A(G140), .B(n1223), .Z(G42) );
NOR2_X1 U884 ( .A1(KEYINPUT19), .A2(n1201), .ZN(n1223) );
NAND3_X1 U885 ( .A1(n1021), .A2(n1048), .A3(n1224), .ZN(n1201) );
XOR2_X1 U886 ( .A(G137), .B(n1207), .Z(G39) );
AND3_X1 U887 ( .A1(n1221), .A2(n1021), .A3(n1037), .ZN(n1207) );
XOR2_X1 U888 ( .A(n1225), .B(n1226), .Z(G36) );
NAND3_X1 U889 ( .A1(n1021), .A2(n1183), .A3(n1222), .ZN(n1226) );
INV_X1 U890 ( .A(n1216), .ZN(n1222) );
INV_X1 U891 ( .A(n1083), .ZN(n1021) );
XOR2_X1 U892 ( .A(G131), .B(n1206), .Z(G33) );
NOR3_X1 U893 ( .A1(n1216), .A2(n1083), .A3(n1055), .ZN(n1206) );
NAND2_X1 U894 ( .A1(n1069), .A2(n1227), .ZN(n1083) );
NAND3_X1 U895 ( .A1(n1048), .A2(n1214), .A3(n1038), .ZN(n1216) );
XOR2_X1 U896 ( .A(G128), .B(n1205), .Z(G30) );
AND3_X1 U897 ( .A1(n1183), .A2(n1193), .A3(n1221), .ZN(n1205) );
AND4_X1 U898 ( .A1(n1048), .A2(n1228), .A3(n1214), .A4(n1229), .ZN(n1221) );
XOR2_X1 U899 ( .A(G101), .B(n1230), .Z(G3) );
NOR4_X1 U900 ( .A1(KEYINPUT10), .A2(n1190), .A3(n1064), .A4(n1032), .ZN(n1230) );
XOR2_X1 U901 ( .A(n1215), .B(n1231), .Z(G27) );
NAND2_X1 U902 ( .A1(KEYINPUT1), .A2(G125), .ZN(n1231) );
NAND3_X1 U903 ( .A1(n1224), .A2(n1193), .A3(n1036), .ZN(n1215) );
INV_X1 U904 ( .A(n1057), .ZN(n1036) );
AND3_X1 U905 ( .A1(n1232), .A2(n1214), .A3(n1056), .ZN(n1224) );
NAND2_X1 U906 ( .A1(n1233), .A2(n1029), .ZN(n1214) );
XOR2_X1 U907 ( .A(KEYINPUT53), .B(n1234), .Z(n1233) );
NOR4_X1 U908 ( .A1(G900), .A2(n1235), .A3(n1236), .A4(n1092), .ZN(n1234) );
XOR2_X1 U909 ( .A(n1237), .B(n1238), .Z(G24) );
XOR2_X1 U910 ( .A(KEYINPUT18), .B(G122), .Z(n1238) );
NAND3_X1 U911 ( .A1(n1239), .A2(n1027), .A3(n1200), .ZN(n1237) );
NAND2_X1 U912 ( .A1(n1240), .A2(n1241), .ZN(n1027) );
NAND2_X1 U913 ( .A1(n1232), .A2(n1242), .ZN(n1241) );
OR3_X1 U914 ( .A1(n1229), .A2(n1228), .A3(n1242), .ZN(n1240) );
XOR2_X1 U915 ( .A(KEYINPUT3), .B(n1199), .Z(n1239) );
AND2_X1 U916 ( .A1(n1077), .A2(n1243), .ZN(n1199) );
XOR2_X1 U917 ( .A(n1182), .B(n1244), .Z(G21) );
NOR2_X1 U918 ( .A1(KEYINPUT11), .A2(n1245), .ZN(n1244) );
AND4_X1 U919 ( .A1(n1200), .A2(n1037), .A3(n1228), .A4(n1229), .ZN(n1182) );
INV_X1 U920 ( .A(n1246), .ZN(n1228) );
XOR2_X1 U921 ( .A(G116), .B(n1181), .Z(G18) );
AND2_X1 U922 ( .A1(n1198), .A2(n1183), .ZN(n1181) );
NOR2_X1 U923 ( .A1(n1243), .A2(n1247), .ZN(n1183) );
XNOR2_X1 U924 ( .A(G113), .B(n1248), .ZN(G15) );
NAND2_X1 U925 ( .A1(n1198), .A2(n1056), .ZN(n1248) );
INV_X1 U926 ( .A(n1055), .ZN(n1056) );
NAND2_X1 U927 ( .A1(n1247), .A2(n1243), .ZN(n1055) );
AND2_X1 U928 ( .A1(n1200), .A2(n1038), .ZN(n1198) );
INV_X1 U929 ( .A(n1064), .ZN(n1038) );
NAND2_X1 U930 ( .A1(n1249), .A2(n1229), .ZN(n1064) );
XOR2_X1 U931 ( .A(n1242), .B(n1246), .Z(n1249) );
INV_X1 U932 ( .A(KEYINPUT63), .ZN(n1242) );
NOR3_X1 U933 ( .A1(n1066), .A2(n1194), .A3(n1057), .ZN(n1200) );
NAND2_X1 U934 ( .A1(n1045), .A2(n1250), .ZN(n1057) );
INV_X1 U935 ( .A(n1195), .ZN(n1194) );
INV_X1 U936 ( .A(n1193), .ZN(n1066) );
XOR2_X1 U937 ( .A(G110), .B(n1180), .Z(G12) );
NOR3_X1 U938 ( .A1(n1190), .A2(n1062), .A3(n1032), .ZN(n1180) );
INV_X1 U939 ( .A(n1037), .ZN(n1032) );
NOR2_X1 U940 ( .A1(n1077), .A2(n1243), .ZN(n1037) );
NAND2_X1 U941 ( .A1(n1088), .A2(n1251), .ZN(n1243) );
OR2_X1 U942 ( .A1(n1082), .A2(n1081), .ZN(n1251) );
NAND2_X1 U943 ( .A1(n1081), .A2(n1082), .ZN(n1088) );
XOR2_X1 U944 ( .A(G475), .B(KEYINPUT15), .Z(n1082) );
NOR2_X1 U945 ( .A1(n1134), .A2(n1252), .ZN(n1081) );
XNOR2_X1 U946 ( .A(n1253), .B(n1254), .ZN(n1134) );
XOR2_X1 U947 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U948 ( .A(G113), .B(G104), .Z(n1256) );
XOR2_X1 U949 ( .A(G125), .B(G122), .Z(n1255) );
XOR2_X1 U950 ( .A(n1257), .B(n1258), .Z(n1253) );
XOR2_X1 U951 ( .A(n1259), .B(n1260), .Z(n1258) );
NOR2_X1 U952 ( .A1(KEYINPUT12), .A2(n1166), .ZN(n1260) );
AND2_X1 U953 ( .A1(G214), .A2(n1261), .ZN(n1259) );
XNOR2_X1 U954 ( .A(n1262), .B(n1263), .ZN(n1257) );
NAND2_X1 U955 ( .A1(KEYINPUT59), .A2(n1104), .ZN(n1262) );
INV_X1 U956 ( .A(n1247), .ZN(n1077) );
XOR2_X1 U957 ( .A(n1264), .B(G478), .Z(n1247) );
OR2_X1 U958 ( .A1(n1130), .A2(n1252), .ZN(n1264) );
XNOR2_X1 U959 ( .A(n1265), .B(n1266), .ZN(n1130) );
XOR2_X1 U960 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U961 ( .A(G122), .B(G116), .Z(n1268) );
XOR2_X1 U962 ( .A(G134), .B(G128), .Z(n1267) );
XOR2_X1 U963 ( .A(n1269), .B(n1270), .Z(n1265) );
XOR2_X1 U964 ( .A(n1271), .B(G107), .Z(n1269) );
NAND2_X1 U965 ( .A1(G217), .A2(n1272), .ZN(n1271) );
INV_X1 U966 ( .A(n1232), .ZN(n1062) );
NOR2_X1 U967 ( .A1(n1229), .A2(n1246), .ZN(n1232) );
XNOR2_X1 U968 ( .A(n1273), .B(n1078), .ZN(n1246) );
NAND2_X1 U969 ( .A1(G217), .A2(n1274), .ZN(n1078) );
XNOR2_X1 U970 ( .A(n1080), .B(KEYINPUT30), .ZN(n1273) );
NOR2_X1 U971 ( .A1(n1125), .A2(n1252), .ZN(n1080) );
INV_X1 U972 ( .A(n1275), .ZN(n1252) );
NAND2_X1 U973 ( .A1(n1276), .A2(n1277), .ZN(n1125) );
NAND2_X1 U974 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U975 ( .A(KEYINPUT7), .B(n1280), .Z(n1278) );
NAND2_X1 U976 ( .A1(n1281), .A2(n1282), .ZN(n1276) );
INV_X1 U977 ( .A(n1279), .ZN(n1282) );
XOR2_X1 U978 ( .A(n1283), .B(n1284), .Z(n1279) );
XNOR2_X1 U979 ( .A(G110), .B(n1285), .ZN(n1284) );
NAND2_X1 U980 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
OR2_X1 U981 ( .A1(n1103), .A2(n1288), .ZN(n1287) );
XOR2_X1 U982 ( .A(n1289), .B(KEYINPUT52), .Z(n1286) );
NAND2_X1 U983 ( .A1(n1288), .A2(n1103), .ZN(n1289) );
XOR2_X1 U984 ( .A(n1166), .B(n1218), .Z(n1103) );
INV_X1 U985 ( .A(G140), .ZN(n1166) );
XOR2_X1 U986 ( .A(n1245), .B(G128), .Z(n1283) );
INV_X1 U987 ( .A(G119), .ZN(n1245) );
XOR2_X1 U988 ( .A(KEYINPUT33), .B(n1280), .Z(n1281) );
AND2_X1 U989 ( .A1(n1290), .A2(n1291), .ZN(n1280) );
NAND3_X1 U990 ( .A1(G221), .A2(G137), .A3(n1272), .ZN(n1291) );
NAND2_X1 U991 ( .A1(n1292), .A2(n1293), .ZN(n1290) );
NAND2_X1 U992 ( .A1(n1272), .A2(G221), .ZN(n1293) );
AND2_X1 U993 ( .A1(G234), .A2(n1092), .ZN(n1272) );
XNOR2_X1 U994 ( .A(G137), .B(KEYINPUT43), .ZN(n1292) );
NAND2_X1 U995 ( .A1(n1086), .A2(n1087), .ZN(n1229) );
NAND3_X1 U996 ( .A1(n1275), .A2(n1294), .A3(n1295), .ZN(n1087) );
XOR2_X1 U997 ( .A(KEYINPUT2), .B(G472), .Z(n1294) );
NAND2_X1 U998 ( .A1(n1296), .A2(n1297), .ZN(n1086) );
NAND2_X1 U999 ( .A1(n1295), .A2(n1275), .ZN(n1297) );
XOR2_X1 U1000 ( .A(n1147), .B(n1298), .Z(n1295) );
XNOR2_X1 U1001 ( .A(n1299), .B(n1139), .ZN(n1298) );
XOR2_X1 U1002 ( .A(n1300), .B(n1301), .Z(n1139) );
NAND2_X1 U1003 ( .A1(n1261), .A2(G210), .ZN(n1300) );
NOR2_X1 U1004 ( .A1(G953), .A2(G237), .ZN(n1261) );
NAND2_X1 U1005 ( .A1(KEYINPUT23), .A2(n1149), .ZN(n1299) );
INV_X1 U1006 ( .A(n1158), .ZN(n1149) );
XOR2_X1 U1007 ( .A(n1302), .B(n1303), .Z(n1147) );
XOR2_X1 U1008 ( .A(n1304), .B(n1171), .Z(n1303) );
XNOR2_X1 U1009 ( .A(G113), .B(KEYINPUT13), .ZN(n1302) );
XNOR2_X1 U1010 ( .A(G472), .B(KEYINPUT2), .ZN(n1296) );
NAND3_X1 U1011 ( .A1(n1193), .A2(n1195), .A3(n1048), .ZN(n1190) );
AND2_X1 U1012 ( .A1(n1250), .A2(n1031), .ZN(n1048) );
INV_X1 U1013 ( .A(n1045), .ZN(n1031) );
XOR2_X1 U1014 ( .A(n1305), .B(G469), .Z(n1045) );
NAND2_X1 U1015 ( .A1(n1275), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1016 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1017 ( .A(n1309), .B(n1157), .Z(n1308) );
XOR2_X1 U1018 ( .A(n1102), .B(n1310), .Z(n1157) );
NAND2_X1 U1019 ( .A1(n1311), .A2(n1312), .ZN(n1102) );
NAND2_X1 U1020 ( .A1(n1263), .A2(n1313), .ZN(n1312) );
NAND2_X1 U1021 ( .A1(G128), .A2(n1314), .ZN(n1313) );
OR2_X1 U1022 ( .A1(KEYINPUT46), .A2(KEYINPUT49), .ZN(n1314) );
NAND3_X1 U1023 ( .A1(n1315), .A2(n1316), .A3(KEYINPUT49), .ZN(n1311) );
OR2_X1 U1024 ( .A1(G128), .A2(KEYINPUT46), .ZN(n1316) );
NAND2_X1 U1025 ( .A1(G128), .A2(n1317), .ZN(n1315) );
OR2_X1 U1026 ( .A1(n1263), .A2(KEYINPUT46), .ZN(n1317) );
XOR2_X1 U1027 ( .A(n1318), .B(n1165), .Z(n1309) );
AND2_X1 U1028 ( .A1(G227), .A2(n1092), .ZN(n1165) );
NAND2_X1 U1029 ( .A1(KEYINPUT4), .A2(G110), .ZN(n1318) );
XOR2_X1 U1030 ( .A(n1319), .B(n1320), .Z(n1307) );
NOR2_X1 U1031 ( .A1(KEYINPUT22), .A2(n1158), .ZN(n1320) );
XOR2_X1 U1032 ( .A(n1104), .B(n1321), .Z(n1158) );
NOR2_X1 U1033 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NOR3_X1 U1034 ( .A1(KEYINPUT27), .A2(G137), .A3(n1225), .ZN(n1323) );
NOR2_X1 U1035 ( .A1(n1100), .A2(n1324), .ZN(n1322) );
INV_X1 U1036 ( .A(KEYINPUT27), .ZN(n1324) );
XNOR2_X1 U1037 ( .A(n1225), .B(G137), .ZN(n1100) );
INV_X1 U1038 ( .A(G134), .ZN(n1225) );
INV_X1 U1039 ( .A(G131), .ZN(n1104) );
XOR2_X1 U1040 ( .A(n1301), .B(G140), .Z(n1319) );
INV_X1 U1041 ( .A(G101), .ZN(n1301) );
XOR2_X1 U1042 ( .A(KEYINPUT41), .B(n1046), .Z(n1250) );
INV_X1 U1043 ( .A(n1033), .ZN(n1046) );
NAND2_X1 U1044 ( .A1(G221), .A2(n1274), .ZN(n1033) );
NAND2_X1 U1045 ( .A1(G234), .A2(n1236), .ZN(n1274) );
NAND2_X1 U1046 ( .A1(n1029), .A2(n1325), .ZN(n1195) );
OR4_X1 U1047 ( .A1(n1092), .A2(n1236), .A3(n1235), .A4(G898), .ZN(n1325) );
INV_X1 U1048 ( .A(n1035), .ZN(n1029) );
NOR3_X1 U1049 ( .A1(n1017), .A2(n1235), .A3(n1219), .ZN(n1035) );
INV_X1 U1050 ( .A(G952), .ZN(n1219) );
AND2_X1 U1051 ( .A1(G237), .A2(G234), .ZN(n1235) );
XNOR2_X1 U1052 ( .A(n1092), .B(KEYINPUT21), .ZN(n1017) );
INV_X1 U1053 ( .A(G953), .ZN(n1092) );
NOR2_X1 U1054 ( .A1(n1069), .A2(n1068), .ZN(n1193) );
INV_X1 U1055 ( .A(n1227), .ZN(n1068) );
NAND2_X1 U1056 ( .A1(G214), .A2(n1326), .ZN(n1227) );
XNOR2_X1 U1057 ( .A(n1327), .B(n1174), .ZN(n1069) );
NAND2_X1 U1058 ( .A1(G210), .A2(n1326), .ZN(n1174) );
NAND2_X1 U1059 ( .A1(n1328), .A2(n1236), .ZN(n1326) );
INV_X1 U1060 ( .A(G237), .ZN(n1328) );
NAND2_X1 U1061 ( .A1(n1329), .A2(n1275), .ZN(n1327) );
XOR2_X1 U1062 ( .A(n1236), .B(KEYINPUT45), .Z(n1275) );
INV_X1 U1063 ( .A(G902), .ZN(n1236) );
XOR2_X1 U1064 ( .A(n1170), .B(n1330), .Z(n1329) );
NOR2_X1 U1065 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1066 ( .A(KEYINPUT25), .B(n1333), .Z(n1332) );
NOR2_X1 U1067 ( .A1(n1171), .A2(n1218), .ZN(n1333) );
INV_X1 U1068 ( .A(G125), .ZN(n1218) );
NOR2_X1 U1069 ( .A1(G125), .A2(n1334), .ZN(n1331) );
INV_X1 U1070 ( .A(n1171), .ZN(n1334) );
XNOR2_X1 U1071 ( .A(G128), .B(n1263), .ZN(n1171) );
XOR2_X1 U1072 ( .A(n1270), .B(n1288), .Z(n1263) );
XNOR2_X1 U1073 ( .A(G146), .B(KEYINPUT35), .ZN(n1288) );
XOR2_X1 U1074 ( .A(G143), .B(KEYINPUT58), .Z(n1270) );
XOR2_X1 U1075 ( .A(n1335), .B(n1119), .Z(n1170) );
XNOR2_X1 U1076 ( .A(n1336), .B(G113), .ZN(n1119) );
NAND2_X1 U1077 ( .A1(KEYINPUT14), .A2(n1304), .ZN(n1336) );
XOR2_X1 U1078 ( .A(G116), .B(G119), .Z(n1304) );
XOR2_X1 U1079 ( .A(n1117), .B(n1337), .Z(n1335) );
NOR2_X1 U1080 ( .A1(G953), .A2(n1110), .ZN(n1337) );
INV_X1 U1081 ( .A(G224), .ZN(n1110) );
XOR2_X1 U1082 ( .A(n1338), .B(n1159), .Z(n1117) );
XOR2_X1 U1083 ( .A(G101), .B(G110), .Z(n1159) );
XOR2_X1 U1084 ( .A(n1339), .B(n1340), .Z(n1338) );
NOR2_X1 U1085 ( .A1(KEYINPUT44), .A2(n1310), .ZN(n1340) );
XNOR2_X1 U1086 ( .A(G104), .B(G107), .ZN(n1310) );
INV_X1 U1087 ( .A(G122), .ZN(n1339) );
endmodule


