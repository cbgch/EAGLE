//Key = 1011100100111000001100100110010100110100010000011110010101001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;

XNOR2_X1 U735 ( .A(G107), .B(n1006), .ZN(G9) );
NOR2_X1 U736 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U737 ( .A1(n1009), .A2(n1010), .A3(G953), .A4(n1011), .ZN(n1008) );
NOR3_X1 U738 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
NOR2_X1 U739 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U740 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U742 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U743 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U744 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U745 ( .A1(n1027), .A2(n1028), .ZN(n1019) );
NOR2_X1 U746 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U747 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR3_X1 U748 ( .A1(n1028), .A2(n1033), .A3(n1022), .ZN(n1015) );
NOR2_X1 U749 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U750 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1009) );
NAND3_X1 U751 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1037) );
XOR2_X1 U752 ( .A(KEYINPUT13), .B(n1042), .Z(n1039) );
NAND2_X1 U753 ( .A1(n1043), .A2(n1042), .ZN(n1036) );
NOR4_X1 U754 ( .A1(n1012), .A2(n1018), .A3(n1028), .A4(n1022), .ZN(n1042) );
XOR2_X1 U755 ( .A(n1044), .B(KEYINPUT22), .Z(n1043) );
NOR3_X1 U756 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1007) );
AND4_X1 U757 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1011) );
NOR4_X1 U758 ( .A1(n1026), .A2(n1049), .A3(n1022), .A4(n1050), .ZN(n1048) );
XOR2_X1 U759 ( .A(G475), .B(n1051), .Z(n1050) );
NOR2_X1 U760 ( .A1(KEYINPUT51), .A2(n1052), .ZN(n1051) );
INV_X1 U761 ( .A(n1053), .ZN(n1022) );
NOR2_X1 U762 ( .A1(n1054), .A2(n1041), .ZN(n1047) );
INV_X1 U763 ( .A(n1055), .ZN(n1041) );
XOR2_X1 U764 ( .A(n1056), .B(n1057), .Z(n1046) );
NOR2_X1 U765 ( .A1(n1058), .A2(KEYINPUT1), .ZN(n1057) );
XNOR2_X1 U766 ( .A(KEYINPUT47), .B(n1059), .ZN(n1045) );
XOR2_X1 U767 ( .A(n1060), .B(n1061), .Z(G72) );
XOR2_X1 U768 ( .A(n1062), .B(n1063), .Z(n1061) );
NOR2_X1 U769 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XOR2_X1 U770 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U771 ( .A1(G900), .A2(n1068), .ZN(n1064) );
XOR2_X1 U772 ( .A(n1069), .B(KEYINPUT54), .Z(n1068) );
NAND2_X1 U773 ( .A1(n1069), .A2(n1070), .ZN(n1062) );
NAND2_X1 U774 ( .A1(G953), .A2(n1071), .ZN(n1060) );
NAND2_X1 U775 ( .A1(G900), .A2(G227), .ZN(n1071) );
XOR2_X1 U776 ( .A(n1072), .B(n1073), .Z(G69) );
NOR2_X1 U777 ( .A1(n1074), .A2(n1069), .ZN(n1073) );
AND2_X1 U778 ( .A1(G224), .A2(G898), .ZN(n1074) );
NAND2_X1 U779 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
NAND2_X1 U780 ( .A1(n1077), .A2(n1069), .ZN(n1076) );
XOR2_X1 U781 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U782 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
XOR2_X1 U783 ( .A(n1006), .B(KEYINPUT8), .Z(n1080) );
NAND3_X1 U784 ( .A1(n1079), .A2(G898), .A3(G953), .ZN(n1075) );
NOR2_X1 U785 ( .A1(KEYINPUT16), .A2(n1082), .ZN(n1079) );
NOR2_X1 U786 ( .A1(n1083), .A2(n1084), .ZN(G66) );
XOR2_X1 U787 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U788 ( .A1(KEYINPUT11), .A2(n1087), .ZN(n1086) );
NAND2_X1 U789 ( .A1(n1088), .A2(n1089), .ZN(n1085) );
NOR2_X1 U790 ( .A1(n1083), .A2(n1090), .ZN(G63) );
XOR2_X1 U791 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U792 ( .A1(n1088), .A2(G478), .ZN(n1091) );
NOR2_X1 U793 ( .A1(n1083), .A2(n1093), .ZN(G60) );
XOR2_X1 U794 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U795 ( .A1(n1088), .A2(G475), .ZN(n1094) );
XOR2_X1 U796 ( .A(n1096), .B(n1097), .Z(G6) );
NOR2_X1 U797 ( .A1(n1083), .A2(n1098), .ZN(G57) );
XOR2_X1 U798 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U799 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U800 ( .A(n1103), .B(n1104), .Z(n1099) );
NOR2_X1 U801 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U802 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U803 ( .A1(KEYINPUT14), .A2(n1109), .ZN(n1107) );
NOR2_X1 U804 ( .A1(G101), .A2(KEYINPUT36), .ZN(n1109) );
NOR2_X1 U805 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
NOR2_X1 U806 ( .A1(n1112), .A2(KEYINPUT36), .ZN(n1110) );
NOR2_X1 U807 ( .A1(KEYINPUT14), .A2(n1113), .ZN(n1112) );
NAND2_X1 U808 ( .A1(n1088), .A2(G472), .ZN(n1103) );
NOR3_X1 U809 ( .A1(n1083), .A2(n1114), .A3(n1115), .ZN(G54) );
NOR2_X1 U810 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U811 ( .A(n1118), .B(n1119), .Z(n1117) );
AND2_X1 U812 ( .A1(n1120), .A2(KEYINPUT34), .ZN(n1119) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1122), .ZN(n1114) );
XOR2_X1 U814 ( .A(n1118), .B(n1123), .Z(n1122) );
NOR2_X1 U815 ( .A1(n1124), .A2(n1120), .ZN(n1123) );
XNOR2_X1 U816 ( .A(n1125), .B(n1126), .ZN(n1120) );
NAND2_X1 U817 ( .A1(KEYINPUT49), .A2(n1127), .ZN(n1125) );
INV_X1 U818 ( .A(KEYINPUT34), .ZN(n1124) );
XOR2_X1 U819 ( .A(n1128), .B(n1129), .Z(n1118) );
XOR2_X1 U820 ( .A(G140), .B(G110), .Z(n1129) );
XOR2_X1 U821 ( .A(n1130), .B(n1131), .Z(n1128) );
NAND2_X1 U822 ( .A1(n1088), .A2(G469), .ZN(n1130) );
INV_X1 U823 ( .A(n1116), .ZN(n1121) );
NOR3_X1 U824 ( .A1(n1083), .A2(n1132), .A3(n1133), .ZN(G51) );
NOR2_X1 U825 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U826 ( .A(KEYINPUT4), .B(n1136), .Z(n1134) );
NOR2_X1 U827 ( .A1(n1082), .A2(n1137), .ZN(n1132) );
XOR2_X1 U828 ( .A(KEYINPUT15), .B(n1136), .Z(n1137) );
XNOR2_X1 U829 ( .A(n1138), .B(n1139), .ZN(n1136) );
XOR2_X1 U830 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U831 ( .A1(KEYINPUT57), .A2(n1142), .ZN(n1141) );
NAND2_X1 U832 ( .A1(KEYINPUT55), .A2(n1143), .ZN(n1140) );
XNOR2_X1 U833 ( .A(n1144), .B(n1101), .ZN(n1138) );
NAND2_X1 U834 ( .A1(n1088), .A2(n1056), .ZN(n1144) );
NOR2_X1 U835 ( .A1(n1145), .A2(n1038), .ZN(n1088) );
AND3_X1 U836 ( .A1(n1081), .A2(n1006), .A3(n1146), .ZN(n1038) );
INV_X1 U837 ( .A(n1070), .ZN(n1146) );
NAND4_X1 U838 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1070) );
NOR4_X1 U839 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
INV_X1 U840 ( .A(n1155), .ZN(n1154) );
NAND2_X1 U841 ( .A1(n1156), .A2(n1157), .ZN(n1149) );
NAND2_X1 U842 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U843 ( .A1(n1160), .A2(n1030), .ZN(n1159) );
XOR2_X1 U844 ( .A(n1161), .B(KEYINPUT40), .Z(n1158) );
NAND3_X1 U845 ( .A1(n1034), .A2(n1162), .A3(n1163), .ZN(n1147) );
NAND3_X1 U846 ( .A1(n1164), .A2(n1165), .A3(n1034), .ZN(n1006) );
AND4_X1 U847 ( .A1(n1097), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1081) );
AND4_X1 U848 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1168) );
NAND3_X1 U849 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1167) );
XOR2_X1 U850 ( .A(KEYINPUT32), .B(n1053), .Z(n1174) );
NAND3_X1 U851 ( .A1(n1164), .A2(n1165), .A3(n1035), .ZN(n1097) );
NOR2_X1 U852 ( .A1(n1069), .A2(G952), .ZN(n1083) );
XNOR2_X1 U853 ( .A(G146), .B(n1148), .ZN(G48) );
NAND3_X1 U854 ( .A1(n1035), .A2(n1162), .A3(n1163), .ZN(n1148) );
INV_X1 U855 ( .A(n1176), .ZN(n1163) );
XOR2_X1 U856 ( .A(n1177), .B(n1155), .Z(G45) );
NAND3_X1 U857 ( .A1(n1024), .A2(n1178), .A3(n1179), .ZN(n1155) );
NOR3_X1 U858 ( .A1(n1180), .A2(n1181), .A3(n1044), .ZN(n1179) );
XOR2_X1 U859 ( .A(n1182), .B(n1183), .Z(G42) );
NAND3_X1 U860 ( .A1(n1184), .A2(n1030), .A3(n1160), .ZN(n1183) );
XOR2_X1 U861 ( .A(KEYINPUT59), .B(n1156), .Z(n1184) );
XNOR2_X1 U862 ( .A(G137), .B(n1185), .ZN(G39) );
NAND2_X1 U863 ( .A1(KEYINPUT50), .A2(n1153), .ZN(n1185) );
NOR3_X1 U864 ( .A1(n1176), .A2(n1014), .A3(n1018), .ZN(n1153) );
XOR2_X1 U865 ( .A(n1186), .B(n1187), .Z(G36) );
NAND2_X1 U866 ( .A1(KEYINPUT31), .A2(n1152), .ZN(n1187) );
AND4_X1 U867 ( .A1(n1024), .A2(n1156), .A3(n1178), .A4(n1034), .ZN(n1152) );
INV_X1 U868 ( .A(n1014), .ZN(n1156) );
XOR2_X1 U869 ( .A(G131), .B(n1188), .Z(G33) );
NOR2_X1 U870 ( .A1(n1014), .A2(n1161), .ZN(n1188) );
NAND2_X1 U871 ( .A1(n1175), .A2(n1178), .ZN(n1161) );
INV_X1 U872 ( .A(n1189), .ZN(n1175) );
NAND2_X1 U873 ( .A1(n1040), .A2(n1055), .ZN(n1014) );
XNOR2_X1 U874 ( .A(n1190), .B(KEYINPUT46), .ZN(n1040) );
XOR2_X1 U875 ( .A(G128), .B(n1191), .Z(G30) );
NOR3_X1 U876 ( .A1(n1192), .A2(n1193), .A3(n1176), .ZN(n1191) );
NAND3_X1 U877 ( .A1(n1194), .A2(n1195), .A3(n1178), .ZN(n1176) );
AND2_X1 U878 ( .A1(n1030), .A2(n1196), .ZN(n1178) );
XOR2_X1 U879 ( .A(KEYINPUT62), .B(n1162), .Z(n1192) );
XOR2_X1 U880 ( .A(n1111), .B(n1166), .Z(G3) );
NAND3_X1 U881 ( .A1(n1024), .A2(n1165), .A3(n1197), .ZN(n1166) );
XOR2_X1 U882 ( .A(G125), .B(n1151), .Z(G27) );
AND3_X1 U883 ( .A1(n1053), .A2(n1162), .A3(n1160), .ZN(n1151) );
AND4_X1 U884 ( .A1(n1198), .A2(n1035), .A3(n1196), .A4(n1195), .ZN(n1160) );
NAND2_X1 U885 ( .A1(n1012), .A2(n1199), .ZN(n1196) );
NAND4_X1 U886 ( .A1(G953), .A2(G902), .A3(n1200), .A4(n1201), .ZN(n1199) );
INV_X1 U887 ( .A(G900), .ZN(n1201) );
XNOR2_X1 U888 ( .A(G122), .B(n1172), .ZN(G24) );
NAND4_X1 U889 ( .A1(n1202), .A2(n1203), .A3(n1164), .A4(n1204), .ZN(n1172) );
INV_X1 U890 ( .A(n1028), .ZN(n1164) );
NAND2_X1 U891 ( .A1(n1025), .A2(n1198), .ZN(n1028) );
XOR2_X1 U892 ( .A(n1205), .B(n1171), .Z(G21) );
NAND4_X1 U893 ( .A1(n1203), .A2(n1197), .A3(n1194), .A4(n1195), .ZN(n1171) );
XOR2_X1 U894 ( .A(n1206), .B(n1207), .Z(G18) );
XOR2_X1 U895 ( .A(KEYINPUT28), .B(G116), .Z(n1207) );
NAND2_X1 U896 ( .A1(KEYINPUT53), .A2(n1170), .ZN(n1206) );
NAND3_X1 U897 ( .A1(n1024), .A2(n1034), .A3(n1203), .ZN(n1170) );
INV_X1 U898 ( .A(n1208), .ZN(n1203) );
INV_X1 U899 ( .A(n1193), .ZN(n1034) );
NAND2_X1 U900 ( .A1(n1180), .A2(n1204), .ZN(n1193) );
XOR2_X1 U901 ( .A(n1209), .B(n1210), .Z(G15) );
NOR2_X1 U902 ( .A1(n1189), .A2(n1208), .ZN(n1210) );
NAND2_X1 U903 ( .A1(n1173), .A2(n1053), .ZN(n1208) );
NAND2_X1 U904 ( .A1(n1024), .A2(n1035), .ZN(n1189) );
NOR2_X1 U905 ( .A1(n1204), .A2(n1180), .ZN(n1035) );
INV_X1 U906 ( .A(n1181), .ZN(n1204) );
AND2_X1 U907 ( .A1(n1025), .A2(n1194), .ZN(n1024) );
XOR2_X1 U908 ( .A(n1026), .B(KEYINPUT21), .Z(n1194) );
INV_X1 U909 ( .A(n1198), .ZN(n1026) );
INV_X1 U910 ( .A(n1195), .ZN(n1025) );
NOR2_X1 U911 ( .A1(KEYINPUT20), .A2(n1211), .ZN(n1209) );
XOR2_X1 U912 ( .A(n1212), .B(n1169), .Z(G12) );
NAND4_X1 U913 ( .A1(n1197), .A2(n1165), .A3(n1198), .A4(n1195), .ZN(n1169) );
NAND2_X1 U914 ( .A1(n1213), .A2(n1059), .ZN(n1195) );
NAND2_X1 U915 ( .A1(n1089), .A2(n1214), .ZN(n1059) );
OR2_X1 U916 ( .A1(n1087), .A2(G902), .ZN(n1214) );
XNOR2_X1 U917 ( .A(n1054), .B(KEYINPUT56), .ZN(n1213) );
NOR3_X1 U918 ( .A1(n1089), .A2(G902), .A3(n1087), .ZN(n1054) );
XOR2_X1 U919 ( .A(n1215), .B(n1216), .Z(n1087) );
XOR2_X1 U920 ( .A(G110), .B(n1217), .Z(n1216) );
NOR2_X1 U921 ( .A1(KEYINPUT52), .A2(n1218), .ZN(n1217) );
XOR2_X1 U922 ( .A(n1219), .B(n1220), .Z(n1218) );
NAND3_X1 U923 ( .A1(n1221), .A2(n1069), .A3(G221), .ZN(n1219) );
XOR2_X1 U924 ( .A(n1222), .B(n1223), .Z(n1215) );
NOR2_X1 U925 ( .A1(KEYINPUT33), .A2(n1224), .ZN(n1223) );
XOR2_X1 U926 ( .A(n1066), .B(n1225), .Z(n1224) );
NOR2_X1 U927 ( .A1(G146), .A2(KEYINPUT9), .ZN(n1225) );
INV_X1 U928 ( .A(n1226), .ZN(n1066) );
NAND3_X1 U929 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1222) );
NAND2_X1 U930 ( .A1(n1230), .A2(n1205), .ZN(n1229) );
INV_X1 U931 ( .A(G119), .ZN(n1205) );
NAND3_X1 U932 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1230) );
NAND2_X1 U933 ( .A1(KEYINPUT43), .A2(n1234), .ZN(n1233) );
OR2_X1 U934 ( .A1(G128), .A2(KEYINPUT35), .ZN(n1232) );
NAND2_X1 U935 ( .A1(KEYINPUT35), .A2(n1235), .ZN(n1231) );
NAND2_X1 U936 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U937 ( .A1(KEYINPUT58), .A2(n1238), .ZN(n1237) );
NAND4_X1 U938 ( .A1(n1236), .A2(n1234), .A3(G119), .A4(n1238), .ZN(n1228) );
INV_X1 U939 ( .A(KEYINPUT43), .ZN(n1238) );
INV_X1 U940 ( .A(KEYINPUT58), .ZN(n1234) );
NAND2_X1 U941 ( .A1(KEYINPUT43), .A2(n1239), .ZN(n1227) );
NAND2_X1 U942 ( .A1(n1236), .A2(n1240), .ZN(n1239) );
NAND2_X1 U943 ( .A1(KEYINPUT58), .A2(G119), .ZN(n1240) );
INV_X1 U944 ( .A(G128), .ZN(n1236) );
AND2_X1 U945 ( .A1(G217), .A2(n1241), .ZN(n1089) );
XOR2_X1 U946 ( .A(n1242), .B(G472), .Z(n1198) );
NAND2_X1 U947 ( .A1(n1243), .A2(n1145), .ZN(n1242) );
XOR2_X1 U948 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U949 ( .A(n1113), .B(n1102), .Z(n1245) );
XOR2_X1 U950 ( .A(n1246), .B(n1116), .Z(n1102) );
INV_X1 U951 ( .A(n1108), .ZN(n1113) );
NAND3_X1 U952 ( .A1(n1247), .A2(n1069), .A3(G210), .ZN(n1108) );
XOR2_X1 U953 ( .A(n1248), .B(n1249), .Z(n1244) );
NOR2_X1 U954 ( .A1(KEYINPUT30), .A2(n1250), .ZN(n1249) );
XOR2_X1 U955 ( .A(n1101), .B(KEYINPUT42), .Z(n1250) );
XOR2_X1 U956 ( .A(n1111), .B(KEYINPUT7), .Z(n1248) );
AND2_X1 U957 ( .A1(n1173), .A2(n1030), .ZN(n1165) );
NAND2_X1 U958 ( .A1(n1251), .A2(n1252), .ZN(n1030) );
NAND3_X1 U959 ( .A1(n1031), .A2(n1032), .A3(n1253), .ZN(n1252) );
INV_X1 U960 ( .A(KEYINPUT61), .ZN(n1253) );
NAND2_X1 U961 ( .A1(KEYINPUT61), .A2(n1053), .ZN(n1251) );
NOR2_X1 U962 ( .A1(n1031), .A2(n1254), .ZN(n1053) );
INV_X1 U963 ( .A(n1032), .ZN(n1254) );
NAND2_X1 U964 ( .A1(G221), .A2(n1241), .ZN(n1032) );
NAND2_X1 U965 ( .A1(G234), .A2(n1145), .ZN(n1241) );
XNOR2_X1 U966 ( .A(n1255), .B(G469), .ZN(n1031) );
NAND3_X1 U967 ( .A1(n1256), .A2(n1257), .A3(n1145), .ZN(n1255) );
NAND2_X1 U968 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
INV_X1 U969 ( .A(KEYINPUT6), .ZN(n1259) );
XNOR2_X1 U970 ( .A(n1260), .B(n1261), .ZN(n1258) );
NAND2_X1 U971 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
NAND4_X1 U972 ( .A1(n1263), .A2(n1262), .A3(n1261), .A4(KEYINPUT6), .ZN(n1256) );
XOR2_X1 U973 ( .A(n1264), .B(n1067), .Z(n1261) );
XNOR2_X1 U974 ( .A(n1126), .B(n1116), .ZN(n1067) );
XOR2_X1 U975 ( .A(n1265), .B(n1220), .Z(n1116) );
XOR2_X1 U976 ( .A(G137), .B(KEYINPUT24), .Z(n1220) );
XOR2_X1 U977 ( .A(G131), .B(n1186), .Z(n1265) );
INV_X1 U978 ( .A(G134), .ZN(n1186) );
XNOR2_X1 U979 ( .A(n1266), .B(n1267), .ZN(n1126) );
XOR2_X1 U980 ( .A(n1177), .B(G146), .Z(n1266) );
XNOR2_X1 U981 ( .A(n1127), .B(KEYINPUT19), .ZN(n1264) );
XNOR2_X1 U982 ( .A(n1268), .B(n1269), .ZN(n1127) );
NOR2_X1 U983 ( .A1(G107), .A2(KEYINPUT38), .ZN(n1269) );
XOR2_X1 U984 ( .A(n1096), .B(G101), .Z(n1268) );
NAND2_X1 U985 ( .A1(n1270), .A2(n1271), .ZN(n1262) );
XOR2_X1 U986 ( .A(n1272), .B(G140), .Z(n1271) );
XNOR2_X1 U987 ( .A(KEYINPUT17), .B(n1131), .ZN(n1270) );
NAND2_X1 U988 ( .A1(n1273), .A2(n1274), .ZN(n1263) );
XOR2_X1 U989 ( .A(n1182), .B(n1272), .Z(n1274) );
NAND2_X1 U990 ( .A1(KEYINPUT60), .A2(n1212), .ZN(n1272) );
INV_X1 U991 ( .A(G140), .ZN(n1182) );
XOR2_X1 U992 ( .A(KEYINPUT17), .B(n1131), .Z(n1273) );
AND2_X1 U993 ( .A1(G227), .A2(n1069), .ZN(n1131) );
AND2_X1 U994 ( .A1(n1162), .A2(n1275), .ZN(n1173) );
NAND2_X1 U995 ( .A1(n1012), .A2(n1276), .ZN(n1275) );
NAND4_X1 U996 ( .A1(G953), .A2(G902), .A3(n1200), .A4(n1277), .ZN(n1276) );
INV_X1 U997 ( .A(G898), .ZN(n1277) );
NAND3_X1 U998 ( .A1(n1200), .A2(n1069), .A3(G952), .ZN(n1012) );
NAND2_X1 U999 ( .A1(G237), .A2(G234), .ZN(n1200) );
INV_X1 U1000 ( .A(n1044), .ZN(n1162) );
NAND2_X1 U1001 ( .A1(n1190), .A2(n1055), .ZN(n1044) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1278), .ZN(n1055) );
XOR2_X1 U1003 ( .A(n1279), .B(n1056), .Z(n1190) );
AND2_X1 U1004 ( .A1(G210), .A2(n1278), .ZN(n1056) );
NAND2_X1 U1005 ( .A1(n1247), .A2(n1145), .ZN(n1278) );
XNOR2_X1 U1006 ( .A(n1058), .B(KEYINPUT0), .ZN(n1279) );
AND2_X1 U1007 ( .A1(n1280), .A2(n1145), .ZN(n1058) );
XOR2_X1 U1008 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U1009 ( .A(n1082), .B(n1142), .Z(n1282) );
NAND2_X1 U1010 ( .A1(G224), .A2(n1069), .ZN(n1142) );
INV_X1 U1011 ( .A(n1135), .ZN(n1082) );
XOR2_X1 U1012 ( .A(n1283), .B(n1284), .Z(n1135) );
XOR2_X1 U1013 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U1014 ( .A(G110), .B(G107), .Z(n1286) );
XOR2_X1 U1015 ( .A(KEYINPUT3), .B(G122), .Z(n1285) );
XOR2_X1 U1016 ( .A(n1246), .B(n1287), .Z(n1283) );
XOR2_X1 U1017 ( .A(n1096), .B(n1288), .Z(n1287) );
NAND2_X1 U1018 ( .A1(KEYINPUT29), .A2(n1111), .ZN(n1288) );
INV_X1 U1019 ( .A(G101), .ZN(n1111) );
XOR2_X1 U1020 ( .A(n1211), .B(n1289), .Z(n1246) );
XOR2_X1 U1021 ( .A(G119), .B(G116), .Z(n1289) );
INV_X1 U1022 ( .A(G113), .ZN(n1211) );
XOR2_X1 U1023 ( .A(n1143), .B(n1290), .Z(n1281) );
NOR2_X1 U1024 ( .A1(KEYINPUT45), .A2(n1101), .ZN(n1290) );
XOR2_X1 U1025 ( .A(n1291), .B(n1267), .Z(n1101) );
XOR2_X1 U1026 ( .A(G128), .B(KEYINPUT18), .Z(n1267) );
NAND3_X1 U1027 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1291) );
OR2_X1 U1028 ( .A1(n1295), .A2(G146), .ZN(n1294) );
NAND3_X1 U1029 ( .A1(G146), .A2(n1295), .A3(n1177), .ZN(n1293) );
NAND2_X1 U1030 ( .A1(G143), .A2(n1296), .ZN(n1292) );
NAND2_X1 U1031 ( .A1(n1297), .A2(n1295), .ZN(n1296) );
INV_X1 U1032 ( .A(KEYINPUT44), .ZN(n1295) );
XNOR2_X1 U1033 ( .A(G146), .B(KEYINPUT41), .ZN(n1297) );
INV_X1 U1034 ( .A(n1018), .ZN(n1197) );
NAND2_X1 U1035 ( .A1(n1181), .A2(n1180), .ZN(n1018) );
INV_X1 U1036 ( .A(n1202), .ZN(n1180) );
XNOR2_X1 U1037 ( .A(G475), .B(n1298), .ZN(n1202) );
NOR2_X1 U1038 ( .A1(n1299), .A2(KEYINPUT39), .ZN(n1298) );
INV_X1 U1039 ( .A(n1052), .ZN(n1299) );
NAND2_X1 U1040 ( .A1(n1095), .A2(n1145), .ZN(n1052) );
XOR2_X1 U1041 ( .A(n1300), .B(n1301), .Z(n1095) );
XOR2_X1 U1042 ( .A(G146), .B(n1302), .Z(n1301) );
NOR2_X1 U1043 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XOR2_X1 U1044 ( .A(n1305), .B(KEYINPUT25), .Z(n1304) );
NAND2_X1 U1045 ( .A1(n1306), .A2(n1096), .ZN(n1305) );
INV_X1 U1046 ( .A(G104), .ZN(n1096) );
NOR2_X1 U1047 ( .A1(n1306), .A2(n1307), .ZN(n1303) );
XOR2_X1 U1048 ( .A(KEYINPUT37), .B(G104), .Z(n1307) );
XOR2_X1 U1049 ( .A(G113), .B(n1308), .Z(n1306) );
XOR2_X1 U1050 ( .A(KEYINPUT12), .B(G122), .Z(n1308) );
XOR2_X1 U1051 ( .A(n1309), .B(n1226), .Z(n1300) );
XNOR2_X1 U1052 ( .A(n1143), .B(G140), .ZN(n1226) );
INV_X1 U1053 ( .A(G125), .ZN(n1143) );
NAND2_X1 U1054 ( .A1(n1310), .A2(KEYINPUT63), .ZN(n1309) );
XOR2_X1 U1055 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U1056 ( .A(G131), .B(n1313), .Z(n1312) );
NOR2_X1 U1057 ( .A1(KEYINPUT23), .A2(n1177), .ZN(n1313) );
NAND3_X1 U1058 ( .A1(n1247), .A2(n1069), .A3(n1314), .ZN(n1311) );
XNOR2_X1 U1059 ( .A(G214), .B(KEYINPUT26), .ZN(n1314) );
INV_X1 U1060 ( .A(G237), .ZN(n1247) );
XNOR2_X1 U1061 ( .A(n1049), .B(KEYINPUT5), .ZN(n1181) );
XNOR2_X1 U1062 ( .A(n1315), .B(G478), .ZN(n1049) );
NAND2_X1 U1063 ( .A1(n1092), .A2(n1145), .ZN(n1315) );
INV_X1 U1064 ( .A(G902), .ZN(n1145) );
XNOR2_X1 U1065 ( .A(n1316), .B(n1317), .ZN(n1092) );
AND3_X1 U1066 ( .A1(G217), .A2(n1069), .A3(n1221), .ZN(n1317) );
XNOR2_X1 U1067 ( .A(G234), .B(KEYINPUT48), .ZN(n1221) );
INV_X1 U1068 ( .A(G953), .ZN(n1069) );
NAND2_X1 U1069 ( .A1(n1318), .A2(KEYINPUT2), .ZN(n1316) );
XOR2_X1 U1070 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1071 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1072 ( .A(G128), .B(G122), .Z(n1322) );
XOR2_X1 U1073 ( .A(KEYINPUT27), .B(G134), .Z(n1321) );
XOR2_X1 U1074 ( .A(n1323), .B(n1324), .Z(n1319) );
XOR2_X1 U1075 ( .A(G116), .B(G107), .Z(n1324) );
NAND2_X1 U1076 ( .A1(KEYINPUT10), .A2(n1177), .ZN(n1323) );
INV_X1 U1077 ( .A(G143), .ZN(n1177) );
INV_X1 U1078 ( .A(G110), .ZN(n1212) );
endmodule


