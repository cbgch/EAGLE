//Key = 1111101110000111110100011001010010001100000001110100111110011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;

XNOR2_X1 U721 ( .A(G107), .B(n981), .ZN(G9) );
NOR2_X1 U722 ( .A1(n982), .A2(n983), .ZN(G75) );
NOR4_X1 U723 ( .A1(G953), .A2(n984), .A3(n985), .A4(n986), .ZN(n983) );
NOR2_X1 U724 ( .A1(n987), .A2(n988), .ZN(n985) );
NOR2_X1 U725 ( .A1(n989), .A2(n990), .ZN(n987) );
NOR2_X1 U726 ( .A1(n991), .A2(n992), .ZN(n990) );
NOR2_X1 U727 ( .A1(n993), .A2(n994), .ZN(n991) );
NOR2_X1 U728 ( .A1(n995), .A2(n996), .ZN(n994) );
NOR2_X1 U729 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR2_X1 U730 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR2_X1 U731 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U732 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U733 ( .A1(n1005), .A2(n1006), .ZN(n997) );
NOR2_X1 U734 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR2_X1 U735 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR3_X1 U736 ( .A1(n1006), .A2(n1011), .A3(n1000), .ZN(n993) );
NOR2_X1 U737 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR3_X1 U738 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1012) );
INV_X1 U739 ( .A(n1017), .ZN(n1016) );
NOR4_X1 U740 ( .A1(n1018), .A2(n1000), .A3(n996), .A4(n1006), .ZN(n989) );
NOR2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR3_X1 U742 ( .A1(n984), .A2(G953), .A3(G952), .ZN(n982) );
AND4_X1 U743 ( .A1(n1009), .A2(n1004), .A3(n1021), .A4(n1022), .ZN(n984) );
NOR4_X1 U744 ( .A1(n1023), .A2(n1024), .A3(n992), .A4(n1025), .ZN(n1022) );
XOR2_X1 U745 ( .A(n1026), .B(n1027), .Z(n1025) );
XNOR2_X1 U746 ( .A(KEYINPUT43), .B(n1028), .ZN(n1027) );
NOR2_X1 U747 ( .A1(KEYINPUT33), .A2(n1029), .ZN(n1028) );
INV_X1 U748 ( .A(n1030), .ZN(n992) );
NOR2_X1 U749 ( .A1(n1031), .A2(n1032), .ZN(n1024) );
NOR2_X1 U750 ( .A1(G472), .A2(n1033), .ZN(n1023) );
XOR2_X1 U751 ( .A(n1032), .B(KEYINPUT17), .Z(n1033) );
XOR2_X1 U752 ( .A(n1034), .B(KEYINPUT4), .Z(n1032) );
INV_X1 U753 ( .A(n1035), .ZN(n1009) );
XOR2_X1 U754 ( .A(n1036), .B(n1037), .Z(G72) );
NAND2_X1 U755 ( .A1(G953), .A2(n1038), .ZN(n1037) );
NAND2_X1 U756 ( .A1(G900), .A2(G227), .ZN(n1038) );
NAND2_X1 U757 ( .A1(KEYINPUT19), .A2(n1039), .ZN(n1036) );
XOR2_X1 U758 ( .A(n1040), .B(n1041), .Z(n1039) );
NOR2_X1 U759 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n1044), .ZN(n1043) );
NOR2_X1 U761 ( .A1(n1045), .A2(n1046), .ZN(n1040) );
XOR2_X1 U762 ( .A(n1047), .B(n1048), .Z(n1046) );
XOR2_X1 U763 ( .A(G140), .B(n1049), .Z(n1048) );
NOR2_X1 U764 ( .A1(G125), .A2(KEYINPUT18), .ZN(n1049) );
XOR2_X1 U765 ( .A(n1050), .B(n1051), .Z(n1047) );
NAND2_X1 U766 ( .A1(KEYINPUT16), .A2(n1052), .ZN(n1050) );
XOR2_X1 U767 ( .A(n1053), .B(n1054), .Z(G69) );
XOR2_X1 U768 ( .A(n1055), .B(n1056), .Z(n1054) );
NOR2_X1 U769 ( .A1(n1057), .A2(n1044), .ZN(n1056) );
NOR2_X1 U770 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U771 ( .A1(n1060), .A2(n1061), .ZN(n1055) );
XOR2_X1 U772 ( .A(n1062), .B(n1063), .Z(n1061) );
NAND3_X1 U773 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1062) );
OR2_X1 U774 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U775 ( .A1(KEYINPUT38), .A2(n1069), .ZN(n1065) );
NAND2_X1 U776 ( .A1(n1070), .A2(n1068), .ZN(n1069) );
XNOR2_X1 U777 ( .A(KEYINPUT27), .B(n1067), .ZN(n1070) );
NAND2_X1 U778 ( .A1(n1071), .A2(n1072), .ZN(n1064) );
INV_X1 U779 ( .A(KEYINPUT38), .ZN(n1072) );
NAND2_X1 U780 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
OR2_X1 U781 ( .A1(n1067), .A2(KEYINPUT27), .ZN(n1074) );
NAND3_X1 U782 ( .A1(n1067), .A2(n1068), .A3(KEYINPUT27), .ZN(n1073) );
XOR2_X1 U783 ( .A(n1075), .B(KEYINPUT35), .Z(n1060) );
NAND2_X1 U784 ( .A1(n1076), .A2(n1059), .ZN(n1075) );
NAND2_X1 U785 ( .A1(n1044), .A2(n1077), .ZN(n1053) );
NOR2_X1 U786 ( .A1(n1078), .A2(n1079), .ZN(G66) );
XNOR2_X1 U787 ( .A(n1080), .B(n1081), .ZN(n1079) );
NOR2_X1 U788 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U789 ( .A1(n1078), .A2(n1084), .ZN(G63) );
XOR2_X1 U790 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND3_X1 U791 ( .A1(n1087), .A2(G478), .A3(KEYINPUT45), .ZN(n1085) );
NOR2_X1 U792 ( .A1(n1078), .A2(n1088), .ZN(G60) );
XOR2_X1 U793 ( .A(n1089), .B(n1090), .Z(n1088) );
NAND3_X1 U794 ( .A1(G475), .A2(G902), .A3(n1091), .ZN(n1089) );
XOR2_X1 U795 ( .A(n986), .B(KEYINPUT58), .Z(n1091) );
XNOR2_X1 U796 ( .A(G104), .B(n1092), .ZN(G6) );
NOR2_X1 U797 ( .A1(n1078), .A2(n1093), .ZN(G57) );
XOR2_X1 U798 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U799 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U800 ( .A1(KEYINPUT52), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U801 ( .A(n1099), .B(n1100), .ZN(n1094) );
NOR3_X1 U802 ( .A1(n1083), .A2(KEYINPUT41), .A3(n1031), .ZN(n1100) );
NAND2_X1 U803 ( .A1(KEYINPUT56), .A2(n1101), .ZN(n1099) );
NOR2_X1 U804 ( .A1(n1078), .A2(n1102), .ZN(G54) );
XOR2_X1 U805 ( .A(n1103), .B(n1104), .Z(n1102) );
AND2_X1 U806 ( .A1(G469), .A2(n1087), .ZN(n1104) );
INV_X1 U807 ( .A(n1083), .ZN(n1087) );
NAND2_X1 U808 ( .A1(n1105), .A2(KEYINPUT13), .ZN(n1103) );
XOR2_X1 U809 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U810 ( .A(n1051), .B(n1108), .Z(n1107) );
XNOR2_X1 U811 ( .A(n1109), .B(n1110), .ZN(n1108) );
NOR2_X1 U812 ( .A1(KEYINPUT34), .A2(n1111), .ZN(n1110) );
XOR2_X1 U813 ( .A(n1112), .B(n1113), .Z(n1106) );
NOR2_X1 U814 ( .A1(n1078), .A2(n1114), .ZN(G51) );
XOR2_X1 U815 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U816 ( .A1(n1029), .A2(n1083), .ZN(n1116) );
NAND2_X1 U817 ( .A1(G902), .A2(n986), .ZN(n1083) );
NAND2_X1 U818 ( .A1(n1042), .A2(n1117), .ZN(n986) );
INV_X1 U819 ( .A(n1077), .ZN(n1117) );
NAND4_X1 U820 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1077) );
AND4_X1 U821 ( .A1(n1092), .A2(n981), .A3(n1122), .A4(n1123), .ZN(n1121) );
NAND3_X1 U822 ( .A1(n1019), .A2(n1124), .A3(n1125), .ZN(n981) );
NAND3_X1 U823 ( .A1(n1125), .A2(n1124), .A3(n1020), .ZN(n1092) );
NOR2_X1 U824 ( .A1(n1126), .A2(n1127), .ZN(n1120) );
NOR2_X1 U825 ( .A1(n1000), .A2(n1128), .ZN(n1127) );
AND2_X1 U826 ( .A1(n1129), .A2(n1130), .ZN(n1042) );
NOR4_X1 U827 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1130) );
AND3_X1 U828 ( .A1(n1135), .A2(n1019), .A3(n1136), .ZN(n1134) );
INV_X1 U829 ( .A(n1137), .ZN(n1132) );
INV_X1 U830 ( .A(n1138), .ZN(n1131) );
AND4_X1 U831 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1129) );
NOR2_X1 U832 ( .A1(n1143), .A2(n1144), .ZN(n1115) );
XOR2_X1 U833 ( .A(KEYINPUT22), .B(n1145), .Z(n1144) );
AND2_X1 U834 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U835 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
XOR2_X1 U836 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U837 ( .A(G125), .B(n1150), .ZN(n1148) );
NOR2_X1 U838 ( .A1(n1044), .A2(G952), .ZN(n1078) );
NAND2_X1 U839 ( .A1(n1151), .A2(n1152), .ZN(G48) );
NAND2_X1 U840 ( .A1(G146), .A2(n1142), .ZN(n1152) );
XOR2_X1 U841 ( .A(KEYINPUT6), .B(n1153), .Z(n1151) );
NOR2_X1 U842 ( .A1(G146), .A2(n1142), .ZN(n1153) );
NAND3_X1 U843 ( .A1(n1002), .A2(n1020), .A3(n1154), .ZN(n1142) );
XNOR2_X1 U844 ( .A(G143), .B(n1141), .ZN(G45) );
NAND4_X1 U845 ( .A1(n1002), .A2(n1135), .A3(n1155), .A4(n1156), .ZN(n1141) );
XOR2_X1 U846 ( .A(G140), .B(n1133), .Z(G42) );
AND3_X1 U847 ( .A1(n1157), .A2(n1013), .A3(n1136), .ZN(n1133) );
XNOR2_X1 U848 ( .A(G137), .B(n1140), .ZN(G39) );
NAND3_X1 U849 ( .A1(n1154), .A2(n1030), .A3(n1136), .ZN(n1140) );
XNOR2_X1 U850 ( .A(G134), .B(n1158), .ZN(G36) );
NAND4_X1 U851 ( .A1(n1159), .A2(n1160), .A3(n1019), .A4(n1161), .ZN(n1158) );
AND2_X1 U852 ( .A1(n1136), .A2(n1008), .ZN(n1161) );
XNOR2_X1 U853 ( .A(KEYINPUT12), .B(n1162), .ZN(n1159) );
XOR2_X1 U854 ( .A(n1139), .B(n1163), .Z(G33) );
NOR2_X1 U855 ( .A1(G131), .A2(KEYINPUT28), .ZN(n1163) );
NAND3_X1 U856 ( .A1(n1136), .A2(n1020), .A3(n1135), .ZN(n1139) );
AND3_X1 U857 ( .A1(n1013), .A2(n1160), .A3(n1008), .ZN(n1135) );
INV_X1 U858 ( .A(n1006), .ZN(n1136) );
NAND2_X1 U859 ( .A1(n1164), .A2(n1004), .ZN(n1006) );
INV_X1 U860 ( .A(n1003), .ZN(n1164) );
XNOR2_X1 U861 ( .A(G128), .B(n1137), .ZN(G30) );
NAND3_X1 U862 ( .A1(n1002), .A2(n1019), .A3(n1154), .ZN(n1137) );
AND4_X1 U863 ( .A1(n1013), .A2(n1035), .A3(n1010), .A4(n1160), .ZN(n1154) );
INV_X1 U864 ( .A(n1162), .ZN(n1013) );
XOR2_X1 U865 ( .A(n1126), .B(n1165), .Z(G3) );
NOR2_X1 U866 ( .A1(KEYINPUT9), .A2(n1166), .ZN(n1165) );
AND3_X1 U867 ( .A1(n1030), .A2(n1125), .A3(n1008), .ZN(n1126) );
XNOR2_X1 U868 ( .A(G125), .B(n1138), .ZN(G27) );
NAND3_X1 U869 ( .A1(n1002), .A2(n1021), .A3(n1157), .ZN(n1138) );
AND4_X1 U870 ( .A1(n1167), .A2(n1020), .A3(n1035), .A4(n1160), .ZN(n1157) );
NAND2_X1 U871 ( .A1(n988), .A2(n1168), .ZN(n1160) );
NAND3_X1 U872 ( .A1(G902), .A2(n1169), .A3(n1045), .ZN(n1168) );
NOR2_X1 U873 ( .A1(n1170), .A2(G900), .ZN(n1045) );
XNOR2_X1 U874 ( .A(n1171), .B(n1172), .ZN(G24) );
NOR2_X1 U875 ( .A1(n1128), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U876 ( .A(KEYINPUT36), .B(n1000), .ZN(n1173) );
INV_X1 U877 ( .A(n1124), .ZN(n1000) );
NOR2_X1 U878 ( .A1(n1010), .A2(n1035), .ZN(n1124) );
NAND3_X1 U879 ( .A1(n1155), .A2(n1156), .A3(n1174), .ZN(n1128) );
XNOR2_X1 U880 ( .A(G119), .B(n1118), .ZN(G21) );
NAND4_X1 U881 ( .A1(n1174), .A2(n1030), .A3(n1035), .A4(n1010), .ZN(n1118) );
XNOR2_X1 U882 ( .A(G116), .B(n1119), .ZN(G18) );
NAND3_X1 U883 ( .A1(n1008), .A2(n1019), .A3(n1174), .ZN(n1119) );
AND3_X1 U884 ( .A1(n1021), .A2(n1175), .A3(n1002), .ZN(n1174) );
XOR2_X1 U885 ( .A(n1176), .B(KEYINPUT2), .Z(n1002) );
NOR2_X1 U886 ( .A1(n1156), .A2(n1177), .ZN(n1019) );
XOR2_X1 U887 ( .A(G113), .B(n1178), .Z(G15) );
NOR2_X1 U888 ( .A1(KEYINPUT26), .A2(n1123), .ZN(n1178) );
NAND4_X1 U889 ( .A1(n1008), .A2(n1020), .A3(n1179), .A4(n1021), .ZN(n1123) );
INV_X1 U890 ( .A(n996), .ZN(n1021) );
NAND3_X1 U891 ( .A1(n1014), .A2(n1180), .A3(n1017), .ZN(n996) );
NOR2_X1 U892 ( .A1(n1181), .A2(n1176), .ZN(n1179) );
AND2_X1 U893 ( .A1(n1177), .A2(n1156), .ZN(n1020) );
INV_X1 U894 ( .A(n1155), .ZN(n1177) );
NOR2_X1 U895 ( .A1(n1035), .A2(n1167), .ZN(n1008) );
XOR2_X1 U896 ( .A(G110), .B(n1182), .Z(G12) );
NOR2_X1 U897 ( .A1(KEYINPUT11), .A2(n1122), .ZN(n1182) );
NAND4_X1 U898 ( .A1(n1030), .A2(n1125), .A3(n1167), .A4(n1035), .ZN(n1122) );
XOR2_X1 U899 ( .A(n1183), .B(n1082), .Z(n1035) );
NAND2_X1 U900 ( .A1(G217), .A2(n1184), .ZN(n1082) );
NAND2_X1 U901 ( .A1(n1080), .A2(n1185), .ZN(n1183) );
XNOR2_X1 U902 ( .A(n1186), .B(n1187), .ZN(n1080) );
XOR2_X1 U903 ( .A(n1188), .B(n1189), .Z(n1187) );
XNOR2_X1 U904 ( .A(n1190), .B(G119), .ZN(n1189) );
INV_X1 U905 ( .A(G128), .ZN(n1190) );
XOR2_X1 U906 ( .A(KEYINPUT57), .B(G137), .Z(n1188) );
XOR2_X1 U907 ( .A(n1191), .B(n1192), .Z(n1186) );
AND3_X1 U908 ( .A1(G221), .A2(n1044), .A3(G234), .ZN(n1192) );
XNOR2_X1 U909 ( .A(G110), .B(n1193), .ZN(n1191) );
NOR2_X1 U910 ( .A1(KEYINPUT31), .A2(n1194), .ZN(n1193) );
XOR2_X1 U911 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U912 ( .A(G140), .B(n1197), .ZN(n1196) );
NOR2_X1 U913 ( .A1(KEYINPUT30), .A2(n1198), .ZN(n1195) );
XNOR2_X1 U914 ( .A(n1199), .B(KEYINPUT1), .ZN(n1198) );
INV_X1 U915 ( .A(n1010), .ZN(n1167) );
XNOR2_X1 U916 ( .A(n1034), .B(n1200), .ZN(n1010) );
XNOR2_X1 U917 ( .A(KEYINPUT5), .B(n1031), .ZN(n1200) );
INV_X1 U918 ( .A(G472), .ZN(n1031) );
NAND2_X1 U919 ( .A1(n1201), .A2(n1185), .ZN(n1034) );
XOR2_X1 U920 ( .A(n1097), .B(n1202), .Z(n1201) );
XOR2_X1 U921 ( .A(n1203), .B(n1101), .Z(n1202) );
XOR2_X1 U922 ( .A(n1204), .B(G113), .Z(n1101) );
NAND2_X1 U923 ( .A1(n1205), .A2(KEYINPUT8), .ZN(n1203) );
XOR2_X1 U924 ( .A(n1098), .B(KEYINPUT29), .Z(n1205) );
XNOR2_X1 U925 ( .A(n1206), .B(n1166), .ZN(n1098) );
NAND3_X1 U926 ( .A1(n1207), .A2(n1044), .A3(G210), .ZN(n1206) );
XOR2_X1 U927 ( .A(n1111), .B(n1149), .Z(n1097) );
NOR3_X1 U928 ( .A1(n1176), .A2(n1181), .A3(n1162), .ZN(n1125) );
NAND2_X1 U929 ( .A1(n1014), .A2(n1208), .ZN(n1162) );
NAND2_X1 U930 ( .A1(n1017), .A2(n1180), .ZN(n1208) );
INV_X1 U931 ( .A(n1015), .ZN(n1180) );
NOR3_X1 U932 ( .A1(n1209), .A2(G902), .A3(n1210), .ZN(n1015) );
NAND2_X1 U933 ( .A1(n1210), .A2(n1211), .ZN(n1017) );
OR2_X1 U934 ( .A1(n1209), .A2(G902), .ZN(n1211) );
XOR2_X1 U935 ( .A(n1111), .B(n1212), .Z(n1209) );
XOR2_X1 U936 ( .A(n1213), .B(n1214), .Z(n1212) );
NAND3_X1 U937 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
OR2_X1 U938 ( .A1(n1051), .A2(KEYINPUT37), .ZN(n1217) );
OR3_X1 U939 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1216) );
INV_X1 U940 ( .A(KEYINPUT37), .ZN(n1218) );
NAND2_X1 U941 ( .A1(n1220), .A2(n1219), .ZN(n1215) );
NAND2_X1 U942 ( .A1(KEYINPUT14), .A2(n1051), .ZN(n1219) );
XOR2_X1 U943 ( .A(n1113), .B(KEYINPUT23), .Z(n1220) );
XOR2_X1 U944 ( .A(n1221), .B(n1222), .Z(n1113) );
XNOR2_X1 U945 ( .A(G101), .B(G107), .ZN(n1221) );
NAND2_X1 U946 ( .A1(n1223), .A2(n1224), .ZN(n1213) );
OR2_X1 U947 ( .A1(n1109), .A2(n1225), .ZN(n1224) );
XOR2_X1 U948 ( .A(n1226), .B(KEYINPUT48), .Z(n1223) );
NAND2_X1 U949 ( .A1(n1225), .A2(n1109), .ZN(n1226) );
NAND2_X1 U950 ( .A1(G227), .A2(n1044), .ZN(n1109) );
XNOR2_X1 U951 ( .A(n1112), .B(KEYINPUT50), .ZN(n1225) );
XNOR2_X1 U952 ( .A(G110), .B(G140), .ZN(n1112) );
XOR2_X1 U953 ( .A(n1052), .B(KEYINPUT15), .Z(n1111) );
XOR2_X1 U954 ( .A(G131), .B(n1227), .Z(n1052) );
XOR2_X1 U955 ( .A(G137), .B(G134), .Z(n1227) );
XOR2_X1 U956 ( .A(G469), .B(KEYINPUT25), .Z(n1210) );
NAND2_X1 U957 ( .A1(n1228), .A2(n1184), .ZN(n1014) );
NAND2_X1 U958 ( .A1(n1229), .A2(n1185), .ZN(n1184) );
XNOR2_X1 U959 ( .A(G221), .B(KEYINPUT0), .ZN(n1228) );
INV_X1 U960 ( .A(n1175), .ZN(n1181) );
NAND2_X1 U961 ( .A1(n988), .A2(n1230), .ZN(n1175) );
NAND4_X1 U962 ( .A1(G902), .A2(n1076), .A3(n1169), .A4(n1059), .ZN(n1230) );
INV_X1 U963 ( .A(G898), .ZN(n1059) );
INV_X1 U964 ( .A(n1170), .ZN(n1076) );
XOR2_X1 U965 ( .A(n1044), .B(KEYINPUT62), .Z(n1170) );
NAND3_X1 U966 ( .A1(n1169), .A2(n1044), .A3(n1231), .ZN(n988) );
XNOR2_X1 U967 ( .A(G952), .B(KEYINPUT60), .ZN(n1231) );
NAND2_X1 U968 ( .A1(G237), .A2(n1229), .ZN(n1169) );
XNOR2_X1 U969 ( .A(G234), .B(KEYINPUT24), .ZN(n1229) );
NAND2_X1 U970 ( .A1(n1003), .A2(n1004), .ZN(n1176) );
NAND2_X1 U971 ( .A1(G214), .A2(n1232), .ZN(n1004) );
XOR2_X1 U972 ( .A(n1026), .B(n1029), .Z(n1003) );
NAND2_X1 U973 ( .A1(G210), .A2(n1232), .ZN(n1029) );
NAND2_X1 U974 ( .A1(n1233), .A2(n1207), .ZN(n1232) );
XNOR2_X1 U975 ( .A(KEYINPUT53), .B(n1185), .ZN(n1233) );
NAND2_X1 U976 ( .A1(n1234), .A2(n1185), .ZN(n1026) );
XOR2_X1 U977 ( .A(n1146), .B(n1235), .Z(n1234) );
XOR2_X1 U978 ( .A(n1150), .B(n1236), .Z(n1235) );
NOR2_X1 U979 ( .A1(KEYINPUT44), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U980 ( .A(n1238), .B(n1197), .ZN(n1237) );
NAND2_X1 U981 ( .A1(KEYINPUT54), .A2(n1149), .ZN(n1238) );
XNOR2_X1 U982 ( .A(n1051), .B(KEYINPUT7), .ZN(n1149) );
XOR2_X1 U983 ( .A(n1239), .B(n1240), .Z(n1051) );
INV_X1 U984 ( .A(n1199), .ZN(n1240) );
NOR2_X1 U985 ( .A1(n1058), .A2(G953), .ZN(n1150) );
INV_X1 U986 ( .A(G224), .ZN(n1058) );
XNOR2_X1 U987 ( .A(n1241), .B(n1242), .ZN(n1146) );
XOR2_X1 U988 ( .A(n1068), .B(n1063), .Z(n1242) );
XNOR2_X1 U989 ( .A(G110), .B(n1243), .ZN(n1063) );
NOR2_X1 U990 ( .A1(G122), .A2(KEYINPUT63), .ZN(n1243) );
XOR2_X1 U991 ( .A(n1244), .B(n1245), .Z(n1068) );
XNOR2_X1 U992 ( .A(KEYINPUT20), .B(n1166), .ZN(n1245) );
INV_X1 U993 ( .A(G101), .ZN(n1166) );
NAND2_X1 U994 ( .A1(n1246), .A2(n1247), .ZN(n1244) );
NAND2_X1 U995 ( .A1(n1222), .A2(n1248), .ZN(n1247) );
XOR2_X1 U996 ( .A(KEYINPUT55), .B(n1249), .Z(n1246) );
NOR2_X1 U997 ( .A1(n1222), .A2(n1248), .ZN(n1249) );
INV_X1 U998 ( .A(G107), .ZN(n1248) );
INV_X1 U999 ( .A(n1067), .ZN(n1241) );
XNOR2_X1 U1000 ( .A(n1250), .B(G113), .ZN(n1067) );
NAND2_X1 U1001 ( .A1(KEYINPUT47), .A2(n1204), .ZN(n1250) );
XOR2_X1 U1002 ( .A(G116), .B(n1251), .Z(n1204) );
XOR2_X1 U1003 ( .A(KEYINPUT51), .B(G119), .Z(n1251) );
NOR2_X1 U1004 ( .A1(n1155), .A2(n1156), .ZN(n1030) );
XNOR2_X1 U1005 ( .A(n1252), .B(G475), .ZN(n1156) );
NAND2_X1 U1006 ( .A1(n1253), .A2(n1185), .ZN(n1252) );
XNOR2_X1 U1007 ( .A(n1090), .B(KEYINPUT46), .ZN(n1253) );
XNOR2_X1 U1008 ( .A(n1254), .B(n1255), .ZN(n1090) );
XNOR2_X1 U1009 ( .A(n1222), .B(n1256), .ZN(n1255) );
XNOR2_X1 U1010 ( .A(n1257), .B(n1199), .ZN(n1256) );
XOR2_X1 U1011 ( .A(G146), .B(KEYINPUT42), .Z(n1199) );
NAND2_X1 U1012 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND4_X1 U1013 ( .A1(G214), .A2(G143), .A3(n1207), .A4(n1044), .ZN(n1259) );
NAND2_X1 U1014 ( .A1(n1260), .A2(n1261), .ZN(n1258) );
NAND3_X1 U1015 ( .A1(n1207), .A2(n1044), .A3(G214), .ZN(n1261) );
INV_X1 U1016 ( .A(G953), .ZN(n1044) );
INV_X1 U1017 ( .A(G237), .ZN(n1207) );
XNOR2_X1 U1018 ( .A(G143), .B(KEYINPUT10), .ZN(n1260) );
XNOR2_X1 U1019 ( .A(G104), .B(KEYINPUT49), .ZN(n1222) );
XOR2_X1 U1020 ( .A(n1262), .B(n1263), .Z(n1254) );
XNOR2_X1 U1021 ( .A(G131), .B(n1264), .ZN(n1263) );
NAND3_X1 U1022 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1264) );
NAND2_X1 U1023 ( .A1(G113), .A2(n1268), .ZN(n1267) );
OR3_X1 U1024 ( .A1(n1268), .A2(G113), .A3(n1171), .ZN(n1266) );
INV_X1 U1025 ( .A(KEYINPUT32), .ZN(n1268) );
NAND2_X1 U1026 ( .A1(n1269), .A2(n1171), .ZN(n1265) );
NAND2_X1 U1027 ( .A1(n1270), .A2(KEYINPUT32), .ZN(n1269) );
XNOR2_X1 U1028 ( .A(G113), .B(KEYINPUT39), .ZN(n1270) );
NAND2_X1 U1029 ( .A1(n1271), .A2(KEYINPUT3), .ZN(n1262) );
XOR2_X1 U1030 ( .A(n1272), .B(G140), .Z(n1271) );
NAND2_X1 U1031 ( .A1(KEYINPUT61), .A2(n1197), .ZN(n1272) );
INV_X1 U1032 ( .A(G125), .ZN(n1197) );
XNOR2_X1 U1033 ( .A(n1273), .B(G478), .ZN(n1155) );
NAND2_X1 U1034 ( .A1(n1086), .A2(n1185), .ZN(n1273) );
INV_X1 U1035 ( .A(G902), .ZN(n1185) );
XNOR2_X1 U1036 ( .A(n1274), .B(n1275), .ZN(n1086) );
XOR2_X1 U1037 ( .A(G116), .B(n1276), .Z(n1275) );
XNOR2_X1 U1038 ( .A(G134), .B(n1171), .ZN(n1276) );
INV_X1 U1039 ( .A(G122), .ZN(n1171) );
XOR2_X1 U1040 ( .A(n1277), .B(n1278), .Z(n1274) );
NOR3_X1 U1041 ( .A1(n1279), .A2(G953), .A3(n1280), .ZN(n1278) );
INV_X1 U1042 ( .A(G217), .ZN(n1280) );
XOR2_X1 U1043 ( .A(KEYINPUT59), .B(G234), .Z(n1279) );
XNOR2_X1 U1044 ( .A(G107), .B(n1281), .ZN(n1277) );
NOR2_X1 U1045 ( .A1(KEYINPUT40), .A2(n1239), .ZN(n1281) );
XNOR2_X1 U1046 ( .A(G128), .B(G143), .ZN(n1239) );
endmodule


