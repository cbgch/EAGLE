//Key = 1101111110001000010000011010011011100001111011101000010110100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380;

XNOR2_X1 U761 ( .A(G107), .B(n1054), .ZN(G9) );
NAND3_X1 U762 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(G75) );
NOR3_X1 U764 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR3_X1 U765 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NOR3_X1 U766 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
AND4_X1 U767 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1055), .ZN(n1068) );
NOR3_X1 U768 ( .A1(n1069), .A2(n1072), .A3(n1073), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR3_X1 U771 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
NOR2_X1 U772 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XNOR2_X1 U773 ( .A(KEYINPUT32), .B(n1083), .ZN(n1082) );
NOR2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1078) );
NOR3_X1 U775 ( .A1(n1085), .A2(n1086), .A3(n1083), .ZN(n1074) );
XOR2_X1 U776 ( .A(n1087), .B(KEYINPUT0), .Z(n1066) );
NAND4_X1 U777 ( .A1(n1070), .A2(n1088), .A3(n1089), .A4(n1071), .ZN(n1087) );
NAND3_X1 U778 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1060) );
NAND3_X1 U779 ( .A1(n1055), .A2(n1093), .A3(n1070), .ZN(n1092) );
NOR2_X1 U780 ( .A1(n1073), .A2(n1085), .ZN(n1070) );
NAND2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND4_X1 U782 ( .A1(n1064), .A2(n1086), .A3(n1089), .A4(n1096), .ZN(n1095) );
NOR2_X1 U783 ( .A1(n1076), .A2(KEYINPUT9), .ZN(n1086) );
INV_X1 U784 ( .A(n1097), .ZN(n1094) );
NOR3_X1 U785 ( .A1(n1098), .A2(G953), .A3(G952), .ZN(n1058) );
INV_X1 U786 ( .A(n1090), .ZN(n1098) );
NAND4_X1 U787 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1090) );
NOR4_X1 U788 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1102) );
NOR2_X1 U789 ( .A1(n1107), .A2(n1108), .ZN(n1101) );
NOR2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U791 ( .A(G478), .B(KEYINPUT36), .ZN(n1110) );
INV_X1 U792 ( .A(n1111), .ZN(n1107) );
XNOR2_X1 U793 ( .A(KEYINPUT44), .B(n1089), .ZN(n1100) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(n1099) );
NOR2_X1 U795 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U796 ( .A1(KEYINPUT11), .A2(n1116), .ZN(n1115) );
AND2_X1 U797 ( .A1(KEYINPUT25), .A2(n1116), .ZN(n1114) );
INV_X1 U798 ( .A(n1117), .ZN(n1116) );
XOR2_X1 U799 ( .A(n1118), .B(n1119), .Z(G72) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR3_X1 U801 ( .A1(n1122), .A2(KEYINPUT16), .A3(G953), .ZN(n1121) );
NOR2_X1 U802 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
XNOR2_X1 U803 ( .A(n1125), .B(n1126), .ZN(n1124) );
NAND2_X1 U804 ( .A1(KEYINPUT23), .A2(n1127), .ZN(n1125) );
XOR2_X1 U805 ( .A(n1128), .B(n1129), .Z(n1127) );
XNOR2_X1 U806 ( .A(n1130), .B(n1131), .ZN(n1129) );
NOR2_X1 U807 ( .A1(G900), .A2(n1091), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1132), .A2(n1091), .ZN(n1118) );
AND2_X1 U809 ( .A1(G227), .A2(G900), .ZN(n1132) );
XOR2_X1 U810 ( .A(n1133), .B(n1134), .Z(G69) );
XOR2_X1 U811 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U812 ( .A1(n1137), .A2(n1091), .ZN(n1136) );
XOR2_X1 U813 ( .A(n1138), .B(KEYINPUT45), .Z(n1137) );
NAND2_X1 U814 ( .A1(G898), .A2(G224), .ZN(n1138) );
NAND3_X1 U815 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1135) );
NAND2_X1 U816 ( .A1(G953), .A2(n1142), .ZN(n1141) );
NAND2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
NAND2_X1 U818 ( .A1(n1091), .A2(n1145), .ZN(n1133) );
NAND2_X1 U819 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U820 ( .A(KEYINPUT57), .B(n1148), .Z(n1147) );
NOR2_X1 U821 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1151), .A2(n1152), .ZN(G66) );
XOR2_X1 U823 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR3_X1 U824 ( .A1(n1155), .A2(KEYINPUT49), .A3(n1156), .ZN(n1153) );
NOR2_X1 U825 ( .A1(n1151), .A2(n1157), .ZN(G63) );
NOR2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U827 ( .A(n1160), .B(KEYINPUT5), .Z(n1159) );
NAND2_X1 U828 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U829 ( .A1(n1161), .A2(n1162), .ZN(n1158) );
NOR2_X1 U830 ( .A1(n1155), .A2(n1163), .ZN(n1162) );
NOR2_X1 U831 ( .A1(n1151), .A2(n1164), .ZN(G60) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U833 ( .A1(n1167), .A2(n1155), .ZN(n1165) );
XNOR2_X1 U834 ( .A(n1149), .B(n1168), .ZN(G6) );
XNOR2_X1 U835 ( .A(KEYINPUT62), .B(n1169), .ZN(n1168) );
NOR2_X1 U836 ( .A1(n1151), .A2(n1170), .ZN(G57) );
XNOR2_X1 U837 ( .A(n1171), .B(n1172), .ZN(n1170) );
XNOR2_X1 U838 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR2_X1 U839 ( .A1(KEYINPUT54), .A2(n1175), .ZN(n1174) );
XOR2_X1 U840 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U841 ( .A1(n1178), .A2(n1155), .ZN(n1176) );
NOR2_X1 U842 ( .A1(n1151), .A2(n1179), .ZN(G54) );
XOR2_X1 U843 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U844 ( .A(n1182), .B(n1183), .Z(n1181) );
NOR2_X1 U845 ( .A1(n1184), .A2(n1155), .ZN(n1183) );
NOR2_X1 U846 ( .A1(KEYINPUT51), .A2(n1185), .ZN(n1182) );
NOR3_X1 U847 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
NOR2_X1 U848 ( .A1(KEYINPUT24), .A2(n1189), .ZN(n1188) );
NOR3_X1 U849 ( .A1(n1131), .A2(n1190), .A3(n1191), .ZN(n1187) );
NOR2_X1 U850 ( .A1(n1192), .A2(n1193), .ZN(n1186) );
NOR2_X1 U851 ( .A1(n1194), .A2(n1191), .ZN(n1192) );
INV_X1 U852 ( .A(KEYINPUT24), .ZN(n1191) );
XNOR2_X1 U853 ( .A(n1189), .B(KEYINPUT35), .ZN(n1194) );
XOR2_X1 U854 ( .A(n1195), .B(n1196), .Z(n1180) );
NOR2_X1 U855 ( .A1(n1151), .A2(n1197), .ZN(G51) );
XOR2_X1 U856 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U857 ( .A1(n1117), .A2(n1155), .ZN(n1199) );
NAND2_X1 U858 ( .A1(G902), .A2(n1062), .ZN(n1155) );
NAND4_X1 U859 ( .A1(n1200), .A2(n1122), .A3(n1201), .A4(n1146), .ZN(n1062) );
AND3_X1 U860 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1146) );
NAND2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U862 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U863 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U864 ( .A1(n1211), .A2(n1088), .ZN(n1207) );
INV_X1 U865 ( .A(n1150), .ZN(n1201) );
NAND2_X1 U866 ( .A1(n1212), .A2(n1213), .ZN(n1150) );
NAND2_X1 U867 ( .A1(n1056), .A2(n1214), .ZN(n1213) );
NAND2_X1 U868 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U869 ( .A1(n1055), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U870 ( .A(KEYINPUT18), .B(n1081), .ZN(n1217) );
INV_X1 U871 ( .A(n1057), .ZN(n1081) );
AND4_X1 U872 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1122) );
NOR4_X1 U873 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
NOR2_X1 U874 ( .A1(n1226), .A2(n1227), .ZN(n1220) );
INV_X1 U875 ( .A(n1228), .ZN(n1227) );
NOR3_X1 U876 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1226) );
XNOR2_X1 U877 ( .A(n1211), .B(KEYINPUT20), .ZN(n1230) );
XNOR2_X1 U878 ( .A(n1149), .B(KEYINPUT10), .ZN(n1200) );
AND3_X1 U879 ( .A1(n1055), .A2(n1056), .A3(n1211), .ZN(n1149) );
NAND2_X1 U880 ( .A1(n1232), .A2(KEYINPUT55), .ZN(n1198) );
XNOR2_X1 U881 ( .A(n1233), .B(n1234), .ZN(n1232) );
XNOR2_X1 U882 ( .A(n1235), .B(n1236), .ZN(n1233) );
NOR2_X1 U883 ( .A1(KEYINPUT50), .A2(n1237), .ZN(n1236) );
NOR2_X1 U884 ( .A1(n1091), .A2(G952), .ZN(n1151) );
XOR2_X1 U885 ( .A(n1218), .B(n1238), .Z(G48) );
XNOR2_X1 U886 ( .A(G146), .B(KEYINPUT2), .ZN(n1238) );
NAND3_X1 U887 ( .A1(n1210), .A2(n1239), .A3(n1211), .ZN(n1218) );
XNOR2_X1 U888 ( .A(n1219), .B(n1240), .ZN(G45) );
NOR2_X1 U889 ( .A1(KEYINPUT31), .A2(n1241), .ZN(n1240) );
NAND4_X1 U890 ( .A1(n1088), .A2(n1239), .A3(n1104), .A4(n1242), .ZN(n1219) );
XOR2_X1 U891 ( .A(n1243), .B(n1244), .Z(G42) );
XOR2_X1 U892 ( .A(KEYINPUT21), .B(G140), .Z(n1244) );
AND2_X1 U893 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
XNOR2_X1 U894 ( .A(n1225), .B(n1247), .ZN(G39) );
NAND2_X1 U895 ( .A1(KEYINPUT41), .A2(G137), .ZN(n1247) );
AND3_X1 U896 ( .A1(n1245), .A2(n1210), .A3(n1209), .ZN(n1225) );
XOR2_X1 U897 ( .A(n1248), .B(n1249), .Z(G36) );
XOR2_X1 U898 ( .A(KEYINPUT34), .B(G134), .Z(n1249) );
NOR2_X1 U899 ( .A1(n1224), .A2(KEYINPUT22), .ZN(n1248) );
AND3_X1 U900 ( .A1(n1245), .A2(n1057), .A3(n1088), .ZN(n1224) );
XOR2_X1 U901 ( .A(G131), .B(n1223), .Z(G33) );
AND3_X1 U902 ( .A1(n1088), .A2(n1245), .A3(n1211), .ZN(n1223) );
INV_X1 U903 ( .A(n1231), .ZN(n1245) );
NAND4_X1 U904 ( .A1(n1096), .A2(n1250), .A3(n1069), .A4(n1251), .ZN(n1231) );
XOR2_X1 U905 ( .A(G128), .B(n1222), .Z(G30) );
AND3_X1 U906 ( .A1(n1239), .A2(n1057), .A3(n1210), .ZN(n1222) );
AND2_X1 U907 ( .A1(n1252), .A2(n1251), .ZN(n1239) );
XNOR2_X1 U908 ( .A(G101), .B(n1212), .ZN(G3) );
NAND3_X1 U909 ( .A1(n1088), .A2(n1056), .A3(n1209), .ZN(n1212) );
AND2_X1 U910 ( .A1(n1252), .A2(n1253), .ZN(n1056) );
XNOR2_X1 U911 ( .A(G125), .B(n1228), .ZN(G27) );
NAND3_X1 U912 ( .A1(n1246), .A2(n1251), .A3(n1097), .ZN(n1228) );
NAND2_X1 U913 ( .A1(n1073), .A2(n1254), .ZN(n1251) );
NAND4_X1 U914 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1256), .ZN(n1254) );
INV_X1 U915 ( .A(G900), .ZN(n1256) );
NOR2_X1 U916 ( .A1(n1229), .A2(n1084), .ZN(n1246) );
XNOR2_X1 U917 ( .A(G122), .B(n1202), .ZN(G24) );
NAND4_X1 U918 ( .A1(n1205), .A2(n1055), .A3(n1104), .A4(n1242), .ZN(n1202) );
INV_X1 U919 ( .A(n1083), .ZN(n1055) );
NAND2_X1 U920 ( .A1(n1257), .A2(n1258), .ZN(n1083) );
XNOR2_X1 U921 ( .A(G119), .B(n1259), .ZN(G21) );
NAND4_X1 U922 ( .A1(KEYINPUT48), .A2(n1205), .A3(n1209), .A4(n1210), .ZN(n1259) );
AND2_X1 U923 ( .A1(n1106), .A2(n1103), .ZN(n1210) );
XNOR2_X1 U924 ( .A(G116), .B(n1203), .ZN(G18) );
NAND3_X1 U925 ( .A1(n1088), .A2(n1057), .A3(n1205), .ZN(n1203) );
NOR2_X1 U926 ( .A1(n1104), .A2(n1260), .ZN(n1057) );
XNOR2_X1 U927 ( .A(G113), .B(n1261), .ZN(G15) );
NAND4_X1 U928 ( .A1(KEYINPUT6), .A2(n1205), .A3(n1211), .A4(n1088), .ZN(n1261) );
AND2_X1 U929 ( .A1(n1106), .A2(n1258), .ZN(n1088) );
XNOR2_X1 U930 ( .A(n1103), .B(KEYINPUT27), .ZN(n1258) );
INV_X1 U931 ( .A(n1084), .ZN(n1211) );
NAND2_X1 U932 ( .A1(n1260), .A2(n1104), .ZN(n1084) );
INV_X1 U933 ( .A(n1242), .ZN(n1260) );
AND2_X1 U934 ( .A1(n1097), .A2(n1253), .ZN(n1205) );
NOR3_X1 U935 ( .A1(n1105), .A2(n1096), .A3(n1069), .ZN(n1097) );
XNOR2_X1 U936 ( .A(n1262), .B(n1263), .ZN(G12) );
NOR4_X1 U937 ( .A1(KEYINPUT43), .A2(n1264), .A3(n1265), .A4(n1215), .ZN(n1263) );
INV_X1 U938 ( .A(n1079), .ZN(n1215) );
NOR2_X1 U939 ( .A1(n1229), .A2(n1085), .ZN(n1079) );
INV_X1 U940 ( .A(n1209), .ZN(n1085) );
NOR2_X1 U941 ( .A1(n1242), .A2(n1104), .ZN(n1209) );
XOR2_X1 U942 ( .A(n1266), .B(n1167), .Z(n1104) );
INV_X1 U943 ( .A(G475), .ZN(n1167) );
OR2_X1 U944 ( .A1(n1166), .A2(G902), .ZN(n1266) );
XNOR2_X1 U945 ( .A(n1267), .B(n1268), .ZN(n1166) );
XOR2_X1 U946 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U947 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U948 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U949 ( .A(n1275), .B(KEYINPUT46), .Z(n1274) );
NAND2_X1 U950 ( .A1(G104), .A2(n1276), .ZN(n1275) );
NOR2_X1 U951 ( .A1(G104), .A2(n1276), .ZN(n1273) );
XNOR2_X1 U952 ( .A(G113), .B(n1277), .ZN(n1276) );
XNOR2_X1 U953 ( .A(KEYINPUT30), .B(n1278), .ZN(n1277) );
NAND3_X1 U954 ( .A1(n1279), .A2(n1091), .A3(G214), .ZN(n1271) );
NAND2_X1 U955 ( .A1(n1280), .A2(KEYINPUT29), .ZN(n1269) );
XNOR2_X1 U956 ( .A(G146), .B(n1126), .ZN(n1280) );
XOR2_X1 U957 ( .A(n1281), .B(n1282), .Z(n1267) );
NOR2_X1 U958 ( .A1(KEYINPUT37), .A2(n1241), .ZN(n1282) );
NAND2_X1 U959 ( .A1(n1283), .A2(n1111), .ZN(n1242) );
NAND2_X1 U960 ( .A1(n1109), .A2(n1163), .ZN(n1111) );
OR2_X1 U961 ( .A1(n1163), .A2(n1109), .ZN(n1283) );
NOR2_X1 U962 ( .A1(n1161), .A2(G902), .ZN(n1109) );
AND2_X1 U963 ( .A1(n1284), .A2(n1285), .ZN(n1161) );
NAND2_X1 U964 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U965 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U966 ( .A1(G217), .A2(n1290), .ZN(n1286) );
XOR2_X1 U967 ( .A(n1291), .B(KEYINPUT52), .Z(n1284) );
NAND4_X1 U968 ( .A1(n1288), .A2(G217), .A3(n1290), .A4(n1289), .ZN(n1291) );
NAND2_X1 U969 ( .A1(n1292), .A2(n1293), .ZN(n1289) );
XOR2_X1 U970 ( .A(n1294), .B(n1295), .Z(n1292) );
XOR2_X1 U971 ( .A(n1296), .B(KEYINPUT61), .Z(n1288) );
NAND2_X1 U972 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
INV_X1 U973 ( .A(n1293), .ZN(n1298) );
XNOR2_X1 U974 ( .A(n1299), .B(n1300), .ZN(n1293) );
XOR2_X1 U975 ( .A(G116), .B(G107), .Z(n1300) );
NAND2_X1 U976 ( .A1(KEYINPUT53), .A2(G122), .ZN(n1299) );
XNOR2_X1 U977 ( .A(n1294), .B(n1295), .ZN(n1297) );
NOR2_X1 U978 ( .A1(n1301), .A2(G134), .ZN(n1294) );
INV_X1 U979 ( .A(KEYINPUT39), .ZN(n1301) );
INV_X1 U980 ( .A(G478), .ZN(n1163) );
NAND2_X1 U981 ( .A1(n1257), .A2(n1103), .ZN(n1229) );
NAND3_X1 U982 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1103) );
NAND2_X1 U983 ( .A1(n1305), .A2(n1154), .ZN(n1304) );
OR3_X1 U984 ( .A1(n1154), .A2(n1305), .A3(G902), .ZN(n1303) );
NOR2_X1 U985 ( .A1(n1156), .A2(G234), .ZN(n1305) );
INV_X1 U986 ( .A(G217), .ZN(n1156) );
XNOR2_X1 U987 ( .A(n1306), .B(n1307), .ZN(n1154) );
XOR2_X1 U988 ( .A(G137), .B(n1308), .Z(n1307) );
NOR2_X1 U989 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U990 ( .A(n1311), .B(KEYINPUT17), .Z(n1310) );
NAND2_X1 U991 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NOR2_X1 U992 ( .A1(n1312), .A2(n1313), .ZN(n1309) );
XNOR2_X1 U993 ( .A(G110), .B(n1314), .ZN(n1313) );
XOR2_X1 U994 ( .A(G128), .B(G119), .Z(n1314) );
XNOR2_X1 U995 ( .A(n1315), .B(n1316), .ZN(n1312) );
NOR2_X1 U996 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
AND3_X1 U997 ( .A1(KEYINPUT47), .A2(n1319), .A3(G140), .ZN(n1318) );
NOR2_X1 U998 ( .A1(KEYINPUT47), .A2(n1126), .ZN(n1317) );
XNOR2_X1 U999 ( .A(n1319), .B(G140), .ZN(n1126) );
INV_X1 U1000 ( .A(G146), .ZN(n1315) );
NAND2_X1 U1001 ( .A1(G221), .A2(n1290), .ZN(n1306) );
AND2_X1 U1002 ( .A1(G234), .A2(n1091), .ZN(n1290) );
NAND2_X1 U1003 ( .A1(G902), .A2(G217), .ZN(n1302) );
INV_X1 U1004 ( .A(n1106), .ZN(n1257) );
XOR2_X1 U1005 ( .A(n1320), .B(n1178), .Z(n1106) );
INV_X1 U1006 ( .A(G472), .ZN(n1178) );
NAND2_X1 U1007 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U1008 ( .A(n1177), .B(n1323), .Z(n1321) );
XNOR2_X1 U1009 ( .A(n1173), .B(n1324), .ZN(n1323) );
NOR2_X1 U1010 ( .A1(KEYINPUT60), .A2(n1171), .ZN(n1324) );
NAND3_X1 U1011 ( .A1(n1279), .A2(n1091), .A3(G210), .ZN(n1171) );
XNOR2_X1 U1012 ( .A(n1325), .B(KEYINPUT7), .ZN(n1279) );
XNOR2_X1 U1013 ( .A(n1326), .B(n1327), .ZN(n1177) );
XNOR2_X1 U1014 ( .A(n1328), .B(n1189), .ZN(n1326) );
INV_X1 U1015 ( .A(n1252), .ZN(n1265) );
NOR3_X1 U1016 ( .A1(n1089), .A2(n1096), .A3(n1105), .ZN(n1252) );
INV_X1 U1017 ( .A(n1250), .ZN(n1105) );
NOR2_X1 U1018 ( .A1(n1064), .A2(n1076), .ZN(n1250) );
INV_X1 U1019 ( .A(n1071), .ZN(n1076) );
NAND2_X1 U1020 ( .A1(G221), .A2(n1329), .ZN(n1071) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1322), .ZN(n1329) );
AND2_X1 U1022 ( .A1(G214), .A2(n1330), .ZN(n1064) );
INV_X1 U1023 ( .A(n1063), .ZN(n1096) );
XOR2_X1 U1024 ( .A(n1112), .B(n1117), .Z(n1063) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1330), .ZN(n1117) );
NAND2_X1 U1026 ( .A1(n1325), .A2(n1322), .ZN(n1330) );
INV_X1 U1027 ( .A(G237), .ZN(n1325) );
NAND3_X1 U1028 ( .A1(n1331), .A2(n1322), .A3(n1332), .ZN(n1112) );
XOR2_X1 U1029 ( .A(KEYINPUT1), .B(n1333), .Z(n1332) );
NOR2_X1 U1030 ( .A1(n1235), .A2(n1334), .ZN(n1333) );
NAND2_X1 U1031 ( .A1(n1235), .A2(n1334), .ZN(n1331) );
NAND3_X1 U1032 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
NAND2_X1 U1033 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
OR3_X1 U1034 ( .A1(n1339), .A2(n1338), .A3(n1340), .ZN(n1336) );
NAND2_X1 U1035 ( .A1(n1341), .A2(n1342), .ZN(n1338) );
NAND2_X1 U1036 ( .A1(KEYINPUT8), .A2(n1234), .ZN(n1342) );
XNOR2_X1 U1037 ( .A(n1319), .B(n1131), .ZN(n1234) );
INV_X1 U1038 ( .A(G125), .ZN(n1319) );
OR3_X1 U1039 ( .A1(n1131), .A2(G125), .A3(KEYINPUT8), .ZN(n1341) );
NAND2_X1 U1040 ( .A1(KEYINPUT33), .A2(n1343), .ZN(n1339) );
INV_X1 U1041 ( .A(n1237), .ZN(n1343) );
NAND2_X1 U1042 ( .A1(n1237), .A2(n1340), .ZN(n1335) );
INV_X1 U1043 ( .A(KEYINPUT26), .ZN(n1340) );
NAND2_X1 U1044 ( .A1(G224), .A2(n1091), .ZN(n1237) );
AND2_X1 U1045 ( .A1(n1344), .A2(n1140), .ZN(n1235) );
OR2_X1 U1046 ( .A1(n1144), .A2(n1143), .ZN(n1140) );
NAND2_X1 U1047 ( .A1(n1345), .A2(n1143), .ZN(n1344) );
XOR2_X1 U1048 ( .A(n1346), .B(n1328), .Z(n1143) );
XOR2_X1 U1049 ( .A(G113), .B(n1347), .Z(n1328) );
XOR2_X1 U1050 ( .A(G119), .B(G116), .Z(n1347) );
NAND3_X1 U1051 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1346) );
NAND2_X1 U1052 ( .A1(G101), .A2(n1351), .ZN(n1350) );
NAND2_X1 U1053 ( .A1(KEYINPUT38), .A2(n1352), .ZN(n1349) );
NAND2_X1 U1054 ( .A1(n1353), .A2(n1173), .ZN(n1352) );
XNOR2_X1 U1055 ( .A(KEYINPUT3), .B(n1354), .ZN(n1353) );
NAND2_X1 U1056 ( .A1(n1355), .A2(n1356), .ZN(n1348) );
INV_X1 U1057 ( .A(KEYINPUT38), .ZN(n1356) );
NAND2_X1 U1058 ( .A1(n1357), .A2(n1358), .ZN(n1355) );
NAND3_X1 U1059 ( .A1(KEYINPUT3), .A2(n1173), .A3(n1354), .ZN(n1358) );
OR2_X1 U1060 ( .A1(n1354), .A2(KEYINPUT3), .ZN(n1357) );
XOR2_X1 U1061 ( .A(n1144), .B(KEYINPUT59), .Z(n1345) );
NAND3_X1 U1062 ( .A1(n1359), .A2(n1360), .A3(n1361), .ZN(n1144) );
NAND2_X1 U1063 ( .A1(n1362), .A2(n1262), .ZN(n1361) );
NAND2_X1 U1064 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XNOR2_X1 U1065 ( .A(KEYINPUT56), .B(n1278), .ZN(n1363) );
NAND3_X1 U1066 ( .A1(G110), .A2(n1278), .A3(n1364), .ZN(n1360) );
INV_X1 U1067 ( .A(KEYINPUT15), .ZN(n1364) );
INV_X1 U1068 ( .A(G122), .ZN(n1278) );
NAND2_X1 U1069 ( .A1(KEYINPUT15), .A2(G122), .ZN(n1359) );
INV_X1 U1070 ( .A(n1069), .ZN(n1089) );
XOR2_X1 U1071 ( .A(n1365), .B(n1184), .Z(n1069) );
INV_X1 U1072 ( .A(G469), .ZN(n1184) );
NAND2_X1 U1073 ( .A1(n1366), .A2(n1322), .ZN(n1365) );
INV_X1 U1074 ( .A(G902), .ZN(n1322) );
XOR2_X1 U1075 ( .A(n1195), .B(n1367), .Z(n1366) );
XOR2_X1 U1076 ( .A(n1368), .B(KEYINPUT63), .Z(n1367) );
NAND2_X1 U1077 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
OR2_X1 U1078 ( .A1(n1196), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1079 ( .A(n1372), .B(KEYINPUT28), .Z(n1369) );
NAND2_X1 U1080 ( .A1(n1371), .A2(n1196), .ZN(n1372) );
XOR2_X1 U1081 ( .A(n1327), .B(KEYINPUT12), .Z(n1196) );
XNOR2_X1 U1082 ( .A(n1130), .B(n1373), .ZN(n1327) );
NOR2_X1 U1083 ( .A1(KEYINPUT19), .A2(n1128), .ZN(n1373) );
XNOR2_X1 U1084 ( .A(G134), .B(G137), .ZN(n1128) );
XOR2_X1 U1085 ( .A(n1281), .B(KEYINPUT14), .Z(n1130) );
XNOR2_X1 U1086 ( .A(G131), .B(KEYINPUT13), .ZN(n1281) );
XOR2_X1 U1087 ( .A(n1374), .B(n1190), .Z(n1371) );
INV_X1 U1088 ( .A(n1193), .ZN(n1190) );
XOR2_X1 U1089 ( .A(n1375), .B(n1173), .Z(n1193) );
INV_X1 U1090 ( .A(G101), .ZN(n1173) );
NAND3_X1 U1091 ( .A1(n1376), .A2(n1377), .A3(KEYINPUT4), .ZN(n1375) );
NAND2_X1 U1092 ( .A1(KEYINPUT42), .A2(n1354), .ZN(n1377) );
INV_X1 U1093 ( .A(n1351), .ZN(n1354) );
XOR2_X1 U1094 ( .A(G104), .B(G107), .Z(n1351) );
OR3_X1 U1095 ( .A1(n1169), .A2(G107), .A3(KEYINPUT42), .ZN(n1376) );
INV_X1 U1096 ( .A(G104), .ZN(n1169) );
NAND2_X1 U1097 ( .A1(KEYINPUT58), .A2(n1131), .ZN(n1374) );
INV_X1 U1098 ( .A(n1189), .ZN(n1131) );
XOR2_X1 U1099 ( .A(G146), .B(n1295), .Z(n1189) );
XNOR2_X1 U1100 ( .A(G128), .B(n1241), .ZN(n1295) );
INV_X1 U1101 ( .A(G143), .ZN(n1241) );
XOR2_X1 U1102 ( .A(n1378), .B(n1379), .Z(n1195) );
XNOR2_X1 U1103 ( .A(G140), .B(n1262), .ZN(n1379) );
NAND2_X1 U1104 ( .A1(G227), .A2(n1091), .ZN(n1378) );
XOR2_X1 U1105 ( .A(n1253), .B(KEYINPUT40), .Z(n1264) );
NAND2_X1 U1106 ( .A1(n1073), .A2(n1380), .ZN(n1253) );
NAND4_X1 U1107 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1142), .ZN(n1380) );
INV_X1 U1108 ( .A(G898), .ZN(n1142) );
NAND3_X1 U1109 ( .A1(n1255), .A2(n1091), .A3(G952), .ZN(n1073) );
INV_X1 U1110 ( .A(G953), .ZN(n1091) );
NAND2_X1 U1111 ( .A1(G237), .A2(G234), .ZN(n1255) );
INV_X1 U1112 ( .A(G110), .ZN(n1262) );
endmodule


