//Key = 0010101110010101011010100000101010001011111010111101011000110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358;

XNOR2_X1 U736 ( .A(G107), .B(n1025), .ZN(G9) );
NOR2_X1 U737 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR3_X1 U738 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NOR2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR4_X1 U740 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1031) );
NOR2_X1 U741 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR4_X1 U742 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1037) );
NOR2_X1 U743 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U744 ( .A1(KEYINPUT14), .A2(n1045), .ZN(n1041) );
NOR2_X1 U745 ( .A1(KEYINPUT55), .A2(n1046), .ZN(n1040) );
NOR2_X1 U746 ( .A1(n1047), .A2(n1048), .ZN(n1039) );
NOR2_X1 U747 ( .A1(n1049), .A2(n1050), .ZN(n1035) );
INV_X1 U748 ( .A(KEYINPUT55), .ZN(n1050) );
NOR2_X1 U749 ( .A1(n1046), .A2(n1038), .ZN(n1049) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1034) );
INV_X1 U751 ( .A(KEYINPUT14), .ZN(n1052) );
NOR2_X1 U752 ( .A1(n1045), .A2(n1038), .ZN(n1051) );
INV_X1 U753 ( .A(n1053), .ZN(n1038) );
NOR4_X1 U754 ( .A1(n1054), .A2(n1055), .A3(n1043), .A4(n1047), .ZN(n1033) );
NOR2_X1 U755 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
XOR2_X1 U756 ( .A(KEYINPUT19), .B(n1058), .Z(n1057) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U758 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1028) );
NAND4_X1 U759 ( .A1(n1053), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1063) );
NAND2_X1 U760 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U761 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1055), .ZN(n1053) );
INV_X1 U763 ( .A(n1072), .ZN(n1071) );
NOR3_X1 U764 ( .A1(n1073), .A2(G953), .A3(G952), .ZN(n1026) );
INV_X1 U765 ( .A(n1061), .ZN(n1073) );
NAND4_X1 U766 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1061) );
NOR4_X1 U767 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1070), .ZN(n1077) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1059), .ZN(n1078) );
NAND2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U770 ( .A(G475), .B(KEYINPUT32), .ZN(n1082) );
NOR3_X1 U771 ( .A1(n1084), .A2(n1085), .A3(n1060), .ZN(n1076) );
XOR2_X1 U772 ( .A(n1086), .B(KEYINPUT13), .Z(n1085) );
XNOR2_X1 U773 ( .A(n1087), .B(n1088), .ZN(n1084) );
XNOR2_X1 U774 ( .A(n1089), .B(KEYINPUT21), .ZN(n1075) );
XOR2_X1 U775 ( .A(n1090), .B(G472), .Z(n1074) );
XOR2_X1 U776 ( .A(n1091), .B(n1092), .Z(G72) );
XOR2_X1 U777 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U778 ( .A1(n1095), .A2(n1062), .ZN(n1094) );
NOR2_X1 U779 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U780 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1100), .A2(n1097), .ZN(n1099) );
XOR2_X1 U782 ( .A(n1101), .B(n1102), .Z(n1098) );
XNOR2_X1 U783 ( .A(n1103), .B(n1104), .ZN(n1102) );
XNOR2_X1 U784 ( .A(n1105), .B(n1106), .ZN(n1101) );
NOR2_X1 U785 ( .A1(KEYINPUT34), .A2(n1107), .ZN(n1106) );
NAND2_X1 U786 ( .A1(n1062), .A2(n1108), .ZN(n1091) );
NAND2_X1 U787 ( .A1(n1109), .A2(n1110), .ZN(G69) );
NAND2_X1 U788 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U789 ( .A(n1113), .B(n1114), .Z(n1109) );
NOR2_X1 U790 ( .A1(G953), .A2(n1115), .ZN(n1114) );
NOR3_X1 U791 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
XNOR2_X1 U792 ( .A(KEYINPUT23), .B(n1119), .ZN(n1118) );
XNOR2_X1 U793 ( .A(n1120), .B(KEYINPUT25), .ZN(n1117) );
NAND3_X1 U794 ( .A1(n1121), .A2(n1025), .A3(n1122), .ZN(n1116) );
INV_X1 U795 ( .A(n1123), .ZN(n1121) );
NAND2_X1 U796 ( .A1(n1124), .A2(n1125), .ZN(n1113) );
XOR2_X1 U797 ( .A(KEYINPUT6), .B(n1111), .Z(n1125) );
AND2_X1 U798 ( .A1(G953), .A2(n1126), .ZN(n1111) );
NAND2_X1 U799 ( .A1(G898), .A2(G224), .ZN(n1126) );
INV_X1 U800 ( .A(n1112), .ZN(n1124) );
NAND2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(n1112) );
NAND2_X1 U802 ( .A1(n1100), .A2(n1129), .ZN(n1128) );
XOR2_X1 U803 ( .A(n1130), .B(n1131), .Z(n1127) );
XNOR2_X1 U804 ( .A(n1132), .B(n1133), .ZN(n1130) );
NAND2_X1 U805 ( .A1(KEYINPUT53), .A2(n1134), .ZN(n1133) );
NAND2_X1 U806 ( .A1(KEYINPUT22), .A2(n1135), .ZN(n1132) );
NOR2_X1 U807 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XNOR2_X1 U808 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U809 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U810 ( .A1(n1136), .A2(n1142), .ZN(G63) );
XOR2_X1 U811 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U812 ( .A1(n1087), .A2(n1141), .ZN(n1144) );
INV_X1 U813 ( .A(G478), .ZN(n1087) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1145), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1146), .B(n1147), .ZN(n1145) );
AND2_X1 U816 ( .A1(G475), .A2(n1148), .ZN(n1147) );
XNOR2_X1 U817 ( .A(G104), .B(n1119), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1136), .A2(n1149), .ZN(G57) );
NOR3_X1 U819 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1149) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
AND3_X1 U821 ( .A1(n1154), .A2(n1153), .A3(n1155), .ZN(n1151) );
INV_X1 U822 ( .A(KEYINPUT60), .ZN(n1154) );
NOR2_X1 U823 ( .A1(n1155), .A2(n1156), .ZN(n1150) );
NOR2_X1 U824 ( .A1(KEYINPUT60), .A2(n1157), .ZN(n1156) );
XNOR2_X1 U825 ( .A(KEYINPUT24), .B(n1153), .ZN(n1157) );
NAND2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
NAND2_X1 U827 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U828 ( .A1(n1148), .A2(G472), .ZN(n1161) );
INV_X1 U829 ( .A(n1162), .ZN(n1160) );
NAND3_X1 U830 ( .A1(n1148), .A2(G472), .A3(n1162), .ZN(n1158) );
XNOR2_X1 U831 ( .A(n1163), .B(n1164), .ZN(n1162) );
XNOR2_X1 U832 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U833 ( .A1(KEYINPUT48), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U834 ( .A(n1168), .B(KEYINPUT3), .ZN(n1163) );
AND2_X1 U835 ( .A1(n1169), .A2(n1170), .ZN(n1155) );
NAND2_X1 U836 ( .A1(n1171), .A2(G101), .ZN(n1170) );
XOR2_X1 U837 ( .A(n1172), .B(KEYINPUT12), .Z(n1169) );
OR2_X1 U838 ( .A1(G101), .A2(n1171), .ZN(n1172) );
NOR2_X1 U839 ( .A1(n1136), .A2(n1173), .ZN(G54) );
XOR2_X1 U840 ( .A(n1174), .B(n1175), .Z(n1173) );
AND2_X1 U841 ( .A1(G469), .A2(n1148), .ZN(n1175) );
INV_X1 U842 ( .A(n1141), .ZN(n1148) );
NAND3_X1 U843 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1174) );
NAND2_X1 U844 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
OR3_X1 U845 ( .A1(n1180), .A2(n1179), .A3(n1181), .ZN(n1177) );
INV_X1 U846 ( .A(KEYINPUT51), .ZN(n1181) );
XOR2_X1 U847 ( .A(n1103), .B(n1182), .Z(n1179) );
XNOR2_X1 U848 ( .A(n1168), .B(n1183), .ZN(n1182) );
NAND2_X1 U849 ( .A1(KEYINPUT59), .A2(n1184), .ZN(n1180) );
OR2_X1 U850 ( .A1(n1184), .A2(KEYINPUT51), .ZN(n1176) );
XNOR2_X1 U851 ( .A(n1185), .B(KEYINPUT44), .ZN(n1184) );
NOR2_X1 U852 ( .A1(n1136), .A2(n1186), .ZN(G51) );
XOR2_X1 U853 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U854 ( .A1(n1189), .A2(n1141), .ZN(n1188) );
NAND2_X1 U855 ( .A1(G902), .A2(n1030), .ZN(n1141) );
NAND4_X1 U856 ( .A1(n1120), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1030) );
AND3_X1 U857 ( .A1(n1119), .A2(n1025), .A3(n1122), .ZN(n1192) );
OR3_X1 U858 ( .A1(n1043), .A2(n1193), .A3(n1044), .ZN(n1025) );
INV_X1 U859 ( .A(n1065), .ZN(n1043) );
OR2_X1 U860 ( .A1(n1045), .A2(n1193), .ZN(n1119) );
NAND2_X1 U861 ( .A1(n1194), .A2(n1065), .ZN(n1045) );
XNOR2_X1 U862 ( .A(n1123), .B(KEYINPUT63), .ZN(n1191) );
INV_X1 U863 ( .A(n1108), .ZN(n1190) );
NAND4_X1 U864 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1108) );
NOR4_X1 U865 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NAND2_X1 U866 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
NAND2_X1 U867 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U868 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U869 ( .A1(n1209), .A2(n1210), .ZN(n1205) );
AND4_X1 U870 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1120) );
NOR2_X1 U871 ( .A1(n1215), .A2(n1216), .ZN(n1187) );
XOR2_X1 U872 ( .A(KEYINPUT0), .B(n1217), .Z(n1216) );
NOR2_X1 U873 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NOR2_X1 U874 ( .A1(n1220), .A2(n1221), .ZN(n1215) );
XNOR2_X1 U875 ( .A(n1218), .B(KEYINPUT10), .ZN(n1221) );
INV_X1 U876 ( .A(n1219), .ZN(n1220) );
NOR2_X1 U877 ( .A1(n1062), .A2(G952), .ZN(n1136) );
XNOR2_X1 U878 ( .A(G146), .B(n1195), .ZN(G48) );
NAND3_X1 U879 ( .A1(n1194), .A2(n1210), .A3(n1209), .ZN(n1195) );
INV_X1 U880 ( .A(n1222), .ZN(n1209) );
XNOR2_X1 U881 ( .A(G143), .B(n1196), .ZN(G45) );
NAND4_X1 U882 ( .A1(n1208), .A2(n1210), .A3(n1223), .A4(n1224), .ZN(n1196) );
XOR2_X1 U883 ( .A(n1225), .B(n1226), .Z(G42) );
XOR2_X1 U884 ( .A(KEYINPUT46), .B(G140), .Z(n1226) );
NAND2_X1 U885 ( .A1(KEYINPUT38), .A2(n1202), .ZN(n1225) );
AND4_X1 U886 ( .A1(n1056), .A2(n1227), .A3(n1194), .A4(n1228), .ZN(n1202) );
NOR2_X1 U887 ( .A1(n1048), .A2(n1032), .ZN(n1228) );
XNOR2_X1 U888 ( .A(n1201), .B(n1229), .ZN(G39) );
NAND2_X1 U889 ( .A1(KEYINPUT41), .A2(G137), .ZN(n1229) );
NOR3_X1 U890 ( .A1(n1032), .A2(n1047), .A3(n1222), .ZN(n1201) );
XOR2_X1 U891 ( .A(G134), .B(n1230), .Z(G36) );
NOR4_X1 U892 ( .A1(KEYINPUT9), .A2(n1044), .A3(n1231), .A4(n1032), .ZN(n1230) );
XOR2_X1 U893 ( .A(G131), .B(n1200), .Z(G33) );
AND3_X1 U894 ( .A1(n1208), .A2(n1194), .A3(n1207), .ZN(n1200) );
INV_X1 U895 ( .A(n1032), .ZN(n1207) );
NAND2_X1 U896 ( .A1(n1069), .A2(n1232), .ZN(n1032) );
XOR2_X1 U897 ( .A(KEYINPUT8), .B(n1070), .Z(n1232) );
INV_X1 U898 ( .A(n1231), .ZN(n1208) );
NAND3_X1 U899 ( .A1(n1056), .A2(n1227), .A3(n1233), .ZN(n1231) );
XOR2_X1 U900 ( .A(G128), .B(n1234), .Z(G30) );
NOR3_X1 U901 ( .A1(n1235), .A2(n1044), .A3(n1222), .ZN(n1234) );
NAND4_X1 U902 ( .A1(n1236), .A2(n1056), .A3(n1089), .A4(n1227), .ZN(n1222) );
INV_X1 U903 ( .A(n1203), .ZN(n1044) );
XNOR2_X1 U904 ( .A(KEYINPUT2), .B(n1067), .ZN(n1235) );
INV_X1 U905 ( .A(n1210), .ZN(n1067) );
XOR2_X1 U906 ( .A(n1122), .B(n1237), .Z(G3) );
NAND2_X1 U907 ( .A1(KEYINPUT39), .A2(G101), .ZN(n1237) );
OR2_X1 U908 ( .A1(n1046), .A2(n1193), .ZN(n1122) );
NAND2_X1 U909 ( .A1(n1064), .A2(n1233), .ZN(n1046) );
XOR2_X1 U910 ( .A(G125), .B(n1199), .Z(G27) );
AND4_X1 U911 ( .A1(n1238), .A2(n1194), .A3(n1239), .A4(n1072), .ZN(n1199) );
AND2_X1 U912 ( .A1(n1227), .A2(n1210), .ZN(n1239) );
NAND2_X1 U913 ( .A1(n1055), .A2(n1240), .ZN(n1227) );
NAND4_X1 U914 ( .A1(n1100), .A2(G902), .A3(n1241), .A4(n1097), .ZN(n1240) );
INV_X1 U915 ( .A(G900), .ZN(n1097) );
INV_X1 U916 ( .A(n1048), .ZN(n1238) );
XNOR2_X1 U917 ( .A(G122), .B(n1211), .ZN(G24) );
NAND4_X1 U918 ( .A1(n1242), .A2(n1065), .A3(n1223), .A4(n1224), .ZN(n1211) );
NOR2_X1 U919 ( .A1(n1089), .A2(n1236), .ZN(n1065) );
XNOR2_X1 U920 ( .A(G119), .B(n1243), .ZN(G21) );
NAND2_X1 U921 ( .A1(KEYINPUT42), .A2(n1244), .ZN(n1243) );
INV_X1 U922 ( .A(n1212), .ZN(n1244) );
NAND4_X1 U923 ( .A1(n1064), .A2(n1242), .A3(n1236), .A4(n1089), .ZN(n1212) );
INV_X1 U924 ( .A(n1245), .ZN(n1236) );
XNOR2_X1 U925 ( .A(n1213), .B(n1246), .ZN(G18) );
NOR2_X1 U926 ( .A1(KEYINPUT43), .A2(n1247), .ZN(n1246) );
INV_X1 U927 ( .A(G116), .ZN(n1247) );
NAND3_X1 U928 ( .A1(n1242), .A2(n1203), .A3(n1233), .ZN(n1213) );
NOR2_X1 U929 ( .A1(n1224), .A2(n1248), .ZN(n1203) );
XNOR2_X1 U930 ( .A(G113), .B(n1214), .ZN(G15) );
NAND3_X1 U931 ( .A1(n1194), .A2(n1242), .A3(n1233), .ZN(n1214) );
NOR2_X1 U932 ( .A1(n1245), .A2(n1089), .ZN(n1233) );
AND2_X1 U933 ( .A1(n1072), .A2(n1249), .ZN(n1242) );
NOR2_X1 U934 ( .A1(n1060), .A2(n1250), .ZN(n1072) );
INV_X1 U935 ( .A(n1251), .ZN(n1060) );
AND2_X1 U936 ( .A1(n1248), .A2(n1224), .ZN(n1194) );
NAND2_X1 U937 ( .A1(n1252), .A2(n1253), .ZN(G12) );
NAND2_X1 U938 ( .A1(n1123), .A2(n1254), .ZN(n1253) );
XOR2_X1 U939 ( .A(KEYINPUT4), .B(n1255), .Z(n1252) );
NOR2_X1 U940 ( .A1(n1123), .A2(n1254), .ZN(n1255) );
NOR3_X1 U941 ( .A1(n1047), .A2(n1193), .A3(n1048), .ZN(n1123) );
NAND2_X1 U942 ( .A1(n1245), .A2(n1089), .ZN(n1048) );
XOR2_X1 U943 ( .A(n1256), .B(n1140), .Z(n1089) );
NAND2_X1 U944 ( .A1(G217), .A2(n1257), .ZN(n1140) );
NAND2_X1 U945 ( .A1(n1138), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U946 ( .A(n1259), .B(n1260), .ZN(n1138) );
XNOR2_X1 U947 ( .A(G137), .B(n1261), .ZN(n1260) );
NAND2_X1 U948 ( .A1(KEYINPUT18), .A2(n1262), .ZN(n1261) );
XOR2_X1 U949 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U950 ( .A(G110), .B(n1265), .ZN(n1264) );
NOR2_X1 U951 ( .A1(KEYINPUT57), .A2(n1266), .ZN(n1265) );
XNOR2_X1 U952 ( .A(G119), .B(G128), .ZN(n1266) );
NAND2_X1 U953 ( .A1(n1267), .A2(n1268), .ZN(n1263) );
NAND2_X1 U954 ( .A1(n1104), .A2(G146), .ZN(n1268) );
XOR2_X1 U955 ( .A(KEYINPUT49), .B(n1269), .Z(n1267) );
NOR2_X1 U956 ( .A1(G146), .A2(n1104), .ZN(n1269) );
NAND2_X1 U957 ( .A1(G221), .A2(n1270), .ZN(n1259) );
XNOR2_X1 U958 ( .A(n1090), .B(n1271), .ZN(n1245) );
NOR2_X1 U959 ( .A1(G472), .A2(KEYINPUT26), .ZN(n1271) );
NAND2_X1 U960 ( .A1(n1272), .A2(n1258), .ZN(n1090) );
XOR2_X1 U961 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U962 ( .A(n1135), .B(n1275), .ZN(n1274) );
XNOR2_X1 U963 ( .A(n1171), .B(n1167), .ZN(n1275) );
AND3_X1 U964 ( .A1(n1276), .A2(n1062), .A3(G210), .ZN(n1171) );
INV_X1 U965 ( .A(n1166), .ZN(n1135) );
XOR2_X1 U966 ( .A(n1277), .B(n1278), .Z(n1273) );
NOR2_X1 U967 ( .A1(KEYINPUT27), .A2(n1168), .ZN(n1278) );
INV_X1 U968 ( .A(n1279), .ZN(n1168) );
XNOR2_X1 U969 ( .A(G101), .B(KEYINPUT15), .ZN(n1277) );
NAND2_X1 U970 ( .A1(n1249), .A2(n1056), .ZN(n1193) );
NOR2_X1 U971 ( .A1(n1250), .A2(n1251), .ZN(n1056) );
XOR2_X1 U972 ( .A(n1280), .B(G469), .Z(n1251) );
NAND2_X1 U973 ( .A1(n1281), .A2(n1258), .ZN(n1280) );
XOR2_X1 U974 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U975 ( .A(KEYINPUT7), .B(n1279), .ZN(n1283) );
NAND3_X1 U976 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1279) );
OR2_X1 U977 ( .A1(n1105), .A2(KEYINPUT62), .ZN(n1286) );
NAND4_X1 U978 ( .A1(n1105), .A2(n1287), .A3(KEYINPUT62), .A4(n1288), .ZN(n1285) );
NAND2_X1 U979 ( .A1(n1107), .A2(n1289), .ZN(n1284) );
NAND2_X1 U980 ( .A1(n1105), .A2(n1287), .ZN(n1289) );
INV_X1 U981 ( .A(KEYINPUT37), .ZN(n1287) );
XOR2_X1 U982 ( .A(G134), .B(G137), .Z(n1105) );
XOR2_X1 U983 ( .A(n1290), .B(n1185), .Z(n1282) );
XNOR2_X1 U984 ( .A(n1291), .B(n1292), .ZN(n1185) );
XNOR2_X1 U985 ( .A(n1254), .B(n1293), .ZN(n1292) );
NOR2_X1 U986 ( .A1(G953), .A2(n1096), .ZN(n1293) );
INV_X1 U987 ( .A(G227), .ZN(n1096) );
NAND2_X1 U988 ( .A1(n1294), .A2(n1295), .ZN(n1290) );
NAND2_X1 U989 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XNOR2_X1 U990 ( .A(KEYINPUT17), .B(n1183), .ZN(n1297) );
XNOR2_X1 U991 ( .A(KEYINPUT1), .B(n1167), .ZN(n1296) );
XOR2_X1 U992 ( .A(n1298), .B(KEYINPUT50), .Z(n1294) );
NAND2_X1 U993 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U994 ( .A(KEYINPUT17), .B(n1183), .Z(n1300) );
XNOR2_X1 U995 ( .A(n1301), .B(n1302), .ZN(n1183) );
XNOR2_X1 U996 ( .A(n1303), .B(n1304), .ZN(n1302) );
NOR2_X1 U997 ( .A1(KEYINPUT56), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U998 ( .A(G101), .B(KEYINPUT52), .ZN(n1305) );
NAND2_X1 U999 ( .A1(KEYINPUT36), .A2(n1306), .ZN(n1303) );
INV_X1 U1000 ( .A(G107), .ZN(n1306) );
XNOR2_X1 U1001 ( .A(KEYINPUT1), .B(n1103), .ZN(n1299) );
XOR2_X1 U1002 ( .A(n1059), .B(KEYINPUT47), .Z(n1250) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1257), .ZN(n1059) );
NAND2_X1 U1004 ( .A1(G234), .A2(n1258), .ZN(n1257) );
AND2_X1 U1005 ( .A1(n1210), .A2(n1307), .ZN(n1249) );
NAND2_X1 U1006 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND4_X1 U1007 ( .A1(n1100), .A2(G902), .A3(n1241), .A4(n1129), .ZN(n1309) );
INV_X1 U1008 ( .A(G898), .ZN(n1129) );
XNOR2_X1 U1009 ( .A(G953), .B(KEYINPUT30), .ZN(n1100) );
XOR2_X1 U1010 ( .A(n1055), .B(KEYINPUT61), .Z(n1308) );
NAND3_X1 U1011 ( .A1(n1241), .A2(n1062), .A3(G952), .ZN(n1055) );
NAND2_X1 U1012 ( .A1(G237), .A2(G234), .ZN(n1241) );
NOR2_X1 U1013 ( .A1(n1069), .A2(n1070), .ZN(n1210) );
AND2_X1 U1014 ( .A1(G214), .A2(n1310), .ZN(n1070) );
NOR2_X1 U1015 ( .A1(n1311), .A2(n1079), .ZN(n1069) );
NOR2_X1 U1016 ( .A1(n1189), .A2(n1312), .ZN(n1079) );
AND2_X1 U1017 ( .A1(n1313), .A2(n1258), .ZN(n1312) );
XNOR2_X1 U1018 ( .A(KEYINPUT11), .B(n1080), .ZN(n1311) );
AND3_X1 U1019 ( .A1(n1189), .A2(n1258), .A3(n1313), .ZN(n1080) );
XNOR2_X1 U1020 ( .A(n1219), .B(n1218), .ZN(n1313) );
AND2_X1 U1021 ( .A1(n1314), .A2(n1315), .ZN(n1218) );
NAND3_X1 U1022 ( .A1(G224), .A2(n1062), .A3(n1316), .ZN(n1315) );
XNOR2_X1 U1023 ( .A(G125), .B(n1103), .ZN(n1316) );
NAND2_X1 U1024 ( .A1(n1317), .A2(n1318), .ZN(n1314) );
NAND2_X1 U1025 ( .A1(G224), .A2(n1062), .ZN(n1318) );
XNOR2_X1 U1026 ( .A(G125), .B(n1167), .ZN(n1317) );
INV_X1 U1027 ( .A(n1103), .ZN(n1167) );
XNOR2_X1 U1028 ( .A(G146), .B(n1319), .ZN(n1103) );
NAND2_X1 U1029 ( .A1(n1320), .A2(n1321), .ZN(n1219) );
NAND2_X1 U1030 ( .A1(n1134), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1031 ( .A(n1323), .B(KEYINPUT33), .Z(n1320) );
OR2_X1 U1032 ( .A1(n1322), .A2(n1134), .ZN(n1323) );
AND2_X1 U1033 ( .A1(n1324), .A2(n1325), .ZN(n1134) );
NAND2_X1 U1034 ( .A1(G122), .A2(n1254), .ZN(n1325) );
INV_X1 U1035 ( .A(G110), .ZN(n1254) );
XOR2_X1 U1036 ( .A(n1326), .B(KEYINPUT16), .Z(n1324) );
NAND2_X1 U1037 ( .A1(G110), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1038 ( .A(n1166), .B(n1131), .Z(n1322) );
XNOR2_X1 U1039 ( .A(n1328), .B(n1301), .ZN(n1131) );
XNOR2_X1 U1040 ( .A(G107), .B(G101), .ZN(n1328) );
XOR2_X1 U1041 ( .A(G113), .B(n1329), .Z(n1166) );
XNOR2_X1 U1042 ( .A(n1330), .B(G116), .ZN(n1329) );
INV_X1 U1043 ( .A(G119), .ZN(n1330) );
NAND2_X1 U1044 ( .A1(G210), .A2(n1310), .ZN(n1189) );
NAND2_X1 U1045 ( .A1(n1276), .A2(n1258), .ZN(n1310) );
INV_X1 U1046 ( .A(n1064), .ZN(n1047) );
NOR2_X1 U1047 ( .A1(n1224), .A2(n1223), .ZN(n1064) );
INV_X1 U1048 ( .A(n1248), .ZN(n1223) );
XOR2_X1 U1049 ( .A(G478), .B(n1331), .Z(n1248) );
NOR2_X1 U1050 ( .A1(n1088), .A2(KEYINPUT45), .ZN(n1331) );
AND2_X1 U1051 ( .A1(n1332), .A2(n1258), .ZN(n1088) );
XOR2_X1 U1052 ( .A(KEYINPUT20), .B(n1143), .Z(n1332) );
AND2_X1 U1053 ( .A1(n1333), .A2(n1334), .ZN(n1143) );
NAND3_X1 U1054 ( .A1(n1270), .A2(n1335), .A3(G217), .ZN(n1334) );
XOR2_X1 U1055 ( .A(n1336), .B(n1337), .Z(n1335) );
NAND2_X1 U1056 ( .A1(n1338), .A2(n1339), .ZN(n1333) );
NAND2_X1 U1057 ( .A1(G217), .A2(n1270), .ZN(n1339) );
AND2_X1 U1058 ( .A1(n1340), .A2(n1062), .ZN(n1270) );
XOR2_X1 U1059 ( .A(KEYINPUT5), .B(G234), .Z(n1340) );
XNOR2_X1 U1060 ( .A(n1337), .B(n1336), .ZN(n1338) );
XNOR2_X1 U1061 ( .A(n1319), .B(n1341), .ZN(n1336) );
NOR2_X1 U1062 ( .A1(G107), .A2(KEYINPUT35), .ZN(n1341) );
XNOR2_X1 U1063 ( .A(G128), .B(G143), .ZN(n1319) );
XOR2_X1 U1064 ( .A(G116), .B(n1342), .Z(n1337) );
XNOR2_X1 U1065 ( .A(G134), .B(n1327), .ZN(n1342) );
NAND2_X1 U1066 ( .A1(n1086), .A2(n1343), .ZN(n1224) );
NAND2_X1 U1067 ( .A1(G475), .A2(n1083), .ZN(n1343) );
OR2_X1 U1068 ( .A1(n1083), .A2(G475), .ZN(n1086) );
NAND2_X1 U1069 ( .A1(n1146), .A2(n1258), .ZN(n1083) );
INV_X1 U1070 ( .A(G902), .ZN(n1258) );
XNOR2_X1 U1071 ( .A(n1344), .B(n1345), .ZN(n1146) );
XNOR2_X1 U1072 ( .A(n1346), .B(n1347), .ZN(n1345) );
XNOR2_X1 U1073 ( .A(G146), .B(n1327), .ZN(n1347) );
INV_X1 U1074 ( .A(G122), .ZN(n1327) );
INV_X1 U1075 ( .A(G113), .ZN(n1346) );
XNOR2_X1 U1076 ( .A(n1348), .B(n1104), .ZN(n1344) );
XOR2_X1 U1077 ( .A(G125), .B(n1291), .Z(n1104) );
XNOR2_X1 U1078 ( .A(G140), .B(KEYINPUT58), .ZN(n1291) );
XOR2_X1 U1079 ( .A(n1349), .B(n1301), .Z(n1348) );
XOR2_X1 U1080 ( .A(G104), .B(KEYINPUT31), .Z(n1301) );
NAND3_X1 U1081 ( .A1(n1350), .A2(n1351), .A3(KEYINPUT40), .ZN(n1349) );
NAND2_X1 U1082 ( .A1(n1107), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1083 ( .A(KEYINPUT54), .B(n1353), .Z(n1350) );
NOR2_X1 U1084 ( .A1(n1107), .A2(n1352), .ZN(n1353) );
NAND2_X1 U1085 ( .A1(n1354), .A2(n1355), .ZN(n1352) );
NAND2_X1 U1086 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1087 ( .A(n1358), .B(KEYINPUT29), .Z(n1354) );
OR2_X1 U1088 ( .A1(n1357), .A2(n1356), .ZN(n1358) );
NAND3_X1 U1089 ( .A1(n1276), .A2(n1062), .A3(G214), .ZN(n1356) );
INV_X1 U1090 ( .A(G953), .ZN(n1062) );
INV_X1 U1091 ( .A(G237), .ZN(n1276) );
INV_X1 U1092 ( .A(G143), .ZN(n1357) );
INV_X1 U1093 ( .A(n1288), .ZN(n1107) );
XOR2_X1 U1094 ( .A(G131), .B(KEYINPUT28), .Z(n1288) );
endmodule


