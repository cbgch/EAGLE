//Key = 1110110100111110110001110011001010100010000100001110010011100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317;

XNOR2_X1 U723 ( .A(G107), .B(n1001), .ZN(G9) );
NAND2_X1 U724 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U725 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR4_X1 U726 ( .A1(n1006), .A2(n1007), .A3(G953), .A4(n1008), .ZN(n1005) );
NOR3_X1 U727 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1007) );
NOR2_X1 U728 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U729 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR2_X1 U731 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NOR2_X1 U732 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U733 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U734 ( .A1(n1024), .A2(n1025), .ZN(n1016) );
NOR2_X1 U735 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U736 ( .A1(KEYINPUT9), .A2(n1028), .ZN(n1026) );
NOR3_X1 U737 ( .A1(n1025), .A2(n1029), .A3(n1019), .ZN(n1012) );
INV_X1 U738 ( .A(n1030), .ZN(n1019) );
NOR2_X1 U739 ( .A1(n1002), .A2(n1031), .ZN(n1029) );
NAND2_X1 U740 ( .A1(n1032), .A2(n1033), .ZN(n1006) );
NAND2_X1 U741 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U742 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U743 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND3_X1 U745 ( .A1(n1043), .A2(n1030), .A3(n1044), .ZN(n1042) );
NAND2_X1 U746 ( .A1(n1045), .A2(n1009), .ZN(n1038) );
NAND3_X1 U747 ( .A1(n1046), .A2(n1047), .A3(KEYINPUT9), .ZN(n1045) );
XOR2_X1 U748 ( .A(n1048), .B(KEYINPUT54), .Z(n1036) );
NAND3_X1 U749 ( .A1(n1049), .A2(n1030), .A3(n1041), .ZN(n1048) );
INV_X1 U750 ( .A(n1009), .ZN(n1041) );
NAND2_X1 U751 ( .A1(KEYINPUT10), .A2(n1050), .ZN(n1009) );
INV_X1 U752 ( .A(n1051), .ZN(n1032) );
NOR3_X1 U753 ( .A1(n1008), .A2(G953), .A3(G952), .ZN(n1004) );
AND4_X1 U754 ( .A1(n1052), .A2(n1053), .A3(n1034), .A4(n1054), .ZN(n1008) );
INV_X1 U755 ( .A(n1025), .ZN(n1034) );
XOR2_X1 U756 ( .A(n1055), .B(KEYINPUT11), .Z(n1053) );
NAND4_X1 U757 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
XNOR2_X1 U758 ( .A(KEYINPUT22), .B(n1060), .ZN(n1059) );
XOR2_X1 U759 ( .A(n1061), .B(G478), .Z(n1056) );
XOR2_X1 U760 ( .A(n1062), .B(G469), .Z(n1052) );
XOR2_X1 U761 ( .A(n1063), .B(n1064), .Z(G72) );
XOR2_X1 U762 ( .A(n1065), .B(n1066), .Z(n1064) );
NOR2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U764 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
INV_X1 U765 ( .A(G900), .ZN(n1070) );
XNOR2_X1 U766 ( .A(G227), .B(KEYINPUT35), .ZN(n1069) );
NOR3_X1 U767 ( .A1(n1071), .A2(KEYINPUT24), .A3(n1072), .ZN(n1065) );
XNOR2_X1 U768 ( .A(G953), .B(KEYINPUT5), .ZN(n1071) );
NOR2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1063) );
XOR2_X1 U770 ( .A(n1075), .B(n1076), .Z(n1074) );
XNOR2_X1 U771 ( .A(n1077), .B(n1078), .ZN(n1076) );
XNOR2_X1 U772 ( .A(KEYINPUT51), .B(n1079), .ZN(n1075) );
NOR2_X1 U773 ( .A1(KEYINPUT31), .A2(n1080), .ZN(n1079) );
XNOR2_X1 U774 ( .A(KEYINPUT62), .B(n1081), .ZN(n1080) );
NAND2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(G69) );
NAND2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NAND2_X1 U778 ( .A1(n1088), .A2(n1085), .ZN(n1087) );
NAND2_X1 U779 ( .A1(G953), .A2(n1089), .ZN(n1085) );
INV_X1 U780 ( .A(n1090), .ZN(n1088) );
INV_X1 U781 ( .A(n1084), .ZN(n1086) );
XNOR2_X1 U782 ( .A(n1091), .B(n1092), .ZN(n1084) );
NOR2_X1 U783 ( .A1(n1090), .A2(n1093), .ZN(n1092) );
XNOR2_X1 U784 ( .A(n1094), .B(n1095), .ZN(n1093) );
NAND3_X1 U785 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1094) );
NAND2_X1 U786 ( .A1(KEYINPUT20), .A2(n1099), .ZN(n1098) );
NAND3_X1 U787 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1097) );
INV_X1 U788 ( .A(KEYINPUT20), .ZN(n1101) );
OR2_X1 U789 ( .A1(n1102), .A2(n1100), .ZN(n1096) );
NOR2_X1 U790 ( .A1(KEYINPUT45), .A2(n1099), .ZN(n1100) );
NAND2_X1 U791 ( .A1(n1068), .A2(n1103), .ZN(n1091) );
NAND2_X1 U792 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XNOR2_X1 U793 ( .A(KEYINPUT53), .B(n1106), .ZN(n1105) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XOR2_X1 U795 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1107), .A2(n1113), .ZN(G63) );
XOR2_X1 U798 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U799 ( .A1(n1111), .A2(G478), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1107), .A2(n1116), .ZN(G60) );
XOR2_X1 U801 ( .A(n1117), .B(n1118), .Z(n1116) );
AND2_X1 U802 ( .A1(G475), .A2(n1111), .ZN(n1118) );
NOR2_X1 U803 ( .A1(KEYINPUT46), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U804 ( .A(G104), .B(n1106), .ZN(G6) );
NOR2_X1 U805 ( .A1(n1107), .A2(n1120), .ZN(G57) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U807 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U808 ( .A1(KEYINPUT56), .A2(n1125), .ZN(n1124) );
NAND2_X1 U809 ( .A1(n1111), .A2(G472), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1107), .A2(n1126), .ZN(G54) );
XOR2_X1 U811 ( .A(n1127), .B(n1128), .Z(n1126) );
XNOR2_X1 U812 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U813 ( .A1(KEYINPUT52), .A2(n1131), .ZN(n1130) );
NAND2_X1 U814 ( .A1(KEYINPUT32), .A2(n1132), .ZN(n1129) );
XNOR2_X1 U815 ( .A(n1133), .B(n1134), .ZN(n1132) );
XNOR2_X1 U816 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR2_X1 U817 ( .A1(KEYINPUT29), .A2(n1137), .ZN(n1136) );
XOR2_X1 U818 ( .A(n1138), .B(n1139), .Z(n1127) );
XNOR2_X1 U819 ( .A(n1140), .B(n1141), .ZN(n1139) );
NAND2_X1 U820 ( .A1(n1111), .A2(G469), .ZN(n1138) );
NOR2_X1 U821 ( .A1(n1107), .A2(n1142), .ZN(G51) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U823 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U824 ( .A(n1147), .B(KEYINPUT33), .Z(n1143) );
NAND2_X1 U825 ( .A1(n1111), .A2(n1148), .ZN(n1147) );
AND2_X1 U826 ( .A1(n1149), .A2(n1051), .ZN(n1111) );
NAND3_X1 U827 ( .A1(n1104), .A2(n1106), .A3(n1072), .ZN(n1051) );
AND4_X1 U828 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1072) );
NOR4_X1 U829 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U832 ( .A(n1162), .B(KEYINPUT40), .Z(n1160) );
NAND2_X1 U833 ( .A1(n1031), .A2(n1003), .ZN(n1106) );
AND4_X1 U834 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1104) );
NOR4_X1 U835 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR2_X1 U836 ( .A1(n1028), .A2(n1171), .ZN(n1170) );
NOR3_X1 U837 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1169) );
NOR2_X1 U838 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
INV_X1 U839 ( .A(KEYINPUT42), .ZN(n1176) );
AND3_X1 U840 ( .A1(n1049), .A2(n1177), .A3(n1161), .ZN(n1175) );
NOR3_X1 U841 ( .A1(n1043), .A2(n1044), .A3(n1015), .ZN(n1049) );
NOR2_X1 U842 ( .A1(KEYINPUT42), .A2(n1178), .ZN(n1173) );
INV_X1 U843 ( .A(n1027), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1179), .A2(n1180), .ZN(n1165) );
NOR2_X1 U845 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND4_X1 U846 ( .A1(n1183), .A2(n1046), .A3(n1040), .A4(n1184), .ZN(n1182) );
INV_X1 U847 ( .A(KEYINPUT36), .ZN(n1181) );
NOR2_X1 U848 ( .A1(KEYINPUT36), .A2(n1185), .ZN(n1179) );
NAND2_X1 U849 ( .A1(n1003), .A2(n1186), .ZN(n1163) );
XOR2_X1 U850 ( .A(KEYINPUT44), .B(n1002), .Z(n1186) );
AND2_X1 U851 ( .A1(n1030), .A2(n1187), .ZN(n1003) );
XNOR2_X1 U852 ( .A(KEYINPUT6), .B(n1188), .ZN(n1149) );
NOR2_X1 U853 ( .A1(n1068), .A2(G952), .ZN(n1107) );
XOR2_X1 U854 ( .A(G146), .B(n1158), .Z(G48) );
AND3_X1 U855 ( .A1(n1189), .A2(n1184), .A3(n1031), .ZN(n1158) );
XNOR2_X1 U856 ( .A(G143), .B(n1150), .ZN(G45) );
NAND4_X1 U857 ( .A1(n1190), .A2(n1191), .A3(n1021), .A4(n1192), .ZN(n1150) );
NOR2_X1 U858 ( .A1(n1193), .A2(n1028), .ZN(n1192) );
XNOR2_X1 U859 ( .A(G140), .B(n1151), .ZN(G42) );
NAND3_X1 U860 ( .A1(n1031), .A2(n1194), .A3(n1027), .ZN(n1151) );
XOR2_X1 U861 ( .A(G137), .B(n1157), .Z(G39) );
AND3_X1 U862 ( .A1(n1194), .A2(n1195), .A3(n1040), .ZN(n1157) );
XNOR2_X1 U863 ( .A(n1156), .B(n1196), .ZN(G36) );
NAND2_X1 U864 ( .A1(KEYINPUT14), .A2(G134), .ZN(n1196) );
AND3_X1 U865 ( .A1(n1194), .A2(n1002), .A3(n1047), .ZN(n1156) );
XNOR2_X1 U866 ( .A(G131), .B(n1197), .ZN(G33) );
NAND2_X1 U867 ( .A1(KEYINPUT30), .A2(n1155), .ZN(n1197) );
AND3_X1 U868 ( .A1(n1031), .A2(n1194), .A3(n1047), .ZN(n1155) );
NOR2_X1 U869 ( .A1(n1193), .A2(n1025), .ZN(n1194) );
NAND2_X1 U870 ( .A1(n1198), .A2(n1023), .ZN(n1025) );
INV_X1 U871 ( .A(n1022), .ZN(n1198) );
XOR2_X1 U872 ( .A(G128), .B(n1154), .Z(G30) );
AND3_X1 U873 ( .A1(n1184), .A2(n1002), .A3(n1189), .ZN(n1154) );
INV_X1 U874 ( .A(n1193), .ZN(n1189) );
NAND3_X1 U875 ( .A1(n1199), .A2(n1054), .A3(n1200), .ZN(n1193) );
AND2_X1 U876 ( .A1(n1195), .A2(n1021), .ZN(n1184) );
INV_X1 U877 ( .A(n1161), .ZN(n1021) );
XNOR2_X1 U878 ( .A(G101), .B(n1201), .ZN(G3) );
NAND2_X1 U879 ( .A1(n1178), .A2(n1202), .ZN(n1201) );
XNOR2_X1 U880 ( .A(KEYINPUT15), .B(n1028), .ZN(n1202) );
INV_X1 U881 ( .A(n1047), .ZN(n1028) );
XOR2_X1 U882 ( .A(G125), .B(n1203), .Z(G27) );
NOR2_X1 U883 ( .A1(n1161), .A2(n1162), .ZN(n1203) );
NAND4_X1 U884 ( .A1(n1046), .A2(n1027), .A3(n1031), .A4(n1200), .ZN(n1162) );
NAND2_X1 U885 ( .A1(n1204), .A2(n1205), .ZN(n1200) );
NAND3_X1 U886 ( .A1(G902), .A2(n1050), .A3(n1073), .ZN(n1205) );
NOR2_X1 U887 ( .A1(n1068), .A2(G900), .ZN(n1073) );
INV_X1 U888 ( .A(n1011), .ZN(n1046) );
XNOR2_X1 U889 ( .A(G122), .B(n1164), .ZN(G24) );
NAND4_X1 U890 ( .A1(n1206), .A2(n1030), .A3(n1190), .A4(n1191), .ZN(n1164) );
NOR2_X1 U891 ( .A1(n1207), .A2(n1208), .ZN(n1030) );
NAND2_X1 U892 ( .A1(n1209), .A2(n1210), .ZN(G21) );
NAND2_X1 U893 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U894 ( .A(KEYINPUT49), .B(n1213), .Z(n1209) );
NOR2_X1 U895 ( .A1(n1211), .A2(n1212), .ZN(n1213) );
INV_X1 U896 ( .A(G119), .ZN(n1212) );
INV_X1 U897 ( .A(n1185), .ZN(n1211) );
NAND3_X1 U898 ( .A1(n1040), .A2(n1195), .A3(n1206), .ZN(n1185) );
NOR2_X1 U899 ( .A1(n1214), .A2(n1057), .ZN(n1195) );
XOR2_X1 U900 ( .A(G116), .B(n1168), .Z(G18) );
AND3_X1 U901 ( .A1(n1047), .A2(n1002), .A3(n1206), .ZN(n1168) );
AND2_X1 U902 ( .A1(n1060), .A2(n1191), .ZN(n1002) );
XNOR2_X1 U903 ( .A(n1215), .B(n1167), .ZN(G15) );
AND3_X1 U904 ( .A1(n1047), .A2(n1031), .A3(n1206), .ZN(n1167) );
NOR3_X1 U905 ( .A1(n1161), .A2(n1183), .A3(n1011), .ZN(n1206) );
NAND2_X1 U906 ( .A1(n1216), .A2(n1054), .ZN(n1011) );
XNOR2_X1 U907 ( .A(KEYINPUT18), .B(n1199), .ZN(n1216) );
AND2_X1 U908 ( .A1(n1217), .A2(n1190), .ZN(n1031) );
NOR2_X1 U909 ( .A1(n1208), .A2(n1057), .ZN(n1047) );
INV_X1 U910 ( .A(n1207), .ZN(n1057) );
INV_X1 U911 ( .A(n1214), .ZN(n1208) );
XNOR2_X1 U912 ( .A(G110), .B(n1218), .ZN(G12) );
NAND2_X1 U913 ( .A1(n1178), .A2(n1027), .ZN(n1218) );
NOR2_X1 U914 ( .A1(n1214), .A2(n1207), .ZN(n1027) );
XNOR2_X1 U915 ( .A(n1219), .B(G472), .ZN(n1207) );
NAND2_X1 U916 ( .A1(n1220), .A2(n1188), .ZN(n1219) );
XNOR2_X1 U917 ( .A(n1121), .B(n1125), .ZN(n1220) );
XNOR2_X1 U918 ( .A(n1221), .B(n1222), .ZN(n1125) );
XNOR2_X1 U919 ( .A(G113), .B(n1223), .ZN(n1222) );
NAND2_X1 U920 ( .A1(KEYINPUT43), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U921 ( .A(n1225), .B(n1081), .ZN(n1221) );
XOR2_X1 U922 ( .A(n1226), .B(G101), .Z(n1121) );
NAND2_X1 U923 ( .A1(G210), .A2(n1227), .ZN(n1226) );
XNOR2_X1 U924 ( .A(n1058), .B(KEYINPUT57), .ZN(n1214) );
XOR2_X1 U925 ( .A(n1228), .B(n1112), .Z(n1058) );
AND2_X1 U926 ( .A1(G217), .A2(n1229), .ZN(n1112) );
NAND2_X1 U927 ( .A1(n1110), .A2(n1188), .ZN(n1228) );
XNOR2_X1 U928 ( .A(n1230), .B(n1231), .ZN(n1110) );
XOR2_X1 U929 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U930 ( .A(G110), .B(n1234), .ZN(n1233) );
NOR2_X1 U931 ( .A1(KEYINPUT19), .A2(n1235), .ZN(n1234) );
XNOR2_X1 U932 ( .A(G119), .B(G128), .ZN(n1235) );
NAND4_X1 U933 ( .A1(KEYINPUT16), .A2(G221), .A3(G234), .A4(n1068), .ZN(n1232) );
XNOR2_X1 U934 ( .A(n1236), .B(n1237), .ZN(n1230) );
NOR2_X1 U935 ( .A1(KEYINPUT3), .A2(n1238), .ZN(n1237) );
INV_X1 U936 ( .A(n1171), .ZN(n1178) );
NAND2_X1 U937 ( .A1(n1040), .A2(n1187), .ZN(n1171) );
NOR4_X1 U938 ( .A1(n1161), .A2(n1183), .A3(n1043), .A4(n1044), .ZN(n1187) );
INV_X1 U939 ( .A(n1054), .ZN(n1044) );
NAND2_X1 U940 ( .A1(G221), .A2(n1229), .ZN(n1054) );
NAND2_X1 U941 ( .A1(G234), .A2(n1188), .ZN(n1229) );
INV_X1 U942 ( .A(n1199), .ZN(n1043) );
NAND2_X1 U943 ( .A1(n1239), .A2(n1240), .ZN(n1199) );
NAND2_X1 U944 ( .A1(G469), .A2(n1062), .ZN(n1240) );
XOR2_X1 U945 ( .A(KEYINPUT12), .B(n1241), .Z(n1239) );
NOR2_X1 U946 ( .A1(G469), .A2(n1062), .ZN(n1241) );
NAND2_X1 U947 ( .A1(n1242), .A2(n1188), .ZN(n1062) );
XOR2_X1 U948 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U949 ( .A(n1245), .B(n1081), .ZN(n1244) );
INV_X1 U950 ( .A(n1133), .ZN(n1081) );
XOR2_X1 U951 ( .A(n1246), .B(n1247), .Z(n1133) );
INV_X1 U952 ( .A(n1236), .ZN(n1247) );
XOR2_X1 U953 ( .A(G137), .B(KEYINPUT25), .Z(n1236) );
XNOR2_X1 U954 ( .A(G131), .B(G134), .ZN(n1246) );
NOR2_X1 U955 ( .A1(n1248), .A2(n1249), .ZN(n1245) );
XOR2_X1 U956 ( .A(n1250), .B(KEYINPUT26), .Z(n1249) );
NAND2_X1 U957 ( .A1(n1251), .A2(n1141), .ZN(n1250) );
XNOR2_X1 U958 ( .A(n1252), .B(KEYINPUT27), .ZN(n1251) );
NOR2_X1 U959 ( .A1(n1141), .A2(n1252), .ZN(n1248) );
XNOR2_X1 U960 ( .A(n1253), .B(n1254), .ZN(n1252) );
XNOR2_X1 U961 ( .A(KEYINPUT55), .B(n1140), .ZN(n1254) );
INV_X1 U962 ( .A(G110), .ZN(n1140) );
NAND2_X1 U963 ( .A1(KEYINPUT34), .A2(n1255), .ZN(n1253) );
AND2_X1 U964 ( .A1(G227), .A2(n1068), .ZN(n1141) );
NOR2_X1 U965 ( .A1(n1256), .A2(n1257), .ZN(n1243) );
AND2_X1 U966 ( .A1(n1137), .A2(n1077), .ZN(n1257) );
NOR2_X1 U967 ( .A1(n1258), .A2(n1137), .ZN(n1256) );
XNOR2_X1 U968 ( .A(n1259), .B(G101), .ZN(n1137) );
NAND2_X1 U969 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND2_X1 U970 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
INV_X1 U971 ( .A(KEYINPUT28), .ZN(n1263) );
NAND3_X1 U972 ( .A1(n1264), .A2(n1265), .A3(KEYINPUT28), .ZN(n1260) );
INV_X1 U973 ( .A(G107), .ZN(n1265) );
XNOR2_X1 U974 ( .A(KEYINPUT17), .B(n1077), .ZN(n1258) );
INV_X1 U975 ( .A(n1135), .ZN(n1077) );
XNOR2_X1 U976 ( .A(n1266), .B(G128), .ZN(n1135) );
NAND2_X1 U977 ( .A1(n1267), .A2(KEYINPUT4), .ZN(n1266) );
XOR2_X1 U978 ( .A(n1268), .B(G146), .Z(n1267) );
NAND2_X1 U979 ( .A1(KEYINPUT50), .A2(n1269), .ZN(n1268) );
INV_X1 U980 ( .A(n1177), .ZN(n1183) );
NAND2_X1 U981 ( .A1(n1204), .A2(n1270), .ZN(n1177) );
NAND3_X1 U982 ( .A1(G902), .A2(n1050), .A3(n1090), .ZN(n1270) );
NOR2_X1 U983 ( .A1(G898), .A2(n1068), .ZN(n1090) );
NAND3_X1 U984 ( .A1(n1050), .A2(n1068), .A3(G952), .ZN(n1204) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1050) );
NAND2_X1 U986 ( .A1(n1022), .A2(n1023), .ZN(n1161) );
NAND2_X1 U987 ( .A1(G214), .A2(n1271), .ZN(n1023) );
XNOR2_X1 U988 ( .A(n1272), .B(n1148), .ZN(n1022) );
AND2_X1 U989 ( .A1(G210), .A2(n1271), .ZN(n1148) );
NAND2_X1 U990 ( .A1(n1273), .A2(n1188), .ZN(n1271) );
INV_X1 U991 ( .A(G237), .ZN(n1273) );
NAND3_X1 U992 ( .A1(n1274), .A2(n1188), .A3(n1275), .ZN(n1272) );
XOR2_X1 U993 ( .A(KEYINPUT13), .B(n1276), .Z(n1275) );
NOR2_X1 U994 ( .A1(n1146), .A2(n1145), .ZN(n1276) );
NAND2_X1 U995 ( .A1(n1146), .A2(n1145), .ZN(n1274) );
XNOR2_X1 U996 ( .A(n1225), .B(n1277), .ZN(n1145) );
XOR2_X1 U997 ( .A(G125), .B(n1278), .Z(n1277) );
NOR2_X1 U998 ( .A1(n1089), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U999 ( .A(KEYINPUT39), .B(n1068), .ZN(n1279) );
INV_X1 U1000 ( .A(G224), .ZN(n1089) );
XOR2_X1 U1001 ( .A(n1280), .B(n1281), .Z(n1225) );
XNOR2_X1 U1002 ( .A(G143), .B(n1282), .ZN(n1281) );
NAND2_X1 U1003 ( .A1(KEYINPUT1), .A2(G146), .ZN(n1282) );
NAND2_X1 U1004 ( .A1(KEYINPUT7), .A2(G128), .ZN(n1280) );
XNOR2_X1 U1005 ( .A(n1102), .B(n1283), .ZN(n1146) );
XNOR2_X1 U1006 ( .A(n1284), .B(n1099), .ZN(n1283) );
XNOR2_X1 U1007 ( .A(n1215), .B(n1224), .ZN(n1099) );
XOR2_X1 U1008 ( .A(G116), .B(G119), .Z(n1224) );
INV_X1 U1009 ( .A(n1095), .ZN(n1284) );
XOR2_X1 U1010 ( .A(G110), .B(n1285), .Z(n1095) );
NOR2_X1 U1011 ( .A1(KEYINPUT60), .A2(n1286), .ZN(n1285) );
XNOR2_X1 U1012 ( .A(n1262), .B(G101), .ZN(n1102) );
XNOR2_X1 U1013 ( .A(G107), .B(n1264), .ZN(n1262) );
INV_X1 U1014 ( .A(n1015), .ZN(n1040) );
NAND2_X1 U1015 ( .A1(n1217), .A2(n1060), .ZN(n1015) );
INV_X1 U1016 ( .A(n1190), .ZN(n1060) );
XNOR2_X1 U1017 ( .A(n1287), .B(G475), .ZN(n1190) );
NAND2_X1 U1018 ( .A1(n1288), .A2(n1119), .ZN(n1287) );
XOR2_X1 U1019 ( .A(n1289), .B(n1290), .Z(n1119) );
XOR2_X1 U1020 ( .A(n1238), .B(n1291), .Z(n1290) );
XOR2_X1 U1021 ( .A(n1286), .B(n1292), .Z(n1291) );
NOR2_X1 U1022 ( .A1(KEYINPUT59), .A2(n1264), .ZN(n1292) );
XNOR2_X1 U1023 ( .A(G104), .B(KEYINPUT38), .ZN(n1264) );
XNOR2_X1 U1024 ( .A(n1078), .B(G146), .ZN(n1238) );
XNOR2_X1 U1025 ( .A(G125), .B(n1255), .ZN(n1078) );
INV_X1 U1026 ( .A(n1131), .ZN(n1255) );
XOR2_X1 U1027 ( .A(G140), .B(KEYINPUT37), .Z(n1131) );
XOR2_X1 U1028 ( .A(n1293), .B(n1294), .Z(n1289) );
XOR2_X1 U1029 ( .A(KEYINPUT58), .B(KEYINPUT41), .Z(n1294) );
XNOR2_X1 U1030 ( .A(n1295), .B(n1215), .ZN(n1293) );
INV_X1 U1031 ( .A(G113), .ZN(n1215) );
NAND2_X1 U1032 ( .A1(n1296), .A2(KEYINPUT2), .ZN(n1295) );
XOR2_X1 U1033 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1034 ( .A(G131), .B(n1299), .Z(n1298) );
AND3_X1 U1035 ( .A1(G214), .A2(n1300), .A3(n1227), .ZN(n1299) );
NOR2_X1 U1036 ( .A1(G953), .A2(G237), .ZN(n1227) );
INV_X1 U1037 ( .A(KEYINPUT47), .ZN(n1300) );
XNOR2_X1 U1038 ( .A(G143), .B(KEYINPUT48), .ZN(n1297) );
XNOR2_X1 U1039 ( .A(G902), .B(KEYINPUT61), .ZN(n1288) );
XOR2_X1 U1040 ( .A(n1191), .B(KEYINPUT0), .Z(n1217) );
NAND3_X1 U1041 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1191) );
NAND2_X1 U1042 ( .A1(KEYINPUT63), .A2(G478), .ZN(n1303) );
OR3_X1 U1043 ( .A1(G478), .A2(KEYINPUT63), .A3(n1061), .ZN(n1302) );
NAND2_X1 U1044 ( .A1(n1304), .A2(n1061), .ZN(n1301) );
NAND2_X1 U1045 ( .A1(n1188), .A2(n1115), .ZN(n1061) );
NAND2_X1 U1046 ( .A1(n1305), .A2(n1306), .ZN(n1115) );
NAND4_X1 U1047 ( .A1(G217), .A2(n1307), .A3(n1308), .A4(n1068), .ZN(n1306) );
XNOR2_X1 U1048 ( .A(n1309), .B(n1310), .ZN(n1307) );
INV_X1 U1049 ( .A(n1311), .ZN(n1310) );
NAND2_X1 U1050 ( .A1(n1312), .A2(n1313), .ZN(n1305) );
NAND3_X1 U1051 ( .A1(n1308), .A2(n1068), .A3(G217), .ZN(n1313) );
INV_X1 U1052 ( .A(G953), .ZN(n1068) );
XOR2_X1 U1053 ( .A(G234), .B(KEYINPUT8), .Z(n1308) );
XNOR2_X1 U1054 ( .A(n1311), .B(n1309), .ZN(n1312) );
XOR2_X1 U1055 ( .A(n1314), .B(n1286), .Z(n1309) );
XNOR2_X1 U1056 ( .A(G122), .B(KEYINPUT23), .ZN(n1286) );
XNOR2_X1 U1057 ( .A(G116), .B(G107), .ZN(n1314) );
XOR2_X1 U1058 ( .A(G128), .B(n1315), .Z(n1311) );
XNOR2_X1 U1059 ( .A(n1269), .B(G134), .ZN(n1315) );
INV_X1 U1060 ( .A(G143), .ZN(n1269) );
INV_X1 U1061 ( .A(G902), .ZN(n1188) );
NAND2_X1 U1062 ( .A1(n1316), .A2(n1317), .ZN(n1304) );
INV_X1 U1063 ( .A(KEYINPUT63), .ZN(n1317) );
XOR2_X1 U1064 ( .A(KEYINPUT21), .B(G478), .Z(n1316) );
endmodule


