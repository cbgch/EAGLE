//Key = 1001011001101101101110000000000111010011000110010111100010111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327;

XNOR2_X1 U727 ( .A(G107), .B(n1011), .ZN(G9) );
NOR2_X1 U728 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR3_X1 U729 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NAND3_X1 U730 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1014) );
NAND2_X1 U731 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U732 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND3_X1 U733 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NAND2_X1 U734 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NAND2_X1 U735 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND3_X1 U736 ( .A1(n1031), .A2(n1032), .A3(n1030), .ZN(n1022) );
NAND2_X1 U737 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NAND2_X1 U738 ( .A1(n1026), .A2(n1035), .ZN(n1034) );
OR2_X1 U739 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U740 ( .A1(n1024), .A2(n1038), .ZN(n1033) );
NAND2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U742 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U743 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U744 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U745 ( .A1(n1047), .A2(n1048), .ZN(n1039) );
NAND2_X1 U746 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
INV_X1 U748 ( .A(n1053), .ZN(n1049) );
INV_X1 U749 ( .A(n1054), .ZN(n1020) );
NOR3_X1 U750 ( .A1(n1055), .A2(G953), .A3(n1056), .ZN(n1012) );
INV_X1 U751 ( .A(n1017), .ZN(n1056) );
NAND4_X1 U752 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1017) );
NOR4_X1 U753 ( .A1(n1045), .A2(n1029), .A3(n1061), .A4(n1062), .ZN(n1060) );
XNOR2_X1 U754 ( .A(G472), .B(n1063), .ZN(n1062) );
NOR2_X1 U755 ( .A1(n1064), .A2(KEYINPUT54), .ZN(n1063) );
XNOR2_X1 U756 ( .A(n1065), .B(KEYINPUT18), .ZN(n1061) );
NOR2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1059) );
XNOR2_X1 U758 ( .A(n1068), .B(n1069), .ZN(n1066) );
NAND2_X1 U759 ( .A1(KEYINPUT44), .A2(n1070), .ZN(n1068) );
XOR2_X1 U760 ( .A(n1071), .B(G469), .Z(n1058) );
XNOR2_X1 U761 ( .A(n1072), .B(n1073), .ZN(n1057) );
XNOR2_X1 U762 ( .A(KEYINPUT48), .B(n1015), .ZN(n1055) );
XOR2_X1 U763 ( .A(n1074), .B(n1075), .Z(G72) );
NOR3_X1 U764 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NOR2_X1 U765 ( .A1(G900), .A2(n1018), .ZN(n1078) );
NOR2_X1 U766 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
XOR2_X1 U767 ( .A(n1081), .B(KEYINPUT9), .Z(n1076) );
NAND2_X1 U768 ( .A1(n1080), .A2(n1079), .ZN(n1081) );
XOR2_X1 U769 ( .A(n1082), .B(n1083), .Z(n1079) );
XOR2_X1 U770 ( .A(G131), .B(n1084), .Z(n1083) );
XNOR2_X1 U771 ( .A(G140), .B(G125), .ZN(n1080) );
NAND2_X1 U772 ( .A1(n1085), .A2(n1086), .ZN(n1074) );
NAND2_X1 U773 ( .A1(n1087), .A2(n1018), .ZN(n1086) );
NAND2_X1 U774 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U775 ( .A(KEYINPUT56), .B(n1090), .ZN(n1089) );
NAND2_X1 U776 ( .A1(G953), .A2(n1091), .ZN(n1085) );
NAND2_X1 U777 ( .A1(G900), .A2(n1092), .ZN(n1091) );
XNOR2_X1 U778 ( .A(KEYINPUT23), .B(n1093), .ZN(n1092) );
XOR2_X1 U779 ( .A(n1094), .B(n1095), .Z(G69) );
XOR2_X1 U780 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XNOR2_X1 U783 ( .A(G953), .B(KEYINPUT13), .ZN(n1100) );
XNOR2_X1 U784 ( .A(n1102), .B(n1103), .ZN(n1098) );
NAND2_X1 U785 ( .A1(n1104), .A2(n1105), .ZN(n1096) );
NAND2_X1 U786 ( .A1(n1106), .A2(G224), .ZN(n1105) );
XNOR2_X1 U787 ( .A(G898), .B(KEYINPUT59), .ZN(n1106) );
XNOR2_X1 U788 ( .A(KEYINPUT37), .B(n1018), .ZN(n1104) );
NOR3_X1 U789 ( .A1(n1107), .A2(KEYINPUT36), .A3(G953), .ZN(n1094) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(G66) );
NOR3_X1 U791 ( .A1(n1072), .A2(n1110), .A3(n1111), .ZN(n1109) );
NOR3_X1 U792 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
INV_X1 U793 ( .A(n1115), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1116), .A2(n1115), .ZN(n1110) );
AND2_X1 U795 ( .A1(n1016), .A2(n1073), .ZN(n1116) );
NOR2_X1 U796 ( .A1(n1108), .A2(n1117), .ZN(G63) );
NOR3_X1 U797 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1117) );
AND2_X1 U798 ( .A1(n1121), .A2(KEYINPUT28), .ZN(n1120) );
NOR3_X1 U799 ( .A1(KEYINPUT28), .A2(n1122), .A3(n1121), .ZN(n1119) );
NOR3_X1 U800 ( .A1(n1114), .A2(KEYINPUT1), .A3(n1123), .ZN(n1122) );
NOR3_X1 U801 ( .A1(n1114), .A2(n1124), .A3(n1123), .ZN(n1118) );
NOR2_X1 U802 ( .A1(n1125), .A2(KEYINPUT28), .ZN(n1124) );
NOR2_X1 U803 ( .A1(KEYINPUT1), .A2(n1126), .ZN(n1125) );
NOR2_X1 U804 ( .A1(n1108), .A2(n1127), .ZN(G60) );
XOR2_X1 U805 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U806 ( .A1(n1130), .A2(n1114), .ZN(n1128) );
XNOR2_X1 U807 ( .A(G104), .B(n1131), .ZN(G6) );
NAND2_X1 U808 ( .A1(KEYINPUT0), .A2(n1132), .ZN(n1131) );
INV_X1 U809 ( .A(n1133), .ZN(n1132) );
NOR2_X1 U810 ( .A1(n1108), .A2(n1134), .ZN(G57) );
XOR2_X1 U811 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U813 ( .A(KEYINPUT46), .B(n1139), .Z(n1138) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
INV_X1 U815 ( .A(n1142), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1143), .A2(n1114), .ZN(n1140) );
NOR3_X1 U817 ( .A1(n1142), .A2(n1143), .A3(n1114), .ZN(n1137) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(n1142) );
NOR2_X1 U819 ( .A1(n1146), .A2(KEYINPUT21), .ZN(n1145) );
XNOR2_X1 U820 ( .A(n1147), .B(G101), .ZN(n1135) );
NOR3_X1 U821 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(G54) );
AND2_X1 U822 ( .A1(KEYINPUT35), .A2(n1108), .ZN(n1150) );
NOR3_X1 U823 ( .A1(KEYINPUT35), .A2(n1018), .A3(n1015), .ZN(n1149) );
INV_X1 U824 ( .A(G952), .ZN(n1015) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1148) );
XNOR2_X1 U826 ( .A(n1153), .B(n1154), .ZN(n1152) );
XNOR2_X1 U827 ( .A(n1155), .B(n1156), .ZN(n1151) );
NAND3_X1 U828 ( .A1(G469), .A2(n1157), .A3(G902), .ZN(n1155) );
XNOR2_X1 U829 ( .A(KEYINPUT63), .B(n1016), .ZN(n1157) );
NOR2_X1 U830 ( .A1(n1108), .A2(n1158), .ZN(G51) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U832 ( .A1(n1070), .A2(n1114), .ZN(n1160) );
NAND2_X1 U833 ( .A1(G902), .A2(n1016), .ZN(n1114) );
NAND3_X1 U834 ( .A1(n1107), .A2(n1090), .A3(n1088), .ZN(n1016) );
AND4_X1 U835 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1088) );
NOR4_X1 U836 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NAND2_X1 U837 ( .A1(n1169), .A2(n1170), .ZN(n1163) );
AND4_X1 U838 ( .A1(n1171), .A2(n1133), .A3(n1172), .A4(n1173), .ZN(n1107) );
AND4_X1 U839 ( .A1(n1174), .A2(n1175), .A3(n1011), .A4(n1176), .ZN(n1173) );
NAND3_X1 U840 ( .A1(n1037), .A2(n1041), .A3(n1177), .ZN(n1011) );
NAND2_X1 U841 ( .A1(KEYINPUT19), .A2(n1178), .ZN(n1172) );
NAND3_X1 U842 ( .A1(n1177), .A2(n1041), .A3(n1036), .ZN(n1133) );
NAND2_X1 U843 ( .A1(n1179), .A2(n1180), .ZN(n1171) );
NAND3_X1 U844 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
XNOR2_X1 U845 ( .A(KEYINPUT49), .B(n1184), .ZN(n1183) );
NAND4_X1 U846 ( .A1(n1185), .A2(n1065), .A3(n1026), .A4(n1186), .ZN(n1182) );
AND2_X1 U847 ( .A1(n1047), .A2(n1041), .ZN(n1026) );
NAND4_X1 U848 ( .A1(n1187), .A2(n1188), .A3(n1047), .A4(n1189), .ZN(n1181) );
INV_X1 U849 ( .A(KEYINPUT19), .ZN(n1188) );
NAND2_X1 U850 ( .A1(KEYINPUT10), .A2(n1190), .ZN(n1159) );
XOR2_X1 U851 ( .A(n1191), .B(n1192), .Z(n1190) );
XNOR2_X1 U852 ( .A(n1193), .B(n1194), .ZN(n1192) );
NOR2_X1 U853 ( .A1(KEYINPUT61), .A2(n1195), .ZN(n1194) );
NOR2_X1 U854 ( .A1(n1018), .A2(G952), .ZN(n1108) );
XNOR2_X1 U855 ( .A(G146), .B(n1196), .ZN(G48) );
NAND2_X1 U856 ( .A1(KEYINPUT15), .A2(n1168), .ZN(n1196) );
AND2_X1 U857 ( .A1(n1036), .A2(n1197), .ZN(n1168) );
NAND3_X1 U858 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(G45) );
OR2_X1 U859 ( .A1(n1161), .A2(KEYINPUT58), .ZN(n1200) );
NAND3_X1 U860 ( .A1(KEYINPUT58), .A2(n1161), .A3(G143), .ZN(n1199) );
NAND2_X1 U861 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
NAND2_X1 U862 ( .A1(KEYINPUT58), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U863 ( .A(KEYINPUT3), .B(n1161), .ZN(n1203) );
NAND4_X1 U864 ( .A1(n1204), .A2(n1179), .A3(n1053), .A4(n1205), .ZN(n1161) );
NOR3_X1 U865 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
XNOR2_X1 U866 ( .A(G140), .B(n1209), .ZN(G42) );
NAND4_X1 U867 ( .A1(n1030), .A2(n1169), .A3(n1210), .A4(n1211), .ZN(n1209) );
XNOR2_X1 U868 ( .A(KEYINPUT2), .B(n1043), .ZN(n1211) );
NOR2_X1 U869 ( .A1(n1029), .A2(n1207), .ZN(n1210) );
XNOR2_X1 U870 ( .A(G137), .B(n1212), .ZN(G39) );
NAND2_X1 U871 ( .A1(KEYINPUT60), .A2(n1167), .ZN(n1212) );
AND2_X1 U872 ( .A1(n1187), .A2(n1170), .ZN(n1167) );
XNOR2_X1 U873 ( .A(G134), .B(n1162), .ZN(G36) );
NAND3_X1 U874 ( .A1(n1170), .A2(n1037), .A3(n1053), .ZN(n1162) );
XOR2_X1 U875 ( .A(G131), .B(n1166), .Z(G33) );
AND3_X1 U876 ( .A1(n1053), .A2(n1170), .A3(n1036), .ZN(n1166) );
AND4_X1 U877 ( .A1(n1030), .A2(n1204), .A3(n1213), .A4(n1032), .ZN(n1170) );
XNOR2_X1 U878 ( .A(n1165), .B(n1214), .ZN(G30) );
NAND2_X1 U879 ( .A1(KEYINPUT12), .A2(G128), .ZN(n1214) );
AND2_X1 U880 ( .A1(n1197), .A2(n1037), .ZN(n1165) );
AND4_X1 U881 ( .A1(n1215), .A2(n1051), .A3(n1216), .A4(n1204), .ZN(n1197) );
NOR2_X1 U882 ( .A1(n1207), .A2(n1027), .ZN(n1216) );
INV_X1 U883 ( .A(n1213), .ZN(n1207) );
XNOR2_X1 U884 ( .A(G101), .B(n1175), .ZN(G3) );
NAND3_X1 U885 ( .A1(n1053), .A2(n1177), .A3(n1024), .ZN(n1175) );
XNOR2_X1 U886 ( .A(G125), .B(n1090), .ZN(G27) );
NAND4_X1 U887 ( .A1(n1047), .A2(n1169), .A3(n1179), .A4(n1213), .ZN(n1090) );
NAND2_X1 U888 ( .A1(n1054), .A2(n1217), .ZN(n1213) );
NAND4_X1 U889 ( .A1(G902), .A2(G953), .A3(n1218), .A4(n1219), .ZN(n1217) );
INV_X1 U890 ( .A(G900), .ZN(n1219) );
AND3_X1 U891 ( .A1(n1051), .A2(n1052), .A3(n1036), .ZN(n1169) );
XNOR2_X1 U892 ( .A(G122), .B(n1220), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1221), .A2(n1222), .A3(n1185), .A4(n1065), .ZN(n1220) );
XNOR2_X1 U894 ( .A(n1041), .B(KEYINPUT39), .ZN(n1221) );
NOR2_X1 U895 ( .A1(n1215), .A2(n1051), .ZN(n1041) );
XOR2_X1 U896 ( .A(G119), .B(n1178), .Z(G21) );
AND2_X1 U897 ( .A1(n1222), .A2(n1187), .ZN(n1178) );
AND3_X1 U898 ( .A1(n1215), .A2(n1051), .A3(n1024), .ZN(n1187) );
INV_X1 U899 ( .A(n1052), .ZN(n1215) );
XNOR2_X1 U900 ( .A(G116), .B(n1223), .ZN(G18) );
NOR2_X1 U901 ( .A1(n1224), .A2(KEYINPUT62), .ZN(n1223) );
NOR2_X1 U902 ( .A1(n1027), .A2(n1184), .ZN(n1224) );
NAND4_X1 U903 ( .A1(n1047), .A2(n1053), .A3(n1037), .A4(n1186), .ZN(n1184) );
NOR2_X1 U904 ( .A1(n1065), .A2(n1206), .ZN(n1037) );
INV_X1 U905 ( .A(n1185), .ZN(n1206) );
XNOR2_X1 U906 ( .A(G113), .B(n1174), .ZN(G15) );
NAND3_X1 U907 ( .A1(n1036), .A2(n1053), .A3(n1222), .ZN(n1174) );
AND3_X1 U908 ( .A1(n1179), .A2(n1186), .A3(n1047), .ZN(n1222) );
AND2_X1 U909 ( .A1(n1046), .A2(n1225), .ZN(n1047) );
NOR2_X1 U910 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
NOR2_X1 U911 ( .A1(n1185), .A2(n1208), .ZN(n1036) );
INV_X1 U912 ( .A(n1065), .ZN(n1208) );
XNOR2_X1 U913 ( .A(n1226), .B(n1227), .ZN(G12) );
NOR2_X1 U914 ( .A1(KEYINPUT34), .A2(n1176), .ZN(n1227) );
NAND4_X1 U915 ( .A1(n1051), .A2(n1024), .A3(n1177), .A4(n1052), .ZN(n1176) );
XOR2_X1 U916 ( .A(n1064), .B(n1228), .Z(n1052) );
NOR2_X1 U917 ( .A1(KEYINPUT11), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U918 ( .A(KEYINPUT8), .B(n1143), .ZN(n1229) );
INV_X1 U919 ( .A(G472), .ZN(n1143) );
AND2_X1 U920 ( .A1(n1230), .A2(n1231), .ZN(n1064) );
XOR2_X1 U921 ( .A(n1232), .B(n1233), .Z(n1230) );
XNOR2_X1 U922 ( .A(n1234), .B(n1235), .ZN(n1233) );
INV_X1 U923 ( .A(n1144), .ZN(n1235) );
XOR2_X1 U924 ( .A(n1236), .B(n1195), .Z(n1144) );
XNOR2_X1 U925 ( .A(G113), .B(n1237), .ZN(n1236) );
NOR2_X1 U926 ( .A1(n1147), .A2(KEYINPUT30), .ZN(n1234) );
AND3_X1 U927 ( .A1(n1238), .A2(n1018), .A3(G210), .ZN(n1147) );
XNOR2_X1 U928 ( .A(n1146), .B(G101), .ZN(n1232) );
NOR3_X1 U929 ( .A1(n1027), .A2(n1189), .A3(n1043), .ZN(n1177) );
INV_X1 U930 ( .A(n1204), .ZN(n1043) );
NOR2_X1 U931 ( .A1(n1046), .A2(n1045), .ZN(n1204) );
INV_X1 U932 ( .A(n1225), .ZN(n1045) );
NAND2_X1 U933 ( .A1(G221), .A2(n1239), .ZN(n1225) );
XNOR2_X1 U934 ( .A(n1071), .B(n1240), .ZN(n1046) );
NOR2_X1 U935 ( .A1(KEYINPUT55), .A2(n1241), .ZN(n1240) );
XOR2_X1 U936 ( .A(KEYINPUT57), .B(G469), .Z(n1241) );
NAND2_X1 U937 ( .A1(n1242), .A2(n1231), .ZN(n1071) );
XOR2_X1 U938 ( .A(n1243), .B(n1154), .Z(n1242) );
XNOR2_X1 U939 ( .A(n1082), .B(n1244), .ZN(n1154) );
XNOR2_X1 U940 ( .A(n1146), .B(n1245), .ZN(n1244) );
NAND3_X1 U941 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1245) );
NAND2_X1 U942 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
OR3_X1 U943 ( .A1(n1250), .A2(n1249), .A3(n1251), .ZN(n1247) );
INV_X1 U944 ( .A(KEYINPUT16), .ZN(n1250) );
NAND2_X1 U945 ( .A1(n1251), .A2(n1252), .ZN(n1246) );
NAND2_X1 U946 ( .A1(KEYINPUT16), .A2(n1253), .ZN(n1252) );
XNOR2_X1 U947 ( .A(KEYINPUT40), .B(n1249), .ZN(n1253) );
XOR2_X1 U948 ( .A(n1254), .B(KEYINPUT53), .Z(n1249) );
XOR2_X1 U949 ( .A(G101), .B(KEYINPUT6), .Z(n1251) );
AND2_X1 U950 ( .A1(n1255), .A2(n1256), .ZN(n1146) );
NAND2_X1 U951 ( .A1(G131), .A2(n1084), .ZN(n1256) );
XOR2_X1 U952 ( .A(KEYINPUT31), .B(n1257), .Z(n1255) );
NOR2_X1 U953 ( .A1(G131), .A2(n1084), .ZN(n1257) );
XOR2_X1 U954 ( .A(G134), .B(G137), .Z(n1084) );
XOR2_X1 U955 ( .A(n1258), .B(n1259), .Z(n1082) );
NOR2_X1 U956 ( .A1(KEYINPUT25), .A2(n1260), .ZN(n1259) );
NOR2_X1 U957 ( .A1(n1261), .A2(n1262), .ZN(n1243) );
NOR3_X1 U958 ( .A1(n1153), .A2(KEYINPUT22), .A3(n1156), .ZN(n1262) );
NAND2_X1 U959 ( .A1(G227), .A2(n1018), .ZN(n1156) );
NOR2_X1 U960 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
INV_X1 U961 ( .A(n1153), .ZN(n1264) );
XOR2_X1 U962 ( .A(G110), .B(G140), .Z(n1153) );
NOR2_X1 U963 ( .A1(KEYINPUT22), .A2(n1093), .ZN(n1263) );
INV_X1 U964 ( .A(G227), .ZN(n1093) );
INV_X1 U965 ( .A(n1186), .ZN(n1189) );
NAND2_X1 U966 ( .A1(n1054), .A2(n1265), .ZN(n1186) );
NAND4_X1 U967 ( .A1(G902), .A2(G953), .A3(n1218), .A4(n1101), .ZN(n1265) );
INV_X1 U968 ( .A(G898), .ZN(n1101) );
NAND3_X1 U969 ( .A1(n1218), .A2(n1018), .A3(n1266), .ZN(n1054) );
XNOR2_X1 U970 ( .A(G952), .B(KEYINPUT33), .ZN(n1266) );
NAND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n1218) );
INV_X1 U972 ( .A(n1179), .ZN(n1027) );
NOR2_X1 U973 ( .A1(n1030), .A2(n1029), .ZN(n1179) );
INV_X1 U974 ( .A(n1032), .ZN(n1029) );
NAND2_X1 U975 ( .A1(G214), .A2(n1267), .ZN(n1032) );
XNOR2_X1 U976 ( .A(n1069), .B(n1070), .ZN(n1030) );
NAND2_X1 U977 ( .A1(G210), .A2(n1267), .ZN(n1070) );
NAND2_X1 U978 ( .A1(n1238), .A2(n1231), .ZN(n1267) );
NAND2_X1 U979 ( .A1(n1268), .A2(n1231), .ZN(n1069) );
XOR2_X1 U980 ( .A(n1269), .B(n1191), .Z(n1268) );
XNOR2_X1 U981 ( .A(n1102), .B(n1270), .ZN(n1191) );
XNOR2_X1 U982 ( .A(n1271), .B(n1272), .ZN(n1270) );
NOR2_X1 U983 ( .A1(KEYINPUT7), .A2(n1103), .ZN(n1272) );
XOR2_X1 U984 ( .A(G113), .B(n1273), .Z(n1103) );
NOR2_X1 U985 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
AND3_X1 U986 ( .A1(KEYINPUT4), .A2(n1276), .A3(G116), .ZN(n1275) );
NOR2_X1 U987 ( .A1(KEYINPUT4), .A2(n1237), .ZN(n1274) );
XNOR2_X1 U988 ( .A(G116), .B(n1276), .ZN(n1237) );
XOR2_X1 U989 ( .A(n1277), .B(n1278), .Z(n1102) );
XNOR2_X1 U990 ( .A(n1226), .B(n1279), .ZN(n1278) );
XNOR2_X1 U991 ( .A(KEYINPUT50), .B(n1280), .ZN(n1279) );
XNOR2_X1 U992 ( .A(n1254), .B(n1281), .ZN(n1277) );
INV_X1 U993 ( .A(G101), .ZN(n1281) );
XNOR2_X1 U994 ( .A(G107), .B(n1282), .ZN(n1254) );
XNOR2_X1 U995 ( .A(n1283), .B(n1195), .ZN(n1269) );
XOR2_X1 U996 ( .A(n1258), .B(n1260), .Z(n1195) );
XNOR2_X1 U997 ( .A(G146), .B(G143), .ZN(n1258) );
NAND2_X1 U998 ( .A1(KEYINPUT47), .A2(n1193), .ZN(n1283) );
NAND2_X1 U999 ( .A1(n1284), .A2(G224), .ZN(n1193) );
XNOR2_X1 U1000 ( .A(G953), .B(KEYINPUT24), .ZN(n1284) );
NOR2_X1 U1001 ( .A1(n1185), .A2(n1065), .ZN(n1024) );
XOR2_X1 U1002 ( .A(n1285), .B(n1130), .Z(n1065) );
INV_X1 U1003 ( .A(G475), .ZN(n1130) );
OR2_X1 U1004 ( .A1(n1129), .A2(G902), .ZN(n1285) );
XNOR2_X1 U1005 ( .A(n1286), .B(n1287), .ZN(n1129) );
XOR2_X1 U1006 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U1007 ( .A(n1280), .B(G113), .ZN(n1289) );
INV_X1 U1008 ( .A(G122), .ZN(n1280) );
XNOR2_X1 U1009 ( .A(KEYINPUT43), .B(n1271), .ZN(n1288) );
INV_X1 U1010 ( .A(G125), .ZN(n1271) );
XNOR2_X1 U1011 ( .A(n1282), .B(n1290), .ZN(n1286) );
XOR2_X1 U1012 ( .A(n1291), .B(n1292), .Z(n1290) );
NOR2_X1 U1013 ( .A1(KEYINPUT45), .A2(n1293), .ZN(n1291) );
XOR2_X1 U1014 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U1015 ( .A(G131), .B(n1296), .Z(n1295) );
AND3_X1 U1016 ( .A1(G214), .A2(n1018), .A3(n1238), .ZN(n1296) );
INV_X1 U1017 ( .A(G237), .ZN(n1238) );
NAND2_X1 U1018 ( .A1(KEYINPUT38), .A2(G143), .ZN(n1294) );
XOR2_X1 U1019 ( .A(G104), .B(KEYINPUT17), .Z(n1282) );
XOR2_X1 U1020 ( .A(n1067), .B(KEYINPUT27), .Z(n1185) );
XOR2_X1 U1021 ( .A(n1297), .B(n1123), .Z(n1067) );
INV_X1 U1022 ( .A(G478), .ZN(n1123) );
NAND2_X1 U1023 ( .A1(n1126), .A2(n1231), .ZN(n1297) );
INV_X1 U1024 ( .A(n1121), .ZN(n1126) );
XNOR2_X1 U1025 ( .A(n1298), .B(n1299), .ZN(n1121) );
XOR2_X1 U1026 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U1027 ( .A(n1302), .B(n1303), .Z(n1301) );
NAND2_X1 U1028 ( .A1(KEYINPUT32), .A2(G116), .ZN(n1303) );
NAND2_X1 U1029 ( .A1(n1304), .A2(n1305), .ZN(n1302) );
NAND2_X1 U1030 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1031 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U1032 ( .A1(n1202), .A2(n1310), .ZN(n1309) );
INV_X1 U1033 ( .A(G143), .ZN(n1202) );
INV_X1 U1034 ( .A(n1260), .ZN(n1306) );
NAND2_X1 U1035 ( .A1(G143), .A2(n1311), .ZN(n1304) );
NAND2_X1 U1036 ( .A1(n1310), .A2(n1312), .ZN(n1311) );
NAND2_X1 U1037 ( .A1(n1260), .A2(n1308), .ZN(n1312) );
INV_X1 U1038 ( .A(KEYINPUT29), .ZN(n1308) );
INV_X1 U1039 ( .A(KEYINPUT42), .ZN(n1310) );
AND2_X1 U1040 ( .A1(n1313), .A2(G217), .ZN(n1300) );
XOR2_X1 U1041 ( .A(n1314), .B(n1315), .Z(n1298) );
XOR2_X1 U1042 ( .A(KEYINPUT51), .B(G134), .Z(n1315) );
XNOR2_X1 U1043 ( .A(G107), .B(G122), .ZN(n1314) );
XNOR2_X1 U1044 ( .A(n1072), .B(n1316), .ZN(n1051) );
NOR2_X1 U1045 ( .A1(n1073), .A2(KEYINPUT41), .ZN(n1316) );
INV_X1 U1046 ( .A(n1113), .ZN(n1073) );
NAND2_X1 U1047 ( .A1(G217), .A2(n1239), .ZN(n1113) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1231), .ZN(n1239) );
INV_X1 U1049 ( .A(G902), .ZN(n1231) );
NOR2_X1 U1050 ( .A1(n1115), .A2(G902), .ZN(n1072) );
XNOR2_X1 U1051 ( .A(n1317), .B(n1318), .ZN(n1115) );
XNOR2_X1 U1052 ( .A(n1319), .B(n1292), .ZN(n1318) );
XOR2_X1 U1053 ( .A(G146), .B(G140), .Z(n1292) );
NAND3_X1 U1054 ( .A1(n1313), .A2(G221), .A3(KEYINPUT52), .ZN(n1319) );
AND2_X1 U1055 ( .A1(G234), .A2(n1018), .ZN(n1313) );
INV_X1 U1056 ( .A(G953), .ZN(n1018) );
XOR2_X1 U1057 ( .A(n1320), .B(n1321), .Z(n1317) );
XNOR2_X1 U1058 ( .A(G137), .B(n1322), .ZN(n1321) );
NAND2_X1 U1059 ( .A1(n1323), .A2(KEYINPUT20), .ZN(n1322) );
XNOR2_X1 U1060 ( .A(G125), .B(KEYINPUT26), .ZN(n1323) );
NAND2_X1 U1061 ( .A1(n1324), .A2(n1325), .ZN(n1320) );
NAND2_X1 U1062 ( .A1(G110), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1063 ( .A(KEYINPUT5), .B(n1327), .Z(n1324) );
NOR2_X1 U1064 ( .A1(G110), .A2(n1326), .ZN(n1327) );
XNOR2_X1 U1065 ( .A(n1276), .B(n1260), .ZN(n1326) );
XOR2_X1 U1066 ( .A(G128), .B(KEYINPUT14), .Z(n1260) );
INV_X1 U1067 ( .A(G119), .ZN(n1276) );
INV_X1 U1068 ( .A(G110), .ZN(n1226) );
endmodule


