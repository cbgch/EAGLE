//Key = 1001110011111000110000111101000101111110011001000110101011001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296;

XNOR2_X1 U721 ( .A(G107), .B(n986), .ZN(G9) );
NOR2_X1 U722 ( .A1(n987), .A2(n988), .ZN(G75) );
XOR2_X1 U723 ( .A(n989), .B(KEYINPUT50), .Z(n988) );
NAND4_X1 U724 ( .A1(n990), .A2(G952), .A3(n991), .A4(n992), .ZN(n989) );
NOR4_X1 U725 ( .A1(G953), .A2(n993), .A3(n994), .A4(n995), .ZN(n992) );
NOR2_X1 U726 ( .A1(n996), .A2(n997), .ZN(n995) );
INV_X1 U727 ( .A(KEYINPUT29), .ZN(n997) );
NOR3_X1 U728 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n996) );
NOR2_X1 U729 ( .A1(n1001), .A2(n998), .ZN(n994) );
NOR2_X1 U730 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U731 ( .A1(n1004), .A2(n1000), .ZN(n1003) );
NOR2_X1 U732 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U733 ( .A1(KEYINPUT29), .A2(n999), .ZN(n1006) );
AND2_X1 U734 ( .A1(n1007), .A2(n1008), .ZN(n999) );
NAND3_X1 U735 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
NAND3_X1 U736 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1007) );
NAND2_X1 U737 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NAND3_X1 U738 ( .A1(n1017), .A2(n1018), .A3(n1010), .ZN(n1012) );
NAND3_X1 U739 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND3_X1 U740 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1017) );
NOR2_X1 U741 ( .A1(n1015), .A2(n1025), .ZN(n1005) );
NOR2_X1 U742 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
XOR2_X1 U746 ( .A(KEYINPUT42), .B(n1034), .Z(n1033) );
NOR3_X1 U747 ( .A1(n1019), .A2(n1020), .A3(n1035), .ZN(n1030) );
NOR2_X1 U748 ( .A1(n1036), .A2(n1016), .ZN(n1026) );
NOR3_X1 U749 ( .A1(n1016), .A2(n1037), .A3(n1029), .ZN(n1002) );
INV_X1 U750 ( .A(n1014), .ZN(n1029) );
INV_X1 U751 ( .A(n1011), .ZN(n1016) );
NOR2_X1 U752 ( .A1(n1035), .A2(n1032), .ZN(n1011) );
INV_X1 U753 ( .A(n1023), .ZN(n1032) );
NOR3_X1 U754 ( .A1(n1038), .A2(G953), .A3(n993), .ZN(n987) );
AND4_X1 U755 ( .A1(n1014), .A2(n1021), .A3(n1039), .A4(n1040), .ZN(n993) );
NOR4_X1 U756 ( .A1(n1041), .A2(n1015), .A3(n1042), .A4(n1043), .ZN(n1040) );
NOR2_X1 U757 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
XNOR2_X1 U758 ( .A(n1046), .B(KEYINPUT46), .ZN(n1045) );
INV_X1 U759 ( .A(n1047), .ZN(n1044) );
XNOR2_X1 U760 ( .A(n1048), .B(G469), .ZN(n1039) );
XOR2_X1 U761 ( .A(KEYINPUT14), .B(G952), .Z(n1038) );
XOR2_X1 U762 ( .A(n1049), .B(n1050), .Z(G72) );
XOR2_X1 U763 ( .A(n1051), .B(n1052), .Z(n1050) );
NOR2_X1 U764 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
XOR2_X1 U765 ( .A(KEYINPUT40), .B(n1055), .Z(n1054) );
NOR2_X1 U766 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U767 ( .A1(n1058), .A2(n1059), .ZN(n1051) );
NAND2_X1 U768 ( .A1(n1060), .A2(n1057), .ZN(n1059) );
XOR2_X1 U769 ( .A(n1061), .B(n1062), .Z(n1058) );
XOR2_X1 U770 ( .A(n1063), .B(n1064), .Z(n1062) );
NAND2_X1 U771 ( .A1(KEYINPUT25), .A2(n1065), .ZN(n1063) );
XOR2_X1 U772 ( .A(n1066), .B(n1067), .Z(n1061) );
XNOR2_X1 U773 ( .A(G134), .B(n1068), .ZN(n1067) );
NOR2_X1 U774 ( .A1(KEYINPUT15), .A2(n1069), .ZN(n1068) );
INV_X1 U775 ( .A(G137), .ZN(n1069) );
NAND2_X1 U776 ( .A1(KEYINPUT31), .A2(G131), .ZN(n1066) );
NAND2_X1 U777 ( .A1(n1053), .A2(n1070), .ZN(n1049) );
XOR2_X1 U778 ( .A(n1071), .B(n1072), .Z(G69) );
NOR2_X1 U779 ( .A1(n1073), .A2(n1053), .ZN(n1072) );
AND2_X1 U780 ( .A1(G224), .A2(G898), .ZN(n1073) );
NAND2_X1 U781 ( .A1(n1074), .A2(n1075), .ZN(n1071) );
NAND3_X1 U782 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
XOR2_X1 U783 ( .A(KEYINPUT36), .B(n1079), .Z(n1076) );
NAND2_X1 U784 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
NAND2_X1 U785 ( .A1(n1078), .A2(n1077), .ZN(n1080) );
INV_X1 U786 ( .A(n1081), .ZN(n1077) );
AND2_X1 U787 ( .A1(n1053), .A2(n1082), .ZN(n1079) );
NAND3_X1 U788 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NOR2_X1 U789 ( .A1(n1086), .A2(n1087), .ZN(G66) );
XOR2_X1 U790 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND3_X1 U791 ( .A1(n1046), .A2(G902), .A3(n1090), .ZN(n1088) );
XOR2_X1 U792 ( .A(n1091), .B(KEYINPUT28), .Z(n1090) );
NOR2_X1 U793 ( .A1(n1086), .A2(n1092), .ZN(G63) );
XNOR2_X1 U794 ( .A(n1093), .B(n1094), .ZN(n1092) );
AND2_X1 U795 ( .A1(G478), .A2(n1095), .ZN(n1093) );
NOR2_X1 U796 ( .A1(n1096), .A2(n1097), .ZN(G60) );
XOR2_X1 U797 ( .A(n1098), .B(n1099), .Z(n1097) );
AND2_X1 U798 ( .A1(G475), .A2(n1095), .ZN(n1099) );
NAND2_X1 U799 ( .A1(KEYINPUT60), .A2(n1100), .ZN(n1098) );
NOR2_X1 U800 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
XNOR2_X1 U801 ( .A(KEYINPUT11), .B(n1053), .ZN(n1102) );
XNOR2_X1 U802 ( .A(KEYINPUT45), .B(G952), .ZN(n1101) );
XNOR2_X1 U803 ( .A(G104), .B(n1084), .ZN(G6) );
NOR2_X1 U804 ( .A1(n1086), .A2(n1103), .ZN(G57) );
XOR2_X1 U805 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U806 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U807 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U808 ( .A(n1110), .B(n1111), .Z(n1104) );
XNOR2_X1 U809 ( .A(KEYINPUT32), .B(n1112), .ZN(n1111) );
NAND3_X1 U810 ( .A1(n1095), .A2(G472), .A3(KEYINPUT16), .ZN(n1110) );
INV_X1 U811 ( .A(n1113), .ZN(n1095) );
NOR2_X1 U812 ( .A1(n1086), .A2(n1114), .ZN(G54) );
XOR2_X1 U813 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U814 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U815 ( .A1(n1119), .A2(n1113), .ZN(n1118) );
NOR2_X1 U816 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
XOR2_X1 U817 ( .A(n1122), .B(KEYINPUT56), .Z(n1121) );
NAND2_X1 U818 ( .A1(n1123), .A2(n1109), .ZN(n1122) );
NOR2_X1 U819 ( .A1(n1123), .A2(n1109), .ZN(n1120) );
XNOR2_X1 U820 ( .A(n1124), .B(n1125), .ZN(n1123) );
XNOR2_X1 U821 ( .A(n1126), .B(KEYINPUT43), .ZN(n1125) );
NAND2_X1 U822 ( .A1(KEYINPUT9), .A2(n1127), .ZN(n1126) );
NOR2_X1 U823 ( .A1(n1086), .A2(n1128), .ZN(G51) );
XNOR2_X1 U824 ( .A(n1078), .B(n1129), .ZN(n1128) );
XOR2_X1 U825 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U826 ( .A1(n1132), .A2(n1113), .ZN(n1131) );
NAND2_X1 U827 ( .A1(G902), .A2(n1091), .ZN(n1113) );
NAND2_X1 U828 ( .A1(n1133), .A2(n990), .ZN(n1091) );
AND3_X1 U829 ( .A1(n1134), .A2(n1083), .A3(n1085), .ZN(n990) );
AND4_X1 U830 ( .A1(n1135), .A2(n986), .A3(n1136), .A4(n1137), .ZN(n1085) );
AND3_X1 U831 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
NAND3_X1 U832 ( .A1(n1023), .A2(n1141), .A3(n1009), .ZN(n986) );
NAND4_X1 U833 ( .A1(n1142), .A2(n1143), .A3(n1014), .A4(n1034), .ZN(n1083) );
XOR2_X1 U834 ( .A(n1144), .B(KEYINPUT63), .Z(n1142) );
XNOR2_X1 U835 ( .A(KEYINPUT3), .B(n1084), .ZN(n1134) );
NAND3_X1 U836 ( .A1(n1023), .A2(n1141), .A3(n1145), .ZN(n1084) );
XNOR2_X1 U837 ( .A(n991), .B(KEYINPUT62), .ZN(n1133) );
INV_X1 U838 ( .A(n1070), .ZN(n991) );
NAND4_X1 U839 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1070) );
AND4_X1 U840 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1149) );
NAND2_X1 U841 ( .A1(n1154), .A2(n1155), .ZN(n1148) );
NAND2_X1 U842 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U843 ( .A1(n1021), .A2(n1158), .ZN(n1157) );
NAND3_X1 U844 ( .A1(n1009), .A2(n1159), .A3(n1160), .ZN(n1146) );
XOR2_X1 U845 ( .A(KEYINPUT1), .B(n1034), .Z(n1159) );
NOR2_X1 U846 ( .A1(n1161), .A2(n1162), .ZN(n1130) );
XOR2_X1 U847 ( .A(KEYINPUT55), .B(n1163), .Z(n1162) );
NOR2_X1 U848 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
AND2_X1 U849 ( .A1(n1165), .A2(n1164), .ZN(n1161) );
XNOR2_X1 U850 ( .A(n1166), .B(KEYINPUT6), .ZN(n1165) );
AND2_X1 U851 ( .A1(G953), .A2(n1167), .ZN(n1086) );
XOR2_X1 U852 ( .A(KEYINPUT45), .B(G952), .Z(n1167) );
XNOR2_X1 U853 ( .A(G146), .B(n1147), .ZN(G48) );
NAND2_X1 U854 ( .A1(n1168), .A2(n1145), .ZN(n1147) );
XNOR2_X1 U855 ( .A(G143), .B(n1153), .ZN(G45) );
OR2_X1 U856 ( .A1(n1169), .A2(n1170), .ZN(n1153) );
XNOR2_X1 U857 ( .A(G140), .B(n1171), .ZN(G42) );
NAND3_X1 U858 ( .A1(n1021), .A2(n1172), .A3(n1154), .ZN(n1171) );
INV_X1 U859 ( .A(n1173), .ZN(n1154) );
XNOR2_X1 U860 ( .A(KEYINPUT53), .B(n1037), .ZN(n1172) );
XNOR2_X1 U861 ( .A(G137), .B(n1152), .ZN(G39) );
NAND3_X1 U862 ( .A1(n1014), .A2(n1021), .A3(n1160), .ZN(n1152) );
XNOR2_X1 U863 ( .A(G134), .B(n1151), .ZN(G36) );
NAND3_X1 U864 ( .A1(n1021), .A2(n1009), .A3(n1174), .ZN(n1151) );
XOR2_X1 U865 ( .A(n1150), .B(n1175), .Z(G33) );
XNOR2_X1 U866 ( .A(KEYINPUT22), .B(n1176), .ZN(n1175) );
NAND3_X1 U867 ( .A1(n1174), .A2(n1021), .A3(n1145), .ZN(n1150) );
INV_X1 U868 ( .A(n1035), .ZN(n1021) );
NAND2_X1 U869 ( .A1(n1022), .A2(n1177), .ZN(n1035) );
INV_X1 U870 ( .A(n1170), .ZN(n1174) );
NAND2_X1 U871 ( .A1(n1143), .A2(n1178), .ZN(n1170) );
XNOR2_X1 U872 ( .A(G128), .B(n1179), .ZN(G30) );
NAND2_X1 U873 ( .A1(n1168), .A2(n1009), .ZN(n1179) );
AND2_X1 U874 ( .A1(n1160), .A2(n1034), .ZN(n1168) );
NOR4_X1 U875 ( .A1(n1019), .A2(n1037), .A3(n1180), .A4(n1181), .ZN(n1160) );
NAND2_X1 U876 ( .A1(n1182), .A2(n1183), .ZN(G3) );
NAND2_X1 U877 ( .A1(n1184), .A2(n1112), .ZN(n1183) );
XOR2_X1 U878 ( .A(KEYINPUT27), .B(n1185), .Z(n1182) );
NOR2_X1 U879 ( .A1(n1184), .A2(n1112), .ZN(n1185) );
AND4_X1 U880 ( .A1(n1143), .A2(n1014), .A3(n1034), .A4(n1144), .ZN(n1184) );
NOR3_X1 U881 ( .A1(n1037), .A2(n1020), .A3(n1019), .ZN(n1143) );
INV_X1 U882 ( .A(n1158), .ZN(n1037) );
XNOR2_X1 U883 ( .A(G125), .B(n1186), .ZN(G27) );
NAND3_X1 U884 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
NAND2_X1 U885 ( .A1(KEYINPUT12), .A2(n1173), .ZN(n1188) );
NAND2_X1 U886 ( .A1(n1190), .A2(n1178), .ZN(n1173) );
NAND2_X1 U887 ( .A1(n1191), .A2(n1192), .ZN(n1187) );
INV_X1 U888 ( .A(KEYINPUT12), .ZN(n1192) );
NAND2_X1 U889 ( .A1(n1180), .A2(n1190), .ZN(n1191) );
NOR3_X1 U890 ( .A1(n1193), .A2(n1181), .A3(n1036), .ZN(n1190) );
INV_X1 U891 ( .A(n1178), .ZN(n1180) );
NAND2_X1 U892 ( .A1(n998), .A2(n1194), .ZN(n1178) );
NAND4_X1 U893 ( .A1(n1060), .A2(G902), .A3(n1195), .A4(n1057), .ZN(n1194) );
INV_X1 U894 ( .A(G900), .ZN(n1057) );
XNOR2_X1 U895 ( .A(G122), .B(n1138), .ZN(G24) );
NAND4_X1 U896 ( .A1(n1144), .A2(n1010), .A3(n1023), .A4(n1196), .ZN(n1138) );
NOR2_X1 U897 ( .A1(n1169), .A2(n1000), .ZN(n1196) );
INV_X1 U898 ( .A(n1197), .ZN(n1000) );
NAND3_X1 U899 ( .A1(n1198), .A2(n1199), .A3(n1034), .ZN(n1169) );
NOR2_X1 U900 ( .A1(n1020), .A2(n1193), .ZN(n1023) );
XOR2_X1 U901 ( .A(n1140), .B(n1200), .Z(G21) );
XOR2_X1 U902 ( .A(KEYINPUT34), .B(G119), .Z(n1200) );
NAND3_X1 U903 ( .A1(n1014), .A2(n1020), .A3(n1201), .ZN(n1140) );
XNOR2_X1 U904 ( .A(G116), .B(n1202), .ZN(G18) );
NAND2_X1 U905 ( .A1(KEYINPUT4), .A2(n1203), .ZN(n1202) );
INV_X1 U906 ( .A(n1139), .ZN(n1203) );
NAND3_X1 U907 ( .A1(n1009), .A2(n1181), .A3(n1201), .ZN(n1139) );
NOR2_X1 U908 ( .A1(n1199), .A2(n1204), .ZN(n1009) );
XNOR2_X1 U909 ( .A(G113), .B(n1136), .ZN(G15) );
NAND3_X1 U910 ( .A1(n1145), .A2(n1181), .A3(n1201), .ZN(n1136) );
AND3_X1 U911 ( .A1(n1193), .A2(n1144), .A3(n1189), .ZN(n1201) );
INV_X1 U912 ( .A(n1156), .ZN(n1189) );
NAND3_X1 U913 ( .A1(n1034), .A2(n1010), .A3(n1197), .ZN(n1156) );
INV_X1 U914 ( .A(n1019), .ZN(n1193) );
INV_X1 U915 ( .A(n1036), .ZN(n1145) );
NAND2_X1 U916 ( .A1(n1204), .A2(n1199), .ZN(n1036) );
INV_X1 U917 ( .A(n1198), .ZN(n1204) );
XNOR2_X1 U918 ( .A(G110), .B(n1135), .ZN(G12) );
NAND4_X1 U919 ( .A1(n1014), .A2(n1141), .A3(n1019), .A4(n1020), .ZN(n1135) );
INV_X1 U920 ( .A(n1181), .ZN(n1020) );
NOR2_X1 U921 ( .A1(n1205), .A2(n1041), .ZN(n1181) );
NOR2_X1 U922 ( .A1(n1047), .A2(n1046), .ZN(n1041) );
AND2_X1 U923 ( .A1(n1046), .A2(n1047), .ZN(n1205) );
NAND2_X1 U924 ( .A1(n1089), .A2(n1206), .ZN(n1047) );
XOR2_X1 U925 ( .A(n1207), .B(n1208), .Z(n1089) );
XNOR2_X1 U926 ( .A(n1209), .B(n1210), .ZN(n1208) );
XOR2_X1 U927 ( .A(n1211), .B(n1212), .Z(n1210) );
NAND2_X1 U928 ( .A1(G221), .A2(n1213), .ZN(n1211) );
XOR2_X1 U929 ( .A(n1214), .B(n1215), .Z(n1207) );
NOR2_X1 U930 ( .A1(KEYINPUT13), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U931 ( .A(n1217), .B(n1218), .ZN(n1216) );
INV_X1 U932 ( .A(n1219), .ZN(n1218) );
NAND2_X1 U933 ( .A1(n1220), .A2(KEYINPUT52), .ZN(n1217) );
XNOR2_X1 U934 ( .A(G125), .B(KEYINPUT44), .ZN(n1220) );
XNOR2_X1 U935 ( .A(G128), .B(G137), .ZN(n1214) );
AND2_X1 U936 ( .A1(G217), .A2(n1221), .ZN(n1046) );
XOR2_X1 U937 ( .A(n1043), .B(KEYINPUT33), .Z(n1019) );
XNOR2_X1 U938 ( .A(n1222), .B(G472), .ZN(n1043) );
NAND2_X1 U939 ( .A1(n1223), .A2(n1206), .ZN(n1222) );
XNOR2_X1 U940 ( .A(n1106), .B(n1224), .ZN(n1223) );
XOR2_X1 U941 ( .A(n1225), .B(n1226), .Z(n1224) );
NAND2_X1 U942 ( .A1(KEYINPUT57), .A2(n1112), .ZN(n1226) );
INV_X1 U943 ( .A(G101), .ZN(n1112) );
NAND2_X1 U944 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
NAND2_X1 U945 ( .A1(n1109), .A2(n1108), .ZN(n1228) );
XOR2_X1 U946 ( .A(n1229), .B(KEYINPUT39), .Z(n1227) );
OR2_X1 U947 ( .A1(n1108), .A2(n1109), .ZN(n1229) );
XNOR2_X1 U948 ( .A(n1230), .B(n1231), .ZN(n1106) );
XOR2_X1 U949 ( .A(G113), .B(n1232), .Z(n1231) );
NOR2_X1 U950 ( .A1(KEYINPUT30), .A2(n1233), .ZN(n1232) );
XNOR2_X1 U951 ( .A(G116), .B(G119), .ZN(n1233) );
NAND2_X1 U952 ( .A1(G210), .A2(n1234), .ZN(n1230) );
AND3_X1 U953 ( .A1(n1034), .A2(n1144), .A3(n1158), .ZN(n1141) );
NOR2_X1 U954 ( .A1(n1197), .A2(n1015), .ZN(n1158) );
INV_X1 U955 ( .A(n1010), .ZN(n1015) );
NAND2_X1 U956 ( .A1(G221), .A2(n1221), .ZN(n1010) );
NAND2_X1 U957 ( .A1(G234), .A2(n1206), .ZN(n1221) );
XOR2_X1 U958 ( .A(n1235), .B(n1119), .Z(n1197) );
INV_X1 U959 ( .A(G469), .ZN(n1119) );
NAND2_X1 U960 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U961 ( .A1(KEYINPUT23), .A2(n1048), .ZN(n1237) );
OR2_X1 U962 ( .A1(KEYINPUT41), .A2(n1048), .ZN(n1236) );
AND2_X1 U963 ( .A1(n1238), .A2(n1206), .ZN(n1048) );
XOR2_X1 U964 ( .A(n1239), .B(n1240), .Z(n1238) );
XNOR2_X1 U965 ( .A(n1241), .B(n1065), .ZN(n1240) );
INV_X1 U966 ( .A(n1127), .ZN(n1065) );
XOR2_X1 U967 ( .A(n1242), .B(n1243), .Z(n1127) );
NOR2_X1 U968 ( .A1(G128), .A2(KEYINPUT19), .ZN(n1243) );
XNOR2_X1 U969 ( .A(n1115), .B(n1124), .ZN(n1241) );
XNOR2_X1 U970 ( .A(n1244), .B(n1245), .ZN(n1124) );
XOR2_X1 U971 ( .A(n1219), .B(n1246), .Z(n1115) );
XOR2_X1 U972 ( .A(G110), .B(n1247), .Z(n1246) );
NOR2_X1 U973 ( .A1(G953), .A2(n1056), .ZN(n1247) );
INV_X1 U974 ( .A(G227), .ZN(n1056) );
XOR2_X1 U975 ( .A(n1248), .B(n1109), .Z(n1239) );
XOR2_X1 U976 ( .A(n1249), .B(n1176), .Z(n1109) );
INV_X1 U977 ( .A(G131), .ZN(n1176) );
NAND3_X1 U978 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1249) );
NAND2_X1 U979 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
OR3_X1 U980 ( .A1(n1254), .A2(n1253), .A3(KEYINPUT2), .ZN(n1251) );
XOR2_X1 U981 ( .A(G134), .B(KEYINPUT58), .Z(n1253) );
OR2_X1 U982 ( .A1(G137), .A2(KEYINPUT47), .ZN(n1254) );
NAND2_X1 U983 ( .A1(KEYINPUT2), .A2(G137), .ZN(n1250) );
XNOR2_X1 U984 ( .A(KEYINPUT49), .B(KEYINPUT38), .ZN(n1248) );
NAND2_X1 U985 ( .A1(n998), .A2(n1255), .ZN(n1144) );
NAND3_X1 U986 ( .A1(G902), .A2(n1195), .A3(n1081), .ZN(n1255) );
NOR2_X1 U987 ( .A1(n1256), .A2(G898), .ZN(n1081) );
INV_X1 U988 ( .A(n1060), .ZN(n1256) );
XNOR2_X1 U989 ( .A(G953), .B(KEYINPUT10), .ZN(n1060) );
NAND3_X1 U990 ( .A1(n1195), .A2(n1053), .A3(G952), .ZN(n998) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1195) );
NOR2_X1 U992 ( .A1(n1022), .A2(n1024), .ZN(n1034) );
INV_X1 U993 ( .A(n1177), .ZN(n1024) );
NAND2_X1 U994 ( .A1(n1257), .A2(n1258), .ZN(n1177) );
XOR2_X1 U995 ( .A(KEYINPUT21), .B(G214), .Z(n1257) );
XNOR2_X1 U996 ( .A(n1259), .B(n1132), .ZN(n1022) );
NAND2_X1 U997 ( .A1(G210), .A2(n1258), .ZN(n1132) );
NAND2_X1 U998 ( .A1(n1260), .A2(n1206), .ZN(n1258) );
INV_X1 U999 ( .A(G237), .ZN(n1260) );
NAND2_X1 U1000 ( .A1(n1261), .A2(n1206), .ZN(n1259) );
XNOR2_X1 U1001 ( .A(n1078), .B(n1262), .ZN(n1261) );
XOR2_X1 U1002 ( .A(n1263), .B(n1164), .Z(n1262) );
XNOR2_X1 U1003 ( .A(G125), .B(n1108), .ZN(n1164) );
XOR2_X1 U1004 ( .A(G128), .B(n1242), .Z(n1108) );
XOR2_X1 U1005 ( .A(G146), .B(G143), .Z(n1242) );
NAND2_X1 U1006 ( .A1(KEYINPUT54), .A2(n1264), .ZN(n1263) );
XNOR2_X1 U1007 ( .A(KEYINPUT26), .B(n1166), .ZN(n1264) );
NAND2_X1 U1008 ( .A1(G224), .A2(n1053), .ZN(n1166) );
XNOR2_X1 U1009 ( .A(n1265), .B(n1266), .ZN(n1078) );
XOR2_X1 U1010 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U1011 ( .A(KEYINPUT24), .B(G113), .Z(n1268) );
XOR2_X1 U1012 ( .A(n1269), .B(n1212), .Z(n1265) );
XOR2_X1 U1013 ( .A(G110), .B(G119), .Z(n1212) );
NAND2_X1 U1014 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U1015 ( .A1(n1272), .A2(n1245), .ZN(n1271) );
INV_X1 U1016 ( .A(n1273), .ZN(n1245) );
XOR2_X1 U1017 ( .A(KEYINPUT0), .B(n1244), .Z(n1272) );
NAND2_X1 U1018 ( .A1(n1244), .A2(n1273), .ZN(n1270) );
XOR2_X1 U1019 ( .A(G104), .B(G101), .Z(n1244) );
NOR2_X1 U1020 ( .A1(n1198), .A2(n1199), .ZN(n1014) );
XNOR2_X1 U1021 ( .A(n1274), .B(G475), .ZN(n1199) );
NAND2_X1 U1022 ( .A1(n1100), .A2(n1206), .ZN(n1274) );
XOR2_X1 U1023 ( .A(n1275), .B(n1276), .Z(n1100) );
XNOR2_X1 U1024 ( .A(n1277), .B(n1278), .ZN(n1276) );
NOR2_X1 U1025 ( .A1(KEYINPUT7), .A2(n1279), .ZN(n1278) );
XOR2_X1 U1026 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U1027 ( .A(n1282), .B(n1283), .ZN(n1281) );
NOR2_X1 U1028 ( .A1(KEYINPUT20), .A2(n1284), .ZN(n1283) );
XOR2_X1 U1029 ( .A(n1064), .B(n1285), .Z(n1284) );
XNOR2_X1 U1030 ( .A(n1286), .B(KEYINPUT37), .ZN(n1285) );
NAND2_X1 U1031 ( .A1(KEYINPUT8), .A2(n1287), .ZN(n1286) );
XOR2_X1 U1032 ( .A(KEYINPUT59), .B(n1209), .Z(n1287) );
XOR2_X1 U1033 ( .A(G146), .B(KEYINPUT5), .Z(n1209) );
XNOR2_X1 U1034 ( .A(G125), .B(n1219), .ZN(n1064) );
XOR2_X1 U1035 ( .A(G140), .B(KEYINPUT17), .Z(n1219) );
NAND3_X1 U1036 ( .A1(G214), .A2(n1234), .A3(KEYINPUT61), .ZN(n1282) );
NOR2_X1 U1037 ( .A1(G953), .A2(G237), .ZN(n1234) );
XNOR2_X1 U1038 ( .A(G131), .B(G143), .ZN(n1280) );
INV_X1 U1039 ( .A(G104), .ZN(n1277) );
XNOR2_X1 U1040 ( .A(G122), .B(G113), .ZN(n1275) );
XNOR2_X1 U1041 ( .A(n1288), .B(G478), .ZN(n1198) );
NAND2_X1 U1042 ( .A1(n1094), .A2(n1289), .ZN(n1288) );
XNOR2_X1 U1043 ( .A(KEYINPUT35), .B(n1206), .ZN(n1289) );
INV_X1 U1044 ( .A(G902), .ZN(n1206) );
XOR2_X1 U1045 ( .A(n1290), .B(n1291), .Z(n1094) );
XOR2_X1 U1046 ( .A(n1292), .B(n1293), .Z(n1291) );
NOR2_X1 U1047 ( .A1(G134), .A2(KEYINPUT48), .ZN(n1293) );
AND2_X1 U1048 ( .A1(n1213), .A2(G217), .ZN(n1292) );
AND2_X1 U1049 ( .A1(G234), .A2(n1053), .ZN(n1213) );
INV_X1 U1050 ( .A(G953), .ZN(n1053) );
XOR2_X1 U1051 ( .A(n1294), .B(n1295), .Z(n1290) );
NOR2_X1 U1052 ( .A1(KEYINPUT51), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U1053 ( .A(n1267), .B(n1273), .ZN(n1296) );
XOR2_X1 U1054 ( .A(G107), .B(KEYINPUT18), .Z(n1273) );
XOR2_X1 U1055 ( .A(G116), .B(G122), .Z(n1267) );
XNOR2_X1 U1056 ( .A(G128), .B(G143), .ZN(n1294) );
endmodule


