//Key = 0101000110110110101100000100010000101100101101001001010010111011


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
n2292, n2293, n2294, n2295, n2296, n2297, n2298;

OR2_X1 U1281 ( .A1(n2298), .A2(n1723), .ZN(U280) );
OR2_X1 U1282 ( .A1(n1873), .A2(STATO_REG_0__SCAN_IN), .ZN(n1722) );
INV_X2 U1283 ( .A(n1722), .ZN(n1723) );
INV_X2 U1284 ( .A(U280), .ZN(n1724) );
NOR3_X2 U1285 ( .A1(n1872), .A2(n2205), .A3(n2297), .ZN(n1953) );
XOR2_X1 U1286 ( .A(n1725), .B(KEYINPUT43), .Z(U375) );
NAND2_X1 U1287 ( .A1(n1726), .A2(n1727), .ZN(U344) );
NAND2_X1 U1288 ( .A1(DATA_IN_7_), .A2(n1728), .ZN(n1727) );
NAND2_X1 U1289 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1729), .ZN(n1726) );
NAND2_X1 U1290 ( .A1(n1730), .A2(n1731), .ZN(U343) );
NAND2_X1 U1291 ( .A1(n1732), .A2(DATA_IN_6_), .ZN(n1731) );
XOR2_X1 U1292 ( .A(n1728), .B(KEYINPUT35), .Z(n1732) );
NAND2_X1 U1293 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1729), .ZN(n1730) );
NAND2_X1 U1294 ( .A1(n1733), .A2(n1734), .ZN(U342) );
NAND2_X1 U1295 ( .A1(DATA_IN_5_), .A2(n1728), .ZN(n1734) );
NAND2_X1 U1296 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1729), .ZN(n1733) );
NAND2_X1 U1297 ( .A1(n1735), .A2(n1736), .ZN(U341) );
NAND2_X1 U1298 ( .A1(DATA_IN_4_), .A2(n1728), .ZN(n1736) );
NAND2_X1 U1299 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1729), .ZN(n1735) );
NAND2_X1 U1300 ( .A1(n1737), .A2(n1738), .ZN(U340) );
NAND2_X1 U1301 ( .A1(DATA_IN_3_), .A2(n1728), .ZN(n1738) );
NAND2_X1 U1302 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1729), .ZN(n1737) );
NAND2_X1 U1303 ( .A1(n1739), .A2(n1740), .ZN(U339) );
NAND2_X1 U1304 ( .A1(n1741), .A2(DATA_IN_2_), .ZN(n1740) );
XOR2_X1 U1305 ( .A(n1728), .B(KEYINPUT2), .Z(n1741) );
NAND2_X1 U1306 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1729), .ZN(n1739) );
NAND2_X1 U1307 ( .A1(n1742), .A2(n1743), .ZN(U338) );
NAND2_X1 U1308 ( .A1(DATA_IN_1_), .A2(n1728), .ZN(n1743) );
NAND2_X1 U1309 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1729), .ZN(n1742) );
NAND2_X1 U1310 ( .A1(n1744), .A2(n1745), .ZN(U337) );
NAND2_X1 U1311 ( .A1(n1746), .A2(n1728), .ZN(n1745) );
NAND2_X1 U1312 ( .A1(n1747), .A2(n1748), .ZN(n1728) );
NAND2_X1 U1313 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1749), .ZN(n1748) );
XOR2_X1 U1314 ( .A(STATO_REG_0__SCAN_IN), .B(KEYINPUT45), .Z(n1747) );
XOR2_X1 U1315 ( .A(KEYINPUT24), .B(DATA_IN_0_), .Z(n1746) );
NAND2_X1 U1316 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1729), .ZN(n1744) );
NAND2_X1 U1317 ( .A1(n1725), .A2(n1750), .ZN(n1729) );
NAND2_X1 U1318 ( .A1(n1751), .A2(n1752), .ZN(n1750) );
NAND2_X1 U1319 ( .A1(n1753), .A2(n1754), .ZN(U336) );
NAND2_X1 U1320 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1755), .ZN(n1754) );
NAND2_X1 U1321 ( .A1(n1756), .A2(DATA_IN_7_), .ZN(n1753) );
NAND2_X1 U1322 ( .A1(n1757), .A2(n1758), .ZN(U335) );
NAND2_X1 U1323 ( .A1(n1756), .A2(DATA_IN_6_), .ZN(n1758) );
XOR2_X1 U1324 ( .A(n1759), .B(KEYINPUT15), .Z(n1757) );
NAND2_X1 U1325 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1755), .ZN(n1759) );
NAND2_X1 U1326 ( .A1(n1760), .A2(n1761), .ZN(U334) );
NAND2_X1 U1327 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1755), .ZN(n1761) );
NAND2_X1 U1328 ( .A1(n1756), .A2(DATA_IN_5_), .ZN(n1760) );
NAND2_X1 U1329 ( .A1(n1762), .A2(n1763), .ZN(U333) );
NAND2_X1 U1330 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1755), .ZN(n1763) );
NAND2_X1 U1331 ( .A1(n1756), .A2(DATA_IN_4_), .ZN(n1762) );
NAND2_X1 U1332 ( .A1(n1764), .A2(n1765), .ZN(U332) );
NAND2_X1 U1333 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1755), .ZN(n1765) );
NAND2_X1 U1334 ( .A1(n1756), .A2(DATA_IN_3_), .ZN(n1764) );
NAND2_X1 U1335 ( .A1(n1766), .A2(n1767), .ZN(U331) );
NAND2_X1 U1336 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1755), .ZN(n1767) );
NAND2_X1 U1337 ( .A1(n1756), .A2(DATA_IN_2_), .ZN(n1766) );
NAND2_X1 U1338 ( .A1(n1768), .A2(n1769), .ZN(U330) );
NAND2_X1 U1339 ( .A1(n1756), .A2(DATA_IN_1_), .ZN(n1769) );
XOR2_X1 U1340 ( .A(KEYINPUT56), .B(n1770), .Z(n1768) );
AND2_X1 U1341 ( .A1(n1755), .A2(RMIN_REG_1__SCAN_IN), .ZN(n1770) );
NAND2_X1 U1342 ( .A1(n1771), .A2(n1772), .ZN(U329) );
NAND2_X1 U1343 ( .A1(n1773), .A2(n1755), .ZN(n1772) );
NAND2_X1 U1344 ( .A1(n1725), .A2(n1774), .ZN(n1755) );
NAND2_X1 U1345 ( .A1(n1775), .A2(n1752), .ZN(n1774) );
XNOR2_X1 U1346 ( .A(KEYINPUT7), .B(n1776), .ZN(n1775) );
XOR2_X1 U1347 ( .A(RMIN_REG_0__SCAN_IN), .B(KEYINPUT4), .Z(n1773) );
NAND2_X1 U1348 ( .A1(n1756), .A2(DATA_IN_0_), .ZN(n1771) );
AND2_X1 U1349 ( .A1(n1777), .A2(n1725), .ZN(n1756) );
NAND2_X1 U1350 ( .A1(n1752), .A2(n1776), .ZN(n1777) );
NAND2_X1 U1351 ( .A1(n1751), .A2(n1778), .ZN(n1776) );
NAND2_X1 U1352 ( .A1(n1779), .A2(n1780), .ZN(n1778) );
NAND3_X1 U1353 ( .A1(n1781), .A2(n1782), .A3(n1783), .ZN(n1780) );
NAND2_X1 U1354 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1784), .ZN(n1783) );
NAND3_X1 U1355 ( .A1(n1785), .A2(n1786), .A3(n1787), .ZN(n1782) );
NAND2_X1 U1356 ( .A1(n1788), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1787) );
XOR2_X1 U1357 ( .A(n1789), .B(KEYINPUT50), .Z(n1788) );
NAND3_X1 U1358 ( .A1(n1790), .A2(n1791), .A3(n1792), .ZN(n1786) );
NAND2_X1 U1359 ( .A1(DATA_IN_5_), .A2(n1793), .ZN(n1792) );
NAND3_X1 U1360 ( .A1(n1794), .A2(n1795), .A3(n1796), .ZN(n1791) );
NAND2_X1 U1361 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1797), .ZN(n1796) );
NAND3_X1 U1362 ( .A1(n1798), .A2(n1799), .A3(n1800), .ZN(n1795) );
NAND2_X1 U1363 ( .A1(DATA_IN_3_), .A2(n1801), .ZN(n1800) );
NAND3_X1 U1364 ( .A1(n1802), .A2(n1803), .A3(n1804), .ZN(n1799) );
NAND2_X1 U1365 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1805), .ZN(n1804) );
NAND2_X1 U1366 ( .A1(n1806), .A2(n1807), .ZN(n1805) );
NAND2_X1 U1367 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1808), .ZN(n1807) );
XOR2_X1 U1368 ( .A(n1809), .B(KEYINPUT3), .Z(n1806) );
NAND3_X1 U1369 ( .A1(n1808), .A2(n1809), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1803) );
NAND2_X1 U1370 ( .A1(n1810), .A2(n1811), .ZN(n1802) );
XOR2_X1 U1371 ( .A(n1812), .B(KEYINPUT34), .Z(n1810) );
NAND2_X1 U1372 ( .A1(DATA_IN_2_), .A2(n1812), .ZN(n1798) );
NAND2_X1 U1373 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1813), .ZN(n1794) );
NAND2_X1 U1374 ( .A1(DATA_IN_4_), .A2(n1814), .ZN(n1790) );
NAND2_X1 U1375 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1815), .ZN(n1785) );
XOR2_X1 U1376 ( .A(KEYINPUT58), .B(DATA_IN_5_), .Z(n1815) );
NAND2_X1 U1377 ( .A1(n1816), .A2(DATA_IN_6_), .ZN(n1781) );
XOR2_X1 U1378 ( .A(n1817), .B(KEYINPUT17), .Z(n1816) );
NAND2_X1 U1379 ( .A1(DATA_IN_7_), .A2(n1818), .ZN(n1779) );
INV_X1 U1380 ( .A(n1749), .ZN(n1751) );
NAND2_X1 U1381 ( .A1(n1819), .A2(n1820), .ZN(n1749) );
NAND2_X1 U1382 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1784), .ZN(n1820) );
NAND3_X1 U1383 ( .A1(n1821), .A2(n1822), .A3(n1823), .ZN(n1819) );
NAND2_X1 U1384 ( .A1(DATA_IN_7_), .A2(n1824), .ZN(n1823) );
NAND3_X1 U1385 ( .A1(n1825), .A2(n1826), .A3(n1827), .ZN(n1822) );
NAND2_X1 U1386 ( .A1(DATA_IN_6_), .A2(n1828), .ZN(n1827) );
NAND3_X1 U1387 ( .A1(n1829), .A2(n1830), .A3(n1831), .ZN(n1826) );
NAND2_X1 U1388 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1797), .ZN(n1831) );
NAND3_X1 U1389 ( .A1(n1832), .A2(n1833), .A3(n1834), .ZN(n1830) );
NAND2_X1 U1390 ( .A1(DATA_IN_4_), .A2(n1835), .ZN(n1834) );
NAND3_X1 U1391 ( .A1(n1836), .A2(n1837), .A3(n1838), .ZN(n1833) );
XOR2_X1 U1392 ( .A(n1839), .B(KEYINPUT32), .Z(n1838) );
NAND2_X1 U1393 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1813), .ZN(n1839) );
NAND3_X1 U1394 ( .A1(n1840), .A2(n1841), .A3(n1842), .ZN(n1837) );
NAND2_X1 U1395 ( .A1(DATA_IN_2_), .A2(n1843), .ZN(n1842) );
NAND3_X1 U1396 ( .A1(n1844), .A2(n1845), .A3(n1846), .ZN(n1841) );
XOR2_X1 U1397 ( .A(n1808), .B(KEYINPUT11), .Z(n1846) );
NAND2_X1 U1398 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1809), .ZN(n1845) );
XOR2_X1 U1399 ( .A(RMAX_REG_0__SCAN_IN), .B(KEYINPUT19), .Z(n1844) );
NAND2_X1 U1400 ( .A1(DATA_IN_1_), .A2(n1847), .ZN(n1840) );
NAND2_X1 U1401 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1811), .ZN(n1836) );
NAND2_X1 U1402 ( .A1(DATA_IN_3_), .A2(n1848), .ZN(n1832) );
NAND2_X1 U1403 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1849), .ZN(n1829) );
XOR2_X1 U1404 ( .A(KEYINPUT14), .B(DATA_IN_5_), .Z(n1849) );
NAND2_X1 U1405 ( .A1(DATA_IN_5_), .A2(n1850), .ZN(n1825) );
NAND2_X1 U1406 ( .A1(n1851), .A2(n1789), .ZN(n1821) );
INV_X1 U1407 ( .A(DATA_IN_6_), .ZN(n1789) );
XOR2_X1 U1408 ( .A(RMAX_REG_6__SCAN_IN), .B(KEYINPUT54), .Z(n1851) );
NAND2_X1 U1409 ( .A1(n1852), .A2(n1853), .ZN(U328) );
NAND2_X1 U1410 ( .A1(n1854), .A2(DATA_IN_7_), .ZN(n1853) );
NAND2_X1 U1411 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1855), .ZN(n1852) );
NAND2_X1 U1412 ( .A1(n1856), .A2(n1857), .ZN(U327) );
NAND2_X1 U1413 ( .A1(n1854), .A2(DATA_IN_6_), .ZN(n1857) );
NAND2_X1 U1414 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1855), .ZN(n1856) );
NAND2_X1 U1415 ( .A1(n1858), .A2(n1859), .ZN(U326) );
NAND2_X1 U1416 ( .A1(n1854), .A2(DATA_IN_5_), .ZN(n1859) );
NAND2_X1 U1417 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1855), .ZN(n1858) );
NAND2_X1 U1418 ( .A1(n1860), .A2(n1861), .ZN(U325) );
NAND2_X1 U1419 ( .A1(n1854), .A2(DATA_IN_4_), .ZN(n1861) );
NAND2_X1 U1420 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1855), .ZN(n1860) );
NAND2_X1 U1421 ( .A1(n1862), .A2(n1863), .ZN(U324) );
NAND2_X1 U1422 ( .A1(n1854), .A2(DATA_IN_3_), .ZN(n1863) );
NAND2_X1 U1423 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1855), .ZN(n1862) );
NAND2_X1 U1424 ( .A1(n1864), .A2(n1865), .ZN(U323) );
NAND2_X1 U1425 ( .A1(n1854), .A2(DATA_IN_2_), .ZN(n1865) );
NAND2_X1 U1426 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1855), .ZN(n1864) );
NAND2_X1 U1427 ( .A1(n1866), .A2(n1867), .ZN(U322) );
NAND2_X1 U1428 ( .A1(n1854), .A2(DATA_IN_1_), .ZN(n1867) );
NAND2_X1 U1429 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1855), .ZN(n1866) );
NAND2_X1 U1430 ( .A1(n1868), .A2(n1869), .ZN(U321) );
NAND2_X1 U1431 ( .A1(n1854), .A2(DATA_IN_0_), .ZN(n1869) );
AND2_X1 U1432 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1870), .ZN(n1854) );
NAND2_X1 U1433 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1855), .ZN(n1868) );
NAND2_X1 U1434 ( .A1(n1871), .A2(n1870), .ZN(n1855) );
NAND2_X1 U1435 ( .A1(n1752), .A2(n1872), .ZN(n1870) );
XNOR2_X1 U1436 ( .A(KEYINPUT8), .B(n1725), .ZN(n1871) );
NAND2_X1 U1437 ( .A1(n1873), .A2(n1752), .ZN(n1725) );
NAND2_X1 U1438 ( .A1(n1874), .A2(n1875), .ZN(U320) );
NAND2_X1 U1439 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1724), .ZN(n1875) );
NAND2_X1 U1440 ( .A1(n1723), .A2(DATA_IN_7_), .ZN(n1874) );
NAND2_X1 U1441 ( .A1(n1876), .A2(n1877), .ZN(U319) );
NAND2_X1 U1442 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1724), .ZN(n1877) );
NAND2_X1 U1443 ( .A1(n1723), .A2(DATA_IN_6_), .ZN(n1876) );
NAND2_X1 U1444 ( .A1(n1878), .A2(n1879), .ZN(U318) );
NAND2_X1 U1445 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1724), .ZN(n1879) );
NAND2_X1 U1446 ( .A1(n1723), .A2(DATA_IN_5_), .ZN(n1878) );
NAND2_X1 U1447 ( .A1(n1880), .A2(n1881), .ZN(U317) );
NAND2_X1 U1448 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1724), .ZN(n1881) );
NAND2_X1 U1449 ( .A1(n1723), .A2(DATA_IN_4_), .ZN(n1880) );
NAND2_X1 U1450 ( .A1(n1882), .A2(n1883), .ZN(U316) );
NAND2_X1 U1451 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1724), .ZN(n1883) );
NAND2_X1 U1452 ( .A1(n1723), .A2(DATA_IN_3_), .ZN(n1882) );
NAND2_X1 U1453 ( .A1(n1884), .A2(n1885), .ZN(U315) );
NAND2_X1 U1454 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1724), .ZN(n1885) );
NAND2_X1 U1455 ( .A1(n1723), .A2(DATA_IN_2_), .ZN(n1884) );
NAND2_X1 U1456 ( .A1(n1886), .A2(n1887), .ZN(U314) );
NAND2_X1 U1457 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1724), .ZN(n1887) );
NAND2_X1 U1458 ( .A1(n1723), .A2(DATA_IN_1_), .ZN(n1886) );
NAND2_X1 U1459 ( .A1(n1888), .A2(n1889), .ZN(U313) );
NAND2_X1 U1460 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1724), .ZN(n1889) );
NAND2_X1 U1461 ( .A1(n1723), .A2(DATA_IN_0_), .ZN(n1888) );
NAND2_X1 U1462 ( .A1(n1890), .A2(n1891), .ZN(U312) );
NAND2_X1 U1463 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1724), .ZN(n1891) );
NAND2_X1 U1464 ( .A1(n1723), .A2(REG1_REG_7__SCAN_IN), .ZN(n1890) );
NAND2_X1 U1465 ( .A1(n1892), .A2(n1893), .ZN(U311) );
NAND2_X1 U1466 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1724), .ZN(n1893) );
NAND2_X1 U1467 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1723), .ZN(n1892) );
NAND2_X1 U1468 ( .A1(n1894), .A2(n1895), .ZN(U310) );
NAND2_X1 U1469 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1724), .ZN(n1895) );
NAND2_X1 U1470 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1723), .ZN(n1894) );
NAND2_X1 U1471 ( .A1(n1896), .A2(n1897), .ZN(U309) );
NAND2_X1 U1472 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1724), .ZN(n1897) );
NAND2_X1 U1473 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1723), .ZN(n1896) );
NAND2_X1 U1474 ( .A1(n1898), .A2(n1899), .ZN(U308) );
NAND2_X1 U1475 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1724), .ZN(n1899) );
XOR2_X1 U1476 ( .A(KEYINPUT63), .B(n1900), .Z(n1898) );
AND2_X1 U1477 ( .A1(n1723), .A2(REG1_REG_3__SCAN_IN), .ZN(n1900) );
NAND2_X1 U1478 ( .A1(n1901), .A2(n1902), .ZN(U307) );
NAND2_X1 U1479 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1724), .ZN(n1902) );
NAND2_X1 U1480 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1723), .ZN(n1901) );
NAND2_X1 U1481 ( .A1(n1903), .A2(n1904), .ZN(U306) );
NAND2_X1 U1482 ( .A1(n1905), .A2(n1724), .ZN(n1904) );
XOR2_X1 U1483 ( .A(REG2_REG_1__SCAN_IN), .B(KEYINPUT44), .Z(n1905) );
NAND2_X1 U1484 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1723), .ZN(n1903) );
NAND2_X1 U1485 ( .A1(n1906), .A2(n1907), .ZN(U305) );
NAND2_X1 U1486 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1724), .ZN(n1907) );
NAND2_X1 U1487 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1723), .ZN(n1906) );
NAND2_X1 U1488 ( .A1(n1908), .A2(n1909), .ZN(U304) );
NAND2_X1 U1489 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1724), .ZN(n1909) );
NAND2_X1 U1490 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1723), .ZN(n1908) );
NAND2_X1 U1491 ( .A1(n1910), .A2(n1911), .ZN(U303) );
NAND2_X1 U1492 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1724), .ZN(n1911) );
NAND2_X1 U1493 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1723), .ZN(n1910) );
NAND2_X1 U1494 ( .A1(n1912), .A2(n1913), .ZN(U302) );
NAND2_X1 U1495 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1724), .ZN(n1913) );
NAND2_X1 U1496 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1723), .ZN(n1912) );
NAND2_X1 U1497 ( .A1(n1914), .A2(n1915), .ZN(U301) );
NAND2_X1 U1498 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1724), .ZN(n1915) );
NAND2_X1 U1499 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1723), .ZN(n1914) );
NAND2_X1 U1500 ( .A1(n1916), .A2(n1917), .ZN(U300) );
NAND2_X1 U1501 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1724), .ZN(n1917) );
NAND2_X1 U1502 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1723), .ZN(n1916) );
NAND2_X1 U1503 ( .A1(n1918), .A2(n1919), .ZN(U299) );
NAND2_X1 U1504 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1724), .ZN(n1919) );
NAND2_X1 U1505 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1723), .ZN(n1918) );
NAND2_X1 U1506 ( .A1(n1920), .A2(n1921), .ZN(U298) );
NAND2_X1 U1507 ( .A1(n1922), .A2(n1723), .ZN(n1921) );
XNOR2_X1 U1508 ( .A(REG2_REG_1__SCAN_IN), .B(KEYINPUT36), .ZN(n1922) );
NAND2_X1 U1509 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1724), .ZN(n1920) );
NAND2_X1 U1510 ( .A1(n1923), .A2(n1924), .ZN(U297) );
NAND2_X1 U1511 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1724), .ZN(n1924) );
NAND2_X1 U1512 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1723), .ZN(n1923) );
NAND2_X1 U1513 ( .A1(n1925), .A2(n1926), .ZN(U296) );
NAND2_X1 U1514 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1724), .ZN(n1926) );
NAND2_X1 U1515 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1723), .ZN(n1925) );
NAND2_X1 U1516 ( .A1(n1927), .A2(n1928), .ZN(U295) );
NAND2_X1 U1517 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1724), .ZN(n1928) );
NAND2_X1 U1518 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1723), .ZN(n1927) );
NAND2_X1 U1519 ( .A1(n1929), .A2(n1930), .ZN(U294) );
NAND2_X1 U1520 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1724), .ZN(n1930) );
XOR2_X1 U1521 ( .A(KEYINPUT13), .B(n1931), .Z(n1929) );
AND2_X1 U1522 ( .A1(n1723), .A2(REG3_REG_5__SCAN_IN), .ZN(n1931) );
NAND2_X1 U1523 ( .A1(n1932), .A2(n1933), .ZN(U293) );
NAND2_X1 U1524 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1724), .ZN(n1933) );
NAND2_X1 U1525 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1723), .ZN(n1932) );
NAND2_X1 U1526 ( .A1(n1934), .A2(n1935), .ZN(U292) );
NAND2_X1 U1527 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1724), .ZN(n1935) );
XOR2_X1 U1528 ( .A(KEYINPUT10), .B(n1936), .Z(n1934) );
AND2_X1 U1529 ( .A1(n1723), .A2(REG3_REG_3__SCAN_IN), .ZN(n1936) );
NAND2_X1 U1530 ( .A1(n1937), .A2(n1938), .ZN(U291) );
NAND2_X1 U1531 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1724), .ZN(n1938) );
NAND2_X1 U1532 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1723), .ZN(n1937) );
NAND2_X1 U1533 ( .A1(n1939), .A2(n1940), .ZN(U290) );
NAND2_X1 U1534 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1724), .ZN(n1940) );
NAND2_X1 U1535 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1723), .ZN(n1939) );
NAND2_X1 U1536 ( .A1(n1941), .A2(n1942), .ZN(U289) );
NAND2_X1 U1537 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1724), .ZN(n1942) );
NAND2_X1 U1538 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1723), .ZN(n1941) );
NAND4_X1 U1539 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .ZN(U288));
NAND2_X1 U1540 ( .A1(n1947), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1946) );
NOR2_X1 U1541 ( .A1(n1948), .A2(n1949), .ZN(n1945) );
AND3_X1 U1542 ( .A1(n1950), .A2(n1951), .A3(n1952), .ZN(n1949) );
NAND2_X1 U1543 ( .A1(n1953), .A2(REG4_REG_7__SCAN_IN), .ZN(n1944) );
NAND2_X1 U1544 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1724), .ZN(n1943) );
NAND4_X1 U1545 ( .A1(n1954), .A2(n1955), .A3(n1956), .A4(n1957), .ZN(U287));
NOR3_X1 U1546 ( .A1(n1958), .A2(n1948), .A3(n1959), .ZN(n1957) );
NOR3_X1 U1547 ( .A1(n1960), .A2(n1961), .A3(n1962), .ZN(n1959) );
AND3_X1 U1548 ( .A1(n1961), .A2(n1960), .A3(n1963), .ZN(n1948) );
NAND2_X1 U1549 ( .A1(n1964), .A2(n1965), .ZN(n1960) );
OR2_X1 U1550 ( .A1(n1966), .A2(n1967), .ZN(n1965) );
NOR2_X1 U1551 ( .A1(n1968), .A2(n1969), .ZN(n1958) );
XOR2_X1 U1552 ( .A(KEYINPUT51), .B(n1947), .Z(n1969) );
INV_X1 U1553 ( .A(RLAST_REG_6__SCAN_IN), .ZN(n1968) );
XOR2_X1 U1554 ( .A(n1970), .B(KEYINPUT5), .Z(n1956) );
NAND2_X1 U1555 ( .A1(n1971), .A2(n1952), .ZN(n1970) );
XOR2_X1 U1556 ( .A(n1951), .B(n1972), .Z(n1971) );
NOR2_X1 U1557 ( .A1(n1950), .A2(KEYINPUT28), .ZN(n1972) );
NAND2_X1 U1558 ( .A1(n1953), .A2(REG4_REG_6__SCAN_IN), .ZN(n1955) );
NAND2_X1 U1559 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1724), .ZN(n1954) );
NAND4_X1 U1560 ( .A1(n1973), .A2(n1974), .A3(n1975), .A4(n1976), .ZN(U286));
NOR3_X1 U1561 ( .A1(n1977), .A2(n1978), .A3(n1979), .ZN(n1976) );
NOR2_X1 U1562 ( .A1(n1962), .A2(n1980), .ZN(n1979) );
XOR2_X1 U1563 ( .A(n1964), .B(n1981), .Z(n1980) );
NOR3_X1 U1564 ( .A1(n1966), .A2(KEYINPUT49), .A3(n1967), .ZN(n1981) );
NOR2_X1 U1565 ( .A1(n1982), .A2(n1983), .ZN(n1967) );
XOR2_X1 U1566 ( .A(n1961), .B(KEYINPUT33), .Z(n1966) );
NOR2_X1 U1567 ( .A1(n1984), .A2(n1985), .ZN(n1961) );
NOR3_X1 U1568 ( .A1(n1986), .A2(n1987), .A3(n1988), .ZN(n1978) );
NOR3_X1 U1569 ( .A1(n1989), .A2(n1990), .A3(n1950), .ZN(n1987) );
XNOR2_X1 U1570 ( .A(KEYINPUT61), .B(n1951), .ZN(n1986) );
NAND2_X1 U1571 ( .A1(n1990), .A2(n1991), .ZN(n1951) );
OR2_X1 U1572 ( .A1(n1989), .A2(n1950), .ZN(n1991) );
NOR2_X1 U1573 ( .A1(n1992), .A2(n1985), .ZN(n1950) );
NOR2_X1 U1574 ( .A1(n1982), .A2(n1993), .ZN(n1989) );
NOR2_X1 U1575 ( .A1(n1994), .A2(n1995), .ZN(n1977) );
XOR2_X1 U1576 ( .A(REG4_REG_5__SCAN_IN), .B(KEYINPUT29), .Z(n1995) );
INV_X1 U1577 ( .A(n1953), .ZN(n1994) );
NAND2_X1 U1578 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1724), .ZN(n1975) );
NAND2_X1 U1579 ( .A1(n1996), .A2(n1985), .ZN(n1974) );
INV_X1 U1580 ( .A(n1982), .ZN(n1985) );
NAND2_X1 U1581 ( .A1(n1997), .A2(n1998), .ZN(n1982) );
NAND3_X1 U1582 ( .A1(n1999), .A2(n2000), .A3(n2001), .ZN(n1998) );
XOR2_X1 U1583 ( .A(n2002), .B(n2003), .Z(n2001) );
NAND2_X1 U1584 ( .A1(n2004), .A2(n2005), .ZN(n2000) );
NAND3_X1 U1585 ( .A1(n2004), .A2(n2006), .A3(n2007), .ZN(n1997) );
XOR2_X1 U1586 ( .A(n2002), .B(n2008), .Z(n2007) );
NOR2_X1 U1587 ( .A1(KEYINPUT57), .A2(n2003), .ZN(n2008) );
NAND2_X1 U1588 ( .A1(n2009), .A2(n2010), .ZN(n2003) );
NAND2_X1 U1589 ( .A1(DATA_IN_6_), .A2(n2011), .ZN(n2010) );
NAND2_X1 U1590 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2009) );
NAND3_X1 U1591 ( .A1(n2012), .A2(n2013), .A3(n2014), .ZN(n2002) );
OR2_X1 U1592 ( .A1(n2015), .A2(REG4_REG_6__SCAN_IN), .ZN(n2014) );
NAND3_X1 U1593 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2015), .A3(n2011), .ZN(n2013) );
NAND2_X1 U1594 ( .A1(RESTART), .A2(n2016), .ZN(n2012) );
NAND2_X1 U1595 ( .A1(n1817), .A2(n2015), .ZN(n2016) );
INV_X1 U1596 ( .A(KEYINPUT52), .ZN(n2015) );
NAND2_X1 U1597 ( .A1(n2017), .A2(n1999), .ZN(n2006) );
NAND2_X1 U1598 ( .A1(n2018), .A2(n2019), .ZN(n1999) );
INV_X1 U1599 ( .A(n2005), .ZN(n2017) );
NAND2_X1 U1600 ( .A1(n2020), .A2(n2021), .ZN(n2004) );
NAND2_X1 U1601 ( .A1(n1947), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1973) );
NAND4_X1 U1602 ( .A1(n2022), .A2(n2023), .A3(n2024), .A4(n2025), .ZN(U285));
NOR3_X1 U1603 ( .A1(n2026), .A2(n2027), .A3(n2028), .ZN(n2025) );
NOR3_X1 U1604 ( .A1(n1988), .A2(n1990), .A3(n2029), .ZN(n2028) );
NOR2_X1 U1605 ( .A1(n2030), .A2(n2031), .ZN(n2029) );
AND2_X1 U1606 ( .A1(n2030), .A2(n2031), .ZN(n1990) );
NAND2_X1 U1607 ( .A1(n1992), .A2(n2032), .ZN(n2031) );
NAND2_X1 U1608 ( .A1(n2033), .A2(n2034), .ZN(n2032) );
INV_X1 U1609 ( .A(n1993), .ZN(n1992) );
NOR2_X1 U1610 ( .A1(n2033), .A2(n2034), .ZN(n1993) );
NOR3_X1 U1611 ( .A1(n1962), .A2(n1964), .A3(n2035), .ZN(n2027) );
NOR2_X1 U1612 ( .A1(n2036), .A2(n2037), .ZN(n2035) );
AND2_X1 U1613 ( .A1(n2038), .A2(n2039), .ZN(n2036) );
AND3_X1 U1614 ( .A1(n2037), .A2(n2038), .A3(n2039), .ZN(n1964) );
NAND2_X1 U1615 ( .A1(n1984), .A2(n2040), .ZN(n2037) );
NAND2_X1 U1616 ( .A1(n2041), .A2(n2034), .ZN(n2040) );
NAND2_X1 U1617 ( .A1(n2042), .A2(n2043), .ZN(n2041) );
INV_X1 U1618 ( .A(n2044), .ZN(n2042) );
INV_X1 U1619 ( .A(n1983), .ZN(n1984) );
NOR3_X1 U1620 ( .A1(n2045), .A2(n2044), .A3(n2034), .ZN(n1983) );
AND2_X1 U1621 ( .A1(n2034), .A2(n1996), .ZN(n2026) );
NAND2_X1 U1622 ( .A1(n2046), .A2(n2047), .ZN(n2034) );
NAND2_X1 U1623 ( .A1(n2048), .A2(n2005), .ZN(n2047) );
XOR2_X1 U1624 ( .A(KEYINPUT25), .B(n2049), .Z(n2046) );
NOR2_X1 U1625 ( .A1(n2048), .A2(n2005), .ZN(n2049) );
NAND2_X1 U1626 ( .A1(n2050), .A2(n2051), .ZN(n2005) );
NAND2_X1 U1627 ( .A1(n2052), .A2(n2053), .ZN(n2051) );
OR2_X1 U1628 ( .A1(n2054), .A2(n2055), .ZN(n2053) );
NAND2_X1 U1629 ( .A1(n2055), .A2(n2054), .ZN(n2050) );
XOR2_X1 U1630 ( .A(n2018), .B(n2019), .Z(n2048) );
INV_X1 U1631 ( .A(n2020), .ZN(n2019) );
NAND2_X1 U1632 ( .A1(n2056), .A2(n2057), .ZN(n2020) );
NAND2_X1 U1633 ( .A1(DATA_IN_5_), .A2(n2011), .ZN(n2057) );
NAND2_X1 U1634 ( .A1(RESTART), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2056) );
INV_X1 U1635 ( .A(n2021), .ZN(n2018) );
NAND3_X1 U1636 ( .A1(n2058), .A2(n2059), .A3(n2060), .ZN(n2021) );
NAND2_X1 U1637 ( .A1(RESTART), .A2(n2061), .ZN(n2060) );
NAND2_X1 U1638 ( .A1(KEYINPUT18), .A2(n1793), .ZN(n2061) );
NAND3_X1 U1639 ( .A1(KEYINPUT18), .A2(n2011), .A3(REG4_REG_5__SCAN_IN), .ZN(n2059) );
OR2_X1 U1640 ( .A1(KEYINPUT18), .A2(REG4_REG_5__SCAN_IN), .ZN(n2058) );
NAND2_X1 U1641 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1724), .ZN(n2024) );
NAND2_X1 U1642 ( .A1(n1947), .A2(RLAST_REG_4__SCAN_IN), .ZN(n2023) );
NAND2_X1 U1643 ( .A1(n1953), .A2(REG4_REG_4__SCAN_IN), .ZN(n2022) );
NAND4_X1 U1644 ( .A1(n2062), .A2(n2063), .A3(n2064), .A4(n2065), .ZN(U284));
NOR3_X1 U1645 ( .A1(n2066), .A2(n2067), .A3(n2068), .ZN(n2065) );
NOR2_X1 U1646 ( .A1(n1962), .A2(n2069), .ZN(n2068) );
XNOR2_X1 U1647 ( .A(n2039), .B(n2038), .ZN(n2069) );
NAND2_X1 U1648 ( .A1(n2070), .A2(n2071), .ZN(n2038) );
NAND2_X1 U1649 ( .A1(n2043), .A2(n2072), .ZN(n2071) );
XOR2_X1 U1650 ( .A(n2044), .B(n2073), .Z(n2070) );
NOR2_X1 U1651 ( .A1(n2043), .A2(n2072), .ZN(n2073) );
INV_X1 U1652 ( .A(KEYINPUT53), .ZN(n2072) );
NOR3_X1 U1653 ( .A1(n1988), .A2(n2030), .A3(n2074), .ZN(n2067) );
NOR2_X1 U1654 ( .A1(n2075), .A2(n2076), .ZN(n2074) );
AND2_X1 U1655 ( .A1(n2075), .A2(n2076), .ZN(n2030) );
NAND2_X1 U1656 ( .A1(n2033), .A2(n2077), .ZN(n2076) );
NAND2_X1 U1657 ( .A1(n2045), .A2(n2078), .ZN(n2077) );
OR2_X1 U1658 ( .A1(n2078), .A2(n2045), .ZN(n2033) );
NOR2_X1 U1659 ( .A1(n2043), .A2(n2079), .ZN(n2066) );
INV_X1 U1660 ( .A(n2045), .ZN(n2043) );
NAND2_X1 U1661 ( .A1(n2080), .A2(n2081), .ZN(n2045) );
NAND2_X1 U1662 ( .A1(n2082), .A2(n2083), .ZN(n2081) );
NAND2_X1 U1663 ( .A1(n2084), .A2(n2085), .ZN(n2082) );
NAND2_X1 U1664 ( .A1(n2086), .A2(n2087), .ZN(n2085) );
XOR2_X1 U1665 ( .A(n2054), .B(n2052), .Z(n2084) );
NAND3_X1 U1666 ( .A1(n2088), .A2(n2087), .A3(n2055), .ZN(n2080) );
INV_X1 U1667 ( .A(n2083), .ZN(n2055) );
NAND2_X1 U1668 ( .A1(n2089), .A2(n2090), .ZN(n2083) );
NAND2_X1 U1669 ( .A1(n2091), .A2(n2092), .ZN(n2090) );
NAND2_X1 U1670 ( .A1(n2093), .A2(n2094), .ZN(n2092) );
XOR2_X1 U1671 ( .A(n2095), .B(KEYINPUT20), .Z(n2089) );
OR2_X1 U1672 ( .A1(n2094), .A2(n2093), .ZN(n2095) );
NAND2_X1 U1673 ( .A1(n2096), .A2(n2097), .ZN(n2087) );
NAND2_X1 U1674 ( .A1(n2098), .A2(n2054), .ZN(n2097) );
XOR2_X1 U1675 ( .A(KEYINPUT16), .B(n2099), .Z(n2096) );
NOR2_X1 U1676 ( .A1(n2098), .A2(n2054), .ZN(n2099) );
NAND2_X1 U1677 ( .A1(n2100), .A2(n2101), .ZN(n2054) );
NAND2_X1 U1678 ( .A1(RESTART), .A2(n1835), .ZN(n2101) );
NAND2_X1 U1679 ( .A1(n1797), .A2(n2011), .ZN(n2100) );
INV_X1 U1680 ( .A(n2052), .ZN(n2098) );
NAND2_X1 U1681 ( .A1(n2102), .A2(n2103), .ZN(n2052) );
NAND2_X1 U1682 ( .A1(RESTART), .A2(n1814), .ZN(n2103) );
NAND2_X1 U1683 ( .A1(n2104), .A2(n2011), .ZN(n2102) );
INV_X1 U1684 ( .A(n2086), .ZN(n2088) );
XNOR2_X1 U1685 ( .A(KEYINPUT59), .B(KEYINPUT46), .ZN(n2086) );
NAND2_X1 U1686 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1724), .ZN(n2064) );
NAND2_X1 U1687 ( .A1(n1947), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2063) );
NAND2_X1 U1688 ( .A1(n1953), .A2(REG4_REG_3__SCAN_IN), .ZN(n2062) );
NAND4_X1 U1689 ( .A1(n2105), .A2(n2106), .A3(n2107), .A4(n2108), .ZN(U283));
NOR3_X1 U1690 ( .A1(n2109), .A2(n2110), .A3(n2111), .ZN(n2108) );
NOR3_X1 U1691 ( .A1(n1988), .A2(n2075), .A3(n2112), .ZN(n2111) );
NOR2_X1 U1692 ( .A1(n2113), .A2(n2114), .ZN(n2112) );
AND2_X1 U1693 ( .A1(n2115), .A2(n2116), .ZN(n2113) );
AND3_X1 U1694 ( .A1(n2116), .A2(n2115), .A3(n2117), .ZN(n2075) );
XOR2_X1 U1695 ( .A(n2114), .B(KEYINPUT26), .Z(n2117) );
NAND3_X1 U1696 ( .A1(n2118), .A2(n2119), .A3(n2120), .ZN(n2114) );
NAND2_X1 U1697 ( .A1(n2121), .A2(n2122), .ZN(n2120) );
XOR2_X1 U1698 ( .A(KEYINPUT12), .B(n2123), .Z(n2121) );
NAND3_X1 U1699 ( .A1(n2123), .A2(n2124), .A3(n2125), .ZN(n2119) );
OR2_X1 U1700 ( .A1(n2125), .A2(n2078), .ZN(n2118) );
NAND2_X1 U1701 ( .A1(n2124), .A2(n2126), .ZN(n2078) );
XOR2_X1 U1702 ( .A(n2122), .B(KEYINPUT62), .Z(n2124) );
INV_X1 U1703 ( .A(KEYINPUT1), .ZN(n2125) );
NOR3_X1 U1704 ( .A1(n1962), .A2(n2039), .A3(n2127), .ZN(n2110) );
NOR2_X1 U1705 ( .A1(n2128), .A2(n2129), .ZN(n2127) );
NOR2_X1 U1706 ( .A1(n2130), .A2(n2131), .ZN(n2128) );
AND3_X1 U1707 ( .A1(n2132), .A2(n2115), .A3(n2129), .ZN(n2039) );
NAND2_X1 U1708 ( .A1(n2044), .A2(n2133), .ZN(n2129) );
NAND2_X1 U1709 ( .A1(n2123), .A2(n2122), .ZN(n2133) );
INV_X1 U1710 ( .A(n2126), .ZN(n2123) );
NAND2_X1 U1711 ( .A1(n2134), .A2(n2126), .ZN(n2044) );
NOR2_X1 U1712 ( .A1(n2126), .A2(n2079), .ZN(n2109) );
XNOR2_X1 U1713 ( .A(n2135), .B(n2094), .ZN(n2126) );
NAND3_X1 U1714 ( .A1(n2136), .A2(n2137), .A3(n2138), .ZN(n2094) );
NAND2_X1 U1715 ( .A1(n2139), .A2(n1801), .ZN(n2138) );
NAND2_X1 U1716 ( .A1(REG4_REG_3__SCAN_IN), .A2(n2011), .ZN(n2139) );
OR2_X1 U1717 ( .A1(n2011), .A2(KEYINPUT60), .ZN(n2137) );
NAND3_X1 U1718 ( .A1(n2140), .A2(n2011), .A3(KEYINPUT60), .ZN(n2136) );
NAND2_X1 U1719 ( .A1(n2141), .A2(n2142), .ZN(n2135) );
NAND2_X1 U1720 ( .A1(n2093), .A2(n2143), .ZN(n2142) );
NAND2_X1 U1721 ( .A1(n2091), .A2(n2144), .ZN(n2141) );
NAND2_X1 U1722 ( .A1(KEYINPUT37), .A2(n2093), .ZN(n2144) );
AND3_X1 U1723 ( .A1(n2145), .A2(n2146), .A3(n2147), .ZN(n2093) );
NAND2_X1 U1724 ( .A1(KEYINPUT47), .A2(n1813), .ZN(n2147) );
NAND3_X1 U1725 ( .A1(DATA_IN_3_), .A2(n2148), .A3(n2011), .ZN(n2146) );
NAND2_X1 U1726 ( .A1(RESTART), .A2(n2149), .ZN(n2145) );
NAND2_X1 U1727 ( .A1(n2148), .A2(n1848), .ZN(n2149) );
INV_X1 U1728 ( .A(KEYINPUT47), .ZN(n2148) );
INV_X1 U1729 ( .A(n2143), .ZN(n2091) );
NAND2_X1 U1730 ( .A1(n2150), .A2(n2151), .ZN(n2143) );
NAND2_X1 U1731 ( .A1(n2152), .A2(n2153), .ZN(n2151) );
NAND2_X1 U1732 ( .A1(n2154), .A2(n2155), .ZN(n2153) );
NAND2_X1 U1733 ( .A1(n2156), .A2(n2157), .ZN(n2150) );
NAND2_X1 U1734 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1724), .ZN(n2107) );
NAND2_X1 U1735 ( .A1(n1947), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2106) );
NAND2_X1 U1736 ( .A1(n1953), .A2(REG4_REG_2__SCAN_IN), .ZN(n2105) );
NAND4_X1 U1737 ( .A1(n2158), .A2(n2159), .A3(n2160), .A4(n2161), .ZN(U282));
NOR3_X1 U1738 ( .A1(n2162), .A2(n2163), .A3(n2164), .ZN(n2161) );
NOR2_X1 U1739 ( .A1(n2165), .A2(n1962), .ZN(n2164) );
INV_X1 U1740 ( .A(n1963), .ZN(n1962) );
NOR2_X1 U1741 ( .A1(n2166), .A2(n2167), .ZN(n2165) );
XOR2_X1 U1742 ( .A(KEYINPUT22), .B(n2168), .Z(n2167) );
NOR2_X1 U1743 ( .A1(n2130), .A2(n2132), .ZN(n2168) );
NOR2_X1 U1744 ( .A1(n2131), .A2(n2115), .ZN(n2166) );
INV_X1 U1745 ( .A(n2132), .ZN(n2131) );
NAND2_X1 U1746 ( .A1(n2122), .A2(n2169), .ZN(n2132) );
NAND2_X1 U1747 ( .A1(n2170), .A2(n2171), .ZN(n2169) );
NOR2_X1 U1748 ( .A1(n2172), .A2(n1988), .ZN(n2163) );
XOR2_X1 U1749 ( .A(n2116), .B(n2130), .Z(n2172) );
INV_X1 U1750 ( .A(n2115), .ZN(n2130) );
NAND2_X1 U1751 ( .A1(n2122), .A2(n2173), .ZN(n2116) );
NAND2_X1 U1752 ( .A1(n2174), .A2(n2171), .ZN(n2173) );
XOR2_X1 U1753 ( .A(n2170), .B(KEYINPUT0), .Z(n2174) );
INV_X1 U1754 ( .A(n2134), .ZN(n2122) );
NOR2_X1 U1755 ( .A1(n2171), .A2(n2170), .ZN(n2134) );
AND2_X1 U1756 ( .A1(n2170), .A2(n1996), .ZN(n2162) );
NAND2_X1 U1757 ( .A1(n2175), .A2(n2176), .ZN(n2170) );
NAND2_X1 U1758 ( .A1(n2177), .A2(n2157), .ZN(n2176) );
NAND2_X1 U1759 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
OR2_X1 U1760 ( .A1(n2152), .A2(n2155), .ZN(n2179) );
XOR2_X1 U1761 ( .A(n2180), .B(KEYINPUT21), .Z(n2178) );
NAND2_X1 U1762 ( .A1(n2155), .A2(n2181), .ZN(n2180) );
XOR2_X1 U1763 ( .A(n2152), .B(KEYINPUT27), .Z(n2181) );
NAND2_X1 U1764 ( .A1(n2182), .A2(n2154), .ZN(n2175) );
INV_X1 U1765 ( .A(n2157), .ZN(n2154) );
NAND2_X1 U1766 ( .A1(n2183), .A2(n2184), .ZN(n2157) );
NAND2_X1 U1767 ( .A1(n2185), .A2(n2186), .ZN(n2184) );
XOR2_X1 U1768 ( .A(n2152), .B(n2155), .Z(n2182) );
INV_X1 U1769 ( .A(n2156), .ZN(n2155) );
NAND2_X1 U1770 ( .A1(n2187), .A2(n2188), .ZN(n2156) );
NAND2_X1 U1771 ( .A1(RESTART), .A2(n1843), .ZN(n2188) );
NAND2_X1 U1772 ( .A1(n1811), .A2(n2011), .ZN(n2187) );
NAND2_X1 U1773 ( .A1(n2189), .A2(n2190), .ZN(n2152) );
NAND2_X1 U1774 ( .A1(RESTART), .A2(n1812), .ZN(n2190) );
NAND2_X1 U1775 ( .A1(n2191), .A2(n2011), .ZN(n2189) );
NAND2_X1 U1776 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1724), .ZN(n2160) );
NAND2_X1 U1777 ( .A1(n1947), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2159) );
NAND2_X1 U1778 ( .A1(n1953), .A2(REG4_REG_1__SCAN_IN), .ZN(n2158) );
NAND4_X1 U1779 ( .A1(n2192), .A2(n2193), .A3(n2194), .A4(n2195), .ZN(U281));
NAND2_X1 U1780 ( .A1(n1996), .A2(n2196), .ZN(n2195) );
INV_X1 U1781 ( .A(n2079), .ZN(n1996) );
NAND4_X1 U1782 ( .A1(STATO_REG_1__SCAN_IN), .A2(U280), .A3(n2197), .A4(n2198), .ZN(n2079) );
NAND2_X1 U1783 ( .A1(n2199), .A2(n2011), .ZN(n2198) );
NAND3_X1 U1784 ( .A1(n2200), .A2(n2201), .A3(ENABLE), .ZN(n2199) );
INV_X1 U1785 ( .A(AVERAGE), .ZN(n2201) );
NAND2_X1 U1786 ( .A1(n2202), .A2(RESTART), .ZN(n2197) );
NOR2_X1 U1787 ( .A1(n2203), .A2(n2204), .ZN(n2194) );
AND2_X1 U1788 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1947), .ZN(n2204) );
NOR2_X1 U1789 ( .A1(n2205), .A2(ENABLE), .ZN(n1947) );
NOR2_X1 U1790 ( .A1(n2206), .A2(n2115), .ZN(n2203) );
NAND2_X1 U1791 ( .A1(n2171), .A2(n2207), .ZN(n2115) );
NAND2_X1 U1792 ( .A1(n2208), .A2(n2196), .ZN(n2207) );
OR2_X1 U1793 ( .A1(n2196), .A2(n2208), .ZN(n2171) );
NAND2_X1 U1794 ( .A1(n2209), .A2(n2210), .ZN(n2208) );
NAND2_X1 U1795 ( .A1(n2211), .A2(n2212), .ZN(n2210) );
NAND2_X1 U1796 ( .A1(n2213), .A2(n2214), .ZN(n2211) );
NAND2_X1 U1797 ( .A1(KEYINPUT55), .A2(n2215), .ZN(n2214) );
OR2_X1 U1798 ( .A1(n2216), .A2(KEYINPUT55), .ZN(n2213) );
NAND2_X1 U1799 ( .A1(n2217), .A2(n2216), .ZN(n2209) );
NOR2_X1 U1800 ( .A1(n2218), .A2(KEYINPUT38), .ZN(n2216) );
NAND3_X1 U1801 ( .A1(n2219), .A2(n2220), .A3(n2221), .ZN(n2196) );
XOR2_X1 U1802 ( .A(n2222), .B(KEYINPUT30), .Z(n2221) );
OR2_X1 U1803 ( .A1(n2186), .A2(n2185), .ZN(n2222) );
NAND3_X1 U1804 ( .A1(n2185), .A2(n2186), .A3(n2183), .ZN(n2220) );
NAND3_X1 U1805 ( .A1(n2215), .A2(n2223), .A3(n2212), .ZN(n2185) );
INV_X1 U1806 ( .A(n2217), .ZN(n2212) );
OR2_X1 U1807 ( .A1(n2183), .A2(n2186), .ZN(n2219) );
NAND3_X1 U1808 ( .A1(n2224), .A2(n2225), .A3(n2226), .ZN(n2186) );
NAND2_X1 U1809 ( .A1(n2227), .A2(n1847), .ZN(n2226) );
NAND2_X1 U1810 ( .A1(DATA_IN_1_), .A2(n2011), .ZN(n2227) );
OR3_X1 U1811 ( .A1(DATA_IN_1_), .A2(KEYINPUT9), .A3(RESTART), .ZN(n2225) );
NAND2_X1 U1812 ( .A1(KEYINPUT9), .A2(RESTART), .ZN(n2224) );
OR2_X1 U1813 ( .A1(n2223), .A2(n2228), .ZN(n2183) );
NOR2_X1 U1814 ( .A1(n2217), .A2(n2218), .ZN(n2228) );
INV_X1 U1815 ( .A(n2215), .ZN(n2218) );
NAND3_X1 U1816 ( .A1(n2229), .A2(n2230), .A3(n2231), .ZN(n2215) );
NAND2_X1 U1817 ( .A1(KEYINPUT23), .A2(n2232), .ZN(n2231) );
OR3_X1 U1818 ( .A1(n2232), .A2(KEYINPUT23), .A3(n2011), .ZN(n2230) );
INV_X1 U1819 ( .A(RMIN_REG_0__SCAN_IN), .ZN(n2232) );
NAND2_X1 U1820 ( .A1(n2233), .A2(n2011), .ZN(n2229) );
OR2_X1 U1821 ( .A1(REG4_REG_0__SCAN_IN), .A2(KEYINPUT23), .ZN(n2233) );
NAND2_X1 U1822 ( .A1(n2234), .A2(n2235), .ZN(n2217) );
OR2_X1 U1823 ( .A1(n2011), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2235) );
NAND2_X1 U1824 ( .A1(n1808), .A2(n2011), .ZN(n2234) );
INV_X1 U1825 ( .A(DATA_IN_0_), .ZN(n1808) );
NAND3_X1 U1826 ( .A1(n2236), .A2(n2237), .A3(n2238), .ZN(n2223) );
NAND2_X1 U1827 ( .A1(KEYINPUT41), .A2(n2239), .ZN(n2238) );
NAND3_X1 U1828 ( .A1(REG4_REG_1__SCAN_IN), .A2(n2240), .A3(n2011), .ZN(n2237) );
NAND2_X1 U1829 ( .A1(RESTART), .A2(n2241), .ZN(n2236) );
NAND2_X1 U1830 ( .A1(n2242), .A2(n2240), .ZN(n2241) );
INV_X1 U1831 ( .A(KEYINPUT41), .ZN(n2240) );
NOR2_X1 U1832 ( .A1(n1963), .A2(n1952), .ZN(n2206) );
INV_X1 U1833 ( .A(n1988), .ZN(n1952) );
NAND4_X1 U1834 ( .A1(n2202), .A2(RESTART), .A3(STATO_REG_1__SCAN_IN), .A4(
U280), .ZN(n1988) );
XOR2_X1 U1835 ( .A(n2243), .B(KEYINPUT40), .Z(n2202) );
NAND2_X1 U1836 ( .A1(n2244), .A2(n2245), .ZN(n2243) );
NAND2_X1 U1837 ( .A1(n2246), .A2(n2247), .ZN(n2245) );
NAND2_X1 U1838 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2247) );
NAND2_X1 U1839 ( .A1(n2248), .A2(n2249), .ZN(n2246) );
NAND2_X1 U1840 ( .A1(RMIN_REG_6__SCAN_IN), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2249) );
NAND3_X1 U1841 ( .A1(n2250), .A2(n2251), .A3(n2252), .ZN(n2248) );
NAND2_X1 U1842 ( .A1(n1828), .A2(n1817), .ZN(n2252) );
INV_X1 U1843 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1817) );
INV_X1 U1844 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1828) );
NAND3_X1 U1845 ( .A1(n2253), .A2(n2254), .A3(n2255), .ZN(n2251) );
NAND2_X1 U1846 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2255) );
NAND3_X1 U1847 ( .A1(n2256), .A2(n2257), .A3(n2258), .ZN(n2254) );
NAND2_X1 U1848 ( .A1(n1835), .A2(n1814), .ZN(n2258) );
INV_X1 U1849 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1814) );
INV_X1 U1850 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1835) );
NAND3_X1 U1851 ( .A1(n2259), .A2(n2260), .A3(n2261), .ZN(n2257) );
NAND2_X1 U1852 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2261) );
NAND3_X1 U1853 ( .A1(n2262), .A2(n2263), .A3(n2264), .ZN(n2260) );
NAND2_X1 U1854 ( .A1(n1843), .A2(n1812), .ZN(n2264) );
INV_X1 U1855 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1812) );
INV_X1 U1856 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1843) );
NAND2_X1 U1857 ( .A1(n2265), .A2(n2266), .ZN(n2263) );
NAND2_X1 U1858 ( .A1(RMIN_REG_1__SCAN_IN), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2266) );
NAND2_X1 U1859 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2265) );
NAND2_X1 U1860 ( .A1(n1847), .A2(n2242), .ZN(n2262) );
INV_X1 U1861 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n2242) );
INV_X1 U1862 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1847) );
NAND2_X1 U1863 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2259) );
NAND2_X1 U1864 ( .A1(n1848), .A2(n1801), .ZN(n2256) );
INV_X1 U1865 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1801) );
INV_X1 U1866 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1848) );
NAND2_X1 U1867 ( .A1(n2267), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2253) );
XOR2_X1 U1868 ( .A(n1850), .B(KEYINPUT42), .Z(n2267) );
NAND2_X1 U1869 ( .A1(n1850), .A2(n1793), .ZN(n2250) );
INV_X1 U1870 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1793) );
INV_X1 U1871 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1850) );
NAND2_X1 U1872 ( .A1(n1824), .A2(n1818), .ZN(n2244) );
INV_X1 U1873 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1818) );
INV_X1 U1874 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1824) );
NOR4_X1 U1875 ( .A1(n1872), .A2(n2205), .A3(n2200), .A4(AVERAGE), .ZN(n1963));
NAND2_X1 U1876 ( .A1(n2268), .A2(n2269), .ZN(n2200) );
NAND2_X1 U1877 ( .A1(n2270), .A2(n2271), .ZN(n2269) );
INV_X1 U1878 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2271) );
OR2_X1 U1879 ( .A1(n2272), .A2(n1784), .ZN(n2270) );
NAND2_X1 U1880 ( .A1(n2272), .A2(n1784), .ZN(n2268) );
INV_X1 U1881 ( .A(DATA_IN_7_), .ZN(n1784) );
NAND2_X1 U1882 ( .A1(n2273), .A2(n2274), .ZN(n2272) );
NAND2_X1 U1883 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2275), .ZN(n2274) );
OR2_X1 U1884 ( .A1(n2276), .A2(DATA_IN_6_), .ZN(n2275) );
NAND2_X1 U1885 ( .A1(DATA_IN_6_), .A2(n2276), .ZN(n2273) );
NAND2_X1 U1886 ( .A1(n2277), .A2(n2278), .ZN(n2276) );
NAND2_X1 U1887 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2278) );
XOR2_X1 U1888 ( .A(n2279), .B(KEYINPUT6), .Z(n2277) );
NAND2_X1 U1889 ( .A1(n2280), .A2(n2281), .ZN(n2279) );
NAND2_X1 U1890 ( .A1(n2282), .A2(n2283), .ZN(n2281) );
NAND3_X1 U1891 ( .A1(n2284), .A2(n2285), .A3(n2286), .ZN(n2283) );
NAND2_X1 U1892 ( .A1(n1797), .A2(n2104), .ZN(n2286) );
INV_X1 U1893 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2104) );
INV_X1 U1894 ( .A(DATA_IN_4_), .ZN(n1797) );
NAND3_X1 U1895 ( .A1(n2287), .A2(n2288), .A3(n2289), .ZN(n2285) );
NAND2_X1 U1896 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2289) );
NAND3_X1 U1897 ( .A1(n2290), .A2(n2291), .A3(n2292), .ZN(n2288) );
NAND2_X1 U1898 ( .A1(n1811), .A2(n2191), .ZN(n2292) );
INV_X1 U1899 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2191) );
INV_X1 U1900 ( .A(DATA_IN_2_), .ZN(n1811) );
NAND2_X1 U1901 ( .A1(n2293), .A2(n2294), .ZN(n2291) );
NAND2_X1 U1902 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2294) );
XOR2_X1 U1903 ( .A(n2295), .B(KEYINPUT39), .Z(n2293) );
NAND2_X1 U1904 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2295) );
NAND2_X1 U1905 ( .A1(n1809), .A2(n2239), .ZN(n2290) );
INV_X1 U1906 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2239) );
INV_X1 U1907 ( .A(DATA_IN_1_), .ZN(n1809) );
NAND2_X1 U1908 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2287) );
NAND2_X1 U1909 ( .A1(n1813), .A2(n2140), .ZN(n2284) );
INV_X1 U1910 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2140) );
INV_X1 U1911 ( .A(DATA_IN_3_), .ZN(n1813) );
NAND2_X1 U1912 ( .A1(DATA_IN_4_), .A2(n2296), .ZN(n2282) );
XOR2_X1 U1913 ( .A(REG4_REG_4__SCAN_IN), .B(KEYINPUT31), .Z(n2296) );
OR2_X1 U1914 ( .A1(DATA_IN_5_), .A2(REG4_REG_5__SCAN_IN), .ZN(n2280) );
NAND2_X1 U1915 ( .A1(n1953), .A2(REG4_REG_0__SCAN_IN), .ZN(n2193) );
XOR2_X1 U1916 ( .A(AVERAGE), .B(KEYINPUT48), .Z(n2297) );
NAND3_X1 U1917 ( .A1(U280), .A2(n2011), .A3(STATO_REG_1__SCAN_IN), .ZN(n2205) );
INV_X1 U1918 ( .A(RESTART), .ZN(n2011) );
INV_X1 U1919 ( .A(ENABLE), .ZN(n1872) );
NAND2_X1 U1920 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1724), .ZN(n2192) );
INV_X1 U1921 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1873) );
NOR2_X1 U1922 ( .A1(n1752), .A2(STATO_REG_1__SCAN_IN), .ZN(n2298) );
INV_X1 U1923 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1752) );
endmodule


