//Key = 1111000101000110000000100001001111011010001110100101101001111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372;

XOR2_X1 U752 ( .A(G107), .B(n1041), .Z(G9) );
NOR2_X1 U753 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1044), .A2(n1045), .A3(G953), .A4(n1046), .ZN(n1043) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U762 ( .A(n1061), .ZN(n1060) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1057) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1053) );
NOR2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR3_X1 U769 ( .A1(n1071), .A2(n1074), .A3(n1056), .ZN(n1049) );
NAND3_X1 U770 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1044) );
XOR2_X1 U771 ( .A(n1078), .B(KEYINPUT6), .Z(n1077) );
NAND4_X1 U772 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1078) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1056), .ZN(n1081) );
INV_X1 U774 ( .A(n1048), .ZN(n1080) );
XOR2_X1 U775 ( .A(n1084), .B(KEYINPUT22), .Z(n1075) );
NOR3_X1 U776 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1042) );
AND4_X1 U777 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1046) );
NOR4_X1 U778 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1088) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U780 ( .A(n1095), .B(KEYINPUT14), .Z(n1089) );
NAND2_X1 U781 ( .A1(G469), .A2(n1096), .ZN(n1095) );
NOR3_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1079), .ZN(n1087) );
NOR2_X1 U783 ( .A1(G469), .A2(n1096), .ZN(n1097) );
XOR2_X1 U784 ( .A(n1099), .B(n1100), .Z(n1086) );
NOR2_X1 U785 ( .A1(G478), .A2(KEYINPUT16), .ZN(n1100) );
XOR2_X1 U786 ( .A(n1101), .B(n1102), .Z(n1085) );
NOR2_X1 U787 ( .A1(n1103), .A2(KEYINPUT61), .ZN(n1102) );
XOR2_X1 U788 ( .A(n1104), .B(n1105), .Z(G72) );
NOR2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
AND2_X1 U790 ( .A1(G227), .A2(G900), .ZN(n1106) );
NOR2_X1 U791 ( .A1(KEYINPUT19), .A2(n1108), .ZN(n1104) );
XOR2_X1 U792 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U793 ( .A1(n1111), .A2(KEYINPUT24), .ZN(n1110) );
NOR2_X1 U794 ( .A1(G953), .A2(n1112), .ZN(n1111) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1114) );
XNOR2_X1 U797 ( .A(n1117), .B(KEYINPUT60), .ZN(n1116) );
NAND2_X1 U798 ( .A1(KEYINPUT52), .A2(n1118), .ZN(n1117) );
XOR2_X1 U799 ( .A(n1119), .B(n1120), .Z(n1115) );
NOR2_X1 U800 ( .A1(G900), .A2(n1107), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(G69) );
NOR2_X1 U802 ( .A1(n1123), .A2(n1107), .ZN(n1122) );
AND2_X1 U803 ( .A1(G224), .A2(G898), .ZN(n1123) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
NAND2_X1 U805 ( .A1(n1126), .A2(n1107), .ZN(n1125) );
XOR2_X1 U806 ( .A(n1076), .B(n1127), .Z(n1126) );
OR3_X1 U807 ( .A1(n1128), .A2(n1127), .A3(n1107), .ZN(n1124) );
XNOR2_X1 U808 ( .A(n1129), .B(KEYINPUT53), .ZN(n1127) );
NOR3_X1 U809 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1133), .A2(G953), .A3(G952), .ZN(n1132) );
INV_X1 U811 ( .A(KEYINPUT45), .ZN(n1133) );
NOR2_X1 U812 ( .A1(KEYINPUT45), .A2(n1134), .ZN(n1131) );
XOR2_X1 U813 ( .A(n1135), .B(n1136), .Z(n1130) );
NAND2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(G63) );
NOR3_X1 U816 ( .A1(n1099), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR3_X1 U817 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
NOR2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
NOR2_X1 U819 ( .A1(n1148), .A2(n1145), .ZN(n1147) );
INV_X1 U820 ( .A(G478), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1084), .A2(n1149), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1139), .A2(n1150), .ZN(G60) );
XOR2_X1 U823 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U824 ( .A1(n1137), .A2(G475), .ZN(n1151) );
XNOR2_X1 U825 ( .A(G104), .B(n1153), .ZN(G6) );
NOR2_X1 U826 ( .A1(n1139), .A2(n1154), .ZN(G57) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U828 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U829 ( .A1(n1137), .A2(G472), .ZN(n1157) );
XOR2_X1 U830 ( .A(n1159), .B(n1160), .Z(n1155) );
XOR2_X1 U831 ( .A(G101), .B(n1161), .Z(n1160) );
NAND2_X1 U832 ( .A1(n1162), .A2(n1163), .ZN(n1159) );
NAND2_X1 U833 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U834 ( .A1(KEYINPUT42), .A2(n1166), .ZN(n1165) );
NAND2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1162) );
NAND2_X1 U837 ( .A1(n1168), .A2(n1171), .ZN(n1170) );
NAND2_X1 U838 ( .A1(KEYINPUT42), .A2(n1172), .ZN(n1171) );
INV_X1 U839 ( .A(n1164), .ZN(n1172) );
XOR2_X1 U840 ( .A(n1118), .B(KEYINPUT54), .Z(n1164) );
INV_X1 U841 ( .A(KEYINPUT41), .ZN(n1168) );
NOR3_X1 U842 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(G54) );
AND3_X1 U843 ( .A1(KEYINPUT39), .A2(G953), .A3(G952), .ZN(n1175) );
NOR2_X1 U844 ( .A1(KEYINPUT39), .A2(n1134), .ZN(n1174) );
INV_X1 U845 ( .A(n1139), .ZN(n1134) );
XOR2_X1 U846 ( .A(n1176), .B(n1177), .Z(n1173) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(n1177) );
NAND2_X1 U848 ( .A1(n1137), .A2(G469), .ZN(n1178) );
XOR2_X1 U849 ( .A(n1180), .B(n1181), .Z(n1176) );
NOR2_X1 U850 ( .A1(G110), .A2(KEYINPUT10), .ZN(n1181) );
NOR2_X1 U851 ( .A1(n1139), .A2(n1182), .ZN(G51) );
XOR2_X1 U852 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U853 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND2_X1 U854 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U855 ( .A1(n1137), .A2(n1101), .ZN(n1185) );
INV_X1 U856 ( .A(n1144), .ZN(n1137) );
NAND2_X1 U857 ( .A1(G902), .A2(n1189), .ZN(n1144) );
NAND2_X1 U858 ( .A1(n1076), .A2(n1112), .ZN(n1189) );
INV_X1 U859 ( .A(n1084), .ZN(n1112) );
NAND4_X1 U860 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1084) );
AND4_X1 U861 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NOR2_X1 U862 ( .A1(n1198), .A2(n1199), .ZN(n1192) );
NOR4_X1 U863 ( .A1(n1200), .A2(n1201), .A3(n1052), .A4(n1202), .ZN(n1199) );
NAND3_X1 U864 ( .A1(n1072), .A2(n1067), .A3(n1063), .ZN(n1201) );
INV_X1 U865 ( .A(KEYINPUT55), .ZN(n1200) );
NOR2_X1 U866 ( .A1(KEYINPUT55), .A2(n1203), .ZN(n1198) );
NAND3_X1 U867 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1190) );
NAND2_X1 U868 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
INV_X1 U869 ( .A(n1149), .ZN(n1076) );
NAND4_X1 U870 ( .A1(n1209), .A2(n1153), .A3(n1210), .A4(n1211), .ZN(n1149) );
NOR4_X1 U871 ( .A1(n1212), .A2(n1041), .A3(n1213), .A4(n1214), .ZN(n1211) );
AND3_X1 U872 ( .A1(n1215), .A2(n1216), .A3(n1072), .ZN(n1041) );
NOR3_X1 U873 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1210) );
NOR2_X1 U874 ( .A1(n1074), .A2(n1220), .ZN(n1219) );
XNOR2_X1 U875 ( .A(KEYINPUT58), .B(n1221), .ZN(n1220) );
NOR4_X1 U876 ( .A1(n1204), .A2(n1222), .A3(n1071), .A4(n1223), .ZN(n1218) );
INV_X1 U877 ( .A(KEYINPUT12), .ZN(n1223) );
NAND3_X1 U878 ( .A1(n1224), .A2(n1225), .A3(n1090), .ZN(n1222) );
NOR2_X1 U879 ( .A1(KEYINPUT12), .A2(n1226), .ZN(n1217) );
NAND3_X1 U880 ( .A1(n1215), .A2(n1216), .A3(n1073), .ZN(n1153) );
NAND3_X1 U881 ( .A1(n1215), .A2(n1227), .A3(n1228), .ZN(n1209) );
XOR2_X1 U882 ( .A(KEYINPUT56), .B(n1063), .Z(n1227) );
NOR2_X1 U883 ( .A1(n1107), .A2(G952), .ZN(n1139) );
NAND2_X1 U884 ( .A1(n1229), .A2(n1230), .ZN(G48) );
NAND2_X1 U885 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U886 ( .A(KEYINPUT30), .B(n1233), .Z(n1229) );
NOR2_X1 U887 ( .A1(n1231), .A2(n1232), .ZN(n1233) );
AND3_X1 U888 ( .A1(n1234), .A2(n1204), .A3(n1235), .ZN(n1231) );
XNOR2_X1 U889 ( .A(n1206), .B(KEYINPUT9), .ZN(n1235) );
XOR2_X1 U890 ( .A(n1236), .B(n1191), .Z(G45) );
NAND4_X1 U891 ( .A1(n1237), .A2(n1204), .A3(n1224), .A4(n1090), .ZN(n1191) );
NAND2_X1 U892 ( .A1(n1238), .A2(n1239), .ZN(G42) );
NAND2_X1 U893 ( .A1(G140), .A2(n1240), .ZN(n1239) );
NAND2_X1 U894 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
OR2_X1 U895 ( .A1(KEYINPUT11), .A2(KEYINPUT49), .ZN(n1242) );
NAND3_X1 U896 ( .A1(n1243), .A2(n1244), .A3(KEYINPUT49), .ZN(n1238) );
OR2_X1 U897 ( .A1(n1241), .A2(KEYINPUT11), .ZN(n1244) );
NAND2_X1 U898 ( .A1(n1241), .A2(n1245), .ZN(n1243) );
OR2_X1 U899 ( .A1(G140), .A2(KEYINPUT11), .ZN(n1245) );
INV_X1 U900 ( .A(n1197), .ZN(n1241) );
NAND3_X1 U901 ( .A1(n1246), .A2(n1062), .A3(n1234), .ZN(n1197) );
XNOR2_X1 U902 ( .A(G137), .B(n1196), .ZN(G39) );
NAND4_X1 U903 ( .A1(n1067), .A2(n1202), .A3(n1206), .A4(n1247), .ZN(n1196) );
NOR2_X1 U904 ( .A1(n1056), .A2(n1052), .ZN(n1247) );
INV_X1 U905 ( .A(n1246), .ZN(n1052) );
INV_X1 U906 ( .A(n1228), .ZN(n1056) );
XNOR2_X1 U907 ( .A(G134), .B(n1203), .ZN(G36) );
NAND3_X1 U908 ( .A1(n1246), .A2(n1072), .A3(n1237), .ZN(n1203) );
AND3_X1 U909 ( .A1(n1067), .A2(n1202), .A3(n1063), .ZN(n1237) );
XNOR2_X1 U910 ( .A(G131), .B(n1195), .ZN(G33) );
NAND3_X1 U911 ( .A1(n1246), .A2(n1063), .A3(n1234), .ZN(n1195) );
INV_X1 U912 ( .A(n1207), .ZN(n1234) );
NAND3_X1 U913 ( .A1(n1067), .A2(n1202), .A3(n1073), .ZN(n1207) );
XOR2_X1 U914 ( .A(n1248), .B(KEYINPUT62), .Z(n1067) );
NOR2_X1 U915 ( .A1(n1083), .A2(n1079), .ZN(n1246) );
INV_X1 U916 ( .A(n1249), .ZN(n1079) );
XOR2_X1 U917 ( .A(G128), .B(n1250), .Z(G30) );
NOR3_X1 U918 ( .A1(n1208), .A2(n1251), .A3(n1074), .ZN(n1250) );
XNOR2_X1 U919 ( .A(n1206), .B(KEYINPUT21), .ZN(n1251) );
NAND3_X1 U920 ( .A1(n1248), .A2(n1202), .A3(n1072), .ZN(n1208) );
XOR2_X1 U921 ( .A(n1252), .B(G101), .Z(G3) );
NAND2_X1 U922 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND3_X1 U923 ( .A1(n1204), .A2(n1255), .A3(n1256), .ZN(n1254) );
INV_X1 U924 ( .A(KEYINPUT7), .ZN(n1256) );
NAND4_X1 U925 ( .A1(n1063), .A2(n1228), .A3(n1248), .A4(n1225), .ZN(n1255) );
NAND4_X1 U926 ( .A1(n1228), .A2(n1215), .A3(n1063), .A4(KEYINPUT7), .ZN(n1253) );
XNOR2_X1 U927 ( .A(G125), .B(n1194), .ZN(G27) );
NAND4_X1 U928 ( .A1(n1073), .A2(n1062), .A3(n1257), .A4(n1061), .ZN(n1194) );
AND2_X1 U929 ( .A1(n1202), .A2(n1204), .ZN(n1257) );
NAND2_X1 U930 ( .A1(n1048), .A2(n1258), .ZN(n1202) );
NAND4_X1 U931 ( .A1(G953), .A2(G902), .A3(n1259), .A4(n1260), .ZN(n1258) );
INV_X1 U932 ( .A(G900), .ZN(n1260) );
XNOR2_X1 U933 ( .A(G122), .B(n1226), .ZN(G24) );
NAND4_X1 U934 ( .A1(n1082), .A2(n1261), .A3(n1224), .A4(n1090), .ZN(n1226) );
INV_X1 U935 ( .A(n1071), .ZN(n1082) );
NAND2_X1 U936 ( .A1(n1061), .A2(n1216), .ZN(n1071) );
INV_X1 U937 ( .A(n1065), .ZN(n1216) );
NAND2_X1 U938 ( .A1(n1262), .A2(n1263), .ZN(n1065) );
XOR2_X1 U939 ( .A(KEYINPUT29), .B(n1264), .Z(n1262) );
NAND2_X1 U940 ( .A1(n1265), .A2(n1266), .ZN(G21) );
NAND2_X1 U941 ( .A1(n1212), .A2(n1267), .ZN(n1266) );
XOR2_X1 U942 ( .A(KEYINPUT13), .B(n1268), .Z(n1265) );
NOR2_X1 U943 ( .A1(n1212), .A2(n1267), .ZN(n1268) );
AND4_X1 U944 ( .A1(n1228), .A2(n1061), .A3(n1206), .A4(n1261), .ZN(n1212) );
AND2_X1 U945 ( .A1(n1269), .A2(n1091), .ZN(n1206) );
XOR2_X1 U946 ( .A(G116), .B(n1270), .Z(G18) );
NOR2_X1 U947 ( .A1(n1074), .A2(n1221), .ZN(n1270) );
NAND4_X1 U948 ( .A1(n1063), .A2(n1061), .A3(n1072), .A4(n1225), .ZN(n1221) );
AND2_X1 U949 ( .A1(n1271), .A2(n1224), .ZN(n1072) );
XOR2_X1 U950 ( .A(G113), .B(n1214), .Z(G15) );
AND4_X1 U951 ( .A1(n1063), .A2(n1073), .A3(n1061), .A4(n1261), .ZN(n1214) );
NOR2_X1 U952 ( .A1(n1068), .A2(n1098), .ZN(n1061) );
INV_X1 U953 ( .A(n1069), .ZN(n1098) );
NOR2_X1 U954 ( .A1(n1224), .A2(n1271), .ZN(n1073) );
AND2_X1 U955 ( .A1(n1269), .A2(n1264), .ZN(n1063) );
XOR2_X1 U956 ( .A(n1091), .B(KEYINPUT27), .Z(n1264) );
XOR2_X1 U957 ( .A(G110), .B(n1213), .Z(G12) );
AND3_X1 U958 ( .A1(n1228), .A2(n1215), .A3(n1062), .ZN(n1213) );
AND2_X1 U959 ( .A1(n1091), .A2(n1263), .ZN(n1062) );
INV_X1 U960 ( .A(n1269), .ZN(n1263) );
XNOR2_X1 U961 ( .A(n1272), .B(n1094), .ZN(n1269) );
NAND2_X1 U962 ( .A1(n1273), .A2(n1274), .ZN(n1094) );
XNOR2_X1 U963 ( .A(n1158), .B(n1275), .ZN(n1273) );
XNOR2_X1 U964 ( .A(n1276), .B(n1277), .ZN(n1275) );
NAND3_X1 U965 ( .A1(KEYINPUT35), .A2(n1278), .A3(n1279), .ZN(n1277) );
XOR2_X1 U966 ( .A(n1280), .B(KEYINPUT40), .Z(n1279) );
OR2_X1 U967 ( .A1(G101), .A2(n1161), .ZN(n1280) );
NAND2_X1 U968 ( .A1(n1161), .A2(G101), .ZN(n1278) );
AND3_X1 U969 ( .A1(n1281), .A2(n1107), .A3(G210), .ZN(n1161) );
NAND2_X1 U970 ( .A1(n1282), .A2(KEYINPUT51), .ZN(n1276) );
XOR2_X1 U971 ( .A(n1169), .B(n1283), .Z(n1282) );
XNOR2_X1 U972 ( .A(n1284), .B(n1285), .ZN(n1158) );
XOR2_X1 U973 ( .A(KEYINPUT0), .B(G119), .Z(n1285) );
XNOR2_X1 U974 ( .A(n1286), .B(n1287), .ZN(n1284) );
NOR2_X1 U975 ( .A1(KEYINPUT25), .A2(n1288), .ZN(n1287) );
NAND2_X1 U976 ( .A1(KEYINPUT36), .A2(n1093), .ZN(n1272) );
INV_X1 U977 ( .A(G472), .ZN(n1093) );
XNOR2_X1 U978 ( .A(n1289), .B(n1138), .ZN(n1091) );
AND2_X1 U979 ( .A1(G217), .A2(n1290), .ZN(n1138) );
NAND2_X1 U980 ( .A1(n1274), .A2(n1135), .ZN(n1289) );
NAND2_X1 U981 ( .A1(n1291), .A2(n1292), .ZN(n1135) );
NAND3_X1 U982 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1292) );
XNOR2_X1 U983 ( .A(n1296), .B(n1297), .ZN(n1293) );
NAND2_X1 U984 ( .A1(n1298), .A2(n1299), .ZN(n1291) );
NAND2_X1 U985 ( .A1(n1295), .A2(n1294), .ZN(n1299) );
NAND2_X1 U986 ( .A1(n1300), .A2(n1301), .ZN(n1294) );
XNOR2_X1 U987 ( .A(n1302), .B(n1303), .ZN(n1301) );
XOR2_X1 U988 ( .A(n1304), .B(KEYINPUT26), .Z(n1295) );
NAND2_X1 U989 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
INV_X1 U990 ( .A(n1300), .ZN(n1306) );
XNOR2_X1 U991 ( .A(n1120), .B(n1307), .ZN(n1300) );
XOR2_X1 U992 ( .A(KEYINPUT33), .B(G146), .Z(n1307) );
XOR2_X1 U993 ( .A(G125), .B(n1308), .Z(n1120) );
XOR2_X1 U994 ( .A(n1302), .B(n1303), .Z(n1305) );
XOR2_X1 U995 ( .A(G110), .B(G128), .Z(n1303) );
NAND2_X1 U996 ( .A1(KEYINPUT46), .A2(n1267), .ZN(n1302) );
XOR2_X1 U997 ( .A(n1296), .B(n1297), .Z(n1298) );
NAND2_X1 U998 ( .A1(KEYINPUT1), .A2(n1309), .ZN(n1297) );
NAND3_X1 U999 ( .A1(G234), .A2(n1107), .A3(G221), .ZN(n1296) );
AND2_X1 U1000 ( .A1(n1248), .A2(n1261), .ZN(n1215) );
AND2_X1 U1001 ( .A1(n1204), .A2(n1225), .ZN(n1261) );
NAND2_X1 U1002 ( .A1(n1048), .A2(n1310), .ZN(n1225) );
NAND4_X1 U1003 ( .A1(G953), .A2(G902), .A3(n1311), .A4(n1128), .ZN(n1310) );
INV_X1 U1004 ( .A(G898), .ZN(n1128) );
XNOR2_X1 U1005 ( .A(KEYINPUT43), .B(n1259), .ZN(n1311) );
NAND3_X1 U1006 ( .A1(n1259), .A2(n1107), .A3(G952), .ZN(n1048) );
NAND2_X1 U1007 ( .A1(G237), .A2(G234), .ZN(n1259) );
INV_X1 U1008 ( .A(n1074), .ZN(n1204) );
NAND2_X1 U1009 ( .A1(n1083), .A2(n1249), .ZN(n1074) );
NAND2_X1 U1010 ( .A1(n1312), .A2(n1313), .ZN(n1249) );
XNOR2_X1 U1011 ( .A(G214), .B(KEYINPUT31), .ZN(n1312) );
XOR2_X1 U1012 ( .A(n1314), .B(n1101), .Z(n1083) );
AND2_X1 U1013 ( .A1(G210), .A2(n1313), .ZN(n1101) );
NAND2_X1 U1014 ( .A1(n1281), .A2(n1274), .ZN(n1313) );
XNOR2_X1 U1015 ( .A(n1103), .B(KEYINPUT3), .ZN(n1314) );
AND2_X1 U1016 ( .A1(n1315), .A2(n1274), .ZN(n1103) );
XOR2_X1 U1017 ( .A(n1316), .B(n1183), .Z(n1315) );
INV_X1 U1018 ( .A(n1129), .ZN(n1183) );
XOR2_X1 U1019 ( .A(n1317), .B(n1318), .Z(n1129) );
XOR2_X1 U1020 ( .A(G122), .B(G110), .Z(n1318) );
XOR2_X1 U1021 ( .A(n1319), .B(n1320), .Z(n1317) );
NAND2_X1 U1022 ( .A1(n1321), .A2(n1322), .ZN(n1319) );
NAND2_X1 U1023 ( .A1(n1323), .A2(n1286), .ZN(n1322) );
XOR2_X1 U1024 ( .A(n1324), .B(KEYINPUT47), .Z(n1321) );
OR2_X1 U1025 ( .A1(n1286), .A2(n1323), .ZN(n1324) );
XNOR2_X1 U1026 ( .A(n1267), .B(n1288), .ZN(n1323) );
INV_X1 U1027 ( .A(G119), .ZN(n1267) );
XOR2_X1 U1028 ( .A(G113), .B(KEYINPUT15), .Z(n1286) );
XOR2_X1 U1029 ( .A(n1325), .B(KEYINPUT28), .Z(n1316) );
NAND2_X1 U1030 ( .A1(n1326), .A2(n1188), .ZN(n1325) );
NAND3_X1 U1031 ( .A1(n1327), .A2(n1107), .A3(G224), .ZN(n1188) );
XOR2_X1 U1032 ( .A(G125), .B(n1167), .Z(n1327) );
INV_X1 U1033 ( .A(n1169), .ZN(n1167) );
XOR2_X1 U1034 ( .A(n1187), .B(KEYINPUT8), .Z(n1326) );
NAND2_X1 U1035 ( .A1(n1328), .A2(n1329), .ZN(n1187) );
NAND2_X1 U1036 ( .A1(G224), .A2(n1107), .ZN(n1329) );
XOR2_X1 U1037 ( .A(n1169), .B(G125), .Z(n1328) );
XNOR2_X1 U1038 ( .A(n1330), .B(n1331), .ZN(n1169) );
NOR2_X1 U1039 ( .A1(KEYINPUT4), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1040 ( .A(n1236), .B(KEYINPUT44), .Z(n1332) );
AND2_X1 U1041 ( .A1(n1068), .A2(n1069), .ZN(n1248) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1290), .ZN(n1069) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1274), .ZN(n1290) );
XOR2_X1 U1044 ( .A(n1096), .B(n1333), .Z(n1068) );
NOR2_X1 U1045 ( .A1(G469), .A2(KEYINPUT5), .ZN(n1333) );
NAND2_X1 U1046 ( .A1(n1334), .A2(n1274), .ZN(n1096) );
XOR2_X1 U1047 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1048 ( .A(G110), .B(n1179), .ZN(n1336) );
XOR2_X1 U1049 ( .A(n1337), .B(n1338), .Z(n1179) );
XOR2_X1 U1050 ( .A(n1283), .B(n1308), .Z(n1338) );
INV_X1 U1051 ( .A(n1118), .ZN(n1283) );
XNOR2_X1 U1052 ( .A(G131), .B(n1339), .ZN(n1118) );
XNOR2_X1 U1053 ( .A(n1309), .B(G134), .ZN(n1339) );
INV_X1 U1054 ( .A(G137), .ZN(n1309) );
XOR2_X1 U1055 ( .A(n1119), .B(n1320), .Z(n1337) );
XNOR2_X1 U1056 ( .A(n1340), .B(n1341), .ZN(n1320) );
XOR2_X1 U1057 ( .A(KEYINPUT48), .B(G107), .Z(n1341) );
XNOR2_X1 U1058 ( .A(G104), .B(G101), .ZN(n1340) );
XOR2_X1 U1059 ( .A(n1342), .B(n1343), .Z(n1119) );
XOR2_X1 U1060 ( .A(KEYINPUT2), .B(n1344), .Z(n1343) );
XOR2_X1 U1061 ( .A(KEYINPUT63), .B(KEYINPUT32), .Z(n1344) );
XOR2_X1 U1062 ( .A(n1236), .B(n1330), .Z(n1342) );
XOR2_X1 U1063 ( .A(G128), .B(G146), .Z(n1330) );
NOR2_X1 U1064 ( .A1(n1345), .A2(n1346), .ZN(n1335) );
NOR2_X1 U1065 ( .A1(KEYINPUT57), .A2(n1347), .ZN(n1346) );
INV_X1 U1066 ( .A(n1180), .ZN(n1347) );
NOR2_X1 U1067 ( .A1(KEYINPUT50), .A2(n1180), .ZN(n1345) );
NAND2_X1 U1068 ( .A1(G227), .A2(n1107), .ZN(n1180) );
NOR2_X1 U1069 ( .A1(n1090), .A2(n1224), .ZN(n1228) );
XNOR2_X1 U1070 ( .A(n1099), .B(n1348), .ZN(n1224) );
NOR2_X1 U1071 ( .A1(G478), .A2(KEYINPUT23), .ZN(n1348) );
NOR2_X1 U1072 ( .A1(n1146), .A2(G902), .ZN(n1099) );
INV_X1 U1073 ( .A(n1143), .ZN(n1146) );
NAND2_X1 U1074 ( .A1(n1349), .A2(n1350), .ZN(n1143) );
OR2_X1 U1075 ( .A1(n1351), .A2(KEYINPUT59), .ZN(n1350) );
XOR2_X1 U1076 ( .A(n1352), .B(n1353), .Z(n1349) );
AND3_X1 U1077 ( .A1(G234), .A2(n1107), .A3(G217), .ZN(n1353) );
NAND2_X1 U1078 ( .A1(KEYINPUT59), .A2(n1351), .ZN(n1352) );
XNOR2_X1 U1079 ( .A(n1354), .B(n1355), .ZN(n1351) );
XOR2_X1 U1080 ( .A(n1288), .B(n1356), .Z(n1355) );
XOR2_X1 U1081 ( .A(G122), .B(G107), .Z(n1356) );
XOR2_X1 U1082 ( .A(G116), .B(KEYINPUT34), .Z(n1288) );
XNOR2_X1 U1083 ( .A(G128), .B(n1357), .ZN(n1354) );
XOR2_X1 U1084 ( .A(G143), .B(G134), .Z(n1357) );
INV_X1 U1085 ( .A(n1271), .ZN(n1090) );
XOR2_X1 U1086 ( .A(n1358), .B(G475), .Z(n1271) );
NAND2_X1 U1087 ( .A1(n1152), .A2(n1274), .ZN(n1358) );
INV_X1 U1088 ( .A(G902), .ZN(n1274) );
XOR2_X1 U1089 ( .A(n1359), .B(n1360), .Z(n1152) );
XOR2_X1 U1090 ( .A(n1361), .B(n1362), .Z(n1360) );
NAND2_X1 U1091 ( .A1(KEYINPUT38), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1092 ( .A(G104), .B(n1364), .Z(n1363) );
XOR2_X1 U1093 ( .A(G122), .B(G113), .Z(n1364) );
NAND2_X1 U1094 ( .A1(n1365), .A2(n1366), .ZN(n1361) );
OR2_X1 U1095 ( .A1(n1236), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1096 ( .A(n1368), .B(KEYINPUT37), .Z(n1365) );
NAND2_X1 U1097 ( .A1(n1236), .A2(n1367), .ZN(n1368) );
NAND3_X1 U1098 ( .A1(n1281), .A2(n1107), .A3(G214), .ZN(n1367) );
INV_X1 U1099 ( .A(G953), .ZN(n1107) );
INV_X1 U1100 ( .A(G237), .ZN(n1281) );
INV_X1 U1101 ( .A(G143), .ZN(n1236) );
XNOR2_X1 U1102 ( .A(G131), .B(n1369), .ZN(n1359) );
NOR2_X1 U1103 ( .A1(KEYINPUT18), .A2(n1370), .ZN(n1369) );
XOR2_X1 U1104 ( .A(n1371), .B(n1372), .Z(n1370) );
NOR2_X1 U1105 ( .A1(KEYINPUT17), .A2(n1308), .ZN(n1372) );
XOR2_X1 U1106 ( .A(G140), .B(KEYINPUT20), .Z(n1308) );
XOR2_X1 U1107 ( .A(G125), .B(n1232), .Z(n1371) );
INV_X1 U1108 ( .A(G146), .ZN(n1232) );
endmodule


