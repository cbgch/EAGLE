//Key = 1100111110010000100110010111101011000011100000110110100011000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296;

XNOR2_X1 U708 ( .A(G107), .B(n983), .ZN(G9) );
NOR2_X1 U709 ( .A1(n984), .A2(n985), .ZN(G75) );
NOR4_X1 U710 ( .A1(n986), .A2(n987), .A3(n988), .A4(n989), .ZN(n985) );
NOR2_X1 U711 ( .A1(n990), .A2(n991), .ZN(n988) );
NOR3_X1 U712 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n990) );
NOR3_X1 U713 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n994) );
NOR2_X1 U714 ( .A1(n998), .A2(n999), .ZN(n996) );
NOR2_X1 U715 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NOR2_X1 U716 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NOR3_X1 U717 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n998) );
INV_X1 U718 ( .A(n1007), .ZN(n995) );
NOR3_X1 U719 ( .A1(n1008), .A2(n1009), .A3(n1001), .ZN(n993) );
NOR2_X1 U720 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR2_X1 U721 ( .A1(KEYINPUT43), .A2(n1012), .ZN(n1010) );
NOR2_X1 U722 ( .A1(n1013), .A2(n1014), .ZN(n992) );
INV_X1 U723 ( .A(KEYINPUT43), .ZN(n1014) );
NOR3_X1 U724 ( .A1(n1008), .A2(n1012), .A3(n1001), .ZN(n1013) );
INV_X1 U725 ( .A(n1015), .ZN(n1008) );
XNOR2_X1 U726 ( .A(KEYINPUT20), .B(n1016), .ZN(n987) );
NAND3_X1 U727 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n986) );
NAND3_X1 U728 ( .A1(n1007), .A2(n1020), .A3(n1015), .ZN(n1019) );
NOR2_X1 U729 ( .A1(n1005), .A2(n997), .ZN(n1015) );
INV_X1 U730 ( .A(n1021), .ZN(n1005) );
NAND2_X1 U731 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NAND2_X1 U732 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U733 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U734 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U735 ( .A1(n1030), .A2(n1031), .ZN(n1022) );
AND3_X1 U736 ( .A1(n1017), .A2(n1018), .A3(n1032), .ZN(n984) );
NAND4_X1 U737 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1017) );
NOR4_X1 U738 ( .A1(n1037), .A2(n1028), .A3(n1038), .A4(n1039), .ZN(n1036) );
XOR2_X1 U739 ( .A(n1040), .B(n1041), .Z(n1038) );
NOR2_X1 U740 ( .A1(n1042), .A2(KEYINPUT12), .ZN(n1041) );
INV_X1 U741 ( .A(n1004), .ZN(n1037) );
NOR2_X1 U742 ( .A1(n1043), .A2(n1044), .ZN(n1035) );
XOR2_X1 U743 ( .A(n1045), .B(n1046), .Z(n1044) );
NOR2_X1 U744 ( .A1(KEYINPUT36), .A2(n1047), .ZN(n1046) );
XOR2_X1 U745 ( .A(n1048), .B(G475), .Z(n1034) );
XOR2_X1 U746 ( .A(n1049), .B(G469), .Z(n1033) );
XOR2_X1 U747 ( .A(n1050), .B(n1051), .Z(G72) );
NOR2_X1 U748 ( .A1(n1052), .A2(n1018), .ZN(n1051) );
NOR2_X1 U749 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U750 ( .A1(n1055), .A2(n1056), .ZN(n1050) );
NAND2_X1 U751 ( .A1(n1057), .A2(n1018), .ZN(n1056) );
XOR2_X1 U752 ( .A(n1058), .B(n1059), .Z(n1057) );
NAND2_X1 U753 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND3_X1 U754 ( .A1(G900), .A2(n1059), .A3(G953), .ZN(n1055) );
XOR2_X1 U755 ( .A(n1062), .B(n1063), .Z(n1059) );
XOR2_X1 U756 ( .A(n1064), .B(n1065), .Z(n1063) );
XOR2_X1 U757 ( .A(n1066), .B(n1067), .Z(n1062) );
XOR2_X1 U758 ( .A(n1068), .B(n1069), .Z(G69) );
XOR2_X1 U759 ( .A(n1070), .B(n1071), .Z(n1069) );
OR2_X1 U760 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U761 ( .A1(KEYINPUT39), .A2(n1074), .ZN(n1070) );
NAND2_X1 U762 ( .A1(n1075), .A2(n1016), .ZN(n1074) );
XOR2_X1 U763 ( .A(n1018), .B(KEYINPUT41), .Z(n1075) );
NAND2_X1 U764 ( .A1(G953), .A2(n1076), .ZN(n1068) );
NAND2_X1 U765 ( .A1(G898), .A2(G224), .ZN(n1076) );
NOR2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(G66) );
XOR2_X1 U767 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR2_X1 U769 ( .A1(n1077), .A2(n1083), .ZN(G63) );
XOR2_X1 U770 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U771 ( .A1(n1081), .A2(G478), .ZN(n1084) );
NOR2_X1 U772 ( .A1(n1077), .A2(n1086), .ZN(G60) );
XOR2_X1 U773 ( .A(n1087), .B(n1088), .Z(n1086) );
XOR2_X1 U774 ( .A(n1089), .B(KEYINPUT56), .Z(n1087) );
NAND2_X1 U775 ( .A1(n1081), .A2(G475), .ZN(n1089) );
XOR2_X1 U776 ( .A(n1090), .B(n1091), .Z(G6) );
NAND2_X1 U777 ( .A1(KEYINPUT30), .A2(G104), .ZN(n1091) );
NAND3_X1 U778 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1090) );
XOR2_X1 U779 ( .A(KEYINPUT60), .B(n1031), .Z(n1093) );
NOR2_X1 U780 ( .A1(n1077), .A2(n1095), .ZN(G57) );
XOR2_X1 U781 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U782 ( .A1(KEYINPUT55), .A2(n1098), .ZN(n1097) );
NAND2_X1 U783 ( .A1(n1099), .A2(n1100), .ZN(n1096) );
NAND2_X1 U784 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U785 ( .A(KEYINPUT6), .B(n1103), .Z(n1099) );
NOR2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1103) );
NAND2_X1 U787 ( .A1(n1081), .A2(G472), .ZN(n1102) );
XNOR2_X1 U788 ( .A(n1104), .B(n1105), .ZN(n1101) );
XOR2_X1 U789 ( .A(n1106), .B(KEYINPUT62), .Z(n1104) );
NOR3_X1 U790 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(G54) );
NOR3_X1 U791 ( .A1(n1110), .A2(n1018), .A3(n1032), .ZN(n1109) );
INV_X1 U792 ( .A(G952), .ZN(n1032) );
AND2_X1 U793 ( .A1(n1110), .A2(n1077), .ZN(n1108) );
INV_X1 U794 ( .A(KEYINPUT15), .ZN(n1110) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(n1107) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U797 ( .A1(n1081), .A2(G469), .ZN(n1113) );
XOR2_X1 U798 ( .A(n1115), .B(n1116), .Z(n1111) );
NOR3_X1 U799 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
AND2_X1 U800 ( .A1(n1120), .A2(KEYINPUT42), .ZN(n1119) );
NOR2_X1 U801 ( .A1(KEYINPUT42), .A2(n1121), .ZN(n1118) );
INV_X1 U802 ( .A(n1122), .ZN(n1121) );
NAND2_X1 U803 ( .A1(KEYINPUT16), .A2(n1123), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1077), .A2(n1124), .ZN(G51) );
XOR2_X1 U805 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U806 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U807 ( .A1(KEYINPUT26), .A2(n1072), .ZN(n1128) );
NAND2_X1 U808 ( .A1(n1081), .A2(G210), .ZN(n1127) );
AND2_X1 U809 ( .A1(G902), .A2(n1129), .ZN(n1081) );
OR2_X1 U810 ( .A1(n989), .A2(n1016), .ZN(n1129) );
NAND4_X1 U811 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1016) );
AND4_X1 U812 ( .A1(n983), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1133) );
NAND3_X1 U813 ( .A1(n1092), .A2(n1031), .A3(n1011), .ZN(n983) );
NAND2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NAND2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U816 ( .A(n1141), .B(KEYINPUT44), .Z(n1139) );
NAND3_X1 U817 ( .A1(n1092), .A2(n1031), .A3(n1094), .ZN(n1130) );
NAND2_X1 U818 ( .A1(n1142), .A2(n1060), .ZN(n989) );
AND4_X1 U819 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1060) );
NOR4_X1 U820 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
NOR3_X1 U821 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR2_X1 U822 ( .A1(KEYINPUT38), .A2(n1154), .ZN(n1153) );
NOR3_X1 U823 ( .A1(n991), .A2(n1031), .A3(n1155), .ZN(n1154) );
INV_X1 U824 ( .A(n1030), .ZN(n991) );
AND2_X1 U825 ( .A1(n1156), .A2(KEYINPUT38), .ZN(n1152) );
NOR3_X1 U826 ( .A1(n1137), .A2(KEYINPUT32), .A3(n1157), .ZN(n1148) );
NOR2_X1 U827 ( .A1(n1158), .A2(n1026), .ZN(n1147) );
NOR2_X1 U828 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U829 ( .A(KEYINPUT34), .B(n1161), .ZN(n1160) );
NOR2_X1 U830 ( .A1(n1157), .A2(n1162), .ZN(n1159) );
INV_X1 U831 ( .A(KEYINPUT32), .ZN(n1162) );
XOR2_X1 U832 ( .A(n1061), .B(KEYINPUT45), .Z(n1142) );
NOR2_X1 U833 ( .A1(n1018), .A2(G952), .ZN(n1077) );
XOR2_X1 U834 ( .A(G146), .B(n1163), .Z(G48) );
NOR2_X1 U835 ( .A1(n1164), .A2(n1026), .ZN(n1163) );
XOR2_X1 U836 ( .A(n1157), .B(KEYINPUT2), .Z(n1164) );
NAND4_X1 U837 ( .A1(n1094), .A2(n1031), .A3(n1165), .A4(n1043), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1155), .A2(n1166), .ZN(n1165) );
INV_X1 U839 ( .A(n1167), .ZN(n1155) );
XOR2_X1 U840 ( .A(G143), .B(n1149), .Z(G45) );
AND4_X1 U841 ( .A1(n1168), .A2(n1003), .A3(n1169), .A4(n1170), .ZN(n1149) );
XNOR2_X1 U842 ( .A(G140), .B(n1061), .ZN(G42) );
NAND3_X1 U843 ( .A1(n1094), .A2(n1171), .A3(n1002), .ZN(n1061) );
XOR2_X1 U844 ( .A(G137), .B(n1172), .Z(G39) );
NOR2_X1 U845 ( .A1(n1156), .A2(n1151), .ZN(n1172) );
XNOR2_X1 U846 ( .A(G134), .B(n1145), .ZN(G36) );
NAND3_X1 U847 ( .A1(n1011), .A2(n1003), .A3(n1171), .ZN(n1145) );
XOR2_X1 U848 ( .A(n1173), .B(n1143), .Z(G33) );
NAND3_X1 U849 ( .A1(n1171), .A2(n1003), .A3(n1094), .ZN(n1143) );
INV_X1 U850 ( .A(n1156), .ZN(n1171) );
NAND3_X1 U851 ( .A1(n1031), .A2(n1167), .A3(n1030), .ZN(n1156) );
NOR2_X1 U852 ( .A1(n1174), .A2(n1028), .ZN(n1030) );
XOR2_X1 U853 ( .A(n1175), .B(n1144), .Z(G30) );
NAND4_X1 U854 ( .A1(n1168), .A2(n1011), .A3(n1043), .A4(n1176), .ZN(n1144) );
AND3_X1 U855 ( .A1(n1137), .A2(n1167), .A3(n1031), .ZN(n1168) );
XOR2_X1 U856 ( .A(n1177), .B(n1131), .Z(G3) );
NAND3_X1 U857 ( .A1(n1137), .A2(n1003), .A3(n1178), .ZN(n1131) );
XOR2_X1 U858 ( .A(G125), .B(n1179), .Z(G27) );
NOR2_X1 U859 ( .A1(n1026), .A2(n1161), .ZN(n1179) );
NAND4_X1 U860 ( .A1(n1024), .A2(n1002), .A3(n1094), .A4(n1167), .ZN(n1161) );
NAND2_X1 U861 ( .A1(n997), .A2(n1180), .ZN(n1167) );
NAND4_X1 U862 ( .A1(G953), .A2(G902), .A3(n1181), .A4(n1054), .ZN(n1180) );
INV_X1 U863 ( .A(G900), .ZN(n1054) );
XOR2_X1 U864 ( .A(n1182), .B(G122), .Z(G24) );
NAND2_X1 U865 ( .A1(KEYINPUT23), .A2(n1136), .ZN(n1182) );
NAND4_X1 U866 ( .A1(n1024), .A2(n1092), .A3(n1169), .A4(n1170), .ZN(n1136) );
AND3_X1 U867 ( .A1(n1137), .A2(n1183), .A3(n1021), .ZN(n1092) );
XNOR2_X1 U868 ( .A(G119), .B(n1135), .ZN(G21) );
OR2_X1 U869 ( .A1(n1184), .A2(n1151), .ZN(n1135) );
NAND3_X1 U870 ( .A1(n1043), .A2(n1176), .A3(n1007), .ZN(n1151) );
NAND2_X1 U871 ( .A1(n1185), .A2(n1186), .ZN(G18) );
NAND2_X1 U872 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U873 ( .A(n1189), .B(n1190), .Z(n1185) );
NOR2_X1 U874 ( .A1(n1026), .A2(n1141), .ZN(n1190) );
NAND4_X1 U875 ( .A1(n1024), .A2(n1011), .A3(n1003), .A4(n1183), .ZN(n1141) );
NOR2_X1 U876 ( .A1(n1170), .A2(n1191), .ZN(n1011) );
INV_X1 U877 ( .A(n1137), .ZN(n1026) );
OR2_X1 U878 ( .A1(n1188), .A2(n1187), .ZN(n1189) );
XOR2_X1 U879 ( .A(G116), .B(KEYINPUT11), .Z(n1187) );
INV_X1 U880 ( .A(KEYINPUT0), .ZN(n1188) );
XOR2_X1 U881 ( .A(n1134), .B(n1192), .Z(G15) );
XOR2_X1 U882 ( .A(KEYINPUT50), .B(G113), .Z(n1192) );
NAND3_X1 U883 ( .A1(n1094), .A2(n1003), .A3(n1193), .ZN(n1134) );
INV_X1 U884 ( .A(n1184), .ZN(n1193) );
NAND3_X1 U885 ( .A1(n1137), .A2(n1183), .A3(n1024), .ZN(n1184) );
INV_X1 U886 ( .A(n1001), .ZN(n1024) );
NAND2_X1 U887 ( .A1(n1194), .A2(n1004), .ZN(n1001) );
XNOR2_X1 U888 ( .A(n1006), .B(KEYINPUT21), .ZN(n1194) );
XNOR2_X1 U889 ( .A(n1195), .B(KEYINPUT49), .ZN(n1006) );
NAND2_X1 U890 ( .A1(n1196), .A2(n1197), .ZN(n1003) );
OR3_X1 U891 ( .A1(n1166), .A2(n1043), .A3(KEYINPUT29), .ZN(n1197) );
NAND2_X1 U892 ( .A1(KEYINPUT29), .A2(n1021), .ZN(n1196) );
NOR2_X1 U893 ( .A1(n1176), .A2(n1043), .ZN(n1021) );
INV_X1 U894 ( .A(n1166), .ZN(n1176) );
INV_X1 U895 ( .A(n1012), .ZN(n1094) );
NAND2_X1 U896 ( .A1(n1191), .A2(n1170), .ZN(n1012) );
XOR2_X1 U897 ( .A(n1198), .B(n1199), .Z(G12) );
NAND2_X1 U898 ( .A1(n1137), .A2(n1200), .ZN(n1199) );
XNOR2_X1 U899 ( .A(KEYINPUT13), .B(n1140), .ZN(n1200) );
NAND2_X1 U900 ( .A1(n1178), .A2(n1002), .ZN(n1140) );
AND2_X1 U901 ( .A1(n1166), .A2(n1043), .ZN(n1002) );
XNOR2_X1 U902 ( .A(n1201), .B(n1082), .ZN(n1043) );
AND2_X1 U903 ( .A1(G217), .A2(n1202), .ZN(n1082) );
NAND2_X1 U904 ( .A1(n1080), .A2(n1203), .ZN(n1201) );
XOR2_X1 U905 ( .A(n1204), .B(n1205), .Z(n1080) );
XOR2_X1 U906 ( .A(G110), .B(n1206), .Z(n1205) );
XOR2_X1 U907 ( .A(G137), .B(G119), .Z(n1206) );
XOR2_X1 U908 ( .A(n1207), .B(n1208), .Z(n1204) );
XOR2_X1 U909 ( .A(n1209), .B(n1210), .Z(n1207) );
NAND2_X1 U910 ( .A1(G221), .A2(n1211), .ZN(n1209) );
XOR2_X1 U911 ( .A(n1212), .B(n1039), .Z(n1166) );
XNOR2_X1 U912 ( .A(n1213), .B(G472), .ZN(n1039) );
NAND2_X1 U913 ( .A1(n1214), .A2(n1203), .ZN(n1213) );
XNOR2_X1 U914 ( .A(n1215), .B(n1098), .ZN(n1214) );
XNOR2_X1 U915 ( .A(n1216), .B(n1177), .ZN(n1098) );
INV_X1 U916 ( .A(G101), .ZN(n1177) );
NAND2_X1 U917 ( .A1(G210), .A2(n1217), .ZN(n1216) );
XOR2_X1 U918 ( .A(n1218), .B(n1219), .Z(n1215) );
INV_X1 U919 ( .A(n1106), .ZN(n1219) );
NAND2_X1 U920 ( .A1(KEYINPUT4), .A2(n1105), .ZN(n1218) );
XNOR2_X1 U921 ( .A(n1220), .B(n1221), .ZN(n1105) );
XNOR2_X1 U922 ( .A(KEYINPUT63), .B(KEYINPUT27), .ZN(n1212) );
AND3_X1 U923 ( .A1(n1031), .A2(n1183), .A3(n1007), .ZN(n1178) );
NOR2_X1 U924 ( .A1(n1169), .A2(n1170), .ZN(n1007) );
NAND2_X1 U925 ( .A1(n1222), .A2(n1223), .ZN(n1170) );
NAND2_X1 U926 ( .A1(n1224), .A2(KEYINPUT3), .ZN(n1223) );
XOR2_X1 U927 ( .A(n1048), .B(n1225), .Z(n1222) );
NOR2_X1 U928 ( .A1(KEYINPUT3), .A2(n1224), .ZN(n1225) );
XNOR2_X1 U929 ( .A(KEYINPUT24), .B(G475), .ZN(n1224) );
OR2_X1 U930 ( .A1(n1088), .A2(G902), .ZN(n1048) );
XNOR2_X1 U931 ( .A(n1226), .B(G122), .ZN(n1088) );
XOR2_X1 U932 ( .A(n1227), .B(n1228), .Z(n1226) );
XOR2_X1 U933 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U934 ( .A(G131), .B(G104), .Z(n1230) );
XOR2_X1 U935 ( .A(KEYINPUT9), .B(G146), .Z(n1229) );
XOR2_X1 U936 ( .A(n1231), .B(n1232), .Z(n1227) );
XOR2_X1 U937 ( .A(n1233), .B(n1234), .Z(n1232) );
NOR2_X1 U938 ( .A1(KEYINPUT17), .A2(n1235), .ZN(n1234) );
AND2_X1 U939 ( .A1(n1217), .A2(G214), .ZN(n1233) );
NOR2_X1 U940 ( .A1(G953), .A2(G237), .ZN(n1217) );
XOR2_X1 U941 ( .A(n1236), .B(n1208), .Z(n1231) );
XOR2_X1 U942 ( .A(n1065), .B(KEYINPUT8), .Z(n1208) );
XOR2_X1 U943 ( .A(G125), .B(G140), .Z(n1065) );
INV_X1 U944 ( .A(n1191), .ZN(n1169) );
XOR2_X1 U945 ( .A(n1047), .B(n1045), .Z(n1191) );
AND2_X1 U946 ( .A1(n1237), .A2(n1085), .ZN(n1045) );
XOR2_X1 U947 ( .A(n1238), .B(n1239), .Z(n1085) );
NOR2_X1 U948 ( .A1(KEYINPUT48), .A2(n1240), .ZN(n1239) );
XOR2_X1 U949 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U950 ( .A(G107), .B(n1243), .Z(n1242) );
XOR2_X1 U951 ( .A(G128), .B(G116), .Z(n1243) );
XOR2_X1 U952 ( .A(n1244), .B(n1245), .Z(n1241) );
XOR2_X1 U953 ( .A(n1246), .B(n1247), .Z(n1244) );
NOR2_X1 U954 ( .A1(KEYINPUT35), .A2(n1236), .ZN(n1247) );
NAND2_X1 U955 ( .A1(n1248), .A2(n1249), .ZN(n1246) );
XNOR2_X1 U956 ( .A(KEYINPUT61), .B(KEYINPUT28), .ZN(n1249) );
XOR2_X1 U957 ( .A(n1250), .B(KEYINPUT14), .Z(n1248) );
INV_X1 U958 ( .A(G122), .ZN(n1250) );
NAND2_X1 U959 ( .A1(n1251), .A2(n1211), .ZN(n1238) );
AND2_X1 U960 ( .A1(G234), .A2(n1018), .ZN(n1211) );
XNOR2_X1 U961 ( .A(G217), .B(KEYINPUT19), .ZN(n1251) );
XOR2_X1 U962 ( .A(n1203), .B(KEYINPUT31), .Z(n1237) );
INV_X1 U963 ( .A(G478), .ZN(n1047) );
NAND2_X1 U964 ( .A1(n1252), .A2(n1253), .ZN(n1183) );
NAND3_X1 U965 ( .A1(G902), .A2(n1181), .A3(n1073), .ZN(n1253) );
NOR2_X1 U966 ( .A1(n1018), .A2(G898), .ZN(n1073) );
XOR2_X1 U967 ( .A(n997), .B(KEYINPUT18), .Z(n1252) );
NAND3_X1 U968 ( .A1(n1181), .A2(n1018), .A3(G952), .ZN(n997) );
NAND2_X1 U969 ( .A1(G237), .A2(G234), .ZN(n1181) );
AND2_X1 U970 ( .A1(n1195), .A2(n1004), .ZN(n1031) );
NAND2_X1 U971 ( .A1(G221), .A2(n1202), .ZN(n1004) );
NAND2_X1 U972 ( .A1(n1254), .A2(n1203), .ZN(n1202) );
XOR2_X1 U973 ( .A(KEYINPUT58), .B(G234), .Z(n1254) );
XNOR2_X1 U974 ( .A(n1255), .B(n1049), .ZN(n1195) );
NAND2_X1 U975 ( .A1(n1256), .A2(n1203), .ZN(n1049) );
XOR2_X1 U976 ( .A(n1257), .B(n1258), .Z(n1256) );
NOR2_X1 U977 ( .A1(n1122), .A2(n1117), .ZN(n1258) );
AND2_X1 U978 ( .A1(n1120), .A2(n1259), .ZN(n1117) );
NAND2_X1 U979 ( .A1(G227), .A2(n1018), .ZN(n1259) );
NOR3_X1 U980 ( .A1(n1120), .A2(G953), .A3(n1053), .ZN(n1122) );
INV_X1 U981 ( .A(G227), .ZN(n1053) );
XOR2_X1 U982 ( .A(G140), .B(G110), .Z(n1120) );
NAND2_X1 U983 ( .A1(n1260), .A2(n1261), .ZN(n1257) );
NAND2_X1 U984 ( .A1(n1114), .A2(n1123), .ZN(n1261) );
XOR2_X1 U985 ( .A(n1262), .B(KEYINPUT51), .Z(n1260) );
OR2_X1 U986 ( .A1(n1123), .A2(n1114), .ZN(n1262) );
XNOR2_X1 U987 ( .A(n1220), .B(KEYINPUT7), .ZN(n1114) );
XNOR2_X1 U988 ( .A(n1064), .B(n1263), .ZN(n1220) );
NOR2_X1 U989 ( .A1(KEYINPUT10), .A2(n1264), .ZN(n1263) );
XOR2_X1 U990 ( .A(n1066), .B(KEYINPUT54), .Z(n1264) );
INV_X1 U991 ( .A(G137), .ZN(n1066) );
XNOR2_X1 U992 ( .A(n1173), .B(n1245), .ZN(n1064) );
XOR2_X1 U993 ( .A(G134), .B(KEYINPUT22), .Z(n1245) );
INV_X1 U994 ( .A(G131), .ZN(n1173) );
XNOR2_X1 U995 ( .A(n1265), .B(n1067), .ZN(n1123) );
XNOR2_X1 U996 ( .A(n1221), .B(KEYINPUT37), .ZN(n1067) );
XOR2_X1 U997 ( .A(n1266), .B(G101), .Z(n1265) );
NAND2_X1 U998 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U999 ( .A1(G107), .A2(n1269), .ZN(n1268) );
XOR2_X1 U1000 ( .A(KEYINPUT33), .B(n1270), .Z(n1267) );
NOR2_X1 U1001 ( .A1(G107), .A2(n1269), .ZN(n1270) );
INV_X1 U1002 ( .A(G104), .ZN(n1269) );
NAND2_X1 U1003 ( .A1(KEYINPUT46), .A2(n1271), .ZN(n1255) );
INV_X1 U1004 ( .A(G469), .ZN(n1271) );
NOR2_X1 U1005 ( .A1(n1029), .A2(n1028), .ZN(n1137) );
AND2_X1 U1006 ( .A1(G214), .A2(n1272), .ZN(n1028) );
INV_X1 U1007 ( .A(n1174), .ZN(n1029) );
NAND3_X1 U1008 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1174) );
OR2_X1 U1009 ( .A1(n1042), .A2(KEYINPUT1), .ZN(n1275) );
NAND3_X1 U1010 ( .A1(KEYINPUT1), .A2(n1042), .A3(n1040), .ZN(n1274) );
NAND2_X1 U1011 ( .A1(n1276), .A2(n1277), .ZN(n1273) );
NAND2_X1 U1012 ( .A1(KEYINPUT1), .A2(n1278), .ZN(n1277) );
XOR2_X1 U1013 ( .A(KEYINPUT59), .B(n1042), .Z(n1278) );
AND2_X1 U1014 ( .A1(n1279), .A2(n1272), .ZN(n1042) );
OR2_X1 U1015 ( .A1(G902), .A2(G237), .ZN(n1272) );
XNOR2_X1 U1016 ( .A(G210), .B(KEYINPUT40), .ZN(n1279) );
INV_X1 U1017 ( .A(n1040), .ZN(n1276) );
NAND2_X1 U1018 ( .A1(n1280), .A2(n1203), .ZN(n1040) );
INV_X1 U1019 ( .A(G902), .ZN(n1203) );
XOR2_X1 U1020 ( .A(n1281), .B(n1125), .Z(n1280) );
XNOR2_X1 U1021 ( .A(n1282), .B(n1221), .ZN(n1125) );
XOR2_X1 U1022 ( .A(n1210), .B(n1236), .Z(n1221) );
XNOR2_X1 U1023 ( .A(G143), .B(KEYINPUT53), .ZN(n1236) );
XNOR2_X1 U1024 ( .A(n1175), .B(G146), .ZN(n1210) );
INV_X1 U1025 ( .A(G128), .ZN(n1175) );
XNOR2_X1 U1026 ( .A(G125), .B(n1283), .ZN(n1282) );
AND2_X1 U1027 ( .A1(n1018), .A2(G224), .ZN(n1283) );
INV_X1 U1028 ( .A(G953), .ZN(n1018) );
NAND2_X1 U1029 ( .A1(KEYINPUT25), .A2(n1072), .ZN(n1281) );
XOR2_X1 U1030 ( .A(n1284), .B(n1285), .Z(n1072) );
XOR2_X1 U1031 ( .A(n1286), .B(n1106), .Z(n1285) );
XOR2_X1 U1032 ( .A(n1235), .B(n1287), .Z(n1106) );
XOR2_X1 U1033 ( .A(G119), .B(G116), .Z(n1287) );
INV_X1 U1034 ( .A(G113), .ZN(n1235) );
NAND2_X1 U1035 ( .A1(KEYINPUT52), .A2(n1288), .ZN(n1286) );
NAND2_X1 U1036 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U1037 ( .A1(G104), .A2(n1291), .ZN(n1290) );
XOR2_X1 U1038 ( .A(KEYINPUT57), .B(n1292), .Z(n1289) );
NOR2_X1 U1039 ( .A1(G104), .A2(n1291), .ZN(n1292) );
XOR2_X1 U1040 ( .A(KEYINPUT47), .B(G107), .Z(n1291) );
XOR2_X1 U1041 ( .A(n1293), .B(G101), .Z(n1284) );
NAND2_X1 U1042 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NAND2_X1 U1043 ( .A1(G122), .A2(n1198), .ZN(n1295) );
XOR2_X1 U1044 ( .A(KEYINPUT5), .B(n1296), .Z(n1294) );
NOR2_X1 U1045 ( .A1(G122), .A2(n1198), .ZN(n1296) );
INV_X1 U1046 ( .A(G110), .ZN(n1198) );
endmodule


