//Key = 0111110101110110111011111101010011001000100111011000110111000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311;

XOR2_X1 U718 ( .A(n984), .B(n985), .Z(G9) );
NOR2_X1 U719 ( .A1(n986), .A2(n987), .ZN(G75) );
XOR2_X1 U720 ( .A(KEYINPUT30), .B(n988), .Z(n987) );
NOR3_X1 U721 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n988) );
NOR3_X1 U722 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n990) );
NOR2_X1 U723 ( .A1(n995), .A2(n996), .ZN(n993) );
NOR2_X1 U724 ( .A1(n997), .A2(n998), .ZN(n996) );
NOR2_X1 U725 ( .A1(n999), .A2(n1000), .ZN(n997) );
NOR2_X1 U726 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NOR2_X1 U727 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U728 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U729 ( .A1(n1007), .A2(n1008), .ZN(n999) );
NOR2_X1 U730 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR2_X1 U731 ( .A1(KEYINPUT31), .A2(n1011), .ZN(n1009) );
NOR3_X1 U732 ( .A1(n1008), .A2(n1012), .A3(n1002), .ZN(n995) );
INV_X1 U733 ( .A(n1013), .ZN(n1002) );
NOR2_X1 U734 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
INV_X1 U736 ( .A(n1018), .ZN(n1008) );
NAND3_X1 U737 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n989) );
NAND4_X1 U738 ( .A1(n1018), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1021) );
NAND2_X1 U739 ( .A1(n1025), .A2(n992), .ZN(n1024) );
NAND3_X1 U740 ( .A1(n1026), .A2(n1027), .A3(KEYINPUT31), .ZN(n1025) );
NAND2_X1 U741 ( .A1(n1028), .A2(n1029), .ZN(n1023) );
NAND2_X1 U742 ( .A1(n1013), .A2(n1030), .ZN(n1029) );
NAND2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
INV_X1 U745 ( .A(n992), .ZN(n1028) );
NOR3_X1 U746 ( .A1(n1035), .A2(G953), .A3(G952), .ZN(n986) );
INV_X1 U747 ( .A(n1019), .ZN(n1035) );
NAND4_X1 U748 ( .A1(n1034), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1019) );
NOR3_X1 U749 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
XOR2_X1 U750 ( .A(n1042), .B(n1043), .Z(n1041) );
NAND2_X1 U751 ( .A1(KEYINPUT10), .A2(n1044), .ZN(n1042) );
XOR2_X1 U752 ( .A(KEYINPUT13), .B(n1045), .Z(n1044) );
NAND3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1017), .ZN(n1039) );
NOR3_X1 U754 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1037) );
NOR3_X1 U755 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NOR2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
INV_X1 U759 ( .A(KEYINPUT57), .ZN(n1059) );
NOR2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1058) );
INV_X1 U761 ( .A(KEYINPUT62), .ZN(n1053) );
NOR2_X1 U762 ( .A1(KEYINPUT57), .A2(n1052), .ZN(n1056) );
XOR2_X1 U763 ( .A(G469), .B(n1060), .Z(n1048) );
XOR2_X1 U764 ( .A(KEYINPUT42), .B(n1061), .Z(n1036) );
NOR2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
AND2_X1 U766 ( .A1(n1064), .A2(G475), .ZN(n1062) );
XOR2_X1 U767 ( .A(n1065), .B(n1066), .Z(G72) );
XOR2_X1 U768 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U769 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U770 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND3_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1071) );
NAND2_X1 U772 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
OR3_X1 U773 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1074) );
INV_X1 U774 ( .A(KEYINPUT32), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1078), .ZN(n1073) );
NAND2_X1 U776 ( .A1(KEYINPUT9), .A2(n1080), .ZN(n1078) );
NOR2_X1 U777 ( .A1(G900), .A2(n1020), .ZN(n1069) );
NAND2_X1 U778 ( .A1(G953), .A2(n1081), .ZN(n1067) );
NAND2_X1 U779 ( .A1(G900), .A2(G227), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1020), .A2(n1082), .ZN(n1065) );
NAND2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(G69) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
OR2_X1 U783 ( .A1(n1020), .A2(G224), .ZN(n1086) );
INV_X1 U784 ( .A(n1087), .ZN(n1085) );
NAND3_X1 U785 ( .A1(G953), .A2(n1088), .A3(n1087), .ZN(n1083) );
XOR2_X1 U786 ( .A(n1089), .B(n1090), .Z(n1087) );
NOR2_X1 U787 ( .A1(n1091), .A2(G953), .ZN(n1090) );
NOR2_X1 U788 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U789 ( .A1(n1094), .A2(n1095), .ZN(n1089) );
NAND2_X1 U790 ( .A1(G953), .A2(n1096), .ZN(n1095) );
XOR2_X1 U791 ( .A(n1097), .B(n1098), .Z(n1094) );
NAND2_X1 U792 ( .A1(KEYINPUT45), .A2(n1099), .ZN(n1097) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1088) );
NOR2_X1 U794 ( .A1(n1100), .A2(n1101), .ZN(G66) );
NOR3_X1 U795 ( .A1(n1045), .A2(n1102), .A3(n1103), .ZN(n1101) );
AND3_X1 U796 ( .A1(n1104), .A2(G217), .A3(n1105), .ZN(n1103) );
NOR2_X1 U797 ( .A1(n1106), .A2(n1104), .ZN(n1102) );
AND2_X1 U798 ( .A1(n991), .A2(G217), .ZN(n1106) );
NOR2_X1 U799 ( .A1(n1100), .A2(n1107), .ZN(G63) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U801 ( .A1(n1105), .A2(G478), .ZN(n1108) );
NOR2_X1 U802 ( .A1(n1100), .A2(n1110), .ZN(G60) );
NOR2_X1 U803 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U804 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U805 ( .A1(n1105), .A2(G475), .ZN(n1114) );
NAND2_X1 U806 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR2_X1 U807 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
INV_X1 U808 ( .A(KEYINPUT34), .ZN(n1116) );
XNOR2_X1 U809 ( .A(G104), .B(n1117), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1118), .A2(KEYINPUT51), .ZN(n1117) );
NOR3_X1 U811 ( .A1(n1011), .A2(n994), .A3(n1119), .ZN(n1118) );
NOR2_X1 U812 ( .A1(n1100), .A2(n1120), .ZN(G57) );
XOR2_X1 U813 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U814 ( .A1(KEYINPUT12), .A2(n1123), .ZN(n1121) );
XOR2_X1 U815 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U816 ( .A(n1080), .B(n1126), .Z(n1125) );
XOR2_X1 U817 ( .A(n1127), .B(n1128), .Z(n1124) );
NOR3_X1 U818 ( .A1(n1129), .A2(KEYINPUT8), .A3(n1130), .ZN(n1128) );
INV_X1 U819 ( .A(G472), .ZN(n1130) );
XOR2_X1 U820 ( .A(n1131), .B(KEYINPUT17), .Z(n1127) );
NOR2_X1 U821 ( .A1(n1100), .A2(n1132), .ZN(G54) );
XOR2_X1 U822 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U823 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR2_X1 U824 ( .A1(n1137), .A2(KEYINPUT58), .ZN(n1136) );
AND2_X1 U825 ( .A1(G469), .A2(n1105), .ZN(n1137) );
INV_X1 U826 ( .A(n1129), .ZN(n1105) );
NAND2_X1 U827 ( .A1(KEYINPUT29), .A2(n1138), .ZN(n1135) );
XOR2_X1 U828 ( .A(KEYINPUT25), .B(G110), .Z(n1138) );
XOR2_X1 U829 ( .A(n1139), .B(n1140), .Z(n1133) );
XOR2_X1 U830 ( .A(G140), .B(n1141), .Z(n1140) );
NOR2_X1 U831 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XOR2_X1 U832 ( .A(n1144), .B(KEYINPUT55), .Z(n1143) );
NAND2_X1 U833 ( .A1(n1080), .A2(n1145), .ZN(n1144) );
NOR2_X1 U834 ( .A1(n1080), .A2(n1145), .ZN(n1142) );
NAND2_X1 U835 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U836 ( .A1(n1148), .A2(n1079), .ZN(n1147) );
XOR2_X1 U837 ( .A(KEYINPUT21), .B(n1149), .Z(n1146) );
NOR2_X1 U838 ( .A1(n1079), .A2(n1148), .ZN(n1149) );
XNOR2_X1 U839 ( .A(KEYINPUT26), .B(n1150), .ZN(n1148) );
NOR2_X1 U840 ( .A1(n1100), .A2(n1151), .ZN(G51) );
NOR2_X1 U841 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U842 ( .A(KEYINPUT50), .B(n1154), .Z(n1153) );
AND2_X1 U843 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U844 ( .A1(n1156), .A2(n1155), .ZN(n1152) );
XNOR2_X1 U845 ( .A(n1157), .B(n1158), .ZN(n1155) );
NAND3_X1 U846 ( .A1(n1159), .A2(n1160), .A3(KEYINPUT40), .ZN(n1157) );
NAND2_X1 U847 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U848 ( .A(KEYINPUT20), .B(n1163), .Z(n1159) );
NOR2_X1 U849 ( .A1(n1162), .A2(n1161), .ZN(n1163) );
XOR2_X1 U850 ( .A(n1164), .B(KEYINPUT19), .Z(n1161) );
NOR2_X1 U851 ( .A1(n1129), .A2(n1051), .ZN(n1156) );
NAND2_X1 U852 ( .A1(G902), .A2(n991), .ZN(n1129) );
OR3_X1 U853 ( .A1(n1093), .A2(n1165), .A3(n1082), .ZN(n991) );
NAND2_X1 U854 ( .A1(n1166), .A2(n1167), .ZN(n1082) );
NOR4_X1 U855 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
AND4_X1 U856 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1166) );
XOR2_X1 U857 ( .A(KEYINPUT15), .B(n1092), .Z(n1165) );
NAND4_X1 U858 ( .A1(n1176), .A2(n1177), .A3(n985), .A4(n1178), .ZN(n1092) );
NAND3_X1 U859 ( .A1(n1027), .A2(n1010), .A3(n1179), .ZN(n985) );
NAND4_X1 U860 ( .A1(n1026), .A2(n1015), .A3(n1180), .A4(n1181), .ZN(n1176) );
XOR2_X1 U861 ( .A(KEYINPUT46), .B(n1004), .Z(n1181) );
NOR2_X1 U862 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
XOR2_X1 U863 ( .A(n994), .B(KEYINPUT59), .Z(n1183) );
INV_X1 U864 ( .A(n1184), .ZN(n1182) );
NAND4_X1 U865 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1093) );
NOR2_X1 U866 ( .A1(n1020), .A2(G952), .ZN(n1100) );
NAND2_X1 U867 ( .A1(n1189), .A2(n1190), .ZN(G48) );
NAND2_X1 U868 ( .A1(G146), .A2(n1175), .ZN(n1190) );
XOR2_X1 U869 ( .A(KEYINPUT2), .B(n1191), .Z(n1189) );
NOR2_X1 U870 ( .A1(G146), .A2(n1175), .ZN(n1191) );
NAND3_X1 U871 ( .A1(n1026), .A2(n1004), .A3(n1192), .ZN(n1175) );
XOR2_X1 U872 ( .A(n1193), .B(n1174), .Z(G45) );
NAND4_X1 U873 ( .A1(n1015), .A2(n1004), .A3(n1194), .A4(n1195), .ZN(n1174) );
AND3_X1 U874 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1195) );
XOR2_X1 U875 ( .A(n1199), .B(G140), .Z(G42) );
NAND2_X1 U876 ( .A1(KEYINPUT63), .A2(n1173), .ZN(n1199) );
NAND3_X1 U877 ( .A1(n1200), .A2(n1015), .A3(n1018), .ZN(n1173) );
XNOR2_X1 U878 ( .A(n1172), .B(n1201), .ZN(G39) );
XOR2_X1 U879 ( .A(KEYINPUT54), .B(G137), .Z(n1201) );
NAND3_X1 U880 ( .A1(n1192), .A2(n1013), .A3(n1018), .ZN(n1172) );
XOR2_X1 U881 ( .A(G134), .B(n1171), .Z(G36) );
AND2_X1 U882 ( .A1(n1202), .A2(n1010), .ZN(n1171) );
XOR2_X1 U883 ( .A(G131), .B(n1170), .Z(G33) );
AND2_X1 U884 ( .A1(n1202), .A2(n1026), .ZN(n1170) );
AND4_X1 U885 ( .A1(n1018), .A2(n1194), .A3(n1015), .A4(n1196), .ZN(n1202) );
NOR2_X1 U886 ( .A1(n1005), .A2(n1040), .ZN(n1018) );
INV_X1 U887 ( .A(n1006), .ZN(n1040) );
XOR2_X1 U888 ( .A(G128), .B(n1169), .Z(G30) );
AND3_X1 U889 ( .A1(n1004), .A2(n1010), .A3(n1192), .ZN(n1169) );
AND4_X1 U890 ( .A1(n1203), .A2(n1033), .A3(n1015), .A4(n1196), .ZN(n1192) );
XNOR2_X1 U891 ( .A(G101), .B(n1178), .ZN(G3) );
NAND3_X1 U892 ( .A1(n1179), .A2(n1013), .A3(n1194), .ZN(n1178) );
XOR2_X1 U893 ( .A(n1204), .B(n1168), .Z(G27) );
AND3_X1 U894 ( .A1(n1200), .A2(n1004), .A3(n1022), .ZN(n1168) );
AND4_X1 U895 ( .A1(n1033), .A2(n1026), .A3(n1034), .A4(n1196), .ZN(n1200) );
NAND2_X1 U896 ( .A1(n992), .A2(n1205), .ZN(n1196) );
NAND4_X1 U897 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1207), .ZN(n1205) );
INV_X1 U898 ( .A(G900), .ZN(n1207) );
NAND2_X1 U899 ( .A1(KEYINPUT4), .A2(n1208), .ZN(n1204) );
XNOR2_X1 U900 ( .A(G122), .B(n1186), .ZN(G24) );
NAND4_X1 U901 ( .A1(n1209), .A2(n1027), .A3(n1198), .A4(n1197), .ZN(n1186) );
INV_X1 U902 ( .A(n994), .ZN(n1027) );
NAND2_X1 U903 ( .A1(n1034), .A2(n1210), .ZN(n994) );
XNOR2_X1 U904 ( .A(G119), .B(n1211), .ZN(G21) );
NAND2_X1 U905 ( .A1(KEYINPUT1), .A2(n1212), .ZN(n1211) );
INV_X1 U906 ( .A(n1185), .ZN(n1212) );
NAND4_X1 U907 ( .A1(n1203), .A2(n1209), .A3(n1033), .A4(n1013), .ZN(n1185) );
XNOR2_X1 U908 ( .A(G116), .B(n1187), .ZN(G18) );
NAND3_X1 U909 ( .A1(n1194), .A2(n1010), .A3(n1209), .ZN(n1187) );
NAND2_X1 U910 ( .A1(n1213), .A2(n1214), .ZN(n1010) );
OR3_X1 U911 ( .A1(n1198), .A2(n1215), .A3(KEYINPUT61), .ZN(n1214) );
NAND2_X1 U912 ( .A1(KEYINPUT61), .A2(n1013), .ZN(n1213) );
XOR2_X1 U913 ( .A(n1216), .B(n1188), .Z(G15) );
NAND3_X1 U914 ( .A1(n1194), .A2(n1026), .A3(n1209), .ZN(n1188) );
AND3_X1 U915 ( .A1(n1004), .A2(n1184), .A3(n1022), .ZN(n1209) );
INV_X1 U916 ( .A(n998), .ZN(n1022) );
NAND2_X1 U917 ( .A1(n1017), .A2(n1217), .ZN(n998) );
INV_X1 U918 ( .A(n1011), .ZN(n1026) );
NAND2_X1 U919 ( .A1(n1215), .A2(n1198), .ZN(n1011) );
INV_X1 U920 ( .A(n1197), .ZN(n1215) );
INV_X1 U921 ( .A(n1031), .ZN(n1194) );
NAND2_X1 U922 ( .A1(n1203), .A2(n1210), .ZN(n1031) );
XOR2_X1 U923 ( .A(n1034), .B(KEYINPUT7), .Z(n1203) );
XNOR2_X1 U924 ( .A(G110), .B(n1177), .ZN(G12) );
NAND4_X1 U925 ( .A1(n1033), .A2(n1179), .A3(n1034), .A4(n1013), .ZN(n1177) );
NOR2_X1 U926 ( .A1(n1197), .A2(n1198), .ZN(n1013) );
NAND2_X1 U927 ( .A1(n1218), .A2(n1219), .ZN(n1198) );
NAND2_X1 U928 ( .A1(G475), .A2(n1064), .ZN(n1219) );
XOR2_X1 U929 ( .A(KEYINPUT56), .B(n1063), .Z(n1218) );
NOR2_X1 U930 ( .A1(n1064), .A2(G475), .ZN(n1063) );
NAND2_X1 U931 ( .A1(n1115), .A2(n1220), .ZN(n1064) );
XOR2_X1 U932 ( .A(n1221), .B(n1222), .Z(n1115) );
XOR2_X1 U933 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U934 ( .A(G113), .B(G104), .Z(n1224) );
XOR2_X1 U935 ( .A(G143), .B(G122), .Z(n1223) );
XNOR2_X1 U936 ( .A(n1225), .B(n1226), .ZN(n1221) );
XOR2_X1 U937 ( .A(n1227), .B(n1228), .Z(n1226) );
NAND2_X1 U938 ( .A1(n1229), .A2(G214), .ZN(n1228) );
NAND2_X1 U939 ( .A1(n1230), .A2(n1231), .ZN(n1227) );
XNOR2_X1 U940 ( .A(KEYINPUT49), .B(KEYINPUT35), .ZN(n1230) );
NAND2_X1 U941 ( .A1(n1232), .A2(n1046), .ZN(n1197) );
NAND3_X1 U942 ( .A1(n1233), .A2(n1220), .A3(n1109), .ZN(n1046) );
INV_X1 U943 ( .A(G478), .ZN(n1233) );
XNOR2_X1 U944 ( .A(KEYINPUT53), .B(n1047), .ZN(n1232) );
NAND2_X1 U945 ( .A1(G478), .A2(n1234), .ZN(n1047) );
NAND2_X1 U946 ( .A1(n1109), .A2(n1220), .ZN(n1234) );
XOR2_X1 U947 ( .A(n1235), .B(n1236), .Z(n1109) );
XOR2_X1 U948 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U949 ( .A(n984), .B(G122), .Z(n1238) );
NAND2_X1 U950 ( .A1(G217), .A2(n1239), .ZN(n1237) );
XOR2_X1 U951 ( .A(n1240), .B(n1241), .Z(n1235) );
XOR2_X1 U952 ( .A(n1242), .B(n1243), .Z(n1240) );
NAND2_X1 U953 ( .A1(KEYINPUT24), .A2(G134), .ZN(n1242) );
XOR2_X1 U954 ( .A(n1244), .B(G472), .Z(n1034) );
NAND2_X1 U955 ( .A1(n1245), .A2(n1220), .ZN(n1244) );
XNOR2_X1 U956 ( .A(n1246), .B(n1122), .ZN(n1245) );
XNOR2_X1 U957 ( .A(n1247), .B(G101), .ZN(n1122) );
NAND2_X1 U958 ( .A1(n1229), .A2(G210), .ZN(n1247) );
NOR2_X1 U959 ( .A1(G953), .A2(G237), .ZN(n1229) );
NAND2_X1 U960 ( .A1(KEYINPUT36), .A2(n1248), .ZN(n1246) );
XOR2_X1 U961 ( .A(n1131), .B(n1249), .Z(n1248) );
NAND3_X1 U962 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1249) );
OR2_X1 U963 ( .A1(n1126), .A2(n1080), .ZN(n1252) );
NAND2_X1 U964 ( .A1(n1253), .A2(n1254), .ZN(n1251) );
INV_X1 U965 ( .A(KEYINPUT16), .ZN(n1254) );
NAND2_X1 U966 ( .A1(n1255), .A2(n1126), .ZN(n1253) );
XOR2_X1 U967 ( .A(KEYINPUT18), .B(n1076), .Z(n1255) );
NAND2_X1 U968 ( .A1(KEYINPUT16), .A2(n1256), .ZN(n1250) );
NAND2_X1 U969 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
OR2_X1 U970 ( .A1(n1080), .A2(KEYINPUT18), .ZN(n1258) );
NAND3_X1 U971 ( .A1(n1126), .A2(n1080), .A3(KEYINPUT18), .ZN(n1257) );
XNOR2_X1 U972 ( .A(n1079), .B(KEYINPUT43), .ZN(n1126) );
NAND3_X1 U973 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1131) );
NAND2_X1 U974 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
OR3_X1 U975 ( .A1(n1263), .A2(n1262), .A3(n1264), .ZN(n1260) );
INV_X1 U976 ( .A(KEYINPUT22), .ZN(n1263) );
NAND2_X1 U977 ( .A1(n1264), .A2(n1265), .ZN(n1259) );
NAND2_X1 U978 ( .A1(KEYINPUT22), .A2(n1266), .ZN(n1265) );
XOR2_X1 U979 ( .A(KEYINPUT47), .B(n1262), .Z(n1266) );
XNOR2_X1 U980 ( .A(n1216), .B(KEYINPUT52), .ZN(n1264) );
INV_X1 U981 ( .A(G113), .ZN(n1216) );
INV_X1 U982 ( .A(n1119), .ZN(n1179) );
NAND3_X1 U983 ( .A1(n1004), .A2(n1184), .A3(n1015), .ZN(n1119) );
AND2_X1 U984 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U985 ( .A1(G221), .A2(n1267), .ZN(n1017) );
INV_X1 U986 ( .A(n1217), .ZN(n1016) );
NAND3_X1 U987 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1217) );
NAND2_X1 U988 ( .A1(KEYINPUT60), .A2(n1060), .ZN(n1270) );
INV_X1 U989 ( .A(n1271), .ZN(n1060) );
OR3_X1 U990 ( .A1(n1272), .A2(KEYINPUT60), .A3(G469), .ZN(n1269) );
NAND2_X1 U991 ( .A1(G469), .A2(n1272), .ZN(n1268) );
NAND2_X1 U992 ( .A1(KEYINPUT23), .A2(n1271), .ZN(n1272) );
NAND2_X1 U993 ( .A1(n1273), .A2(n1220), .ZN(n1271) );
XOR2_X1 U994 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U995 ( .A(n1139), .B(n1276), .Z(n1275) );
NAND2_X1 U996 ( .A1(KEYINPUT14), .A2(n1277), .ZN(n1276) );
INV_X1 U997 ( .A(G140), .ZN(n1277) );
NAND2_X1 U998 ( .A1(n1278), .A2(n1020), .ZN(n1139) );
XOR2_X1 U999 ( .A(KEYINPUT28), .B(G227), .Z(n1278) );
XOR2_X1 U1000 ( .A(G110), .B(n1279), .Z(n1274) );
NOR2_X1 U1001 ( .A1(KEYINPUT38), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U1002 ( .A(n1150), .B(n1281), .ZN(n1280) );
XOR2_X1 U1003 ( .A(n1079), .B(n1076), .Z(n1281) );
INV_X1 U1004 ( .A(n1080), .ZN(n1076) );
XOR2_X1 U1005 ( .A(n1231), .B(n1282), .Z(n1080) );
XOR2_X1 U1006 ( .A(G137), .B(G134), .Z(n1282) );
INV_X1 U1007 ( .A(G131), .ZN(n1231) );
XOR2_X1 U1008 ( .A(G101), .B(n1283), .Z(n1150) );
NOR2_X1 U1009 ( .A1(KEYINPUT37), .A2(n1284), .ZN(n1283) );
XOR2_X1 U1010 ( .A(G104), .B(n984), .Z(n1284) );
INV_X1 U1011 ( .A(G107), .ZN(n984) );
NAND2_X1 U1012 ( .A1(n992), .A2(n1285), .ZN(n1184) );
NAND4_X1 U1013 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1096), .ZN(n1285) );
INV_X1 U1014 ( .A(G898), .ZN(n1096) );
NAND3_X1 U1015 ( .A1(n1206), .A2(n1020), .A3(G952), .ZN(n992) );
NAND2_X1 U1016 ( .A1(G237), .A2(G234), .ZN(n1206) );
AND2_X1 U1017 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1286), .ZN(n1006) );
XOR2_X1 U1019 ( .A(n1287), .B(n1054), .Z(n1005) );
INV_X1 U1020 ( .A(n1051), .ZN(n1054) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1286), .ZN(n1051) );
NAND2_X1 U1022 ( .A1(n1288), .A2(n1220), .ZN(n1286) );
INV_X1 U1023 ( .A(G237), .ZN(n1288) );
XNOR2_X1 U1024 ( .A(n1052), .B(KEYINPUT5), .ZN(n1287) );
AND2_X1 U1025 ( .A1(n1289), .A2(n1220), .ZN(n1052) );
XOR2_X1 U1026 ( .A(n1158), .B(n1290), .Z(n1289) );
XNOR2_X1 U1027 ( .A(n1162), .B(n1164), .ZN(n1290) );
XOR2_X1 U1028 ( .A(n1208), .B(n1079), .Z(n1164) );
XNOR2_X1 U1029 ( .A(G146), .B(n1241), .ZN(n1079) );
XNOR2_X1 U1030 ( .A(G128), .B(n1193), .ZN(n1241) );
INV_X1 U1031 ( .A(G143), .ZN(n1193) );
INV_X1 U1032 ( .A(G125), .ZN(n1208) );
NAND2_X1 U1033 ( .A1(G224), .A2(n1020), .ZN(n1162) );
XOR2_X1 U1034 ( .A(n1098), .B(n1099), .Z(n1158) );
XNOR2_X1 U1035 ( .A(G122), .B(G110), .ZN(n1099) );
XOR2_X1 U1036 ( .A(n1291), .B(n1292), .Z(n1098) );
XOR2_X1 U1037 ( .A(n1262), .B(n1293), .Z(n1292) );
XOR2_X1 U1038 ( .A(n1294), .B(n1295), .Z(n1293) );
NOR2_X1 U1039 ( .A1(G104), .A2(KEYINPUT39), .ZN(n1295) );
NOR2_X1 U1040 ( .A1(G113), .A2(KEYINPUT0), .ZN(n1294) );
XOR2_X1 U1041 ( .A(G119), .B(n1243), .Z(n1262) );
XOR2_X1 U1042 ( .A(G116), .B(KEYINPUT27), .Z(n1243) );
XNOR2_X1 U1043 ( .A(G101), .B(n1296), .ZN(n1291) );
XOR2_X1 U1044 ( .A(KEYINPUT3), .B(G107), .Z(n1296) );
XOR2_X1 U1045 ( .A(n1210), .B(KEYINPUT33), .Z(n1033) );
XNOR2_X1 U1046 ( .A(n1045), .B(n1043), .ZN(n1210) );
AND2_X1 U1047 ( .A1(n1297), .A2(n1267), .ZN(n1043) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1220), .ZN(n1267) );
INV_X1 U1049 ( .A(G902), .ZN(n1220) );
XNOR2_X1 U1050 ( .A(G217), .B(KEYINPUT48), .ZN(n1297) );
NOR2_X1 U1051 ( .A1(n1104), .A2(G902), .ZN(n1045) );
XOR2_X1 U1052 ( .A(n1298), .B(n1299), .Z(n1104) );
XOR2_X1 U1053 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U1054 ( .A(n1302), .B(KEYINPUT44), .Z(n1301) );
INV_X1 U1055 ( .A(G137), .ZN(n1302) );
NAND3_X1 U1056 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1300) );
OR2_X1 U1057 ( .A1(G110), .A2(KEYINPUT11), .ZN(n1305) );
NAND3_X1 U1058 ( .A1(KEYINPUT11), .A2(G110), .A3(n1306), .ZN(n1304) );
INV_X1 U1059 ( .A(n1307), .ZN(n1306) );
NAND2_X1 U1060 ( .A1(n1307), .A2(n1308), .ZN(n1303) );
NAND2_X1 U1061 ( .A1(KEYINPUT11), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1062 ( .A(KEYINPUT41), .B(G110), .Z(n1309) );
XNOR2_X1 U1063 ( .A(G119), .B(G128), .ZN(n1307) );
XOR2_X1 U1064 ( .A(n1310), .B(n1311), .Z(n1298) );
NOR2_X1 U1065 ( .A1(KEYINPUT6), .A2(n1225), .ZN(n1311) );
XOR2_X1 U1066 ( .A(G146), .B(n1072), .Z(n1225) );
XOR2_X1 U1067 ( .A(G125), .B(G140), .Z(n1072) );
NAND2_X1 U1068 ( .A1(n1239), .A2(G221), .ZN(n1310) );
AND2_X1 U1069 ( .A1(G234), .A2(n1020), .ZN(n1239) );
INV_X1 U1070 ( .A(G953), .ZN(n1020) );
endmodule


