//Key = 1000110000001001101110101101100010000001000001011011011011000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346;

XNOR2_X1 U744 ( .A(n1028), .B(n1029), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U746 ( .A1(G953), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR3_X1 U752 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1043) );
NOR2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR2_X1 U755 ( .A1(KEYINPUT62), .A2(n1052), .ZN(n1051) );
NOR2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1046) );
XNOR2_X1 U758 ( .A(KEYINPUT12), .B(n1057), .ZN(n1056) );
NOR2_X1 U759 ( .A1(n1058), .A2(n1057), .ZN(n1045) );
NOR3_X1 U760 ( .A1(n1049), .A2(n1059), .A3(n1057), .ZN(n1041) );
NOR2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR3_X1 U762 ( .A1(n1049), .A2(n1062), .A3(n1044), .ZN(n1037) );
NOR2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U764 ( .A1(n1065), .A2(n1057), .ZN(n1064) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
AND3_X1 U767 ( .A1(KEYINPUT62), .A2(n1040), .A3(n1070), .ZN(n1063) );
NOR3_X1 U768 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1030) );
AND4_X1 U769 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1032) );
NOR4_X1 U770 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
NOR2_X1 U771 ( .A1(n1079), .A2(n1068), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1080), .B(n1081), .Z(n1072) );
NOR2_X1 U773 ( .A1(KEYINPUT43), .A2(n1082), .ZN(n1081) );
XNOR2_X1 U774 ( .A(n1083), .B(KEYINPUT38), .ZN(n1080) );
XNOR2_X1 U775 ( .A(n1084), .B(G478), .ZN(n1071) );
XOR2_X1 U776 ( .A(n1085), .B(n1086), .Z(G72) );
NOR2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
AND2_X1 U778 ( .A1(G227), .A2(G900), .ZN(n1087) );
NAND2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1085) );
NAND3_X1 U780 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
INV_X1 U781 ( .A(n1094), .ZN(n1092) );
OR2_X1 U782 ( .A1(n1091), .A2(n1093), .ZN(n1089) );
NAND3_X1 U783 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1093) );
OR2_X1 U784 ( .A1(n1098), .A2(KEYINPUT32), .ZN(n1097) );
OR3_X1 U785 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1096) );
INV_X1 U786 ( .A(KEYINPUT32), .ZN(n1099) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1100), .ZN(n1095) );
NAND2_X1 U788 ( .A1(n1102), .A2(n1098), .ZN(n1100) );
XNOR2_X1 U789 ( .A(KEYINPUT52), .B(KEYINPUT42), .ZN(n1102) );
XNOR2_X1 U790 ( .A(n1103), .B(n1104), .ZN(n1101) );
XOR2_X1 U791 ( .A(KEYINPUT46), .B(G140), .Z(n1104) );
NAND2_X1 U792 ( .A1(KEYINPUT15), .A2(G125), .ZN(n1103) );
NAND2_X1 U793 ( .A1(n1088), .A2(n1105), .ZN(n1091) );
NAND4_X1 U794 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1105) );
NOR2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U799 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XNOR2_X1 U800 ( .A(n1119), .B(n1120), .ZN(n1116) );
NAND2_X1 U801 ( .A1(KEYINPUT47), .A2(n1121), .ZN(n1119) );
NAND2_X1 U802 ( .A1(G953), .A2(n1122), .ZN(n1114) );
NAND2_X1 U803 ( .A1(G224), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U804 ( .A(KEYINPUT44), .B(n1118), .ZN(n1123) );
NOR2_X1 U805 ( .A1(n1124), .A2(G953), .ZN(n1112) );
NOR2_X1 U806 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XOR2_X1 U807 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U808 ( .A(KEYINPUT9), .B(n1129), .Z(n1128) );
NOR2_X1 U809 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1132), .ZN(G63) );
NOR3_X1 U811 ( .A1(n1084), .A2(n1133), .A3(n1134), .ZN(n1132) );
NOR3_X1 U812 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
AND2_X1 U813 ( .A1(n1135), .A2(n1137), .ZN(n1133) );
NAND2_X1 U814 ( .A1(n1138), .A2(G478), .ZN(n1137) );
XOR2_X1 U815 ( .A(n1034), .B(KEYINPUT63), .Z(n1138) );
INV_X1 U816 ( .A(n1139), .ZN(n1084) );
NOR2_X1 U817 ( .A1(n1125), .A2(n1140), .ZN(G60) );
NOR3_X1 U818 ( .A1(n1083), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR3_X1 U819 ( .A1(n1143), .A2(n1082), .A3(n1131), .ZN(n1142) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
AND2_X1 U821 ( .A1(n1034), .A2(G475), .ZN(n1144) );
XOR2_X1 U822 ( .A(G104), .B(n1146), .Z(G6) );
NOR2_X1 U823 ( .A1(n1125), .A2(n1147), .ZN(G57) );
XOR2_X1 U824 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U825 ( .A(n1150), .B(n1151), .ZN(n1149) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1150) );
NAND2_X1 U827 ( .A1(KEYINPUT56), .A2(n1154), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1148) );
NOR2_X1 U829 ( .A1(n1157), .A2(n1131), .ZN(n1156) );
XOR2_X1 U830 ( .A(n1158), .B(G101), .Z(n1155) );
NAND2_X1 U831 ( .A1(KEYINPUT57), .A2(n1159), .ZN(n1158) );
NOR2_X1 U832 ( .A1(n1125), .A2(n1160), .ZN(G54) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U834 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U835 ( .A1(KEYINPUT25), .A2(n1165), .ZN(n1163) );
XOR2_X1 U836 ( .A(n1166), .B(n1167), .Z(n1161) );
NOR2_X1 U837 ( .A1(n1168), .A2(n1131), .ZN(n1167) );
XNOR2_X1 U838 ( .A(G140), .B(KEYINPUT6), .ZN(n1166) );
AND2_X1 U839 ( .A1(G953), .A2(n1169), .ZN(n1125) );
XOR2_X1 U840 ( .A(KEYINPUT24), .B(G952), .Z(n1169) );
NOR2_X1 U841 ( .A1(n1170), .A2(n1171), .ZN(G51) );
XOR2_X1 U842 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U843 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U844 ( .A1(n1176), .A2(n1131), .ZN(n1175) );
NAND2_X1 U845 ( .A1(G902), .A2(n1034), .ZN(n1131) );
NAND4_X1 U846 ( .A1(n1177), .A2(n1124), .A3(n1178), .A4(n1179), .ZN(n1034) );
AND3_X1 U847 ( .A1(n1180), .A2(n1107), .A3(n1108), .ZN(n1179) );
NAND2_X1 U848 ( .A1(n1181), .A2(n1182), .ZN(n1108) );
XNOR2_X1 U849 ( .A(n1183), .B(KEYINPUT16), .ZN(n1181) );
INV_X1 U850 ( .A(n1110), .ZN(n1180) );
NOR2_X1 U851 ( .A1(n1184), .A2(n1057), .ZN(n1110) );
INV_X1 U852 ( .A(n1185), .ZN(n1184) );
XOR2_X1 U853 ( .A(n1111), .B(KEYINPUT5), .Z(n1178) );
NAND4_X1 U854 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1111) );
NAND2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
XOR2_X1 U856 ( .A(n1192), .B(KEYINPUT22), .Z(n1190) );
NAND2_X1 U857 ( .A1(n1182), .A2(n1193), .ZN(n1186) );
INV_X1 U858 ( .A(n1194), .ZN(n1182) );
AND4_X1 U859 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1124) );
NOR4_X1 U860 ( .A1(n1029), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1198) );
NOR3_X1 U861 ( .A1(n1202), .A2(n1058), .A3(n1203), .ZN(n1201) );
NOR3_X1 U862 ( .A1(n1049), .A2(n1204), .A3(n1205), .ZN(n1200) );
NOR3_X1 U863 ( .A1(n1205), .A2(n1044), .A3(n1058), .ZN(n1029) );
NOR2_X1 U864 ( .A1(n1206), .A2(n1146), .ZN(n1197) );
NOR3_X1 U865 ( .A1(n1205), .A2(n1044), .A3(n1055), .ZN(n1146) );
INV_X1 U866 ( .A(n1207), .ZN(n1044) );
XOR2_X1 U867 ( .A(n1106), .B(KEYINPUT59), .Z(n1177) );
NAND2_X1 U868 ( .A1(KEYINPUT54), .A2(n1208), .ZN(n1174) );
XOR2_X1 U869 ( .A(n1209), .B(n1210), .Z(n1172) );
NOR2_X1 U870 ( .A1(KEYINPUT60), .A2(n1211), .ZN(n1210) );
XOR2_X1 U871 ( .A(n1120), .B(n1121), .Z(n1211) );
NOR2_X1 U872 ( .A1(n1212), .A2(n1213), .ZN(n1170) );
XNOR2_X1 U873 ( .A(G953), .B(KEYINPUT33), .ZN(n1213) );
XNOR2_X1 U874 ( .A(KEYINPUT24), .B(G952), .ZN(n1212) );
XOR2_X1 U875 ( .A(G146), .B(n1214), .Z(G48) );
NOR2_X1 U876 ( .A1(n1055), .A2(n1194), .ZN(n1214) );
XNOR2_X1 U877 ( .A(G143), .B(n1106), .ZN(G45) );
NAND4_X1 U878 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1106) );
NOR2_X1 U879 ( .A1(n1219), .A2(n1202), .ZN(n1218) );
XNOR2_X1 U880 ( .A(G140), .B(n1220), .ZN(G42) );
NAND2_X1 U881 ( .A1(n1221), .A2(n1191), .ZN(n1220) );
XNOR2_X1 U882 ( .A(n1185), .B(KEYINPUT45), .ZN(n1221) );
NOR3_X1 U883 ( .A1(n1222), .A2(n1204), .A3(n1055), .ZN(n1185) );
XOR2_X1 U884 ( .A(G137), .B(n1223), .Z(G39) );
NOR2_X1 U885 ( .A1(KEYINPUT34), .A2(n1107), .ZN(n1223) );
NAND3_X1 U886 ( .A1(n1224), .A2(n1191), .A3(n1225), .ZN(n1107) );
NOR3_X1 U887 ( .A1(n1222), .A2(n1226), .A3(n1227), .ZN(n1225) );
XNOR2_X1 U888 ( .A(G134), .B(n1188), .ZN(G36) );
NAND4_X1 U889 ( .A1(n1060), .A2(n1191), .A3(n1228), .A4(n1193), .ZN(n1188) );
XOR2_X1 U890 ( .A(G131), .B(n1229), .Z(G33) );
NOR2_X1 U891 ( .A1(n1057), .A2(n1192), .ZN(n1229) );
NAND3_X1 U892 ( .A1(n1183), .A2(n1228), .A3(n1060), .ZN(n1192) );
INV_X1 U893 ( .A(n1222), .ZN(n1228) );
NAND2_X1 U894 ( .A1(n1067), .A2(n1215), .ZN(n1222) );
INV_X1 U895 ( .A(n1191), .ZN(n1057) );
NOR2_X1 U896 ( .A1(n1054), .A2(n1075), .ZN(n1191) );
INV_X1 U897 ( .A(n1053), .ZN(n1075) );
XOR2_X1 U898 ( .A(n1079), .B(KEYINPUT3), .Z(n1054) );
XOR2_X1 U899 ( .A(G128), .B(n1230), .Z(G30) );
NOR2_X1 U900 ( .A1(n1058), .A2(n1194), .ZN(n1230) );
NAND4_X1 U901 ( .A1(n1231), .A2(n1232), .A3(n1078), .A4(n1215), .ZN(n1194) );
XOR2_X1 U902 ( .A(G101), .B(n1206), .Z(G3) );
NOR3_X1 U903 ( .A1(n1049), .A2(n1205), .A3(n1202), .ZN(n1206) );
INV_X1 U904 ( .A(n1060), .ZN(n1202) );
NAND2_X1 U905 ( .A1(n1232), .A2(n1233), .ZN(n1205) );
INV_X1 U906 ( .A(n1224), .ZN(n1049) );
XNOR2_X1 U907 ( .A(G125), .B(n1189), .ZN(G27) );
NAND3_X1 U908 ( .A1(n1183), .A2(n1234), .A3(n1235), .ZN(n1189) );
AND3_X1 U909 ( .A1(n1061), .A2(n1215), .A3(n1070), .ZN(n1235) );
NAND2_X1 U910 ( .A1(n1236), .A2(n1237), .ZN(n1215) );
NAND3_X1 U911 ( .A1(G902), .A2(n1238), .A3(n1094), .ZN(n1237) );
NOR2_X1 U912 ( .A1(n1088), .A2(G900), .ZN(n1094) );
XNOR2_X1 U913 ( .A(KEYINPUT20), .B(n1036), .ZN(n1236) );
XOR2_X1 U914 ( .A(n1199), .B(n1239), .Z(G24) );
NOR2_X1 U915 ( .A1(KEYINPUT17), .A2(n1240), .ZN(n1239) );
AND4_X1 U916 ( .A1(n1241), .A2(n1207), .A3(n1217), .A4(n1216), .ZN(n1199) );
NAND2_X1 U917 ( .A1(n1242), .A2(n1243), .ZN(n1207) );
OR2_X1 U918 ( .A1(n1204), .A2(KEYINPUT28), .ZN(n1243) );
INV_X1 U919 ( .A(n1061), .ZN(n1204) );
NAND3_X1 U920 ( .A1(n1227), .A2(n1226), .A3(KEYINPUT28), .ZN(n1242) );
XOR2_X1 U921 ( .A(n1195), .B(n1244), .Z(G21) );
XNOR2_X1 U922 ( .A(G119), .B(KEYINPUT23), .ZN(n1244) );
NAND4_X1 U923 ( .A1(n1241), .A2(n1224), .A3(n1231), .A4(n1078), .ZN(n1195) );
XNOR2_X1 U924 ( .A(G116), .B(n1245), .ZN(G18) );
NAND3_X1 U925 ( .A1(n1241), .A2(n1246), .A3(n1060), .ZN(n1245) );
XNOR2_X1 U926 ( .A(KEYINPUT29), .B(n1058), .ZN(n1246) );
INV_X1 U927 ( .A(n1193), .ZN(n1058) );
NOR2_X1 U928 ( .A1(n1216), .A2(n1247), .ZN(n1193) );
XOR2_X1 U929 ( .A(n1196), .B(n1248), .Z(G15) );
XOR2_X1 U930 ( .A(KEYINPUT53), .B(G113), .Z(n1248) );
NAND3_X1 U931 ( .A1(n1183), .A2(n1241), .A3(n1060), .ZN(n1196) );
NOR2_X1 U932 ( .A1(n1227), .A2(n1078), .ZN(n1060) );
INV_X1 U933 ( .A(n1203), .ZN(n1241) );
NAND3_X1 U934 ( .A1(n1070), .A2(n1233), .A3(n1234), .ZN(n1203) );
INV_X1 U935 ( .A(n1040), .ZN(n1234) );
NAND2_X1 U936 ( .A1(n1249), .A2(n1069), .ZN(n1040) );
XNOR2_X1 U937 ( .A(n1068), .B(KEYINPUT2), .ZN(n1249) );
INV_X1 U938 ( .A(n1055), .ZN(n1183) );
NAND2_X1 U939 ( .A1(n1247), .A2(n1216), .ZN(n1055) );
INV_X1 U940 ( .A(n1217), .ZN(n1247) );
XNOR2_X1 U941 ( .A(G110), .B(n1250), .ZN(G12) );
NAND4_X1 U942 ( .A1(n1251), .A2(n1224), .A3(n1061), .A4(n1232), .ZN(n1250) );
INV_X1 U943 ( .A(n1219), .ZN(n1232) );
NAND2_X1 U944 ( .A1(n1067), .A2(n1070), .ZN(n1219) );
INV_X1 U945 ( .A(n1052), .ZN(n1070) );
NAND2_X1 U946 ( .A1(n1252), .A2(n1079), .ZN(n1052) );
XOR2_X1 U947 ( .A(n1253), .B(n1176), .Z(n1079) );
NAND2_X1 U948 ( .A1(G210), .A2(n1254), .ZN(n1176) );
NAND2_X1 U949 ( .A1(n1255), .A2(n1136), .ZN(n1253) );
XOR2_X1 U950 ( .A(n1256), .B(n1208), .Z(n1255) );
XNOR2_X1 U951 ( .A(G125), .B(n1151), .ZN(n1208) );
XNOR2_X1 U952 ( .A(n1257), .B(n1209), .ZN(n1256) );
NAND2_X1 U953 ( .A1(G224), .A2(n1088), .ZN(n1209) );
NAND2_X1 U954 ( .A1(n1258), .A2(KEYINPUT27), .ZN(n1257) );
XNOR2_X1 U955 ( .A(n1121), .B(n1120), .ZN(n1258) );
XOR2_X1 U956 ( .A(n1153), .B(n1259), .Z(n1120) );
XNOR2_X1 U957 ( .A(n1240), .B(G110), .ZN(n1259) );
NAND2_X1 U958 ( .A1(n1260), .A2(n1261), .ZN(n1121) );
NAND2_X1 U959 ( .A1(n1262), .A2(G107), .ZN(n1261) );
NAND2_X1 U960 ( .A1(n1263), .A2(n1028), .ZN(n1260) );
XNOR2_X1 U961 ( .A(n1262), .B(KEYINPUT35), .ZN(n1263) );
XNOR2_X1 U962 ( .A(KEYINPUT4), .B(n1053), .ZN(n1252) );
NAND2_X1 U963 ( .A1(G214), .A2(n1254), .ZN(n1053) );
NAND2_X1 U964 ( .A1(n1264), .A2(n1136), .ZN(n1254) );
NOR2_X1 U965 ( .A1(n1265), .A2(n1076), .ZN(n1067) );
INV_X1 U966 ( .A(n1069), .ZN(n1076) );
NAND2_X1 U967 ( .A1(G221), .A2(n1266), .ZN(n1069) );
INV_X1 U968 ( .A(n1068), .ZN(n1265) );
XOR2_X1 U969 ( .A(n1267), .B(n1168), .Z(n1068) );
INV_X1 U970 ( .A(G469), .ZN(n1168) );
NAND2_X1 U971 ( .A1(n1268), .A2(n1136), .ZN(n1267) );
XOR2_X1 U972 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U973 ( .A(n1164), .B(n1165), .ZN(n1270) );
XOR2_X1 U974 ( .A(n1271), .B(n1272), .Z(n1164) );
XOR2_X1 U975 ( .A(n1262), .B(n1098), .Z(n1272) );
XOR2_X1 U976 ( .A(n1273), .B(n1274), .Z(n1098) );
XNOR2_X1 U977 ( .A(n1275), .B(n1276), .ZN(n1274) );
NAND2_X1 U978 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
OR2_X1 U979 ( .A1(n1279), .A2(G146), .ZN(n1278) );
XOR2_X1 U980 ( .A(n1280), .B(KEYINPUT36), .Z(n1277) );
NAND2_X1 U981 ( .A1(G146), .A2(n1279), .ZN(n1280) );
INV_X1 U982 ( .A(G143), .ZN(n1279) );
XOR2_X1 U983 ( .A(G104), .B(G101), .Z(n1262) );
XOR2_X1 U984 ( .A(n1281), .B(n1282), .Z(n1271) );
XNOR2_X1 U985 ( .A(KEYINPUT10), .B(n1028), .ZN(n1282) );
NAND2_X1 U986 ( .A1(G227), .A2(n1088), .ZN(n1281) );
XOR2_X1 U987 ( .A(n1283), .B(G140), .Z(n1269) );
XNOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT30), .ZN(n1283) );
NOR2_X1 U989 ( .A1(n1226), .A2(n1231), .ZN(n1061) );
INV_X1 U990 ( .A(n1227), .ZN(n1231) );
XOR2_X1 U991 ( .A(n1077), .B(KEYINPUT51), .Z(n1227) );
XOR2_X1 U992 ( .A(n1284), .B(n1157), .Z(n1077) );
INV_X1 U993 ( .A(G472), .ZN(n1157) );
NAND2_X1 U994 ( .A1(n1285), .A2(n1136), .ZN(n1284) );
XOR2_X1 U995 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U996 ( .A(G101), .B(n1154), .ZN(n1287) );
AND3_X1 U997 ( .A1(G210), .A2(n1264), .A3(n1288), .ZN(n1154) );
XNOR2_X1 U998 ( .A(G953), .B(KEYINPUT58), .ZN(n1288) );
NAND2_X1 U999 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
NAND2_X1 U1000 ( .A1(n1291), .A2(n1153), .ZN(n1290) );
XOR2_X1 U1001 ( .A(n1292), .B(KEYINPUT41), .Z(n1289) );
OR2_X1 U1002 ( .A1(n1153), .A2(n1291), .ZN(n1292) );
AND2_X1 U1003 ( .A1(n1293), .A2(n1294), .ZN(n1291) );
NAND2_X1 U1004 ( .A1(n1151), .A2(n1159), .ZN(n1294) );
XOR2_X1 U1005 ( .A(n1295), .B(KEYINPUT7), .Z(n1293) );
OR2_X1 U1006 ( .A1(n1159), .A2(n1151), .ZN(n1295) );
XOR2_X1 U1007 ( .A(n1296), .B(n1297), .Z(n1151) );
XOR2_X1 U1008 ( .A(G128), .B(n1298), .Z(n1297) );
NOR2_X1 U1009 ( .A1(G146), .A2(KEYINPUT1), .ZN(n1298) );
XNOR2_X1 U1010 ( .A(G143), .B(KEYINPUT37), .ZN(n1296) );
XOR2_X1 U1011 ( .A(G137), .B(n1276), .Z(n1159) );
XOR2_X1 U1012 ( .A(G131), .B(G134), .Z(n1276) );
XOR2_X1 U1013 ( .A(G113), .B(n1299), .Z(n1153) );
XOR2_X1 U1014 ( .A(G119), .B(G116), .Z(n1299) );
INV_X1 U1015 ( .A(n1078), .ZN(n1226) );
XOR2_X1 U1016 ( .A(n1300), .B(n1130), .Z(n1078) );
NAND2_X1 U1017 ( .A1(G217), .A2(n1266), .ZN(n1130) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1136), .ZN(n1266) );
OR2_X1 U1019 ( .A1(n1127), .A2(G902), .ZN(n1300) );
XNOR2_X1 U1020 ( .A(n1301), .B(n1302), .ZN(n1127) );
XOR2_X1 U1021 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1022 ( .A(n1165), .B(n1305), .ZN(n1304) );
AND3_X1 U1023 ( .A1(G221), .A2(n1088), .A3(G234), .ZN(n1305) );
INV_X1 U1024 ( .A(G110), .ZN(n1165) );
NOR2_X1 U1025 ( .A1(G119), .A2(KEYINPUT8), .ZN(n1303) );
XOR2_X1 U1026 ( .A(n1306), .B(n1273), .Z(n1301) );
XOR2_X1 U1027 ( .A(G137), .B(G128), .Z(n1273) );
NOR2_X1 U1028 ( .A1(n1217), .A2(n1216), .ZN(n1224) );
NAND3_X1 U1029 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1216) );
NAND2_X1 U1030 ( .A1(KEYINPUT40), .A2(n1083), .ZN(n1309) );
NAND3_X1 U1031 ( .A1(n1310), .A2(n1311), .A3(G475), .ZN(n1308) );
INV_X1 U1032 ( .A(n1083), .ZN(n1310) );
NAND2_X1 U1033 ( .A1(n1312), .A2(n1082), .ZN(n1307) );
INV_X1 U1034 ( .A(G475), .ZN(n1082) );
NAND2_X1 U1035 ( .A1(n1313), .A2(n1311), .ZN(n1312) );
INV_X1 U1036 ( .A(KEYINPUT40), .ZN(n1311) );
XNOR2_X1 U1037 ( .A(n1083), .B(KEYINPUT61), .ZN(n1313) );
NOR2_X1 U1038 ( .A1(n1145), .A2(G902), .ZN(n1083) );
INV_X1 U1039 ( .A(n1143), .ZN(n1145) );
XNOR2_X1 U1040 ( .A(n1314), .B(n1315), .ZN(n1143) );
XOR2_X1 U1041 ( .A(G104), .B(n1316), .Z(n1315) );
NOR2_X1 U1042 ( .A1(KEYINPUT11), .A2(n1317), .ZN(n1316) );
XOR2_X1 U1043 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1044 ( .A(n1320), .B(n1321), .Z(n1319) );
AND3_X1 U1045 ( .A1(G214), .A2(n1088), .A3(n1264), .ZN(n1321) );
INV_X1 U1046 ( .A(G237), .ZN(n1264) );
NAND2_X1 U1047 ( .A1(n1322), .A2(KEYINPUT0), .ZN(n1320) );
XOR2_X1 U1048 ( .A(n1306), .B(KEYINPUT14), .Z(n1322) );
XNOR2_X1 U1049 ( .A(G125), .B(n1323), .ZN(n1306) );
XOR2_X1 U1050 ( .A(G146), .B(G140), .Z(n1323) );
XNOR2_X1 U1051 ( .A(G131), .B(G143), .ZN(n1318) );
NAND2_X1 U1052 ( .A1(KEYINPUT39), .A2(n1324), .ZN(n1314) );
XNOR2_X1 U1053 ( .A(n1240), .B(G113), .ZN(n1324) );
XOR2_X1 U1054 ( .A(G478), .B(n1325), .Z(n1217) );
NOR2_X1 U1055 ( .A1(KEYINPUT31), .A2(n1326), .ZN(n1325) );
XNOR2_X1 U1056 ( .A(KEYINPUT19), .B(n1139), .ZN(n1326) );
NAND2_X1 U1057 ( .A1(n1136), .A2(n1135), .ZN(n1139) );
NAND2_X1 U1058 ( .A1(n1327), .A2(n1328), .ZN(n1135) );
NAND4_X1 U1059 ( .A1(G234), .A2(G217), .A3(n1329), .A4(n1088), .ZN(n1328) );
XOR2_X1 U1060 ( .A(n1330), .B(KEYINPUT55), .Z(n1327) );
NAND2_X1 U1061 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND3_X1 U1062 ( .A1(G217), .A2(n1088), .A3(G234), .ZN(n1332) );
INV_X1 U1063 ( .A(n1329), .ZN(n1331) );
XNOR2_X1 U1064 ( .A(n1333), .B(n1334), .ZN(n1329) );
XNOR2_X1 U1065 ( .A(n1028), .B(n1335), .ZN(n1334) );
NOR2_X1 U1066 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1067 ( .A(KEYINPUT21), .B(n1338), .Z(n1337) );
NOR2_X1 U1068 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
AND2_X1 U1069 ( .A1(n1340), .A2(n1339), .ZN(n1336) );
XOR2_X1 U1070 ( .A(G134), .B(KEYINPUT26), .Z(n1339) );
NAND2_X1 U1071 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
OR2_X1 U1072 ( .A1(n1343), .A2(G128), .ZN(n1342) );
XOR2_X1 U1073 ( .A(n1344), .B(KEYINPUT13), .Z(n1341) );
NAND2_X1 U1074 ( .A1(G128), .A2(n1343), .ZN(n1344) );
XOR2_X1 U1075 ( .A(G143), .B(KEYINPUT50), .Z(n1343) );
INV_X1 U1076 ( .A(G107), .ZN(n1028) );
XNOR2_X1 U1077 ( .A(G116), .B(n1345), .ZN(n1333) );
XNOR2_X1 U1078 ( .A(KEYINPUT18), .B(n1240), .ZN(n1345) );
INV_X1 U1079 ( .A(G122), .ZN(n1240) );
INV_X1 U1080 ( .A(G902), .ZN(n1136) );
XOR2_X1 U1081 ( .A(n1233), .B(KEYINPUT49), .Z(n1251) );
NAND2_X1 U1082 ( .A1(n1036), .A2(n1346), .ZN(n1233) );
NAND4_X1 U1083 ( .A1(G953), .A2(G902), .A3(n1238), .A4(n1118), .ZN(n1346) );
INV_X1 U1084 ( .A(G898), .ZN(n1118) );
NAND3_X1 U1085 ( .A1(n1238), .A2(n1088), .A3(G952), .ZN(n1036) );
INV_X1 U1086 ( .A(G953), .ZN(n1088) );
NAND2_X1 U1087 ( .A1(G237), .A2(G234), .ZN(n1238) );
endmodule


