//Key = 0101001000001001001100000110101101111110100011001000011000110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308;

XOR2_X1 U713 ( .A(n984), .B(n985), .Z(G9) );
NOR2_X1 U714 ( .A1(KEYINPUT4), .A2(n986), .ZN(n985) );
XOR2_X1 U715 ( .A(KEYINPUT24), .B(G107), .Z(n986) );
NOR2_X1 U716 ( .A1(n987), .A2(n988), .ZN(G75) );
XOR2_X1 U717 ( .A(KEYINPUT22), .B(n989), .Z(n988) );
AND3_X1 U718 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n989) );
NOR4_X1 U719 ( .A1(n993), .A2(n994), .A3(n995), .A4(n992), .ZN(n987) );
INV_X1 U720 ( .A(G952), .ZN(n992) );
NOR2_X1 U721 ( .A1(n996), .A2(n997), .ZN(n995) );
NOR2_X1 U722 ( .A1(n998), .A2(n999), .ZN(n996) );
XOR2_X1 U723 ( .A(KEYINPUT63), .B(n1000), .Z(n999) );
NOR4_X1 U724 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
XOR2_X1 U725 ( .A(n1005), .B(KEYINPUT17), .Z(n1001) );
NOR3_X1 U726 ( .A1(n1004), .A2(n1006), .A3(n1005), .ZN(n998) );
NOR2_X1 U727 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NOR2_X1 U728 ( .A1(n1002), .A2(n1009), .ZN(n1008) );
NOR2_X1 U729 ( .A1(n1010), .A2(n1011), .ZN(n1007) );
NOR2_X1 U730 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NAND3_X1 U731 ( .A1(n990), .A2(n991), .A3(n1014), .ZN(n993) );
NAND4_X1 U732 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1014) );
NOR2_X1 U733 ( .A1(n1011), .A2(n1002), .ZN(n1018) );
INV_X1 U734 ( .A(n1004), .ZN(n1017) );
NAND2_X1 U735 ( .A1(n1019), .A2(n1005), .ZN(n1016) );
NAND2_X1 U736 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U737 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
INV_X1 U738 ( .A(n997), .ZN(n1020) );
NAND3_X1 U739 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1015) );
NAND2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
INV_X1 U741 ( .A(n1029), .ZN(n1024) );
NAND4_X1 U742 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n990) );
NOR4_X1 U743 ( .A1(n1002), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1033) );
XOR2_X1 U744 ( .A(KEYINPUT11), .B(n1037), .Z(n1036) );
XOR2_X1 U745 ( .A(KEYINPUT27), .B(n1038), .Z(n1035) );
XOR2_X1 U746 ( .A(KEYINPUT47), .B(n1039), .Z(n1034) );
NOR2_X1 U747 ( .A1(G469), .A2(n1040), .ZN(n1039) );
NOR2_X1 U748 ( .A1(n1027), .A2(n1041), .ZN(n1032) );
AND2_X1 U749 ( .A1(n1040), .A2(G469), .ZN(n1041) );
XOR2_X1 U750 ( .A(G472), .B(n1042), .Z(n1031) );
NOR2_X1 U751 ( .A1(n1043), .A2(KEYINPUT57), .ZN(n1042) );
XOR2_X1 U752 ( .A(KEYINPUT1), .B(n1022), .Z(n1030) );
NAND3_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(G72) );
NAND2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
OR3_X1 U755 ( .A1(n1048), .A2(n1047), .A3(n1049), .ZN(n1045) );
INV_X1 U756 ( .A(KEYINPUT44), .ZN(n1048) );
NAND2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1044) );
NAND2_X1 U758 ( .A1(KEYINPUT44), .A2(n1051), .ZN(n1050) );
XNOR2_X1 U759 ( .A(KEYINPUT7), .B(n1047), .ZN(n1051) );
NAND2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1047) );
NAND2_X1 U761 ( .A1(G227), .A2(n1054), .ZN(n1053) );
XOR2_X1 U762 ( .A(KEYINPUT8), .B(G900), .Z(n1054) );
XOR2_X1 U763 ( .A(KEYINPUT10), .B(G953), .Z(n1052) );
XNOR2_X1 U764 ( .A(n1055), .B(n1056), .ZN(n1049) );
NOR2_X1 U765 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
XOR2_X1 U766 ( .A(n1059), .B(n1060), .Z(n1058) );
XOR2_X1 U767 ( .A(n1061), .B(n1062), .Z(n1060) );
XOR2_X1 U768 ( .A(n1063), .B(n1064), .Z(n1059) );
NOR2_X1 U769 ( .A1(KEYINPUT9), .A2(n1065), .ZN(n1064) );
NOR2_X1 U770 ( .A1(G900), .A2(n991), .ZN(n1057) );
NAND2_X1 U771 ( .A1(n1066), .A2(n991), .ZN(n1055) );
XOR2_X1 U772 ( .A(KEYINPUT15), .B(n1067), .Z(n1066) );
XOR2_X1 U773 ( .A(n1068), .B(n1069), .Z(G69) );
NOR2_X1 U774 ( .A1(n1070), .A2(n991), .ZN(n1069) );
NOR2_X1 U775 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U776 ( .A1(KEYINPUT49), .A2(n1073), .ZN(n1068) );
XOR2_X1 U777 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U778 ( .A1(n1076), .A2(G953), .ZN(n1075) );
NOR2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U780 ( .A(KEYINPUT33), .B(n1079), .Z(n1078) );
NAND2_X1 U781 ( .A1(n1080), .A2(n1081), .ZN(n1074) );
NAND2_X1 U782 ( .A1(G953), .A2(n1072), .ZN(n1081) );
XOR2_X1 U783 ( .A(n1082), .B(n1083), .Z(n1080) );
XOR2_X1 U784 ( .A(G122), .B(n1084), .Z(n1083) );
NOR2_X1 U785 ( .A1(KEYINPUT16), .A2(n1085), .ZN(n1084) );
XOR2_X1 U786 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U787 ( .A1(n1088), .A2(n1089), .ZN(G66) );
XOR2_X1 U788 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U789 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR2_X1 U790 ( .A1(n1088), .A2(n1094), .ZN(G63) );
XOR2_X1 U791 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND3_X1 U792 ( .A1(n1097), .A2(n1098), .A3(G478), .ZN(n1095) );
NAND2_X1 U793 ( .A1(KEYINPUT40), .A2(n1093), .ZN(n1098) );
NAND2_X1 U794 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
INV_X1 U795 ( .A(KEYINPUT40), .ZN(n1100) );
OR2_X1 U796 ( .A1(n994), .A2(n1101), .ZN(n1099) );
NOR2_X1 U797 ( .A1(n1088), .A2(n1102), .ZN(G60) );
XNOR2_X1 U798 ( .A(n1103), .B(n1104), .ZN(n1102) );
NOR2_X1 U799 ( .A1(n1105), .A2(n1093), .ZN(n1104) );
INV_X1 U800 ( .A(G475), .ZN(n1105) );
XOR2_X1 U801 ( .A(G104), .B(n1106), .Z(G6) );
NOR2_X1 U802 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U803 ( .A1(n1088), .A2(n1109), .ZN(G57) );
XOR2_X1 U804 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U805 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR2_X1 U806 ( .A1(n1114), .A2(n1093), .ZN(n1113) );
INV_X1 U807 ( .A(G472), .ZN(n1114) );
XOR2_X1 U808 ( .A(n1115), .B(n1116), .Z(n1110) );
XNOR2_X1 U809 ( .A(n1117), .B(KEYINPUT0), .ZN(n1116) );
NAND2_X1 U810 ( .A1(KEYINPUT28), .A2(n1118), .ZN(n1117) );
NAND2_X1 U811 ( .A1(KEYINPUT35), .A2(n1119), .ZN(n1115) );
INV_X1 U812 ( .A(n1120), .ZN(n1119) );
NOR2_X1 U813 ( .A1(n1088), .A2(n1121), .ZN(G54) );
XOR2_X1 U814 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U815 ( .A1(n1124), .A2(n1093), .ZN(n1123) );
NAND3_X1 U816 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1122) );
NAND2_X1 U817 ( .A1(KEYINPUT56), .A2(n1128), .ZN(n1127) );
NAND3_X1 U818 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1126) );
INV_X1 U819 ( .A(KEYINPUT56), .ZN(n1130) );
OR2_X1 U820 ( .A1(n1131), .A2(n1129), .ZN(n1125) );
NOR2_X1 U821 ( .A1(n1132), .A2(n1128), .ZN(n1129) );
XNOR2_X1 U822 ( .A(n1133), .B(n1134), .ZN(n1128) );
XOR2_X1 U823 ( .A(KEYINPUT60), .B(n1135), .Z(n1134) );
INV_X1 U824 ( .A(KEYINPUT61), .ZN(n1132) );
NOR2_X1 U825 ( .A1(n1088), .A2(n1136), .ZN(G51) );
XNOR2_X1 U826 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U827 ( .A1(n1139), .A2(n1093), .ZN(n1138) );
NAND2_X1 U828 ( .A1(G902), .A2(n994), .ZN(n1093) );
NAND3_X1 U829 ( .A1(n1079), .A2(n1067), .A3(n1140), .ZN(n994) );
XOR2_X1 U830 ( .A(n1077), .B(KEYINPUT59), .Z(n1140) );
NAND4_X1 U831 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1077) );
OR2_X1 U832 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
NAND2_X1 U833 ( .A1(n1147), .A2(n1029), .ZN(n1141) );
XOR2_X1 U834 ( .A(n1148), .B(KEYINPUT31), .Z(n1147) );
NAND3_X1 U835 ( .A1(n1026), .A2(n1149), .A3(n1150), .ZN(n1148) );
XOR2_X1 U836 ( .A(KEYINPUT54), .B(n1151), .Z(n1149) );
AND4_X1 U837 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1067) );
NOR4_X1 U838 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NOR3_X1 U839 ( .A1(n1005), .A2(n1160), .A3(n1161), .ZN(n1159) );
INV_X1 U840 ( .A(n1162), .ZN(n1158) );
NAND2_X1 U841 ( .A1(n1163), .A2(n1164), .ZN(n1153) );
NAND2_X1 U842 ( .A1(n1165), .A2(n1146), .ZN(n1164) );
XOR2_X1 U843 ( .A(KEYINPUT58), .B(n1012), .Z(n1165) );
INV_X1 U844 ( .A(n1166), .ZN(n1163) );
NAND2_X1 U845 ( .A1(n1150), .A2(n1167), .ZN(n1152) );
AND3_X1 U846 ( .A1(n1168), .A2(n984), .A3(n1169), .ZN(n1079) );
NAND2_X1 U847 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XNOR2_X1 U848 ( .A(KEYINPUT13), .B(n1108), .ZN(n1171) );
NAND3_X1 U849 ( .A1(n1013), .A2(n1172), .A3(n1173), .ZN(n1108) );
NOR3_X1 U850 ( .A1(n1174), .A2(n1151), .A3(n1022), .ZN(n1173) );
NAND3_X1 U851 ( .A1(n1012), .A2(n1172), .A3(n1175), .ZN(n984) );
INV_X1 U852 ( .A(n1176), .ZN(n1012) );
NAND3_X1 U853 ( .A1(n1175), .A2(n1177), .A3(n1178), .ZN(n1168) );
INV_X1 U854 ( .A(n1002), .ZN(n1178) );
NAND2_X1 U855 ( .A1(n1003), .A2(n1009), .ZN(n1177) );
INV_X1 U856 ( .A(n1179), .ZN(n1175) );
NOR2_X1 U857 ( .A1(n991), .A2(G952), .ZN(n1088) );
XOR2_X1 U858 ( .A(n1180), .B(n1181), .Z(G48) );
NOR2_X1 U859 ( .A1(KEYINPUT52), .A2(n1182), .ZN(n1181) );
NOR2_X1 U860 ( .A1(n1146), .A2(n1166), .ZN(n1180) );
XNOR2_X1 U861 ( .A(G143), .B(n1183), .ZN(G45) );
NAND2_X1 U862 ( .A1(KEYINPUT26), .A2(n1184), .ZN(n1183) );
INV_X1 U863 ( .A(n1154), .ZN(n1184) );
NAND3_X1 U864 ( .A1(n1029), .A2(n1185), .A3(n1186), .ZN(n1154) );
NOR3_X1 U865 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
XOR2_X1 U866 ( .A(n1190), .B(n1162), .Z(G42) );
NAND3_X1 U867 ( .A1(n1167), .A2(n1013), .A3(n1191), .ZN(n1162) );
XOR2_X1 U868 ( .A(G137), .B(n1157), .Z(G39) );
AND2_X1 U869 ( .A1(n1192), .A2(n1167), .ZN(n1157) );
XNOR2_X1 U870 ( .A(G134), .B(n1193), .ZN(G36) );
NAND3_X1 U871 ( .A1(n1150), .A2(n1194), .A3(n1195), .ZN(n1193) );
XOR2_X1 U872 ( .A(n997), .B(KEYINPUT30), .Z(n1195) );
XOR2_X1 U873 ( .A(G131), .B(n1156), .Z(G33) );
AND3_X1 U874 ( .A1(n1167), .A2(n1013), .A3(n1185), .ZN(n1156) );
NOR2_X1 U875 ( .A1(n997), .A2(n1187), .ZN(n1167) );
INV_X1 U876 ( .A(n1194), .ZN(n1187) );
NAND2_X1 U877 ( .A1(n1028), .A2(n1196), .ZN(n997) );
XOR2_X1 U878 ( .A(n1197), .B(n1198), .Z(G30) );
NOR2_X1 U879 ( .A1(KEYINPUT2), .A2(n1199), .ZN(n1198) );
NOR2_X1 U880 ( .A1(n1176), .A2(n1166), .ZN(n1197) );
NAND4_X1 U881 ( .A1(n1029), .A2(n1194), .A3(n1200), .A4(n1038), .ZN(n1166) );
NOR3_X1 U882 ( .A1(n1160), .A2(n1022), .A3(n1174), .ZN(n1194) );
INV_X1 U883 ( .A(n1201), .ZN(n1022) );
XOR2_X1 U884 ( .A(G101), .B(n1202), .Z(G3) );
NOR4_X1 U885 ( .A1(KEYINPUT42), .A2(n1179), .A3(n1002), .A4(n1003), .ZN(n1202) );
XOR2_X1 U886 ( .A(G125), .B(n1203), .Z(G27) );
NOR3_X1 U887 ( .A1(n1204), .A2(n1160), .A3(n1161), .ZN(n1203) );
NAND3_X1 U888 ( .A1(n1191), .A2(n1013), .A3(n1029), .ZN(n1161) );
INV_X1 U889 ( .A(n1009), .ZN(n1191) );
AND2_X1 U890 ( .A1(n1004), .A2(n1205), .ZN(n1160) );
NAND4_X1 U891 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1207), .ZN(n1205) );
INV_X1 U892 ( .A(G900), .ZN(n1207) );
XOR2_X1 U893 ( .A(KEYINPUT25), .B(n1026), .Z(n1204) );
INV_X1 U894 ( .A(n1005), .ZN(n1026) );
XOR2_X1 U895 ( .A(n1208), .B(n1143), .Z(G24) );
NAND4_X1 U896 ( .A1(n1209), .A2(n1172), .A3(n1210), .A4(n1211), .ZN(n1143) );
INV_X1 U897 ( .A(n1011), .ZN(n1172) );
NAND2_X1 U898 ( .A1(n1212), .A2(n1213), .ZN(n1011) );
XOR2_X1 U899 ( .A(n1214), .B(n1144), .Z(G21) );
NAND2_X1 U900 ( .A1(n1209), .A2(n1192), .ZN(n1144) );
NOR3_X1 U901 ( .A1(n1213), .A2(n1212), .A3(n1002), .ZN(n1192) );
XOR2_X1 U902 ( .A(G116), .B(n1215), .Z(G18) );
AND2_X1 U903 ( .A1(n1150), .A2(n1209), .ZN(n1215) );
AND2_X1 U904 ( .A1(n1216), .A2(n1029), .ZN(n1209) );
XOR2_X1 U905 ( .A(n1107), .B(KEYINPUT12), .Z(n1029) );
INV_X1 U906 ( .A(n1170), .ZN(n1107) );
NOR2_X1 U907 ( .A1(n1003), .A2(n1176), .ZN(n1150) );
NAND2_X1 U908 ( .A1(n1188), .A2(n1210), .ZN(n1176) );
INV_X1 U909 ( .A(n1189), .ZN(n1210) );
XOR2_X1 U910 ( .A(n1217), .B(n1218), .Z(G15) );
XOR2_X1 U911 ( .A(KEYINPUT51), .B(G113), .Z(n1218) );
NOR2_X1 U912 ( .A1(n1145), .A2(n1219), .ZN(n1217) );
XOR2_X1 U913 ( .A(KEYINPUT6), .B(n1013), .Z(n1219) );
INV_X1 U914 ( .A(n1146), .ZN(n1013) );
NAND2_X1 U915 ( .A1(n1189), .A2(n1220), .ZN(n1146) );
XOR2_X1 U916 ( .A(KEYINPUT20), .B(n1211), .Z(n1220) );
INV_X1 U917 ( .A(n1188), .ZN(n1211) );
NAND3_X1 U918 ( .A1(n1185), .A2(n1170), .A3(n1216), .ZN(n1145) );
NOR2_X1 U919 ( .A1(n1005), .A2(n1151), .ZN(n1216) );
INV_X1 U920 ( .A(n1221), .ZN(n1151) );
NAND2_X1 U921 ( .A1(n1174), .A2(n1201), .ZN(n1005) );
INV_X1 U922 ( .A(n1023), .ZN(n1174) );
INV_X1 U923 ( .A(n1003), .ZN(n1185) );
NAND2_X1 U924 ( .A1(n1212), .A2(n1200), .ZN(n1003) );
XOR2_X1 U925 ( .A(G110), .B(n1222), .Z(G12) );
NOR4_X1 U926 ( .A1(KEYINPUT41), .A2(n1179), .A3(n1002), .A4(n1009), .ZN(n1222) );
NAND2_X1 U927 ( .A1(n1213), .A2(n1038), .ZN(n1009) );
INV_X1 U928 ( .A(n1212), .ZN(n1038) );
XNOR2_X1 U929 ( .A(n1223), .B(n1092), .ZN(n1212) );
NAND2_X1 U930 ( .A1(G217), .A2(n1224), .ZN(n1092) );
OR2_X1 U931 ( .A1(n1091), .A2(G902), .ZN(n1223) );
XNOR2_X1 U932 ( .A(n1225), .B(n1226), .ZN(n1091) );
XOR2_X1 U933 ( .A(G110), .B(n1227), .Z(n1226) );
XOR2_X1 U934 ( .A(G146), .B(G119), .Z(n1227) );
XOR2_X1 U935 ( .A(n1228), .B(n1229), .Z(n1225) );
XOR2_X1 U936 ( .A(n1230), .B(n1063), .Z(n1228) );
NAND2_X1 U937 ( .A1(n1231), .A2(G221), .ZN(n1230) );
INV_X1 U938 ( .A(n1200), .ZN(n1213) );
XOR2_X1 U939 ( .A(n1043), .B(G472), .Z(n1200) );
AND2_X1 U940 ( .A1(n1232), .A2(n1101), .ZN(n1043) );
XOR2_X1 U941 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U942 ( .A(n1235), .B(n1236), .Z(n1233) );
INV_X1 U943 ( .A(n1112), .ZN(n1236) );
XNOR2_X1 U944 ( .A(n1237), .B(n1238), .ZN(n1112) );
XOR2_X1 U945 ( .A(n1239), .B(n1135), .Z(n1238) );
XNOR2_X1 U946 ( .A(n1240), .B(n1061), .ZN(n1135) );
XOR2_X1 U947 ( .A(G131), .B(n1229), .Z(n1061) );
XNOR2_X1 U948 ( .A(G137), .B(n1199), .ZN(n1229) );
NOR2_X1 U949 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
INV_X1 U950 ( .A(G210), .ZN(n1241) );
NAND2_X1 U951 ( .A1(KEYINPUT37), .A2(n1120), .ZN(n1235) );
XOR2_X1 U952 ( .A(n1243), .B(n1087), .Z(n1120) );
XOR2_X1 U953 ( .A(n1244), .B(G119), .Z(n1243) );
NAND2_X1 U954 ( .A1(n1189), .A2(n1188), .ZN(n1002) );
XOR2_X1 U955 ( .A(n1245), .B(G475), .Z(n1188) );
NAND2_X1 U956 ( .A1(n1103), .A2(n1101), .ZN(n1245) );
XNOR2_X1 U957 ( .A(n1246), .B(n1247), .ZN(n1103) );
XOR2_X1 U958 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U959 ( .A(G104), .B(n1250), .ZN(n1249) );
NOR3_X1 U960 ( .A1(n1242), .A2(KEYINPUT39), .A3(n1251), .ZN(n1250) );
INV_X1 U961 ( .A(G214), .ZN(n1251) );
NAND2_X1 U962 ( .A1(n991), .A2(n1252), .ZN(n1242) );
NAND2_X1 U963 ( .A1(n1253), .A2(n1254), .ZN(n1248) );
NAND2_X1 U964 ( .A1(G146), .A2(n1255), .ZN(n1254) );
NAND2_X1 U965 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XNOR2_X1 U966 ( .A(KEYINPUT53), .B(n1258), .ZN(n1256) );
NAND2_X1 U967 ( .A1(n1259), .A2(n1182), .ZN(n1253) );
NAND2_X1 U968 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
OR2_X1 U969 ( .A1(n1258), .A2(KEYINPUT53), .ZN(n1261) );
NAND2_X1 U970 ( .A1(n1063), .A2(KEYINPUT53), .ZN(n1260) );
AND2_X1 U971 ( .A1(n1257), .A2(n1258), .ZN(n1063) );
OR2_X1 U972 ( .A1(n1190), .A2(G125), .ZN(n1258) );
NAND2_X1 U973 ( .A1(G125), .A2(n1190), .ZN(n1257) );
INV_X1 U974 ( .A(G140), .ZN(n1190) );
XOR2_X1 U975 ( .A(n1262), .B(n1263), .Z(n1246) );
XOR2_X1 U976 ( .A(G143), .B(G131), .Z(n1263) );
XOR2_X1 U977 ( .A(n1244), .B(G122), .Z(n1262) );
XOR2_X1 U978 ( .A(n1264), .B(G478), .Z(n1189) );
NAND2_X1 U979 ( .A1(n1096), .A2(n1101), .ZN(n1264) );
XOR2_X1 U980 ( .A(n1265), .B(n1266), .Z(n1096) );
XOR2_X1 U981 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U982 ( .A(G134), .B(G107), .Z(n1268) );
AND3_X1 U983 ( .A1(G217), .A2(n1269), .A3(n1231), .ZN(n1267) );
AND2_X1 U984 ( .A1(G234), .A2(n991), .ZN(n1231) );
INV_X1 U985 ( .A(KEYINPUT14), .ZN(n1269) );
XNOR2_X1 U986 ( .A(n1270), .B(n1271), .ZN(n1265) );
NOR2_X1 U987 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NOR2_X1 U988 ( .A1(n1199), .A2(n1274), .ZN(n1273) );
XOR2_X1 U989 ( .A(KEYINPUT18), .B(G143), .Z(n1274) );
NOR2_X1 U990 ( .A1(G128), .A2(n1275), .ZN(n1272) );
XOR2_X1 U991 ( .A(KEYINPUT23), .B(G143), .Z(n1275) );
NAND4_X1 U992 ( .A1(n1023), .A2(n1170), .A3(n1201), .A4(n1221), .ZN(n1179) );
NAND2_X1 U993 ( .A1(n1276), .A2(n1004), .ZN(n1221) );
NAND3_X1 U994 ( .A1(n1206), .A2(n991), .A3(G952), .ZN(n1004) );
NAND4_X1 U995 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1072), .ZN(n1276) );
INV_X1 U996 ( .A(G898), .ZN(n1072) );
NAND2_X1 U997 ( .A1(G237), .A2(n1277), .ZN(n1206) );
NAND2_X1 U998 ( .A1(G221), .A2(n1224), .ZN(n1201) );
NAND2_X1 U999 ( .A1(n1277), .A2(n1101), .ZN(n1224) );
XOR2_X1 U1000 ( .A(G234), .B(KEYINPUT29), .Z(n1277) );
NOR2_X1 U1001 ( .A1(n1028), .A2(n1027), .ZN(n1170) );
INV_X1 U1002 ( .A(n1196), .ZN(n1027) );
NAND2_X1 U1003 ( .A1(G214), .A2(n1278), .ZN(n1196) );
XOR2_X1 U1004 ( .A(n1037), .B(KEYINPUT45), .Z(n1028) );
XOR2_X1 U1005 ( .A(n1279), .B(n1139), .Z(n1037) );
NAND2_X1 U1006 ( .A1(G210), .A2(n1278), .ZN(n1139) );
NAND2_X1 U1007 ( .A1(n1280), .A2(n1252), .ZN(n1278) );
INV_X1 U1008 ( .A(G237), .ZN(n1252) );
XOR2_X1 U1009 ( .A(KEYINPUT34), .B(G902), .Z(n1280) );
NAND2_X1 U1010 ( .A1(n1137), .A2(n1101), .ZN(n1279) );
XNOR2_X1 U1011 ( .A(n1281), .B(n1282), .ZN(n1137) );
XOR2_X1 U1012 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U1013 ( .A(n1285), .B(n1237), .Z(n1284) );
NOR2_X1 U1014 ( .A1(G953), .A2(n1071), .ZN(n1285) );
INV_X1 U1015 ( .A(G224), .ZN(n1071) );
XOR2_X1 U1016 ( .A(G128), .B(G125), .Z(n1283) );
XOR2_X1 U1017 ( .A(n1086), .B(n1286), .Z(n1281) );
XOR2_X1 U1018 ( .A(n1270), .B(n1287), .Z(n1286) );
INV_X1 U1019 ( .A(n1082), .ZN(n1287) );
XOR2_X1 U1020 ( .A(n1288), .B(KEYINPUT32), .Z(n1082) );
INV_X1 U1021 ( .A(G110), .ZN(n1288) );
XNOR2_X1 U1022 ( .A(n1208), .B(n1087), .ZN(n1270) );
XOR2_X1 U1023 ( .A(G116), .B(KEYINPUT38), .Z(n1087) );
INV_X1 U1024 ( .A(G122), .ZN(n1208) );
XOR2_X1 U1025 ( .A(n1289), .B(n1290), .Z(n1086) );
XOR2_X1 U1026 ( .A(n1234), .B(n1291), .Z(n1290) );
XOR2_X1 U1027 ( .A(n1292), .B(n1293), .Z(n1289) );
NOR2_X1 U1028 ( .A1(KEYINPUT5), .A2(n1214), .ZN(n1293) );
INV_X1 U1029 ( .A(G119), .ZN(n1214) );
NAND2_X1 U1030 ( .A1(KEYINPUT3), .A2(n1244), .ZN(n1292) );
INV_X1 U1031 ( .A(G113), .ZN(n1244) );
XNOR2_X1 U1032 ( .A(n1294), .B(n1040), .ZN(n1023) );
NAND2_X1 U1033 ( .A1(n1295), .A2(n1101), .ZN(n1040) );
INV_X1 U1034 ( .A(G902), .ZN(n1101) );
XOR2_X1 U1035 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1036 ( .A(n1133), .B(n1131), .Z(n1297) );
XOR2_X1 U1037 ( .A(n1298), .B(n1299), .Z(n1131) );
XOR2_X1 U1038 ( .A(G140), .B(G110), .Z(n1299) );
NAND2_X1 U1039 ( .A1(G227), .A2(n991), .ZN(n1298) );
INV_X1 U1040 ( .A(G953), .ZN(n991) );
XOR2_X1 U1041 ( .A(n1300), .B(n1062), .Z(n1133) );
AND2_X1 U1042 ( .A1(n1301), .A2(n1302), .ZN(n1062) );
OR2_X1 U1043 ( .A1(n1237), .A2(KEYINPUT21), .ZN(n1302) );
XOR2_X1 U1044 ( .A(G143), .B(G146), .Z(n1237) );
NAND3_X1 U1045 ( .A1(G143), .A2(n1182), .A3(KEYINPUT21), .ZN(n1301) );
INV_X1 U1046 ( .A(G146), .ZN(n1182) );
XNOR2_X1 U1047 ( .A(n1291), .B(n1303), .ZN(n1300) );
NOR2_X1 U1048 ( .A1(KEYINPUT50), .A2(n1234), .ZN(n1303) );
INV_X1 U1049 ( .A(n1118), .ZN(n1234) );
XNOR2_X1 U1050 ( .A(G101), .B(KEYINPUT55), .ZN(n1118) );
XOR2_X1 U1051 ( .A(G104), .B(G107), .Z(n1291) );
XOR2_X1 U1052 ( .A(n1304), .B(n1305), .Z(n1296) );
XOR2_X1 U1053 ( .A(n1199), .B(KEYINPUT48), .Z(n1305) );
INV_X1 U1054 ( .A(G128), .ZN(n1199) );
NAND2_X1 U1055 ( .A1(n1306), .A2(KEYINPUT36), .ZN(n1304) );
XOR2_X1 U1056 ( .A(n1240), .B(n1307), .Z(n1306) );
XOR2_X1 U1057 ( .A(G137), .B(G131), .Z(n1307) );
XNOR2_X1 U1058 ( .A(KEYINPUT62), .B(n1308), .ZN(n1240) );
NOR2_X1 U1059 ( .A1(KEYINPUT43), .A2(n1065), .ZN(n1308) );
XOR2_X1 U1060 ( .A(G134), .B(KEYINPUT46), .Z(n1065) );
NAND2_X1 U1061 ( .A1(KEYINPUT19), .A2(n1124), .ZN(n1294) );
INV_X1 U1062 ( .A(G469), .ZN(n1124) );
endmodule


