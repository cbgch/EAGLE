//Key = 0011110001110000111010110100001000111111111110101101100101110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351;

XOR2_X1 U744 ( .A(n1022), .B(n1023), .Z(G9) );
NAND2_X1 U745 ( .A1(KEYINPUT44), .A2(n1024), .ZN(n1023) );
XNOR2_X1 U746 ( .A(KEYINPUT26), .B(n1025), .ZN(n1024) );
NAND2_X1 U747 ( .A1(n1026), .A2(n1027), .ZN(n1022) );
XNOR2_X1 U748 ( .A(KEYINPUT15), .B(n1028), .ZN(n1027) );
NOR2_X1 U749 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U750 ( .A1(G953), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1030) );
NOR2_X1 U751 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR3_X1 U752 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1034) );
NOR2_X1 U753 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U754 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U755 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U758 ( .A1(n1049), .A2(n1026), .ZN(n1047) );
NOR2_X1 U759 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U760 ( .A1(n1052), .A2(n1053), .ZN(n1045) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR4_X1 U763 ( .A1(KEYINPUT38), .A2(n1058), .A3(n1059), .A4(n1048), .ZN(n1041) );
NOR3_X1 U764 ( .A1(n1053), .A2(n1060), .A3(n1048), .ZN(n1037) );
NOR2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1063), .A2(n1044), .ZN(n1062) );
NOR2_X1 U767 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND3_X1 U768 ( .A1(KEYINPUT38), .A2(n1066), .A3(n1067), .ZN(n1061) );
NOR4_X1 U769 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1036) );
NOR2_X1 U770 ( .A1(KEYINPUT56), .A2(n1072), .ZN(n1071) );
NOR2_X1 U771 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
AND2_X1 U772 ( .A1(n1044), .A2(KEYINPUT56), .ZN(n1070) );
XNOR2_X1 U773 ( .A(KEYINPUT55), .B(n1048), .ZN(n1069) );
INV_X1 U774 ( .A(n1075), .ZN(n1048) );
NAND2_X1 U775 ( .A1(n1067), .A2(n1058), .ZN(n1068) );
NOR3_X1 U776 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1029) );
AND4_X1 U777 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1031) );
AND4_X1 U778 ( .A1(n1080), .A2(n1081), .A3(n1058), .A4(n1056), .ZN(n1079) );
XOR2_X1 U779 ( .A(n1082), .B(KEYINPUT45), .Z(n1078) );
XNOR2_X1 U780 ( .A(n1083), .B(KEYINPUT58), .ZN(n1076) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(G72) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NAND2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1084) );
NAND3_X1 U785 ( .A1(n1092), .A2(n1087), .A3(n1093), .ZN(n1091) );
INV_X1 U786 ( .A(n1094), .ZN(n1093) );
NAND3_X1 U787 ( .A1(n1095), .A2(n1096), .A3(n1094), .ZN(n1090) );
XOR2_X1 U788 ( .A(n1097), .B(n1098), .Z(n1094) );
NOR2_X1 U789 ( .A1(KEYINPUT50), .A2(n1099), .ZN(n1098) );
XOR2_X1 U790 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U791 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U792 ( .A1(KEYINPUT28), .A2(n1104), .ZN(n1103) );
XNOR2_X1 U793 ( .A(G134), .B(G137), .ZN(n1100) );
NAND2_X1 U794 ( .A1(G953), .A2(n1089), .ZN(n1096) );
XOR2_X1 U795 ( .A(n1092), .B(KEYINPUT25), .Z(n1095) );
XOR2_X1 U796 ( .A(n1105), .B(n1106), .Z(G69) );
XOR2_X1 U797 ( .A(n1107), .B(n1108), .Z(n1106) );
AND2_X1 U798 ( .A1(n1087), .A2(n1109), .ZN(n1108) );
NOR2_X1 U799 ( .A1(KEYINPUT0), .A2(n1110), .ZN(n1107) );
NOR2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XNOR2_X1 U801 ( .A(n1113), .B(KEYINPUT51), .ZN(n1112) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(n1111) );
XNOR2_X1 U803 ( .A(n1116), .B(KEYINPUT20), .ZN(n1114) );
NAND3_X1 U804 ( .A1(G953), .A2(n1117), .A3(KEYINPUT22), .ZN(n1105) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1117) );
NOR2_X1 U806 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U807 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U808 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1118), .A2(n1124), .ZN(G63) );
XOR2_X1 U810 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR3_X1 U811 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1125) );
XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n1033), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n1118), .A2(n1130), .ZN(G60) );
XOR2_X1 U814 ( .A(n1131), .B(n1132), .Z(n1130) );
NAND3_X1 U815 ( .A1(G475), .A2(n1133), .A3(G902), .ZN(n1131) );
XNOR2_X1 U816 ( .A(KEYINPUT23), .B(n1033), .ZN(n1133) );
INV_X1 U817 ( .A(n1134), .ZN(n1033) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(G6) );
NAND2_X1 U819 ( .A1(KEYINPUT16), .A2(G104), .ZN(n1136) );
NAND3_X1 U820 ( .A1(n1137), .A2(n1138), .A3(n1065), .ZN(n1135) );
XNOR2_X1 U821 ( .A(KEYINPUT29), .B(n1139), .ZN(n1138) );
NOR2_X1 U822 ( .A1(n1118), .A2(n1140), .ZN(G57) );
XOR2_X1 U823 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U825 ( .A1(n1122), .A2(G472), .ZN(n1143) );
XNOR2_X1 U826 ( .A(n1145), .B(n1146), .ZN(n1141) );
NOR2_X1 U827 ( .A1(KEYINPUT13), .A2(G101), .ZN(n1146) );
NOR2_X1 U828 ( .A1(KEYINPUT54), .A2(n1147), .ZN(n1145) );
XOR2_X1 U829 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U830 ( .A1(KEYINPUT49), .A2(n1150), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1151), .A2(n1152), .ZN(G54) );
XOR2_X1 U832 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U834 ( .A(n1157), .B(n1158), .ZN(n1156) );
XNOR2_X1 U835 ( .A(KEYINPUT60), .B(n1159), .ZN(n1155) );
XOR2_X1 U836 ( .A(n1160), .B(n1161), .Z(n1153) );
NOR2_X1 U837 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
AND3_X1 U838 ( .A1(KEYINPUT31), .A2(n1102), .A3(n1164), .ZN(n1163) );
NOR2_X1 U839 ( .A1(KEYINPUT31), .A2(n1165), .ZN(n1162) );
XNOR2_X1 U840 ( .A(n1166), .B(n1167), .ZN(n1160) );
NAND2_X1 U841 ( .A1(n1122), .A2(G469), .ZN(n1166) );
XNOR2_X1 U842 ( .A(n1118), .B(KEYINPUT9), .ZN(n1151) );
NOR2_X1 U843 ( .A1(n1118), .A2(n1168), .ZN(G51) );
XOR2_X1 U844 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U845 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U846 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U847 ( .A(n1175), .B(KEYINPUT48), .Z(n1174) );
NAND2_X1 U848 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U849 ( .A(n1178), .B(KEYINPUT21), .Z(n1176) );
NOR2_X1 U850 ( .A1(n1178), .A2(n1177), .ZN(n1173) );
XNOR2_X1 U851 ( .A(n1179), .B(n1180), .ZN(n1177) );
NAND2_X1 U852 ( .A1(n1122), .A2(n1181), .ZN(n1171) );
NOR2_X1 U853 ( .A1(n1129), .A2(n1134), .ZN(n1122) );
NOR2_X1 U854 ( .A1(n1092), .A2(n1109), .ZN(n1134) );
NAND4_X1 U855 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1109) );
AND3_X1 U856 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
NAND2_X1 U857 ( .A1(n1026), .A2(n1189), .ZN(n1184) );
NAND3_X1 U858 ( .A1(n1190), .A2(n1028), .A3(n1191), .ZN(n1189) );
XOR2_X1 U859 ( .A(n1192), .B(KEYINPUT6), .Z(n1191) );
NAND2_X1 U860 ( .A1(n1064), .A2(n1137), .ZN(n1028) );
NAND2_X1 U861 ( .A1(n1065), .A2(n1137), .ZN(n1190) );
AND3_X1 U862 ( .A1(n1066), .A2(n1193), .A3(n1075), .ZN(n1137) );
NAND4_X1 U863 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1092) );
NOR4_X1 U864 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
INV_X1 U865 ( .A(n1202), .ZN(n1199) );
OR2_X1 U866 ( .A1(n1203), .A2(n1139), .ZN(n1196) );
NAND4_X1 U867 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1194) );
NAND2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U869 ( .A1(n1057), .A2(n1040), .ZN(n1206) );
NOR2_X1 U870 ( .A1(n1087), .A2(G952), .ZN(n1118) );
XNOR2_X1 U871 ( .A(n1210), .B(n1201), .ZN(G48) );
AND2_X1 U872 ( .A1(n1065), .A2(n1211), .ZN(n1201) );
XOR2_X1 U873 ( .A(n1212), .B(n1213), .Z(G45) );
NOR2_X1 U874 ( .A1(KEYINPUT53), .A2(n1214), .ZN(n1213) );
NOR2_X1 U875 ( .A1(n1203), .A2(n1215), .ZN(n1212) );
XNOR2_X1 U876 ( .A(KEYINPUT39), .B(n1139), .ZN(n1215) );
NAND3_X1 U877 ( .A1(n1055), .A2(n1066), .A3(n1216), .ZN(n1203) );
NOR3_X1 U878 ( .A1(n1083), .A2(n1217), .A3(n1081), .ZN(n1216) );
XOR2_X1 U879 ( .A(n1218), .B(n1219), .Z(G42) );
NOR2_X1 U880 ( .A1(KEYINPUT24), .A2(n1220), .ZN(n1219) );
AND2_X1 U881 ( .A1(n1204), .A2(n1221), .ZN(n1220) );
XNOR2_X1 U882 ( .A(G140), .B(KEYINPUT63), .ZN(n1218) );
XNOR2_X1 U883 ( .A(G137), .B(n1222), .ZN(G39) );
NAND4_X1 U884 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1058), .ZN(n1222) );
INV_X1 U885 ( .A(n1053), .ZN(n1058) );
NOR2_X1 U886 ( .A1(n1208), .A2(n1217), .ZN(n1225) );
XNOR2_X1 U887 ( .A(n1066), .B(KEYINPUT43), .ZN(n1223) );
XOR2_X1 U888 ( .A(G134), .B(n1200), .Z(G36) );
AND3_X1 U889 ( .A1(n1204), .A2(n1064), .A3(n1055), .ZN(n1200) );
XNOR2_X1 U890 ( .A(G131), .B(n1202), .ZN(G33) );
NAND3_X1 U891 ( .A1(n1055), .A2(n1204), .A3(n1065), .ZN(n1202) );
NOR3_X1 U892 ( .A1(n1059), .A2(n1217), .A3(n1053), .ZN(n1204) );
NAND2_X1 U893 ( .A1(n1226), .A2(n1051), .ZN(n1053) );
INV_X1 U894 ( .A(n1050), .ZN(n1226) );
INV_X1 U895 ( .A(n1227), .ZN(n1217) );
XNOR2_X1 U896 ( .A(n1228), .B(n1198), .ZN(G30) );
AND2_X1 U897 ( .A1(n1211), .A2(n1064), .ZN(n1198) );
AND4_X1 U898 ( .A1(n1227), .A2(n1057), .A3(n1205), .A4(n1229), .ZN(n1211) );
NOR2_X1 U899 ( .A1(n1059), .A2(n1139), .ZN(n1229) );
XNOR2_X1 U900 ( .A(G101), .B(n1230), .ZN(G3) );
NOR2_X1 U901 ( .A1(n1231), .A2(KEYINPUT14), .ZN(n1230) );
INV_X1 U902 ( .A(n1182), .ZN(n1231) );
NAND3_X1 U903 ( .A1(n1067), .A2(n1066), .A3(n1232), .ZN(n1182) );
INV_X1 U904 ( .A(n1040), .ZN(n1067) );
XNOR2_X1 U905 ( .A(G125), .B(n1195), .ZN(G27) );
NAND4_X1 U906 ( .A1(n1221), .A2(n1077), .A3(n1026), .A4(n1227), .ZN(n1195) );
NAND2_X1 U907 ( .A1(n1035), .A2(n1233), .ZN(n1227) );
NAND4_X1 U908 ( .A1(G902), .A2(G953), .A3(n1234), .A4(n1089), .ZN(n1233) );
INV_X1 U909 ( .A(G900), .ZN(n1089) );
NOR3_X1 U910 ( .A1(n1057), .A2(n1056), .A3(n1209), .ZN(n1221) );
XNOR2_X1 U911 ( .A(G122), .B(n1183), .ZN(G24) );
NAND4_X1 U912 ( .A1(n1235), .A2(n1077), .A3(n1236), .A4(n1075), .ZN(n1183) );
NOR2_X1 U913 ( .A1(n1057), .A2(n1205), .ZN(n1075) );
NOR2_X1 U914 ( .A1(n1081), .A2(n1083), .ZN(n1236) );
XOR2_X1 U915 ( .A(G119), .B(n1237), .Z(G21) );
NOR2_X1 U916 ( .A1(n1139), .A2(n1192), .ZN(n1237) );
NAND4_X1 U917 ( .A1(n1224), .A2(n1077), .A3(n1057), .A4(n1193), .ZN(n1192) );
XOR2_X1 U918 ( .A(G116), .B(n1238), .Z(G18) );
NOR2_X1 U919 ( .A1(KEYINPUT27), .A2(n1186), .ZN(n1238) );
NAND3_X1 U920 ( .A1(n1077), .A2(n1064), .A3(n1232), .ZN(n1186) );
NOR2_X1 U921 ( .A1(n1239), .A2(n1083), .ZN(n1064) );
XNOR2_X1 U922 ( .A(G113), .B(n1188), .ZN(G15) );
NAND3_X1 U923 ( .A1(n1065), .A2(n1077), .A3(n1232), .ZN(n1188) );
AND2_X1 U924 ( .A1(n1235), .A2(n1055), .ZN(n1232) );
NOR2_X1 U925 ( .A1(n1205), .A2(n1208), .ZN(n1055) );
INV_X1 U926 ( .A(n1044), .ZN(n1077) );
NAND2_X1 U927 ( .A1(n1240), .A2(n1074), .ZN(n1044) );
INV_X1 U928 ( .A(n1073), .ZN(n1240) );
INV_X1 U929 ( .A(n1209), .ZN(n1065) );
NAND2_X1 U930 ( .A1(n1083), .A2(n1239), .ZN(n1209) );
XNOR2_X1 U931 ( .A(G110), .B(n1187), .ZN(G12) );
NAND4_X1 U932 ( .A1(n1235), .A2(n1224), .A3(n1066), .A4(n1208), .ZN(n1187) );
INV_X1 U933 ( .A(n1057), .ZN(n1208) );
NAND2_X1 U934 ( .A1(n1082), .A2(n1080), .ZN(n1057) );
NAND2_X1 U935 ( .A1(G472), .A2(n1241), .ZN(n1080) );
OR2_X1 U936 ( .A1(n1241), .A2(G472), .ZN(n1082) );
NAND2_X1 U937 ( .A1(n1242), .A2(n1129), .ZN(n1241) );
XOR2_X1 U938 ( .A(n1150), .B(n1243), .Z(n1242) );
XOR2_X1 U939 ( .A(n1149), .B(n1244), .Z(n1243) );
NOR2_X1 U940 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U941 ( .A(n1247), .B(KEYINPUT18), .Z(n1246) );
NAND2_X1 U942 ( .A1(n1144), .A2(G101), .ZN(n1247) );
NOR2_X1 U943 ( .A1(G101), .A2(n1144), .ZN(n1245) );
AND2_X1 U944 ( .A1(n1248), .A2(G210), .ZN(n1144) );
XNOR2_X1 U945 ( .A(n1249), .B(n1180), .ZN(n1149) );
NAND2_X1 U946 ( .A1(n1250), .A2(n1251), .ZN(n1150) );
NAND2_X1 U947 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U948 ( .A(KEYINPUT47), .ZN(n1253) );
NAND3_X1 U949 ( .A1(G113), .A2(n1254), .A3(KEYINPUT47), .ZN(n1250) );
INV_X1 U950 ( .A(n1059), .ZN(n1066) );
NAND2_X1 U951 ( .A1(n1073), .A2(n1074), .ZN(n1059) );
NAND2_X1 U952 ( .A1(G221), .A2(n1255), .ZN(n1074) );
XNOR2_X1 U953 ( .A(n1256), .B(G469), .ZN(n1073) );
NAND2_X1 U954 ( .A1(n1257), .A2(n1129), .ZN(n1256) );
XNOR2_X1 U955 ( .A(n1167), .B(n1258), .ZN(n1257) );
XNOR2_X1 U956 ( .A(n1259), .B(n1165), .ZN(n1258) );
XNOR2_X1 U957 ( .A(n1102), .B(n1164), .ZN(n1165) );
XOR2_X1 U958 ( .A(n1260), .B(n1261), .Z(n1164) );
INV_X1 U959 ( .A(G101), .ZN(n1261) );
NAND3_X1 U960 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1260) );
OR2_X1 U961 ( .A1(n1265), .A2(n1025), .ZN(n1264) );
NAND2_X1 U962 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
INV_X1 U963 ( .A(KEYINPUT35), .ZN(n1267) );
NAND2_X1 U964 ( .A1(n1268), .A2(n1265), .ZN(n1266) );
XNOR2_X1 U965 ( .A(KEYINPUT46), .B(n1025), .ZN(n1268) );
NAND2_X1 U966 ( .A1(KEYINPUT35), .A2(n1269), .ZN(n1262) );
NAND2_X1 U967 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND3_X1 U968 ( .A1(KEYINPUT46), .A2(n1265), .A3(n1025), .ZN(n1271) );
OR2_X1 U969 ( .A1(n1025), .A2(KEYINPUT46), .ZN(n1270) );
NAND2_X1 U970 ( .A1(n1272), .A2(n1273), .ZN(n1102) );
NAND2_X1 U971 ( .A1(G128), .A2(n1274), .ZN(n1273) );
NAND3_X1 U972 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1274) );
NAND2_X1 U973 ( .A1(G146), .A2(n1278), .ZN(n1276) );
NAND2_X1 U974 ( .A1(n1279), .A2(n1210), .ZN(n1275) );
NAND2_X1 U975 ( .A1(n1280), .A2(n1228), .ZN(n1272) );
XNOR2_X1 U976 ( .A(n1279), .B(G146), .ZN(n1280) );
NOR2_X1 U977 ( .A1(n1278), .A2(n1214), .ZN(n1279) );
INV_X1 U978 ( .A(KEYINPUT11), .ZN(n1278) );
NAND3_X1 U979 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1259) );
NAND2_X1 U980 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U981 ( .A1(n1158), .A2(n1286), .ZN(n1285) );
XNOR2_X1 U982 ( .A(G140), .B(n1287), .ZN(n1284) );
OR2_X1 U983 ( .A1(n1158), .A2(KEYINPUT17), .ZN(n1282) );
NAND4_X1 U984 ( .A1(n1288), .A2(n1286), .A3(n1158), .A4(KEYINPUT17), .ZN(n1281) );
NOR2_X1 U985 ( .A1(n1088), .A2(G953), .ZN(n1158) );
INV_X1 U986 ( .A(G227), .ZN(n1088) );
INV_X1 U987 ( .A(KEYINPUT12), .ZN(n1286) );
XNOR2_X1 U988 ( .A(n1287), .B(n1159), .ZN(n1288) );
INV_X1 U989 ( .A(G140), .ZN(n1159) );
NAND2_X1 U990 ( .A1(KEYINPUT59), .A2(n1157), .ZN(n1287) );
INV_X1 U991 ( .A(G110), .ZN(n1157) );
INV_X1 U992 ( .A(n1249), .ZN(n1167) );
XNOR2_X1 U993 ( .A(n1289), .B(n1290), .ZN(n1249) );
XNOR2_X1 U994 ( .A(G134), .B(n1104), .ZN(n1290) );
NAND2_X1 U995 ( .A1(KEYINPUT36), .A2(n1291), .ZN(n1289) );
INV_X1 U996 ( .A(G137), .ZN(n1291) );
NOR2_X1 U997 ( .A1(n1040), .A2(n1056), .ZN(n1224) );
INV_X1 U998 ( .A(n1205), .ZN(n1056) );
XNOR2_X1 U999 ( .A(n1292), .B(n1123), .ZN(n1205) );
AND2_X1 U1000 ( .A1(G217), .A2(n1255), .ZN(n1123) );
NAND2_X1 U1001 ( .A1(G234), .A2(n1129), .ZN(n1255) );
NAND2_X1 U1002 ( .A1(n1121), .A2(n1129), .ZN(n1292) );
XNOR2_X1 U1003 ( .A(n1293), .B(n1294), .ZN(n1121) );
XOR2_X1 U1004 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1005 ( .A(n1297), .B(n1298), .ZN(n1296) );
NAND2_X1 U1006 ( .A1(n1299), .A2(KEYINPUT41), .ZN(n1298) );
XNOR2_X1 U1007 ( .A(G110), .B(n1300), .ZN(n1299) );
XNOR2_X1 U1008 ( .A(n1228), .B(G119), .ZN(n1300) );
NAND2_X1 U1009 ( .A1(KEYINPUT10), .A2(n1097), .ZN(n1297) );
NAND2_X1 U1010 ( .A1(KEYINPUT57), .A2(G137), .ZN(n1295) );
XOR2_X1 U1011 ( .A(n1301), .B(n1302), .Z(n1293) );
XNOR2_X1 U1012 ( .A(KEYINPUT4), .B(n1210), .ZN(n1302) );
NAND3_X1 U1013 ( .A1(G234), .A2(n1087), .A3(G221), .ZN(n1301) );
NAND2_X1 U1014 ( .A1(n1081), .A2(n1083), .ZN(n1040) );
XNOR2_X1 U1015 ( .A(n1303), .B(n1304), .ZN(n1083) );
XNOR2_X1 U1016 ( .A(KEYINPUT5), .B(n1128), .ZN(n1304) );
INV_X1 U1017 ( .A(G478), .ZN(n1128) );
OR2_X1 U1018 ( .A1(n1126), .A2(G902), .ZN(n1303) );
XNOR2_X1 U1019 ( .A(n1305), .B(n1306), .ZN(n1126) );
NOR2_X1 U1020 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XOR2_X1 U1021 ( .A(n1309), .B(KEYINPUT37), .Z(n1308) );
NAND2_X1 U1022 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NOR2_X1 U1023 ( .A1(n1310), .A2(n1311), .ZN(n1307) );
XNOR2_X1 U1024 ( .A(n1025), .B(n1312), .ZN(n1311) );
XNOR2_X1 U1025 ( .A(n1313), .B(G116), .ZN(n1312) );
INV_X1 U1026 ( .A(G107), .ZN(n1025) );
XNOR2_X1 U1027 ( .A(G128), .B(n1314), .ZN(n1310) );
XNOR2_X1 U1028 ( .A(n1214), .B(G134), .ZN(n1314) );
NAND3_X1 U1029 ( .A1(G217), .A2(n1087), .A3(G234), .ZN(n1305) );
INV_X1 U1030 ( .A(n1239), .ZN(n1081) );
XNOR2_X1 U1031 ( .A(n1315), .B(G475), .ZN(n1239) );
NAND2_X1 U1032 ( .A1(n1132), .A2(n1129), .ZN(n1315) );
XNOR2_X1 U1033 ( .A(n1316), .B(n1317), .ZN(n1132) );
XOR2_X1 U1034 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1035 ( .A(n1320), .B(G104), .Z(n1319) );
NAND2_X1 U1036 ( .A1(KEYINPUT62), .A2(n1313), .ZN(n1320) );
NAND2_X1 U1037 ( .A1(n1248), .A2(G214), .ZN(n1318) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1248) );
XOR2_X1 U1039 ( .A(n1321), .B(n1097), .Z(n1316) );
XOR2_X1 U1040 ( .A(G125), .B(G140), .Z(n1097) );
NAND3_X1 U1041 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1321) );
NAND2_X1 U1042 ( .A1(n1325), .A2(n1210), .ZN(n1324) );
XNOR2_X1 U1043 ( .A(n1214), .B(n1326), .ZN(n1325) );
INV_X1 U1044 ( .A(G143), .ZN(n1214) );
NAND3_X1 U1045 ( .A1(G143), .A2(G146), .A3(n1326), .ZN(n1323) );
OR2_X1 U1046 ( .A1(n1277), .A2(n1326), .ZN(n1322) );
XNOR2_X1 U1047 ( .A(G113), .B(n1104), .ZN(n1326) );
INV_X1 U1048 ( .A(G131), .ZN(n1104) );
INV_X1 U1049 ( .A(n1327), .ZN(n1277) );
AND2_X1 U1050 ( .A1(n1026), .A2(n1193), .ZN(n1235) );
NAND2_X1 U1051 ( .A1(n1328), .A2(n1329), .ZN(n1193) );
NAND3_X1 U1052 ( .A1(G902), .A2(n1113), .A3(n1330), .ZN(n1329) );
XOR2_X1 U1053 ( .A(n1234), .B(KEYINPUT33), .Z(n1330) );
AND2_X1 U1054 ( .A1(n1331), .A2(G953), .ZN(n1113) );
XNOR2_X1 U1055 ( .A(G898), .B(KEYINPUT32), .ZN(n1331) );
XOR2_X1 U1056 ( .A(n1035), .B(KEYINPUT7), .Z(n1328) );
NAND3_X1 U1057 ( .A1(n1234), .A2(n1087), .A3(G952), .ZN(n1035) );
NAND2_X1 U1058 ( .A1(G237), .A2(G234), .ZN(n1234) );
INV_X1 U1059 ( .A(n1139), .ZN(n1026) );
NAND2_X1 U1060 ( .A1(n1050), .A2(n1051), .ZN(n1139) );
NAND2_X1 U1061 ( .A1(n1332), .A2(n1333), .ZN(n1051) );
XOR2_X1 U1062 ( .A(KEYINPUT8), .B(G214), .Z(n1332) );
XNOR2_X1 U1063 ( .A(n1334), .B(n1181), .ZN(n1050) );
AND2_X1 U1064 ( .A1(G210), .A2(n1333), .ZN(n1181) );
NAND2_X1 U1065 ( .A1(n1335), .A2(n1129), .ZN(n1333) );
INV_X1 U1066 ( .A(G237), .ZN(n1335) );
NAND2_X1 U1067 ( .A1(n1336), .A2(n1129), .ZN(n1334) );
INV_X1 U1068 ( .A(G902), .ZN(n1129) );
XOR2_X1 U1069 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1070 ( .A(n1178), .B(n1339), .ZN(n1338) );
XNOR2_X1 U1071 ( .A(n1340), .B(KEYINPUT1), .ZN(n1339) );
NAND2_X1 U1072 ( .A1(KEYINPUT52), .A2(n1341), .ZN(n1340) );
XNOR2_X1 U1073 ( .A(KEYINPUT3), .B(n1179), .ZN(n1341) );
INV_X1 U1074 ( .A(G125), .ZN(n1179) );
NAND2_X1 U1075 ( .A1(n1342), .A2(n1087), .ZN(n1178) );
INV_X1 U1076 ( .A(G953), .ZN(n1087) );
XNOR2_X1 U1077 ( .A(G224), .B(KEYINPUT40), .ZN(n1342) );
XOR2_X1 U1078 ( .A(n1169), .B(n1180), .Z(n1337) );
XNOR2_X1 U1079 ( .A(n1343), .B(n1344), .ZN(n1180) );
NOR2_X1 U1080 ( .A1(n1327), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1081 ( .A(n1346), .B(KEYINPUT30), .Z(n1345) );
NAND2_X1 U1082 ( .A1(n1347), .A2(n1210), .ZN(n1346) );
XNOR2_X1 U1083 ( .A(G143), .B(KEYINPUT34), .ZN(n1347) );
NOR2_X1 U1084 ( .A1(n1210), .A2(G143), .ZN(n1327) );
INV_X1 U1085 ( .A(G146), .ZN(n1210) );
NAND2_X1 U1086 ( .A1(KEYINPUT42), .A2(n1228), .ZN(n1343) );
INV_X1 U1087 ( .A(G128), .ZN(n1228) );
XNOR2_X1 U1088 ( .A(n1348), .B(n1349), .ZN(n1169) );
INV_X1 U1089 ( .A(n1116), .ZN(n1349) );
XOR2_X1 U1090 ( .A(n1252), .B(n1350), .Z(n1116) );
XNOR2_X1 U1091 ( .A(n1313), .B(G110), .ZN(n1350) );
INV_X1 U1092 ( .A(G122), .ZN(n1313) );
XOR2_X1 U1093 ( .A(G113), .B(n1254), .Z(n1252) );
XOR2_X1 U1094 ( .A(G116), .B(G119), .Z(n1254) );
NAND2_X1 U1095 ( .A1(KEYINPUT2), .A2(n1115), .ZN(n1348) );
XNOR2_X1 U1096 ( .A(n1351), .B(n1265), .ZN(n1115) );
XOR2_X1 U1097 ( .A(G104), .B(KEYINPUT19), .Z(n1265) );
XNOR2_X1 U1098 ( .A(G101), .B(G107), .ZN(n1351) );
endmodule


