//Key = 0101100010110101111100011110001011110110111011111100100011010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423;

XNOR2_X1 U772 ( .A(G107), .B(n1081), .ZN(G9) );
NAND4_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
OR2_X1 U775 ( .A1(n1088), .A2(KEYINPUT53), .ZN(n1083) );
NAND2_X1 U776 ( .A1(KEYINPUT53), .A2(n1089), .ZN(n1082) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U778 ( .A1(n1092), .A2(n1093), .ZN(G75) );
NOR3_X1 U779 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
NAND3_X1 U780 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1094) );
NAND2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND3_X1 U783 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
NAND2_X1 U784 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
OR3_X1 U785 ( .A1(n1087), .A2(KEYINPUT47), .A3(n1109), .ZN(n1107) );
NAND3_X1 U786 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1104) );
NAND2_X1 U787 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NAND2_X1 U788 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U789 ( .A1(KEYINPUT47), .A2(n1117), .ZN(n1116) );
NAND2_X1 U790 ( .A1(n1118), .A2(n1119), .ZN(n1110) );
NAND2_X1 U791 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U792 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND3_X1 U793 ( .A1(n1113), .A2(n1124), .A3(n1118), .ZN(n1102) );
NAND2_X1 U794 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U795 ( .A1(n1112), .A2(n1127), .ZN(n1126) );
OR2_X1 U796 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U797 ( .A1(n1106), .A2(n1130), .ZN(n1125) );
NAND2_X1 U798 ( .A1(n1090), .A2(n1131), .ZN(n1130) );
NAND2_X1 U799 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
INV_X1 U800 ( .A(n1134), .ZN(n1100) );
NOR3_X1 U801 ( .A1(n1135), .A2(G953), .A3(G952), .ZN(n1092) );
INV_X1 U802 ( .A(n1097), .ZN(n1135) );
NAND4_X1 U803 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1097) );
NOR3_X1 U804 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
XOR2_X1 U805 ( .A(KEYINPUT5), .B(n1143), .Z(n1142) );
NOR2_X1 U806 ( .A1(G478), .A2(n1144), .ZN(n1143) );
XNOR2_X1 U807 ( .A(n1145), .B(n1146), .ZN(n1141) );
NAND3_X1 U808 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1140) );
XOR2_X1 U809 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U810 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
NAND2_X1 U811 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND2_X1 U812 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
OR2_X1 U813 ( .A1(n1157), .A2(n1158), .ZN(n1154) );
INV_X1 U814 ( .A(KEYINPUT46), .ZN(n1157) );
NAND2_X1 U815 ( .A1(n1158), .A2(n1159), .ZN(n1147) );
NOR2_X1 U816 ( .A1(n1160), .A2(KEYINPUT27), .ZN(n1158) );
INV_X1 U817 ( .A(n1156), .ZN(n1160) );
NOR3_X1 U818 ( .A1(n1161), .A2(n1122), .A3(n1132), .ZN(n1138) );
AND2_X1 U819 ( .A1(n1144), .A2(G478), .ZN(n1161) );
XOR2_X1 U820 ( .A(n1162), .B(n1163), .Z(n1137) );
XNOR2_X1 U821 ( .A(n1164), .B(KEYINPUT17), .ZN(n1163) );
XOR2_X1 U822 ( .A(KEYINPUT11), .B(n1165), .Z(n1136) );
XOR2_X1 U823 ( .A(n1166), .B(n1167), .Z(G72) );
XOR2_X1 U824 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U825 ( .A1(G953), .A2(n1170), .ZN(n1169) );
NAND2_X1 U826 ( .A1(G900), .A2(G227), .ZN(n1170) );
NAND2_X1 U827 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
NAND2_X1 U828 ( .A1(G953), .A2(n1173), .ZN(n1172) );
XOR2_X1 U829 ( .A(n1174), .B(n1175), .Z(n1171) );
XOR2_X1 U830 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U831 ( .A1(n1178), .A2(n1179), .ZN(n1174) );
NAND2_X1 U832 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U833 ( .A(KEYINPUT56), .B(n1182), .Z(n1180) );
NAND2_X1 U834 ( .A1(n1182), .A2(G137), .ZN(n1178) );
AND2_X1 U835 ( .A1(n1095), .A2(n1098), .ZN(n1166) );
NAND2_X1 U836 ( .A1(n1183), .A2(n1184), .ZN(G69) );
NAND3_X1 U837 ( .A1(n1185), .A2(n1186), .A3(G953), .ZN(n1184) );
XOR2_X1 U838 ( .A(KEYINPUT33), .B(n1187), .Z(n1183) );
NOR2_X1 U839 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U840 ( .A(n1096), .B(n1186), .Z(n1189) );
NAND2_X1 U841 ( .A1(n1190), .A2(n1191), .ZN(n1186) );
NAND2_X1 U842 ( .A1(G953), .A2(n1192), .ZN(n1191) );
XOR2_X1 U843 ( .A(KEYINPUT14), .B(n1193), .Z(n1190) );
NOR2_X1 U844 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U845 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U846 ( .A(KEYINPUT59), .B(n1198), .Z(n1197) );
NOR2_X1 U847 ( .A1(n1199), .A2(n1198), .ZN(n1194) );
XNOR2_X1 U848 ( .A(n1200), .B(n1201), .ZN(n1198) );
NOR2_X1 U849 ( .A1(KEYINPUT7), .A2(n1202), .ZN(n1201) );
INV_X1 U850 ( .A(n1196), .ZN(n1199) );
AND2_X1 U851 ( .A1(n1185), .A2(G953), .ZN(n1188) );
NAND2_X1 U852 ( .A1(G898), .A2(G224), .ZN(n1185) );
NOR2_X1 U853 ( .A1(n1203), .A2(n1204), .ZN(G66) );
XOR2_X1 U854 ( .A(n1205), .B(n1206), .Z(n1204) );
NAND3_X1 U855 ( .A1(n1207), .A2(n1159), .A3(KEYINPUT32), .ZN(n1205) );
NOR2_X1 U856 ( .A1(n1203), .A2(n1208), .ZN(G63) );
XOR2_X1 U857 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U858 ( .A(KEYINPUT48), .B(n1211), .Z(n1210) );
AND2_X1 U859 ( .A1(G478), .A2(n1207), .ZN(n1211) );
NOR3_X1 U860 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(G60) );
AND2_X1 U861 ( .A1(KEYINPUT61), .A2(n1203), .ZN(n1214) );
NOR3_X1 U862 ( .A1(KEYINPUT61), .A2(G953), .A3(G952), .ZN(n1213) );
XOR2_X1 U863 ( .A(n1215), .B(n1216), .Z(n1212) );
NAND3_X1 U864 ( .A1(n1207), .A2(G475), .A3(KEYINPUT18), .ZN(n1216) );
XOR2_X1 U865 ( .A(G104), .B(n1217), .Z(G6) );
NOR2_X1 U866 ( .A1(n1203), .A2(n1218), .ZN(G57) );
XOR2_X1 U867 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U868 ( .A(G101), .B(n1221), .Z(n1220) );
NOR2_X1 U869 ( .A1(KEYINPUT60), .A2(n1222), .ZN(n1221) );
XOR2_X1 U870 ( .A(n1223), .B(KEYINPUT51), .Z(n1222) );
XNOR2_X1 U871 ( .A(n1224), .B(n1225), .ZN(n1219) );
NOR2_X1 U872 ( .A1(n1151), .A2(n1226), .ZN(n1225) );
INV_X1 U873 ( .A(G472), .ZN(n1151) );
NOR2_X1 U874 ( .A1(n1203), .A2(n1227), .ZN(G54) );
XOR2_X1 U875 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U876 ( .A(n1230), .B(n1231), .Z(n1229) );
NAND2_X1 U877 ( .A1(KEYINPUT10), .A2(n1232), .ZN(n1231) );
NAND2_X1 U878 ( .A1(n1233), .A2(n1234), .ZN(n1230) );
INV_X1 U879 ( .A(n1235), .ZN(n1234) );
XOR2_X1 U880 ( .A(KEYINPUT40), .B(n1236), .Z(n1233) );
XOR2_X1 U881 ( .A(n1237), .B(n1238), .Z(n1228) );
AND2_X1 U882 ( .A1(G469), .A2(n1207), .ZN(n1238) );
INV_X1 U883 ( .A(n1226), .ZN(n1207) );
NAND2_X1 U884 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
XNOR2_X1 U885 ( .A(KEYINPUT25), .B(n1241), .ZN(n1239) );
NOR2_X1 U886 ( .A1(n1203), .A2(n1242), .ZN(G51) );
XOR2_X1 U887 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U888 ( .A(n1245), .B(n1246), .Z(n1244) );
NOR2_X1 U889 ( .A1(n1247), .A2(KEYINPUT22), .ZN(n1245) );
XNOR2_X1 U890 ( .A(n1248), .B(n1249), .ZN(n1243) );
NOR2_X1 U891 ( .A1(n1162), .A2(n1226), .ZN(n1249) );
NAND2_X1 U892 ( .A1(G902), .A2(n1250), .ZN(n1226) );
OR2_X1 U893 ( .A1(n1096), .A2(n1095), .ZN(n1250) );
NAND4_X1 U894 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1095) );
NOR4_X1 U895 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
NOR2_X1 U896 ( .A1(KEYINPUT39), .A2(n1259), .ZN(n1258) );
NOR2_X1 U897 ( .A1(n1260), .A2(n1261), .ZN(n1257) );
NOR2_X1 U898 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
NOR2_X1 U899 ( .A1(KEYINPUT58), .A2(n1264), .ZN(n1263) );
AND4_X1 U900 ( .A1(n1117), .A2(n1112), .A3(n1265), .A4(KEYINPUT39), .ZN(n1262) );
AND4_X1 U901 ( .A1(n1120), .A2(n1129), .A3(n1266), .A4(KEYINPUT58), .ZN(n1256) );
INV_X1 U902 ( .A(n1267), .ZN(n1255) );
NOR3_X1 U903 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1253) );
NAND4_X1 U904 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1096) );
NOR4_X1 U905 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1217), .ZN(n1274) );
NOR4_X1 U906 ( .A1(n1115), .A2(n1278), .A3(n1120), .A4(n1086), .ZN(n1217) );
NAND3_X1 U907 ( .A1(n1084), .A2(n1279), .A3(n1088), .ZN(n1273) );
NAND2_X1 U908 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U909 ( .A1(n1117), .A2(n1106), .ZN(n1281) );
INV_X1 U910 ( .A(n1086), .ZN(n1106) );
NAND2_X1 U911 ( .A1(n1128), .A2(n1118), .ZN(n1280) );
NOR2_X1 U912 ( .A1(n1098), .A2(G952), .ZN(n1203) );
XOR2_X1 U913 ( .A(G146), .B(n1268), .Z(G48) );
AND3_X1 U914 ( .A1(n1282), .A2(n1283), .A3(n1284), .ZN(n1268) );
NAND2_X1 U915 ( .A1(n1285), .A2(n1286), .ZN(G45) );
NAND2_X1 U916 ( .A1(G143), .A2(n1267), .ZN(n1286) );
XOR2_X1 U917 ( .A(KEYINPUT8), .B(n1287), .Z(n1285) );
NOR2_X1 U918 ( .A1(G143), .A2(n1267), .ZN(n1287) );
NAND3_X1 U919 ( .A1(n1288), .A2(n1283), .A3(n1289), .ZN(n1267) );
NOR3_X1 U920 ( .A1(n1290), .A2(n1265), .A3(n1291), .ZN(n1289) );
XNOR2_X1 U921 ( .A(G140), .B(n1251), .ZN(G42) );
NAND3_X1 U922 ( .A1(n1128), .A2(n1084), .A3(n1266), .ZN(n1251) );
XOR2_X1 U923 ( .A(n1181), .B(n1292), .Z(G39) );
NOR2_X1 U924 ( .A1(n1270), .A2(KEYINPUT36), .ZN(n1292) );
AND3_X1 U925 ( .A1(n1284), .A2(n1118), .A3(n1112), .ZN(n1270) );
INV_X1 U926 ( .A(n1108), .ZN(n1112) );
XNOR2_X1 U927 ( .A(n1259), .B(n1293), .ZN(G36) );
NOR2_X1 U928 ( .A1(KEYINPUT31), .A2(n1294), .ZN(n1293) );
INV_X1 U929 ( .A(G134), .ZN(n1294) );
OR4_X1 U930 ( .A1(n1108), .A2(n1261), .A3(n1087), .A4(n1265), .ZN(n1259) );
XOR2_X1 U931 ( .A(n1295), .B(n1296), .Z(G33) );
NOR2_X1 U932 ( .A1(n1261), .A2(n1264), .ZN(n1296) );
INV_X1 U933 ( .A(n1266), .ZN(n1264) );
NOR3_X1 U934 ( .A1(n1115), .A2(n1265), .A3(n1108), .ZN(n1266) );
NAND2_X1 U935 ( .A1(n1297), .A2(n1133), .ZN(n1108) );
XOR2_X1 U936 ( .A(KEYINPUT57), .B(n1132), .Z(n1297) );
XNOR2_X1 U937 ( .A(G131), .B(KEYINPUT15), .ZN(n1295) );
XNOR2_X1 U938 ( .A(G128), .B(n1298), .ZN(G30) );
NOR2_X1 U939 ( .A1(n1269), .A2(KEYINPUT43), .ZN(n1298) );
AND3_X1 U940 ( .A1(n1117), .A2(n1283), .A3(n1284), .ZN(n1269) );
NOR4_X1 U941 ( .A1(n1120), .A2(n1299), .A3(n1300), .A4(n1265), .ZN(n1284) );
XNOR2_X1 U942 ( .A(n1277), .B(n1301), .ZN(G3) );
XOR2_X1 U943 ( .A(n1302), .B(KEYINPUT2), .Z(n1301) );
AND3_X1 U944 ( .A1(n1288), .A2(n1088), .A3(n1118), .ZN(n1277) );
INV_X1 U945 ( .A(n1261), .ZN(n1288) );
NAND2_X1 U946 ( .A1(n1129), .A2(n1084), .ZN(n1261) );
XNOR2_X1 U947 ( .A(G125), .B(n1252), .ZN(G27) );
NAND4_X1 U948 ( .A1(n1128), .A2(n1282), .A3(n1303), .A4(n1113), .ZN(n1252) );
NOR2_X1 U949 ( .A1(n1265), .A2(n1090), .ZN(n1303) );
INV_X1 U950 ( .A(n1283), .ZN(n1090) );
AND2_X1 U951 ( .A1(n1134), .A2(n1304), .ZN(n1265) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1173), .A4(n1305), .ZN(n1304) );
XOR2_X1 U953 ( .A(KEYINPUT3), .B(G900), .Z(n1173) );
XOR2_X1 U954 ( .A(n1306), .B(n1271), .Z(G24) );
NAND3_X1 U955 ( .A1(n1088), .A2(n1113), .A3(n1307), .ZN(n1271) );
NOR3_X1 U956 ( .A1(n1086), .A2(n1291), .A3(n1290), .ZN(n1307) );
NAND2_X1 U957 ( .A1(n1300), .A2(n1299), .ZN(n1086) );
XNOR2_X1 U958 ( .A(G119), .B(n1272), .ZN(G21) );
NAND3_X1 U959 ( .A1(n1118), .A2(n1088), .A3(n1308), .ZN(n1272) );
NOR3_X1 U960 ( .A1(n1109), .A2(n1300), .A3(n1299), .ZN(n1308) );
INV_X1 U961 ( .A(n1309), .ZN(n1299) );
XOR2_X1 U962 ( .A(G116), .B(n1276), .Z(G18) );
AND2_X1 U963 ( .A1(n1310), .A2(n1117), .ZN(n1276) );
INV_X1 U964 ( .A(n1087), .ZN(n1117) );
NAND2_X1 U965 ( .A1(n1291), .A2(n1311), .ZN(n1087) );
XOR2_X1 U966 ( .A(G113), .B(n1275), .Z(G15) );
AND2_X1 U967 ( .A1(n1282), .A2(n1310), .ZN(n1275) );
AND3_X1 U968 ( .A1(n1113), .A2(n1129), .A3(n1088), .ZN(n1310) );
NOR2_X1 U969 ( .A1(n1309), .A2(n1300), .ZN(n1129) );
INV_X1 U970 ( .A(n1109), .ZN(n1113) );
NAND2_X1 U971 ( .A1(n1123), .A2(n1312), .ZN(n1109) );
INV_X1 U972 ( .A(n1115), .ZN(n1282) );
NAND2_X1 U973 ( .A1(n1290), .A2(n1165), .ZN(n1115) );
XOR2_X1 U974 ( .A(n1313), .B(n1314), .Z(G12) );
XNOR2_X1 U975 ( .A(G110), .B(KEYINPUT9), .ZN(n1314) );
NAND4_X1 U976 ( .A1(n1315), .A2(n1128), .A3(n1118), .A4(n1088), .ZN(n1313) );
INV_X1 U977 ( .A(n1278), .ZN(n1088) );
NAND2_X1 U978 ( .A1(n1283), .A2(n1091), .ZN(n1278) );
NAND2_X1 U979 ( .A1(n1134), .A2(n1316), .ZN(n1091) );
NAND4_X1 U980 ( .A1(G953), .A2(G902), .A3(n1305), .A4(n1192), .ZN(n1316) );
INV_X1 U981 ( .A(G898), .ZN(n1192) );
NAND3_X1 U982 ( .A1(n1305), .A2(n1098), .A3(G952), .ZN(n1134) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1305) );
NOR2_X1 U984 ( .A1(n1133), .A2(n1317), .ZN(n1283) );
XNOR2_X1 U985 ( .A(KEYINPUT57), .B(n1132), .ZN(n1317) );
AND2_X1 U986 ( .A1(G214), .A2(n1318), .ZN(n1132) );
XNOR2_X1 U987 ( .A(n1162), .B(n1319), .ZN(n1133) );
NOR2_X1 U988 ( .A1(n1164), .A2(KEYINPUT50), .ZN(n1319) );
AND2_X1 U989 ( .A1(n1320), .A2(n1321), .ZN(n1164) );
XNOR2_X1 U990 ( .A(n1246), .B(n1322), .ZN(n1320) );
XNOR2_X1 U991 ( .A(n1247), .B(n1323), .ZN(n1322) );
NOR2_X1 U992 ( .A1(KEYINPUT6), .A2(n1248), .ZN(n1323) );
NAND2_X1 U993 ( .A1(G224), .A2(n1324), .ZN(n1248) );
AND2_X1 U994 ( .A1(n1325), .A2(n1326), .ZN(n1247) );
NAND2_X1 U995 ( .A1(KEYINPUT55), .A2(n1196), .ZN(n1326) );
XOR2_X1 U996 ( .A(n1327), .B(n1328), .Z(n1325) );
OR2_X1 U997 ( .A1(n1196), .A2(KEYINPUT55), .ZN(n1328) );
XOR2_X1 U998 ( .A(n1329), .B(G110), .Z(n1196) );
NAND2_X1 U999 ( .A1(KEYINPUT1), .A2(n1306), .ZN(n1329) );
NAND2_X1 U1000 ( .A1(n1330), .A2(n1331), .ZN(n1327) );
NAND2_X1 U1001 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XNOR2_X1 U1002 ( .A(KEYINPUT21), .B(n1200), .ZN(n1333) );
XNOR2_X1 U1003 ( .A(n1202), .B(KEYINPUT29), .ZN(n1332) );
XOR2_X1 U1004 ( .A(n1334), .B(KEYINPUT28), .Z(n1330) );
NAND2_X1 U1005 ( .A1(n1200), .A2(n1202), .ZN(n1334) );
XNOR2_X1 U1006 ( .A(n1335), .B(n1336), .ZN(n1202) );
XOR2_X1 U1007 ( .A(G104), .B(G101), .Z(n1336) );
NAND2_X1 U1008 ( .A1(KEYINPUT4), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1009 ( .A(n1338), .B(n1339), .Z(n1200) );
XOR2_X1 U1010 ( .A(G119), .B(G116), .Z(n1339) );
NAND2_X1 U1011 ( .A1(KEYINPUT37), .A2(G113), .ZN(n1338) );
XOR2_X1 U1012 ( .A(n1340), .B(n1341), .Z(n1246) );
XOR2_X1 U1013 ( .A(KEYINPUT38), .B(n1342), .Z(n1341) );
NAND2_X1 U1014 ( .A1(G210), .A2(n1318), .ZN(n1162) );
NAND2_X1 U1015 ( .A1(n1343), .A2(n1344), .ZN(n1318) );
NOR2_X1 U1016 ( .A1(n1311), .A2(n1165), .ZN(n1118) );
INV_X1 U1017 ( .A(n1291), .ZN(n1165) );
XOR2_X1 U1018 ( .A(n1345), .B(G475), .Z(n1291) );
NAND2_X1 U1019 ( .A1(n1321), .A2(n1215), .ZN(n1345) );
NAND3_X1 U1020 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(n1215) );
NAND2_X1 U1021 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1022 ( .A1(n1351), .A2(n1352), .ZN(n1347) );
INV_X1 U1023 ( .A(KEYINPUT42), .ZN(n1352) );
NAND2_X1 U1024 ( .A1(n1353), .A2(n1354), .ZN(n1351) );
XNOR2_X1 U1025 ( .A(KEYINPUT62), .B(n1349), .ZN(n1354) );
NAND2_X1 U1026 ( .A1(KEYINPUT42), .A2(n1355), .ZN(n1346) );
NAND2_X1 U1027 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
OR3_X1 U1028 ( .A1(n1349), .A2(n1350), .A3(KEYINPUT62), .ZN(n1357) );
INV_X1 U1029 ( .A(n1353), .ZN(n1350) );
XOR2_X1 U1030 ( .A(n1358), .B(n1359), .Z(n1353) );
XOR2_X1 U1031 ( .A(G122), .B(G113), .Z(n1359) );
NAND2_X1 U1032 ( .A1(KEYINPUT62), .A2(n1349), .ZN(n1356) );
XOR2_X1 U1033 ( .A(n1360), .B(n1361), .Z(n1349) );
XNOR2_X1 U1034 ( .A(n1362), .B(n1342), .ZN(n1361) );
XOR2_X1 U1035 ( .A(G125), .B(G146), .Z(n1342) );
NAND2_X1 U1036 ( .A1(KEYINPUT16), .A2(n1363), .ZN(n1362) );
XNOR2_X1 U1037 ( .A(G143), .B(n1364), .ZN(n1363) );
NAND2_X1 U1038 ( .A1(G214), .A2(n1365), .ZN(n1364) );
XNOR2_X1 U1039 ( .A(G131), .B(G140), .ZN(n1360) );
INV_X1 U1040 ( .A(n1290), .ZN(n1311) );
XOR2_X1 U1041 ( .A(n1144), .B(n1366), .Z(n1290) );
XOR2_X1 U1042 ( .A(KEYINPUT0), .B(G478), .Z(n1366) );
NAND2_X1 U1043 ( .A1(n1209), .A2(n1321), .ZN(n1144) );
XNOR2_X1 U1044 ( .A(n1367), .B(n1368), .ZN(n1209) );
XOR2_X1 U1045 ( .A(n1340), .B(n1337), .Z(n1368) );
XOR2_X1 U1046 ( .A(n1369), .B(n1370), .Z(n1367) );
NOR2_X1 U1047 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
INV_X1 U1048 ( .A(G217), .ZN(n1372) );
XOR2_X1 U1049 ( .A(n1373), .B(G134), .Z(n1369) );
NAND2_X1 U1050 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
OR2_X1 U1051 ( .A1(n1376), .A2(G116), .ZN(n1375) );
XOR2_X1 U1052 ( .A(n1377), .B(KEYINPUT63), .Z(n1374) );
NAND2_X1 U1053 ( .A1(G116), .A2(n1376), .ZN(n1377) );
XNOR2_X1 U1054 ( .A(n1306), .B(KEYINPUT52), .ZN(n1376) );
INV_X1 U1055 ( .A(G122), .ZN(n1306) );
AND2_X1 U1056 ( .A1(n1300), .A2(n1309), .ZN(n1128) );
XNOR2_X1 U1057 ( .A(n1156), .B(n1159), .ZN(n1309) );
INV_X1 U1058 ( .A(n1153), .ZN(n1159) );
NAND2_X1 U1059 ( .A1(G217), .A2(n1378), .ZN(n1153) );
NAND2_X1 U1060 ( .A1(n1206), .A2(n1321), .ZN(n1156) );
XNOR2_X1 U1061 ( .A(n1379), .B(n1380), .ZN(n1206) );
XOR2_X1 U1062 ( .A(G119), .B(n1381), .Z(n1380) );
XOR2_X1 U1063 ( .A(G137), .B(G128), .Z(n1381) );
XOR2_X1 U1064 ( .A(n1382), .B(n1383), .Z(n1379) );
NOR2_X1 U1065 ( .A1(n1384), .A2(n1371), .ZN(n1383) );
NAND2_X1 U1066 ( .A1(n1324), .A2(G234), .ZN(n1371) );
INV_X1 U1067 ( .A(G221), .ZN(n1384) );
XOR2_X1 U1068 ( .A(n1385), .B(G110), .Z(n1382) );
NAND3_X1 U1069 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n1385) );
NAND2_X1 U1070 ( .A1(n1177), .A2(n1389), .ZN(n1388) );
NAND2_X1 U1071 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
INV_X1 U1072 ( .A(KEYINPUT20), .ZN(n1391) );
XOR2_X1 U1073 ( .A(n1392), .B(KEYINPUT49), .Z(n1390) );
OR3_X1 U1074 ( .A1(n1392), .A2(n1177), .A3(KEYINPUT20), .ZN(n1387) );
XOR2_X1 U1075 ( .A(G125), .B(G140), .Z(n1177) );
NAND2_X1 U1076 ( .A1(KEYINPUT20), .A2(n1392), .ZN(n1386) );
XOR2_X1 U1077 ( .A(n1393), .B(KEYINPUT26), .Z(n1392) );
XOR2_X1 U1078 ( .A(n1394), .B(G472), .Z(n1300) );
NAND2_X1 U1079 ( .A1(KEYINPUT24), .A2(n1150), .ZN(n1394) );
AND2_X1 U1080 ( .A1(n1321), .A2(n1395), .ZN(n1150) );
NAND2_X1 U1081 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
NAND2_X1 U1082 ( .A1(n1398), .A2(n1224), .ZN(n1397) );
XOR2_X1 U1083 ( .A(KEYINPUT19), .B(n1399), .Z(n1396) );
NOR2_X1 U1084 ( .A1(n1224), .A2(n1398), .ZN(n1399) );
XOR2_X1 U1085 ( .A(n1223), .B(G101), .Z(n1398) );
NAND2_X1 U1086 ( .A1(G210), .A2(n1365), .ZN(n1223) );
AND2_X1 U1087 ( .A1(n1324), .A2(n1344), .ZN(n1365) );
INV_X1 U1088 ( .A(G237), .ZN(n1344) );
XNOR2_X1 U1089 ( .A(n1400), .B(n1401), .ZN(n1224) );
XOR2_X1 U1090 ( .A(G113), .B(n1402), .Z(n1401) );
XOR2_X1 U1091 ( .A(G146), .B(G119), .Z(n1402) );
XOR2_X1 U1092 ( .A(n1403), .B(n1404), .Z(n1400) );
NOR2_X1 U1093 ( .A1(n1405), .A2(n1406), .ZN(n1404) );
AND2_X1 U1094 ( .A1(KEYINPUT30), .A2(n1407), .ZN(n1406) );
NOR2_X1 U1095 ( .A1(KEYINPUT34), .A2(n1407), .ZN(n1405) );
INV_X1 U1096 ( .A(G116), .ZN(n1407) );
XOR2_X1 U1097 ( .A(n1232), .B(n1340), .Z(n1403) );
XOR2_X1 U1098 ( .A(G128), .B(G143), .Z(n1340) );
XOR2_X1 U1099 ( .A(n1120), .B(KEYINPUT41), .Z(n1315) );
INV_X1 U1100 ( .A(n1084), .ZN(n1120) );
NOR2_X1 U1101 ( .A1(n1123), .A2(n1122), .ZN(n1084) );
INV_X1 U1102 ( .A(n1312), .ZN(n1122) );
NAND2_X1 U1103 ( .A1(G221), .A2(n1378), .ZN(n1312) );
NAND2_X1 U1104 ( .A1(G234), .A2(n1343), .ZN(n1378) );
INV_X1 U1105 ( .A(G902), .ZN(n1343) );
XNOR2_X1 U1106 ( .A(n1146), .B(n1408), .ZN(n1123) );
NOR2_X1 U1107 ( .A1(n1145), .A2(KEYINPUT12), .ZN(n1408) );
AND2_X1 U1108 ( .A1(n1409), .A2(n1321), .ZN(n1145) );
XOR2_X1 U1109 ( .A(G902), .B(KEYINPUT45), .Z(n1321) );
XOR2_X1 U1110 ( .A(n1410), .B(n1411), .Z(n1409) );
INV_X1 U1111 ( .A(n1232), .ZN(n1411) );
XOR2_X1 U1112 ( .A(n1181), .B(n1182), .Z(n1232) );
XOR2_X1 U1113 ( .A(G131), .B(G134), .Z(n1182) );
INV_X1 U1114 ( .A(G137), .ZN(n1181) );
XOR2_X1 U1115 ( .A(n1412), .B(n1413), .Z(n1410) );
NOR2_X1 U1116 ( .A1(n1236), .A2(n1235), .ZN(n1413) );
NOR2_X1 U1117 ( .A1(n1414), .A2(n1415), .ZN(n1235) );
AND2_X1 U1118 ( .A1(n1415), .A2(n1414), .ZN(n1236) );
NAND2_X1 U1119 ( .A1(G227), .A2(n1324), .ZN(n1414) );
XOR2_X1 U1120 ( .A(n1098), .B(KEYINPUT54), .Z(n1324) );
INV_X1 U1121 ( .A(G953), .ZN(n1098) );
XOR2_X1 U1122 ( .A(G110), .B(G140), .Z(n1415) );
NAND2_X1 U1123 ( .A1(n1240), .A2(n1241), .ZN(n1412) );
NAND2_X1 U1124 ( .A1(n1416), .A2(n1417), .ZN(n1241) );
INV_X1 U1125 ( .A(n1176), .ZN(n1417) );
XOR2_X1 U1126 ( .A(n1418), .B(n1419), .Z(n1416) );
NAND2_X1 U1127 ( .A1(n1176), .A2(n1420), .ZN(n1240) );
XOR2_X1 U1128 ( .A(n1419), .B(n1421), .Z(n1420) );
INV_X1 U1129 ( .A(n1418), .ZN(n1421) );
XOR2_X1 U1130 ( .A(n1358), .B(n1337), .Z(n1418) );
XOR2_X1 U1131 ( .A(G107), .B(KEYINPUT35), .Z(n1337) );
INV_X1 U1132 ( .A(G104), .ZN(n1358) );
AND2_X1 U1133 ( .A1(KEYINPUT44), .A2(n1302), .ZN(n1419) );
INV_X1 U1134 ( .A(G101), .ZN(n1302) );
XOR2_X1 U1135 ( .A(n1422), .B(G128), .Z(n1176) );
NAND2_X1 U1136 ( .A1(n1423), .A2(KEYINPUT23), .ZN(n1422) );
XOR2_X1 U1137 ( .A(G143), .B(n1393), .Z(n1423) );
INV_X1 U1138 ( .A(G146), .ZN(n1393) );
XOR2_X1 U1139 ( .A(G469), .B(KEYINPUT13), .Z(n1146) );
endmodule


