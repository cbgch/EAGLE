//Key = 0110101100101010101101101011110111110111100010111010100111110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327;

XNOR2_X1 U740 ( .A(G107), .B(n1014), .ZN(G9) );
NOR2_X1 U741 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
NOR2_X1 U743 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U744 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U745 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
INV_X1 U746 ( .A(n1027), .ZN(n1026) );
NOR2_X1 U747 ( .A1(n1028), .A2(n1029), .ZN(n1025) );
AND2_X1 U748 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR3_X1 U749 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1023) );
NOR3_X1 U750 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
AND2_X1 U753 ( .A1(n1042), .A2(KEYINPUT31), .ZN(n1040) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1036) );
NOR2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1047), .A2(n1048), .ZN(n1033) );
NOR3_X1 U757 ( .A1(n1049), .A2(KEYINPUT31), .A3(n1039), .ZN(n1048) );
INV_X1 U758 ( .A(n1035), .ZN(n1047) );
NAND3_X1 U759 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1017) );
NAND3_X1 U760 ( .A1(n1053), .A2(n1054), .A3(n1027), .ZN(n1052) );
NOR3_X1 U761 ( .A1(n1039), .A2(n1044), .A3(n1035), .ZN(n1027) );
NAND2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
OR2_X1 U763 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR3_X1 U764 ( .A1(n1059), .A2(G953), .A3(G952), .ZN(n1015) );
INV_X1 U765 ( .A(n1050), .ZN(n1059) );
NAND4_X1 U766 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1050) );
NOR4_X1 U767 ( .A1(n1064), .A2(n1065), .A3(n1022), .A4(n1066), .ZN(n1063) );
XOR2_X1 U768 ( .A(n1067), .B(KEYINPUT16), .Z(n1064) );
NAND3_X1 U769 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NAND2_X1 U770 ( .A1(KEYINPUT20), .A2(n1071), .ZN(n1070) );
OR3_X1 U771 ( .A1(n1072), .A2(KEYINPUT20), .A3(G472), .ZN(n1069) );
NAND2_X1 U772 ( .A1(G472), .A2(n1072), .ZN(n1068) );
NAND2_X1 U773 ( .A1(KEYINPUT47), .A2(n1073), .ZN(n1072) );
NOR3_X1 U774 ( .A1(n1074), .A2(n1075), .A3(n1031), .ZN(n1062) );
NAND2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1061) );
XNOR2_X1 U776 ( .A(n1078), .B(KEYINPUT1), .ZN(n1076) );
NAND2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1060) );
XOR2_X1 U778 ( .A(n1081), .B(n1082), .Z(G72) );
NOR2_X1 U779 ( .A1(n1083), .A2(n1051), .ZN(n1082) );
NOR2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U781 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
NAND2_X1 U782 ( .A1(n1088), .A2(n1051), .ZN(n1087) );
XOR2_X1 U783 ( .A(n1020), .B(n1089), .Z(n1088) );
NAND3_X1 U784 ( .A1(G900), .A2(n1089), .A3(G953), .ZN(n1086) );
XNOR2_X1 U785 ( .A(n1090), .B(n1091), .ZN(n1089) );
XNOR2_X1 U786 ( .A(n1092), .B(n1093), .ZN(n1091) );
XNOR2_X1 U787 ( .A(G125), .B(n1094), .ZN(n1093) );
NAND2_X1 U788 ( .A1(KEYINPUT57), .A2(G140), .ZN(n1094) );
XNOR2_X1 U789 ( .A(n1095), .B(n1096), .ZN(n1090) );
XOR2_X1 U790 ( .A(n1097), .B(n1098), .Z(G69) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U792 ( .A1(G953), .A2(n1101), .ZN(n1100) );
NAND2_X1 U793 ( .A1(n1102), .A2(G224), .ZN(n1101) );
XNOR2_X1 U794 ( .A(G898), .B(KEYINPUT21), .ZN(n1102) );
NAND3_X1 U795 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1099) );
XOR2_X1 U796 ( .A(KEYINPUT2), .B(n1106), .Z(n1105) );
NOR2_X1 U797 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U798 ( .A1(n1108), .A2(n1107), .ZN(n1104) );
XNOR2_X1 U799 ( .A(n1109), .B(n1110), .ZN(n1108) );
XNOR2_X1 U800 ( .A(n1111), .B(KEYINPUT39), .ZN(n1109) );
NAND2_X1 U801 ( .A1(G953), .A2(n1112), .ZN(n1103) );
NOR2_X1 U802 ( .A1(n1113), .A2(G953), .ZN(n1097) );
NOR2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(G66) );
XNOR2_X1 U804 ( .A(n1116), .B(KEYINPUT46), .ZN(n1115) );
NOR3_X1 U805 ( .A1(n1117), .A2(n1079), .A3(n1118), .ZN(n1114) );
NOR2_X1 U806 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1080), .ZN(n1119) );
XOR2_X1 U808 ( .A(n1122), .B(KEYINPUT26), .Z(n1117) );
NAND3_X1 U809 ( .A1(n1120), .A2(n1123), .A3(n1124), .ZN(n1122) );
INV_X1 U810 ( .A(n1080), .ZN(n1123) );
NOR2_X1 U811 ( .A1(n1125), .A2(n1126), .ZN(G63) );
XOR2_X1 U812 ( .A(KEYINPUT8), .B(n1116), .Z(n1126) );
XOR2_X1 U813 ( .A(n1127), .B(n1128), .Z(n1125) );
XOR2_X1 U814 ( .A(KEYINPUT3), .B(n1129), .Z(n1128) );
AND2_X1 U815 ( .A1(G478), .A2(n1124), .ZN(n1129) );
NOR2_X1 U816 ( .A1(n1116), .A2(n1130), .ZN(G60) );
XOR2_X1 U817 ( .A(n1131), .B(n1132), .Z(n1130) );
NAND2_X1 U818 ( .A1(n1124), .A2(G475), .ZN(n1131) );
XNOR2_X1 U819 ( .A(G104), .B(n1133), .ZN(G6) );
NOR2_X1 U820 ( .A1(n1116), .A2(n1134), .ZN(G57) );
XOR2_X1 U821 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U822 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U823 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U824 ( .A(n1141), .B(KEYINPUT7), .Z(n1140) );
NOR2_X1 U825 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
AND3_X1 U826 ( .A1(G210), .A2(n1144), .A3(n1145), .ZN(n1137) );
INV_X1 U827 ( .A(KEYINPUT43), .ZN(n1144) );
XOR2_X1 U828 ( .A(n1146), .B(n1147), .Z(n1135) );
NAND2_X1 U829 ( .A1(n1124), .A2(G472), .ZN(n1146) );
NOR2_X1 U830 ( .A1(n1116), .A2(n1148), .ZN(G54) );
XOR2_X1 U831 ( .A(n1149), .B(n1150), .Z(n1148) );
AND2_X1 U832 ( .A1(G469), .A2(n1124), .ZN(n1150) );
NAND2_X1 U833 ( .A1(n1151), .A2(KEYINPUT52), .ZN(n1149) );
XOR2_X1 U834 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U835 ( .A(n1154), .B(n1155), .ZN(n1153) );
NAND3_X1 U836 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1154) );
OR2_X1 U837 ( .A1(n1092), .A2(KEYINPUT14), .ZN(n1158) );
NAND3_X1 U838 ( .A1(KEYINPUT14), .A2(n1092), .A3(n1159), .ZN(n1157) );
NAND2_X1 U839 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
NAND2_X1 U840 ( .A1(n1162), .A2(KEYINPUT14), .ZN(n1161) );
XNOR2_X1 U841 ( .A(n1163), .B(KEYINPUT5), .ZN(n1162) );
NOR2_X1 U842 ( .A1(n1116), .A2(n1164), .ZN(G51) );
XOR2_X1 U843 ( .A(n1165), .B(n1166), .Z(n1164) );
AND2_X1 U844 ( .A1(n1078), .A2(n1124), .ZN(n1166) );
NOR2_X1 U845 ( .A1(n1167), .A2(n1121), .ZN(n1124) );
AND2_X1 U846 ( .A1(n1113), .A2(n1168), .ZN(n1121) );
XNOR2_X1 U847 ( .A(KEYINPUT13), .B(n1020), .ZN(n1168) );
NAND4_X1 U848 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1020) );
AND4_X1 U849 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172) );
NOR2_X1 U850 ( .A1(n1177), .A2(n1178), .ZN(n1171) );
NAND2_X1 U851 ( .A1(n1029), .A2(n1179), .ZN(n1169) );
XOR2_X1 U852 ( .A(KEYINPUT15), .B(n1180), .Z(n1179) );
INV_X1 U853 ( .A(n1018), .ZN(n1113) );
NAND4_X1 U854 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1018) );
AND4_X1 U855 ( .A1(n1014), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1184) );
NAND3_X1 U856 ( .A1(n1045), .A2(n1188), .A3(n1189), .ZN(n1014) );
AND2_X1 U857 ( .A1(n1190), .A2(n1133), .ZN(n1183) );
NAND3_X1 U858 ( .A1(n1189), .A2(n1188), .A3(n1046), .ZN(n1133) );
NAND2_X1 U859 ( .A1(n1191), .A2(KEYINPUT19), .ZN(n1165) );
XNOR2_X1 U860 ( .A(n1192), .B(n1193), .ZN(n1191) );
NOR2_X1 U861 ( .A1(n1051), .A2(G952), .ZN(n1116) );
XOR2_X1 U862 ( .A(G146), .B(n1177), .Z(G48) );
AND3_X1 U863 ( .A1(n1046), .A2(n1029), .A3(n1194), .ZN(n1177) );
XNOR2_X1 U864 ( .A(G143), .B(n1170), .ZN(G45) );
NAND4_X1 U865 ( .A1(n1195), .A2(n1029), .A3(n1042), .A4(n1196), .ZN(n1170) );
NOR3_X1 U866 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
XNOR2_X1 U867 ( .A(G140), .B(n1176), .ZN(G42) );
NAND3_X1 U868 ( .A1(n1046), .A2(n1041), .A3(n1200), .ZN(n1176) );
XOR2_X1 U869 ( .A(G137), .B(n1178), .Z(G39) );
AND3_X1 U870 ( .A1(n1053), .A2(n1201), .A3(n1194), .ZN(n1178) );
INV_X1 U871 ( .A(n1032), .ZN(n1053) );
XNOR2_X1 U872 ( .A(G134), .B(n1175), .ZN(G36) );
NAND3_X1 U873 ( .A1(n1042), .A2(n1045), .A3(n1200), .ZN(n1175) );
XNOR2_X1 U874 ( .A(G131), .B(n1174), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1042), .A2(n1046), .A3(n1200), .ZN(n1174) );
NOR3_X1 U876 ( .A1(n1055), .A2(n1198), .A3(n1032), .ZN(n1200) );
NAND2_X1 U877 ( .A1(n1030), .A2(n1202), .ZN(n1032) );
INV_X1 U878 ( .A(n1203), .ZN(n1198) );
XNOR2_X1 U879 ( .A(G128), .B(n1204), .ZN(G30) );
NAND2_X1 U880 ( .A1(n1180), .A2(n1029), .ZN(n1204) );
AND2_X1 U881 ( .A1(n1194), .A2(n1045), .ZN(n1180) );
AND4_X1 U882 ( .A1(n1205), .A2(n1206), .A3(n1195), .A4(n1203), .ZN(n1194) );
XNOR2_X1 U883 ( .A(G101), .B(n1190), .ZN(G3) );
NAND3_X1 U884 ( .A1(n1201), .A2(n1188), .A3(n1042), .ZN(n1190) );
XNOR2_X1 U885 ( .A(G125), .B(n1173), .ZN(G27) );
NAND3_X1 U886 ( .A1(n1046), .A2(n1041), .A3(n1207), .ZN(n1173) );
AND3_X1 U887 ( .A1(n1208), .A2(n1203), .A3(n1029), .ZN(n1207) );
NAND2_X1 U888 ( .A1(n1209), .A2(n1035), .ZN(n1203) );
XOR2_X1 U889 ( .A(n1210), .B(KEYINPUT25), .Z(n1209) );
NAND4_X1 U890 ( .A1(G953), .A2(G902), .A3(n1211), .A4(n1085), .ZN(n1210) );
INV_X1 U891 ( .A(G900), .ZN(n1085) );
NAND2_X1 U892 ( .A1(n1212), .A2(n1213), .ZN(G24) );
NAND2_X1 U893 ( .A1(G122), .A2(n1181), .ZN(n1213) );
XOR2_X1 U894 ( .A(KEYINPUT63), .B(n1214), .Z(n1212) );
NOR2_X1 U895 ( .A1(G122), .A2(n1181), .ZN(n1214) );
NAND4_X1 U896 ( .A1(n1215), .A2(n1189), .A3(n1065), .A4(n1066), .ZN(n1181) );
INV_X1 U897 ( .A(n1044), .ZN(n1189) );
NAND2_X1 U898 ( .A1(n1216), .A2(n1217), .ZN(n1044) );
XNOR2_X1 U899 ( .A(n1218), .B(KEYINPUT32), .ZN(n1216) );
XOR2_X1 U900 ( .A(n1182), .B(n1219), .Z(G21) );
NAND2_X1 U901 ( .A1(KEYINPUT58), .A2(G119), .ZN(n1219) );
NAND4_X1 U902 ( .A1(n1206), .A2(n1215), .A3(n1205), .A4(n1201), .ZN(n1182) );
XNOR2_X1 U903 ( .A(G116), .B(n1187), .ZN(G18) );
NAND3_X1 U904 ( .A1(n1215), .A2(n1045), .A3(n1042), .ZN(n1187) );
AND2_X1 U905 ( .A1(n1220), .A2(n1066), .ZN(n1045) );
XNOR2_X1 U906 ( .A(KEYINPUT34), .B(n1197), .ZN(n1220) );
XNOR2_X1 U907 ( .A(G113), .B(n1186), .ZN(G15) );
NAND3_X1 U908 ( .A1(n1215), .A2(n1046), .A3(n1042), .ZN(n1186) );
INV_X1 U909 ( .A(n1049), .ZN(n1042) );
NAND2_X1 U910 ( .A1(n1206), .A2(n1217), .ZN(n1049) );
XNOR2_X1 U911 ( .A(n1218), .B(KEYINPUT42), .ZN(n1206) );
AND2_X1 U912 ( .A1(n1221), .A2(n1065), .ZN(n1046) );
XNOR2_X1 U913 ( .A(n1066), .B(KEYINPUT36), .ZN(n1221) );
AND2_X1 U914 ( .A1(n1208), .A2(n1222), .ZN(n1215) );
INV_X1 U915 ( .A(n1022), .ZN(n1208) );
NAND2_X1 U916 ( .A1(n1223), .A2(n1058), .ZN(n1022) );
XOR2_X1 U917 ( .A(n1185), .B(n1224), .Z(G12) );
XNOR2_X1 U918 ( .A(KEYINPUT10), .B(n1155), .ZN(n1224) );
NAND3_X1 U919 ( .A1(n1041), .A2(n1188), .A3(n1201), .ZN(n1185) );
INV_X1 U920 ( .A(n1039), .ZN(n1201) );
NAND2_X1 U921 ( .A1(n1199), .A2(n1225), .ZN(n1039) );
XNOR2_X1 U922 ( .A(KEYINPUT6), .B(n1197), .ZN(n1225) );
INV_X1 U923 ( .A(n1065), .ZN(n1197) );
XNOR2_X1 U924 ( .A(n1226), .B(G475), .ZN(n1065) );
NAND2_X1 U925 ( .A1(n1132), .A2(n1167), .ZN(n1226) );
XNOR2_X1 U926 ( .A(n1227), .B(n1228), .ZN(n1132) );
XOR2_X1 U927 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U928 ( .A(n1231), .B(G140), .ZN(n1230) );
XOR2_X1 U929 ( .A(KEYINPUT9), .B(G146), .Z(n1229) );
XOR2_X1 U930 ( .A(n1232), .B(n1233), .Z(n1227) );
XNOR2_X1 U931 ( .A(n1193), .B(n1234), .ZN(n1233) );
NOR2_X1 U932 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U933 ( .A(n1237), .B(KEYINPUT22), .Z(n1236) );
NAND2_X1 U934 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XNOR2_X1 U935 ( .A(G104), .B(KEYINPUT12), .ZN(n1238) );
NOR2_X1 U936 ( .A1(G104), .A2(n1239), .ZN(n1235) );
XNOR2_X1 U937 ( .A(n1240), .B(n1241), .ZN(n1239) );
XOR2_X1 U938 ( .A(n1242), .B(n1243), .Z(n1232) );
AND2_X1 U939 ( .A1(n1145), .A2(G214), .ZN(n1243) );
NAND2_X1 U940 ( .A1(KEYINPUT18), .A2(n1095), .ZN(n1242) );
INV_X1 U941 ( .A(n1066), .ZN(n1199) );
XNOR2_X1 U942 ( .A(n1244), .B(G478), .ZN(n1066) );
OR2_X1 U943 ( .A1(n1127), .A2(G902), .ZN(n1244) );
XNOR2_X1 U944 ( .A(n1245), .B(n1246), .ZN(n1127) );
XOR2_X1 U945 ( .A(n1247), .B(n1248), .Z(n1246) );
XNOR2_X1 U946 ( .A(n1249), .B(n1250), .ZN(n1248) );
NAND2_X1 U947 ( .A1(KEYINPUT37), .A2(G143), .ZN(n1250) );
NAND2_X1 U948 ( .A1(KEYINPUT40), .A2(n1251), .ZN(n1249) );
XNOR2_X1 U949 ( .A(G116), .B(n1252), .ZN(n1251) );
NAND2_X1 U950 ( .A1(KEYINPUT29), .A2(n1240), .ZN(n1252) );
INV_X1 U951 ( .A(G122), .ZN(n1240) );
NAND3_X1 U952 ( .A1(G234), .A2(n1051), .A3(G217), .ZN(n1247) );
XNOR2_X1 U953 ( .A(G107), .B(n1253), .ZN(n1245) );
XNOR2_X1 U954 ( .A(G134), .B(n1254), .ZN(n1253) );
AND2_X1 U955 ( .A1(n1195), .A2(n1222), .ZN(n1188) );
AND2_X1 U956 ( .A1(n1029), .A2(n1255), .ZN(n1222) );
NAND2_X1 U957 ( .A1(n1035), .A2(n1256), .ZN(n1255) );
NAND4_X1 U958 ( .A1(G953), .A2(G902), .A3(n1211), .A4(n1112), .ZN(n1256) );
INV_X1 U959 ( .A(G898), .ZN(n1112) );
NAND3_X1 U960 ( .A1(n1211), .A2(n1051), .A3(G952), .ZN(n1035) );
NAND2_X1 U961 ( .A1(G237), .A2(G234), .ZN(n1211) );
NOR2_X1 U962 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
INV_X1 U963 ( .A(n1202), .ZN(n1031) );
NAND2_X1 U964 ( .A1(G214), .A2(n1257), .ZN(n1202) );
NOR2_X1 U965 ( .A1(n1074), .A2(n1258), .ZN(n1030) );
AND2_X1 U966 ( .A1(n1259), .A2(n1077), .ZN(n1258) );
XNOR2_X1 U967 ( .A(n1078), .B(KEYINPUT35), .ZN(n1259) );
NOR2_X1 U968 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
AND2_X1 U969 ( .A1(G210), .A2(n1257), .ZN(n1078) );
NAND2_X1 U970 ( .A1(n1260), .A2(n1167), .ZN(n1257) );
INV_X1 U971 ( .A(G237), .ZN(n1260) );
NAND2_X1 U972 ( .A1(n1261), .A2(n1167), .ZN(n1077) );
XOR2_X1 U973 ( .A(n1262), .B(n1192), .Z(n1261) );
XOR2_X1 U974 ( .A(n1263), .B(n1264), .Z(n1192) );
XOR2_X1 U975 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U976 ( .A(n1267), .B(n1268), .ZN(n1266) );
NOR2_X1 U977 ( .A1(KEYINPUT54), .A2(n1269), .ZN(n1268) );
INV_X1 U978 ( .A(n1111), .ZN(n1269) );
NOR2_X1 U979 ( .A1(KEYINPUT0), .A2(n1107), .ZN(n1267) );
XNOR2_X1 U980 ( .A(n1155), .B(G122), .ZN(n1107) );
NAND2_X1 U981 ( .A1(G224), .A2(n1051), .ZN(n1265) );
XOR2_X1 U982 ( .A(n1142), .B(n1110), .Z(n1263) );
XNOR2_X1 U983 ( .A(n1270), .B(G101), .ZN(n1110) );
NAND3_X1 U984 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
NAND2_X1 U985 ( .A1(KEYINPUT49), .A2(G107), .ZN(n1273) );
OR3_X1 U986 ( .A1(n1274), .A2(KEYINPUT49), .A3(n1275), .ZN(n1272) );
NAND2_X1 U987 ( .A1(n1275), .A2(n1274), .ZN(n1271) );
NAND2_X1 U988 ( .A1(KEYINPUT48), .A2(n1276), .ZN(n1274) );
XOR2_X1 U989 ( .A(G104), .B(KEYINPUT53), .Z(n1275) );
NAND2_X1 U990 ( .A1(KEYINPUT59), .A2(n1277), .ZN(n1262) );
XNOR2_X1 U991 ( .A(KEYINPUT55), .B(n1193), .ZN(n1277) );
INV_X1 U992 ( .A(n1055), .ZN(n1195) );
NAND2_X1 U993 ( .A1(n1278), .A2(n1057), .ZN(n1055) );
INV_X1 U994 ( .A(n1223), .ZN(n1057) );
XOR2_X1 U995 ( .A(n1279), .B(G469), .Z(n1223) );
NAND2_X1 U996 ( .A1(n1280), .A2(n1167), .ZN(n1279) );
XOR2_X1 U997 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U998 ( .A(n1152), .B(n1159), .ZN(n1282) );
INV_X1 U999 ( .A(n1160), .ZN(n1159) );
XNOR2_X1 U1000 ( .A(n1283), .B(n1284), .ZN(n1160) );
XNOR2_X1 U1001 ( .A(n1276), .B(G101), .ZN(n1284) );
INV_X1 U1002 ( .A(G107), .ZN(n1276) );
NAND2_X1 U1003 ( .A1(KEYINPUT50), .A2(n1285), .ZN(n1283) );
INV_X1 U1004 ( .A(G104), .ZN(n1285) );
XOR2_X1 U1005 ( .A(n1143), .B(n1286), .Z(n1152) );
XNOR2_X1 U1006 ( .A(n1287), .B(n1288), .ZN(n1286) );
NOR2_X1 U1007 ( .A1(G953), .A2(n1084), .ZN(n1288) );
INV_X1 U1008 ( .A(G227), .ZN(n1084) );
XNOR2_X1 U1009 ( .A(n1289), .B(n1290), .ZN(n1281) );
NAND2_X1 U1010 ( .A1(KEYINPUT62), .A2(n1092), .ZN(n1290) );
INV_X1 U1011 ( .A(n1163), .ZN(n1092) );
XNOR2_X1 U1012 ( .A(n1291), .B(n1292), .ZN(n1163) );
XNOR2_X1 U1013 ( .A(G143), .B(n1293), .ZN(n1292) );
NAND2_X1 U1014 ( .A1(KEYINPUT33), .A2(G146), .ZN(n1293) );
NAND2_X1 U1015 ( .A1(KEYINPUT38), .A2(n1254), .ZN(n1291) );
NAND2_X1 U1016 ( .A1(KEYINPUT56), .A2(n1155), .ZN(n1289) );
INV_X1 U1017 ( .A(G110), .ZN(n1155) );
XOR2_X1 U1018 ( .A(n1058), .B(KEYINPUT30), .Z(n1278) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1294), .ZN(n1058) );
AND2_X1 U1020 ( .A1(n1205), .A2(n1218), .ZN(n1041) );
AND2_X1 U1021 ( .A1(n1295), .A2(n1296), .ZN(n1218) );
NAND2_X1 U1022 ( .A1(n1071), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1023 ( .A(KEYINPUT61), .B(n1298), .Z(n1295) );
NOR2_X1 U1024 ( .A1(n1071), .A2(n1297), .ZN(n1298) );
INV_X1 U1025 ( .A(G472), .ZN(n1297) );
INV_X1 U1026 ( .A(n1073), .ZN(n1071) );
NAND2_X1 U1027 ( .A1(n1299), .A2(n1167), .ZN(n1073) );
XOR2_X1 U1028 ( .A(n1147), .B(n1300), .Z(n1299) );
XOR2_X1 U1029 ( .A(n1301), .B(n1302), .Z(n1300) );
NAND3_X1 U1030 ( .A1(G210), .A2(n1145), .A3(KEYINPUT28), .ZN(n1302) );
NOR2_X1 U1031 ( .A1(G953), .A2(G237), .ZN(n1145) );
NAND2_X1 U1032 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
OR2_X1 U1033 ( .A1(n1143), .A2(n1142), .ZN(n1304) );
XOR2_X1 U1034 ( .A(n1141), .B(KEYINPUT41), .Z(n1303) );
NAND2_X1 U1035 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XNOR2_X1 U1036 ( .A(n1095), .B(n1305), .ZN(n1143) );
NOR2_X1 U1037 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
AND3_X1 U1038 ( .A1(KEYINPUT51), .A2(n1308), .A3(G134), .ZN(n1307) );
NOR2_X1 U1039 ( .A1(KEYINPUT51), .A2(n1096), .ZN(n1306) );
XNOR2_X1 U1040 ( .A(G134), .B(n1308), .ZN(n1096) );
INV_X1 U1041 ( .A(G137), .ZN(n1308) );
XOR2_X1 U1042 ( .A(G131), .B(KEYINPUT60), .Z(n1095) );
XOR2_X1 U1043 ( .A(n1309), .B(n1310), .Z(n1142) );
XNOR2_X1 U1044 ( .A(G146), .B(n1231), .ZN(n1310) );
INV_X1 U1045 ( .A(G143), .ZN(n1231) );
NAND2_X1 U1046 ( .A1(KEYINPUT24), .A2(G128), .ZN(n1309) );
XNOR2_X1 U1047 ( .A(n1311), .B(n1111), .ZN(n1147) );
XNOR2_X1 U1048 ( .A(n1312), .B(n1241), .ZN(n1111) );
XOR2_X1 U1049 ( .A(G113), .B(KEYINPUT45), .Z(n1241) );
XNOR2_X1 U1050 ( .A(G116), .B(G119), .ZN(n1312) );
INV_X1 U1051 ( .A(G101), .ZN(n1311) );
XNOR2_X1 U1052 ( .A(n1217), .B(KEYINPUT11), .ZN(n1205) );
NOR2_X1 U1053 ( .A1(n1313), .A2(n1075), .ZN(n1217) );
NOR2_X1 U1054 ( .A1(n1080), .A2(n1079), .ZN(n1075) );
AND2_X1 U1055 ( .A1(n1314), .A2(n1080), .ZN(n1313) );
NAND2_X1 U1056 ( .A1(G217), .A2(n1294), .ZN(n1080) );
NAND2_X1 U1057 ( .A1(G234), .A2(n1167), .ZN(n1294) );
INV_X1 U1058 ( .A(G902), .ZN(n1167) );
XOR2_X1 U1059 ( .A(KEYINPUT23), .B(n1079), .Z(n1314) );
NOR2_X1 U1060 ( .A1(n1120), .A2(G902), .ZN(n1079) );
XOR2_X1 U1061 ( .A(n1315), .B(n1316), .Z(n1120) );
XOR2_X1 U1062 ( .A(G137), .B(n1317), .Z(n1316) );
AND3_X1 U1063 ( .A1(G234), .A2(n1051), .A3(G221), .ZN(n1317) );
INV_X1 U1064 ( .A(G953), .ZN(n1051) );
NAND2_X1 U1065 ( .A1(n1318), .A2(KEYINPUT27), .ZN(n1315) );
XOR2_X1 U1066 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1067 ( .A(n1193), .B(n1321), .ZN(n1320) );
XOR2_X1 U1068 ( .A(KEYINPUT4), .B(G146), .Z(n1321) );
INV_X1 U1069 ( .A(G125), .ZN(n1193) );
XOR2_X1 U1070 ( .A(n1322), .B(n1323), .Z(n1319) );
XNOR2_X1 U1071 ( .A(G110), .B(n1324), .ZN(n1323) );
NAND2_X1 U1072 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
OR2_X1 U1073 ( .A1(n1254), .A2(G119), .ZN(n1326) );
XOR2_X1 U1074 ( .A(n1327), .B(KEYINPUT17), .Z(n1325) );
NAND2_X1 U1075 ( .A1(G119), .A2(n1254), .ZN(n1327) );
INV_X1 U1076 ( .A(G128), .ZN(n1254) );
NAND2_X1 U1077 ( .A1(KEYINPUT44), .A2(n1287), .ZN(n1322) );
INV_X1 U1078 ( .A(G140), .ZN(n1287) );
endmodule


