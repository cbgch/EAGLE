//Key = 0110100100010010000010001011010111101000100101110100000110101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339;

XOR2_X1 U731 ( .A(n1013), .B(n1014), .Z(G9) );
NAND2_X1 U732 ( .A1(KEYINPUT11), .A2(n1015), .ZN(n1013) );
NOR2_X1 U733 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U734 ( .A1(G953), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1017) );
NOR2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U737 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR2_X1 U738 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U739 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U741 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U743 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U744 ( .A1(n1039), .A2(n1040), .ZN(n1031) );
NOR2_X1 U745 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR3_X1 U747 ( .A1(n1034), .A2(n1045), .A3(n1040), .ZN(n1027) );
NOR2_X1 U748 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR4_X1 U750 ( .A1(n1050), .A2(n1040), .A3(n1034), .A4(n1030), .ZN(n1023) );
INV_X1 U751 ( .A(n1051), .ZN(n1034) );
INV_X1 U752 ( .A(n1052), .ZN(n1040) );
NOR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
NOR3_X1 U754 ( .A1(n1018), .A2(G953), .A3(G952), .ZN(n1016) );
AND2_X1 U755 ( .A1(n1055), .A2(n1056), .ZN(n1018) );
NOR4_X1 U756 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
XNOR2_X1 U757 ( .A(n1061), .B(n1062), .ZN(n1059) );
NAND2_X1 U758 ( .A1(KEYINPUT58), .A2(n1063), .ZN(n1061) );
XNOR2_X1 U759 ( .A(n1064), .B(KEYINPUT45), .ZN(n1058) );
NOR4_X1 U760 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1055) );
XNOR2_X1 U761 ( .A(G475), .B(n1069), .ZN(n1068) );
NAND2_X1 U762 ( .A1(KEYINPUT56), .A2(n1070), .ZN(n1069) );
XOR2_X1 U763 ( .A(n1071), .B(n1072), .Z(n1067) );
XNOR2_X1 U764 ( .A(KEYINPUT40), .B(n1073), .ZN(n1072) );
NOR2_X1 U765 ( .A1(KEYINPUT42), .A2(n1074), .ZN(n1073) );
INV_X1 U766 ( .A(n1075), .ZN(n1074) );
NOR2_X1 U767 ( .A1(n1076), .A2(n1077), .ZN(n1066) );
INV_X1 U768 ( .A(KEYINPUT50), .ZN(n1077) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR2_X1 U770 ( .A1(KEYINPUT50), .A2(n1051), .ZN(n1065) );
XOR2_X1 U771 ( .A(n1080), .B(n1081), .Z(G72) );
NOR2_X1 U772 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U773 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U774 ( .A(n1086), .B(n1087), .ZN(n1085) );
XOR2_X1 U775 ( .A(n1088), .B(n1089), .Z(n1084) );
NOR2_X1 U776 ( .A1(KEYINPUT12), .A2(G134), .ZN(n1089) );
XNOR2_X1 U777 ( .A(G125), .B(KEYINPUT6), .ZN(n1088) );
NAND3_X1 U778 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1080) );
INV_X1 U779 ( .A(n1082), .ZN(n1091) );
NOR2_X1 U780 ( .A1(n1093), .A2(G900), .ZN(n1082) );
OR2_X1 U781 ( .A1(n1093), .A2(G227), .ZN(n1090) );
XOR2_X1 U782 ( .A(n1094), .B(n1095), .Z(G69) );
XOR2_X1 U783 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U785 ( .A(KEYINPUT30), .B(n1093), .ZN(n1099) );
NAND2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
NAND2_X1 U787 ( .A1(G953), .A2(n1102), .ZN(n1101) );
XNOR2_X1 U788 ( .A(n1103), .B(n1104), .ZN(n1100) );
XNOR2_X1 U789 ( .A(n1105), .B(n1106), .ZN(n1104) );
NAND2_X1 U790 ( .A1(G953), .A2(n1107), .ZN(n1094) );
NAND2_X1 U791 ( .A1(G898), .A2(G224), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XNOR2_X1 U793 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U794 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U795 ( .A1(n1108), .A2(n1114), .ZN(G63) );
NOR3_X1 U796 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
AND3_X1 U797 ( .A1(n1118), .A2(G478), .A3(n1119), .ZN(n1117) );
NOR2_X1 U798 ( .A1(n1120), .A2(n1118), .ZN(n1116) );
AND2_X1 U799 ( .A1(n1020), .A2(G478), .ZN(n1120) );
NOR2_X1 U800 ( .A1(n1108), .A2(n1121), .ZN(G60) );
XOR2_X1 U801 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U802 ( .A1(n1124), .A2(n1113), .ZN(n1122) );
XOR2_X1 U803 ( .A(G104), .B(n1125), .Z(G6) );
NOR2_X1 U804 ( .A1(n1108), .A2(n1126), .ZN(G57) );
XOR2_X1 U805 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U806 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR3_X1 U807 ( .A1(KEYINPUT17), .A2(n1131), .A3(n1132), .ZN(n1130) );
NOR2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U809 ( .A(n1135), .B(KEYINPUT38), .Z(n1134) );
AND2_X1 U810 ( .A1(n1135), .A2(n1133), .ZN(n1131) );
XOR2_X1 U811 ( .A(n1136), .B(n1137), .Z(n1133) );
XNOR2_X1 U812 ( .A(KEYINPUT20), .B(n1138), .ZN(n1136) );
NOR2_X1 U813 ( .A1(KEYINPUT59), .A2(n1139), .ZN(n1138) );
NAND2_X1 U814 ( .A1(n1119), .A2(G472), .ZN(n1135) );
NAND2_X1 U815 ( .A1(KEYINPUT60), .A2(n1140), .ZN(n1127) );
NOR3_X1 U816 ( .A1(n1108), .A2(n1141), .A3(n1142), .ZN(G54) );
AND4_X1 U817 ( .A1(n1143), .A2(KEYINPUT26), .A3(G469), .A4(n1119), .ZN(n1142) );
INV_X1 U818 ( .A(n1113), .ZN(n1119) );
NOR2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NOR3_X1 U820 ( .A1(n1113), .A2(n1145), .A3(n1146), .ZN(n1144) );
NOR2_X1 U821 ( .A1(KEYINPUT26), .A2(n1147), .ZN(n1145) );
NOR2_X1 U822 ( .A1(KEYINPUT21), .A2(n1148), .ZN(n1143) );
INV_X1 U823 ( .A(n1147), .ZN(n1148) );
XNOR2_X1 U824 ( .A(n1149), .B(KEYINPUT4), .ZN(n1147) );
NOR2_X1 U825 ( .A1(n1108), .A2(n1150), .ZN(G51) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U827 ( .A1(n1075), .A2(n1113), .ZN(n1152) );
NAND2_X1 U828 ( .A1(G902), .A2(n1020), .ZN(n1113) );
NAND2_X1 U829 ( .A1(n1098), .A2(n1092), .ZN(n1020) );
AND2_X1 U830 ( .A1(n1153), .A2(n1154), .ZN(n1092) );
NOR4_X1 U831 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
NOR4_X1 U832 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1153) );
NOR2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR3_X1 U834 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1161) );
XNOR2_X1 U835 ( .A(n1042), .B(KEYINPUT15), .ZN(n1166) );
NOR2_X1 U836 ( .A1(n1168), .A2(n1169), .ZN(n1160) );
XNOR2_X1 U837 ( .A(n1170), .B(KEYINPUT18), .ZN(n1168) );
INV_X1 U838 ( .A(n1171), .ZN(n1159) );
AND2_X1 U839 ( .A1(n1172), .A2(n1173), .ZN(n1098) );
NOR4_X1 U840 ( .A1(n1174), .A2(n1014), .A3(n1175), .A4(n1125), .ZN(n1173) );
AND2_X1 U841 ( .A1(n1054), .A2(n1176), .ZN(n1125) );
NOR4_X1 U842 ( .A1(n1177), .A2(n1026), .A3(n1178), .A4(n1179), .ZN(n1175) );
NAND2_X1 U843 ( .A1(n1180), .A2(n1036), .ZN(n1177) );
XOR2_X1 U844 ( .A(n1181), .B(KEYINPUT37), .Z(n1180) );
AND2_X1 U845 ( .A1(n1053), .A2(n1176), .ZN(n1014) );
AND4_X1 U846 ( .A1(n1042), .A2(n1052), .A3(n1047), .A4(n1181), .ZN(n1176) );
AND4_X1 U847 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1172) );
NAND2_X1 U848 ( .A1(n1186), .A2(KEYINPUT1), .ZN(n1151) );
XOR2_X1 U849 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U850 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U851 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
AND3_X1 U852 ( .A1(KEYINPUT44), .A2(n1193), .A3(G125), .ZN(n1192) );
NOR2_X1 U853 ( .A1(KEYINPUT44), .A2(n1194), .ZN(n1191) );
XNOR2_X1 U854 ( .A(G125), .B(n1193), .ZN(n1194) );
XOR2_X1 U855 ( .A(KEYINPUT51), .B(n1195), .Z(n1187) );
NOR2_X1 U856 ( .A1(n1093), .A2(G952), .ZN(n1108) );
XOR2_X1 U857 ( .A(n1157), .B(n1196), .Z(G48) );
NOR2_X1 U858 ( .A1(KEYINPUT0), .A2(n1197), .ZN(n1196) );
AND3_X1 U859 ( .A1(n1054), .A2(n1047), .A3(n1198), .ZN(n1157) );
XNOR2_X1 U860 ( .A(G143), .B(n1171), .ZN(G45) );
NAND3_X1 U861 ( .A1(n1199), .A2(n1036), .A3(n1200), .ZN(n1171) );
NOR3_X1 U862 ( .A1(n1178), .A2(n1201), .A3(n1202), .ZN(n1200) );
XNOR2_X1 U863 ( .A(n1203), .B(n1158), .ZN(G42) );
AND4_X1 U864 ( .A1(n1204), .A2(n1064), .A3(n1054), .A4(n1205), .ZN(n1158) );
NOR2_X1 U865 ( .A1(n1206), .A2(n1030), .ZN(n1205) );
XOR2_X1 U866 ( .A(G137), .B(n1207), .Z(G39) );
NOR2_X1 U867 ( .A1(n1030), .A2(n1169), .ZN(n1207) );
NAND2_X1 U868 ( .A1(n1198), .A2(n1208), .ZN(n1169) );
INV_X1 U869 ( .A(n1170), .ZN(n1030) );
XOR2_X1 U870 ( .A(G134), .B(n1156), .Z(G36) );
AND3_X1 U871 ( .A1(n1053), .A2(n1042), .A3(n1209), .ZN(n1156) );
NAND3_X1 U872 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(G33) );
NAND4_X1 U873 ( .A1(n1209), .A2(n1054), .A3(n1042), .A4(n1213), .ZN(n1212) );
NAND2_X1 U874 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U875 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U876 ( .A1(KEYINPUT25), .A2(n1216), .ZN(n1211) );
NAND3_X1 U877 ( .A1(n1218), .A2(n1214), .A3(G131), .ZN(n1210) );
INV_X1 U878 ( .A(KEYINPUT25), .ZN(n1214) );
NAND4_X1 U879 ( .A1(n1209), .A2(n1054), .A3(n1042), .A4(n1217), .ZN(n1218) );
INV_X1 U880 ( .A(KEYINPUT28), .ZN(n1217) );
INV_X1 U881 ( .A(n1165), .ZN(n1209) );
NAND3_X1 U882 ( .A1(n1036), .A2(n1219), .A3(n1170), .ZN(n1165) );
NOR2_X1 U883 ( .A1(n1048), .A2(n1057), .ZN(n1170) );
XOR2_X1 U884 ( .A(n1220), .B(KEYINPUT39), .Z(n1048) );
XNOR2_X1 U885 ( .A(n1221), .B(n1155), .ZN(G30) );
AND3_X1 U886 ( .A1(n1053), .A2(n1047), .A3(n1198), .ZN(n1155) );
NOR3_X1 U887 ( .A1(n1037), .A2(n1204), .A3(n1206), .ZN(n1198) );
INV_X1 U888 ( .A(n1199), .ZN(n1206) );
NOR2_X1 U889 ( .A1(n1179), .A2(n1163), .ZN(n1199) );
INV_X1 U890 ( .A(n1219), .ZN(n1163) );
XNOR2_X1 U891 ( .A(G101), .B(n1222), .ZN(G3) );
NAND2_X1 U892 ( .A1(n1223), .A2(n1047), .ZN(n1222) );
XOR2_X1 U893 ( .A(n1224), .B(KEYINPUT34), .Z(n1223) );
NAND2_X1 U894 ( .A1(n1225), .A2(n1036), .ZN(n1224) );
XNOR2_X1 U895 ( .A(n1226), .B(n1227), .ZN(G27) );
NOR2_X1 U896 ( .A1(n1164), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U897 ( .A(KEYINPUT41), .B(n1219), .ZN(n1228) );
NAND2_X1 U898 ( .A1(n1022), .A2(n1229), .ZN(n1219) );
NAND2_X1 U899 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
INV_X1 U900 ( .A(G900), .ZN(n1231) );
NAND3_X1 U901 ( .A1(n1054), .A2(n1051), .A3(n1232), .ZN(n1164) );
XOR2_X1 U902 ( .A(G122), .B(n1174), .Z(G24) );
AND4_X1 U903 ( .A1(n1233), .A2(n1052), .A3(n1234), .A4(n1235), .ZN(n1174) );
NOR2_X1 U904 ( .A1(n1038), .A2(n1064), .ZN(n1052) );
XNOR2_X1 U905 ( .A(G119), .B(n1185), .ZN(G21) );
NAND4_X1 U906 ( .A1(n1208), .A2(n1233), .A3(n1064), .A4(n1038), .ZN(n1185) );
NAND2_X1 U907 ( .A1(n1236), .A2(n1237), .ZN(G18) );
NAND2_X1 U908 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XOR2_X1 U909 ( .A(KEYINPUT33), .B(n1240), .Z(n1236) );
NOR2_X1 U910 ( .A1(n1238), .A2(n1239), .ZN(n1240) );
INV_X1 U911 ( .A(G116), .ZN(n1239) );
INV_X1 U912 ( .A(n1184), .ZN(n1238) );
NAND3_X1 U913 ( .A1(n1233), .A2(n1053), .A3(n1036), .ZN(n1184) );
NOR2_X1 U914 ( .A1(n1235), .A2(n1202), .ZN(n1053) );
XNOR2_X1 U915 ( .A(G113), .B(n1183), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1036), .A2(n1233), .A3(n1054), .ZN(n1183) );
INV_X1 U917 ( .A(n1167), .ZN(n1054) );
NAND2_X1 U918 ( .A1(n1241), .A2(n1235), .ZN(n1167) );
INV_X1 U919 ( .A(n1201), .ZN(n1235) );
AND3_X1 U920 ( .A1(n1047), .A2(n1181), .A3(n1051), .ZN(n1233) );
NOR2_X1 U921 ( .A1(n1044), .A2(n1078), .ZN(n1051) );
NOR2_X1 U922 ( .A1(n1064), .A2(n1204), .ZN(n1036) );
INV_X1 U923 ( .A(n1038), .ZN(n1204) );
XNOR2_X1 U924 ( .A(G110), .B(n1182), .ZN(G12) );
NAND2_X1 U925 ( .A1(n1225), .A2(n1232), .ZN(n1182) );
NOR3_X1 U926 ( .A1(n1038), .A2(n1037), .A3(n1178), .ZN(n1232) );
INV_X1 U927 ( .A(n1047), .ZN(n1178) );
NOR2_X1 U928 ( .A1(n1242), .A2(n1057), .ZN(n1047) );
INV_X1 U929 ( .A(n1049), .ZN(n1057) );
NAND2_X1 U930 ( .A1(G214), .A2(n1243), .ZN(n1049) );
INV_X1 U931 ( .A(n1220), .ZN(n1242) );
XOR2_X1 U932 ( .A(n1244), .B(n1075), .Z(n1220) );
NAND2_X1 U933 ( .A1(G210), .A2(n1243), .ZN(n1075) );
NAND2_X1 U934 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
XNOR2_X1 U935 ( .A(G902), .B(KEYINPUT13), .ZN(n1245) );
XOR2_X1 U936 ( .A(n1071), .B(KEYINPUT8), .Z(n1244) );
NAND2_X1 U937 ( .A1(n1247), .A2(n1248), .ZN(n1071) );
XOR2_X1 U938 ( .A(n1249), .B(n1250), .Z(n1247) );
XOR2_X1 U939 ( .A(n1195), .B(n1251), .Z(n1250) );
NOR2_X1 U940 ( .A1(KEYINPUT54), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U941 ( .A(n1226), .B(n1193), .ZN(n1252) );
XOR2_X1 U942 ( .A(G128), .B(n1253), .Z(n1193) );
INV_X1 U943 ( .A(G125), .ZN(n1226) );
AND2_X1 U944 ( .A1(G224), .A2(n1254), .ZN(n1195) );
NAND2_X1 U945 ( .A1(KEYINPUT47), .A2(n1255), .ZN(n1249) );
XOR2_X1 U946 ( .A(KEYINPUT24), .B(n1189), .Z(n1255) );
XNOR2_X1 U947 ( .A(n1256), .B(n1105), .ZN(n1189) );
XOR2_X1 U948 ( .A(G110), .B(n1257), .Z(n1105) );
XOR2_X1 U949 ( .A(KEYINPUT63), .B(G122), .Z(n1257) );
NAND3_X1 U950 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1256) );
NAND2_X1 U951 ( .A1(KEYINPUT3), .A2(n1261), .ZN(n1260) );
NAND3_X1 U952 ( .A1(n1106), .A2(n1262), .A3(n1263), .ZN(n1259) );
INV_X1 U953 ( .A(n1103), .ZN(n1263) );
NAND2_X1 U954 ( .A1(n1103), .A2(n1264), .ZN(n1258) );
NAND2_X1 U955 ( .A1(n1265), .A2(n1262), .ZN(n1264) );
INV_X1 U956 ( .A(KEYINPUT3), .ZN(n1262) );
XNOR2_X1 U957 ( .A(KEYINPUT62), .B(n1106), .ZN(n1265) );
INV_X1 U958 ( .A(n1261), .ZN(n1106) );
XNOR2_X1 U959 ( .A(n1266), .B(n1267), .ZN(n1261) );
NOR2_X1 U960 ( .A1(KEYINPUT22), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U961 ( .A(G101), .B(KEYINPUT55), .ZN(n1266) );
XNOR2_X1 U962 ( .A(n1269), .B(n1270), .ZN(n1103) );
NAND2_X1 U963 ( .A1(KEYINPUT7), .A2(n1271), .ZN(n1269) );
INV_X1 U964 ( .A(G113), .ZN(n1271) );
INV_X1 U965 ( .A(n1064), .ZN(n1037) );
XNOR2_X1 U966 ( .A(n1272), .B(n1273), .ZN(n1064) );
NOR2_X1 U967 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XNOR2_X1 U968 ( .A(KEYINPUT2), .B(n1112), .ZN(n1275) );
NAND2_X1 U969 ( .A1(n1110), .A2(n1248), .ZN(n1272) );
XNOR2_X1 U970 ( .A(n1276), .B(n1277), .ZN(n1110) );
XOR2_X1 U971 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U972 ( .A(G110), .B(G146), .ZN(n1279) );
NAND3_X1 U973 ( .A1(G234), .A2(n1254), .A3(G221), .ZN(n1278) );
XNOR2_X1 U974 ( .A(n1280), .B(n1281), .ZN(n1276) );
XOR2_X1 U975 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U976 ( .A(n1060), .B(KEYINPUT16), .Z(n1038) );
XNOR2_X1 U977 ( .A(n1284), .B(G472), .ZN(n1060) );
NAND2_X1 U978 ( .A1(n1285), .A2(n1248), .ZN(n1284) );
XOR2_X1 U979 ( .A(n1129), .B(n1286), .Z(n1285) );
XNOR2_X1 U980 ( .A(n1287), .B(n1140), .ZN(n1286) );
NAND2_X1 U981 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U982 ( .A1(n1139), .A2(n1137), .ZN(n1289) );
XOR2_X1 U983 ( .A(n1290), .B(KEYINPUT10), .Z(n1288) );
OR2_X1 U984 ( .A1(n1137), .A2(n1139), .ZN(n1290) );
XNOR2_X1 U985 ( .A(n1270), .B(G113), .ZN(n1139) );
XOR2_X1 U986 ( .A(G116), .B(n1282), .Z(n1270) );
XOR2_X1 U987 ( .A(G119), .B(KEYINPUT53), .Z(n1282) );
XNOR2_X1 U988 ( .A(n1291), .B(n1292), .ZN(n1137) );
XOR2_X1 U989 ( .A(KEYINPUT35), .B(n1253), .Z(n1292) );
XNOR2_X1 U990 ( .A(n1197), .B(n1293), .ZN(n1253) );
NOR2_X1 U991 ( .A1(G143), .A2(KEYINPUT61), .ZN(n1293) );
INV_X1 U992 ( .A(G146), .ZN(n1197) );
NAND3_X1 U993 ( .A1(n1254), .A2(n1246), .A3(G210), .ZN(n1129) );
AND3_X1 U994 ( .A1(n1042), .A2(n1181), .A3(n1208), .ZN(n1225) );
INV_X1 U995 ( .A(n1026), .ZN(n1208) );
NAND2_X1 U996 ( .A1(n1201), .A2(n1241), .ZN(n1026) );
XNOR2_X1 U997 ( .A(n1234), .B(KEYINPUT57), .ZN(n1241) );
INV_X1 U998 ( .A(n1202), .ZN(n1234) );
XOR2_X1 U999 ( .A(n1294), .B(n1063), .Z(n1202) );
INV_X1 U1000 ( .A(G478), .ZN(n1063) );
NAND2_X1 U1001 ( .A1(KEYINPUT32), .A2(n1062), .ZN(n1294) );
INV_X1 U1002 ( .A(n1115), .ZN(n1062) );
NOR2_X1 U1003 ( .A1(n1118), .A2(G902), .ZN(n1115) );
XNOR2_X1 U1004 ( .A(n1295), .B(n1296), .ZN(n1118) );
XNOR2_X1 U1005 ( .A(n1015), .B(n1297), .ZN(n1296) );
NOR3_X1 U1006 ( .A1(n1298), .A2(n1112), .A3(n1299), .ZN(n1297) );
INV_X1 U1007 ( .A(G217), .ZN(n1112) );
XOR2_X1 U1008 ( .A(KEYINPUT43), .B(n1254), .Z(n1298) );
INV_X1 U1009 ( .A(G107), .ZN(n1015) );
XNOR2_X1 U1010 ( .A(n1300), .B(n1301), .ZN(n1295) );
NAND2_X1 U1011 ( .A1(n1302), .A2(KEYINPUT14), .ZN(n1301) );
XNOR2_X1 U1012 ( .A(G116), .B(G122), .ZN(n1302) );
NAND2_X1 U1013 ( .A1(KEYINPUT29), .A2(n1303), .ZN(n1300) );
XNOR2_X1 U1014 ( .A(n1221), .B(n1304), .ZN(n1303) );
XNOR2_X1 U1015 ( .A(n1305), .B(G134), .ZN(n1304) );
XOR2_X1 U1016 ( .A(n1070), .B(n1124), .Z(n1201) );
INV_X1 U1017 ( .A(G475), .ZN(n1124) );
NOR2_X1 U1018 ( .A1(n1123), .A2(G902), .ZN(n1070) );
XNOR2_X1 U1019 ( .A(n1306), .B(n1307), .ZN(n1123) );
XOR2_X1 U1020 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1021 ( .A(n1310), .B(n1311), .ZN(n1309) );
NOR2_X1 U1022 ( .A1(KEYINPUT23), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1023 ( .A(n1313), .B(n1314), .Z(n1312) );
XNOR2_X1 U1024 ( .A(G143), .B(KEYINPUT52), .ZN(n1314) );
NAND3_X1 U1025 ( .A1(n1254), .A2(n1246), .A3(G214), .ZN(n1313) );
INV_X1 U1026 ( .A(G237), .ZN(n1246) );
NAND2_X1 U1027 ( .A1(KEYINPUT36), .A2(G146), .ZN(n1310) );
NOR2_X1 U1028 ( .A1(n1315), .A2(n1316), .ZN(n1308) );
NOR3_X1 U1029 ( .A1(KEYINPUT46), .A2(G125), .A3(n1203), .ZN(n1316) );
NOR2_X1 U1030 ( .A1(n1283), .A2(n1317), .ZN(n1315) );
INV_X1 U1031 ( .A(KEYINPUT46), .ZN(n1317) );
XNOR2_X1 U1032 ( .A(n1203), .B(G125), .ZN(n1283) );
XOR2_X1 U1033 ( .A(n1318), .B(n1319), .Z(n1306) );
XNOR2_X1 U1034 ( .A(n1216), .B(G122), .ZN(n1319) );
XNOR2_X1 U1035 ( .A(G104), .B(G113), .ZN(n1318) );
NAND2_X1 U1036 ( .A1(n1022), .A2(n1320), .ZN(n1181) );
NAND2_X1 U1037 ( .A1(n1230), .A2(n1102), .ZN(n1320) );
INV_X1 U1038 ( .A(G898), .ZN(n1102) );
AND3_X1 U1039 ( .A1(n1321), .A2(n1322), .A3(G953), .ZN(n1230) );
XNOR2_X1 U1040 ( .A(KEYINPUT5), .B(n1248), .ZN(n1321) );
NAND3_X1 U1041 ( .A1(n1322), .A2(n1093), .A3(G952), .ZN(n1022) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1322) );
INV_X1 U1043 ( .A(n1179), .ZN(n1042) );
NAND2_X1 U1044 ( .A1(n1323), .A2(n1044), .ZN(n1179) );
NAND2_X1 U1045 ( .A1(n1079), .A2(n1324), .ZN(n1044) );
NAND2_X1 U1046 ( .A1(G469), .A2(n1325), .ZN(n1324) );
NAND2_X1 U1047 ( .A1(n1326), .A2(n1248), .ZN(n1325) );
NAND3_X1 U1048 ( .A1(n1146), .A2(n1248), .A3(n1326), .ZN(n1079) );
XNOR2_X1 U1049 ( .A(KEYINPUT31), .B(n1149), .ZN(n1326) );
XOR2_X1 U1050 ( .A(n1327), .B(n1328), .Z(n1149) );
XOR2_X1 U1051 ( .A(n1329), .B(n1330), .Z(n1328) );
XNOR2_X1 U1052 ( .A(G110), .B(n1140), .ZN(n1330) );
INV_X1 U1053 ( .A(G101), .ZN(n1140) );
XOR2_X1 U1054 ( .A(KEYINPUT9), .B(KEYINPUT48), .Z(n1329) );
XOR2_X1 U1055 ( .A(n1331), .B(n1332), .Z(n1327) );
XOR2_X1 U1056 ( .A(n1333), .B(n1268), .Z(n1332) );
XNOR2_X1 U1057 ( .A(G104), .B(G107), .ZN(n1268) );
NAND2_X1 U1058 ( .A1(G227), .A2(n1254), .ZN(n1333) );
XNOR2_X1 U1059 ( .A(n1093), .B(KEYINPUT27), .ZN(n1254) );
INV_X1 U1060 ( .A(G953), .ZN(n1093) );
XNOR2_X1 U1061 ( .A(n1291), .B(n1334), .ZN(n1331) );
INV_X1 U1062 ( .A(n1086), .ZN(n1334) );
XOR2_X1 U1063 ( .A(n1335), .B(n1203), .Z(n1086) );
INV_X1 U1064 ( .A(G140), .ZN(n1203) );
NAND2_X1 U1065 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
NAND2_X1 U1066 ( .A1(G146), .A2(n1305), .ZN(n1337) );
XOR2_X1 U1067 ( .A(KEYINPUT49), .B(n1338), .Z(n1336) );
NOR2_X1 U1068 ( .A1(G146), .A2(n1305), .ZN(n1338) );
INV_X1 U1069 ( .A(G143), .ZN(n1305) );
XNOR2_X1 U1070 ( .A(n1087), .B(G134), .ZN(n1291) );
XNOR2_X1 U1071 ( .A(n1216), .B(n1280), .ZN(n1087) );
XNOR2_X1 U1072 ( .A(G137), .B(n1221), .ZN(n1280) );
INV_X1 U1073 ( .A(G128), .ZN(n1221) );
INV_X1 U1074 ( .A(G131), .ZN(n1216) );
INV_X1 U1075 ( .A(G902), .ZN(n1248) );
INV_X1 U1076 ( .A(G469), .ZN(n1146) );
XNOR2_X1 U1077 ( .A(n1078), .B(KEYINPUT19), .ZN(n1323) );
INV_X1 U1078 ( .A(n1043), .ZN(n1078) );
NAND2_X1 U1079 ( .A1(G221), .A2(n1339), .ZN(n1043) );
INV_X1 U1080 ( .A(n1274), .ZN(n1339) );
NOR2_X1 U1081 ( .A1(n1299), .A2(G902), .ZN(n1274) );
INV_X1 U1082 ( .A(G234), .ZN(n1299) );
endmodule


