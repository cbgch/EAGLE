//Key = 0000110000100000011100100011111111000011010111000001101101000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428;

NAND2_X1 U787 ( .A1(n1083), .A2(n1084), .ZN(G9) );
NAND2_X1 U788 ( .A1(G107), .A2(n1085), .ZN(n1084) );
XOR2_X1 U789 ( .A(n1086), .B(KEYINPUT20), .Z(n1083) );
OR2_X1 U790 ( .A1(n1085), .A2(G107), .ZN(n1086) );
NAND3_X1 U791 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
NOR2_X1 U792 ( .A1(n1090), .A2(n1091), .ZN(G75) );
NOR4_X1 U793 ( .A1(G953), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1091) );
NOR2_X1 U794 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NOR2_X1 U795 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NOR2_X1 U796 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
INV_X1 U797 ( .A(n1101), .ZN(n1100) );
NOR2_X1 U798 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
NOR2_X1 U799 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR3_X1 U800 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1104) );
NOR3_X1 U801 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1108) );
XNOR2_X1 U802 ( .A(KEYINPUT31), .B(n1112), .ZN(n1109) );
NOR2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1106) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
NOR3_X1 U806 ( .A1(n1112), .A2(n1119), .A3(n1114), .ZN(n1102) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
AND2_X1 U808 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NOR4_X1 U809 ( .A1(n1124), .A2(n1105), .A3(n1114), .A4(n1112), .ZN(n1097) );
NOR2_X1 U810 ( .A1(n1087), .A2(n1125), .ZN(n1124) );
NOR3_X1 U811 ( .A1(n1092), .A2(G953), .A3(G952), .ZN(n1090) );
AND4_X1 U812 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1092) );
NOR4_X1 U813 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1129) );
NAND3_X1 U814 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1130) );
NAND2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(n1135) );
INV_X1 U817 ( .A(n1141), .ZN(n1140) );
XNOR2_X1 U818 ( .A(KEYINPUT34), .B(n1142), .ZN(n1139) );
NOR3_X1 U819 ( .A1(n1117), .A2(n1143), .A3(n1144), .ZN(n1128) );
XOR2_X1 U820 ( .A(n1145), .B(KEYINPUT44), .Z(n1143) );
XOR2_X1 U821 ( .A(n1146), .B(KEYINPUT6), .Z(n1127) );
XNOR2_X1 U822 ( .A(G472), .B(n1147), .ZN(n1126) );
NOR2_X1 U823 ( .A1(KEYINPUT49), .A2(n1148), .ZN(n1147) );
NAND2_X1 U824 ( .A1(n1149), .A2(n1150), .ZN(G72) );
NAND2_X1 U825 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND2_X1 U826 ( .A1(G953), .A2(n1153), .ZN(n1152) );
NAND2_X1 U827 ( .A1(G900), .A2(G227), .ZN(n1153) );
NAND2_X1 U828 ( .A1(n1154), .A2(n1155), .ZN(n1149) );
INV_X1 U829 ( .A(n1151), .ZN(n1155) );
NOR2_X1 U830 ( .A1(KEYINPUT60), .A2(n1156), .ZN(n1151) );
NOR3_X1 U831 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
NOR2_X1 U832 ( .A1(KEYINPUT54), .A2(n1160), .ZN(n1159) );
NOR3_X1 U833 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1158) );
NOR2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1157) );
NOR2_X1 U835 ( .A1(n1163), .A2(n1166), .ZN(n1165) );
XOR2_X1 U836 ( .A(KEYINPUT7), .B(n1167), .Z(n1166) );
NOR2_X1 U837 ( .A1(n1160), .A2(G953), .ZN(n1167) );
INV_X1 U838 ( .A(KEYINPUT54), .ZN(n1163) );
INV_X1 U839 ( .A(n1162), .ZN(n1164) );
NAND2_X1 U840 ( .A1(n1168), .A2(n1169), .ZN(n1162) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1168) );
XNOR2_X1 U842 ( .A(G125), .B(n1172), .ZN(n1171) );
XNOR2_X1 U843 ( .A(KEYINPUT56), .B(KEYINPUT17), .ZN(n1172) );
XNOR2_X1 U844 ( .A(n1173), .B(n1174), .ZN(n1170) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1173) );
NOR2_X1 U846 ( .A1(G140), .A2(KEYINPUT9), .ZN(n1176) );
NAND2_X1 U847 ( .A1(n1169), .A2(n1177), .ZN(n1154) );
OR2_X1 U848 ( .A1(n1178), .A2(G227), .ZN(n1177) );
INV_X1 U849 ( .A(n1179), .ZN(n1169) );
NAND2_X1 U850 ( .A1(n1180), .A2(n1181), .ZN(G69) );
NAND2_X1 U851 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
OR2_X1 U852 ( .A1(n1178), .A2(G224), .ZN(n1183) );
NAND3_X1 U853 ( .A1(G953), .A2(n1184), .A3(n1185), .ZN(n1180) );
INV_X1 U854 ( .A(n1182), .ZN(n1185) );
XNOR2_X1 U855 ( .A(n1186), .B(n1187), .ZN(n1182) );
NOR2_X1 U856 ( .A1(n1188), .A2(G953), .ZN(n1187) );
NOR3_X1 U857 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1188) );
INV_X1 U858 ( .A(n1192), .ZN(n1190) );
NAND3_X1 U859 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1186) );
NAND2_X1 U860 ( .A1(G953), .A2(n1196), .ZN(n1193) );
NAND2_X1 U861 ( .A1(G898), .A2(G224), .ZN(n1184) );
NOR2_X1 U862 ( .A1(n1197), .A2(n1198), .ZN(G66) );
XOR2_X1 U863 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U864 ( .A1(n1142), .A2(n1201), .ZN(n1199) );
NOR2_X1 U865 ( .A1(n1197), .A2(n1202), .ZN(G63) );
XNOR2_X1 U866 ( .A(n1203), .B(n1204), .ZN(n1202) );
NOR2_X1 U867 ( .A1(n1205), .A2(n1201), .ZN(n1204) );
NOR2_X1 U868 ( .A1(n1197), .A2(n1206), .ZN(G60) );
XOR2_X1 U869 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U870 ( .A1(n1209), .A2(n1201), .ZN(n1207) );
XOR2_X1 U871 ( .A(n1210), .B(n1211), .Z(G6) );
XNOR2_X1 U872 ( .A(G104), .B(KEYINPUT13), .ZN(n1211) );
NAND3_X1 U873 ( .A1(n1089), .A2(n1212), .A3(n1125), .ZN(n1210) );
XNOR2_X1 U874 ( .A(KEYINPUT62), .B(n1105), .ZN(n1212) );
NOR2_X1 U875 ( .A1(n1197), .A2(n1213), .ZN(G57) );
XOR2_X1 U876 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U877 ( .A(n1216), .B(n1217), .Z(n1215) );
NOR2_X1 U878 ( .A1(n1218), .A2(n1201), .ZN(n1217) );
NAND2_X1 U879 ( .A1(KEYINPUT19), .A2(n1219), .ZN(n1216) );
NOR2_X1 U880 ( .A1(n1197), .A2(n1220), .ZN(G54) );
XOR2_X1 U881 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U882 ( .A(n1223), .B(n1224), .ZN(n1222) );
XNOR2_X1 U883 ( .A(n1225), .B(n1226), .ZN(n1224) );
NAND2_X1 U884 ( .A1(KEYINPUT18), .A2(n1227), .ZN(n1226) );
NAND2_X1 U885 ( .A1(KEYINPUT43), .A2(n1228), .ZN(n1225) );
XNOR2_X1 U886 ( .A(n1229), .B(n1230), .ZN(n1228) );
NAND2_X1 U887 ( .A1(KEYINPUT32), .A2(n1231), .ZN(n1229) );
XOR2_X1 U888 ( .A(n1232), .B(n1233), .Z(n1221) );
XNOR2_X1 U889 ( .A(n1234), .B(n1235), .ZN(n1233) );
NOR3_X1 U890 ( .A1(n1201), .A2(KEYINPUT35), .A3(n1236), .ZN(n1232) );
NOR2_X1 U891 ( .A1(n1197), .A2(n1237), .ZN(G51) );
XOR2_X1 U892 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U893 ( .A(n1240), .B(n1241), .Z(n1239) );
NOR2_X1 U894 ( .A1(KEYINPUT47), .A2(n1242), .ZN(n1241) );
NOR2_X1 U895 ( .A1(n1243), .A2(n1201), .ZN(n1240) );
NAND2_X1 U896 ( .A1(G902), .A2(n1094), .ZN(n1201) );
NAND4_X1 U897 ( .A1(n1244), .A2(n1160), .A3(n1245), .A4(n1192), .ZN(n1094) );
INV_X1 U898 ( .A(n1189), .ZN(n1245) );
NAND2_X1 U899 ( .A1(n1246), .A2(n1247), .ZN(n1189) );
NAND2_X1 U900 ( .A1(n1089), .A2(n1248), .ZN(n1247) );
NAND2_X1 U901 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NAND2_X1 U902 ( .A1(n1087), .A2(n1251), .ZN(n1250) );
XNOR2_X1 U903 ( .A(KEYINPUT53), .B(n1105), .ZN(n1251) );
INV_X1 U904 ( .A(n1088), .ZN(n1105) );
NAND2_X1 U905 ( .A1(n1125), .A2(n1088), .ZN(n1249) );
INV_X1 U906 ( .A(n1161), .ZN(n1160) );
NAND4_X1 U907 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1161) );
NOR4_X1 U908 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1255) );
AND2_X1 U909 ( .A1(n1260), .A2(n1261), .ZN(n1254) );
NAND3_X1 U910 ( .A1(n1101), .A2(n1262), .A3(n1263), .ZN(n1252) );
XNOR2_X1 U911 ( .A(KEYINPUT36), .B(n1114), .ZN(n1262) );
XOR2_X1 U912 ( .A(n1191), .B(KEYINPUT30), .Z(n1244) );
NAND4_X1 U913 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1191) );
NAND4_X1 U914 ( .A1(n1268), .A2(n1269), .A3(n1125), .A4(n1270), .ZN(n1264) );
AND2_X1 U915 ( .A1(n1271), .A2(n1121), .ZN(n1270) );
OR2_X1 U916 ( .A1(n1107), .A2(KEYINPUT8), .ZN(n1269) );
NAND2_X1 U917 ( .A1(KEYINPUT8), .A2(n1272), .ZN(n1268) );
OR2_X1 U918 ( .A1(n1112), .A2(n1273), .ZN(n1272) );
XOR2_X1 U919 ( .A(n1274), .B(n1275), .Z(n1238) );
NOR2_X1 U920 ( .A1(n1178), .A2(G952), .ZN(n1197) );
XNOR2_X1 U921 ( .A(G146), .B(n1253), .ZN(G48) );
NAND3_X1 U922 ( .A1(n1125), .A2(n1273), .A3(n1263), .ZN(n1253) );
XNOR2_X1 U923 ( .A(G143), .B(n1261), .ZN(G45) );
NAND4_X1 U924 ( .A1(n1116), .A2(n1273), .A3(n1121), .A4(n1276), .ZN(n1261) );
AND3_X1 U925 ( .A1(n1277), .A2(n1278), .A3(n1279), .ZN(n1276) );
XNOR2_X1 U926 ( .A(G140), .B(n1260), .ZN(G42) );
NAND3_X1 U927 ( .A1(n1280), .A2(n1116), .A3(n1281), .ZN(n1260) );
NAND2_X1 U928 ( .A1(n1282), .A2(n1283), .ZN(G39) );
NAND3_X1 U929 ( .A1(n1280), .A2(n1101), .A3(n1284), .ZN(n1283) );
NOR3_X1 U930 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1284) );
AND2_X1 U931 ( .A1(G137), .A2(KEYINPUT26), .ZN(n1287) );
NOR2_X1 U932 ( .A1(G137), .A2(n1288), .ZN(n1286) );
NAND3_X1 U933 ( .A1(G137), .A2(n1289), .A3(KEYINPUT26), .ZN(n1282) );
NAND4_X1 U934 ( .A1(n1263), .A2(n1280), .A3(n1101), .A4(n1288), .ZN(n1289) );
INV_X1 U935 ( .A(KEYINPUT1), .ZN(n1288) );
XNOR2_X1 U936 ( .A(G134), .B(n1290), .ZN(G36) );
NOR2_X1 U937 ( .A1(n1257), .A2(KEYINPUT59), .ZN(n1290) );
AND3_X1 U938 ( .A1(n1087), .A2(n1279), .A3(n1291), .ZN(n1257) );
XNOR2_X1 U939 ( .A(n1292), .B(n1256), .ZN(G33) );
AND3_X1 U940 ( .A1(n1291), .A2(n1279), .A3(n1125), .ZN(n1256) );
AND3_X1 U941 ( .A1(n1280), .A2(n1116), .A3(n1121), .ZN(n1291) );
INV_X1 U942 ( .A(n1114), .ZN(n1280) );
NAND2_X1 U943 ( .A1(n1293), .A2(n1111), .ZN(n1114) );
XNOR2_X1 U944 ( .A(KEYINPUT58), .B(n1110), .ZN(n1293) );
INV_X1 U945 ( .A(n1294), .ZN(n1110) );
XNOR2_X1 U946 ( .A(n1295), .B(n1259), .ZN(G30) );
AND3_X1 U947 ( .A1(n1087), .A2(n1273), .A3(n1263), .ZN(n1259) );
INV_X1 U948 ( .A(n1285), .ZN(n1263) );
NAND4_X1 U949 ( .A1(n1116), .A2(n1296), .A3(n1279), .A4(n1122), .ZN(n1285) );
XNOR2_X1 U950 ( .A(G101), .B(n1246), .ZN(G3) );
NAND3_X1 U951 ( .A1(n1101), .A2(n1089), .A3(n1121), .ZN(n1246) );
XOR2_X1 U952 ( .A(G125), .B(n1258), .Z(G27) );
AND2_X1 U953 ( .A1(n1107), .A2(n1281), .ZN(n1258) );
AND4_X1 U954 ( .A1(n1123), .A2(n1125), .A3(n1279), .A4(n1122), .ZN(n1281) );
NAND2_X1 U955 ( .A1(n1096), .A2(n1297), .ZN(n1279) );
NAND3_X1 U956 ( .A1(G902), .A2(n1298), .A3(n1179), .ZN(n1297) );
NOR2_X1 U957 ( .A1(n1178), .A2(G900), .ZN(n1179) );
NAND2_X1 U958 ( .A1(n1299), .A2(n1300), .ZN(G24) );
NAND2_X1 U959 ( .A1(G122), .A2(n1265), .ZN(n1300) );
XOR2_X1 U960 ( .A(n1301), .B(KEYINPUT37), .Z(n1299) );
OR2_X1 U961 ( .A1(n1265), .A2(G122), .ZN(n1301) );
NAND4_X1 U962 ( .A1(n1302), .A2(n1088), .A3(n1277), .A4(n1278), .ZN(n1265) );
NOR2_X1 U963 ( .A1(n1122), .A2(n1296), .ZN(n1088) );
XOR2_X1 U964 ( .A(n1266), .B(n1303), .Z(G21) );
NAND2_X1 U965 ( .A1(KEYINPUT51), .A2(G119), .ZN(n1303) );
NAND4_X1 U966 ( .A1(n1302), .A2(n1101), .A3(n1296), .A4(n1122), .ZN(n1266) );
XNOR2_X1 U967 ( .A(G116), .B(n1267), .ZN(G18) );
NAND2_X1 U968 ( .A1(n1304), .A2(n1087), .ZN(n1267) );
NOR2_X1 U969 ( .A1(n1278), .A2(n1305), .ZN(n1087) );
XNOR2_X1 U970 ( .A(G113), .B(n1306), .ZN(G15) );
NAND2_X1 U971 ( .A1(n1304), .A2(n1125), .ZN(n1306) );
AND2_X1 U972 ( .A1(n1307), .A2(n1278), .ZN(n1125) );
XNOR2_X1 U973 ( .A(KEYINPUT33), .B(n1305), .ZN(n1307) );
INV_X1 U974 ( .A(n1277), .ZN(n1305) );
AND2_X1 U975 ( .A1(n1302), .A2(n1121), .ZN(n1304) );
NOR2_X1 U976 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
AND2_X1 U977 ( .A1(n1107), .A2(n1271), .ZN(n1302) );
NOR2_X1 U978 ( .A1(n1112), .A2(n1308), .ZN(n1107) );
INV_X1 U979 ( .A(n1273), .ZN(n1308) );
NAND2_X1 U980 ( .A1(n1309), .A2(n1310), .ZN(n1112) );
XNOR2_X1 U981 ( .A(n1133), .B(KEYINPUT15), .ZN(n1309) );
XNOR2_X1 U982 ( .A(n1192), .B(n1311), .ZN(G12) );
NOR2_X1 U983 ( .A1(KEYINPUT46), .A2(n1234), .ZN(n1311) );
NAND4_X1 U984 ( .A1(n1101), .A2(n1089), .A3(n1123), .A4(n1122), .ZN(n1192) );
NAND2_X1 U985 ( .A1(n1146), .A2(n1312), .ZN(n1122) );
OR2_X1 U986 ( .A1(n1142), .A2(n1141), .ZN(n1312) );
NAND2_X1 U987 ( .A1(n1141), .A2(n1142), .ZN(n1146) );
NAND2_X1 U988 ( .A1(G217), .A2(n1313), .ZN(n1142) );
NOR2_X1 U989 ( .A1(n1200), .A2(G902), .ZN(n1141) );
XNOR2_X1 U990 ( .A(n1314), .B(n1315), .ZN(n1200) );
XNOR2_X1 U991 ( .A(n1316), .B(n1317), .ZN(n1315) );
NAND2_X1 U992 ( .A1(KEYINPUT41), .A2(n1318), .ZN(n1316) );
XOR2_X1 U993 ( .A(n1319), .B(n1320), .Z(n1314) );
NOR2_X1 U994 ( .A1(KEYINPUT14), .A2(n1321), .ZN(n1320) );
XOR2_X1 U995 ( .A(n1322), .B(n1323), .Z(n1321) );
NAND2_X1 U996 ( .A1(KEYINPUT38), .A2(n1324), .ZN(n1323) );
NAND3_X1 U997 ( .A1(G221), .A2(G234), .A3(n1325), .ZN(n1322) );
XNOR2_X1 U998 ( .A(G128), .B(G110), .ZN(n1319) );
INV_X1 U999 ( .A(n1296), .ZN(n1123) );
XOR2_X1 U1000 ( .A(n1148), .B(n1218), .Z(n1296) );
INV_X1 U1001 ( .A(G472), .ZN(n1218) );
NAND2_X1 U1002 ( .A1(n1326), .A2(n1327), .ZN(n1148) );
XNOR2_X1 U1003 ( .A(n1219), .B(n1328), .ZN(n1326) );
XOR2_X1 U1004 ( .A(n1214), .B(KEYINPUT55), .Z(n1328) );
XNOR2_X1 U1005 ( .A(n1329), .B(n1330), .ZN(n1214) );
XNOR2_X1 U1006 ( .A(n1223), .B(n1331), .ZN(n1329) );
AND2_X1 U1007 ( .A1(n1332), .A2(n1333), .ZN(n1219) );
NAND2_X1 U1008 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1009 ( .A1(n1336), .A2(G210), .ZN(n1334) );
NAND3_X1 U1010 ( .A1(n1336), .A2(G210), .A3(G101), .ZN(n1332) );
AND3_X1 U1011 ( .A1(n1273), .A2(n1271), .A3(n1116), .ZN(n1089) );
NOR2_X1 U1012 ( .A1(n1310), .A2(n1133), .ZN(n1116) );
INV_X1 U1013 ( .A(n1118), .ZN(n1133) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1313), .ZN(n1118) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1327), .ZN(n1313) );
INV_X1 U1016 ( .A(n1117), .ZN(n1310) );
XOR2_X1 U1017 ( .A(n1337), .B(n1236), .Z(n1117) );
INV_X1 U1018 ( .A(G469), .ZN(n1236) );
NAND4_X1 U1019 ( .A1(n1338), .A2(n1327), .A3(n1339), .A4(n1340), .ZN(n1337) );
NAND4_X1 U1020 ( .A1(n1341), .A2(n1342), .A3(n1343), .A4(n1344), .ZN(n1340) );
INV_X1 U1021 ( .A(KEYINPUT61), .ZN(n1344) );
NOR2_X1 U1022 ( .A1(KEYINPUT0), .A2(n1345), .ZN(n1343) );
INV_X1 U1023 ( .A(n1346), .ZN(n1345) );
NAND2_X1 U1024 ( .A1(KEYINPUT61), .A2(n1347), .ZN(n1339) );
NAND2_X1 U1025 ( .A1(n1348), .A2(n1349), .ZN(n1338) );
NAND2_X1 U1026 ( .A1(n1341), .A2(n1346), .ZN(n1349) );
NAND2_X1 U1027 ( .A1(n1350), .A2(n1174), .ZN(n1346) );
INV_X1 U1028 ( .A(n1223), .ZN(n1174) );
XNOR2_X1 U1029 ( .A(n1231), .B(n1230), .ZN(n1350) );
XOR2_X1 U1030 ( .A(n1351), .B(KEYINPUT21), .Z(n1341) );
NAND2_X1 U1031 ( .A1(n1352), .A2(n1223), .ZN(n1351) );
XOR2_X1 U1032 ( .A(G131), .B(n1353), .Z(n1223) );
XNOR2_X1 U1033 ( .A(n1324), .B(G134), .ZN(n1353) );
INV_X1 U1034 ( .A(G137), .ZN(n1324) );
XNOR2_X1 U1035 ( .A(n1231), .B(n1354), .ZN(n1352) );
INV_X1 U1036 ( .A(n1230), .ZN(n1354) );
XNOR2_X1 U1037 ( .A(n1355), .B(n1356), .ZN(n1230) );
XNOR2_X1 U1038 ( .A(n1335), .B(n1357), .ZN(n1356) );
NOR2_X1 U1039 ( .A1(G104), .A2(KEYINPUT16), .ZN(n1357) );
INV_X1 U1040 ( .A(G101), .ZN(n1335) );
XNOR2_X1 U1041 ( .A(G107), .B(KEYINPUT2), .ZN(n1355) );
XNOR2_X1 U1042 ( .A(n1175), .B(KEYINPUT39), .ZN(n1231) );
NAND2_X1 U1043 ( .A1(n1358), .A2(n1359), .ZN(n1175) );
NAND2_X1 U1044 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
XOR2_X1 U1045 ( .A(KEYINPUT28), .B(n1362), .Z(n1358) );
NOR2_X1 U1046 ( .A1(n1360), .A2(n1361), .ZN(n1362) );
XNOR2_X1 U1047 ( .A(n1295), .B(KEYINPUT24), .ZN(n1361) );
XNOR2_X1 U1048 ( .A(G143), .B(n1363), .ZN(n1360) );
NOR2_X1 U1049 ( .A1(G146), .A2(KEYINPUT23), .ZN(n1363) );
OR2_X1 U1050 ( .A1(n1347), .A2(KEYINPUT0), .ZN(n1348) );
INV_X1 U1051 ( .A(n1342), .ZN(n1347) );
XNOR2_X1 U1052 ( .A(n1364), .B(n1235), .ZN(n1342) );
AND2_X1 U1053 ( .A1(G227), .A2(n1325), .ZN(n1235) );
XNOR2_X1 U1054 ( .A(G140), .B(G110), .ZN(n1364) );
NAND2_X1 U1055 ( .A1(n1096), .A2(n1365), .ZN(n1271) );
NAND4_X1 U1056 ( .A1(G902), .A2(G953), .A3(n1298), .A4(n1196), .ZN(n1365) );
INV_X1 U1057 ( .A(G898), .ZN(n1196) );
NAND3_X1 U1058 ( .A1(n1298), .A2(n1178), .A3(G952), .ZN(n1096) );
INV_X1 U1059 ( .A(G953), .ZN(n1178) );
NAND2_X1 U1060 ( .A1(G237), .A2(G234), .ZN(n1298) );
NOR2_X1 U1061 ( .A1(n1131), .A2(n1294), .ZN(n1273) );
NOR2_X1 U1062 ( .A1(n1366), .A2(n1132), .ZN(n1294) );
NOR2_X1 U1063 ( .A1(n1138), .A2(n1137), .ZN(n1132) );
AND2_X1 U1064 ( .A1(n1367), .A2(n1137), .ZN(n1366) );
INV_X1 U1065 ( .A(n1243), .ZN(n1137) );
NAND2_X1 U1066 ( .A1(G210), .A2(n1368), .ZN(n1243) );
XOR2_X1 U1067 ( .A(n1138), .B(KEYINPUT42), .Z(n1367) );
NAND3_X1 U1068 ( .A1(n1369), .A2(n1327), .A3(n1370), .ZN(n1138) );
XOR2_X1 U1069 ( .A(KEYINPUT45), .B(n1371), .Z(n1370) );
NOR2_X1 U1070 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
XOR2_X1 U1071 ( .A(KEYINPUT29), .B(n1374), .Z(n1373) );
XOR2_X1 U1072 ( .A(n1274), .B(KEYINPUT22), .Z(n1372) );
OR2_X1 U1073 ( .A1(n1274), .A2(n1374), .ZN(n1369) );
XOR2_X1 U1074 ( .A(n1375), .B(n1275), .Z(n1374) );
NAND2_X1 U1075 ( .A1(G224), .A2(n1325), .ZN(n1275) );
NAND3_X1 U1076 ( .A1(n1376), .A2(n1377), .A3(KEYINPUT52), .ZN(n1375) );
NAND2_X1 U1077 ( .A1(KEYINPUT5), .A2(n1242), .ZN(n1377) );
XNOR2_X1 U1078 ( .A(n1378), .B(G125), .ZN(n1242) );
OR3_X1 U1079 ( .A1(n1330), .A2(G125), .A3(KEYINPUT5), .ZN(n1376) );
INV_X1 U1080 ( .A(n1378), .ZN(n1330) );
XOR2_X1 U1081 ( .A(G146), .B(n1379), .Z(n1378) );
NAND3_X1 U1082 ( .A1(n1380), .A2(n1381), .A3(n1194), .ZN(n1274) );
NAND2_X1 U1083 ( .A1(n1382), .A2(n1383), .ZN(n1194) );
NAND2_X1 U1084 ( .A1(KEYINPUT40), .A2(n1384), .ZN(n1381) );
NAND3_X1 U1085 ( .A1(n1385), .A2(n1386), .A3(n1387), .ZN(n1384) );
INV_X1 U1086 ( .A(n1382), .ZN(n1387) );
NOR2_X1 U1087 ( .A1(n1331), .A2(n1388), .ZN(n1382) );
NAND2_X1 U1088 ( .A1(n1383), .A2(n1389), .ZN(n1386) );
NAND3_X1 U1089 ( .A1(n1390), .A2(n1331), .A3(n1388), .ZN(n1385) );
OR2_X1 U1090 ( .A1(n1195), .A2(KEYINPUT40), .ZN(n1380) );
AND2_X1 U1091 ( .A1(n1391), .A2(n1392), .ZN(n1195) );
NAND3_X1 U1092 ( .A1(n1388), .A2(n1390), .A3(n1393), .ZN(n1392) );
INV_X1 U1093 ( .A(n1331), .ZN(n1393) );
NAND2_X1 U1094 ( .A1(n1394), .A2(n1331), .ZN(n1391) );
XNOR2_X1 U1095 ( .A(n1395), .B(n1396), .ZN(n1331) );
XNOR2_X1 U1096 ( .A(KEYINPUT10), .B(n1318), .ZN(n1396) );
INV_X1 U1097 ( .A(G119), .ZN(n1318) );
XNOR2_X1 U1098 ( .A(G116), .B(G113), .ZN(n1395) );
XNOR2_X1 U1099 ( .A(n1388), .B(n1383), .ZN(n1394) );
INV_X1 U1100 ( .A(n1390), .ZN(n1383) );
XNOR2_X1 U1101 ( .A(n1397), .B(n1398), .ZN(n1390) );
NOR2_X1 U1102 ( .A1(G107), .A2(KEYINPUT50), .ZN(n1398) );
XNOR2_X1 U1103 ( .A(G101), .B(G104), .ZN(n1397) );
INV_X1 U1104 ( .A(n1389), .ZN(n1388) );
NAND2_X1 U1105 ( .A1(n1399), .A2(n1400), .ZN(n1389) );
NAND2_X1 U1106 ( .A1(n1401), .A2(n1234), .ZN(n1400) );
XOR2_X1 U1107 ( .A(KEYINPUT4), .B(n1402), .Z(n1399) );
NOR2_X1 U1108 ( .A1(n1234), .A2(n1401), .ZN(n1402) );
XOR2_X1 U1109 ( .A(KEYINPUT48), .B(G122), .Z(n1401) );
INV_X1 U1110 ( .A(G110), .ZN(n1234) );
INV_X1 U1111 ( .A(n1111), .ZN(n1131) );
NAND2_X1 U1112 ( .A1(G214), .A2(n1368), .ZN(n1111) );
NAND2_X1 U1113 ( .A1(n1403), .A2(n1327), .ZN(n1368) );
NOR2_X1 U1114 ( .A1(n1277), .A2(n1278), .ZN(n1101) );
NAND2_X1 U1115 ( .A1(n1145), .A2(n1134), .ZN(n1278) );
NAND2_X1 U1116 ( .A1(G475), .A2(n1404), .ZN(n1134) );
INV_X1 U1117 ( .A(n1405), .ZN(n1404) );
NAND2_X1 U1118 ( .A1(n1405), .A2(n1209), .ZN(n1145) );
INV_X1 U1119 ( .A(G475), .ZN(n1209) );
NOR2_X1 U1120 ( .A1(n1208), .A2(G902), .ZN(n1405) );
XNOR2_X1 U1121 ( .A(n1406), .B(n1407), .ZN(n1208) );
NOR2_X1 U1122 ( .A1(KEYINPUT12), .A2(n1408), .ZN(n1407) );
XOR2_X1 U1123 ( .A(n1409), .B(n1410), .Z(n1408) );
XNOR2_X1 U1124 ( .A(n1292), .B(n1411), .ZN(n1410) );
NOR2_X1 U1125 ( .A1(G143), .A2(KEYINPUT25), .ZN(n1411) );
INV_X1 U1126 ( .A(G131), .ZN(n1292) );
XNOR2_X1 U1127 ( .A(n1412), .B(n1413), .ZN(n1409) );
INV_X1 U1128 ( .A(n1317), .ZN(n1413) );
XOR2_X1 U1129 ( .A(G125), .B(n1414), .Z(n1317) );
XNOR2_X1 U1130 ( .A(G146), .B(n1227), .ZN(n1414) );
INV_X1 U1131 ( .A(G140), .ZN(n1227) );
NAND2_X1 U1132 ( .A1(n1336), .A2(G214), .ZN(n1412) );
AND2_X1 U1133 ( .A1(n1325), .A2(n1403), .ZN(n1336) );
INV_X1 U1134 ( .A(G237), .ZN(n1403) );
NAND2_X1 U1135 ( .A1(n1415), .A2(n1416), .ZN(n1406) );
NAND2_X1 U1136 ( .A1(G104), .A2(n1417), .ZN(n1416) );
XOR2_X1 U1137 ( .A(KEYINPUT63), .B(n1418), .Z(n1415) );
NOR2_X1 U1138 ( .A1(G104), .A2(n1417), .ZN(n1418) );
XOR2_X1 U1139 ( .A(G122), .B(G113), .Z(n1417) );
XOR2_X1 U1140 ( .A(n1144), .B(KEYINPUT3), .Z(n1277) );
XOR2_X1 U1141 ( .A(n1419), .B(n1205), .Z(n1144) );
INV_X1 U1142 ( .A(G478), .ZN(n1205) );
NAND2_X1 U1143 ( .A1(n1327), .A2(n1203), .ZN(n1419) );
NAND2_X1 U1144 ( .A1(n1420), .A2(n1421), .ZN(n1203) );
NAND2_X1 U1145 ( .A1(n1422), .A2(n1423), .ZN(n1421) );
XOR2_X1 U1146 ( .A(KEYINPUT27), .B(n1424), .Z(n1420) );
NOR2_X1 U1147 ( .A1(n1422), .A2(n1423), .ZN(n1424) );
XOR2_X1 U1148 ( .A(n1425), .B(n1426), .Z(n1423) );
XOR2_X1 U1149 ( .A(G134), .B(G107), .Z(n1426) );
XOR2_X1 U1150 ( .A(n1427), .B(n1379), .Z(n1425) );
XNOR2_X1 U1151 ( .A(n1295), .B(G143), .ZN(n1379) );
INV_X1 U1152 ( .A(G128), .ZN(n1295) );
NAND2_X1 U1153 ( .A1(KEYINPUT57), .A2(n1428), .ZN(n1427) );
XOR2_X1 U1154 ( .A(G122), .B(G116), .Z(n1428) );
AND3_X1 U1155 ( .A1(n1325), .A2(G234), .A3(G217), .ZN(n1422) );
XNOR2_X1 U1156 ( .A(G953), .B(KEYINPUT11), .ZN(n1325) );
INV_X1 U1157 ( .A(G902), .ZN(n1327) );
endmodule


