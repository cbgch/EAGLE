//Key = 0101011000100101111010101000011010110101000000011001010110101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338;

XNOR2_X1 U741 ( .A(G107), .B(n1018), .ZN(G9) );
NOR2_X1 U742 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U743 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1020) );
NOR3_X1 U744 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
NOR2_X1 U745 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U747 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR3_X1 U748 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1032) );
AND3_X1 U749 ( .A1(KEYINPUT49), .A2(n1033), .A3(n1037), .ZN(n1028) );
NAND3_X1 U750 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1033) );
NAND2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
XNOR2_X1 U752 ( .A(KEYINPUT33), .B(n1035), .ZN(n1042) );
OR2_X1 U753 ( .A1(n1043), .A2(KEYINPUT49), .ZN(n1038) );
NOR4_X1 U754 ( .A1(n1044), .A2(n1045), .A3(n1035), .A4(n1031), .ZN(n1023) );
NOR2_X1 U755 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1027), .ZN(n1047) );
NOR2_X1 U757 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U758 ( .A1(n1051), .A2(n1025), .ZN(n1046) );
INV_X1 U759 ( .A(n1052), .ZN(n1025) );
NOR2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NAND3_X1 U761 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1021) );
NAND3_X1 U762 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
XOR2_X1 U763 ( .A(n1061), .B(KEYINPUT58), .Z(n1060) );
NAND4_X1 U764 ( .A1(n1040), .A2(n1062), .A3(n1052), .A4(n1063), .ZN(n1061) );
INV_X1 U765 ( .A(n1031), .ZN(n1040) );
NOR3_X1 U766 ( .A1(n1064), .A2(G953), .A3(G952), .ZN(n1019) );
INV_X1 U767 ( .A(n1055), .ZN(n1064) );
NAND4_X1 U768 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1055) );
NOR4_X1 U769 ( .A1(n1059), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1068) );
XOR2_X1 U770 ( .A(n1072), .B(KEYINPUT53), .Z(n1070) );
NOR2_X1 U771 ( .A1(n1073), .A2(n1074), .ZN(n1069) );
NOR2_X1 U772 ( .A1(n1045), .A2(n1075), .ZN(n1067) );
XNOR2_X1 U773 ( .A(n1076), .B(n1077), .ZN(n1066) );
NOR2_X1 U774 ( .A1(KEYINPUT45), .A2(n1078), .ZN(n1077) );
XOR2_X1 U775 ( .A(n1079), .B(n1080), .Z(n1065) );
NOR2_X1 U776 ( .A1(KEYINPUT19), .A2(n1081), .ZN(n1080) );
XOR2_X1 U777 ( .A(n1082), .B(n1083), .Z(G72) );
NOR2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U779 ( .A1(G227), .A2(n1056), .ZN(n1084) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1082) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U782 ( .A(KEYINPUT27), .B(n1085), .Z(n1089) );
XOR2_X1 U783 ( .A(n1090), .B(n1091), .Z(n1088) );
XNOR2_X1 U784 ( .A(KEYINPUT18), .B(n1092), .ZN(n1091) );
XOR2_X1 U785 ( .A(n1093), .B(n1094), .Z(n1090) );
NAND2_X1 U786 ( .A1(n1056), .A2(n1095), .ZN(n1086) );
XOR2_X1 U787 ( .A(n1096), .B(n1097), .Z(G69) );
XOR2_X1 U788 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U789 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U791 ( .A1(KEYINPUT54), .A2(n1104), .ZN(n1103) );
NOR2_X1 U792 ( .A1(G898), .A2(n1056), .ZN(n1100) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1098) );
XNOR2_X1 U794 ( .A(G953), .B(KEYINPUT10), .ZN(n1106) );
NOR3_X1 U795 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1105) );
XNOR2_X1 U796 ( .A(KEYINPUT63), .B(n1110), .ZN(n1107) );
NOR2_X1 U797 ( .A1(n1111), .A2(n1056), .ZN(n1096) );
AND2_X1 U798 ( .A1(G224), .A2(G898), .ZN(n1111) );
NOR2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(G66) );
NOR3_X1 U800 ( .A1(n1076), .A2(n1114), .A3(n1115), .ZN(n1113) );
NOR3_X1 U801 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
AND2_X1 U802 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NAND3_X1 U803 ( .A1(n1119), .A2(G217), .A3(n1120), .ZN(n1116) );
XOR2_X1 U804 ( .A(n1022), .B(KEYINPUT52), .Z(n1120) );
XOR2_X1 U805 ( .A(n1121), .B(KEYINPUT26), .Z(n1119) );
NOR2_X1 U806 ( .A1(n1112), .A2(n1122), .ZN(G63) );
XNOR2_X1 U807 ( .A(n1123), .B(n1124), .ZN(n1122) );
AND2_X1 U808 ( .A1(G478), .A2(n1125), .ZN(n1124) );
NOR2_X1 U809 ( .A1(n1112), .A2(n1126), .ZN(G60) );
XOR2_X1 U810 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND3_X1 U811 ( .A1(n1125), .A2(n1129), .A3(KEYINPUT34), .ZN(n1127) );
XNOR2_X1 U812 ( .A(KEYINPUT9), .B(n1074), .ZN(n1129) );
XNOR2_X1 U813 ( .A(G104), .B(n1110), .ZN(G6) );
NOR2_X1 U814 ( .A1(n1112), .A2(n1130), .ZN(G57) );
XOR2_X1 U815 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U816 ( .A(n1133), .B(n1134), .ZN(n1132) );
XNOR2_X1 U817 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR3_X1 U818 ( .A1(n1137), .A2(KEYINPUT41), .A3(n1138), .ZN(n1136) );
NAND2_X1 U819 ( .A1(KEYINPUT60), .A2(n1139), .ZN(n1135) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(n1131) );
XNOR2_X1 U821 ( .A(n1142), .B(n1143), .ZN(n1141) );
NAND2_X1 U822 ( .A1(KEYINPUT5), .A2(n1144), .ZN(n1142) );
XNOR2_X1 U823 ( .A(n1145), .B(KEYINPUT35), .ZN(n1140) );
NOR2_X1 U824 ( .A1(n1112), .A2(n1146), .ZN(G54) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U826 ( .A(n1149), .B(n1093), .Z(n1148) );
XNOR2_X1 U827 ( .A(n1133), .B(n1150), .ZN(n1093) );
NAND2_X1 U828 ( .A1(n1151), .A2(KEYINPUT61), .ZN(n1149) );
XNOR2_X1 U829 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR2_X1 U830 ( .A1(KEYINPUT0), .A2(n1154), .ZN(n1153) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1147) );
XNOR2_X1 U832 ( .A(n1157), .B(n1158), .ZN(n1156) );
AND2_X1 U833 ( .A1(G469), .A2(n1125), .ZN(n1155) );
INV_X1 U834 ( .A(n1137), .ZN(n1125) );
NOR2_X1 U835 ( .A1(n1112), .A2(n1159), .ZN(G51) );
XOR2_X1 U836 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U837 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U838 ( .A1(n1079), .A2(n1137), .ZN(n1163) );
NAND2_X1 U839 ( .A1(G902), .A2(n1022), .ZN(n1137) );
OR4_X1 U840 ( .A1(n1164), .A2(n1095), .A3(n1109), .A4(n1165), .ZN(n1022) );
INV_X1 U841 ( .A(n1110), .ZN(n1165) );
NAND3_X1 U842 ( .A1(n1166), .A2(n1052), .A3(n1054), .ZN(n1110) );
NAND2_X1 U843 ( .A1(n1018), .A2(n1167), .ZN(n1109) );
NAND2_X1 U844 ( .A1(n1063), .A2(n1168), .ZN(n1167) );
NAND2_X1 U845 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND4_X1 U846 ( .A1(KEYINPUT40), .A2(n1171), .A3(n1050), .A4(n1172), .ZN(n1170) );
NAND2_X1 U847 ( .A1(n1166), .A2(n1173), .ZN(n1169) );
NAND2_X1 U848 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND2_X1 U849 ( .A1(n1050), .A2(n1176), .ZN(n1175) );
INV_X1 U850 ( .A(KEYINPUT40), .ZN(n1176) );
NAND3_X1 U851 ( .A1(n1053), .A2(n1052), .A3(n1166), .ZN(n1018) );
NAND4_X1 U852 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1095) );
NOR3_X1 U853 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
INV_X1 U854 ( .A(n1184), .ZN(n1181) );
NAND2_X1 U855 ( .A1(n1185), .A2(n1186), .ZN(n1179) );
NAND2_X1 U856 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND3_X1 U857 ( .A1(n1075), .A2(n1189), .A3(n1190), .ZN(n1188) );
NAND2_X1 U858 ( .A1(n1191), .A2(n1053), .ZN(n1187) );
NAND4_X1 U859 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1177) );
NAND2_X1 U860 ( .A1(n1071), .A2(n1196), .ZN(n1195) );
NAND3_X1 U861 ( .A1(n1197), .A2(n1063), .A3(n1191), .ZN(n1196) );
XNOR2_X1 U862 ( .A(KEYINPUT28), .B(n1198), .ZN(n1197) );
NAND2_X1 U863 ( .A1(n1199), .A2(n1200), .ZN(n1194) );
NAND3_X1 U864 ( .A1(n1062), .A2(n1201), .A3(n1054), .ZN(n1200) );
XOR2_X1 U865 ( .A(KEYINPUT12), .B(n1190), .Z(n1201) );
XNOR2_X1 U866 ( .A(n1108), .B(KEYINPUT17), .ZN(n1164) );
NAND4_X1 U867 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1108) );
NOR2_X1 U868 ( .A1(n1206), .A2(n1207), .ZN(n1162) );
XOR2_X1 U869 ( .A(KEYINPUT8), .B(n1208), .Z(n1207) );
NOR2_X1 U870 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XNOR2_X1 U871 ( .A(n1211), .B(KEYINPUT31), .ZN(n1210) );
INV_X1 U872 ( .A(n1212), .ZN(n1209) );
NOR2_X1 U873 ( .A1(n1211), .A2(n1212), .ZN(n1206) );
XNOR2_X1 U874 ( .A(n1213), .B(KEYINPUT30), .ZN(n1212) );
XNOR2_X1 U875 ( .A(n1214), .B(n1215), .ZN(n1211) );
NOR2_X1 U876 ( .A1(n1145), .A2(KEYINPUT46), .ZN(n1215) );
NOR2_X1 U877 ( .A1(n1056), .A2(G952), .ZN(n1112) );
XNOR2_X1 U878 ( .A(G146), .B(n1178), .ZN(G48) );
NAND4_X1 U879 ( .A1(n1216), .A2(n1054), .A3(n1190), .A4(n1041), .ZN(n1178) );
XNOR2_X1 U880 ( .A(G143), .B(n1217), .ZN(G45) );
NAND4_X1 U881 ( .A1(n1218), .A2(KEYINPUT56), .A3(n1219), .A4(n1185), .ZN(n1217) );
NOR2_X1 U882 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XNOR2_X1 U883 ( .A(n1190), .B(KEYINPUT16), .ZN(n1218) );
XNOR2_X1 U884 ( .A(G140), .B(n1184), .ZN(G42) );
NAND4_X1 U885 ( .A1(n1049), .A2(n1191), .A3(n1222), .A4(n1054), .ZN(n1184) );
AND2_X1 U886 ( .A1(n1193), .A2(n1041), .ZN(n1222) );
XNOR2_X1 U887 ( .A(G137), .B(n1223), .ZN(G39) );
NAND4_X1 U888 ( .A1(KEYINPUT32), .A2(n1191), .A3(n1224), .A4(n1216), .ZN(n1223) );
NOR2_X1 U889 ( .A1(n1027), .A2(n1198), .ZN(n1224) );
INV_X1 U890 ( .A(n1063), .ZN(n1027) );
XNOR2_X1 U891 ( .A(G134), .B(n1225), .ZN(G36) );
NAND3_X1 U892 ( .A1(n1053), .A2(n1226), .A3(n1185), .ZN(n1225) );
XNOR2_X1 U893 ( .A(KEYINPUT38), .B(n1035), .ZN(n1226) );
XOR2_X1 U894 ( .A(G131), .B(n1183), .Z(G33) );
AND3_X1 U895 ( .A1(n1191), .A2(n1054), .A3(n1185), .ZN(n1183) );
AND3_X1 U896 ( .A1(n1041), .A2(n1193), .A3(n1050), .ZN(n1185) );
INV_X1 U897 ( .A(n1198), .ZN(n1041) );
INV_X1 U898 ( .A(n1035), .ZN(n1191) );
NAND2_X1 U899 ( .A1(n1058), .A2(n1227), .ZN(n1035) );
NAND2_X1 U900 ( .A1(n1228), .A2(n1229), .ZN(G30) );
NAND2_X1 U901 ( .A1(G128), .A2(n1230), .ZN(n1229) );
XOR2_X1 U902 ( .A(n1231), .B(KEYINPUT2), .Z(n1228) );
NAND2_X1 U903 ( .A1(n1182), .A2(n1232), .ZN(n1231) );
INV_X1 U904 ( .A(n1230), .ZN(n1182) );
NAND3_X1 U905 ( .A1(n1053), .A2(n1172), .A3(n1216), .ZN(n1230) );
AND3_X1 U906 ( .A1(n1192), .A2(n1193), .A3(n1071), .ZN(n1216) );
XNOR2_X1 U907 ( .A(G101), .B(n1233), .ZN(G3) );
NAND4_X1 U908 ( .A1(KEYINPUT48), .A2(n1050), .A3(n1166), .A4(n1063), .ZN(n1233) );
XNOR2_X1 U909 ( .A(G125), .B(n1234), .ZN(G27) );
NAND4_X1 U910 ( .A1(n1037), .A2(n1049), .A3(n1235), .A4(n1193), .ZN(n1234) );
NAND2_X1 U911 ( .A1(n1031), .A2(n1236), .ZN(n1193) );
NAND3_X1 U912 ( .A1(G902), .A2(n1237), .A3(n1085), .ZN(n1236) );
NOR2_X1 U913 ( .A1(G900), .A2(n1056), .ZN(n1085) );
XOR2_X1 U914 ( .A(KEYINPUT62), .B(n1054), .Z(n1235) );
INV_X1 U915 ( .A(n1043), .ZN(n1037) );
XOR2_X1 U916 ( .A(n1202), .B(n1238), .Z(G24) );
NOR2_X1 U917 ( .A1(G122), .A2(KEYINPUT57), .ZN(n1238) );
NAND4_X1 U918 ( .A1(n1239), .A2(n1052), .A3(n1075), .A4(n1189), .ZN(n1202) );
NOR2_X1 U919 ( .A1(n1192), .A2(n1071), .ZN(n1052) );
XNOR2_X1 U920 ( .A(G119), .B(n1203), .ZN(G21) );
NAND4_X1 U921 ( .A1(n1239), .A2(n1063), .A3(n1071), .A4(n1192), .ZN(n1203) );
XNOR2_X1 U922 ( .A(G116), .B(n1204), .ZN(G18) );
NAND3_X1 U923 ( .A1(n1050), .A2(n1053), .A3(n1239), .ZN(n1204) );
AND2_X1 U924 ( .A1(n1240), .A2(n1075), .ZN(n1053) );
XNOR2_X1 U925 ( .A(n1220), .B(KEYINPUT6), .ZN(n1240) );
XNOR2_X1 U926 ( .A(G113), .B(n1205), .ZN(G15) );
NAND3_X1 U927 ( .A1(n1050), .A2(n1054), .A3(n1239), .ZN(n1205) );
NOR2_X1 U928 ( .A1(n1043), .A2(n1171), .ZN(n1239) );
INV_X1 U929 ( .A(n1241), .ZN(n1171) );
NAND2_X1 U930 ( .A1(n1062), .A2(n1190), .ZN(n1043) );
INV_X1 U931 ( .A(n1045), .ZN(n1062) );
NAND2_X1 U932 ( .A1(n1242), .A2(n1034), .ZN(n1045) );
INV_X1 U933 ( .A(n1036), .ZN(n1242) );
NOR2_X1 U934 ( .A1(n1192), .A2(n1199), .ZN(n1050) );
XNOR2_X1 U935 ( .A(G110), .B(n1243), .ZN(G12) );
NAND4_X1 U936 ( .A1(KEYINPUT24), .A2(n1049), .A3(n1166), .A4(n1063), .ZN(n1243) );
NAND2_X1 U937 ( .A1(n1244), .A2(n1245), .ZN(n1063) );
NAND2_X1 U938 ( .A1(n1054), .A2(n1246), .ZN(n1245) );
INV_X1 U939 ( .A(KEYINPUT6), .ZN(n1246) );
NOR2_X1 U940 ( .A1(n1075), .A2(n1220), .ZN(n1054) );
NAND3_X1 U941 ( .A1(n1220), .A2(n1221), .A3(KEYINPUT6), .ZN(n1244) );
INV_X1 U942 ( .A(n1075), .ZN(n1221) );
XNOR2_X1 U943 ( .A(n1247), .B(G478), .ZN(n1075) );
NAND2_X1 U944 ( .A1(n1123), .A2(n1118), .ZN(n1247) );
XNOR2_X1 U945 ( .A(n1248), .B(KEYINPUT4), .ZN(n1123) );
XOR2_X1 U946 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U947 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U948 ( .A(n1232), .B(G122), .ZN(n1252) );
XNOR2_X1 U949 ( .A(KEYINPUT29), .B(n1253), .ZN(n1251) );
INV_X1 U950 ( .A(G143), .ZN(n1253) );
XOR2_X1 U951 ( .A(n1254), .B(n1255), .Z(n1249) );
XOR2_X1 U952 ( .A(n1256), .B(n1257), .Z(n1255) );
NAND2_X1 U953 ( .A1(KEYINPUT39), .A2(n1258), .ZN(n1257) );
INV_X1 U954 ( .A(G134), .ZN(n1258) );
NAND2_X1 U955 ( .A1(G217), .A2(n1259), .ZN(n1256) );
XNOR2_X1 U956 ( .A(G116), .B(G107), .ZN(n1254) );
INV_X1 U957 ( .A(n1189), .ZN(n1220) );
NAND2_X1 U958 ( .A1(n1072), .A2(n1260), .ZN(n1189) );
NAND2_X1 U959 ( .A1(G475), .A2(n1261), .ZN(n1260) );
NAND2_X1 U960 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
INV_X1 U961 ( .A(G475), .ZN(n1074) );
INV_X1 U962 ( .A(n1261), .ZN(n1073) );
NAND2_X1 U963 ( .A1(n1128), .A2(n1118), .ZN(n1261) );
XNOR2_X1 U964 ( .A(n1262), .B(n1263), .ZN(n1128) );
XOR2_X1 U965 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U966 ( .A(G104), .B(n1266), .ZN(n1265) );
NOR2_X1 U967 ( .A1(G140), .A2(KEYINPUT59), .ZN(n1266) );
XNOR2_X1 U968 ( .A(G113), .B(G131), .ZN(n1264) );
XOR2_X1 U969 ( .A(n1267), .B(n1094), .Z(n1262) );
XNOR2_X1 U970 ( .A(n1214), .B(n1268), .ZN(n1094) );
XOR2_X1 U971 ( .A(n1269), .B(n1270), .Z(n1267) );
AND3_X1 U972 ( .A1(G214), .A2(n1056), .A3(n1271), .ZN(n1270) );
NAND2_X1 U973 ( .A1(KEYINPUT47), .A2(G122), .ZN(n1269) );
AND2_X1 U974 ( .A1(n1172), .A2(n1241), .ZN(n1166) );
NAND2_X1 U975 ( .A1(n1031), .A2(n1272), .ZN(n1241) );
NAND4_X1 U976 ( .A1(G953), .A2(G902), .A3(n1237), .A4(n1273), .ZN(n1272) );
INV_X1 U977 ( .A(G898), .ZN(n1273) );
NAND3_X1 U978 ( .A1(n1237), .A2(n1056), .A3(G952), .ZN(n1031) );
NAND2_X1 U979 ( .A1(G234), .A2(n1274), .ZN(n1237) );
XNOR2_X1 U980 ( .A(KEYINPUT11), .B(n1271), .ZN(n1274) );
AND2_X1 U981 ( .A1(n1190), .A2(n1275), .ZN(n1172) );
XNOR2_X1 U982 ( .A(KEYINPUT23), .B(n1198), .ZN(n1275) );
NAND2_X1 U983 ( .A1(n1036), .A2(n1034), .ZN(n1198) );
NAND2_X1 U984 ( .A1(G221), .A2(n1121), .ZN(n1034) );
XNOR2_X1 U985 ( .A(n1276), .B(G469), .ZN(n1036) );
NAND2_X1 U986 ( .A1(n1277), .A2(n1118), .ZN(n1276) );
XOR2_X1 U987 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U988 ( .A(n1152), .B(n1154), .Z(n1279) );
XNOR2_X1 U989 ( .A(n1139), .B(n1280), .ZN(n1154) );
XNOR2_X1 U990 ( .A(G107), .B(n1281), .ZN(n1280) );
INV_X1 U991 ( .A(G104), .ZN(n1281) );
XOR2_X1 U992 ( .A(n1092), .B(n1282), .Z(n1152) );
NAND2_X1 U993 ( .A1(KEYINPUT37), .A2(n1232), .ZN(n1092) );
XOR2_X1 U994 ( .A(n1283), .B(n1133), .Z(n1278) );
NAND2_X1 U995 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U996 ( .A1(n1158), .A2(n1286), .ZN(n1285) );
XOR2_X1 U997 ( .A(n1287), .B(KEYINPUT42), .Z(n1284) );
OR2_X1 U998 ( .A1(n1286), .A2(n1158), .ZN(n1287) );
AND2_X1 U999 ( .A1(G227), .A2(n1056), .ZN(n1158) );
XOR2_X1 U1000 ( .A(n1288), .B(n1157), .Z(n1286) );
NAND2_X1 U1001 ( .A1(KEYINPUT3), .A2(n1150), .ZN(n1288) );
INV_X1 U1002 ( .A(G140), .ZN(n1150) );
NOR2_X1 U1003 ( .A1(n1058), .A2(n1059), .ZN(n1190) );
INV_X1 U1004 ( .A(n1227), .ZN(n1059) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1289), .ZN(n1227) );
XNOR2_X1 U1006 ( .A(n1081), .B(n1079), .ZN(n1058) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1289), .ZN(n1079) );
NAND2_X1 U1008 ( .A1(n1290), .A2(n1271), .ZN(n1289) );
NAND2_X1 U1009 ( .A1(n1291), .A2(n1118), .ZN(n1081) );
XNOR2_X1 U1010 ( .A(n1160), .B(n1292), .ZN(n1291) );
XOR2_X1 U1011 ( .A(n1213), .B(n1293), .Z(n1292) );
NAND2_X1 U1012 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NAND2_X1 U1013 ( .A1(n1214), .A2(n1296), .ZN(n1295) );
XOR2_X1 U1014 ( .A(KEYINPUT13), .B(n1297), .Z(n1294) );
NOR2_X1 U1015 ( .A1(n1214), .A2(n1296), .ZN(n1297) );
NAND2_X1 U1016 ( .A1(n1298), .A2(G224), .ZN(n1213) );
XNOR2_X1 U1017 ( .A(G953), .B(KEYINPUT21), .ZN(n1298) );
XNOR2_X1 U1018 ( .A(n1102), .B(n1299), .ZN(n1160) );
NOR2_X1 U1019 ( .A1(KEYINPUT36), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U1020 ( .A(n1104), .B(KEYINPUT14), .ZN(n1300) );
XOR2_X1 U1021 ( .A(G110), .B(G122), .Z(n1104) );
XNOR2_X1 U1022 ( .A(n1301), .B(n1144), .ZN(n1102) );
XNOR2_X1 U1023 ( .A(n1302), .B(n1139), .ZN(n1301) );
INV_X1 U1024 ( .A(G101), .ZN(n1139) );
NAND2_X1 U1025 ( .A1(n1303), .A2(KEYINPUT1), .ZN(n1302) );
XNOR2_X1 U1026 ( .A(G107), .B(n1304), .ZN(n1303) );
NOR2_X1 U1027 ( .A1(G104), .A2(KEYINPUT43), .ZN(n1304) );
INV_X1 U1028 ( .A(n1174), .ZN(n1049) );
NAND2_X1 U1029 ( .A1(n1199), .A2(n1192), .ZN(n1174) );
XNOR2_X1 U1030 ( .A(n1076), .B(n1078), .ZN(n1192) );
NAND2_X1 U1031 ( .A1(G217), .A2(n1121), .ZN(n1078) );
NAND2_X1 U1032 ( .A1(G234), .A2(n1290), .ZN(n1121) );
XNOR2_X1 U1033 ( .A(n1118), .B(KEYINPUT20), .ZN(n1290) );
AND2_X1 U1034 ( .A1(n1117), .A2(n1118), .ZN(n1076) );
XOR2_X1 U1035 ( .A(n1305), .B(n1306), .Z(n1117) );
XOR2_X1 U1036 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1037 ( .A(n1309), .B(n1157), .ZN(n1308) );
INV_X1 U1038 ( .A(G110), .ZN(n1157) );
NAND2_X1 U1039 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND2_X1 U1040 ( .A1(G119), .A2(n1232), .ZN(n1311) );
XOR2_X1 U1041 ( .A(n1312), .B(KEYINPUT7), .Z(n1310) );
NAND2_X1 U1042 ( .A1(G128), .A2(n1313), .ZN(n1312) );
XNOR2_X1 U1043 ( .A(G137), .B(G140), .ZN(n1307) );
XOR2_X1 U1044 ( .A(n1214), .B(n1314), .Z(n1305) );
XOR2_X1 U1045 ( .A(n1315), .B(n1316), .Z(n1314) );
NAND2_X1 U1046 ( .A1(KEYINPUT51), .A2(n1317), .ZN(n1316) );
NAND2_X1 U1047 ( .A1(n1259), .A2(G221), .ZN(n1315) );
AND2_X1 U1048 ( .A1(G234), .A2(n1056), .ZN(n1259) );
XNOR2_X1 U1049 ( .A(G125), .B(KEYINPUT55), .ZN(n1214) );
INV_X1 U1050 ( .A(n1071), .ZN(n1199) );
XOR2_X1 U1051 ( .A(n1318), .B(n1138), .Z(n1071) );
INV_X1 U1052 ( .A(G472), .ZN(n1138) );
NAND4_X1 U1053 ( .A1(n1319), .A2(n1118), .A3(n1320), .A4(n1321), .ZN(n1318) );
OR2_X1 U1054 ( .A1(n1322), .A2(KEYINPUT15), .ZN(n1321) );
NAND4_X1 U1055 ( .A1(n1323), .A2(n1324), .A3(n1322), .A4(KEYINPUT15), .ZN(n1320) );
XNOR2_X1 U1056 ( .A(n1325), .B(n1326), .ZN(n1323) );
INV_X1 U1057 ( .A(G902), .ZN(n1118) );
NAND2_X1 U1058 ( .A1(n1327), .A2(n1328), .ZN(n1319) );
NAND2_X1 U1059 ( .A1(n1322), .A2(n1324), .ZN(n1328) );
INV_X1 U1060 ( .A(KEYINPUT50), .ZN(n1324) );
XNOR2_X1 U1061 ( .A(n1143), .B(G101), .ZN(n1322) );
NAND3_X1 U1062 ( .A1(n1271), .A2(n1056), .A3(G210), .ZN(n1143) );
INV_X1 U1063 ( .A(G953), .ZN(n1056) );
INV_X1 U1064 ( .A(G237), .ZN(n1271) );
XNOR2_X1 U1065 ( .A(n1326), .B(n1144), .ZN(n1327) );
INV_X1 U1066 ( .A(n1325), .ZN(n1144) );
XOR2_X1 U1067 ( .A(G113), .B(n1329), .Z(n1325) );
XNOR2_X1 U1068 ( .A(n1313), .B(G116), .ZN(n1329) );
INV_X1 U1069 ( .A(G119), .ZN(n1313) );
XNOR2_X1 U1070 ( .A(n1330), .B(n1145), .ZN(n1326) );
INV_X1 U1071 ( .A(n1296), .ZN(n1145) );
NAND3_X1 U1072 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1296) );
NAND2_X1 U1073 ( .A1(KEYINPUT44), .A2(n1232), .ZN(n1333) );
NAND3_X1 U1074 ( .A1(G128), .A2(n1334), .A3(n1268), .ZN(n1332) );
NAND2_X1 U1075 ( .A1(n1282), .A2(n1335), .ZN(n1331) );
NAND2_X1 U1076 ( .A1(n1336), .A2(n1334), .ZN(n1335) );
INV_X1 U1077 ( .A(KEYINPUT44), .ZN(n1334) );
XNOR2_X1 U1078 ( .A(KEYINPUT25), .B(n1232), .ZN(n1336) );
INV_X1 U1079 ( .A(G128), .ZN(n1232) );
INV_X1 U1080 ( .A(n1268), .ZN(n1282) );
XNOR2_X1 U1081 ( .A(G143), .B(n1317), .ZN(n1268) );
INV_X1 U1082 ( .A(G146), .ZN(n1317) );
NAND2_X1 U1083 ( .A1(KEYINPUT22), .A2(n1133), .ZN(n1330) );
XNOR2_X1 U1084 ( .A(G131), .B(n1337), .ZN(n1133) );
XNOR2_X1 U1085 ( .A(n1338), .B(G134), .ZN(n1337) );
INV_X1 U1086 ( .A(G137), .ZN(n1338) );
endmodule


