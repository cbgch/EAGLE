//Key = 1101101100110110101100111100001010101110101011010100111001011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366;

XOR2_X1 U739 ( .A(G107), .B(n1024), .Z(G9) );
NOR2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR4_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
NOR2_X1 U742 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR3_X1 U745 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1033) );
XOR2_X1 U746 ( .A(n1036), .B(KEYINPUT46), .Z(n1039) );
NAND3_X1 U747 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1027) );
NAND3_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NAND3_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1044) );
NAND2_X1 U750 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
OR2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
INV_X1 U752 ( .A(n1032), .ZN(n1049) );
NAND3_X1 U753 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1032) );
NAND3_X1 U754 ( .A1(n1056), .A2(n1057), .A3(n1055), .ZN(n1047) );
NAND3_X1 U755 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NAND2_X1 U756 ( .A1(n1053), .A2(n1061), .ZN(n1060) );
NAND2_X1 U757 ( .A1(n1054), .A2(n1062), .ZN(n1059) );
NAND2_X1 U758 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U759 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
INV_X1 U760 ( .A(n1067), .ZN(n1063) );
NAND2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1058) );
INV_X1 U762 ( .A(KEYINPUT33), .ZN(n1069) );
NAND2_X1 U763 ( .A1(KEYINPUT33), .A2(n1070), .ZN(n1046) );
NAND3_X1 U764 ( .A1(n1068), .A2(n1056), .A3(n1055), .ZN(n1070) );
INV_X1 U765 ( .A(n1071), .ZN(n1055) );
NOR3_X1 U766 ( .A1(n1072), .A2(G953), .A3(G952), .ZN(n1025) );
INV_X1 U767 ( .A(n1040), .ZN(n1072) );
NAND4_X1 U768 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1040) );
NOR4_X1 U769 ( .A1(n1077), .A2(n1078), .A3(n1065), .A4(n1079), .ZN(n1076) );
NOR2_X1 U770 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
INV_X1 U771 ( .A(n1082), .ZN(n1077) );
NOR2_X1 U772 ( .A1(n1036), .A2(n1083), .ZN(n1075) );
XOR2_X1 U773 ( .A(n1084), .B(n1085), .Z(n1074) );
XNOR2_X1 U774 ( .A(G469), .B(KEYINPUT22), .ZN(n1085) );
XOR2_X1 U775 ( .A(n1086), .B(n1087), .Z(n1073) );
XOR2_X1 U776 ( .A(n1088), .B(KEYINPUT38), .Z(n1087) );
XOR2_X1 U777 ( .A(n1089), .B(n1090), .Z(G72) );
XOR2_X1 U778 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U779 ( .A1(G953), .A2(n1093), .ZN(n1092) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U783 ( .A1(KEYINPUT48), .A2(n1098), .ZN(n1096) );
XOR2_X1 U784 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U785 ( .A1(KEYINPUT43), .A2(n1101), .ZN(n1100) );
XOR2_X1 U786 ( .A(KEYINPUT42), .B(n1102), .Z(n1101) );
NOR3_X1 U787 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1099) );
NOR2_X1 U788 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR3_X1 U789 ( .A1(G131), .A2(n1108), .A3(n1109), .ZN(n1104) );
INV_X1 U790 ( .A(n1107), .ZN(n1109) );
NAND2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
XNOR2_X1 U792 ( .A(G134), .B(KEYINPUT16), .ZN(n1110) );
INV_X1 U793 ( .A(n1112), .ZN(n1103) );
XOR2_X1 U794 ( .A(n1113), .B(KEYINPUT62), .Z(n1094) );
NAND2_X1 U795 ( .A1(G953), .A2(n1114), .ZN(n1113) );
NOR2_X1 U796 ( .A1(n1115), .A2(G953), .ZN(n1089) );
NAND2_X1 U797 ( .A1(n1116), .A2(n1117), .ZN(G69) );
NAND2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U799 ( .A1(G953), .A2(n1120), .ZN(n1119) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1120) );
INV_X1 U801 ( .A(n1121), .ZN(n1118) );
NAND2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U804 ( .A1(G953), .A2(n1125), .ZN(n1124) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1121) );
NOR2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U807 ( .A(n1041), .B(KEYINPUT61), .Z(n1129) );
NAND4_X1 U808 ( .A1(n1130), .A2(n1123), .A3(n1131), .A4(n1132), .ZN(n1126) );
OR3_X1 U809 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
NAND2_X1 U810 ( .A1(n1136), .A2(n1135), .ZN(n1131) );
XOR2_X1 U811 ( .A(n1134), .B(n1137), .Z(n1136) );
XNOR2_X1 U812 ( .A(KEYINPUT6), .B(n1133), .ZN(n1137) );
INV_X1 U813 ( .A(n1138), .ZN(n1123) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U815 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U816 ( .A1(n1081), .A2(n1143), .ZN(n1141) );
NOR2_X1 U817 ( .A1(n1139), .A2(n1144), .ZN(G63) );
XOR2_X1 U818 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND3_X1 U819 ( .A1(n1147), .A2(G478), .A3(KEYINPUT36), .ZN(n1145) );
NOR2_X1 U820 ( .A1(n1139), .A2(n1148), .ZN(G60) );
XNOR2_X1 U821 ( .A(n1149), .B(n1150), .ZN(n1148) );
AND2_X1 U822 ( .A1(G475), .A2(n1147), .ZN(n1150) );
NAND2_X1 U823 ( .A1(n1151), .A2(n1152), .ZN(G6) );
OR2_X1 U824 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U825 ( .A(n1155), .B(KEYINPUT20), .Z(n1151) );
NAND2_X1 U826 ( .A1(n1154), .A2(n1153), .ZN(n1155) );
XOR2_X1 U827 ( .A(G104), .B(KEYINPUT5), .Z(n1154) );
NOR2_X1 U828 ( .A1(n1139), .A2(n1156), .ZN(G57) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U830 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U831 ( .A1(G472), .A2(n1147), .ZN(n1159) );
INV_X1 U832 ( .A(n1143), .ZN(n1147) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1157) );
NAND2_X1 U834 ( .A1(KEYINPUT60), .A2(n1163), .ZN(n1162) );
NAND2_X1 U835 ( .A1(n1164), .A2(KEYINPUT11), .ZN(n1161) );
XOR2_X1 U836 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U837 ( .A1(n1139), .A2(n1167), .ZN(G54) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
XNOR2_X1 U839 ( .A(n1170), .B(n1171), .ZN(n1169) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1168) );
XOR2_X1 U841 ( .A(KEYINPUT57), .B(n1174), .Z(n1173) );
NAND3_X1 U842 ( .A1(G469), .A2(n1175), .A3(n1176), .ZN(n1172) );
XOR2_X1 U843 ( .A(n1177), .B(KEYINPUT14), .Z(n1176) );
NOR2_X1 U844 ( .A1(n1139), .A2(n1178), .ZN(G51) );
XOR2_X1 U845 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U846 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U847 ( .A1(n1086), .A2(n1143), .ZN(n1181) );
NAND2_X1 U848 ( .A1(G902), .A2(n1175), .ZN(n1143) );
NAND2_X1 U849 ( .A1(n1115), .A2(n1128), .ZN(n1175) );
INV_X1 U850 ( .A(n1030), .ZN(n1128) );
NAND4_X1 U851 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1030) );
NOR4_X1 U852 ( .A1(n1187), .A2(n1188), .A3(n1024), .A4(n1189), .ZN(n1186) );
INV_X1 U853 ( .A(n1153), .ZN(n1189) );
NAND3_X1 U854 ( .A1(n1190), .A2(n1054), .A3(n1051), .ZN(n1153) );
AND3_X1 U855 ( .A1(n1054), .A2(n1052), .A3(n1190), .ZN(n1024) );
NAND2_X1 U856 ( .A1(KEYINPUT37), .A2(n1191), .ZN(n1185) );
NAND3_X1 U857 ( .A1(n1192), .A2(n1193), .A3(n1053), .ZN(n1183) );
NAND3_X1 U858 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1193) );
NAND2_X1 U859 ( .A1(n1051), .A2(n1061), .ZN(n1196) );
NAND3_X1 U860 ( .A1(n1197), .A2(n1198), .A3(n1054), .ZN(n1195) );
INV_X1 U861 ( .A(KEYINPUT37), .ZN(n1198) );
NAND2_X1 U862 ( .A1(n1199), .A2(n1056), .ZN(n1194) );
INV_X1 U863 ( .A(n1028), .ZN(n1115) );
NAND4_X1 U864 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1028) );
NOR4_X1 U865 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
NAND2_X1 U866 ( .A1(n1051), .A2(n1208), .ZN(n1202) );
NAND2_X1 U867 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND3_X1 U868 ( .A1(n1199), .A2(n1211), .A3(n1067), .ZN(n1210) );
NAND2_X1 U869 ( .A1(n1212), .A2(n1213), .ZN(n1209) );
XOR2_X1 U870 ( .A(KEYINPUT27), .B(n1214), .Z(n1213) );
NOR2_X1 U871 ( .A1(n1041), .A2(G952), .ZN(n1139) );
XOR2_X1 U872 ( .A(n1215), .B(n1216), .Z(G48) );
XOR2_X1 U873 ( .A(n1217), .B(KEYINPUT26), .Z(n1216) );
NAND4_X1 U874 ( .A1(n1067), .A2(KEYINPUT18), .A3(n1218), .A4(n1199), .ZN(n1215) );
NOR2_X1 U875 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XNOR2_X1 U876 ( .A(G143), .B(n1200), .ZN(G45) );
NAND4_X1 U877 ( .A1(n1067), .A2(n1221), .A3(n1211), .A4(n1061), .ZN(n1200) );
XOR2_X1 U878 ( .A(G140), .B(n1222), .Z(G42) );
NOR3_X1 U879 ( .A1(n1223), .A2(n1224), .A3(n1219), .ZN(n1222) );
XOR2_X1 U880 ( .A(n1111), .B(n1201), .Z(G39) );
NAND3_X1 U881 ( .A1(n1199), .A2(n1056), .A3(n1212), .ZN(n1201) );
XOR2_X1 U882 ( .A(G134), .B(n1207), .Z(G36) );
AND3_X1 U883 ( .A1(n1052), .A2(n1061), .A3(n1212), .ZN(n1207) );
INV_X1 U884 ( .A(n1223), .ZN(n1212) );
XOR2_X1 U885 ( .A(G131), .B(n1206), .Z(G33) );
NOR3_X1 U886 ( .A1(n1219), .A2(n1225), .A3(n1223), .ZN(n1206) );
NAND4_X1 U887 ( .A1(n1067), .A2(n1045), .A3(n1043), .A4(n1226), .ZN(n1223) );
INV_X1 U888 ( .A(n1038), .ZN(n1043) );
XOR2_X1 U889 ( .A(n1078), .B(KEYINPUT52), .Z(n1045) );
INV_X1 U890 ( .A(n1037), .ZN(n1078) );
XNOR2_X1 U891 ( .A(n1227), .B(KEYINPUT24), .ZN(n1067) );
XOR2_X1 U892 ( .A(G128), .B(n1205), .Z(G30) );
AND4_X1 U893 ( .A1(n1199), .A2(n1211), .A3(n1052), .A4(n1227), .ZN(n1205) );
XOR2_X1 U894 ( .A(n1163), .B(n1228), .Z(G3) );
NOR2_X1 U895 ( .A1(n1188), .A2(KEYINPUT35), .ZN(n1228) );
AND3_X1 U896 ( .A1(n1190), .A2(n1061), .A3(n1056), .ZN(n1188) );
INV_X1 U897 ( .A(G101), .ZN(n1163) );
XOR2_X1 U898 ( .A(G125), .B(n1204), .Z(G27) );
AND3_X1 U899 ( .A1(n1068), .A2(n1051), .A3(n1211), .ZN(n1204) );
INV_X1 U900 ( .A(n1220), .ZN(n1211) );
NAND2_X1 U901 ( .A1(n1229), .A2(n1226), .ZN(n1220) );
NAND2_X1 U902 ( .A1(n1071), .A2(n1230), .ZN(n1226) );
NAND4_X1 U903 ( .A1(G953), .A2(G902), .A3(n1231), .A4(n1114), .ZN(n1230) );
INV_X1 U904 ( .A(G900), .ZN(n1114) );
NOR2_X1 U905 ( .A1(n1224), .A2(n1232), .ZN(n1068) );
INV_X1 U906 ( .A(n1214), .ZN(n1224) );
NAND2_X1 U907 ( .A1(n1233), .A2(n1234), .ZN(G24) );
NAND2_X1 U908 ( .A1(n1191), .A2(n1235), .ZN(n1234) );
INV_X1 U909 ( .A(n1236), .ZN(n1191) );
XOR2_X1 U910 ( .A(n1237), .B(KEYINPUT58), .Z(n1233) );
NAND2_X1 U911 ( .A1(G122), .A2(n1236), .ZN(n1237) );
NAND4_X1 U912 ( .A1(n1221), .A2(n1053), .A3(n1054), .A4(n1192), .ZN(n1236) );
INV_X1 U913 ( .A(n1197), .ZN(n1221) );
NAND2_X1 U914 ( .A1(n1238), .A2(n1239), .ZN(n1197) );
XOR2_X1 U915 ( .A(n1240), .B(n1241), .Z(G21) );
XNOR2_X1 U916 ( .A(G119), .B(KEYINPUT56), .ZN(n1241) );
NAND3_X1 U917 ( .A1(n1242), .A2(n1199), .A3(n1243), .ZN(n1240) );
NOR3_X1 U918 ( .A1(n1232), .A2(n1244), .A3(n1036), .ZN(n1243) );
INV_X1 U919 ( .A(n1056), .ZN(n1036) );
AND2_X1 U920 ( .A1(n1071), .A2(n1245), .ZN(n1244) );
AND2_X1 U921 ( .A1(n1083), .A2(n1246), .ZN(n1199) );
XOR2_X1 U922 ( .A(n1035), .B(KEYINPUT49), .Z(n1242) );
XOR2_X1 U923 ( .A(n1187), .B(n1247), .Z(G18) );
NOR2_X1 U924 ( .A1(KEYINPUT15), .A2(n1248), .ZN(n1247) );
INV_X1 U925 ( .A(G116), .ZN(n1248) );
AND4_X1 U926 ( .A1(n1053), .A2(n1052), .A3(n1192), .A4(n1061), .ZN(n1187) );
NOR2_X1 U927 ( .A1(n1238), .A2(n1249), .ZN(n1052) );
XOR2_X1 U928 ( .A(n1250), .B(n1251), .Z(G15) );
NAND3_X1 U929 ( .A1(KEYINPUT47), .A2(n1051), .A3(n1252), .ZN(n1251) );
NOR3_X1 U930 ( .A1(n1253), .A2(n1225), .A3(n1254), .ZN(n1252) );
XOR2_X1 U931 ( .A(n1232), .B(KEYINPUT28), .Z(n1254) );
INV_X1 U932 ( .A(n1053), .ZN(n1232) );
NOR2_X1 U933 ( .A1(n1255), .A2(n1065), .ZN(n1053) );
INV_X1 U934 ( .A(n1061), .ZN(n1225) );
NAND2_X1 U935 ( .A1(n1256), .A2(n1257), .ZN(n1061) );
NAND2_X1 U936 ( .A1(n1054), .A2(n1258), .ZN(n1257) );
INV_X1 U937 ( .A(KEYINPUT3), .ZN(n1258) );
NOR2_X1 U938 ( .A1(n1246), .A2(n1083), .ZN(n1054) );
NAND3_X1 U939 ( .A1(n1259), .A2(n1083), .A3(KEYINPUT3), .ZN(n1256) );
INV_X1 U940 ( .A(n1219), .ZN(n1051) );
NAND2_X1 U941 ( .A1(n1249), .A2(n1238), .ZN(n1219) );
XNOR2_X1 U942 ( .A(G110), .B(n1184), .ZN(G12) );
NAND3_X1 U943 ( .A1(n1056), .A2(n1190), .A3(n1214), .ZN(n1184) );
NOR2_X1 U944 ( .A1(n1083), .A2(n1259), .ZN(n1214) );
INV_X1 U945 ( .A(n1246), .ZN(n1259) );
NAND3_X1 U946 ( .A1(n1260), .A2(n1261), .A3(n1082), .ZN(n1246) );
NAND2_X1 U947 ( .A1(n1080), .A2(n1081), .ZN(n1082) );
NAND2_X1 U948 ( .A1(n1081), .A2(n1262), .ZN(n1261) );
OR3_X1 U949 ( .A1(n1081), .A2(n1080), .A3(n1262), .ZN(n1260) );
INV_X1 U950 ( .A(KEYINPUT53), .ZN(n1262) );
NOR2_X1 U951 ( .A1(n1142), .A2(G902), .ZN(n1080) );
XNOR2_X1 U952 ( .A(n1263), .B(n1264), .ZN(n1142) );
XOR2_X1 U953 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U954 ( .A(G119), .B(G110), .Z(n1266) );
XOR2_X1 U955 ( .A(KEYINPUT25), .B(G128), .Z(n1265) );
XOR2_X1 U956 ( .A(n1267), .B(n1268), .Z(n1263) );
XOR2_X1 U957 ( .A(n1269), .B(n1270), .Z(n1268) );
NAND3_X1 U958 ( .A1(G234), .A2(n1041), .A3(G221), .ZN(n1270) );
NAND2_X1 U959 ( .A1(KEYINPUT0), .A2(n1111), .ZN(n1269) );
XNOR2_X1 U960 ( .A(n1271), .B(n1272), .ZN(n1267) );
NAND2_X1 U961 ( .A1(G217), .A2(n1273), .ZN(n1081) );
XNOR2_X1 U962 ( .A(n1274), .B(G472), .ZN(n1083) );
NAND2_X1 U963 ( .A1(n1275), .A2(n1177), .ZN(n1274) );
XOR2_X1 U964 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U965 ( .A(n1278), .B(n1160), .ZN(n1277) );
XNOR2_X1 U966 ( .A(n1279), .B(n1280), .ZN(n1160) );
XOR2_X1 U967 ( .A(n1281), .B(G113), .Z(n1279) );
NAND2_X1 U968 ( .A1(n1282), .A2(G210), .ZN(n1281) );
NAND3_X1 U969 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1278) );
NAND2_X1 U970 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U971 ( .A1(n1288), .A2(n1289), .ZN(n1284) );
INV_X1 U972 ( .A(KEYINPUT19), .ZN(n1289) );
NAND2_X1 U973 ( .A1(n1166), .A2(n1290), .ZN(n1288) );
XOR2_X1 U974 ( .A(KEYINPUT17), .B(n1165), .Z(n1290) );
INV_X1 U975 ( .A(n1287), .ZN(n1165) );
INV_X1 U976 ( .A(n1286), .ZN(n1166) );
NAND2_X1 U977 ( .A1(KEYINPUT19), .A2(n1291), .ZN(n1283) );
NAND2_X1 U978 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
OR3_X1 U979 ( .A1(n1287), .A2(n1286), .A3(KEYINPUT17), .ZN(n1293) );
NAND2_X1 U980 ( .A1(KEYINPUT17), .A2(n1287), .ZN(n1292) );
XOR2_X1 U981 ( .A(KEYINPUT9), .B(G101), .Z(n1276) );
AND2_X1 U982 ( .A1(n1192), .A2(n1227), .ZN(n1190) );
NOR2_X1 U983 ( .A1(n1065), .A2(n1066), .ZN(n1227) );
INV_X1 U984 ( .A(n1255), .ZN(n1066) );
NAND2_X1 U985 ( .A1(n1294), .A2(n1295), .ZN(n1255) );
NAND2_X1 U986 ( .A1(G469), .A2(n1084), .ZN(n1295) );
XOR2_X1 U987 ( .A(KEYINPUT7), .B(n1296), .Z(n1294) );
NOR2_X1 U988 ( .A1(G469), .A2(n1084), .ZN(n1296) );
NAND2_X1 U989 ( .A1(n1297), .A2(n1177), .ZN(n1084) );
XOR2_X1 U990 ( .A(n1170), .B(n1298), .Z(n1297) );
NOR2_X1 U991 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NOR3_X1 U992 ( .A1(n1174), .A2(n1171), .A3(n1301), .ZN(n1300) );
INV_X1 U993 ( .A(n1302), .ZN(n1174) );
NOR2_X1 U994 ( .A1(n1303), .A2(n1302), .ZN(n1299) );
NAND2_X1 U995 ( .A1(G227), .A2(n1041), .ZN(n1302) );
NOR2_X1 U996 ( .A1(n1171), .A2(n1301), .ZN(n1303) );
INV_X1 U997 ( .A(KEYINPUT34), .ZN(n1301) );
XNOR2_X1 U998 ( .A(G140), .B(G110), .ZN(n1171) );
XOR2_X1 U999 ( .A(n1304), .B(n1305), .Z(n1170) );
XOR2_X1 U1000 ( .A(n1287), .B(n1306), .Z(n1305) );
XNOR2_X1 U1001 ( .A(KEYINPUT39), .B(KEYINPUT12), .ZN(n1306) );
NAND3_X1 U1002 ( .A1(n1307), .A2(n1308), .A3(n1112), .ZN(n1287) );
NAND2_X1 U1003 ( .A1(G131), .A2(n1108), .ZN(n1112) );
NOR2_X1 U1004 ( .A1(n1111), .A2(G134), .ZN(n1108) );
NAND2_X1 U1005 ( .A1(n1309), .A2(n1111), .ZN(n1308) );
INV_X1 U1006 ( .A(G137), .ZN(n1111) );
XOR2_X1 U1007 ( .A(n1106), .B(G134), .Z(n1309) );
NAND3_X1 U1008 ( .A1(G134), .A2(n1106), .A3(G137), .ZN(n1307) );
XOR2_X1 U1009 ( .A(n1102), .B(n1310), .Z(n1304) );
XNOR2_X1 U1010 ( .A(n1311), .B(n1312), .ZN(n1102) );
NAND2_X1 U1011 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
XNOR2_X1 U1012 ( .A(KEYINPUT59), .B(KEYINPUT13), .ZN(n1313) );
AND2_X1 U1013 ( .A1(G221), .A2(n1273), .ZN(n1065) );
NAND2_X1 U1014 ( .A1(n1315), .A2(n1177), .ZN(n1273) );
INV_X1 U1015 ( .A(n1253), .ZN(n1192) );
NAND2_X1 U1016 ( .A1(n1229), .A2(n1316), .ZN(n1253) );
NAND2_X1 U1017 ( .A1(n1071), .A2(n1245), .ZN(n1316) );
NAND3_X1 U1018 ( .A1(G902), .A2(n1231), .A3(n1138), .ZN(n1245) );
NOR2_X1 U1019 ( .A1(n1041), .A2(G898), .ZN(n1138) );
NAND3_X1 U1020 ( .A1(n1231), .A2(n1041), .A3(G952), .ZN(n1071) );
NAND2_X1 U1021 ( .A1(G237), .A2(n1315), .ZN(n1231) );
XNOR2_X1 U1022 ( .A(G234), .B(KEYINPUT40), .ZN(n1315) );
INV_X1 U1023 ( .A(n1035), .ZN(n1229) );
NAND2_X1 U1024 ( .A1(n1038), .A2(n1037), .ZN(n1035) );
NAND2_X1 U1025 ( .A1(G214), .A2(n1317), .ZN(n1037) );
XNOR2_X1 U1026 ( .A(n1318), .B(n1088), .ZN(n1038) );
NAND2_X1 U1027 ( .A1(n1319), .A2(n1320), .ZN(n1088) );
XOR2_X1 U1028 ( .A(KEYINPUT1), .B(G902), .Z(n1320) );
XNOR2_X1 U1029 ( .A(n1182), .B(n1321), .ZN(n1319) );
NOR2_X1 U1030 ( .A1(KEYINPUT63), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U1031 ( .A(n1179), .B(KEYINPUT51), .ZN(n1322) );
XNOR2_X1 U1032 ( .A(n1286), .B(G125), .ZN(n1179) );
XNOR2_X1 U1033 ( .A(n1312), .B(n1323), .ZN(n1286) );
NOR2_X1 U1034 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
AND3_X1 U1035 ( .A1(KEYINPUT2), .A2(n1217), .A3(G143), .ZN(n1325) );
NOR2_X1 U1036 ( .A1(KEYINPUT2), .A2(n1314), .ZN(n1324) );
XOR2_X1 U1037 ( .A(G143), .B(G146), .Z(n1314) );
XOR2_X1 U1038 ( .A(G128), .B(KEYINPUT55), .Z(n1312) );
XNOR2_X1 U1039 ( .A(n1326), .B(n1327), .ZN(n1182) );
NOR2_X1 U1040 ( .A1(G953), .A2(n1125), .ZN(n1327) );
INV_X1 U1041 ( .A(G224), .ZN(n1125) );
NAND3_X1 U1042 ( .A1(n1328), .A2(n1329), .A3(n1130), .ZN(n1326) );
NAND3_X1 U1043 ( .A1(n1134), .A2(n1133), .A3(n1310), .ZN(n1130) );
NAND2_X1 U1044 ( .A1(n1135), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1045 ( .A(n1331), .B(n1332), .Z(n1330) );
INV_X1 U1046 ( .A(n1310), .ZN(n1135) );
NAND2_X1 U1047 ( .A1(n1333), .A2(n1310), .ZN(n1328) );
XOR2_X1 U1048 ( .A(n1334), .B(n1335), .Z(n1310) );
XOR2_X1 U1049 ( .A(G104), .B(G101), .Z(n1335) );
XNOR2_X1 U1050 ( .A(G107), .B(KEYINPUT8), .ZN(n1334) );
NAND2_X1 U1051 ( .A1(n1336), .A2(n1337), .ZN(n1333) );
NAND2_X1 U1052 ( .A1(n1331), .A2(n1332), .ZN(n1337) );
INV_X1 U1053 ( .A(n1134), .ZN(n1332) );
NOR2_X1 U1054 ( .A1(n1133), .A2(KEYINPUT29), .ZN(n1331) );
NAND2_X1 U1055 ( .A1(n1338), .A2(n1339), .ZN(n1133) );
NAND2_X1 U1056 ( .A1(n1340), .A2(n1250), .ZN(n1339) );
XOR2_X1 U1057 ( .A(KEYINPUT4), .B(n1341), .Z(n1338) );
NOR2_X1 U1058 ( .A1(n1250), .A2(n1340), .ZN(n1341) );
XOR2_X1 U1059 ( .A(KEYINPUT10), .B(n1280), .Z(n1340) );
XOR2_X1 U1060 ( .A(G116), .B(G119), .Z(n1280) );
INV_X1 U1061 ( .A(G113), .ZN(n1250) );
NAND2_X1 U1062 ( .A1(KEYINPUT29), .A2(n1134), .ZN(n1336) );
XOR2_X1 U1063 ( .A(G110), .B(G122), .Z(n1134) );
NAND2_X1 U1064 ( .A1(KEYINPUT23), .A2(n1086), .ZN(n1318) );
NAND2_X1 U1065 ( .A1(G210), .A2(n1317), .ZN(n1086) );
NAND2_X1 U1066 ( .A1(n1342), .A2(n1343), .ZN(n1317) );
INV_X1 U1067 ( .A(G237), .ZN(n1343) );
XOR2_X1 U1068 ( .A(KEYINPUT45), .B(G902), .Z(n1342) );
NOR2_X1 U1069 ( .A1(n1239), .A2(n1238), .ZN(n1056) );
XNOR2_X1 U1070 ( .A(n1344), .B(G475), .ZN(n1238) );
NAND2_X1 U1071 ( .A1(n1149), .A2(n1177), .ZN(n1344) );
XNOR2_X1 U1072 ( .A(n1345), .B(n1346), .ZN(n1149) );
XOR2_X1 U1073 ( .A(n1271), .B(n1347), .Z(n1346) );
XOR2_X1 U1074 ( .A(n1348), .B(n1349), .Z(n1347) );
NAND2_X1 U1075 ( .A1(n1282), .A2(G214), .ZN(n1349) );
NOR2_X1 U1076 ( .A1(G953), .A2(G237), .ZN(n1282) );
NAND2_X1 U1077 ( .A1(n1350), .A2(n1351), .ZN(n1348) );
NAND2_X1 U1078 ( .A1(G104), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1079 ( .A(KEYINPUT44), .B(n1353), .Z(n1350) );
NOR2_X1 U1080 ( .A1(G104), .A2(n1352), .ZN(n1353) );
XOR2_X1 U1081 ( .A(G122), .B(G113), .Z(n1352) );
XNOR2_X1 U1082 ( .A(n1217), .B(KEYINPUT54), .ZN(n1271) );
INV_X1 U1083 ( .A(G146), .ZN(n1217) );
XOR2_X1 U1084 ( .A(n1354), .B(n1355), .Z(n1345) );
XOR2_X1 U1085 ( .A(KEYINPUT32), .B(G143), .Z(n1355) );
XOR2_X1 U1086 ( .A(n1106), .B(n1356), .Z(n1354) );
NOR2_X1 U1087 ( .A1(KEYINPUT50), .A2(n1357), .ZN(n1356) );
XNOR2_X1 U1088 ( .A(n1272), .B(KEYINPUT41), .ZN(n1357) );
XOR2_X1 U1089 ( .A(n1097), .B(KEYINPUT21), .Z(n1272) );
XOR2_X1 U1090 ( .A(G125), .B(G140), .Z(n1097) );
INV_X1 U1091 ( .A(G131), .ZN(n1106) );
INV_X1 U1092 ( .A(n1249), .ZN(n1239) );
XOR2_X1 U1093 ( .A(n1358), .B(G478), .Z(n1249) );
NAND2_X1 U1094 ( .A1(n1146), .A2(n1177), .ZN(n1358) );
INV_X1 U1095 ( .A(G902), .ZN(n1177) );
XNOR2_X1 U1096 ( .A(n1359), .B(n1360), .ZN(n1146) );
XOR2_X1 U1097 ( .A(n1361), .B(n1362), .Z(n1360) );
XOR2_X1 U1098 ( .A(n1363), .B(n1364), .Z(n1362) );
AND3_X1 U1099 ( .A1(G217), .A2(n1041), .A3(G234), .ZN(n1364) );
INV_X1 U1100 ( .A(G953), .ZN(n1041) );
NAND2_X1 U1101 ( .A1(KEYINPUT30), .A2(G116), .ZN(n1363) );
XOR2_X1 U1102 ( .A(G107), .B(n1235), .Z(n1361) );
INV_X1 U1103 ( .A(G122), .ZN(n1235) );
XOR2_X1 U1104 ( .A(n1365), .B(n1366), .Z(n1359) );
XOR2_X1 U1105 ( .A(KEYINPUT31), .B(G143), .Z(n1366) );
XNOR2_X1 U1106 ( .A(G128), .B(G134), .ZN(n1365) );
endmodule


