//Key = 0101100010111110000101010101010111010000001111111110001101000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434;

XOR2_X1 U788 ( .A(n1080), .B(n1081), .Z(G9) );
XNOR2_X1 U789 ( .A(G107), .B(KEYINPUT15), .ZN(n1081) );
NOR2_X1 U790 ( .A1(n1082), .A2(n1083), .ZN(G75) );
NOR4_X1 U791 ( .A1(G953), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1083) );
NOR2_X1 U792 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U793 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR3_X1 U794 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NOR2_X1 U795 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U796 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U797 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NOR2_X1 U798 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U799 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U800 ( .A1(n1104), .A2(n1105), .ZN(n1098) );
NOR2_X1 U801 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U802 ( .A1(n1108), .A2(n1105), .ZN(n1094) );
NOR2_X1 U803 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR3_X1 U804 ( .A1(n1111), .A2(n1101), .A3(n1112), .ZN(n1109) );
NOR4_X1 U805 ( .A1(n1113), .A2(n1105), .A3(n1097), .A4(n1101), .ZN(n1089) );
NOR2_X1 U806 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U807 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
XNOR2_X1 U808 ( .A(KEYINPUT0), .B(n1118), .ZN(n1117) );
NOR3_X1 U809 ( .A1(n1084), .A2(G953), .A3(G952), .ZN(n1082) );
AND4_X1 U810 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1084) );
NOR4_X1 U811 ( .A1(n1123), .A2(n1092), .A3(n1124), .A4(n1125), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1126), .A2(n1127), .ZN(n1121) );
XNOR2_X1 U813 ( .A(KEYINPUT5), .B(n1128), .ZN(n1127) );
XNOR2_X1 U814 ( .A(G469), .B(n1129), .ZN(n1126) );
XNOR2_X1 U815 ( .A(n1130), .B(n1131), .ZN(n1120) );
NOR2_X1 U816 ( .A1(KEYINPUT62), .A2(n1132), .ZN(n1131) );
XNOR2_X1 U817 ( .A(n1133), .B(n1134), .ZN(n1119) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(G72) );
NOR2_X1 U819 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U820 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U821 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U822 ( .A(G131), .B(n1143), .ZN(n1142) );
XOR2_X1 U823 ( .A(n1144), .B(n1145), .Z(n1139) );
XOR2_X1 U824 ( .A(n1146), .B(n1147), .Z(n1144) );
NOR2_X1 U825 ( .A1(G125), .A2(KEYINPUT28), .ZN(n1147) );
NAND3_X1 U826 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1146) );
NAND2_X1 U827 ( .A1(KEYINPUT20), .A2(n1151), .ZN(n1150) );
NAND2_X1 U828 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U829 ( .A1(G134), .A2(n1154), .ZN(n1153) );
NAND4_X1 U830 ( .A1(n1152), .A2(n1155), .A3(KEYINPUT32), .A4(G134), .ZN(n1149) );
NAND2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(n1148) );
NAND3_X1 U832 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1156) );
NAND2_X1 U833 ( .A1(KEYINPUT32), .A2(KEYINPUT20), .ZN(n1160) );
OR2_X1 U834 ( .A1(G137), .A2(KEYINPUT4), .ZN(n1159) );
NAND2_X1 U835 ( .A1(KEYINPUT4), .A2(n1161), .ZN(n1158) );
NAND2_X1 U836 ( .A1(n1152), .A2(n1162), .ZN(n1161) );
NAND2_X1 U837 ( .A1(n1155), .A2(n1154), .ZN(n1162) );
INV_X1 U838 ( .A(KEYINPUT32), .ZN(n1154) );
INV_X1 U839 ( .A(KEYINPUT20), .ZN(n1155) );
NOR2_X1 U840 ( .A1(G900), .A2(n1163), .ZN(n1137) );
XOR2_X1 U841 ( .A(n1164), .B(n1165), .Z(n1135) );
NOR2_X1 U842 ( .A1(G953), .A2(n1166), .ZN(n1165) );
XNOR2_X1 U843 ( .A(n1167), .B(KEYINPUT10), .ZN(n1166) );
NAND2_X1 U844 ( .A1(KEYINPUT47), .A2(n1168), .ZN(n1164) );
NAND2_X1 U845 ( .A1(G953), .A2(n1169), .ZN(n1168) );
NAND2_X1 U846 ( .A1(G900), .A2(n1170), .ZN(n1169) );
XOR2_X1 U847 ( .A(KEYINPUT22), .B(G227), .Z(n1170) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(G69) );
NOR2_X1 U849 ( .A1(KEYINPUT39), .A2(n1173), .ZN(n1172) );
XOR2_X1 U850 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U851 ( .A1(n1163), .A2(n1176), .ZN(n1175) );
NAND2_X1 U852 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND4_X1 U853 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1174) );
NAND4_X1 U854 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
INV_X1 U855 ( .A(n1187), .ZN(n1186) );
NAND4_X1 U856 ( .A1(n1185), .A2(n1184), .A3(n1188), .A4(n1187), .ZN(n1181) );
XOR2_X1 U857 ( .A(n1183), .B(KEYINPUT29), .Z(n1188) );
NAND2_X1 U858 ( .A1(G953), .A2(n1189), .ZN(n1180) );
NAND2_X1 U859 ( .A1(n1190), .A2(n1191), .ZN(n1179) );
NAND2_X1 U860 ( .A1(n1192), .A2(n1184), .ZN(n1191) );
INV_X1 U861 ( .A(KEYINPUT63), .ZN(n1184) );
XOR2_X1 U862 ( .A(n1183), .B(n1193), .Z(n1192) );
AND2_X1 U863 ( .A1(n1187), .A2(KEYINPUT29), .ZN(n1193) );
INV_X1 U864 ( .A(n1185), .ZN(n1190) );
NAND2_X1 U865 ( .A1(G953), .A2(n1194), .ZN(n1171) );
NAND2_X1 U866 ( .A1(G898), .A2(G224), .ZN(n1194) );
NOR2_X1 U867 ( .A1(n1195), .A2(n1196), .ZN(G66) );
NOR3_X1 U868 ( .A1(n1130), .A2(n1197), .A3(n1198), .ZN(n1196) );
NOR3_X1 U869 ( .A1(n1199), .A2(n1132), .A3(n1200), .ZN(n1198) );
INV_X1 U870 ( .A(n1201), .ZN(n1199) );
NOR2_X1 U871 ( .A1(n1202), .A2(n1201), .ZN(n1197) );
NOR2_X1 U872 ( .A1(n1203), .A2(n1132), .ZN(n1202) );
NOR2_X1 U873 ( .A1(n1195), .A2(n1204), .ZN(G63) );
XNOR2_X1 U874 ( .A(n1205), .B(n1206), .ZN(n1204) );
AND2_X1 U875 ( .A1(G478), .A2(n1207), .ZN(n1205) );
NOR2_X1 U876 ( .A1(n1195), .A2(n1208), .ZN(G60) );
XNOR2_X1 U877 ( .A(n1209), .B(n1210), .ZN(n1208) );
NAND2_X1 U878 ( .A1(KEYINPUT23), .A2(n1211), .ZN(n1209) );
NAND3_X1 U879 ( .A1(n1212), .A2(n1213), .A3(G475), .ZN(n1211) );
NAND2_X1 U880 ( .A1(KEYINPUT33), .A2(n1200), .ZN(n1213) );
INV_X1 U881 ( .A(n1207), .ZN(n1200) );
NAND2_X1 U882 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
INV_X1 U883 ( .A(KEYINPUT33), .ZN(n1215) );
NAND2_X1 U884 ( .A1(n1203), .A2(G902), .ZN(n1214) );
XNOR2_X1 U885 ( .A(G104), .B(n1216), .ZN(G6) );
NOR2_X1 U886 ( .A1(n1195), .A2(n1217), .ZN(G57) );
XOR2_X1 U887 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U888 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U889 ( .A(G101), .B(n1222), .Z(n1221) );
NOR2_X1 U890 ( .A1(KEYINPUT18), .A2(n1223), .ZN(n1220) );
XOR2_X1 U891 ( .A(n1224), .B(n1225), .Z(n1218) );
NAND2_X1 U892 ( .A1(n1207), .A2(G472), .ZN(n1224) );
NOR2_X1 U893 ( .A1(n1195), .A2(n1226), .ZN(G54) );
XNOR2_X1 U894 ( .A(n1227), .B(n1228), .ZN(n1226) );
XOR2_X1 U895 ( .A(n1229), .B(n1230), .Z(n1228) );
NOR2_X1 U896 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U897 ( .A(KEYINPUT17), .B(n1233), .Z(n1232) );
NOR2_X1 U898 ( .A1(n1223), .A2(n1234), .ZN(n1233) );
XOR2_X1 U899 ( .A(n1235), .B(KEYINPUT9), .Z(n1234) );
NAND3_X1 U900 ( .A1(n1207), .A2(G469), .A3(KEYINPUT31), .ZN(n1229) );
NOR2_X1 U901 ( .A1(n1195), .A2(n1236), .ZN(G51) );
XOR2_X1 U902 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U903 ( .A(n1239), .B(n1240), .ZN(n1238) );
NAND2_X1 U904 ( .A1(n1207), .A2(n1241), .ZN(n1239) );
NOR2_X1 U905 ( .A1(n1242), .A2(n1203), .ZN(n1207) );
INV_X1 U906 ( .A(n1086), .ZN(n1203) );
NAND3_X1 U907 ( .A1(n1167), .A2(n1178), .A3(n1177), .ZN(n1086) );
AND4_X1 U908 ( .A1(n1216), .A2(n1243), .A3(n1080), .A4(n1244), .ZN(n1177) );
AND2_X1 U909 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND4_X1 U910 ( .A1(n1247), .A2(n1248), .A3(n1106), .A4(n1249), .ZN(n1080) );
NAND4_X1 U911 ( .A1(n1107), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1216) );
NAND2_X1 U912 ( .A1(n1250), .A2(n1251), .ZN(n1178) );
NAND2_X1 U913 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND4_X1 U914 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1253) );
INV_X1 U915 ( .A(KEYINPUT42), .ZN(n1257) );
NAND2_X1 U916 ( .A1(n1248), .A2(n1258), .ZN(n1252) );
NAND3_X1 U917 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1258) );
NAND2_X1 U918 ( .A1(n1106), .A2(n1103), .ZN(n1261) );
NAND2_X1 U919 ( .A1(KEYINPUT42), .A2(n1254), .ZN(n1260) );
NAND2_X1 U920 ( .A1(n1262), .A2(n1249), .ZN(n1259) );
AND4_X1 U921 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1167) );
NOR4_X1 U922 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1266) );
NAND2_X1 U923 ( .A1(n1271), .A2(n1272), .ZN(n1265) );
NAND2_X1 U924 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND4_X1 U925 ( .A1(n1275), .A2(n1118), .A3(n1110), .A4(n1116), .ZN(n1274) );
XOR2_X1 U926 ( .A(n1276), .B(KEYINPUT16), .Z(n1275) );
NAND2_X1 U927 ( .A1(n1277), .A2(n1106), .ZN(n1273) );
NAND3_X1 U928 ( .A1(n1262), .A2(n1103), .A3(n1277), .ZN(n1263) );
NOR2_X1 U929 ( .A1(n1163), .A2(G952), .ZN(n1195) );
XNOR2_X1 U930 ( .A(n1264), .B(n1278), .ZN(G48) );
NOR2_X1 U931 ( .A1(KEYINPUT40), .A2(n1279), .ZN(n1278) );
NAND3_X1 U932 ( .A1(n1271), .A2(n1107), .A3(n1277), .ZN(n1264) );
NAND2_X1 U933 ( .A1(n1280), .A2(n1281), .ZN(G45) );
NAND2_X1 U934 ( .A1(G143), .A2(n1282), .ZN(n1281) );
XOR2_X1 U935 ( .A(KEYINPUT27), .B(n1283), .Z(n1280) );
NOR2_X1 U936 ( .A1(G143), .A2(n1282), .ZN(n1283) );
NAND4_X1 U937 ( .A1(n1284), .A2(n1276), .A3(n1103), .A4(n1285), .ZN(n1282) );
NOR2_X1 U938 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XNOR2_X1 U939 ( .A(KEYINPUT41), .B(n1256), .ZN(n1284) );
XOR2_X1 U940 ( .A(G140), .B(n1270), .Z(G42) );
AND3_X1 U941 ( .A1(n1102), .A2(n1107), .A3(n1288), .ZN(n1270) );
XNOR2_X1 U942 ( .A(n1152), .B(n1289), .ZN(G39) );
NOR2_X1 U943 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XNOR2_X1 U944 ( .A(n1157), .B(n1269), .ZN(G36) );
AND3_X1 U945 ( .A1(n1106), .A2(n1103), .A3(n1288), .ZN(n1269) );
XOR2_X1 U946 ( .A(G131), .B(n1268), .Z(G33) );
AND2_X1 U947 ( .A1(n1288), .A2(n1254), .ZN(n1268) );
INV_X1 U948 ( .A(n1291), .ZN(n1288) );
NAND4_X1 U949 ( .A1(n1118), .A2(n1247), .A3(n1276), .A4(n1116), .ZN(n1291) );
XNOR2_X1 U950 ( .A(G128), .B(n1292), .ZN(G30) );
NAND4_X1 U951 ( .A1(n1293), .A2(KEYINPUT21), .A3(n1277), .A4(n1106), .ZN(n1292) );
AND3_X1 U952 ( .A1(n1115), .A2(n1276), .A3(n1247), .ZN(n1277) );
XNOR2_X1 U953 ( .A(n1271), .B(KEYINPUT25), .ZN(n1293) );
INV_X1 U954 ( .A(n1294), .ZN(n1271) );
XNOR2_X1 U955 ( .A(G101), .B(n1243), .ZN(G3) );
NAND3_X1 U956 ( .A1(n1248), .A2(n1103), .A3(n1110), .ZN(n1243) );
XOR2_X1 U957 ( .A(G125), .B(n1267), .Z(G27) );
AND4_X1 U958 ( .A1(n1115), .A2(n1276), .A3(n1107), .A4(n1295), .ZN(n1267) );
NOR2_X1 U959 ( .A1(n1097), .A2(n1296), .ZN(n1295) );
NAND2_X1 U960 ( .A1(n1088), .A2(n1297), .ZN(n1276) );
NAND4_X1 U961 ( .A1(G953), .A2(G902), .A3(n1298), .A4(n1299), .ZN(n1297) );
INV_X1 U962 ( .A(G900), .ZN(n1299) );
NAND2_X1 U963 ( .A1(n1300), .A2(n1301), .ZN(G24) );
NAND3_X1 U964 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1301) );
INV_X1 U965 ( .A(KEYINPUT37), .ZN(n1304) );
NAND2_X1 U966 ( .A1(G122), .A2(KEYINPUT12), .ZN(n1303) );
NAND2_X1 U967 ( .A1(n1305), .A2(n1306), .ZN(n1302) );
NAND4_X1 U968 ( .A1(n1115), .A2(n1249), .A3(n1262), .A4(n1307), .ZN(n1305) );
NOR3_X1 U969 ( .A1(n1308), .A2(n1097), .A3(n1309), .ZN(n1307) );
INV_X1 U970 ( .A(KEYINPUT12), .ZN(n1309) );
XNOR2_X1 U971 ( .A(KEYINPUT51), .B(n1255), .ZN(n1308) );
NAND2_X1 U972 ( .A1(n1310), .A2(n1311), .ZN(n1300) );
NAND4_X1 U973 ( .A1(n1312), .A2(n1313), .A3(n1250), .A4(n1314), .ZN(n1311) );
NOR2_X1 U974 ( .A1(n1105), .A2(n1287), .ZN(n1314) );
INV_X1 U975 ( .A(n1262), .ZN(n1287) );
NOR2_X1 U976 ( .A1(n1315), .A2(n1128), .ZN(n1262) );
INV_X1 U977 ( .A(n1249), .ZN(n1105) );
NAND2_X1 U978 ( .A1(n1316), .A2(n1317), .ZN(n1249) );
NAND2_X1 U979 ( .A1(n1103), .A2(n1318), .ZN(n1317) );
OR3_X1 U980 ( .A1(n1319), .A2(n1125), .A3(n1318), .ZN(n1316) );
INV_X1 U981 ( .A(KEYINPUT46), .ZN(n1318) );
OR2_X1 U982 ( .A1(n1248), .A2(KEYINPUT51), .ZN(n1313) );
NAND2_X1 U983 ( .A1(KEYINPUT51), .A2(n1320), .ZN(n1312) );
OR2_X1 U984 ( .A1(n1255), .A2(n1256), .ZN(n1320) );
NAND2_X1 U985 ( .A1(n1321), .A2(n1306), .ZN(n1310) );
NAND2_X1 U986 ( .A1(KEYINPUT37), .A2(KEYINPUT12), .ZN(n1321) );
NAND2_X1 U987 ( .A1(n1322), .A2(n1323), .ZN(G21) );
OR2_X1 U988 ( .A1(n1246), .A2(G119), .ZN(n1323) );
XOR2_X1 U989 ( .A(n1324), .B(KEYINPUT2), .Z(n1322) );
NAND2_X1 U990 ( .A1(G119), .A2(n1246), .ZN(n1324) );
OR3_X1 U991 ( .A1(n1097), .A2(n1325), .A3(n1290), .ZN(n1246) );
OR2_X1 U992 ( .A1(n1294), .A2(n1101), .ZN(n1290) );
NAND2_X1 U993 ( .A1(n1326), .A2(n1125), .ZN(n1294) );
INV_X1 U994 ( .A(n1250), .ZN(n1097) );
XNOR2_X1 U995 ( .A(G116), .B(n1327), .ZN(G18) );
NAND4_X1 U996 ( .A1(n1328), .A2(n1255), .A3(n1103), .A4(n1329), .ZN(n1327) );
AND2_X1 U997 ( .A1(n1106), .A2(n1250), .ZN(n1329) );
NOR2_X1 U998 ( .A1(n1128), .A2(n1124), .ZN(n1106) );
INV_X1 U999 ( .A(n1315), .ZN(n1124) );
XNOR2_X1 U1000 ( .A(KEYINPUT38), .B(n1256), .ZN(n1328) );
INV_X1 U1001 ( .A(n1115), .ZN(n1256) );
XNOR2_X1 U1002 ( .A(G113), .B(n1330), .ZN(G15) );
NAND3_X1 U1003 ( .A1(n1254), .A2(n1248), .A3(n1250), .ZN(n1330) );
NOR2_X1 U1004 ( .A1(n1112), .A2(n1123), .ZN(n1250) );
AND2_X1 U1005 ( .A1(n1107), .A2(n1103), .ZN(n1254) );
NOR2_X1 U1006 ( .A1(n1331), .A2(n1319), .ZN(n1103) );
NOR2_X1 U1007 ( .A1(n1315), .A2(n1332), .ZN(n1107) );
XNOR2_X1 U1008 ( .A(G110), .B(n1245), .ZN(G12) );
NAND3_X1 U1009 ( .A1(n1110), .A2(n1248), .A3(n1102), .ZN(n1245) );
INV_X1 U1010 ( .A(n1296), .ZN(n1102) );
NAND2_X1 U1011 ( .A1(n1331), .A2(n1326), .ZN(n1296) );
XNOR2_X1 U1012 ( .A(n1319), .B(KEYINPUT14), .ZN(n1326) );
XNOR2_X1 U1013 ( .A(n1333), .B(n1132), .ZN(n1319) );
NAND2_X1 U1014 ( .A1(G217), .A2(n1334), .ZN(n1132) );
XNOR2_X1 U1015 ( .A(n1130), .B(KEYINPUT45), .ZN(n1333) );
NOR2_X1 U1016 ( .A1(n1201), .A2(G902), .ZN(n1130) );
XNOR2_X1 U1017 ( .A(n1335), .B(n1336), .ZN(n1201) );
XOR2_X1 U1018 ( .A(n1337), .B(n1338), .Z(n1336) );
NAND2_X1 U1019 ( .A1(n1339), .A2(G221), .ZN(n1338) );
NAND2_X1 U1020 ( .A1(n1340), .A2(n1341), .ZN(n1337) );
OR2_X1 U1021 ( .A1(n1342), .A2(n1279), .ZN(n1341) );
XOR2_X1 U1022 ( .A(n1343), .B(KEYINPUT60), .Z(n1340) );
NAND2_X1 U1023 ( .A1(n1342), .A2(n1279), .ZN(n1343) );
INV_X1 U1024 ( .A(G146), .ZN(n1279) );
XOR2_X1 U1025 ( .A(G125), .B(n1145), .Z(n1342) );
XOR2_X1 U1026 ( .A(n1344), .B(n1345), .Z(n1335) );
XNOR2_X1 U1027 ( .A(n1152), .B(G110), .ZN(n1345) );
NAND2_X1 U1028 ( .A1(n1346), .A2(n1347), .ZN(n1344) );
NAND2_X1 U1029 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1030 ( .A(KEYINPUT8), .B(n1350), .Z(n1346) );
NOR2_X1 U1031 ( .A1(n1349), .A2(n1348), .ZN(n1350) );
XNOR2_X1 U1032 ( .A(KEYINPUT58), .B(G128), .ZN(n1348) );
INV_X1 U1033 ( .A(n1125), .ZN(n1331) );
XNOR2_X1 U1034 ( .A(n1351), .B(G472), .ZN(n1125) );
NAND2_X1 U1035 ( .A1(n1352), .A2(n1242), .ZN(n1351) );
XOR2_X1 U1036 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1037 ( .A(n1225), .B(n1355), .ZN(n1354) );
XNOR2_X1 U1038 ( .A(n1356), .B(n1357), .ZN(n1225) );
XOR2_X1 U1039 ( .A(n1358), .B(G113), .Z(n1356) );
NAND2_X1 U1040 ( .A1(KEYINPUT54), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1041 ( .A(n1360), .B(n1222), .Z(n1353) );
AND3_X1 U1042 ( .A1(G210), .A2(n1361), .A3(n1362), .ZN(n1222) );
XNOR2_X1 U1043 ( .A(G953), .B(KEYINPUT30), .ZN(n1362) );
NAND2_X1 U1044 ( .A1(KEYINPUT57), .A2(G101), .ZN(n1360) );
INV_X1 U1045 ( .A(n1325), .ZN(n1248) );
NAND2_X1 U1046 ( .A1(n1115), .A2(n1255), .ZN(n1325) );
NAND2_X1 U1047 ( .A1(n1088), .A2(n1363), .ZN(n1255) );
NAND4_X1 U1048 ( .A1(G953), .A2(G902), .A3(n1298), .A4(n1189), .ZN(n1363) );
INV_X1 U1049 ( .A(G898), .ZN(n1189) );
NAND3_X1 U1050 ( .A1(n1298), .A2(n1163), .A3(G952), .ZN(n1088) );
NAND2_X1 U1051 ( .A1(G237), .A2(G234), .ZN(n1298) );
NOR2_X1 U1052 ( .A1(n1118), .A2(n1092), .ZN(n1115) );
INV_X1 U1053 ( .A(n1116), .ZN(n1092) );
NAND2_X1 U1054 ( .A1(G214), .A2(n1364), .ZN(n1116) );
INV_X1 U1055 ( .A(n1091), .ZN(n1118) );
XOR2_X1 U1056 ( .A(n1241), .B(n1365), .Z(n1091) );
NOR2_X1 U1057 ( .A1(KEYINPUT56), .A2(n1133), .ZN(n1365) );
NAND2_X1 U1058 ( .A1(n1366), .A2(n1242), .ZN(n1133) );
XOR2_X1 U1059 ( .A(n1367), .B(n1368), .Z(n1366) );
NAND2_X1 U1060 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
NAND2_X1 U1061 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
INV_X1 U1062 ( .A(KEYINPUT3), .ZN(n1372) );
XNOR2_X1 U1063 ( .A(n1373), .B(n1374), .ZN(n1371) );
NOR2_X1 U1064 ( .A1(n1357), .A2(n1375), .ZN(n1374) );
NAND2_X1 U1065 ( .A1(KEYINPUT3), .A2(n1237), .ZN(n1369) );
XNOR2_X1 U1066 ( .A(n1376), .B(n1377), .ZN(n1237) );
INV_X1 U1067 ( .A(n1373), .ZN(n1377) );
XNOR2_X1 U1068 ( .A(n1378), .B(n1379), .ZN(n1373) );
XNOR2_X1 U1069 ( .A(n1185), .B(n1187), .ZN(n1379) );
XOR2_X1 U1070 ( .A(G107), .B(n1380), .Z(n1187) );
XOR2_X1 U1071 ( .A(G110), .B(n1306), .Z(n1185) );
XOR2_X1 U1072 ( .A(n1183), .B(KEYINPUT19), .Z(n1378) );
XNOR2_X1 U1073 ( .A(n1381), .B(n1359), .ZN(n1183) );
XOR2_X1 U1074 ( .A(G116), .B(n1349), .Z(n1359) );
XNOR2_X1 U1075 ( .A(G119), .B(KEYINPUT13), .ZN(n1349) );
NAND2_X1 U1076 ( .A1(KEYINPUT1), .A2(G113), .ZN(n1381) );
XNOR2_X1 U1077 ( .A(n1357), .B(n1375), .ZN(n1376) );
XOR2_X1 U1078 ( .A(G125), .B(KEYINPUT44), .Z(n1375) );
XNOR2_X1 U1079 ( .A(G128), .B(n1382), .ZN(n1357) );
NAND2_X1 U1080 ( .A1(KEYINPUT35), .A2(n1240), .ZN(n1367) );
NAND2_X1 U1081 ( .A1(G224), .A2(n1163), .ZN(n1240) );
INV_X1 U1082 ( .A(n1134), .ZN(n1241) );
NAND2_X1 U1083 ( .A1(G210), .A2(n1364), .ZN(n1134) );
NAND2_X1 U1084 ( .A1(n1361), .A2(n1242), .ZN(n1364) );
NOR2_X1 U1085 ( .A1(n1101), .A2(n1286), .ZN(n1110) );
INV_X1 U1086 ( .A(n1247), .ZN(n1286) );
NOR2_X1 U1087 ( .A1(n1383), .A2(n1123), .ZN(n1247) );
INV_X1 U1088 ( .A(n1111), .ZN(n1123) );
NAND2_X1 U1089 ( .A1(G221), .A2(n1334), .ZN(n1111) );
NAND2_X1 U1090 ( .A1(G234), .A2(n1242), .ZN(n1334) );
INV_X1 U1091 ( .A(n1112), .ZN(n1383) );
XNOR2_X1 U1092 ( .A(n1129), .B(n1384), .ZN(n1112) );
NOR2_X1 U1093 ( .A1(KEYINPUT52), .A2(n1385), .ZN(n1384) );
INV_X1 U1094 ( .A(G469), .ZN(n1385) );
NAND3_X1 U1095 ( .A1(n1386), .A2(n1242), .A3(n1387), .ZN(n1129) );
NAND2_X1 U1096 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NAND2_X1 U1097 ( .A1(n1390), .A2(n1391), .ZN(n1388) );
NAND3_X1 U1098 ( .A1(n1392), .A2(n1393), .A3(n1235), .ZN(n1391) );
NAND2_X1 U1099 ( .A1(KEYINPUT43), .A2(n1394), .ZN(n1393) );
NAND2_X1 U1100 ( .A1(n1395), .A2(n1355), .ZN(n1394) );
INV_X1 U1101 ( .A(n1227), .ZN(n1395) );
OR2_X1 U1102 ( .A1(n1227), .A2(KEYINPUT43), .ZN(n1392) );
NAND2_X1 U1103 ( .A1(n1231), .A2(n1227), .ZN(n1390) );
AND2_X1 U1104 ( .A1(n1223), .A2(n1235), .ZN(n1231) );
NAND2_X1 U1105 ( .A1(n1396), .A2(n1397), .ZN(n1386) );
NAND2_X1 U1106 ( .A1(n1235), .A2(n1389), .ZN(n1397) );
INV_X1 U1107 ( .A(KEYINPUT36), .ZN(n1389) );
XOR2_X1 U1108 ( .A(n1398), .B(n1380), .Z(n1235) );
XNOR2_X1 U1109 ( .A(n1399), .B(G101), .ZN(n1380) );
XNOR2_X1 U1110 ( .A(n1400), .B(n1141), .ZN(n1398) );
NOR2_X1 U1111 ( .A1(KEYINPUT34), .A2(n1382), .ZN(n1141) );
XNOR2_X1 U1112 ( .A(n1401), .B(n1227), .ZN(n1396) );
XOR2_X1 U1113 ( .A(n1145), .B(n1402), .Z(n1227) );
XOR2_X1 U1114 ( .A(G110), .B(n1403), .Z(n1402) );
AND2_X1 U1115 ( .A1(n1163), .A2(G227), .ZN(n1403) );
NAND2_X1 U1116 ( .A1(KEYINPUT43), .A2(n1223), .ZN(n1401) );
INV_X1 U1117 ( .A(n1355), .ZN(n1223) );
XNOR2_X1 U1118 ( .A(n1404), .B(G131), .ZN(n1355) );
NAND3_X1 U1119 ( .A1(n1405), .A2(n1406), .A3(n1407), .ZN(n1404) );
OR2_X1 U1120 ( .A1(n1152), .A2(n1408), .ZN(n1407) );
NAND3_X1 U1121 ( .A1(n1408), .A2(n1152), .A3(KEYINPUT11), .ZN(n1406) );
INV_X1 U1122 ( .A(G137), .ZN(n1152) );
NOR2_X1 U1123 ( .A1(G134), .A2(KEYINPUT59), .ZN(n1408) );
OR2_X1 U1124 ( .A1(n1157), .A2(KEYINPUT11), .ZN(n1405) );
NAND2_X1 U1125 ( .A1(n1128), .A2(n1315), .ZN(n1101) );
XNOR2_X1 U1126 ( .A(n1409), .B(n1410), .ZN(n1315) );
XOR2_X1 U1127 ( .A(KEYINPUT55), .B(G475), .Z(n1410) );
NAND2_X1 U1128 ( .A1(n1210), .A2(n1242), .ZN(n1409) );
INV_X1 U1129 ( .A(G902), .ZN(n1242) );
XNOR2_X1 U1130 ( .A(n1411), .B(n1412), .ZN(n1210) );
XNOR2_X1 U1131 ( .A(n1413), .B(n1382), .ZN(n1412) );
XNOR2_X1 U1132 ( .A(G143), .B(G146), .ZN(n1382) );
AND3_X1 U1133 ( .A1(G214), .A2(n1163), .A3(n1361), .ZN(n1413) );
INV_X1 U1134 ( .A(G237), .ZN(n1361) );
XOR2_X1 U1135 ( .A(n1414), .B(n1415), .Z(n1411) );
NOR2_X1 U1136 ( .A1(G131), .A2(KEYINPUT24), .ZN(n1415) );
XOR2_X1 U1137 ( .A(n1416), .B(n1417), .Z(n1414) );
NOR2_X1 U1138 ( .A1(KEYINPUT61), .A2(n1418), .ZN(n1417) );
XOR2_X1 U1139 ( .A(n1419), .B(n1420), .Z(n1418) );
XNOR2_X1 U1140 ( .A(n1306), .B(G113), .ZN(n1420) );
INV_X1 U1141 ( .A(G122), .ZN(n1306) );
NOR2_X1 U1142 ( .A1(KEYINPUT7), .A2(n1399), .ZN(n1419) );
INV_X1 U1143 ( .A(G104), .ZN(n1399) );
NAND2_X1 U1144 ( .A1(n1421), .A2(n1422), .ZN(n1416) );
NAND2_X1 U1145 ( .A1(n1423), .A2(n1424), .ZN(n1422) );
XOR2_X1 U1146 ( .A(KEYINPUT26), .B(n1145), .Z(n1424) );
XNOR2_X1 U1147 ( .A(G125), .B(KEYINPUT6), .ZN(n1423) );
NAND2_X1 U1148 ( .A1(n1425), .A2(n1426), .ZN(n1421) );
XNOR2_X1 U1149 ( .A(KEYINPUT26), .B(n1145), .ZN(n1426) );
XOR2_X1 U1150 ( .A(G140), .B(KEYINPUT50), .Z(n1145) );
XNOR2_X1 U1151 ( .A(G125), .B(KEYINPUT48), .ZN(n1425) );
INV_X1 U1152 ( .A(n1332), .ZN(n1128) );
XNOR2_X1 U1153 ( .A(n1427), .B(G478), .ZN(n1332) );
NAND2_X1 U1154 ( .A1(n1428), .A2(n1206), .ZN(n1427) );
XOR2_X1 U1155 ( .A(n1429), .B(n1430), .Z(n1206) );
XOR2_X1 U1156 ( .A(n1431), .B(n1432), .Z(n1430) );
XNOR2_X1 U1157 ( .A(n1157), .B(G122), .ZN(n1432) );
INV_X1 U1158 ( .A(G134), .ZN(n1157) );
XOR2_X1 U1159 ( .A(KEYINPUT49), .B(G143), .Z(n1431) );
XOR2_X1 U1160 ( .A(n1433), .B(n1400), .Z(n1429) );
XNOR2_X1 U1161 ( .A(G107), .B(n1143), .ZN(n1400) );
INV_X1 U1162 ( .A(G128), .ZN(n1143) );
XOR2_X1 U1163 ( .A(n1434), .B(G116), .Z(n1433) );
NAND2_X1 U1164 ( .A1(G217), .A2(n1339), .ZN(n1434) );
AND2_X1 U1165 ( .A1(G234), .A2(n1163), .ZN(n1339) );
INV_X1 U1166 ( .A(G953), .ZN(n1163) );
XNOR2_X1 U1167 ( .A(G902), .B(KEYINPUT53), .ZN(n1428) );
endmodule


