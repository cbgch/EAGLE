//Key = 1110001011110001110100100000011011000010101111100001111111011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305;

XOR2_X1 U725 ( .A(n999), .B(n1000), .Z(G9) );
XNOR2_X1 U726 ( .A(G107), .B(KEYINPUT39), .ZN(n1000) );
NAND3_X1 U727 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(G75) );
NOR3_X1 U728 ( .A1(n1004), .A2(G953), .A3(n1005), .ZN(n1003) );
NOR4_X1 U729 ( .A1(n1006), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n1005) );
NAND4_X1 U730 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1006) );
OR2_X1 U731 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND3_X1 U732 ( .A1(n1016), .A2(n1017), .A3(n1014), .ZN(n1012) );
NOR3_X1 U733 ( .A1(n1018), .A2(n1019), .A3(n1009), .ZN(n1004) );
NAND3_X1 U734 ( .A1(n1020), .A2(n1014), .A3(n1015), .ZN(n1018) );
NAND2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U736 ( .A1(n1010), .A2(n1023), .ZN(n1022) );
NAND3_X1 U737 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1021) );
OR2_X1 U738 ( .A1(n1027), .A2(n1010), .ZN(n1025) );
NAND3_X1 U739 ( .A1(n1028), .A2(n1029), .A3(n1027), .ZN(n1024) );
NAND3_X1 U740 ( .A1(n1030), .A2(n1027), .A3(n1010), .ZN(n1002) );
NAND2_X1 U741 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND4_X1 U742 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
NOR2_X1 U743 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
XOR2_X1 U744 ( .A(n1039), .B(KEYINPUT33), .Z(n1038) );
XNOR2_X1 U745 ( .A(n1040), .B(n1041), .ZN(n1034) );
NAND2_X1 U746 ( .A1(KEYINPUT30), .A2(n1042), .ZN(n1040) );
XOR2_X1 U747 ( .A(n1043), .B(n1044), .Z(n1033) );
XOR2_X1 U748 ( .A(KEYINPUT38), .B(G469), .Z(n1044) );
NAND2_X1 U749 ( .A1(KEYINPUT17), .A2(n1045), .ZN(n1043) );
NAND4_X1 U750 ( .A1(n1046), .A2(n1011), .A3(n1026), .A4(n1015), .ZN(n1031) );
INV_X1 U751 ( .A(n1019), .ZN(n1011) );
XNOR2_X1 U752 ( .A(n1047), .B(KEYINPUT9), .ZN(n1046) );
XOR2_X1 U753 ( .A(n1048), .B(n1049), .Z(G72) );
XOR2_X1 U754 ( .A(n1050), .B(n1051), .Z(n1049) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
AND2_X1 U756 ( .A1(G227), .A2(G900), .ZN(n1052) );
NAND3_X1 U757 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1050) );
XOR2_X1 U758 ( .A(n1057), .B(KEYINPUT50), .Z(n1056) );
OR2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U760 ( .A1(G953), .A2(n1060), .ZN(n1055) );
NAND2_X1 U761 ( .A1(n1059), .A2(n1058), .ZN(n1054) );
XNOR2_X1 U762 ( .A(n1061), .B(n1062), .ZN(n1058) );
XOR2_X1 U763 ( .A(n1063), .B(n1064), .Z(n1062) );
NOR2_X1 U764 ( .A1(KEYINPUT34), .A2(n1065), .ZN(n1063) );
XOR2_X1 U765 ( .A(n1066), .B(n1067), .Z(n1061) );
NOR2_X1 U766 ( .A1(KEYINPUT4), .A2(n1068), .ZN(n1067) );
INV_X1 U767 ( .A(n1069), .ZN(n1068) );
XNOR2_X1 U768 ( .A(G131), .B(KEYINPUT3), .ZN(n1066) );
NAND2_X1 U769 ( .A1(n1053), .A2(n1070), .ZN(n1048) );
XOR2_X1 U770 ( .A(n1071), .B(n1072), .Z(G69) );
NOR2_X1 U771 ( .A1(n1073), .A2(n1053), .ZN(n1072) );
AND2_X1 U772 ( .A1(G224), .A2(G898), .ZN(n1073) );
NAND2_X1 U773 ( .A1(n1074), .A2(KEYINPUT63), .ZN(n1071) );
XOR2_X1 U774 ( .A(n1075), .B(n1076), .Z(n1074) );
AND2_X1 U775 ( .A1(n1077), .A2(n1053), .ZN(n1076) );
NAND2_X1 U776 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
NAND2_X1 U777 ( .A1(G953), .A2(n1080), .ZN(n1079) );
XOR2_X1 U778 ( .A(n1081), .B(n1082), .Z(n1078) );
XOR2_X1 U779 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U780 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U781 ( .A1(KEYINPUT27), .A2(n1087), .ZN(n1085) );
XOR2_X1 U782 ( .A(n1088), .B(G110), .Z(n1081) );
XNOR2_X1 U783 ( .A(KEYINPUT51), .B(KEYINPUT37), .ZN(n1088) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(G66) );
XOR2_X1 U785 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U786 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
XNOR2_X1 U787 ( .A(KEYINPUT7), .B(n1095), .ZN(n1094) );
NOR4_X1 U788 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(G63) );
NOR3_X1 U789 ( .A1(n1100), .A2(G953), .A3(G952), .ZN(n1099) );
AND2_X1 U790 ( .A1(n1100), .A2(n1089), .ZN(n1098) );
INV_X1 U791 ( .A(KEYINPUT21), .ZN(n1100) );
NOR4_X1 U792 ( .A1(n1101), .A2(n1102), .A3(KEYINPUT36), .A4(n1103), .ZN(n1097) );
INV_X1 U793 ( .A(n1104), .ZN(n1101) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1096) );
NOR3_X1 U795 ( .A1(n1102), .A2(n1106), .A3(n1103), .ZN(n1105) );
AND2_X1 U796 ( .A1(n1107), .A2(KEYINPUT36), .ZN(n1106) );
NOR2_X1 U797 ( .A1(KEYINPUT13), .A2(n1107), .ZN(n1104) );
NOR2_X1 U798 ( .A1(n1089), .A2(n1108), .ZN(G60) );
XOR2_X1 U799 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U800 ( .A1(n1093), .A2(G475), .ZN(n1109) );
NAND3_X1 U801 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(G6) );
NAND2_X1 U802 ( .A1(G104), .A2(n1114), .ZN(n1113) );
NAND2_X1 U803 ( .A1(KEYINPUT20), .A2(n1115), .ZN(n1112) );
NAND2_X1 U804 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
INV_X1 U805 ( .A(n1114), .ZN(n1117) );
XNOR2_X1 U806 ( .A(KEYINPUT61), .B(G104), .ZN(n1116) );
NAND2_X1 U807 ( .A1(n1118), .A2(n1119), .ZN(n1111) );
INV_X1 U808 ( .A(KEYINPUT20), .ZN(n1119) );
NAND2_X1 U809 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
OR3_X1 U810 ( .A1(n1114), .A2(G104), .A3(KEYINPUT61), .ZN(n1121) );
NAND2_X1 U811 ( .A1(KEYINPUT61), .A2(G104), .ZN(n1120) );
NOR2_X1 U812 ( .A1(n1089), .A2(n1122), .ZN(G57) );
XOR2_X1 U813 ( .A(n1123), .B(n1124), .Z(n1122) );
XNOR2_X1 U814 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR3_X1 U815 ( .A1(n1102), .A2(KEYINPUT41), .A3(n1127), .ZN(n1126) );
INV_X1 U816 ( .A(n1093), .ZN(n1102) );
XOR2_X1 U817 ( .A(n1128), .B(n1129), .Z(n1123) );
NAND2_X1 U818 ( .A1(KEYINPUT15), .A2(n1130), .ZN(n1128) );
NOR2_X1 U819 ( .A1(n1089), .A2(n1131), .ZN(G54) );
XOR2_X1 U820 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U821 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U822 ( .A1(KEYINPUT56), .A2(n1136), .ZN(n1135) );
NAND2_X1 U823 ( .A1(n1093), .A2(G469), .ZN(n1134) );
NOR2_X1 U824 ( .A1(n1089), .A2(n1137), .ZN(G51) );
XOR2_X1 U825 ( .A(n1138), .B(n1139), .Z(n1137) );
XNOR2_X1 U826 ( .A(n1140), .B(n1069), .ZN(n1139) );
NAND2_X1 U827 ( .A1(n1093), .A2(n1042), .ZN(n1140) );
NOR2_X1 U828 ( .A1(n1141), .A2(n1001), .ZN(n1093) );
NOR2_X1 U829 ( .A1(n1077), .A2(n1070), .ZN(n1001) );
NAND4_X1 U830 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1070) );
NOR4_X1 U831 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
NAND2_X1 U832 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
NAND2_X1 U833 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U834 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XNOR2_X1 U835 ( .A(n1156), .B(KEYINPUT40), .ZN(n1154) );
NAND2_X1 U836 ( .A1(n1010), .A2(n1157), .ZN(n1152) );
NAND2_X1 U837 ( .A1(n1158), .A2(n1159), .ZN(n1077) );
AND4_X1 U838 ( .A1(n999), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1159) );
NAND3_X1 U839 ( .A1(n1015), .A2(n1163), .A3(n1164), .ZN(n999) );
AND4_X1 U840 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1114), .ZN(n1158) );
NAND3_X1 U841 ( .A1(n1164), .A2(n1015), .A3(n1155), .ZN(n1114) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1138) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U844 ( .A1(G125), .A2(KEYINPUT5), .ZN(n1171) );
NAND2_X1 U845 ( .A1(KEYINPUT59), .A2(n1172), .ZN(n1168) );
NOR2_X1 U846 ( .A1(n1053), .A2(G952), .ZN(n1089) );
XNOR2_X1 U847 ( .A(G146), .B(n1142), .ZN(G48) );
NAND3_X1 U848 ( .A1(n1155), .A2(n1157), .A3(n1173), .ZN(n1142) );
XNOR2_X1 U849 ( .A(G143), .B(n1143), .ZN(G45) );
NAND4_X1 U850 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1143) );
XNOR2_X1 U851 ( .A(n1177), .B(n1178), .ZN(G42) );
NOR3_X1 U852 ( .A1(n1179), .A2(n1017), .A3(n1028), .ZN(n1178) );
INV_X1 U853 ( .A(n1156), .ZN(n1017) );
XNOR2_X1 U854 ( .A(G137), .B(n1180), .ZN(G39) );
NAND4_X1 U855 ( .A1(KEYINPUT57), .A2(n1150), .A3(n1010), .A4(n1157), .ZN(n1180) );
INV_X1 U856 ( .A(n1179), .ZN(n1150) );
XNOR2_X1 U857 ( .A(n1181), .B(n1149), .ZN(G36) );
NOR3_X1 U858 ( .A1(n1029), .A2(n1016), .A3(n1179), .ZN(n1149) );
INV_X1 U859 ( .A(n1163), .ZN(n1029) );
XNOR2_X1 U860 ( .A(n1182), .B(n1148), .ZN(G33) );
NOR3_X1 U861 ( .A1(n1028), .A2(n1016), .A3(n1179), .ZN(n1148) );
NAND4_X1 U862 ( .A1(n1183), .A2(n1023), .A3(n1014), .A4(n1184), .ZN(n1179) );
INV_X1 U863 ( .A(n1174), .ZN(n1016) );
XOR2_X1 U864 ( .A(G128), .B(n1147), .Z(G30) );
AND3_X1 U865 ( .A1(n1163), .A2(n1157), .A3(n1173), .ZN(n1147) );
AND3_X1 U866 ( .A1(n1047), .A2(n1184), .A3(n1023), .ZN(n1173) );
XNOR2_X1 U867 ( .A(G101), .B(n1167), .ZN(G3) );
NAND3_X1 U868 ( .A1(n1164), .A2(n1174), .A3(n1010), .ZN(n1167) );
XOR2_X1 U869 ( .A(n1146), .B(n1185), .Z(G27) );
NOR2_X1 U870 ( .A1(KEYINPUT31), .A2(n1186), .ZN(n1185) );
AND4_X1 U871 ( .A1(n1026), .A2(n1156), .A3(n1155), .A4(n1187), .ZN(n1146) );
AND3_X1 U872 ( .A1(n1047), .A2(n1184), .A3(n1027), .ZN(n1187) );
NAND2_X1 U873 ( .A1(n1188), .A2(n1019), .ZN(n1184) );
NAND2_X1 U874 ( .A1(n1189), .A2(n1060), .ZN(n1188) );
XOR2_X1 U875 ( .A(KEYINPUT10), .B(G900), .Z(n1060) );
XNOR2_X1 U876 ( .A(G122), .B(n1166), .ZN(G24) );
NAND4_X1 U877 ( .A1(n1190), .A2(n1015), .A3(n1175), .A4(n1176), .ZN(n1166) );
XNOR2_X1 U878 ( .A(G119), .B(n1165), .ZN(G21) );
NAND3_X1 U879 ( .A1(n1010), .A2(n1157), .A3(n1190), .ZN(n1165) );
NAND2_X1 U880 ( .A1(n1191), .A2(n1192), .ZN(n1157) );
NAND2_X1 U881 ( .A1(n1156), .A2(n1193), .ZN(n1192) );
NAND3_X1 U882 ( .A1(n1194), .A2(n1195), .A3(KEYINPUT42), .ZN(n1191) );
NAND2_X1 U883 ( .A1(n1196), .A2(n1197), .ZN(G18) );
OR2_X1 U884 ( .A1(n1162), .A2(G116), .ZN(n1197) );
XOR2_X1 U885 ( .A(n1198), .B(KEYINPUT24), .Z(n1196) );
NAND2_X1 U886 ( .A1(G116), .A2(n1162), .ZN(n1198) );
NAND3_X1 U887 ( .A1(n1163), .A2(n1174), .A3(n1190), .ZN(n1162) );
NOR2_X1 U888 ( .A1(n1175), .A2(n1199), .ZN(n1163) );
XNOR2_X1 U889 ( .A(G113), .B(n1161), .ZN(G15) );
NAND3_X1 U890 ( .A1(n1155), .A2(n1174), .A3(n1190), .ZN(n1161) );
AND3_X1 U891 ( .A1(n1200), .A2(n1027), .A3(n1026), .ZN(n1190) );
NAND2_X1 U892 ( .A1(n1201), .A2(n1202), .ZN(n1174) );
NAND2_X1 U893 ( .A1(n1015), .A2(n1193), .ZN(n1202) );
INV_X1 U894 ( .A(KEYINPUT42), .ZN(n1193) );
NOR2_X1 U895 ( .A1(n1194), .A2(n1195), .ZN(n1015) );
NAND3_X1 U896 ( .A1(n1036), .A2(n1195), .A3(KEYINPUT42), .ZN(n1201) );
INV_X1 U897 ( .A(n1028), .ZN(n1155) );
NAND2_X1 U898 ( .A1(n1199), .A2(n1175), .ZN(n1028) );
INV_X1 U899 ( .A(n1176), .ZN(n1199) );
XOR2_X1 U900 ( .A(n1160), .B(n1203), .Z(G12) );
XOR2_X1 U901 ( .A(KEYINPUT60), .B(G110), .Z(n1203) );
NAND3_X1 U902 ( .A1(n1010), .A2(n1164), .A3(n1156), .ZN(n1160) );
NOR2_X1 U903 ( .A1(n1036), .A2(n1195), .ZN(n1156) );
XOR2_X1 U904 ( .A(n1039), .B(KEYINPUT19), .Z(n1195) );
XNOR2_X1 U905 ( .A(n1204), .B(n1127), .ZN(n1039) );
INV_X1 U906 ( .A(G472), .ZN(n1127) );
NAND2_X1 U907 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XNOR2_X1 U908 ( .A(n1129), .B(n1207), .ZN(n1205) );
XOR2_X1 U909 ( .A(KEYINPUT46), .B(n1208), .Z(n1207) );
NOR2_X1 U910 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U911 ( .A(n1211), .B(KEYINPUT45), .Z(n1210) );
NAND2_X1 U912 ( .A1(n1130), .A2(G101), .ZN(n1211) );
NOR2_X1 U913 ( .A1(G101), .A2(n1130), .ZN(n1209) );
AND3_X1 U914 ( .A1(n1212), .A2(n1053), .A3(G210), .ZN(n1130) );
XNOR2_X1 U915 ( .A(n1213), .B(n1214), .ZN(n1129) );
XNOR2_X1 U916 ( .A(G119), .B(n1215), .ZN(n1214) );
XNOR2_X1 U917 ( .A(n1216), .B(n1217), .ZN(n1213) );
INV_X1 U918 ( .A(n1194), .ZN(n1036) );
XNOR2_X1 U919 ( .A(n1218), .B(n1219), .ZN(n1194) );
NOR2_X1 U920 ( .A1(n1220), .A2(n1095), .ZN(n1219) );
INV_X1 U921 ( .A(G217), .ZN(n1095) );
NOR2_X1 U922 ( .A1(G902), .A2(n1221), .ZN(n1220) );
NAND2_X1 U923 ( .A1(n1206), .A2(n1092), .ZN(n1218) );
XNOR2_X1 U924 ( .A(n1222), .B(n1223), .ZN(n1092) );
XOR2_X1 U925 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U926 ( .A(n1226), .B(n1227), .ZN(n1225) );
NAND2_X1 U927 ( .A1(KEYINPUT1), .A2(n1065), .ZN(n1227) );
NAND2_X1 U928 ( .A1(KEYINPUT53), .A2(n1177), .ZN(n1226) );
XNOR2_X1 U929 ( .A(G110), .B(G125), .ZN(n1224) );
XOR2_X1 U930 ( .A(n1228), .B(n1229), .Z(n1222) );
XNOR2_X1 U931 ( .A(n1230), .B(n1231), .ZN(n1229) );
NOR2_X1 U932 ( .A1(G146), .A2(KEYINPUT26), .ZN(n1230) );
XOR2_X1 U933 ( .A(n1232), .B(n1233), .Z(n1228) );
NOR2_X1 U934 ( .A1(G119), .A2(KEYINPUT47), .ZN(n1233) );
NAND2_X1 U935 ( .A1(n1234), .A2(G221), .ZN(n1232) );
AND2_X1 U936 ( .A1(n1023), .A2(n1200), .ZN(n1164) );
AND2_X1 U937 ( .A1(n1047), .A2(n1235), .ZN(n1200) );
NAND2_X1 U938 ( .A1(n1236), .A2(n1019), .ZN(n1235) );
NAND3_X1 U939 ( .A1(n1237), .A2(n1053), .A3(G952), .ZN(n1019) );
NAND2_X1 U940 ( .A1(n1189), .A2(n1080), .ZN(n1236) );
XOR2_X1 U941 ( .A(KEYINPUT54), .B(G898), .Z(n1080) );
AND3_X1 U942 ( .A1(n1238), .A2(n1237), .A3(G953), .ZN(n1189) );
NAND2_X1 U943 ( .A1(G237), .A2(G234), .ZN(n1237) );
XNOR2_X1 U944 ( .A(KEYINPUT62), .B(n1141), .ZN(n1238) );
NOR2_X1 U945 ( .A1(n1183), .A2(n1037), .ZN(n1047) );
INV_X1 U946 ( .A(n1014), .ZN(n1037) );
NAND2_X1 U947 ( .A1(G214), .A2(n1239), .ZN(n1014) );
INV_X1 U948 ( .A(n1009), .ZN(n1183) );
XNOR2_X1 U949 ( .A(n1041), .B(n1042), .ZN(n1009) );
AND2_X1 U950 ( .A1(G210), .A2(n1239), .ZN(n1042) );
NAND2_X1 U951 ( .A1(n1212), .A2(n1141), .ZN(n1239) );
NAND2_X1 U952 ( .A1(n1206), .A2(n1240), .ZN(n1041) );
XOR2_X1 U953 ( .A(n1241), .B(n1242), .Z(n1240) );
XNOR2_X1 U954 ( .A(n1243), .B(n1170), .ZN(n1242) );
NAND2_X1 U955 ( .A1(n1244), .A2(n1245), .ZN(n1170) );
NAND2_X1 U956 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U957 ( .A(KEYINPUT44), .B(n1248), .Z(n1244) );
NOR2_X1 U958 ( .A1(n1246), .A2(n1247), .ZN(n1248) );
XOR2_X1 U959 ( .A(n1249), .B(n1087), .Z(n1247) );
AND2_X1 U960 ( .A1(n1250), .A2(n1251), .ZN(n1087) );
NAND2_X1 U961 ( .A1(n1252), .A2(n1217), .ZN(n1251) );
XNOR2_X1 U962 ( .A(n1215), .B(n1253), .ZN(n1252) );
NAND2_X1 U963 ( .A1(G113), .A2(n1254), .ZN(n1250) );
XNOR2_X1 U964 ( .A(G116), .B(n1253), .ZN(n1254) );
NOR2_X1 U965 ( .A1(G119), .A2(KEYINPUT25), .ZN(n1253) );
XNOR2_X1 U966 ( .A(n1083), .B(n1255), .ZN(n1249) );
XNOR2_X1 U967 ( .A(n1256), .B(n1257), .ZN(n1083) );
NAND2_X1 U968 ( .A1(KEYINPUT29), .A2(n1125), .ZN(n1256) );
INV_X1 U969 ( .A(G101), .ZN(n1125) );
XOR2_X1 U970 ( .A(G110), .B(n1258), .Z(n1246) );
XNOR2_X1 U971 ( .A(KEYINPUT0), .B(n1259), .ZN(n1258) );
NAND2_X1 U972 ( .A1(KEYINPUT11), .A2(n1069), .ZN(n1243) );
XNOR2_X1 U973 ( .A(G125), .B(n1172), .ZN(n1241) );
AND2_X1 U974 ( .A1(G224), .A2(n1053), .ZN(n1172) );
NOR2_X1 U975 ( .A1(n1026), .A2(n1008), .ZN(n1023) );
INV_X1 U976 ( .A(n1027), .ZN(n1008) );
NAND2_X1 U977 ( .A1(G221), .A2(n1260), .ZN(n1027) );
NAND2_X1 U978 ( .A1(G234), .A2(n1141), .ZN(n1260) );
INV_X1 U979 ( .A(G902), .ZN(n1141) );
INV_X1 U980 ( .A(n1007), .ZN(n1026) );
XNOR2_X1 U981 ( .A(n1045), .B(G469), .ZN(n1007) );
NAND2_X1 U982 ( .A1(n1261), .A2(n1206), .ZN(n1045) );
XOR2_X1 U983 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U984 ( .A(KEYINPUT58), .B(KEYINPUT49), .Z(n1263) );
XNOR2_X1 U985 ( .A(n1264), .B(n1136), .ZN(n1262) );
XOR2_X1 U986 ( .A(n1265), .B(n1266), .Z(n1136) );
XOR2_X1 U987 ( .A(G110), .B(n1267), .Z(n1266) );
AND2_X1 U988 ( .A1(n1053), .A2(G227), .ZN(n1267) );
XNOR2_X1 U989 ( .A(G140), .B(KEYINPUT28), .ZN(n1265) );
NAND2_X1 U990 ( .A1(n1268), .A2(KEYINPUT43), .ZN(n1264) );
XOR2_X1 U991 ( .A(n1132), .B(KEYINPUT16), .Z(n1268) );
XOR2_X1 U992 ( .A(n1216), .B(n1269), .Z(n1132) );
XNOR2_X1 U993 ( .A(G101), .B(n1270), .ZN(n1269) );
NAND3_X1 U994 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1270) );
NAND2_X1 U995 ( .A1(KEYINPUT23), .A2(G104), .ZN(n1273) );
NAND3_X1 U996 ( .A1(n1255), .A2(n1274), .A3(G107), .ZN(n1272) );
NAND2_X1 U997 ( .A1(n1275), .A2(n1257), .ZN(n1271) );
NAND2_X1 U998 ( .A1(n1276), .A2(n1274), .ZN(n1275) );
INV_X1 U999 ( .A(KEYINPUT23), .ZN(n1274) );
XNOR2_X1 U1000 ( .A(KEYINPUT52), .B(n1255), .ZN(n1276) );
XOR2_X1 U1001 ( .A(n1277), .B(n1278), .Z(n1216) );
XNOR2_X1 U1002 ( .A(n1065), .B(G131), .ZN(n1278) );
INV_X1 U1003 ( .A(G137), .ZN(n1065) );
XNOR2_X1 U1004 ( .A(n1069), .B(n1064), .ZN(n1277) );
XNOR2_X1 U1005 ( .A(n1181), .B(KEYINPUT55), .ZN(n1064) );
INV_X1 U1006 ( .A(G134), .ZN(n1181) );
XOR2_X1 U1007 ( .A(n1279), .B(n1280), .Z(n1069) );
XNOR2_X1 U1008 ( .A(G146), .B(n1231), .ZN(n1280) );
NOR2_X1 U1009 ( .A1(n1176), .A2(n1175), .ZN(n1010) );
XNOR2_X1 U1010 ( .A(n1281), .B(G475), .ZN(n1175) );
NAND2_X1 U1011 ( .A1(n1110), .A2(n1206), .ZN(n1281) );
XNOR2_X1 U1012 ( .A(n1086), .B(n1282), .ZN(n1110) );
XNOR2_X1 U1013 ( .A(n1217), .B(n1283), .ZN(n1282) );
NOR2_X1 U1014 ( .A1(KEYINPUT18), .A2(n1284), .ZN(n1283) );
XOR2_X1 U1015 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U1016 ( .A(n1287), .B(n1059), .ZN(n1286) );
XNOR2_X1 U1017 ( .A(n1186), .B(n1177), .ZN(n1059) );
INV_X1 U1018 ( .A(G140), .ZN(n1177) );
INV_X1 U1019 ( .A(G125), .ZN(n1186) );
AND3_X1 U1020 ( .A1(G214), .A2(n1053), .A3(n1212), .ZN(n1287) );
INV_X1 U1021 ( .A(G237), .ZN(n1212) );
INV_X1 U1022 ( .A(G953), .ZN(n1053) );
XOR2_X1 U1023 ( .A(n1288), .B(n1289), .Z(n1285) );
XNOR2_X1 U1024 ( .A(G146), .B(n1182), .ZN(n1289) );
INV_X1 U1025 ( .A(G131), .ZN(n1182) );
NAND2_X1 U1026 ( .A1(KEYINPUT22), .A2(n1279), .ZN(n1288) );
INV_X1 U1027 ( .A(G113), .ZN(n1217) );
XNOR2_X1 U1028 ( .A(G122), .B(n1255), .ZN(n1086) );
INV_X1 U1029 ( .A(G104), .ZN(n1255) );
XOR2_X1 U1030 ( .A(n1290), .B(n1103), .Z(n1176) );
INV_X1 U1031 ( .A(G478), .ZN(n1103) );
NAND2_X1 U1032 ( .A1(n1291), .A2(n1206), .ZN(n1290) );
XNOR2_X1 U1033 ( .A(G902), .B(KEYINPUT12), .ZN(n1206) );
INV_X1 U1034 ( .A(n1107), .ZN(n1291) );
XNOR2_X1 U1035 ( .A(n1292), .B(n1293), .ZN(n1107) );
AND2_X1 U1036 ( .A1(G217), .A2(n1234), .ZN(n1293) );
NOR2_X1 U1037 ( .A1(n1221), .A2(G953), .ZN(n1234) );
INV_X1 U1038 ( .A(G234), .ZN(n1221) );
NAND2_X1 U1039 ( .A1(n1294), .A2(KEYINPUT8), .ZN(n1292) );
XOR2_X1 U1040 ( .A(n1295), .B(n1296), .Z(n1294) );
NOR2_X1 U1041 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U1042 ( .A(n1299), .B(KEYINPUT32), .Z(n1298) );
NAND2_X1 U1043 ( .A1(n1231), .A2(n1300), .ZN(n1299) );
NOR2_X1 U1044 ( .A1(n1231), .A2(n1300), .ZN(n1297) );
INV_X1 U1045 ( .A(n1279), .ZN(n1300) );
XOR2_X1 U1046 ( .A(G143), .B(KEYINPUT6), .Z(n1279) );
XNOR2_X1 U1047 ( .A(G128), .B(KEYINPUT14), .ZN(n1231) );
XNOR2_X1 U1048 ( .A(G134), .B(n1301), .ZN(n1295) );
NOR2_X1 U1049 ( .A1(KEYINPUT48), .A2(n1302), .ZN(n1301) );
XNOR2_X1 U1050 ( .A(n1257), .B(n1303), .ZN(n1302) );
NOR2_X1 U1051 ( .A1(KEYINPUT35), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U1052 ( .A(n1215), .B(n1305), .ZN(n1304) );
XNOR2_X1 U1053 ( .A(KEYINPUT2), .B(n1259), .ZN(n1305) );
INV_X1 U1054 ( .A(G122), .ZN(n1259) );
INV_X1 U1055 ( .A(G116), .ZN(n1215) );
INV_X1 U1056 ( .A(G107), .ZN(n1257) );
endmodule


