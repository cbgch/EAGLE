//Key = 0100100100100110010101010001010011000010111100100110111011111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369;

XOR2_X1 U747 ( .A(G107), .B(n1040), .Z(G9) );
NOR2_X1 U748 ( .A1(KEYINPUT39), .A2(n1041), .ZN(n1040) );
NOR2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U750 ( .A1(G953), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1043) );
NOR2_X1 U751 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U753 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
INV_X1 U754 ( .A(n1053), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1051) );
NOR4_X1 U756 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
NOR3_X1 U757 ( .A1(n1060), .A2(KEYINPUT63), .A3(n1061), .ZN(n1057) );
NOR2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1056) );
NOR2_X1 U759 ( .A1(KEYINPUT63), .A2(n1061), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1054) );
NOR2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U762 ( .A1(n1068), .A2(n1058), .ZN(n1067) );
NOR2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U764 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U765 ( .A1(n1073), .A2(n1059), .ZN(n1066) );
NOR2_X1 U766 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR4_X1 U767 ( .A1(n1076), .A2(n1058), .A3(n1059), .A4(n1065), .ZN(n1049) );
INV_X1 U768 ( .A(n1077), .ZN(n1065) );
INV_X1 U769 ( .A(n1078), .ZN(n1058) );
NOR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1076) );
NOR3_X1 U771 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n1042) );
AND4_X1 U772 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1044) );
NOR4_X1 U773 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
XNOR2_X1 U774 ( .A(n1089), .B(n1090), .ZN(n1088) );
NAND2_X1 U775 ( .A1(KEYINPUT38), .A2(n1091), .ZN(n1089) );
NOR2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1087) );
NOR2_X1 U777 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
INV_X1 U778 ( .A(n1096), .ZN(n1095) );
NOR2_X1 U779 ( .A1(KEYINPUT16), .A2(n1097), .ZN(n1094) );
NOR2_X1 U780 ( .A1(KEYINPUT6), .A2(n1098), .ZN(n1097) );
NOR2_X1 U781 ( .A1(G478), .A2(n1099), .ZN(n1092) );
NOR2_X1 U782 ( .A1(n1100), .A2(KEYINPUT6), .ZN(n1099) );
NOR2_X1 U783 ( .A1(KEYINPUT16), .A2(n1096), .ZN(n1100) );
XNOR2_X1 U784 ( .A(n1101), .B(KEYINPUT45), .ZN(n1096) );
NOR3_X1 U785 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1086) );
NOR2_X1 U786 ( .A1(KEYINPUT1), .A2(n1105), .ZN(n1104) );
AND4_X1 U787 ( .A1(n1105), .A2(KEYINPUT21), .A3(n1106), .A4(KEYINPUT1), .ZN(n1103) );
NOR2_X1 U788 ( .A1(n1107), .A2(n1106), .ZN(n1102) );
AND2_X1 U789 ( .A1(n1105), .A2(KEYINPUT21), .ZN(n1107) );
XNOR2_X1 U790 ( .A(n1108), .B(n1109), .ZN(n1083) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(G72) );
NAND2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U793 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
XOR2_X1 U794 ( .A(n1117), .B(KEYINPUT22), .Z(n1114) );
OR2_X1 U795 ( .A1(n1117), .A2(n1116), .ZN(n1112) );
XOR2_X1 U796 ( .A(n1118), .B(n1119), .Z(n1116) );
XOR2_X1 U797 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U798 ( .A(G131), .B(G137), .ZN(n1121) );
NAND2_X1 U799 ( .A1(n1122), .A2(KEYINPUT42), .ZN(n1120) );
XNOR2_X1 U800 ( .A(G134), .B(KEYINPUT5), .ZN(n1122) );
XOR2_X1 U801 ( .A(n1123), .B(n1124), .Z(n1118) );
NOR3_X1 U802 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
NOR2_X1 U803 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
AND3_X1 U804 ( .A1(n1129), .A2(n1128), .A3(KEYINPUT41), .ZN(n1126) );
AND2_X1 U805 ( .A1(KEYINPUT52), .A2(n1130), .ZN(n1128) );
NOR2_X1 U806 ( .A1(KEYINPUT41), .A2(n1130), .ZN(n1125) );
NAND2_X1 U807 ( .A1(n1131), .A2(n1132), .ZN(n1117) );
NAND2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U809 ( .A1(n1115), .A2(n1135), .ZN(n1110) );
OR2_X1 U810 ( .A1(n1131), .A2(G227), .ZN(n1135) );
INV_X1 U811 ( .A(n1136), .ZN(n1115) );
NAND3_X1 U812 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(G69) );
NAND2_X1 U813 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
OR3_X1 U814 ( .A1(n1140), .A2(n1141), .A3(G953), .ZN(n1138) );
NAND2_X1 U815 ( .A1(n1142), .A2(G953), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U817 ( .A1(n1140), .A2(n1145), .ZN(n1144) );
NAND2_X1 U818 ( .A1(G224), .A2(n1146), .ZN(n1143) );
NAND2_X1 U819 ( .A1(G898), .A2(n1140), .ZN(n1146) );
NAND3_X1 U820 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1140) );
XOR2_X1 U821 ( .A(n1150), .B(KEYINPUT12), .Z(n1149) );
NAND2_X1 U822 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
OR2_X1 U823 ( .A1(n1152), .A2(n1151), .ZN(n1148) );
XNOR2_X1 U824 ( .A(n1153), .B(KEYINPUT43), .ZN(n1152) );
NAND2_X1 U825 ( .A1(G953), .A2(n1154), .ZN(n1147) );
NOR2_X1 U826 ( .A1(n1155), .A2(n1156), .ZN(G66) );
NOR3_X1 U827 ( .A1(n1108), .A2(n1157), .A3(n1158), .ZN(n1156) );
NOR3_X1 U828 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
NOR2_X1 U829 ( .A1(n1162), .A2(n1163), .ZN(n1157) );
AND2_X1 U830 ( .A1(n1046), .A2(G217), .ZN(n1162) );
NOR2_X1 U831 ( .A1(n1155), .A2(n1164), .ZN(G63) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U833 ( .A(n1167), .B(KEYINPUT19), .ZN(n1166) );
NAND2_X1 U834 ( .A1(KEYINPUT29), .A2(n1168), .ZN(n1167) );
NOR2_X1 U835 ( .A1(n1098), .A2(n1161), .ZN(n1165) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1169), .ZN(G60) );
XNOR2_X1 U837 ( .A(n1170), .B(n1171), .ZN(n1169) );
NAND2_X1 U838 ( .A1(KEYINPUT7), .A2(n1172), .ZN(n1170) );
NAND2_X1 U839 ( .A1(n1173), .A2(G475), .ZN(n1172) );
XNOR2_X1 U840 ( .A(G104), .B(n1174), .ZN(G6) );
NOR2_X1 U841 ( .A1(n1155), .A2(n1175), .ZN(G57) );
XNOR2_X1 U842 ( .A(n1176), .B(n1177), .ZN(n1175) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
AND3_X1 U844 ( .A1(n1180), .A2(G472), .A3(n1173), .ZN(n1179) );
INV_X1 U845 ( .A(n1161), .ZN(n1173) );
NOR2_X1 U846 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
XOR2_X1 U847 ( .A(KEYINPUT62), .B(n1182), .Z(n1181) );
NOR2_X1 U848 ( .A1(n1106), .A2(n1161), .ZN(n1182) );
XNOR2_X1 U849 ( .A(n1183), .B(n1184), .ZN(n1180) );
NOR2_X1 U850 ( .A1(KEYINPUT35), .A2(n1185), .ZN(n1184) );
NOR2_X1 U851 ( .A1(n1155), .A2(n1186), .ZN(G54) );
XOR2_X1 U852 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U853 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U854 ( .A1(n1091), .A2(n1161), .ZN(n1189) );
XOR2_X1 U855 ( .A(n1191), .B(n1192), .Z(n1187) );
XOR2_X1 U856 ( .A(KEYINPUT34), .B(n1193), .Z(n1192) );
NOR4_X1 U857 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NOR2_X1 U858 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR3_X1 U859 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1195) );
NOR2_X1 U860 ( .A1(n1129), .A2(n1198), .ZN(n1202) );
INV_X1 U861 ( .A(KEYINPUT27), .ZN(n1198) );
NOR3_X1 U862 ( .A1(G110), .A2(KEYINPUT27), .A3(n1203), .ZN(n1194) );
NOR2_X1 U863 ( .A1(KEYINPUT28), .A2(n1204), .ZN(n1191) );
NOR2_X1 U864 ( .A1(n1155), .A2(n1205), .ZN(G51) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U866 ( .A(n1185), .B(n1208), .ZN(n1207) );
XOR2_X1 U867 ( .A(n1209), .B(n1210), .Z(n1206) );
NOR2_X1 U868 ( .A1(n1211), .A2(n1161), .ZN(n1210) );
NAND2_X1 U869 ( .A1(G902), .A2(n1046), .ZN(n1161) );
NAND3_X1 U870 ( .A1(n1212), .A2(n1133), .A3(n1213), .ZN(n1046) );
XNOR2_X1 U871 ( .A(n1134), .B(KEYINPUT61), .ZN(n1213) );
AND4_X1 U872 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1134) );
AND4_X1 U873 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1133) );
INV_X1 U874 ( .A(n1141), .ZN(n1212) );
NAND4_X1 U875 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1141) );
AND4_X1 U876 ( .A1(n1174), .A2(n1041), .A3(n1226), .A4(n1227), .ZN(n1225) );
NAND4_X1 U877 ( .A1(n1079), .A2(n1078), .A3(n1070), .A4(n1228), .ZN(n1041) );
NAND4_X1 U878 ( .A1(n1080), .A2(n1078), .A3(n1070), .A4(n1228), .ZN(n1174) );
NOR2_X1 U879 ( .A1(n1229), .A2(n1230), .ZN(n1224) );
NOR2_X1 U880 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U881 ( .A1(KEYINPUT10), .A2(n1233), .ZN(n1209) );
NOR2_X1 U882 ( .A1(n1131), .A2(G952), .ZN(n1155) );
XNOR2_X1 U883 ( .A(G146), .B(n1234), .ZN(G48) );
NAND2_X1 U884 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND2_X1 U885 ( .A1(KEYINPUT49), .A2(n1218), .ZN(n1236) );
NAND2_X1 U886 ( .A1(KEYINPUT44), .A2(n1237), .ZN(n1235) );
INV_X1 U887 ( .A(n1218), .ZN(n1237) );
NAND3_X1 U888 ( .A1(n1080), .A2(n1070), .A3(n1238), .ZN(n1218) );
XOR2_X1 U889 ( .A(G143), .B(n1239), .Z(G45) );
NOR2_X1 U890 ( .A1(KEYINPUT48), .A2(n1219), .ZN(n1239) );
NAND3_X1 U891 ( .A1(n1240), .A2(n1074), .A3(n1241), .ZN(n1219) );
NOR3_X1 U892 ( .A1(n1231), .A2(n1242), .A3(n1243), .ZN(n1241) );
XNOR2_X1 U893 ( .A(G140), .B(n1220), .ZN(G42) );
NAND2_X1 U894 ( .A1(n1244), .A2(n1075), .ZN(n1220) );
XNOR2_X1 U895 ( .A(G137), .B(n1221), .ZN(G39) );
NAND3_X1 U896 ( .A1(n1053), .A2(n1082), .A3(n1238), .ZN(n1221) );
XNOR2_X1 U897 ( .A(G134), .B(n1215), .ZN(G36) );
NAND4_X1 U898 ( .A1(n1240), .A2(n1074), .A3(n1082), .A4(n1079), .ZN(n1215) );
XNOR2_X1 U899 ( .A(n1216), .B(n1245), .ZN(G33) );
NOR2_X1 U900 ( .A1(KEYINPUT51), .A2(n1246), .ZN(n1245) );
NAND2_X1 U901 ( .A1(n1244), .A2(n1074), .ZN(n1216) );
AND3_X1 U902 ( .A1(n1080), .A2(n1082), .A3(n1240), .ZN(n1244) );
INV_X1 U903 ( .A(n1059), .ZN(n1082) );
NAND2_X1 U904 ( .A1(n1247), .A2(n1072), .ZN(n1059) );
INV_X1 U905 ( .A(n1071), .ZN(n1247) );
XNOR2_X1 U906 ( .A(G128), .B(n1217), .ZN(G30) );
NAND3_X1 U907 ( .A1(n1079), .A2(n1070), .A3(n1238), .ZN(n1217) );
AND3_X1 U908 ( .A1(n1248), .A2(n1249), .A3(n1240), .ZN(n1238) );
NOR3_X1 U909 ( .A1(n1250), .A2(n1085), .A3(n1060), .ZN(n1240) );
INV_X1 U910 ( .A(n1063), .ZN(n1060) );
OR2_X1 U911 ( .A1(n1251), .A2(n1074), .ZN(n1249) );
NAND2_X1 U912 ( .A1(n1252), .A2(n1251), .ZN(n1248) );
INV_X1 U913 ( .A(KEYINPUT20), .ZN(n1251) );
NAND2_X1 U914 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U915 ( .A(G101), .B(n1229), .Z(G3) );
AND4_X1 U916 ( .A1(n1053), .A2(n1074), .A3(n1070), .A4(n1228), .ZN(n1229) );
XNOR2_X1 U917 ( .A(G125), .B(n1255), .ZN(G27) );
NAND2_X1 U918 ( .A1(KEYINPUT59), .A2(n1256), .ZN(n1255) );
INV_X1 U919 ( .A(n1214), .ZN(n1256) );
NAND4_X1 U920 ( .A1(n1075), .A2(n1077), .A3(n1257), .A4(n1080), .ZN(n1214) );
NOR2_X1 U921 ( .A1(n1250), .A2(n1231), .ZN(n1257) );
AND2_X1 U922 ( .A1(n1048), .A2(n1258), .ZN(n1250) );
NAND3_X1 U923 ( .A1(G902), .A2(n1259), .A3(n1136), .ZN(n1258) );
NOR2_X1 U924 ( .A1(G900), .A2(n1131), .ZN(n1136) );
XOR2_X1 U925 ( .A(n1222), .B(n1260), .Z(G24) );
XNOR2_X1 U926 ( .A(G122), .B(KEYINPUT9), .ZN(n1260) );
NAND4_X1 U927 ( .A1(n1261), .A2(n1078), .A3(n1262), .A4(n1263), .ZN(n1222) );
NOR2_X1 U928 ( .A1(n1253), .A2(n1254), .ZN(n1078) );
XNOR2_X1 U929 ( .A(G119), .B(n1223), .ZN(G21) );
NAND4_X1 U930 ( .A1(n1264), .A2(n1053), .A3(n1254), .A4(n1261), .ZN(n1223) );
XNOR2_X1 U931 ( .A(KEYINPUT20), .B(n1265), .ZN(n1264) );
XNOR2_X1 U932 ( .A(G116), .B(n1266), .ZN(G18) );
NOR2_X1 U933 ( .A1(n1267), .A2(KEYINPUT0), .ZN(n1266) );
INV_X1 U934 ( .A(n1227), .ZN(n1267) );
NAND3_X1 U935 ( .A1(n1261), .A2(n1079), .A3(n1074), .ZN(n1227) );
NOR2_X1 U936 ( .A1(n1263), .A2(n1243), .ZN(n1079) );
INV_X1 U937 ( .A(n1262), .ZN(n1243) );
XNOR2_X1 U938 ( .A(G113), .B(n1226), .ZN(G15) );
NAND3_X1 U939 ( .A1(n1261), .A2(n1080), .A3(n1074), .ZN(n1226) );
NOR2_X1 U940 ( .A1(n1268), .A2(n1253), .ZN(n1074) );
INV_X1 U941 ( .A(n1265), .ZN(n1253) );
NOR2_X1 U942 ( .A1(n1262), .A2(n1242), .ZN(n1080) );
INV_X1 U943 ( .A(n1263), .ZN(n1242) );
AND3_X1 U944 ( .A1(n1070), .A2(n1269), .A3(n1077), .ZN(n1261) );
NOR2_X1 U945 ( .A1(n1063), .A2(n1085), .ZN(n1077) );
INV_X1 U946 ( .A(n1061), .ZN(n1085) );
XNOR2_X1 U947 ( .A(G110), .B(n1270), .ZN(G12) );
NAND2_X1 U948 ( .A1(n1271), .A2(n1070), .ZN(n1270) );
INV_X1 U949 ( .A(n1231), .ZN(n1070) );
NAND2_X1 U950 ( .A1(n1071), .A2(n1072), .ZN(n1231) );
NAND2_X1 U951 ( .A1(G214), .A2(n1272), .ZN(n1072) );
XOR2_X1 U952 ( .A(n1273), .B(n1211), .Z(n1071) );
NAND2_X1 U953 ( .A1(G210), .A2(n1272), .ZN(n1211) );
NAND2_X1 U954 ( .A1(n1274), .A2(n1275), .ZN(n1272) );
NAND3_X1 U955 ( .A1(n1276), .A2(n1275), .A3(n1277), .ZN(n1273) );
NAND3_X1 U956 ( .A1(n1278), .A2(n1185), .A3(KEYINPUT57), .ZN(n1277) );
XOR2_X1 U957 ( .A(n1279), .B(n1233), .Z(n1278) );
NOR2_X1 U958 ( .A1(KEYINPUT11), .A2(n1208), .ZN(n1279) );
INV_X1 U959 ( .A(n1280), .ZN(n1208) );
NAND2_X1 U960 ( .A1(n1281), .A2(n1282), .ZN(n1276) );
NAND2_X1 U961 ( .A1(KEYINPUT57), .A2(n1185), .ZN(n1282) );
XOR2_X1 U962 ( .A(n1283), .B(n1233), .Z(n1281) );
XNOR2_X1 U963 ( .A(n1153), .B(n1284), .ZN(n1233) );
XNOR2_X1 U964 ( .A(KEYINPUT58), .B(n1151), .ZN(n1284) );
XNOR2_X1 U965 ( .A(G122), .B(G110), .ZN(n1151) );
XOR2_X1 U966 ( .A(n1285), .B(n1286), .Z(n1153) );
XOR2_X1 U967 ( .A(KEYINPUT18), .B(n1287), .Z(n1286) );
NOR2_X1 U968 ( .A1(KEYINPUT26), .A2(n1288), .ZN(n1287) );
XOR2_X1 U969 ( .A(n1289), .B(n1290), .Z(n1285) );
NOR2_X1 U970 ( .A1(KEYINPUT11), .A2(n1280), .ZN(n1283) );
XOR2_X1 U971 ( .A(n1291), .B(n1130), .Z(n1280) );
INV_X1 U972 ( .A(G125), .ZN(n1130) );
NAND2_X1 U973 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U974 ( .A(KEYINPUT24), .B(n1145), .ZN(n1292) );
INV_X1 U975 ( .A(G224), .ZN(n1145) );
XOR2_X1 U976 ( .A(n1232), .B(KEYINPUT50), .Z(n1271) );
NAND3_X1 U977 ( .A1(n1053), .A2(n1228), .A3(n1075), .ZN(n1232) );
NOR2_X1 U978 ( .A1(n1265), .A2(n1254), .ZN(n1075) );
INV_X1 U979 ( .A(n1268), .ZN(n1254) );
XOR2_X1 U980 ( .A(n1294), .B(n1105), .Z(n1268) );
NAND2_X1 U981 ( .A1(n1295), .A2(n1275), .ZN(n1105) );
XOR2_X1 U982 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U983 ( .A(KEYINPUT3), .B(n1298), .ZN(n1297) );
INV_X1 U984 ( .A(n1185), .ZN(n1298) );
XNOR2_X1 U985 ( .A(n1299), .B(n1300), .ZN(n1185) );
NOR2_X1 U986 ( .A1(G128), .A2(KEYINPUT2), .ZN(n1300) );
XOR2_X1 U987 ( .A(n1301), .B(G143), .Z(n1299) );
NAND2_X1 U988 ( .A1(KEYINPUT54), .A2(n1302), .ZN(n1301) );
XNOR2_X1 U989 ( .A(n1183), .B(n1303), .ZN(n1296) );
INV_X1 U990 ( .A(n1176), .ZN(n1303) );
XOR2_X1 U991 ( .A(G101), .B(n1304), .Z(n1176) );
AND2_X1 U992 ( .A1(n1305), .A2(G210), .ZN(n1304) );
XOR2_X1 U993 ( .A(n1289), .B(n1306), .Z(n1183) );
XNOR2_X1 U994 ( .A(n1288), .B(n1204), .ZN(n1306) );
INV_X1 U995 ( .A(G119), .ZN(n1288) );
XNOR2_X1 U996 ( .A(G113), .B(G116), .ZN(n1289) );
NAND2_X1 U997 ( .A1(KEYINPUT13), .A2(n1106), .ZN(n1294) );
INV_X1 U998 ( .A(G472), .ZN(n1106) );
NAND2_X1 U999 ( .A1(n1307), .A2(n1308), .ZN(n1265) );
NAND2_X1 U1000 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XNOR2_X1 U1001 ( .A(n1108), .B(KEYINPUT55), .ZN(n1309) );
NAND2_X1 U1002 ( .A1(n1311), .A2(n1109), .ZN(n1307) );
INV_X1 U1003 ( .A(n1310), .ZN(n1109) );
NAND2_X1 U1004 ( .A1(n1312), .A2(G217), .ZN(n1310) );
XOR2_X1 U1005 ( .A(n1313), .B(KEYINPUT30), .Z(n1312) );
XNOR2_X1 U1006 ( .A(KEYINPUT15), .B(n1314), .ZN(n1311) );
INV_X1 U1007 ( .A(n1108), .ZN(n1314) );
NOR2_X1 U1008 ( .A1(n1163), .A2(G902), .ZN(n1108) );
INV_X1 U1009 ( .A(n1159), .ZN(n1163) );
XNOR2_X1 U1010 ( .A(n1315), .B(n1316), .ZN(n1159) );
XNOR2_X1 U1011 ( .A(n1317), .B(n1318), .ZN(n1316) );
XNOR2_X1 U1012 ( .A(n1302), .B(n1319), .ZN(n1318) );
NOR2_X1 U1013 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
INV_X1 U1014 ( .A(G221), .ZN(n1321) );
XOR2_X1 U1015 ( .A(n1322), .B(n1323), .Z(n1315) );
NOR2_X1 U1016 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
XOR2_X1 U1017 ( .A(n1326), .B(KEYINPUT23), .Z(n1325) );
NAND2_X1 U1018 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
XNOR2_X1 U1019 ( .A(n1329), .B(n1200), .ZN(n1327) );
XNOR2_X1 U1020 ( .A(KEYINPUT40), .B(KEYINPUT25), .ZN(n1329) );
NOR2_X1 U1021 ( .A1(G110), .A2(n1328), .ZN(n1324) );
XNOR2_X1 U1022 ( .A(G119), .B(n1330), .ZN(n1328) );
XOR2_X1 U1023 ( .A(KEYINPUT32), .B(G128), .Z(n1330) );
XNOR2_X1 U1024 ( .A(G137), .B(KEYINPUT60), .ZN(n1322) );
AND3_X1 U1025 ( .A1(n1269), .A2(n1061), .A3(n1063), .ZN(n1228) );
XOR2_X1 U1026 ( .A(n1090), .B(n1091), .Z(n1063) );
INV_X1 U1027 ( .A(G469), .ZN(n1091) );
NAND2_X1 U1028 ( .A1(n1331), .A2(n1275), .ZN(n1090) );
XOR2_X1 U1029 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1030 ( .A(KEYINPUT46), .B(n1334), .Z(n1333) );
NOR3_X1 U1031 ( .A1(n1335), .A2(n1336), .A3(n1196), .ZN(n1334) );
NOR3_X1 U1032 ( .A1(G110), .A2(G140), .A3(n1203), .ZN(n1196) );
INV_X1 U1033 ( .A(n1199), .ZN(n1336) );
NAND2_X1 U1034 ( .A1(n1337), .A2(G140), .ZN(n1199) );
XNOR2_X1 U1035 ( .A(n1201), .B(G110), .ZN(n1337) );
NOR3_X1 U1036 ( .A1(n1200), .A2(G140), .A3(n1201), .ZN(n1335) );
INV_X1 U1037 ( .A(n1203), .ZN(n1201) );
NAND2_X1 U1038 ( .A1(G227), .A2(n1293), .ZN(n1203) );
INV_X1 U1039 ( .A(G110), .ZN(n1200) );
XNOR2_X1 U1040 ( .A(n1190), .B(n1204), .ZN(n1332) );
XNOR2_X1 U1041 ( .A(n1338), .B(G131), .ZN(n1204) );
NAND2_X1 U1042 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NAND2_X1 U1043 ( .A1(G137), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1044 ( .A(n1342), .B(KEYINPUT36), .Z(n1339) );
OR2_X1 U1045 ( .A1(n1341), .A2(G137), .ZN(n1342) );
XNOR2_X1 U1046 ( .A(n1123), .B(n1290), .ZN(n1190) );
XNOR2_X1 U1047 ( .A(n1343), .B(n1344), .ZN(n1290) );
XNOR2_X1 U1048 ( .A(G101), .B(G104), .ZN(n1343) );
XOR2_X1 U1049 ( .A(n1345), .B(G128), .Z(n1123) );
NAND2_X1 U1050 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
NAND2_X1 U1051 ( .A1(G143), .A2(n1302), .ZN(n1347) );
XOR2_X1 U1052 ( .A(KEYINPUT17), .B(n1348), .Z(n1346) );
NOR2_X1 U1053 ( .A1(G143), .A2(n1302), .ZN(n1348) );
NAND2_X1 U1054 ( .A1(G221), .A2(n1313), .ZN(n1061) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1275), .ZN(n1313) );
NAND2_X1 U1056 ( .A1(n1048), .A2(n1349), .ZN(n1269) );
NAND4_X1 U1057 ( .A1(G902), .A2(G953), .A3(n1259), .A4(n1154), .ZN(n1349) );
INV_X1 U1058 ( .A(G898), .ZN(n1154) );
NAND3_X1 U1059 ( .A1(n1259), .A2(n1131), .A3(G952), .ZN(n1048) );
NAND2_X1 U1060 ( .A1(G237), .A2(G234), .ZN(n1259) );
NOR2_X1 U1061 ( .A1(n1262), .A2(n1263), .ZN(n1053) );
XNOR2_X1 U1062 ( .A(n1081), .B(KEYINPUT37), .ZN(n1263) );
XOR2_X1 U1063 ( .A(n1350), .B(G475), .Z(n1081) );
NAND2_X1 U1064 ( .A1(n1171), .A2(n1275), .ZN(n1350) );
XNOR2_X1 U1065 ( .A(n1351), .B(n1352), .ZN(n1171) );
XOR2_X1 U1066 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1067 ( .A(n1355), .B(n1356), .ZN(n1354) );
NOR2_X1 U1068 ( .A1(G104), .A2(KEYINPUT8), .ZN(n1356) );
NOR2_X1 U1069 ( .A1(KEYINPUT47), .A2(n1357), .ZN(n1355) );
XNOR2_X1 U1070 ( .A(n1358), .B(n1359), .ZN(n1357) );
INV_X1 U1071 ( .A(n1302), .ZN(n1359) );
XOR2_X1 U1072 ( .A(G146), .B(KEYINPUT4), .Z(n1302) );
NAND2_X1 U1073 ( .A1(KEYINPUT33), .A2(n1317), .ZN(n1358) );
XNOR2_X1 U1074 ( .A(G125), .B(n1129), .ZN(n1317) );
INV_X1 U1075 ( .A(G140), .ZN(n1129) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1305), .ZN(n1353) );
AND2_X1 U1077 ( .A1(n1293), .A2(n1274), .ZN(n1305) );
INV_X1 U1078 ( .A(G237), .ZN(n1274) );
XOR2_X1 U1079 ( .A(n1360), .B(n1361), .Z(n1351) );
XNOR2_X1 U1080 ( .A(G143), .B(n1246), .ZN(n1361) );
INV_X1 U1081 ( .A(G131), .ZN(n1246) );
XNOR2_X1 U1082 ( .A(G113), .B(G122), .ZN(n1360) );
XOR2_X1 U1083 ( .A(n1101), .B(n1098), .Z(n1262) );
INV_X1 U1084 ( .A(G478), .ZN(n1098) );
NAND2_X1 U1085 ( .A1(n1168), .A2(n1275), .ZN(n1101) );
INV_X1 U1086 ( .A(G902), .ZN(n1275) );
XNOR2_X1 U1087 ( .A(n1362), .B(n1363), .ZN(n1168) );
NOR2_X1 U1088 ( .A1(KEYINPUT31), .A2(n1364), .ZN(n1363) );
XOR2_X1 U1089 ( .A(n1365), .B(n1366), .Z(n1364) );
XNOR2_X1 U1090 ( .A(n1367), .B(n1344), .ZN(n1366) );
XOR2_X1 U1091 ( .A(G107), .B(KEYINPUT56), .Z(n1344) );
NAND2_X1 U1092 ( .A1(n1368), .A2(KEYINPUT53), .ZN(n1367) );
XNOR2_X1 U1093 ( .A(G128), .B(n1369), .ZN(n1368) );
XNOR2_X1 U1094 ( .A(G143), .B(n1341), .ZN(n1369) );
INV_X1 U1095 ( .A(G134), .ZN(n1341) );
XNOR2_X1 U1096 ( .A(G116), .B(G122), .ZN(n1365) );
OR2_X1 U1097 ( .A1(n1160), .A2(n1320), .ZN(n1362) );
NAND2_X1 U1098 ( .A1(G234), .A2(n1293), .ZN(n1320) );
XNOR2_X1 U1099 ( .A(n1131), .B(KEYINPUT14), .ZN(n1293) );
INV_X1 U1100 ( .A(G953), .ZN(n1131) );
INV_X1 U1101 ( .A(G217), .ZN(n1160) );
endmodule


