//Key = 1111100001000110110001101011110110011010001001100000101111101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321;

XNOR2_X1 U730 ( .A(G107), .B(n1000), .ZN(G9) );
NOR2_X1 U731 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR4_X1 U732 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1002) );
XOR2_X1 U733 ( .A(n1007), .B(KEYINPUT7), .Z(n1006) );
NAND3_X1 U734 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NAND4_X1 U735 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
NOR2_X1 U736 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND3_X1 U737 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1009) );
NAND2_X1 U738 ( .A1(n1012), .A2(n1020), .ZN(n1008) );
NAND3_X1 U739 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1020) );
NAND3_X1 U740 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
INV_X1 U741 ( .A(n1027), .ZN(n1026) );
NAND4_X1 U742 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1022) );
INV_X1 U743 ( .A(KEYINPUT6), .ZN(n1031) );
NOR3_X1 U744 ( .A1(n1015), .A2(n1032), .A3(n1033), .ZN(n1030) );
NAND2_X1 U745 ( .A1(KEYINPUT6), .A2(n1019), .ZN(n1021) );
INV_X1 U746 ( .A(n1034), .ZN(n1019) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1034), .ZN(n1005) );
NAND2_X1 U748 ( .A1(n1025), .A2(n1036), .ZN(n1034) );
NAND3_X1 U749 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1003) );
NAND2_X1 U750 ( .A1(n1012), .A2(n1040), .ZN(n1039) );
NAND2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U752 ( .A1(n1036), .A2(n1043), .A3(n1029), .ZN(n1042) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1013), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NAND2_X1 U756 ( .A1(n1025), .A2(n1049), .ZN(n1041) );
AND3_X1 U757 ( .A1(n1047), .A2(n1013), .A3(n1029), .ZN(n1025) );
INV_X1 U758 ( .A(n1016), .ZN(n1029) );
AND3_X1 U759 ( .A1(n1037), .A2(n1038), .A3(n1050), .ZN(n1001) );
NAND4_X1 U760 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1037) );
NOR2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U762 ( .A(KEYINPUT34), .B(n1018), .Z(n1056) );
XOR2_X1 U763 ( .A(G475), .B(n1057), .Z(n1055) );
XOR2_X1 U764 ( .A(n1058), .B(KEYINPUT56), .Z(n1053) );
NAND4_X1 U765 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1027), .ZN(n1058) );
XOR2_X1 U766 ( .A(n1062), .B(n1063), .Z(n1060) );
XNOR2_X1 U767 ( .A(n1064), .B(KEYINPUT13), .ZN(n1063) );
XNOR2_X1 U768 ( .A(n1065), .B(G469), .ZN(n1059) );
XOR2_X1 U769 ( .A(KEYINPUT16), .B(n1066), .Z(n1052) );
XOR2_X1 U770 ( .A(n1067), .B(n1068), .Z(G72) );
XOR2_X1 U771 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR3_X1 U772 ( .A1(n1071), .A2(KEYINPUT40), .A3(n1072), .ZN(n1070) );
XOR2_X1 U773 ( .A(n1073), .B(n1074), .Z(n1071) );
XNOR2_X1 U774 ( .A(n1075), .B(n1076), .ZN(n1074) );
NOR2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U776 ( .A(KEYINPUT33), .B(n1079), .Z(n1078) );
NOR2_X1 U777 ( .A1(G125), .A2(n1080), .ZN(n1079) );
NOR2_X1 U778 ( .A1(G140), .A2(n1081), .ZN(n1077) );
XOR2_X1 U779 ( .A(n1082), .B(n1083), .Z(n1073) );
XOR2_X1 U780 ( .A(KEYINPUT4), .B(G128), .Z(n1083) );
NOR2_X1 U781 ( .A1(n1084), .A2(n1085), .ZN(n1069) );
XOR2_X1 U782 ( .A(KEYINPUT44), .B(G953), .Z(n1085) );
NOR2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1088), .A2(n1038), .ZN(n1067) );
AND2_X1 U785 ( .A1(G227), .A2(G900), .ZN(n1088) );
NAND2_X1 U786 ( .A1(n1089), .A2(n1090), .ZN(G69) );
NAND2_X1 U787 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U788 ( .A1(G953), .A2(n1093), .ZN(n1092) );
NAND3_X1 U789 ( .A1(G953), .A2(n1094), .A3(n1095), .ZN(n1089) );
INV_X1 U790 ( .A(n1091), .ZN(n1095) );
NOR2_X1 U791 ( .A1(KEYINPUT50), .A2(n1096), .ZN(n1091) );
XOR2_X1 U792 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U793 ( .A1(n1099), .A2(G953), .ZN(n1098) );
NAND3_X1 U794 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1097) );
XOR2_X1 U795 ( .A(KEYINPUT45), .B(n1103), .Z(n1102) );
NOR2_X1 U796 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U797 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
XNOR2_X1 U798 ( .A(n1106), .B(n1107), .ZN(n1105) );
XNOR2_X1 U799 ( .A(n1108), .B(KEYINPUT47), .ZN(n1107) );
NAND2_X1 U800 ( .A1(n1109), .A2(KEYINPUT1), .ZN(n1108) );
XOR2_X1 U801 ( .A(n1110), .B(KEYINPUT54), .Z(n1109) );
NAND2_X1 U802 ( .A1(G953), .A2(n1111), .ZN(n1100) );
NAND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1094) );
NOR2_X1 U804 ( .A1(n1112), .A2(n1113), .ZN(G66) );
XOR2_X1 U805 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U806 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U807 ( .A1(KEYINPUT2), .A2(n1118), .ZN(n1114) );
NOR2_X1 U808 ( .A1(n1112), .A2(n1119), .ZN(G63) );
XNOR2_X1 U809 ( .A(n1120), .B(n1121), .ZN(n1119) );
AND2_X1 U810 ( .A1(G478), .A2(n1122), .ZN(n1121) );
NOR2_X1 U811 ( .A1(n1112), .A2(n1123), .ZN(G60) );
NOR3_X1 U812 ( .A1(n1057), .A2(n1124), .A3(n1125), .ZN(n1123) );
AND3_X1 U813 ( .A1(n1126), .A2(G475), .A3(n1122), .ZN(n1125) );
NOR2_X1 U814 ( .A1(n1127), .A2(n1126), .ZN(n1124) );
AND2_X1 U815 ( .A1(n1004), .A2(G475), .ZN(n1127) );
XOR2_X1 U816 ( .A(n1128), .B(n1129), .Z(G6) );
NOR3_X1 U817 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(G57) );
AND2_X1 U818 ( .A1(KEYINPUT29), .A2(n1112), .ZN(n1132) );
NOR3_X1 U819 ( .A1(KEYINPUT29), .A2(n1038), .A3(n1050), .ZN(n1131) );
INV_X1 U820 ( .A(G952), .ZN(n1050) );
XOR2_X1 U821 ( .A(n1133), .B(n1134), .Z(n1130) );
NOR2_X1 U822 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
XNOR2_X1 U823 ( .A(KEYINPUT8), .B(KEYINPUT60), .ZN(n1136) );
XOR2_X1 U824 ( .A(n1137), .B(n1138), .Z(n1135) );
XNOR2_X1 U825 ( .A(KEYINPUT17), .B(n1139), .ZN(n1138) );
NOR2_X1 U826 ( .A1(n1140), .A2(KEYINPUT43), .ZN(n1139) );
AND2_X1 U827 ( .A1(G472), .A2(n1122), .ZN(n1140) );
NOR2_X1 U828 ( .A1(n1141), .A2(n1142), .ZN(G54) );
XOR2_X1 U829 ( .A(KEYINPUT59), .B(n1112), .Z(n1142) );
XOR2_X1 U830 ( .A(n1143), .B(n1144), .Z(n1141) );
XOR2_X1 U831 ( .A(n1145), .B(n1146), .Z(n1144) );
AND2_X1 U832 ( .A1(G469), .A2(n1122), .ZN(n1146) );
INV_X1 U833 ( .A(n1117), .ZN(n1122) );
NAND3_X1 U834 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1145) );
INV_X1 U835 ( .A(n1150), .ZN(n1149) );
OR2_X1 U836 ( .A1(n1151), .A2(KEYINPUT0), .ZN(n1148) );
NAND3_X1 U837 ( .A1(n1151), .A2(n1152), .A3(KEYINPUT0), .ZN(n1147) );
NOR2_X1 U838 ( .A1(n1112), .A2(n1153), .ZN(G51) );
XNOR2_X1 U839 ( .A(n1154), .B(n1155), .ZN(n1153) );
XOR2_X1 U840 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U841 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
INV_X1 U842 ( .A(n1160), .ZN(n1159) );
NOR2_X1 U843 ( .A1(n1161), .A2(n1162), .ZN(n1158) );
NOR2_X1 U844 ( .A1(n1163), .A2(n1117), .ZN(n1156) );
NAND2_X1 U845 ( .A1(G902), .A2(n1004), .ZN(n1117) );
NAND3_X1 U846 ( .A1(n1099), .A2(n1164), .A3(n1165), .ZN(n1004) );
XNOR2_X1 U847 ( .A(n1086), .B(KEYINPUT19), .ZN(n1165) );
INV_X1 U848 ( .A(n1087), .ZN(n1164) );
NAND4_X1 U849 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1087) );
NOR4_X1 U850 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
INV_X1 U851 ( .A(n1174), .ZN(n1173) );
NAND3_X1 U852 ( .A1(n1011), .A2(n1175), .A3(n1176), .ZN(n1168) );
XOR2_X1 U853 ( .A(KEYINPUT49), .B(n1036), .Z(n1175) );
AND4_X1 U854 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1099) );
AND4_X1 U855 ( .A1(n1181), .A2(n1000), .A3(n1182), .A4(n1183), .ZN(n1180) );
NAND3_X1 U856 ( .A1(n1011), .A2(n1012), .A3(n1184), .ZN(n1000) );
NOR3_X1 U857 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1179) );
NOR3_X1 U858 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
NOR4_X1 U859 ( .A1(n1191), .A2(n1192), .A3(n1032), .A4(n1193), .ZN(n1189) );
INV_X1 U860 ( .A(n1194), .ZN(n1191) );
INV_X1 U861 ( .A(KEYINPUT30), .ZN(n1188) );
NOR4_X1 U862 ( .A1(KEYINPUT30), .A2(n1032), .A3(n1195), .A4(n1193), .ZN(n1186) );
XOR2_X1 U863 ( .A(n1196), .B(KEYINPUT22), .Z(n1193) );
INV_X1 U864 ( .A(n1129), .ZN(n1185) );
NAND3_X1 U865 ( .A1(n1184), .A2(n1012), .A3(n1046), .ZN(n1129) );
XNOR2_X1 U866 ( .A(n1064), .B(KEYINPUT51), .ZN(n1163) );
NOR2_X1 U867 ( .A1(n1038), .A2(G952), .ZN(n1112) );
XOR2_X1 U868 ( .A(n1197), .B(n1166), .Z(G48) );
NAND3_X1 U869 ( .A1(n1046), .A2(n1049), .A3(n1198), .ZN(n1166) );
XOR2_X1 U870 ( .A(n1199), .B(n1167), .Z(G45) );
NAND4_X1 U871 ( .A1(n1200), .A2(n1176), .A3(n1049), .A4(n1201), .ZN(n1167) );
XOR2_X1 U872 ( .A(G140), .B(n1172), .Z(G42) );
AND3_X1 U873 ( .A1(n1202), .A2(n1048), .A3(n1036), .ZN(n1172) );
NAND2_X1 U874 ( .A1(n1203), .A2(n1204), .ZN(G39) );
NAND2_X1 U875 ( .A1(n1086), .A2(n1205), .ZN(n1204) );
XOR2_X1 U876 ( .A(KEYINPUT35), .B(n1206), .Z(n1203) );
NOR2_X1 U877 ( .A1(n1086), .A2(n1205), .ZN(n1206) );
AND3_X1 U878 ( .A1(n1198), .A2(n1047), .A3(n1036), .ZN(n1086) );
XOR2_X1 U879 ( .A(G134), .B(n1207), .Z(G36) );
NOR4_X1 U880 ( .A1(KEYINPUT48), .A2(n1208), .A3(n1015), .A4(n1209), .ZN(n1207) );
XOR2_X1 U881 ( .A(n1210), .B(n1174), .Z(G33) );
NAND3_X1 U882 ( .A1(n1036), .A2(n1046), .A3(n1176), .ZN(n1174) );
INV_X1 U883 ( .A(n1209), .ZN(n1176) );
NAND3_X1 U884 ( .A1(n1048), .A2(n1211), .A3(n1196), .ZN(n1209) );
INV_X1 U885 ( .A(n1015), .ZN(n1036) );
NAND2_X1 U886 ( .A1(n1024), .A2(n1027), .ZN(n1015) );
XOR2_X1 U887 ( .A(G128), .B(n1171), .Z(G30) );
AND3_X1 U888 ( .A1(n1011), .A2(n1049), .A3(n1198), .ZN(n1171) );
AND4_X1 U889 ( .A1(n1048), .A2(n1018), .A3(n1066), .A4(n1211), .ZN(n1198) );
XOR2_X1 U890 ( .A(n1212), .B(n1213), .Z(G3) );
XOR2_X1 U891 ( .A(KEYINPUT27), .B(G101), .Z(n1213) );
NAND4_X1 U892 ( .A1(KEYINPUT24), .A2(n1047), .A3(n1196), .A4(n1184), .ZN(n1212) );
XOR2_X1 U893 ( .A(G125), .B(n1170), .Z(G27) );
AND3_X1 U894 ( .A1(n1013), .A2(n1049), .A3(n1202), .ZN(n1170) );
AND4_X1 U895 ( .A1(n1017), .A2(n1046), .A3(n1018), .A4(n1211), .ZN(n1202) );
NAND2_X1 U896 ( .A1(n1016), .A2(n1214), .ZN(n1211) );
NAND3_X1 U897 ( .A1(G902), .A2(n1215), .A3(n1072), .ZN(n1214) );
NOR2_X1 U898 ( .A1(n1038), .A2(G900), .ZN(n1072) );
XNOR2_X1 U899 ( .A(G122), .B(n1177), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1200), .A2(n1216), .A3(n1012), .A4(n1201), .ZN(n1177) );
NOR2_X1 U901 ( .A1(n1066), .A2(n1018), .ZN(n1012) );
NAND2_X1 U902 ( .A1(n1217), .A2(n1218), .ZN(G21) );
OR2_X1 U903 ( .A1(n1219), .A2(G119), .ZN(n1218) );
NAND2_X1 U904 ( .A1(G119), .A2(n1220), .ZN(n1217) );
NAND2_X1 U905 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
OR2_X1 U906 ( .A1(n1178), .A2(KEYINPUT31), .ZN(n1222) );
NAND2_X1 U907 ( .A1(KEYINPUT31), .A2(n1219), .ZN(n1221) );
OR2_X1 U908 ( .A1(KEYINPUT20), .A2(n1178), .ZN(n1219) );
NAND4_X1 U909 ( .A1(n1047), .A2(n1216), .A3(n1018), .A4(n1066), .ZN(n1178) );
XNOR2_X1 U910 ( .A(G116), .B(n1223), .ZN(G18) );
NOR2_X1 U911 ( .A1(n1224), .A2(KEYINPUT25), .ZN(n1223) );
INV_X1 U912 ( .A(n1181), .ZN(n1224) );
NAND3_X1 U913 ( .A1(n1196), .A2(n1011), .A3(n1216), .ZN(n1181) );
INV_X1 U914 ( .A(n1208), .ZN(n1011) );
NAND2_X1 U915 ( .A1(n1225), .A2(n1201), .ZN(n1208) );
XNOR2_X1 U916 ( .A(G113), .B(n1183), .ZN(G15) );
NAND3_X1 U917 ( .A1(n1216), .A2(n1196), .A3(n1046), .ZN(n1183) );
NOR2_X1 U918 ( .A1(n1225), .A2(n1201), .ZN(n1046) );
INV_X1 U919 ( .A(n1051), .ZN(n1201) );
INV_X1 U920 ( .A(n1035), .ZN(n1196) );
NAND2_X1 U921 ( .A1(n1226), .A2(n1066), .ZN(n1035) );
INV_X1 U922 ( .A(n1017), .ZN(n1066) );
AND3_X1 U923 ( .A1(n1049), .A2(n1194), .A3(n1013), .ZN(n1216) );
NOR2_X1 U924 ( .A1(n1033), .A2(n1028), .ZN(n1013) );
INV_X1 U925 ( .A(n1061), .ZN(n1028) );
XNOR2_X1 U926 ( .A(G110), .B(n1182), .ZN(G12) );
NAND4_X1 U927 ( .A1(n1047), .A2(n1184), .A3(n1017), .A4(n1018), .ZN(n1182) );
INV_X1 U928 ( .A(n1226), .ZN(n1018) );
XNOR2_X1 U929 ( .A(n1227), .B(n1116), .ZN(n1226) );
NAND2_X1 U930 ( .A1(G217), .A2(n1228), .ZN(n1116) );
NAND2_X1 U931 ( .A1(n1118), .A2(n1229), .ZN(n1227) );
XOR2_X1 U932 ( .A(n1230), .B(n1231), .Z(n1118) );
XOR2_X1 U933 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U934 ( .A(G137), .B(G110), .Z(n1233) );
XOR2_X1 U935 ( .A(KEYINPUT46), .B(G146), .Z(n1232) );
XOR2_X1 U936 ( .A(n1234), .B(n1235), .Z(n1230) );
XOR2_X1 U937 ( .A(n1236), .B(n1237), .Z(n1235) );
AND3_X1 U938 ( .A1(G221), .A2(n1038), .A3(n1238), .ZN(n1237) );
NOR2_X1 U939 ( .A1(KEYINPUT10), .A2(n1239), .ZN(n1236) );
NOR2_X1 U940 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
XOR2_X1 U941 ( .A(n1242), .B(KEYINPUT14), .Z(n1241) );
NAND2_X1 U942 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U943 ( .A(KEYINPUT23), .B(G119), .Z(n1243) );
NOR2_X1 U944 ( .A1(G119), .A2(n1245), .ZN(n1240) );
XOR2_X1 U945 ( .A(n1244), .B(KEYINPUT37), .Z(n1245) );
INV_X1 U946 ( .A(G128), .ZN(n1244) );
NAND2_X1 U947 ( .A1(n1246), .A2(n1247), .ZN(n1234) );
NAND2_X1 U948 ( .A1(KEYINPUT38), .A2(n1248), .ZN(n1247) );
NAND3_X1 U949 ( .A1(n1249), .A2(n1081), .A3(n1250), .ZN(n1246) );
INV_X1 U950 ( .A(KEYINPUT38), .ZN(n1250) );
XOR2_X1 U951 ( .A(n1251), .B(G472), .Z(n1017) );
NAND2_X1 U952 ( .A1(n1252), .A2(n1229), .ZN(n1251) );
XNOR2_X1 U953 ( .A(n1134), .B(n1137), .ZN(n1252) );
XOR2_X1 U954 ( .A(n1253), .B(n1254), .Z(n1137) );
XOR2_X1 U955 ( .A(KEYINPUT58), .B(n1255), .Z(n1254) );
XOR2_X1 U956 ( .A(n1256), .B(n1257), .Z(n1253) );
XNOR2_X1 U957 ( .A(n1258), .B(G101), .ZN(n1134) );
NAND2_X1 U958 ( .A1(n1259), .A2(G210), .ZN(n1258) );
INV_X1 U959 ( .A(n1195), .ZN(n1184) );
NAND3_X1 U960 ( .A1(n1048), .A2(n1194), .A3(n1049), .ZN(n1195) );
INV_X1 U961 ( .A(n1190), .ZN(n1049) );
NAND2_X1 U962 ( .A1(n1260), .A2(n1027), .ZN(n1190) );
NAND2_X1 U963 ( .A1(G214), .A2(n1261), .ZN(n1027) );
INV_X1 U964 ( .A(n1024), .ZN(n1260) );
XNOR2_X1 U965 ( .A(n1262), .B(n1062), .ZN(n1024) );
NAND2_X1 U966 ( .A1(n1263), .A2(n1229), .ZN(n1062) );
XOR2_X1 U967 ( .A(n1264), .B(n1265), .Z(n1263) );
NAND2_X1 U968 ( .A1(KEYINPUT57), .A2(n1154), .ZN(n1265) );
XOR2_X1 U969 ( .A(n1266), .B(n1106), .Z(n1154) );
XNOR2_X1 U970 ( .A(G104), .B(n1267), .ZN(n1106) );
XOR2_X1 U971 ( .A(n1268), .B(n1255), .Z(n1266) );
INV_X1 U972 ( .A(n1110), .ZN(n1255) );
XNOR2_X1 U973 ( .A(G113), .B(n1269), .ZN(n1110) );
XOR2_X1 U974 ( .A(G119), .B(G116), .Z(n1269) );
NAND2_X1 U975 ( .A1(KEYINPUT26), .A2(n1104), .ZN(n1268) );
XNOR2_X1 U976 ( .A(G110), .B(G122), .ZN(n1104) );
NAND3_X1 U977 ( .A1(n1270), .A2(n1271), .A3(n1160), .ZN(n1264) );
NAND2_X1 U978 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
OR3_X1 U979 ( .A1(n1162), .A2(n1161), .A3(KEYINPUT12), .ZN(n1271) );
XOR2_X1 U980 ( .A(n1272), .B(n1257), .Z(n1162) );
XOR2_X1 U981 ( .A(n1081), .B(G128), .Z(n1272) );
INV_X1 U982 ( .A(G125), .ZN(n1081) );
NAND2_X1 U983 ( .A1(KEYINPUT12), .A2(n1161), .ZN(n1270) );
NOR2_X1 U984 ( .A1(n1093), .A2(G953), .ZN(n1161) );
INV_X1 U985 ( .A(G224), .ZN(n1093) );
NAND2_X1 U986 ( .A1(KEYINPUT36), .A2(n1064), .ZN(n1262) );
AND2_X1 U987 ( .A1(G210), .A2(n1261), .ZN(n1064) );
NAND2_X1 U988 ( .A1(n1273), .A2(n1229), .ZN(n1261) );
INV_X1 U989 ( .A(G237), .ZN(n1273) );
NAND2_X1 U990 ( .A1(n1016), .A2(n1274), .ZN(n1194) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1215), .A4(n1111), .ZN(n1274) );
INV_X1 U992 ( .A(G898), .ZN(n1111) );
NAND3_X1 U993 ( .A1(n1215), .A2(n1038), .A3(G952), .ZN(n1016) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1215) );
INV_X1 U995 ( .A(n1192), .ZN(n1048) );
NAND2_X1 U996 ( .A1(n1033), .A2(n1061), .ZN(n1192) );
NAND2_X1 U997 ( .A1(G221), .A2(n1228), .ZN(n1061) );
NAND2_X1 U998 ( .A1(G234), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U999 ( .A(n1275), .B(n1276), .ZN(n1033) );
NOR2_X1 U1000 ( .A1(KEYINPUT61), .A2(n1065), .ZN(n1276) );
AND2_X1 U1001 ( .A1(n1277), .A2(n1229), .ZN(n1065) );
XOR2_X1 U1002 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U1003 ( .A(KEYINPUT52), .B(n1280), .Z(n1279) );
NOR2_X1 U1004 ( .A1(n1150), .A2(n1281), .ZN(n1280) );
AND2_X1 U1005 ( .A1(n1152), .A2(n1151), .ZN(n1281) );
NOR2_X1 U1006 ( .A1(n1152), .A2(n1151), .ZN(n1150) );
XNOR2_X1 U1007 ( .A(G110), .B(n1080), .ZN(n1151) );
INV_X1 U1008 ( .A(G140), .ZN(n1080) );
NAND2_X1 U1009 ( .A1(G227), .A2(n1038), .ZN(n1152) );
INV_X1 U1010 ( .A(n1143), .ZN(n1278) );
XOR2_X1 U1011 ( .A(n1282), .B(n1283), .Z(n1143) );
XNOR2_X1 U1012 ( .A(n1256), .B(n1267), .ZN(n1283) );
XOR2_X1 U1013 ( .A(G101), .B(G107), .Z(n1267) );
XOR2_X1 U1014 ( .A(n1284), .B(G128), .Z(n1256) );
NAND2_X1 U1015 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND3_X1 U1016 ( .A1(G131), .A2(n1287), .A3(n1288), .ZN(n1286) );
INV_X1 U1017 ( .A(KEYINPUT32), .ZN(n1288) );
NAND2_X1 U1018 ( .A1(n1075), .A2(KEYINPUT32), .ZN(n1285) );
XNOR2_X1 U1019 ( .A(n1210), .B(n1287), .ZN(n1075) );
XNOR2_X1 U1020 ( .A(G134), .B(n1205), .ZN(n1287) );
INV_X1 U1021 ( .A(G137), .ZN(n1205) );
XNOR2_X1 U1022 ( .A(n1289), .B(n1082), .ZN(n1282) );
NAND3_X1 U1023 ( .A1(n1290), .A2(n1291), .A3(KEYINPUT42), .ZN(n1082) );
OR2_X1 U1024 ( .A1(n1257), .A2(KEYINPUT5), .ZN(n1291) );
XNOR2_X1 U1025 ( .A(n1197), .B(G143), .ZN(n1257) );
INV_X1 U1026 ( .A(G146), .ZN(n1197) );
NAND3_X1 U1027 ( .A1(G146), .A2(n1199), .A3(KEYINPUT5), .ZN(n1290) );
NAND2_X1 U1028 ( .A1(KEYINPUT21), .A2(n1128), .ZN(n1289) );
INV_X1 U1029 ( .A(G104), .ZN(n1128) );
XNOR2_X1 U1030 ( .A(G469), .B(KEYINPUT9), .ZN(n1275) );
INV_X1 U1031 ( .A(n1032), .ZN(n1047) );
NAND2_X1 U1032 ( .A1(n1051), .A2(n1225), .ZN(n1032) );
INV_X1 U1033 ( .A(n1200), .ZN(n1225) );
XOR2_X1 U1034 ( .A(n1292), .B(n1293), .Z(n1200) );
NOR2_X1 U1035 ( .A1(KEYINPUT39), .A2(G475), .ZN(n1293) );
XNOR2_X1 U1036 ( .A(n1057), .B(KEYINPUT41), .ZN(n1292) );
NOR2_X1 U1037 ( .A1(n1126), .A2(G902), .ZN(n1057) );
XOR2_X1 U1038 ( .A(n1294), .B(n1295), .Z(n1126) );
XOR2_X1 U1039 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1040 ( .A(G122), .B(G113), .Z(n1297) );
XOR2_X1 U1041 ( .A(KEYINPUT62), .B(G146), .Z(n1296) );
XNOR2_X1 U1042 ( .A(n1298), .B(n1248), .ZN(n1294) );
XNOR2_X1 U1043 ( .A(G125), .B(n1249), .ZN(n1248) );
XOR2_X1 U1044 ( .A(G140), .B(KEYINPUT11), .Z(n1249) );
XOR2_X1 U1045 ( .A(n1299), .B(G104), .Z(n1298) );
NAND3_X1 U1046 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1299) );
NAND2_X1 U1047 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
INV_X1 U1048 ( .A(KEYINPUT28), .ZN(n1304) );
NAND3_X1 U1049 ( .A1(KEYINPUT28), .A2(n1305), .A3(n1210), .ZN(n1301) );
OR2_X1 U1050 ( .A1(n1210), .A2(n1305), .ZN(n1300) );
NOR2_X1 U1051 ( .A1(n1306), .A2(n1303), .ZN(n1305) );
XNOR2_X1 U1052 ( .A(n1307), .B(G143), .ZN(n1303) );
NAND2_X1 U1053 ( .A1(n1259), .A2(G214), .ZN(n1307) );
NOR2_X1 U1054 ( .A1(G953), .A2(G237), .ZN(n1259) );
INV_X1 U1055 ( .A(KEYINPUT55), .ZN(n1306) );
INV_X1 U1056 ( .A(G131), .ZN(n1210) );
XOR2_X1 U1057 ( .A(n1308), .B(G478), .Z(n1051) );
NAND2_X1 U1058 ( .A1(n1120), .A2(n1229), .ZN(n1308) );
INV_X1 U1059 ( .A(G902), .ZN(n1229) );
XNOR2_X1 U1060 ( .A(n1309), .B(n1310), .ZN(n1120) );
NOR2_X1 U1061 ( .A1(KEYINPUT63), .A2(n1311), .ZN(n1310) );
XOR2_X1 U1062 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1063 ( .A(G122), .B(G116), .Z(n1313) );
NAND2_X1 U1064 ( .A1(n1314), .A2(n1315), .ZN(n1312) );
NAND2_X1 U1065 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
XOR2_X1 U1066 ( .A(n1199), .B(G128), .Z(n1316) );
INV_X1 U1067 ( .A(G143), .ZN(n1199) );
NAND2_X1 U1068 ( .A1(n1318), .A2(n1319), .ZN(n1314) );
XNOR2_X1 U1069 ( .A(n1317), .B(n1320), .ZN(n1319) );
XNOR2_X1 U1070 ( .A(KEYINPUT53), .B(KEYINPUT3), .ZN(n1320) );
XOR2_X1 U1071 ( .A(G134), .B(n1321), .Z(n1317) );
NOR2_X1 U1072 ( .A1(KEYINPUT15), .A2(G107), .ZN(n1321) );
XOR2_X1 U1073 ( .A(G143), .B(G128), .Z(n1318) );
NAND3_X1 U1074 ( .A1(n1238), .A2(n1038), .A3(G217), .ZN(n1309) );
INV_X1 U1075 ( .A(G953), .ZN(n1038) );
XOR2_X1 U1076 ( .A(G234), .B(KEYINPUT18), .Z(n1238) );
endmodule


