//Key = 0111111011101100100001011001010101111010010011110010100011010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372;

XNOR2_X1 U762 ( .A(n1049), .B(n1050), .ZN(G9) );
XOR2_X1 U763 ( .A(KEYINPUT6), .B(G107), .Z(n1050) );
NOR2_X1 U764 ( .A1(n1051), .A2(n1052), .ZN(G75) );
NOR4_X1 U765 ( .A1(n1053), .A2(n1054), .A3(G953), .A4(n1055), .ZN(n1052) );
NOR2_X1 U766 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U767 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR4_X1 U768 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
NOR3_X1 U769 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1061) );
NOR2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U772 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U773 ( .A1(n1073), .A2(n1074), .ZN(n1065) );
NOR2_X1 U774 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1060) );
NOR2_X1 U776 ( .A1(n1079), .A2(n1068), .ZN(n1077) );
XOR2_X1 U777 ( .A(n1074), .B(KEYINPUT26), .Z(n1079) );
NOR3_X1 U778 ( .A1(n1080), .A2(n1064), .A3(n1068), .ZN(n1058) );
NAND3_X1 U779 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
NAND2_X1 U780 ( .A1(n1063), .A2(n1062), .ZN(n1082) );
NAND3_X1 U781 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1081) );
NOR3_X1 U782 ( .A1(n1055), .A2(G953), .A3(G952), .ZN(n1051) );
AND4_X1 U783 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1055) );
NOR3_X1 U784 ( .A1(n1091), .A2(n1064), .A3(n1092), .ZN(n1090) );
NOR2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND3_X1 U786 ( .A1(n1095), .A2(n1072), .A3(n1096), .ZN(n1091) );
NOR3_X1 U787 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1089) );
XOR2_X1 U788 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U789 ( .A1(G472), .A2(KEYINPUT30), .ZN(n1101) );
XOR2_X1 U790 ( .A(n1102), .B(KEYINPUT1), .Z(n1098) );
XOR2_X1 U791 ( .A(n1103), .B(n1104), .Z(n1088) );
XOR2_X1 U792 ( .A(KEYINPUT27), .B(G469), .Z(n1104) );
NAND2_X1 U793 ( .A1(KEYINPUT23), .A2(n1105), .ZN(n1103) );
XNOR2_X1 U794 ( .A(n1106), .B(n1107), .ZN(n1087) );
XOR2_X1 U795 ( .A(n1108), .B(n1109), .Z(G72) );
XOR2_X1 U796 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U798 ( .A1(G953), .A2(n1114), .ZN(n1113) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1112) );
XOR2_X1 U800 ( .A(G125), .B(n1117), .Z(n1116) );
NOR2_X1 U801 ( .A1(KEYINPUT43), .A2(n1118), .ZN(n1117) );
XOR2_X1 U802 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U803 ( .A(G137), .B(n1121), .Z(n1120) );
XOR2_X1 U804 ( .A(n1122), .B(KEYINPUT24), .Z(n1115) );
NAND2_X1 U805 ( .A1(n1123), .A2(G953), .ZN(n1110) );
XOR2_X1 U806 ( .A(n1124), .B(KEYINPUT60), .Z(n1123) );
NAND2_X1 U807 ( .A1(n1125), .A2(G227), .ZN(n1124) );
XOR2_X1 U808 ( .A(n1114), .B(KEYINPUT21), .Z(n1125) );
NOR3_X1 U809 ( .A1(n1126), .A2(KEYINPUT39), .A3(G953), .ZN(n1108) );
XOR2_X1 U810 ( .A(n1127), .B(n1128), .Z(G69) );
NOR2_X1 U811 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U812 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
INV_X1 U813 ( .A(G224), .ZN(n1132) );
XNOR2_X1 U814 ( .A(G898), .B(KEYINPUT32), .ZN(n1131) );
NOR2_X1 U815 ( .A1(KEYINPUT42), .A2(n1133), .ZN(n1127) );
XOR2_X1 U816 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U817 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U818 ( .A1(n1138), .A2(n1139), .ZN(n1134) );
NAND2_X1 U819 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U820 ( .A(KEYINPUT9), .B(G953), .Z(n1138) );
NOR2_X1 U821 ( .A1(n1142), .A2(n1143), .ZN(G66) );
XNOR2_X1 U822 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U824 ( .A1(n1142), .A2(n1148), .ZN(G63) );
XOR2_X1 U825 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U826 ( .A1(n1151), .A2(n1147), .ZN(n1150) );
NOR2_X1 U827 ( .A1(KEYINPUT19), .A2(n1152), .ZN(n1149) );
NOR2_X1 U828 ( .A1(n1142), .A2(n1153), .ZN(G60) );
XOR2_X1 U829 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U830 ( .A1(n1094), .A2(n1147), .ZN(n1154) );
NAND2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(G6) );
OR2_X1 U832 ( .A1(n1158), .A2(G104), .ZN(n1157) );
XOR2_X1 U833 ( .A(n1159), .B(KEYINPUT7), .Z(n1156) );
NAND2_X1 U834 ( .A1(G104), .A2(n1158), .ZN(n1159) );
NOR2_X1 U835 ( .A1(n1142), .A2(n1160), .ZN(G57) );
NOR3_X1 U836 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
NOR2_X1 U837 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
INV_X1 U838 ( .A(n1166), .ZN(n1165) );
NOR2_X1 U839 ( .A1(KEYINPUT49), .A2(n1167), .ZN(n1164) );
XNOR2_X1 U840 ( .A(n1168), .B(KEYINPUT46), .ZN(n1167) );
NOR3_X1 U841 ( .A1(n1166), .A2(KEYINPUT49), .A3(n1168), .ZN(n1162) );
XOR2_X1 U842 ( .A(n1169), .B(n1170), .Z(n1166) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1147), .ZN(n1170) );
INV_X1 U844 ( .A(G472), .ZN(n1171) );
NAND2_X1 U845 ( .A1(n1172), .A2(n1173), .ZN(n1169) );
NAND2_X1 U846 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U847 ( .A(KEYINPUT16), .B(n1176), .Z(n1172) );
NOR2_X1 U848 ( .A1(n1177), .A2(n1175), .ZN(n1176) );
XNOR2_X1 U849 ( .A(n1178), .B(n1179), .ZN(n1175) );
NAND2_X1 U850 ( .A1(KEYINPUT38), .A2(n1180), .ZN(n1178) );
XOR2_X1 U851 ( .A(n1174), .B(KEYINPUT40), .Z(n1177) );
AND2_X1 U852 ( .A1(n1168), .A2(KEYINPUT49), .ZN(n1161) );
AND2_X1 U853 ( .A1(n1181), .A2(n1182), .ZN(n1168) );
NOR2_X1 U854 ( .A1(n1183), .A2(n1184), .ZN(G54) );
XOR2_X1 U855 ( .A(KEYINPUT14), .B(n1142), .Z(n1184) );
XOR2_X1 U856 ( .A(n1185), .B(n1186), .Z(n1183) );
XOR2_X1 U857 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U858 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U859 ( .A1(n1191), .A2(n1147), .ZN(n1190) );
INV_X1 U860 ( .A(G469), .ZN(n1191) );
NAND2_X1 U861 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
NAND2_X1 U862 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U863 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U864 ( .A1(KEYINPUT5), .A2(n1122), .ZN(n1197) );
XOR2_X1 U865 ( .A(n1198), .B(KEYINPUT25), .Z(n1194) );
NAND2_X1 U866 ( .A1(G140), .A2(n1199), .ZN(n1192) );
NAND2_X1 U867 ( .A1(KEYINPUT5), .A2(n1196), .ZN(n1199) );
XOR2_X1 U868 ( .A(G110), .B(KEYINPUT44), .Z(n1196) );
NAND2_X1 U869 ( .A1(KEYINPUT47), .A2(n1200), .ZN(n1187) );
XOR2_X1 U870 ( .A(n1201), .B(n1179), .Z(n1185) );
NAND4_X1 U871 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
NAND3_X1 U872 ( .A1(KEYINPUT50), .A2(n1206), .A3(n1180), .ZN(n1205) );
NAND2_X1 U873 ( .A1(KEYINPUT35), .A2(n1207), .ZN(n1206) );
NAND3_X1 U874 ( .A1(n1208), .A2(n1209), .A3(n1121), .ZN(n1204) );
INV_X1 U875 ( .A(KEYINPUT50), .ZN(n1209) );
NAND2_X1 U876 ( .A1(n1207), .A2(n1210), .ZN(n1208) );
INV_X1 U877 ( .A(KEYINPUT35), .ZN(n1210) );
OR2_X1 U878 ( .A1(n1207), .A2(KEYINPUT56), .ZN(n1203) );
NAND3_X1 U879 ( .A1(n1211), .A2(n1207), .A3(KEYINPUT56), .ZN(n1202) );
XOR2_X1 U880 ( .A(KEYINPUT35), .B(n1180), .Z(n1211) );
NOR2_X1 U881 ( .A1(n1142), .A2(n1212), .ZN(G51) );
XOR2_X1 U882 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U883 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR2_X1 U884 ( .A1(n1107), .A2(n1147), .ZN(n1216) );
NAND2_X1 U885 ( .A1(G902), .A2(n1053), .ZN(n1147) );
NAND3_X1 U886 ( .A1(n1217), .A2(n1126), .A3(n1140), .ZN(n1053) );
AND4_X1 U887 ( .A1(n1158), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1140) );
NOR3_X1 U888 ( .A1(n1221), .A2(n1049), .A3(n1222), .ZN(n1220) );
AND2_X1 U889 ( .A1(n1075), .A2(n1223), .ZN(n1049) );
INV_X1 U890 ( .A(n1224), .ZN(n1221) );
NAND2_X1 U891 ( .A1(n1225), .A2(n1226), .ZN(n1219) );
NAND2_X1 U892 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND3_X1 U893 ( .A1(n1229), .A2(n1230), .A3(n1076), .ZN(n1228) );
NAND2_X1 U894 ( .A1(KEYINPUT61), .A2(n1231), .ZN(n1230) );
NAND2_X1 U895 ( .A1(n1232), .A2(n1233), .ZN(n1229) );
INV_X1 U896 ( .A(KEYINPUT61), .ZN(n1233) );
NAND2_X1 U897 ( .A1(n1234), .A2(n1235), .ZN(n1232) );
INV_X1 U898 ( .A(n1236), .ZN(n1234) );
OR2_X1 U899 ( .A1(n1068), .A2(n1237), .ZN(n1227) );
NAND2_X1 U900 ( .A1(n1076), .A2(n1223), .ZN(n1158) );
NOR2_X1 U901 ( .A1(n1237), .A2(n1062), .ZN(n1223) );
INV_X1 U902 ( .A(n1238), .ZN(n1062) );
AND4_X1 U903 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1126) );
AND4_X1 U904 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242) );
NAND3_X1 U905 ( .A1(n1247), .A2(n1248), .A3(n1083), .ZN(n1239) );
NAND2_X1 U906 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NAND2_X1 U907 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U908 ( .A1(n1225), .A2(n1075), .ZN(n1249) );
XOR2_X1 U909 ( .A(n1141), .B(KEYINPUT54), .Z(n1217) );
NOR3_X1 U910 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1215) );
NOR3_X1 U911 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1255) );
AND2_X1 U912 ( .A1(n1256), .A2(n1258), .ZN(n1254) );
XOR2_X1 U913 ( .A(n1259), .B(KEYINPUT3), .Z(n1258) );
NAND2_X1 U914 ( .A1(n1121), .A2(n1260), .ZN(n1259) );
INV_X1 U915 ( .A(n1261), .ZN(n1253) );
NOR2_X1 U916 ( .A1(KEYINPUT20), .A2(n1262), .ZN(n1213) );
NOR2_X1 U917 ( .A1(n1130), .A2(G952), .ZN(n1142) );
XNOR2_X1 U918 ( .A(G146), .B(n1246), .ZN(G48) );
NAND3_X1 U919 ( .A1(n1263), .A2(n1070), .A3(n1251), .ZN(n1246) );
XNOR2_X1 U920 ( .A(G143), .B(n1245), .ZN(G45) );
NAND4_X1 U921 ( .A1(n1247), .A2(n1225), .A3(n1264), .A4(n1070), .ZN(n1245) );
NOR2_X1 U922 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XOR2_X1 U923 ( .A(n1244), .B(n1267), .Z(G42) );
XOR2_X1 U924 ( .A(KEYINPUT59), .B(G140), .Z(n1267) );
NAND3_X1 U925 ( .A1(n1263), .A2(n1268), .A3(n1083), .ZN(n1244) );
XNOR2_X1 U926 ( .A(G137), .B(n1269), .ZN(G39) );
NAND4_X1 U927 ( .A1(n1083), .A2(n1252), .A3(n1251), .A4(n1270), .ZN(n1269) );
NOR3_X1 U928 ( .A1(n1271), .A2(n1064), .A3(n1086), .ZN(n1270) );
INV_X1 U929 ( .A(n1078), .ZN(n1064) );
XOR2_X1 U930 ( .A(n1272), .B(KEYINPUT8), .Z(n1271) );
XNOR2_X1 U931 ( .A(G134), .B(n1273), .ZN(G36) );
NAND4_X1 U932 ( .A1(n1274), .A2(n1247), .A3(n1075), .A4(n1275), .ZN(n1273) );
XOR2_X1 U933 ( .A(KEYINPUT53), .B(n1083), .Z(n1275) );
XOR2_X1 U934 ( .A(n1084), .B(KEYINPUT57), .Z(n1274) );
NAND3_X1 U935 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(G33) );
NAND2_X1 U936 ( .A1(n1243), .A2(n1279), .ZN(n1278) );
OR3_X1 U937 ( .A1(n1279), .A2(n1243), .A3(n1280), .ZN(n1277) );
INV_X1 U938 ( .A(KEYINPUT13), .ZN(n1279) );
NAND2_X1 U939 ( .A1(n1280), .A2(n1281), .ZN(n1276) );
NAND2_X1 U940 ( .A1(n1282), .A2(KEYINPUT13), .ZN(n1281) );
XOR2_X1 U941 ( .A(n1243), .B(KEYINPUT31), .Z(n1282) );
NAND3_X1 U942 ( .A1(n1263), .A2(n1225), .A3(n1083), .ZN(n1243) );
INV_X1 U943 ( .A(n1074), .ZN(n1083) );
NAND2_X1 U944 ( .A1(n1283), .A2(n1072), .ZN(n1074) );
INV_X1 U945 ( .A(n1084), .ZN(n1225) );
AND2_X1 U946 ( .A1(n1247), .A2(n1076), .ZN(n1263) );
XOR2_X1 U947 ( .A(G131), .B(KEYINPUT55), .Z(n1280) );
XNOR2_X1 U948 ( .A(n1240), .B(n1284), .ZN(G30) );
NOR2_X1 U949 ( .A1(KEYINPUT11), .A2(n1285), .ZN(n1284) );
NAND4_X1 U950 ( .A1(n1251), .A2(n1247), .A3(n1075), .A4(n1070), .ZN(n1240) );
AND3_X1 U951 ( .A1(n1272), .A2(n1078), .A3(n1063), .ZN(n1247) );
XOR2_X1 U952 ( .A(G101), .B(n1286), .Z(G3) );
NOR3_X1 U953 ( .A1(n1084), .A2(n1287), .A3(n1237), .ZN(n1286) );
XOR2_X1 U954 ( .A(n1068), .B(KEYINPUT51), .Z(n1287) );
XOR2_X1 U955 ( .A(n1260), .B(n1288), .Z(G27) );
NAND2_X1 U956 ( .A1(KEYINPUT29), .A2(n1289), .ZN(n1288) );
INV_X1 U957 ( .A(n1241), .ZN(n1289) );
NAND4_X1 U958 ( .A1(n1076), .A2(n1235), .A3(n1268), .A4(n1272), .ZN(n1241) );
NAND2_X1 U959 ( .A1(n1057), .A2(n1290), .ZN(n1272) );
NAND4_X1 U960 ( .A1(G902), .A2(G953), .A3(n1291), .A4(n1114), .ZN(n1290) );
INV_X1 U961 ( .A(G900), .ZN(n1114) );
INV_X1 U962 ( .A(n1085), .ZN(n1268) );
XNOR2_X1 U963 ( .A(G122), .B(n1218), .ZN(G24) );
NAND4_X1 U964 ( .A1(n1292), .A2(n1238), .A3(n1293), .A4(n1294), .ZN(n1218) );
NOR2_X1 U965 ( .A1(n1097), .A2(n1295), .ZN(n1238) );
XOR2_X1 U966 ( .A(n1141), .B(n1296), .Z(G21) );
XOR2_X1 U967 ( .A(n1297), .B(KEYINPUT15), .Z(n1296) );
NAND3_X1 U968 ( .A1(n1292), .A2(n1252), .A3(n1251), .ZN(n1141) );
AND2_X1 U969 ( .A1(n1295), .A2(n1097), .ZN(n1251) );
INV_X1 U970 ( .A(n1068), .ZN(n1252) );
INV_X1 U971 ( .A(n1231), .ZN(n1292) );
XOR2_X1 U972 ( .A(n1298), .B(n1224), .Z(G18) );
NAND2_X1 U973 ( .A1(n1299), .A2(n1075), .ZN(n1224) );
NOR2_X1 U974 ( .A1(n1293), .A2(n1265), .ZN(n1075) );
XOR2_X1 U975 ( .A(G113), .B(n1300), .Z(G15) );
AND2_X1 U976 ( .A1(n1299), .A2(n1076), .ZN(n1300) );
NOR2_X1 U977 ( .A1(n1294), .A2(n1266), .ZN(n1076) );
NOR2_X1 U978 ( .A1(n1084), .A2(n1231), .ZN(n1299) );
NAND2_X1 U979 ( .A1(n1235), .A2(n1236), .ZN(n1231) );
AND3_X1 U980 ( .A1(n1070), .A2(n1078), .A3(n1086), .ZN(n1235) );
NAND2_X1 U981 ( .A1(n1301), .A2(n1295), .ZN(n1084) );
XOR2_X1 U982 ( .A(G110), .B(n1222), .Z(G12) );
NOR3_X1 U983 ( .A1(n1085), .A2(n1237), .A3(n1068), .ZN(n1222) );
NAND2_X1 U984 ( .A1(n1265), .A2(n1266), .ZN(n1068) );
INV_X1 U985 ( .A(n1293), .ZN(n1266) );
NAND3_X1 U986 ( .A1(n1302), .A2(n1303), .A3(n1095), .ZN(n1293) );
NAND2_X1 U987 ( .A1(n1093), .A2(n1094), .ZN(n1095) );
NAND2_X1 U988 ( .A1(n1093), .A2(n1304), .ZN(n1303) );
OR3_X1 U989 ( .A1(n1094), .A2(n1093), .A3(n1304), .ZN(n1302) );
INV_X1 U990 ( .A(KEYINPUT52), .ZN(n1304) );
NOR2_X1 U991 ( .A1(n1155), .A2(G902), .ZN(n1093) );
XNOR2_X1 U992 ( .A(n1305), .B(G146), .ZN(n1155) );
XOR2_X1 U993 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U994 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U995 ( .A(G131), .B(G122), .Z(n1309) );
XOR2_X1 U996 ( .A(G143), .B(G140), .Z(n1308) );
XOR2_X1 U997 ( .A(n1310), .B(n1311), .Z(n1306) );
XNOR2_X1 U998 ( .A(n1312), .B(n1313), .ZN(n1311) );
NOR2_X1 U999 ( .A1(G125), .A2(KEYINPUT0), .ZN(n1313) );
NAND3_X1 U1000 ( .A1(G214), .A2(n1314), .A3(KEYINPUT4), .ZN(n1312) );
XNOR2_X1 U1001 ( .A(G113), .B(G104), .ZN(n1310) );
INV_X1 U1002 ( .A(G475), .ZN(n1094) );
INV_X1 U1003 ( .A(n1294), .ZN(n1265) );
NAND2_X1 U1004 ( .A1(n1096), .A2(n1102), .ZN(n1294) );
NAND3_X1 U1005 ( .A1(n1315), .A2(n1316), .A3(n1152), .ZN(n1102) );
XOR2_X1 U1006 ( .A(KEYINPUT45), .B(G478), .Z(n1315) );
NAND2_X1 U1007 ( .A1(n1317), .A2(n1318), .ZN(n1096) );
NAND2_X1 U1008 ( .A1(n1152), .A2(n1316), .ZN(n1318) );
XOR2_X1 U1009 ( .A(n1319), .B(n1320), .Z(n1152) );
XNOR2_X1 U1010 ( .A(n1321), .B(n1322), .ZN(n1320) );
NOR2_X1 U1011 ( .A1(G107), .A2(KEYINPUT62), .ZN(n1321) );
XOR2_X1 U1012 ( .A(n1323), .B(n1324), .Z(n1319) );
XOR2_X1 U1013 ( .A(G134), .B(n1325), .Z(n1324) );
NOR2_X1 U1014 ( .A1(KEYINPUT22), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1015 ( .A(n1285), .B(G143), .Z(n1326) );
INV_X1 U1016 ( .A(G128), .ZN(n1285) );
NAND2_X1 U1017 ( .A1(G217), .A2(n1327), .ZN(n1323) );
XOR2_X1 U1018 ( .A(n1151), .B(KEYINPUT45), .Z(n1317) );
INV_X1 U1019 ( .A(G478), .ZN(n1151) );
NAND4_X1 U1020 ( .A1(n1070), .A2(n1063), .A3(n1078), .A4(n1236), .ZN(n1237) );
NAND2_X1 U1021 ( .A1(n1057), .A2(n1328), .ZN(n1236) );
NAND3_X1 U1022 ( .A1(n1136), .A2(n1291), .A3(G902), .ZN(n1328) );
NOR2_X1 U1023 ( .A1(n1130), .A2(G898), .ZN(n1136) );
NAND3_X1 U1024 ( .A1(n1291), .A2(n1130), .A3(G952), .ZN(n1057) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1291) );
NAND2_X1 U1026 ( .A1(G221), .A2(n1329), .ZN(n1078) );
INV_X1 U1027 ( .A(n1086), .ZN(n1063) );
XOR2_X1 U1028 ( .A(n1105), .B(n1330), .Z(n1086) );
XOR2_X1 U1029 ( .A(KEYINPUT37), .B(G469), .Z(n1330) );
NAND2_X1 U1030 ( .A1(n1331), .A2(n1316), .ZN(n1105) );
XOR2_X1 U1031 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1032 ( .A(n1207), .B(n1334), .Z(n1333) );
XOR2_X1 U1033 ( .A(n1121), .B(n1335), .Z(n1334) );
XOR2_X1 U1034 ( .A(n1336), .B(n1337), .Z(n1332) );
XNOR2_X1 U1035 ( .A(n1338), .B(KEYINPUT33), .ZN(n1337) );
NAND2_X1 U1036 ( .A1(KEYINPUT41), .A2(n1200), .ZN(n1338) );
AND2_X1 U1037 ( .A1(G227), .A2(n1130), .ZN(n1200) );
NAND2_X1 U1038 ( .A1(KEYINPUT34), .A2(n1179), .ZN(n1336) );
AND2_X1 U1039 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U1040 ( .A1(G214), .A2(n1339), .ZN(n1072) );
INV_X1 U1041 ( .A(n1283), .ZN(n1071) );
XOR2_X1 U1042 ( .A(n1340), .B(n1107), .Z(n1283) );
NAND2_X1 U1043 ( .A1(G210), .A2(n1339), .ZN(n1107) );
NAND2_X1 U1044 ( .A1(n1316), .A2(n1341), .ZN(n1339) );
INV_X1 U1045 ( .A(G237), .ZN(n1341) );
NAND2_X1 U1046 ( .A1(KEYINPUT12), .A2(n1106), .ZN(n1340) );
NAND2_X1 U1047 ( .A1(n1342), .A2(n1316), .ZN(n1106) );
XOR2_X1 U1048 ( .A(n1343), .B(n1262), .Z(n1342) );
INV_X1 U1049 ( .A(n1137), .ZN(n1262) );
XOR2_X1 U1050 ( .A(n1344), .B(n1345), .Z(n1137) );
XOR2_X1 U1051 ( .A(n1207), .B(n1322), .Z(n1345) );
XNOR2_X1 U1052 ( .A(G116), .B(G122), .ZN(n1322) );
XNOR2_X1 U1053 ( .A(n1346), .B(n1347), .ZN(n1207) );
XNOR2_X1 U1054 ( .A(G107), .B(G104), .ZN(n1346) );
XOR2_X1 U1055 ( .A(n1348), .B(n1349), .Z(n1344) );
XOR2_X1 U1056 ( .A(n1198), .B(KEYINPUT63), .Z(n1348) );
XOR2_X1 U1057 ( .A(n1350), .B(KEYINPUT36), .Z(n1343) );
NAND3_X1 U1058 ( .A1(n1351), .A2(n1352), .A3(n1261), .ZN(n1350) );
NAND2_X1 U1059 ( .A1(n1257), .A2(n1256), .ZN(n1261) );
NOR2_X1 U1060 ( .A1(n1260), .A2(n1121), .ZN(n1257) );
NAND2_X1 U1061 ( .A1(n1353), .A2(n1260), .ZN(n1352) );
INV_X1 U1062 ( .A(G125), .ZN(n1260) );
XOR2_X1 U1063 ( .A(n1256), .B(n1180), .Z(n1353) );
NAND3_X1 U1064 ( .A1(n1354), .A2(n1121), .A3(G125), .ZN(n1351) );
INV_X1 U1065 ( .A(n1180), .ZN(n1121) );
INV_X1 U1066 ( .A(n1256), .ZN(n1354) );
NAND2_X1 U1067 ( .A1(G224), .A2(n1130), .ZN(n1256) );
NAND2_X1 U1068 ( .A1(n1355), .A2(n1097), .ZN(n1085) );
INV_X1 U1069 ( .A(n1301), .ZN(n1097) );
XNOR2_X1 U1070 ( .A(n1356), .B(n1146), .ZN(n1301) );
NAND2_X1 U1071 ( .A1(G217), .A2(n1329), .ZN(n1146) );
NAND2_X1 U1072 ( .A1(G234), .A2(n1316), .ZN(n1329) );
NAND2_X1 U1073 ( .A1(n1144), .A2(n1316), .ZN(n1356) );
XNOR2_X1 U1074 ( .A(n1357), .B(n1358), .ZN(n1144) );
XOR2_X1 U1075 ( .A(G119), .B(n1359), .Z(n1358) );
XOR2_X1 U1076 ( .A(G137), .B(G125), .Z(n1359) );
XOR2_X1 U1077 ( .A(n1360), .B(n1335), .Z(n1357) );
XOR2_X1 U1078 ( .A(n1198), .B(n1122), .Z(n1335) );
INV_X1 U1079 ( .A(G140), .ZN(n1122) );
INV_X1 U1080 ( .A(G110), .ZN(n1198) );
XOR2_X1 U1081 ( .A(n1361), .B(n1362), .Z(n1360) );
NAND2_X1 U1082 ( .A1(G221), .A2(n1327), .ZN(n1361) );
AND2_X1 U1083 ( .A1(G234), .A2(n1130), .ZN(n1327) );
INV_X1 U1084 ( .A(G953), .ZN(n1130) );
XOR2_X1 U1085 ( .A(KEYINPUT10), .B(n1295), .Z(n1355) );
XNOR2_X1 U1086 ( .A(n1100), .B(G472), .ZN(n1295) );
NAND2_X1 U1087 ( .A1(n1363), .A2(n1316), .ZN(n1100) );
INV_X1 U1088 ( .A(G902), .ZN(n1316) );
XOR2_X1 U1089 ( .A(n1364), .B(n1365), .Z(n1363) );
XNOR2_X1 U1090 ( .A(n1179), .B(n1174), .ZN(n1365) );
XOR2_X1 U1091 ( .A(n1366), .B(n1349), .Z(n1174) );
XNOR2_X1 U1092 ( .A(G113), .B(n1297), .ZN(n1349) );
INV_X1 U1093 ( .A(G119), .ZN(n1297) );
NAND2_X1 U1094 ( .A1(KEYINPUT2), .A2(n1298), .ZN(n1366) );
INV_X1 U1095 ( .A(G116), .ZN(n1298) );
XOR2_X1 U1096 ( .A(n1119), .B(n1367), .Z(n1179) );
NOR2_X1 U1097 ( .A1(KEYINPUT18), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1098 ( .A(KEYINPUT48), .B(G137), .Z(n1368) );
XOR2_X1 U1099 ( .A(G131), .B(G134), .Z(n1119) );
XOR2_X1 U1100 ( .A(n1180), .B(n1369), .Z(n1364) );
XOR2_X1 U1101 ( .A(n1370), .B(KEYINPUT58), .Z(n1369) );
NAND2_X1 U1102 ( .A1(n1371), .A2(n1181), .ZN(n1370) );
NAND2_X1 U1103 ( .A1(n1347), .A2(n1372), .ZN(n1181) );
XOR2_X1 U1104 ( .A(n1182), .B(KEYINPUT28), .Z(n1371) );
OR2_X1 U1105 ( .A1(n1372), .A2(n1347), .ZN(n1182) );
XNOR2_X1 U1106 ( .A(G101), .B(KEYINPUT17), .ZN(n1347) );
NAND2_X1 U1107 ( .A1(G210), .A2(n1314), .ZN(n1372) );
NOR2_X1 U1108 ( .A1(G953), .A2(G237), .ZN(n1314) );
XNOR2_X1 U1109 ( .A(G143), .B(n1362), .ZN(n1180) );
XOR2_X1 U1110 ( .A(G128), .B(G146), .Z(n1362) );
endmodule


