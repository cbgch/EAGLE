//Key = 0010100100011010011010101111111000101011110111111011111101010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338;

XNOR2_X1 U740 ( .A(G107), .B(n1013), .ZN(G9) );
NAND2_X1 U741 ( .A1(KEYINPUT12), .A2(n1014), .ZN(n1013) );
INV_X1 U742 ( .A(n1015), .ZN(n1014) );
NOR2_X1 U743 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U744 ( .A1(n1018), .A2(n1019), .A3(G953), .A4(n1020), .ZN(n1017) );
NOR2_X1 U745 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
XNOR2_X1 U746 ( .A(KEYINPUT35), .B(n1023), .ZN(n1022) );
NOR2_X1 U747 ( .A1(n1024), .A2(n1025), .ZN(n1021) );
NOR2_X1 U748 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
INV_X1 U749 ( .A(n1028), .ZN(n1027) );
NOR2_X1 U750 ( .A1(n1029), .A2(n1030), .ZN(n1026) );
NOR2_X1 U751 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U752 ( .A1(n1033), .A2(n1034), .ZN(n1029) );
NOR2_X1 U753 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U754 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR2_X1 U755 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR3_X1 U756 ( .A1(n1031), .A2(n1042), .A3(n1043), .ZN(n1035) );
NOR3_X1 U757 ( .A1(n1038), .A2(n1044), .A3(n1045), .ZN(n1043) );
NOR2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U759 ( .A1(n1048), .A2(n1049), .ZN(n1042) );
NOR4_X1 U760 ( .A1(n1050), .A2(n1031), .A3(n1037), .A4(n1051), .ZN(n1024) );
INV_X1 U761 ( .A(n1052), .ZN(n1051) );
INV_X1 U762 ( .A(n1053), .ZN(n1031) );
NOR2_X1 U763 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
NAND2_X1 U764 ( .A1(KEYINPUT36), .A2(n1056), .ZN(n1018) );
NOR3_X1 U765 ( .A1(n1020), .A2(G953), .A3(G952), .ZN(n1016) );
AND4_X1 U766 ( .A1(n1052), .A2(n1048), .A3(n1057), .A4(n1058), .ZN(n1020) );
NOR3_X1 U767 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
XNOR2_X1 U768 ( .A(G475), .B(n1062), .ZN(n1060) );
NOR2_X1 U769 ( .A1(n1063), .A2(KEYINPUT9), .ZN(n1062) );
XOR2_X1 U770 ( .A(n1064), .B(n1065), .Z(n1057) );
XOR2_X1 U771 ( .A(KEYINPUT24), .B(n1066), .Z(n1065) );
NOR2_X1 U772 ( .A1(KEYINPUT3), .A2(G472), .ZN(n1066) );
XOR2_X1 U773 ( .A(n1067), .B(n1068), .Z(G72) );
XOR2_X1 U774 ( .A(n1069), .B(n1070), .Z(n1068) );
NAND2_X1 U775 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U776 ( .A1(G900), .A2(G227), .ZN(n1072) );
NAND2_X1 U777 ( .A1(n1073), .A2(n1074), .ZN(n1069) );
NAND2_X1 U778 ( .A1(G953), .A2(n1075), .ZN(n1074) );
XOR2_X1 U779 ( .A(n1076), .B(n1077), .Z(n1073) );
NAND2_X1 U780 ( .A1(KEYINPUT30), .A2(n1078), .ZN(n1076) );
NOR2_X1 U781 ( .A1(n1079), .A2(G953), .ZN(n1067) );
XOR2_X1 U782 ( .A(n1080), .B(n1081), .Z(G69) );
XOR2_X1 U783 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U784 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
INV_X1 U785 ( .A(n1071), .ZN(n1085) );
XOR2_X1 U786 ( .A(G953), .B(KEYINPUT37), .Z(n1071) );
AND2_X1 U787 ( .A1(G224), .A2(G898), .ZN(n1084) );
NAND2_X1 U788 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
INV_X1 U789 ( .A(n1088), .ZN(n1087) );
XOR2_X1 U790 ( .A(n1089), .B(n1090), .Z(n1086) );
NAND2_X1 U791 ( .A1(n1091), .A2(n1092), .ZN(n1080) );
NAND2_X1 U792 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XNOR2_X1 U793 ( .A(KEYINPUT48), .B(n1095), .ZN(n1094) );
NOR2_X1 U794 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XOR2_X1 U795 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND3_X1 U796 ( .A1(n1100), .A2(G217), .A3(KEYINPUT38), .ZN(n1098) );
NOR2_X1 U797 ( .A1(n1096), .A2(n1101), .ZN(G63) );
XOR2_X1 U798 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND3_X1 U799 ( .A1(n1104), .A2(n1105), .A3(G478), .ZN(n1102) );
NAND2_X1 U800 ( .A1(KEYINPUT41), .A2(n1106), .ZN(n1105) );
NAND2_X1 U801 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
INV_X1 U802 ( .A(KEYINPUT41), .ZN(n1108) );
NAND2_X1 U803 ( .A1(n1056), .A2(G902), .ZN(n1107) );
NOR3_X1 U804 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(G60) );
AND2_X1 U805 ( .A1(KEYINPUT62), .A2(n1096), .ZN(n1111) );
NOR3_X1 U806 ( .A1(KEYINPUT62), .A2(G953), .A3(G952), .ZN(n1110) );
XNOR2_X1 U807 ( .A(n1112), .B(n1113), .ZN(n1109) );
NOR2_X1 U808 ( .A1(n1114), .A2(n1106), .ZN(n1113) );
XNOR2_X1 U809 ( .A(G104), .B(n1115), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1116), .A2(n1117), .ZN(G57) );
XOR2_X1 U811 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U812 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U813 ( .A(G101), .B(n1122), .ZN(n1121) );
AND2_X1 U814 ( .A1(G472), .A2(n1100), .ZN(n1120) );
XOR2_X1 U815 ( .A(n1123), .B(n1124), .Z(n1118) );
NOR2_X1 U816 ( .A1(n1125), .A2(KEYINPUT32), .ZN(n1124) );
INV_X1 U817 ( .A(n1126), .ZN(n1125) );
NAND2_X1 U818 ( .A1(n1127), .A2(n1128), .ZN(n1123) );
NAND2_X1 U819 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
OR3_X1 U820 ( .A1(n1131), .A2(n1132), .A3(n1130), .ZN(n1127) );
INV_X1 U821 ( .A(KEYINPUT15), .ZN(n1130) );
NOR2_X1 U822 ( .A1(n1133), .A2(n1091), .ZN(n1116) );
XNOR2_X1 U823 ( .A(G952), .B(KEYINPUT50), .ZN(n1133) );
NOR2_X1 U824 ( .A1(n1096), .A2(n1134), .ZN(G54) );
XOR2_X1 U825 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U826 ( .A(n1137), .B(n1138), .ZN(n1136) );
XOR2_X1 U827 ( .A(n1139), .B(n1140), .Z(n1135) );
XOR2_X1 U828 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U829 ( .A1(G110), .A2(KEYINPUT58), .ZN(n1142) );
AND2_X1 U830 ( .A1(G469), .A2(n1100), .ZN(n1141) );
NAND2_X1 U831 ( .A1(KEYINPUT28), .A2(n1143), .ZN(n1139) );
NOR2_X1 U832 ( .A1(n1096), .A2(n1144), .ZN(G51) );
XOR2_X1 U833 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U834 ( .A(KEYINPUT19), .B(n1147), .Z(n1146) );
NOR2_X1 U835 ( .A1(n1148), .A2(n1106), .ZN(n1147) );
INV_X1 U836 ( .A(n1100), .ZN(n1106) );
NOR2_X1 U837 ( .A1(n1149), .A2(n1056), .ZN(n1100) );
AND3_X1 U838 ( .A1(n1093), .A2(n1095), .A3(n1079), .ZN(n1056) );
AND4_X1 U839 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1079) );
AND4_X1 U840 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NOR2_X1 U841 ( .A1(n1158), .A2(n1159), .ZN(n1152) );
NOR3_X1 U842 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1159) );
XNOR2_X1 U843 ( .A(KEYINPUT14), .B(n1163), .ZN(n1162) );
NAND3_X1 U844 ( .A1(n1164), .A2(n1165), .A3(n1044), .ZN(n1160) );
XOR2_X1 U845 ( .A(KEYINPUT61), .B(n1166), .Z(n1164) );
AND4_X1 U846 ( .A1(n1115), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1093) );
AND4_X1 U847 ( .A1(n1015), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1169) );
NAND3_X1 U848 ( .A1(n1054), .A2(n1053), .A3(n1173), .ZN(n1015) );
NAND3_X1 U849 ( .A1(n1173), .A2(n1053), .A3(n1055), .ZN(n1115) );
XOR2_X1 U850 ( .A(n1174), .B(n1131), .Z(n1145) );
NOR2_X1 U851 ( .A1(n1091), .A2(G952), .ZN(n1096) );
XNOR2_X1 U852 ( .A(n1175), .B(n1158), .ZN(G48) );
AND3_X1 U853 ( .A1(n1176), .A2(n1055), .A3(n1177), .ZN(n1158) );
XNOR2_X1 U854 ( .A(G143), .B(n1150), .ZN(G45) );
NAND4_X1 U855 ( .A1(n1177), .A2(n1041), .A3(n1059), .A4(n1178), .ZN(n1150) );
INV_X1 U856 ( .A(n1179), .ZN(n1177) );
NAND2_X1 U857 ( .A1(n1180), .A2(n1181), .ZN(G42) );
NAND2_X1 U858 ( .A1(G140), .A2(n1182), .ZN(n1181) );
NAND2_X1 U859 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND2_X1 U860 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
INV_X1 U861 ( .A(KEYINPUT57), .ZN(n1186) );
XOR2_X1 U862 ( .A(n1151), .B(KEYINPUT2), .Z(n1183) );
NAND3_X1 U863 ( .A1(KEYINPUT57), .A2(n1185), .A3(n1187), .ZN(n1180) );
INV_X1 U864 ( .A(G140), .ZN(n1187) );
XOR2_X1 U865 ( .A(n1151), .B(KEYINPUT47), .Z(n1185) );
NAND3_X1 U866 ( .A1(n1055), .A2(n1040), .A3(n1188), .ZN(n1151) );
XNOR2_X1 U867 ( .A(G137), .B(n1157), .ZN(G39) );
NAND3_X1 U868 ( .A1(n1028), .A2(n1188), .A3(n1176), .ZN(n1157) );
XNOR2_X1 U869 ( .A(G134), .B(n1156), .ZN(G36) );
NAND3_X1 U870 ( .A1(n1188), .A2(n1054), .A3(n1041), .ZN(n1156) );
XOR2_X1 U871 ( .A(n1155), .B(n1189), .Z(G33) );
XNOR2_X1 U872 ( .A(G131), .B(KEYINPUT1), .ZN(n1189) );
NAND3_X1 U873 ( .A1(n1188), .A2(n1055), .A3(n1041), .ZN(n1155) );
AND3_X1 U874 ( .A1(n1044), .A2(n1165), .A3(n1052), .ZN(n1188) );
NOR2_X1 U875 ( .A1(n1034), .A2(n1038), .ZN(n1052) );
XOR2_X1 U876 ( .A(n1190), .B(n1191), .Z(G30) );
NOR3_X1 U877 ( .A1(n1179), .A2(n1161), .A3(n1163), .ZN(n1191) );
INV_X1 U878 ( .A(n1054), .ZN(n1161) );
NAND3_X1 U879 ( .A1(n1166), .A2(n1165), .A3(n1044), .ZN(n1179) );
XNOR2_X1 U880 ( .A(G128), .B(KEYINPUT55), .ZN(n1190) );
NAND3_X1 U881 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(G3) );
NAND2_X1 U882 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U883 ( .A1(n1197), .A2(n1198), .ZN(n1193) );
INV_X1 U884 ( .A(KEYINPUT53), .ZN(n1198) );
NAND2_X1 U885 ( .A1(n1199), .A2(G101), .ZN(n1197) );
XNOR2_X1 U886 ( .A(KEYINPUT63), .B(n1195), .ZN(n1199) );
NAND2_X1 U887 ( .A1(KEYINPUT53), .A2(n1200), .ZN(n1192) );
NAND2_X1 U888 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
OR3_X1 U889 ( .A1(n1196), .A2(n1195), .A3(KEYINPUT63), .ZN(n1202) );
NAND2_X1 U890 ( .A1(KEYINPUT63), .A2(n1195), .ZN(n1201) );
INV_X1 U891 ( .A(n1095), .ZN(n1195) );
NAND3_X1 U892 ( .A1(n1041), .A2(n1173), .A3(n1028), .ZN(n1095) );
XOR2_X1 U893 ( .A(G125), .B(n1203), .Z(G27) );
NOR2_X1 U894 ( .A1(KEYINPUT13), .A2(n1154), .ZN(n1203) );
NAND4_X1 U895 ( .A1(n1055), .A2(n1204), .A3(n1040), .A4(n1165), .ZN(n1154) );
NAND2_X1 U896 ( .A1(n1205), .A2(n1206), .ZN(n1165) );
NAND4_X1 U897 ( .A1(G953), .A2(G902), .A3(n1023), .A4(n1075), .ZN(n1206) );
INV_X1 U898 ( .A(G900), .ZN(n1075) );
XNOR2_X1 U899 ( .A(G122), .B(n1167), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1207), .A2(n1053), .A3(n1059), .A4(n1178), .ZN(n1167) );
NOR2_X1 U901 ( .A1(n1061), .A2(n1208), .ZN(n1053) );
XNOR2_X1 U902 ( .A(G119), .B(n1172), .ZN(G21) );
NAND3_X1 U903 ( .A1(n1176), .A2(n1028), .A3(n1207), .ZN(n1172) );
INV_X1 U904 ( .A(n1163), .ZN(n1176) );
NAND2_X1 U905 ( .A1(n1208), .A2(n1061), .ZN(n1163) );
XOR2_X1 U906 ( .A(n1209), .B(G116), .Z(G18) );
NAND2_X1 U907 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND4_X1 U908 ( .A1(n1204), .A2(n1054), .A3(n1212), .A4(n1213), .ZN(n1211) );
NOR2_X1 U909 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
INV_X1 U910 ( .A(n1041), .ZN(n1214) );
OR2_X1 U911 ( .A1(n1168), .A2(n1213), .ZN(n1210) );
INV_X1 U912 ( .A(KEYINPUT22), .ZN(n1213) );
NAND3_X1 U913 ( .A1(n1041), .A2(n1054), .A3(n1207), .ZN(n1168) );
AND2_X1 U914 ( .A1(n1204), .A2(n1215), .ZN(n1207) );
INV_X1 U915 ( .A(n1032), .ZN(n1204) );
NAND2_X1 U916 ( .A1(n1048), .A2(n1166), .ZN(n1032) );
NOR2_X1 U917 ( .A1(n1178), .A2(n1216), .ZN(n1054) );
INV_X1 U918 ( .A(n1059), .ZN(n1216) );
XOR2_X1 U919 ( .A(n1171), .B(n1217), .Z(G15) );
XNOR2_X1 U920 ( .A(G113), .B(KEYINPUT6), .ZN(n1217) );
NAND4_X1 U921 ( .A1(n1218), .A2(n1215), .A3(n1048), .A4(n1219), .ZN(n1171) );
AND2_X1 U922 ( .A1(n1055), .A2(n1041), .ZN(n1219) );
NOR2_X1 U923 ( .A1(n1061), .A2(n1220), .ZN(n1041) );
NOR2_X1 U924 ( .A1(n1059), .A2(n1221), .ZN(n1055) );
INV_X1 U925 ( .A(n1178), .ZN(n1221) );
INV_X1 U926 ( .A(n1037), .ZN(n1048) );
NAND2_X1 U927 ( .A1(n1222), .A2(n1047), .ZN(n1037) );
INV_X1 U928 ( .A(n1046), .ZN(n1222) );
XNOR2_X1 U929 ( .A(n1223), .B(n1224), .ZN(G12) );
NOR2_X1 U930 ( .A1(KEYINPUT49), .A2(n1170), .ZN(n1224) );
NAND3_X1 U931 ( .A1(n1040), .A2(n1173), .A3(n1028), .ZN(n1170) );
NOR2_X1 U932 ( .A1(n1059), .A2(n1178), .ZN(n1028) );
XOR2_X1 U933 ( .A(n1063), .B(n1225), .Z(n1178) );
XNOR2_X1 U934 ( .A(KEYINPUT31), .B(n1114), .ZN(n1225) );
INV_X1 U935 ( .A(G475), .ZN(n1114) );
AND2_X1 U936 ( .A1(n1226), .A2(n1112), .ZN(n1063) );
XNOR2_X1 U937 ( .A(n1227), .B(n1228), .ZN(n1112) );
XOR2_X1 U938 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U939 ( .A(n1231), .B(G113), .ZN(n1230) );
XNOR2_X1 U940 ( .A(n1232), .B(G131), .ZN(n1229) );
XOR2_X1 U941 ( .A(n1233), .B(n1234), .Z(n1227) );
NOR4_X1 U942 ( .A1(KEYINPUT33), .A2(G953), .A3(G237), .A4(n1235), .ZN(n1234) );
INV_X1 U943 ( .A(G214), .ZN(n1235) );
XNOR2_X1 U944 ( .A(n1236), .B(n1237), .ZN(n1233) );
NAND2_X1 U945 ( .A1(n1238), .A2(n1239), .ZN(n1236) );
XOR2_X1 U946 ( .A(n1240), .B(KEYINPUT42), .Z(n1238) );
XNOR2_X1 U947 ( .A(KEYINPUT20), .B(n1241), .ZN(n1226) );
XNOR2_X1 U948 ( .A(n1242), .B(G478), .ZN(n1059) );
NAND2_X1 U949 ( .A1(n1103), .A2(n1241), .ZN(n1242) );
XOR2_X1 U950 ( .A(n1243), .B(n1244), .Z(n1103) );
XNOR2_X1 U951 ( .A(n1245), .B(n1246), .ZN(n1244) );
XOR2_X1 U952 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U953 ( .A1(KEYINPUT23), .A2(n1249), .ZN(n1248) );
XNOR2_X1 U954 ( .A(G128), .B(n1250), .ZN(n1249) );
NAND2_X1 U955 ( .A1(KEYINPUT46), .A2(n1232), .ZN(n1250) );
INV_X1 U956 ( .A(G143), .ZN(n1232) );
NAND2_X1 U957 ( .A1(G217), .A2(n1251), .ZN(n1247) );
XNOR2_X1 U958 ( .A(G107), .B(n1252), .ZN(n1243) );
XNOR2_X1 U959 ( .A(n1231), .B(G116), .ZN(n1252) );
AND3_X1 U960 ( .A1(n1218), .A2(n1215), .A3(n1044), .ZN(n1173) );
AND2_X1 U961 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NAND2_X1 U962 ( .A1(G221), .A2(n1253), .ZN(n1047) );
XNOR2_X1 U963 ( .A(n1254), .B(n1255), .ZN(n1046) );
XOR2_X1 U964 ( .A(KEYINPUT21), .B(G469), .Z(n1255) );
NAND2_X1 U965 ( .A1(n1241), .A2(n1256), .ZN(n1254) );
XOR2_X1 U966 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U967 ( .A(n1259), .B(n1260), .Z(n1258) );
XNOR2_X1 U968 ( .A(G110), .B(KEYINPUT45), .ZN(n1260) );
NAND2_X1 U969 ( .A1(KEYINPUT34), .A2(n1137), .ZN(n1259) );
XOR2_X1 U970 ( .A(n1138), .B(n1261), .Z(n1257) );
NOR2_X1 U971 ( .A1(n1143), .A2(KEYINPUT5), .ZN(n1261) );
AND2_X1 U972 ( .A1(n1262), .A2(n1263), .ZN(n1143) );
NAND2_X1 U973 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XNOR2_X1 U974 ( .A(KEYINPUT43), .B(n1196), .ZN(n1265) );
XNOR2_X1 U975 ( .A(G104), .B(G107), .ZN(n1264) );
NAND2_X1 U976 ( .A1(n1266), .A2(n1267), .ZN(n1262) );
XNOR2_X1 U977 ( .A(n1268), .B(G104), .ZN(n1267) );
INV_X1 U978 ( .A(G107), .ZN(n1268) );
XNOR2_X1 U979 ( .A(G101), .B(KEYINPUT4), .ZN(n1266) );
XNOR2_X1 U980 ( .A(n1078), .B(n1269), .ZN(n1138) );
AND2_X1 U981 ( .A1(n1091), .A2(G227), .ZN(n1269) );
AND2_X1 U982 ( .A1(n1270), .A2(n1271), .ZN(n1078) );
NAND2_X1 U983 ( .A1(n1272), .A2(n1175), .ZN(n1271) );
NAND2_X1 U984 ( .A1(n1273), .A2(G146), .ZN(n1270) );
XOR2_X1 U985 ( .A(KEYINPUT27), .B(n1272), .Z(n1273) );
XNOR2_X1 U986 ( .A(n1274), .B(G143), .ZN(n1272) );
NAND2_X1 U987 ( .A1(n1205), .A2(n1275), .ZN(n1215) );
NAND3_X1 U988 ( .A1(G902), .A2(n1023), .A3(n1088), .ZN(n1275) );
NOR2_X1 U989 ( .A1(n1091), .A2(G898), .ZN(n1088) );
NAND3_X1 U990 ( .A1(n1023), .A2(n1091), .A3(G952), .ZN(n1205) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1023) );
XNOR2_X1 U992 ( .A(n1166), .B(KEYINPUT44), .ZN(n1218) );
NOR2_X1 U993 ( .A1(n1276), .A2(n1038), .ZN(n1166) );
INV_X1 U994 ( .A(n1049), .ZN(n1038) );
NAND2_X1 U995 ( .A1(G214), .A2(n1277), .ZN(n1049) );
INV_X1 U996 ( .A(n1034), .ZN(n1276) );
XOR2_X1 U997 ( .A(n1278), .B(n1148), .Z(n1034) );
NAND2_X1 U998 ( .A1(G210), .A2(n1277), .ZN(n1148) );
NAND2_X1 U999 ( .A1(n1279), .A2(n1149), .ZN(n1277) );
NAND2_X1 U1000 ( .A1(n1280), .A2(n1241), .ZN(n1278) );
XOR2_X1 U1001 ( .A(n1174), .B(n1281), .Z(n1280) );
XNOR2_X1 U1002 ( .A(n1282), .B(KEYINPUT11), .ZN(n1281) );
NAND2_X1 U1003 ( .A1(KEYINPUT26), .A2(n1131), .ZN(n1282) );
XNOR2_X1 U1004 ( .A(n1283), .B(n1284), .ZN(n1131) );
XOR2_X1 U1005 ( .A(n1285), .B(n1286), .Z(n1174) );
XNOR2_X1 U1006 ( .A(n1287), .B(n1090), .ZN(n1286) );
XOR2_X1 U1007 ( .A(n1288), .B(n1223), .Z(n1090) );
NAND2_X1 U1008 ( .A1(KEYINPUT54), .A2(n1231), .ZN(n1288) );
INV_X1 U1009 ( .A(G122), .ZN(n1231) );
NAND2_X1 U1010 ( .A1(G224), .A2(n1091), .ZN(n1287) );
XOR2_X1 U1011 ( .A(n1289), .B(G125), .Z(n1285) );
NAND2_X1 U1012 ( .A1(KEYINPUT40), .A2(n1089), .ZN(n1289) );
XNOR2_X1 U1013 ( .A(n1290), .B(n1291), .ZN(n1089) );
NOR2_X1 U1014 ( .A1(KEYINPUT16), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U1015 ( .A(n1293), .B(n1294), .ZN(n1290) );
NAND2_X1 U1016 ( .A1(n1295), .A2(n1296), .ZN(n1293) );
NAND2_X1 U1017 ( .A1(G101), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1018 ( .A(n1298), .B(KEYINPUT10), .Z(n1295) );
OR2_X1 U1019 ( .A1(n1297), .A2(G101), .ZN(n1298) );
NAND2_X1 U1020 ( .A1(n1299), .A2(n1300), .ZN(n1297) );
NAND2_X1 U1021 ( .A1(n1301), .A2(n1237), .ZN(n1300) );
XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n1302), .Z(n1299) );
NOR2_X1 U1023 ( .A1(n1301), .A2(n1237), .ZN(n1302) );
INV_X1 U1024 ( .A(G104), .ZN(n1237) );
XNOR2_X1 U1025 ( .A(KEYINPUT59), .B(G107), .ZN(n1301) );
AND2_X1 U1026 ( .A1(n1220), .A2(n1061), .ZN(n1040) );
XNOR2_X1 U1027 ( .A(n1303), .B(n1304), .ZN(n1061) );
AND2_X1 U1028 ( .A1(n1253), .A2(G217), .ZN(n1304) );
NAND2_X1 U1029 ( .A1(n1305), .A2(n1149), .ZN(n1253) );
XOR2_X1 U1030 ( .A(KEYINPUT56), .B(G234), .Z(n1305) );
NAND2_X1 U1031 ( .A1(n1099), .A2(n1241), .ZN(n1303) );
XOR2_X1 U1032 ( .A(n1306), .B(n1307), .Z(n1099) );
AND2_X1 U1033 ( .A1(G221), .A2(n1251), .ZN(n1307) );
AND2_X1 U1034 ( .A1(G234), .A2(n1091), .ZN(n1251) );
XOR2_X1 U1035 ( .A(n1308), .B(G137), .Z(n1306) );
NAND2_X1 U1036 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND3_X1 U1037 ( .A1(n1239), .A2(n1240), .A3(n1311), .ZN(n1310) );
XOR2_X1 U1038 ( .A(KEYINPUT7), .B(n1312), .Z(n1309) );
NOR2_X1 U1039 ( .A1(n1313), .A2(n1311), .ZN(n1312) );
NAND3_X1 U1040 ( .A1(n1314), .A2(n1315), .A3(n1316), .ZN(n1311) );
NAND2_X1 U1041 ( .A1(G110), .A2(n1317), .ZN(n1316) );
NAND2_X1 U1042 ( .A1(n1318), .A2(n1319), .ZN(n1315) );
INV_X1 U1043 ( .A(KEYINPUT17), .ZN(n1319) );
NAND2_X1 U1044 ( .A1(n1320), .A2(n1321), .ZN(n1318) );
XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n1223), .ZN(n1321) );
NAND2_X1 U1046 ( .A1(KEYINPUT17), .A2(n1322), .ZN(n1314) );
NAND2_X1 U1047 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND3_X1 U1048 ( .A1(KEYINPUT52), .A2(n1320), .A3(n1223), .ZN(n1324) );
INV_X1 U1049 ( .A(n1317), .ZN(n1320) );
XNOR2_X1 U1050 ( .A(G119), .B(n1284), .ZN(n1317) );
INV_X1 U1051 ( .A(G128), .ZN(n1284) );
OR2_X1 U1052 ( .A1(n1223), .A2(KEYINPUT52), .ZN(n1323) );
AND2_X1 U1053 ( .A1(n1239), .A2(n1240), .ZN(n1313) );
NAND2_X1 U1054 ( .A1(n1077), .A2(G146), .ZN(n1240) );
OR2_X1 U1055 ( .A1(n1077), .A2(G146), .ZN(n1239) );
XOR2_X1 U1056 ( .A(G125), .B(n1325), .Z(n1077) );
INV_X1 U1057 ( .A(n1137), .ZN(n1325) );
XOR2_X1 U1058 ( .A(G140), .B(KEYINPUT25), .Z(n1137) );
INV_X1 U1059 ( .A(n1208), .ZN(n1220) );
XNOR2_X1 U1060 ( .A(n1064), .B(G472), .ZN(n1208) );
NAND2_X1 U1061 ( .A1(n1241), .A2(n1326), .ZN(n1064) );
XOR2_X1 U1062 ( .A(n1129), .B(n1327), .Z(n1326) );
XOR2_X1 U1063 ( .A(n1328), .B(n1329), .Z(n1327) );
NOR2_X1 U1064 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XOR2_X1 U1065 ( .A(n1332), .B(KEYINPUT18), .Z(n1331) );
NAND2_X1 U1066 ( .A1(n1196), .A2(n1126), .ZN(n1332) );
NOR2_X1 U1067 ( .A1(n1196), .A2(n1126), .ZN(n1330) );
NAND3_X1 U1068 ( .A1(n1279), .A2(n1091), .A3(G210), .ZN(n1126) );
INV_X1 U1069 ( .A(G953), .ZN(n1091) );
INV_X1 U1070 ( .A(G237), .ZN(n1279) );
INV_X1 U1071 ( .A(G101), .ZN(n1196) );
NOR2_X1 U1072 ( .A1(KEYINPUT0), .A2(n1122), .ZN(n1328) );
NAND2_X1 U1073 ( .A1(n1333), .A2(n1334), .ZN(n1122) );
NAND2_X1 U1074 ( .A1(n1292), .A2(n1294), .ZN(n1334) );
XOR2_X1 U1075 ( .A(n1335), .B(KEYINPUT8), .Z(n1333) );
OR2_X1 U1076 ( .A1(n1294), .A2(n1292), .ZN(n1335) );
XOR2_X1 U1077 ( .A(G116), .B(n1336), .Z(n1292) );
INV_X1 U1078 ( .A(G119), .ZN(n1336) );
INV_X1 U1079 ( .A(G113), .ZN(n1294) );
XNOR2_X1 U1080 ( .A(n1274), .B(n1283), .ZN(n1129) );
XOR2_X1 U1081 ( .A(G143), .B(n1337), .Z(n1283) );
XNOR2_X1 U1082 ( .A(KEYINPUT29), .B(n1175), .ZN(n1337) );
INV_X1 U1083 ( .A(G146), .ZN(n1175) );
XNOR2_X1 U1084 ( .A(G128), .B(n1132), .ZN(n1274) );
XNOR2_X1 U1085 ( .A(n1338), .B(n1245), .ZN(n1132) );
XOR2_X1 U1086 ( .A(G134), .B(KEYINPUT39), .Z(n1245) );
XNOR2_X1 U1087 ( .A(G131), .B(G137), .ZN(n1338) );
XOR2_X1 U1088 ( .A(n1149), .B(KEYINPUT60), .Z(n1241) );
INV_X1 U1089 ( .A(G902), .ZN(n1149) );
INV_X1 U1090 ( .A(G110), .ZN(n1223) );
endmodule


