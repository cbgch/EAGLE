//Key = 1111010000010111100110111100000101001111101001011100010010100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354;

XNOR2_X1 U746 ( .A(G107), .B(n1027), .ZN(G9) );
NOR2_X1 U747 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U748 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
NOR2_X1 U749 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NAND4_X1 U750 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1030) );
NAND3_X1 U751 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1037) );
XNOR2_X1 U752 ( .A(KEYINPUT30), .B(n1035), .ZN(n1041) );
NAND4_X1 U753 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1035) );
NAND3_X1 U754 ( .A1(n1047), .A2(n1048), .A3(n1043), .ZN(n1036) );
INV_X1 U755 ( .A(n1049), .ZN(n1043) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND4_X1 U757 ( .A1(n1052), .A2(n1046), .A3(n1044), .A4(n1053), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND3_X1 U759 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1047) );
NAND3_X1 U760 ( .A1(n1046), .A2(n1059), .A3(n1045), .ZN(n1057) );
OR2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U762 ( .A1(n1044), .A2(n1062), .ZN(n1056) );
NAND3_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NAND2_X1 U764 ( .A1(n1066), .A2(n1045), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1046), .A2(n1067), .ZN(n1063) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U767 ( .A1(n1052), .A2(n1055), .A3(n1070), .ZN(n1069) );
INV_X1 U768 ( .A(KEYINPUT21), .ZN(n1055) );
INV_X1 U769 ( .A(n1071), .ZN(n1068) );
AND3_X1 U770 ( .A1(n1038), .A2(n1039), .A3(n1072), .ZN(n1028) );
NAND4_X1 U771 ( .A1(n1073), .A2(n1045), .A3(n1074), .A4(n1075), .ZN(n1038) );
NOR4_X1 U772 ( .A1(n1076), .A2(n1077), .A3(n1051), .A4(n1078), .ZN(n1075) );
NOR2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
AND3_X1 U774 ( .A1(KEYINPUT11), .A2(n1081), .A3(n1082), .ZN(n1080) );
NOR2_X1 U775 ( .A1(KEYINPUT11), .A2(n1082), .ZN(n1079) );
XNOR2_X1 U776 ( .A(n1083), .B(n1084), .ZN(n1073) );
XOR2_X1 U777 ( .A(n1085), .B(n1086), .Z(G72) );
XOR2_X1 U778 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U780 ( .A1(G953), .A2(n1091), .ZN(n1090) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(n1089) );
XNOR2_X1 U782 ( .A(n1094), .B(n1095), .ZN(n1093) );
NAND2_X1 U783 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
OR2_X1 U784 ( .A1(n1098), .A2(KEYINPUT60), .ZN(n1097) );
NAND3_X1 U785 ( .A1(G131), .A2(n1099), .A3(KEYINPUT60), .ZN(n1096) );
XNOR2_X1 U786 ( .A(G125), .B(n1100), .ZN(n1092) );
XNOR2_X1 U787 ( .A(KEYINPUT1), .B(n1101), .ZN(n1100) );
INV_X1 U788 ( .A(G140), .ZN(n1101) );
NAND2_X1 U789 ( .A1(G953), .A2(n1102), .ZN(n1087) );
NAND2_X1 U790 ( .A1(n1103), .A2(G227), .ZN(n1102) );
XNOR2_X1 U791 ( .A(G900), .B(KEYINPUT38), .ZN(n1103) );
AND2_X1 U792 ( .A1(n1033), .A2(n1039), .ZN(n1085) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(G69) );
NAND4_X1 U794 ( .A1(G953), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1105) );
NAND2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
NAND2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND3_X1 U797 ( .A1(n1113), .A2(n1106), .A3(G953), .ZN(n1112) );
NAND2_X1 U798 ( .A1(n1108), .A2(n1114), .ZN(n1113) );
INV_X1 U799 ( .A(KEYINPUT4), .ZN(n1108) );
NAND2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U801 ( .A1(G953), .A2(n1106), .ZN(n1115) );
NAND2_X1 U802 ( .A1(G224), .A2(n1116), .ZN(n1106) );
XNOR2_X1 U803 ( .A(KEYINPUT10), .B(n1117), .ZN(n1116) );
INV_X1 U804 ( .A(KEYINPUT6), .ZN(n1114) );
XNOR2_X1 U805 ( .A(n1107), .B(n1118), .ZN(n1109) );
NOR2_X1 U806 ( .A1(G953), .A2(n1119), .ZN(n1118) );
XNOR2_X1 U807 ( .A(KEYINPUT44), .B(n1031), .ZN(n1119) );
NAND2_X1 U808 ( .A1(n1120), .A2(n1121), .ZN(n1107) );
NAND2_X1 U809 ( .A1(G953), .A2(n1117), .ZN(n1121) );
XOR2_X1 U810 ( .A(n1122), .B(n1123), .Z(n1120) );
NOR2_X1 U811 ( .A1(KEYINPUT29), .A2(n1124), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XOR2_X1 U813 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U814 ( .A1(KEYINPUT34), .A2(n1129), .ZN(n1128) );
NAND2_X1 U815 ( .A1(n1130), .A2(n1082), .ZN(n1127) );
NOR2_X1 U816 ( .A1(n1125), .A2(n1131), .ZN(G63) );
XOR2_X1 U817 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U818 ( .A1(n1084), .A2(n1134), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1125), .A2(n1135), .ZN(G60) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
XNOR2_X1 U821 ( .A(KEYINPUT55), .B(n1138), .ZN(n1137) );
AND2_X1 U822 ( .A1(G475), .A2(n1130), .ZN(n1136) );
XOR2_X1 U823 ( .A(G104), .B(n1139), .Z(G6) );
NOR2_X1 U824 ( .A1(KEYINPUT28), .A2(n1140), .ZN(n1139) );
NOR2_X1 U825 ( .A1(n1125), .A2(n1141), .ZN(G57) );
XOR2_X1 U826 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U827 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U828 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U829 ( .A(KEYINPUT7), .B(n1148), .Z(n1147) );
NOR2_X1 U830 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U831 ( .A1(n1098), .A2(n1151), .ZN(n1146) );
AND2_X1 U832 ( .A1(G472), .A2(n1130), .ZN(n1144) );
XNOR2_X1 U833 ( .A(n1152), .B(n1153), .ZN(n1142) );
XNOR2_X1 U834 ( .A(G101), .B(n1154), .ZN(n1153) );
NOR2_X1 U835 ( .A1(n1125), .A2(n1155), .ZN(G54) );
XOR2_X1 U836 ( .A(n1156), .B(n1157), .Z(n1155) );
XNOR2_X1 U837 ( .A(n1158), .B(n1159), .ZN(n1157) );
NAND2_X1 U838 ( .A1(KEYINPUT24), .A2(n1160), .ZN(n1158) );
NAND2_X1 U839 ( .A1(n1130), .A2(G469), .ZN(n1160) );
INV_X1 U840 ( .A(n1134), .ZN(n1130) );
XOR2_X1 U841 ( .A(n1161), .B(n1162), .Z(n1156) );
NOR2_X1 U842 ( .A1(KEYINPUT26), .A2(n1163), .ZN(n1162) );
XOR2_X1 U843 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U844 ( .A(n1149), .B(KEYINPUT22), .ZN(n1165) );
NAND3_X1 U845 ( .A1(G227), .A2(n1039), .A3(KEYINPUT20), .ZN(n1161) );
NOR2_X1 U846 ( .A1(n1166), .A2(n1167), .ZN(G51) );
XOR2_X1 U847 ( .A(KEYINPUT12), .B(n1125), .Z(n1167) );
AND2_X1 U848 ( .A1(n1168), .A2(n1072), .ZN(n1125) );
INV_X1 U849 ( .A(G952), .ZN(n1072) );
XNOR2_X1 U850 ( .A(G953), .B(KEYINPUT63), .ZN(n1168) );
XNOR2_X1 U851 ( .A(n1169), .B(n1170), .ZN(n1166) );
XOR2_X1 U852 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U853 ( .A1(n1173), .A2(n1134), .ZN(n1172) );
NAND2_X1 U854 ( .A1(G902), .A2(n1174), .ZN(n1134) );
OR2_X1 U855 ( .A1(n1031), .A2(n1033), .ZN(n1174) );
NAND2_X1 U856 ( .A1(n1175), .A2(n1176), .ZN(n1033) );
NOR4_X1 U857 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NOR2_X1 U858 ( .A1(KEYINPUT46), .A2(n1181), .ZN(n1179) );
NOR2_X1 U859 ( .A1(n1182), .A2(n1183), .ZN(n1178) );
NOR2_X1 U860 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
AND3_X1 U861 ( .A1(KEYINPUT46), .A2(n1051), .A3(n1186), .ZN(n1185) );
AND3_X1 U862 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1184) );
INV_X1 U863 ( .A(n1190), .ZN(n1177) );
NOR4_X1 U864 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1175) );
AND3_X1 U865 ( .A1(n1186), .A2(n1195), .A3(n1189), .ZN(n1194) );
INV_X1 U866 ( .A(n1196), .ZN(n1192) );
INV_X1 U867 ( .A(n1197), .ZN(n1191) );
NAND2_X1 U868 ( .A1(n1198), .A2(n1199), .ZN(n1031) );
AND4_X1 U869 ( .A1(n1027), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1199) );
NAND3_X1 U870 ( .A1(n1046), .A2(n1060), .A3(n1203), .ZN(n1027) );
NOR4_X1 U871 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1198) );
AND3_X1 U872 ( .A1(n1208), .A2(n1195), .A3(n1046), .ZN(n1207) );
INV_X1 U873 ( .A(n1140), .ZN(n1206) );
NAND3_X1 U874 ( .A1(n1203), .A2(n1046), .A3(n1061), .ZN(n1140) );
NAND2_X1 U875 ( .A1(n1209), .A2(n1210), .ZN(n1171) );
NAND2_X1 U876 ( .A1(n1211), .A2(n1151), .ZN(n1209) );
XNOR2_X1 U877 ( .A(n1212), .B(KEYINPUT37), .ZN(n1211) );
NAND2_X1 U878 ( .A1(n1213), .A2(n1214), .ZN(G48) );
NAND2_X1 U879 ( .A1(n1193), .A2(n1215), .ZN(n1214) );
XOR2_X1 U880 ( .A(KEYINPUT45), .B(n1216), .Z(n1213) );
NOR2_X1 U881 ( .A1(n1193), .A2(n1215), .ZN(n1216) );
AND2_X1 U882 ( .A1(n1217), .A2(n1061), .ZN(n1193) );
XOR2_X1 U883 ( .A(n1218), .B(n1219), .Z(G45) );
NOR3_X1 U884 ( .A1(n1220), .A2(n1221), .A3(n1034), .ZN(n1219) );
XNOR2_X1 U885 ( .A(n1195), .B(KEYINPUT43), .ZN(n1221) );
NAND2_X1 U886 ( .A1(KEYINPUT16), .A2(n1222), .ZN(n1218) );
XNOR2_X1 U887 ( .A(G140), .B(n1190), .ZN(G42) );
NAND4_X1 U888 ( .A1(n1223), .A2(n1061), .A3(n1224), .A4(n1058), .ZN(n1190) );
NAND2_X1 U889 ( .A1(n1225), .A2(n1226), .ZN(G39) );
OR2_X1 U890 ( .A1(n1196), .A2(G137), .ZN(n1226) );
XOR2_X1 U891 ( .A(n1227), .B(KEYINPUT9), .Z(n1225) );
NAND2_X1 U892 ( .A1(G137), .A2(n1196), .ZN(n1227) );
NAND4_X1 U893 ( .A1(n1223), .A2(n1044), .A3(n1058), .A4(n1077), .ZN(n1196) );
NAND2_X1 U894 ( .A1(n1228), .A2(n1229), .ZN(G36) );
OR2_X1 U895 ( .A1(n1197), .A2(G134), .ZN(n1229) );
XOR2_X1 U896 ( .A(n1230), .B(KEYINPUT27), .Z(n1228) );
NAND2_X1 U897 ( .A1(G134), .A2(n1197), .ZN(n1230) );
NAND3_X1 U898 ( .A1(n1058), .A2(n1060), .A3(n1186), .ZN(n1197) );
XNOR2_X1 U899 ( .A(n1231), .B(n1181), .ZN(G33) );
NAND3_X1 U900 ( .A1(n1061), .A2(n1058), .A3(n1186), .ZN(n1181) );
INV_X1 U901 ( .A(n1220), .ZN(n1186) );
NAND3_X1 U902 ( .A1(n1071), .A2(n1188), .A3(n1066), .ZN(n1220) );
INV_X1 U903 ( .A(n1051), .ZN(n1058) );
NAND2_X1 U904 ( .A1(n1040), .A2(n1232), .ZN(n1051) );
XNOR2_X1 U905 ( .A(G131), .B(KEYINPUT33), .ZN(n1231) );
XNOR2_X1 U906 ( .A(n1233), .B(n1180), .ZN(G30) );
AND2_X1 U907 ( .A1(n1217), .A2(n1060), .ZN(n1180) );
AND3_X1 U908 ( .A1(n1189), .A2(n1077), .A3(n1223), .ZN(n1217) );
AND3_X1 U909 ( .A1(n1234), .A2(n1188), .A3(n1071), .ZN(n1223) );
XOR2_X1 U910 ( .A(n1205), .B(n1235), .Z(G3) );
NOR2_X1 U911 ( .A1(KEYINPUT35), .A2(n1236), .ZN(n1235) );
AND3_X1 U912 ( .A1(n1044), .A2(n1203), .A3(n1066), .ZN(n1205) );
XOR2_X1 U913 ( .A(n1237), .B(n1238), .Z(G27) );
NAND2_X1 U914 ( .A1(KEYINPUT23), .A2(G125), .ZN(n1238) );
NAND4_X1 U915 ( .A1(n1239), .A2(n1187), .A3(n1061), .A4(n1188), .ZN(n1237) );
NAND2_X1 U916 ( .A1(n1049), .A2(n1240), .ZN(n1188) );
NAND4_X1 U917 ( .A1(n1241), .A2(G902), .A3(n1242), .A4(n1091), .ZN(n1240) );
INV_X1 U918 ( .A(G900), .ZN(n1091) );
XNOR2_X1 U919 ( .A(G953), .B(KEYINPUT15), .ZN(n1241) );
INV_X1 U920 ( .A(n1064), .ZN(n1187) );
NAND3_X1 U921 ( .A1(n1224), .A2(n1234), .A3(n1045), .ZN(n1064) );
XNOR2_X1 U922 ( .A(n1034), .B(KEYINPUT62), .ZN(n1239) );
XOR2_X1 U923 ( .A(n1243), .B(n1244), .Z(G24) );
NOR2_X1 U924 ( .A1(G122), .A2(KEYINPUT59), .ZN(n1244) );
NAND4_X1 U925 ( .A1(n1245), .A2(n1046), .A3(n1195), .A4(n1246), .ZN(n1243) );
XNOR2_X1 U926 ( .A(KEYINPUT36), .B(n1189), .ZN(n1246) );
NOR2_X1 U927 ( .A1(n1247), .A2(n1077), .ZN(n1046) );
XOR2_X1 U928 ( .A(G119), .B(n1204), .Z(G21) );
AND4_X1 U929 ( .A1(n1208), .A2(n1044), .A3(n1234), .A4(n1077), .ZN(n1204) );
XOR2_X1 U930 ( .A(G116), .B(n1248), .Z(G18) );
NOR2_X1 U931 ( .A1(KEYINPUT61), .A2(n1202), .ZN(n1248) );
NAND3_X1 U932 ( .A1(n1066), .A2(n1060), .A3(n1208), .ZN(n1202) );
AND2_X1 U933 ( .A1(n1189), .A2(n1245), .ZN(n1208) );
INV_X1 U934 ( .A(n1034), .ZN(n1189) );
XOR2_X1 U935 ( .A(n1249), .B(KEYINPUT58), .Z(n1034) );
NAND2_X1 U936 ( .A1(n1250), .A2(n1251), .ZN(n1060) );
OR3_X1 U937 ( .A1(n1252), .A2(n1078), .A3(KEYINPUT51), .ZN(n1251) );
NAND2_X1 U938 ( .A1(KEYINPUT51), .A2(n1195), .ZN(n1250) );
NOR2_X1 U939 ( .A1(n1252), .A2(n1253), .ZN(n1195) );
INV_X1 U940 ( .A(n1078), .ZN(n1253) );
XNOR2_X1 U941 ( .A(G113), .B(n1201), .ZN(G15) );
NAND4_X1 U942 ( .A1(n1066), .A2(n1245), .A3(n1061), .A4(n1249), .ZN(n1201) );
INV_X1 U943 ( .A(n1183), .ZN(n1061) );
NAND2_X1 U944 ( .A1(n1252), .A2(n1078), .ZN(n1183) );
AND2_X1 U945 ( .A1(n1045), .A2(n1254), .ZN(n1245) );
NOR2_X1 U946 ( .A1(n1255), .A2(n1070), .ZN(n1045) );
NOR2_X1 U947 ( .A1(n1247), .A2(n1224), .ZN(n1066) );
XNOR2_X1 U948 ( .A(G110), .B(n1200), .ZN(G12) );
NAND4_X1 U949 ( .A1(n1044), .A2(n1203), .A3(n1224), .A4(n1234), .ZN(n1200) );
XNOR2_X1 U950 ( .A(n1247), .B(KEYINPUT13), .ZN(n1234) );
OR2_X1 U951 ( .A1(n1076), .A2(n1256), .ZN(n1247) );
AND2_X1 U952 ( .A1(n1082), .A2(n1081), .ZN(n1256) );
NOR2_X1 U953 ( .A1(n1081), .A2(n1082), .ZN(n1076) );
AND2_X1 U954 ( .A1(G217), .A2(n1257), .ZN(n1082) );
OR2_X1 U955 ( .A1(n1129), .A2(G902), .ZN(n1081) );
XOR2_X1 U956 ( .A(n1258), .B(n1259), .Z(n1129) );
XOR2_X1 U957 ( .A(n1260), .B(n1261), .Z(n1259) );
XNOR2_X1 U958 ( .A(n1233), .B(G119), .ZN(n1261) );
XNOR2_X1 U959 ( .A(n1215), .B(G137), .ZN(n1260) );
INV_X1 U960 ( .A(G146), .ZN(n1215) );
XOR2_X1 U961 ( .A(n1262), .B(n1159), .Z(n1258) );
XOR2_X1 U962 ( .A(n1263), .B(n1264), .Z(n1262) );
NAND2_X1 U963 ( .A1(n1265), .A2(G221), .ZN(n1263) );
INV_X1 U964 ( .A(n1077), .ZN(n1224) );
XNOR2_X1 U965 ( .A(n1266), .B(G472), .ZN(n1077) );
NAND2_X1 U966 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
XOR2_X1 U967 ( .A(n1269), .B(n1270), .Z(n1267) );
XNOR2_X1 U968 ( .A(G101), .B(n1271), .ZN(n1270) );
NAND2_X1 U969 ( .A1(KEYINPUT40), .A2(n1272), .ZN(n1271) );
XOR2_X1 U970 ( .A(n1154), .B(n1273), .Z(n1272) );
NAND2_X1 U971 ( .A1(n1274), .A2(KEYINPUT5), .ZN(n1273) );
XNOR2_X1 U972 ( .A(n1151), .B(n1098), .ZN(n1274) );
INV_X1 U973 ( .A(n1149), .ZN(n1098) );
NAND3_X1 U974 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1154) );
NAND2_X1 U975 ( .A1(G113), .A2(n1278), .ZN(n1277) );
NAND3_X1 U976 ( .A1(n1279), .A2(n1280), .A3(KEYINPUT31), .ZN(n1276) );
INV_X1 U977 ( .A(n1278), .ZN(n1279) );
NAND2_X1 U978 ( .A1(KEYINPUT56), .A2(n1281), .ZN(n1278) );
OR2_X1 U979 ( .A1(n1281), .A2(KEYINPUT31), .ZN(n1275) );
NAND2_X1 U980 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U981 ( .A1(G119), .A2(n1284), .ZN(n1283) );
XOR2_X1 U982 ( .A(n1285), .B(KEYINPUT32), .Z(n1282) );
OR2_X1 U983 ( .A1(n1284), .A2(G119), .ZN(n1285) );
XOR2_X1 U984 ( .A(G116), .B(KEYINPUT49), .Z(n1284) );
NOR2_X1 U985 ( .A1(KEYINPUT52), .A2(n1152), .ZN(n1269) );
NAND3_X1 U986 ( .A1(n1286), .A2(n1039), .A3(G210), .ZN(n1152) );
AND3_X1 U987 ( .A1(n1249), .A2(n1254), .A3(n1071), .ZN(n1203) );
NOR2_X1 U988 ( .A1(n1052), .A2(n1070), .ZN(n1071) );
INV_X1 U989 ( .A(n1054), .ZN(n1070) );
NAND2_X1 U990 ( .A1(G221), .A2(n1257), .ZN(n1054) );
NAND2_X1 U991 ( .A1(G234), .A2(n1268), .ZN(n1257) );
INV_X1 U992 ( .A(n1255), .ZN(n1052) );
XNOR2_X1 U993 ( .A(n1287), .B(G469), .ZN(n1255) );
NAND2_X1 U994 ( .A1(n1288), .A2(n1268), .ZN(n1287) );
XOR2_X1 U995 ( .A(n1159), .B(n1289), .Z(n1288) );
XOR2_X1 U996 ( .A(n1290), .B(n1291), .Z(n1289) );
NOR2_X1 U997 ( .A1(KEYINPUT57), .A2(n1292), .ZN(n1291) );
INV_X1 U998 ( .A(G227), .ZN(n1292) );
NOR2_X1 U999 ( .A1(n1293), .A2(n1294), .ZN(n1290) );
XOR2_X1 U1000 ( .A(n1295), .B(KEYINPUT0), .Z(n1294) );
NAND2_X1 U1001 ( .A1(n1164), .A2(n1149), .ZN(n1295) );
NOR2_X1 U1002 ( .A1(n1164), .A2(n1149), .ZN(n1293) );
XOR2_X1 U1003 ( .A(G131), .B(n1099), .Z(n1149) );
XOR2_X1 U1004 ( .A(G134), .B(G137), .Z(n1099) );
XOR2_X1 U1005 ( .A(n1296), .B(n1297), .Z(n1164) );
NOR2_X1 U1006 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NOR2_X1 U1007 ( .A1(KEYINPUT41), .A2(n1300), .ZN(n1299) );
NOR2_X1 U1008 ( .A1(KEYINPUT42), .A2(n1301), .ZN(n1298) );
INV_X1 U1009 ( .A(n1300), .ZN(n1301) );
XOR2_X1 U1010 ( .A(G104), .B(n1302), .Z(n1300) );
NOR2_X1 U1011 ( .A1(G107), .A2(KEYINPUT54), .ZN(n1302) );
XNOR2_X1 U1012 ( .A(n1094), .B(G101), .ZN(n1296) );
XOR2_X1 U1013 ( .A(G110), .B(G140), .Z(n1159) );
NAND2_X1 U1014 ( .A1(n1049), .A2(n1303), .ZN(n1254) );
NAND4_X1 U1015 ( .A1(G953), .A2(G902), .A3(n1242), .A4(n1117), .ZN(n1303) );
INV_X1 U1016 ( .A(G898), .ZN(n1117) );
NAND3_X1 U1017 ( .A1(n1242), .A2(n1039), .A3(G952), .ZN(n1049) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1242) );
NOR2_X1 U1019 ( .A1(n1040), .A2(n1042), .ZN(n1249) );
INV_X1 U1020 ( .A(n1232), .ZN(n1042) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1304), .ZN(n1232) );
XNOR2_X1 U1022 ( .A(n1305), .B(n1173), .ZN(n1040) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1304), .ZN(n1173) );
NAND2_X1 U1024 ( .A1(n1286), .A2(n1268), .ZN(n1304) );
NAND3_X1 U1025 ( .A1(n1306), .A2(n1307), .A3(n1268), .ZN(n1305) );
NAND2_X1 U1026 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XNOR2_X1 U1027 ( .A(n1151), .B(n1310), .ZN(n1309) );
INV_X1 U1028 ( .A(n1169), .ZN(n1308) );
NAND2_X1 U1029 ( .A1(n1169), .A2(n1311), .ZN(n1306) );
NAND2_X1 U1030 ( .A1(n1210), .A2(n1312), .ZN(n1311) );
NAND2_X1 U1031 ( .A1(n1151), .A2(n1212), .ZN(n1312) );
INV_X1 U1032 ( .A(n1150), .ZN(n1151) );
NAND2_X1 U1033 ( .A1(n1310), .A2(n1150), .ZN(n1210) );
NAND2_X1 U1034 ( .A1(n1313), .A2(n1314), .ZN(n1150) );
OR3_X1 U1035 ( .A1(n1233), .A2(n1315), .A3(KEYINPUT14), .ZN(n1314) );
INV_X1 U1036 ( .A(G128), .ZN(n1233) );
NAND2_X1 U1037 ( .A1(n1094), .A2(KEYINPUT14), .ZN(n1313) );
XNOR2_X1 U1038 ( .A(G128), .B(n1315), .ZN(n1094) );
INV_X1 U1039 ( .A(n1212), .ZN(n1310) );
XOR2_X1 U1040 ( .A(G125), .B(n1316), .Z(n1212) );
AND2_X1 U1041 ( .A1(n1039), .A2(G224), .ZN(n1316) );
XOR2_X1 U1042 ( .A(n1123), .B(n1124), .Z(n1169) );
AND2_X1 U1043 ( .A1(n1317), .A2(n1318), .ZN(n1124) );
NAND2_X1 U1044 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
INV_X1 U1045 ( .A(G107), .ZN(n1320) );
XOR2_X1 U1046 ( .A(KEYINPUT53), .B(n1321), .Z(n1319) );
NAND2_X1 U1047 ( .A1(n1321), .A2(G107), .ZN(n1317) );
XNOR2_X1 U1048 ( .A(n1236), .B(G104), .ZN(n1321) );
INV_X1 U1049 ( .A(G101), .ZN(n1236) );
XNOR2_X1 U1050 ( .A(n1322), .B(n1323), .ZN(n1123) );
XOR2_X1 U1051 ( .A(G116), .B(n1324), .Z(n1323) );
XOR2_X1 U1052 ( .A(KEYINPUT39), .B(G119), .Z(n1324) );
XOR2_X1 U1053 ( .A(n1325), .B(n1326), .Z(n1322) );
XNOR2_X1 U1054 ( .A(n1327), .B(n1328), .ZN(n1326) );
NOR2_X1 U1055 ( .A1(KEYINPUT18), .A2(n1329), .ZN(n1328) );
INV_X1 U1056 ( .A(G110), .ZN(n1327) );
NAND2_X1 U1057 ( .A1(KEYINPUT2), .A2(n1280), .ZN(n1325) );
INV_X1 U1058 ( .A(G113), .ZN(n1280) );
AND2_X1 U1059 ( .A1(n1330), .A2(n1252), .ZN(n1044) );
XOR2_X1 U1060 ( .A(n1331), .B(n1083), .Z(n1252) );
NAND2_X1 U1061 ( .A1(n1332), .A2(n1268), .ZN(n1083) );
XOR2_X1 U1062 ( .A(KEYINPUT19), .B(n1133), .Z(n1332) );
XNOR2_X1 U1063 ( .A(n1333), .B(n1334), .ZN(n1133) );
XOR2_X1 U1064 ( .A(n1335), .B(n1336), .Z(n1334) );
NAND2_X1 U1065 ( .A1(n1265), .A2(G217), .ZN(n1336) );
AND2_X1 U1066 ( .A1(G234), .A2(n1039), .ZN(n1265) );
NAND2_X1 U1067 ( .A1(KEYINPUT3), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1068 ( .A(n1338), .B(n1339), .Z(n1337) );
XNOR2_X1 U1069 ( .A(n1222), .B(G134), .ZN(n1339) );
NOR2_X1 U1070 ( .A1(G128), .A2(KEYINPUT17), .ZN(n1338) );
XNOR2_X1 U1071 ( .A(G107), .B(n1340), .ZN(n1333) );
XNOR2_X1 U1072 ( .A(n1329), .B(G116), .ZN(n1340) );
NAND2_X1 U1073 ( .A1(KEYINPUT47), .A2(n1084), .ZN(n1331) );
INV_X1 U1074 ( .A(G478), .ZN(n1084) );
XNOR2_X1 U1075 ( .A(n1078), .B(KEYINPUT51), .ZN(n1330) );
XNOR2_X1 U1076 ( .A(n1341), .B(G475), .ZN(n1078) );
NAND2_X1 U1077 ( .A1(n1268), .A2(n1138), .ZN(n1341) );
NAND2_X1 U1078 ( .A1(n1342), .A2(n1343), .ZN(n1138) );
NAND2_X1 U1079 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1080 ( .A(n1346), .B(KEYINPUT50), .Z(n1342) );
OR2_X1 U1081 ( .A1(n1345), .A2(n1344), .ZN(n1346) );
XOR2_X1 U1082 ( .A(G104), .B(n1347), .Z(n1344) );
XNOR2_X1 U1083 ( .A(n1329), .B(G113), .ZN(n1347) );
INV_X1 U1084 ( .A(G122), .ZN(n1329) );
XNOR2_X1 U1085 ( .A(n1348), .B(n1349), .ZN(n1345) );
XOR2_X1 U1086 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1087 ( .A(G140), .B(n1352), .ZN(n1351) );
AND3_X1 U1088 ( .A1(G214), .A2(n1039), .A3(n1286), .ZN(n1352) );
INV_X1 U1089 ( .A(G237), .ZN(n1286) );
INV_X1 U1090 ( .A(G953), .ZN(n1039) );
NAND2_X1 U1091 ( .A1(KEYINPUT48), .A2(n1353), .ZN(n1350) );
XNOR2_X1 U1092 ( .A(KEYINPUT25), .B(n1354), .ZN(n1353) );
INV_X1 U1093 ( .A(G131), .ZN(n1354) );
XOR2_X1 U1094 ( .A(n1315), .B(n1264), .Z(n1348) );
XOR2_X1 U1095 ( .A(G125), .B(KEYINPUT8), .Z(n1264) );
XOR2_X1 U1096 ( .A(n1222), .B(G146), .Z(n1315) );
INV_X1 U1097 ( .A(G143), .ZN(n1222) );
INV_X1 U1098 ( .A(G902), .ZN(n1268) );
endmodule


