//Key = 1110011111110001100100001111011000001100000001000011100001101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368;

NAND2_X1 U762 ( .A1(n1046), .A2(n1047), .ZN(G9) );
OR2_X1 U763 ( .A1(n1048), .A2(G107), .ZN(n1047) );
XOR2_X1 U764 ( .A(n1049), .B(KEYINPUT35), .Z(n1046) );
NAND2_X1 U765 ( .A1(G107), .A2(n1048), .ZN(n1049) );
NOR2_X1 U766 ( .A1(n1050), .A2(n1051), .ZN(G75) );
NOR2_X1 U767 ( .A1(G952), .A2(n1052), .ZN(n1051) );
NOR3_X1 U768 ( .A1(n1053), .A2(n1054), .A3(n1052), .ZN(n1050) );
NAND2_X1 U769 ( .A1(n1055), .A2(n1056), .ZN(n1052) );
NAND4_X1 U770 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR3_X1 U771 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
XOR2_X1 U772 ( .A(n1064), .B(n1065), .Z(n1063) );
XNOR2_X1 U773 ( .A(G472), .B(n1066), .ZN(n1062) );
XNOR2_X1 U774 ( .A(n1067), .B(n1068), .ZN(n1061) );
NOR2_X1 U775 ( .A1(KEYINPUT39), .A2(n1069), .ZN(n1068) );
INV_X1 U776 ( .A(G475), .ZN(n1069) );
NOR2_X1 U777 ( .A1(n1070), .A2(n1071), .ZN(n1054) );
NOR2_X1 U778 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR3_X1 U779 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NOR2_X1 U780 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U781 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U782 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR2_X1 U783 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR2_X1 U784 ( .A1(n1085), .A2(n1086), .ZN(n1077) );
NOR2_X1 U785 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U786 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR3_X1 U787 ( .A1(n1086), .A2(n1091), .A3(n1092), .ZN(n1072) );
NOR4_X1 U788 ( .A1(n1080), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1092) );
AND3_X1 U789 ( .A1(n1074), .A2(n1096), .A3(KEYINPUT59), .ZN(n1095) );
NOR2_X1 U790 ( .A1(n1097), .A2(n1074), .ZN(n1094) );
NOR2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U792 ( .A1(KEYINPUT59), .A2(n1100), .ZN(n1099) );
NOR2_X1 U793 ( .A1(n1101), .A2(n1076), .ZN(n1093) );
NOR2_X1 U794 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
AND2_X1 U795 ( .A1(n1104), .A2(KEYINPUT10), .ZN(n1103) );
NOR2_X1 U796 ( .A1(n1058), .A2(n1105), .ZN(n1091) );
NOR3_X1 U797 ( .A1(n1106), .A2(KEYINPUT10), .A3(n1076), .ZN(n1105) );
XOR2_X1 U798 ( .A(n1107), .B(n1108), .Z(G72) );
NOR2_X1 U799 ( .A1(n1109), .A2(n1055), .ZN(n1108) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U801 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
NAND2_X1 U802 ( .A1(n1114), .A2(n1055), .ZN(n1113) );
XNOR2_X1 U803 ( .A(n1115), .B(n1116), .ZN(n1114) );
NAND3_X1 U804 ( .A1(G900), .A2(n1116), .A3(G953), .ZN(n1112) );
XOR2_X1 U805 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U806 ( .A(n1119), .B(n1120), .ZN(n1118) );
XNOR2_X1 U807 ( .A(n1121), .B(KEYINPUT41), .ZN(n1120) );
NAND2_X1 U808 ( .A1(KEYINPUT26), .A2(G131), .ZN(n1121) );
XOR2_X1 U809 ( .A(n1122), .B(n1123), .Z(n1117) );
XOR2_X1 U810 ( .A(n1124), .B(n1125), .Z(G69) );
NOR2_X1 U811 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U812 ( .A(n1128), .B(KEYINPUT2), .Z(n1127) );
NAND2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U814 ( .A1(n1129), .A2(n1130), .ZN(n1126) );
NAND3_X1 U815 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1130) );
INV_X1 U816 ( .A(n1134), .ZN(n1133) );
NAND2_X1 U817 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
NAND2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1131) );
XOR2_X1 U819 ( .A(KEYINPUT7), .B(n1135), .Z(n1137) );
XNOR2_X1 U820 ( .A(n1139), .B(n1140), .ZN(n1135) );
XOR2_X1 U821 ( .A(n1141), .B(n1142), .Z(n1139) );
AND2_X1 U822 ( .A1(n1055), .A2(n1143), .ZN(n1129) );
NAND2_X1 U823 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U824 ( .A1(G953), .A2(n1146), .ZN(n1124) );
NAND2_X1 U825 ( .A1(G898), .A2(G224), .ZN(n1146) );
NOR3_X1 U826 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(G66) );
AND3_X1 U827 ( .A1(KEYINPUT28), .A2(G953), .A3(G952), .ZN(n1149) );
NOR2_X1 U828 ( .A1(KEYINPUT28), .A2(n1150), .ZN(n1148) );
INV_X1 U829 ( .A(n1151), .ZN(n1150) );
XNOR2_X1 U830 ( .A(n1152), .B(n1153), .ZN(n1147) );
NOR3_X1 U831 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
XOR2_X1 U832 ( .A(n1157), .B(KEYINPUT55), .Z(n1156) );
NOR2_X1 U833 ( .A1(n1151), .A2(n1158), .ZN(G63) );
XOR2_X1 U834 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U835 ( .A1(G478), .A2(n1161), .ZN(n1160) );
NOR2_X1 U836 ( .A1(KEYINPUT13), .A2(n1162), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1151), .A2(n1163), .ZN(G60) );
XOR2_X1 U838 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U839 ( .A1(n1161), .A2(G475), .ZN(n1164) );
XNOR2_X1 U840 ( .A(G104), .B(n1166), .ZN(G6) );
NAND2_X1 U841 ( .A1(n1104), .A2(n1167), .ZN(n1166) );
NOR2_X1 U842 ( .A1(n1151), .A2(n1168), .ZN(G57) );
XOR2_X1 U843 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U844 ( .A(G101), .B(n1171), .Z(n1170) );
NOR2_X1 U845 ( .A1(KEYINPUT3), .A2(n1172), .ZN(n1171) );
XOR2_X1 U846 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U847 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U848 ( .A(n1177), .B(n1178), .Z(n1173) );
NOR2_X1 U849 ( .A1(KEYINPUT12), .A2(n1179), .ZN(n1178) );
NAND2_X1 U850 ( .A1(n1161), .A2(G472), .ZN(n1177) );
NOR2_X1 U851 ( .A1(n1151), .A2(n1180), .ZN(G54) );
XOR2_X1 U852 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND2_X1 U853 ( .A1(n1161), .A2(G469), .ZN(n1182) );
NAND2_X1 U854 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
NAND2_X1 U855 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XNOR2_X1 U856 ( .A(KEYINPUT21), .B(n1187), .ZN(n1186) );
XOR2_X1 U857 ( .A(n1188), .B(KEYINPUT61), .Z(n1183) );
NAND2_X1 U858 ( .A1(n1189), .A2(n1187), .ZN(n1188) );
NAND2_X1 U859 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND2_X1 U860 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U861 ( .A(KEYINPUT25), .B(n1194), .Z(n1190) );
NOR2_X1 U862 ( .A1(n1192), .A2(n1193), .ZN(n1194) );
XNOR2_X1 U863 ( .A(KEYINPUT11), .B(n1195), .ZN(n1193) );
INV_X1 U864 ( .A(n1185), .ZN(n1189) );
XOR2_X1 U865 ( .A(n1196), .B(n1197), .Z(n1185) );
NAND2_X1 U866 ( .A1(KEYINPUT37), .A2(n1198), .ZN(n1196) );
XOR2_X1 U867 ( .A(KEYINPUT53), .B(n1199), .Z(n1198) );
NOR2_X1 U868 ( .A1(n1151), .A2(n1200), .ZN(G51) );
XOR2_X1 U869 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U870 ( .A(n1203), .B(n1204), .Z(n1202) );
XOR2_X1 U871 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U872 ( .A(n1207), .B(n1208), .Z(n1201) );
XNOR2_X1 U873 ( .A(KEYINPUT52), .B(n1209), .ZN(n1208) );
NAND2_X1 U874 ( .A1(n1161), .A2(n1210), .ZN(n1207) );
NOR2_X1 U875 ( .A1(n1157), .A2(n1155), .ZN(n1161) );
INV_X1 U876 ( .A(n1053), .ZN(n1155) );
NAND3_X1 U877 ( .A1(n1115), .A2(n1144), .A3(n1211), .ZN(n1053) );
XNOR2_X1 U878 ( .A(n1145), .B(KEYINPUT16), .ZN(n1211) );
AND4_X1 U879 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1145) );
OR2_X1 U880 ( .A1(n1216), .A2(n1217), .ZN(n1212) );
AND4_X1 U881 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1048), .ZN(n1144) );
NAND2_X1 U882 ( .A1(n1102), .A2(n1167), .ZN(n1048) );
AND2_X1 U883 ( .A1(n1221), .A2(n1222), .ZN(n1167) );
NAND4_X1 U884 ( .A1(n1223), .A2(n1104), .A3(n1224), .A4(n1222), .ZN(n1218) );
AND2_X1 U885 ( .A1(n1225), .A2(n1088), .ZN(n1224) );
XOR2_X1 U886 ( .A(n1226), .B(KEYINPUT18), .Z(n1223) );
AND4_X1 U887 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1115) );
NOR4_X1 U888 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1230) );
NOR3_X1 U889 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1229) );
NOR2_X1 U890 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
AND4_X1 U891 ( .A1(n1238), .A2(n1240), .A3(n1102), .A4(n1241), .ZN(n1236) );
AND2_X1 U892 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
INV_X1 U893 ( .A(KEYINPUT29), .ZN(n1238) );
NOR2_X1 U894 ( .A1(n1244), .A2(n1245), .ZN(n1235) );
XOR2_X1 U895 ( .A(n1246), .B(KEYINPUT43), .Z(n1244) );
NOR2_X1 U896 ( .A1(n1055), .A2(G952), .ZN(n1151) );
XNOR2_X1 U897 ( .A(n1233), .B(n1247), .ZN(G48) );
NOR2_X1 U898 ( .A1(G146), .A2(KEYINPUT63), .ZN(n1247) );
AND3_X1 U899 ( .A1(n1248), .A2(n1104), .A3(n1241), .ZN(n1233) );
XOR2_X1 U900 ( .A(n1249), .B(n1250), .Z(G45) );
XOR2_X1 U901 ( .A(KEYINPUT22), .B(G143), .Z(n1250) );
NOR2_X1 U902 ( .A1(n1245), .A2(n1246), .ZN(n1249) );
NAND4_X1 U903 ( .A1(n1096), .A2(n1248), .A3(n1251), .A4(n1252), .ZN(n1246) );
XOR2_X1 U904 ( .A(n1227), .B(n1253), .Z(G42) );
NAND2_X1 U905 ( .A1(KEYINPUT50), .A2(G140), .ZN(n1253) );
NAND3_X1 U906 ( .A1(n1098), .A2(n1104), .A3(n1254), .ZN(n1227) );
XNOR2_X1 U907 ( .A(n1255), .B(n1228), .ZN(G39) );
NAND2_X1 U908 ( .A1(n1256), .A2(n1254), .ZN(n1228) );
XNOR2_X1 U909 ( .A(G137), .B(KEYINPUT57), .ZN(n1255) );
XOR2_X1 U910 ( .A(G134), .B(n1232), .Z(G36) );
AND3_X1 U911 ( .A1(n1254), .A2(n1102), .A3(n1096), .ZN(n1232) );
XOR2_X1 U912 ( .A(n1257), .B(G131), .Z(G33) );
NAND2_X1 U913 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U914 ( .A1(n1234), .A2(n1260), .ZN(n1259) );
INV_X1 U915 ( .A(KEYINPUT17), .ZN(n1260) );
AND2_X1 U916 ( .A1(n1261), .A2(n1254), .ZN(n1234) );
AND2_X1 U917 ( .A1(n1059), .A2(n1248), .ZN(n1254) );
INV_X1 U918 ( .A(n1086), .ZN(n1059) );
NAND4_X1 U919 ( .A1(n1248), .A2(n1086), .A3(n1261), .A4(KEYINPUT17), .ZN(n1258) );
NAND2_X1 U920 ( .A1(n1262), .A2(n1084), .ZN(n1086) );
XOR2_X1 U921 ( .A(n1263), .B(n1239), .Z(G30) );
NAND3_X1 U922 ( .A1(n1248), .A2(n1102), .A3(n1241), .ZN(n1239) );
NOR3_X1 U923 ( .A1(n1245), .A2(n1057), .A3(n1264), .ZN(n1241) );
AND2_X1 U924 ( .A1(n1088), .A2(n1243), .ZN(n1248) );
XOR2_X1 U925 ( .A(n1265), .B(n1219), .Z(G3) );
NAND3_X1 U926 ( .A1(n1096), .A2(n1221), .A3(n1266), .ZN(n1219) );
XOR2_X1 U927 ( .A(n1267), .B(G125), .Z(G27) );
NAND2_X1 U928 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U929 ( .A1(n1231), .A2(n1270), .ZN(n1269) );
INV_X1 U930 ( .A(KEYINPUT49), .ZN(n1270) );
AND3_X1 U931 ( .A1(n1058), .A2(n1271), .A3(n1098), .ZN(n1231) );
NAND4_X1 U932 ( .A1(n1271), .A2(n1080), .A3(n1098), .A4(KEYINPUT49), .ZN(n1268) );
AND3_X1 U933 ( .A1(n1082), .A2(n1243), .A3(n1104), .ZN(n1271) );
NAND2_X1 U934 ( .A1(n1272), .A2(n1071), .ZN(n1243) );
NAND4_X1 U935 ( .A1(G902), .A2(G953), .A3(n1273), .A4(n1111), .ZN(n1272) );
INV_X1 U936 ( .A(G900), .ZN(n1111) );
XOR2_X1 U937 ( .A(G122), .B(n1274), .Z(G24) );
NOR3_X1 U938 ( .A1(n1216), .A2(KEYINPUT48), .A3(n1217), .ZN(n1274) );
NAND3_X1 U939 ( .A1(n1251), .A2(n1252), .A3(n1222), .ZN(n1216) );
INV_X1 U940 ( .A(n1076), .ZN(n1222) );
NAND2_X1 U941 ( .A1(n1057), .A2(n1264), .ZN(n1076) );
NAND2_X1 U942 ( .A1(n1275), .A2(n1276), .ZN(G21) );
NAND2_X1 U943 ( .A1(G119), .A2(n1213), .ZN(n1276) );
XOR2_X1 U944 ( .A(KEYINPUT36), .B(n1277), .Z(n1275) );
NOR2_X1 U945 ( .A1(G119), .A2(n1213), .ZN(n1277) );
NAND2_X1 U946 ( .A1(n1278), .A2(n1256), .ZN(n1213) );
NOR3_X1 U947 ( .A1(n1264), .A2(n1057), .A3(n1074), .ZN(n1256) );
INV_X1 U948 ( .A(n1266), .ZN(n1074) );
INV_X1 U949 ( .A(n1279), .ZN(n1264) );
XOR2_X1 U950 ( .A(n1214), .B(n1280), .Z(G18) );
NAND2_X1 U951 ( .A1(KEYINPUT27), .A2(G116), .ZN(n1280) );
NAND3_X1 U952 ( .A1(n1096), .A2(n1102), .A3(n1278), .ZN(n1214) );
INV_X1 U953 ( .A(n1217), .ZN(n1278) );
NAND3_X1 U954 ( .A1(n1082), .A2(n1225), .A3(n1058), .ZN(n1217) );
INV_X1 U955 ( .A(n1245), .ZN(n1082) );
AND2_X1 U956 ( .A1(n1281), .A2(n1252), .ZN(n1102) );
INV_X1 U957 ( .A(n1100), .ZN(n1096) );
XOR2_X1 U958 ( .A(n1215), .B(n1282), .Z(G15) );
NAND2_X1 U959 ( .A1(KEYINPUT30), .A2(G113), .ZN(n1282) );
NAND4_X1 U960 ( .A1(n1261), .A2(n1058), .A3(n1226), .A4(n1225), .ZN(n1215) );
INV_X1 U961 ( .A(n1080), .ZN(n1058) );
NAND2_X1 U962 ( .A1(n1283), .A2(n1090), .ZN(n1080) );
NOR2_X1 U963 ( .A1(n1100), .A2(n1106), .ZN(n1261) );
INV_X1 U964 ( .A(n1104), .ZN(n1106) );
NOR2_X1 U965 ( .A1(n1252), .A2(n1281), .ZN(n1104) );
NAND2_X1 U966 ( .A1(n1279), .A2(n1057), .ZN(n1100) );
XOR2_X1 U967 ( .A(n1284), .B(n1220), .Z(G12) );
NAND3_X1 U968 ( .A1(n1098), .A2(n1221), .A3(n1266), .ZN(n1220) );
NOR2_X1 U969 ( .A1(n1252), .A2(n1251), .ZN(n1266) );
INV_X1 U970 ( .A(n1281), .ZN(n1251) );
XOR2_X1 U971 ( .A(n1067), .B(G475), .Z(n1281) );
NAND2_X1 U972 ( .A1(n1165), .A2(n1157), .ZN(n1067) );
XNOR2_X1 U973 ( .A(n1285), .B(n1286), .ZN(n1165) );
XOR2_X1 U974 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U975 ( .A(G131), .B(G104), .Z(n1288) );
AND3_X1 U976 ( .A1(G214), .A2(n1055), .A3(n1289), .ZN(n1287) );
XOR2_X1 U977 ( .A(n1290), .B(n1140), .Z(n1285) );
XNOR2_X1 U978 ( .A(n1291), .B(n1123), .ZN(n1290) );
NAND3_X1 U979 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1252) );
OR2_X1 U980 ( .A1(n1295), .A2(n1065), .ZN(n1294) );
NAND3_X1 U981 ( .A1(n1065), .A2(n1295), .A3(G478), .ZN(n1293) );
NAND2_X1 U982 ( .A1(n1296), .A2(n1064), .ZN(n1292) );
INV_X1 U983 ( .A(G478), .ZN(n1064) );
NAND2_X1 U984 ( .A1(n1297), .A2(n1295), .ZN(n1296) );
INV_X1 U985 ( .A(KEYINPUT44), .ZN(n1295) );
XOR2_X1 U986 ( .A(n1065), .B(KEYINPUT40), .Z(n1297) );
NAND2_X1 U987 ( .A1(n1162), .A2(n1157), .ZN(n1065) );
XOR2_X1 U988 ( .A(n1298), .B(n1299), .Z(n1162) );
XOR2_X1 U989 ( .A(G134), .B(n1300), .Z(n1299) );
XOR2_X1 U990 ( .A(KEYINPUT4), .B(G143), .Z(n1300) );
XOR2_X1 U991 ( .A(n1301), .B(n1302), .Z(n1298) );
XOR2_X1 U992 ( .A(G128), .B(n1303), .Z(n1302) );
AND2_X1 U993 ( .A1(n1304), .A2(G217), .ZN(n1303) );
NAND3_X1 U994 ( .A1(n1305), .A2(n1306), .A3(KEYINPUT19), .ZN(n1301) );
NAND3_X1 U995 ( .A1(G107), .A2(n1307), .A3(n1308), .ZN(n1306) );
INV_X1 U996 ( .A(KEYINPUT58), .ZN(n1308) );
NAND2_X1 U997 ( .A1(n1309), .A2(KEYINPUT58), .ZN(n1305) );
XOR2_X1 U998 ( .A(G107), .B(n1307), .Z(n1309) );
XOR2_X1 U999 ( .A(G116), .B(G122), .Z(n1307) );
AND3_X1 U1000 ( .A1(n1226), .A2(n1225), .A3(n1088), .ZN(n1221) );
INV_X1 U1001 ( .A(n1242), .ZN(n1088) );
NAND2_X1 U1002 ( .A1(n1089), .A2(n1090), .ZN(n1242) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1310), .ZN(n1090) );
INV_X1 U1004 ( .A(n1283), .ZN(n1089) );
XOR2_X1 U1005 ( .A(n1311), .B(G469), .Z(n1283) );
NAND2_X1 U1006 ( .A1(n1312), .A2(n1157), .ZN(n1311) );
XOR2_X1 U1007 ( .A(n1313), .B(n1314), .Z(n1312) );
XOR2_X1 U1008 ( .A(n1197), .B(n1192), .Z(n1314) );
INV_X1 U1009 ( .A(n1179), .ZN(n1192) );
NOR2_X1 U1010 ( .A1(n1110), .A2(G953), .ZN(n1197) );
INV_X1 U1011 ( .A(G227), .ZN(n1110) );
XOR2_X1 U1012 ( .A(n1195), .B(n1199), .Z(n1313) );
XNOR2_X1 U1013 ( .A(G140), .B(n1284), .ZN(n1199) );
XOR2_X1 U1014 ( .A(n1315), .B(n1316), .Z(n1195) );
INV_X1 U1015 ( .A(n1122), .ZN(n1316) );
XOR2_X1 U1016 ( .A(n1317), .B(n1318), .Z(n1122) );
XOR2_X1 U1017 ( .A(n1319), .B(n1320), .Z(n1318) );
NOR2_X1 U1018 ( .A1(KEYINPUT62), .A2(n1263), .ZN(n1320) );
NOR2_X1 U1019 ( .A1(G143), .A2(KEYINPUT20), .ZN(n1319) );
XOR2_X1 U1020 ( .A(n1321), .B(G146), .Z(n1317) );
XNOR2_X1 U1021 ( .A(KEYINPUT9), .B(KEYINPUT46), .ZN(n1321) );
XOR2_X1 U1022 ( .A(n1136), .B(KEYINPUT8), .Z(n1315) );
NAND2_X1 U1023 ( .A1(n1071), .A2(n1322), .ZN(n1225) );
NAND3_X1 U1024 ( .A1(n1134), .A2(n1273), .A3(G902), .ZN(n1322) );
NOR2_X1 U1025 ( .A1(n1055), .A2(G898), .ZN(n1134) );
NAND3_X1 U1026 ( .A1(n1273), .A2(n1055), .A3(n1323), .ZN(n1071) );
XNOR2_X1 U1027 ( .A(G952), .B(KEYINPUT6), .ZN(n1323) );
NAND2_X1 U1028 ( .A1(G237), .A2(G234), .ZN(n1273) );
XOR2_X1 U1029 ( .A(n1245), .B(KEYINPUT15), .Z(n1226) );
NAND2_X1 U1030 ( .A1(n1083), .A2(n1084), .ZN(n1245) );
NAND2_X1 U1031 ( .A1(G214), .A2(n1324), .ZN(n1084) );
INV_X1 U1032 ( .A(n1262), .ZN(n1083) );
XOR2_X1 U1033 ( .A(n1325), .B(n1210), .Z(n1262) );
AND2_X1 U1034 ( .A1(G210), .A2(n1324), .ZN(n1210) );
NAND2_X1 U1035 ( .A1(n1289), .A2(n1157), .ZN(n1324) );
NAND2_X1 U1036 ( .A1(n1326), .A2(n1157), .ZN(n1325) );
XOR2_X1 U1037 ( .A(n1327), .B(n1328), .Z(n1326) );
INV_X1 U1038 ( .A(n1203), .ZN(n1328) );
XOR2_X1 U1039 ( .A(n1329), .B(n1330), .Z(n1203) );
XOR2_X1 U1040 ( .A(n1142), .B(n1140), .Z(n1330) );
XOR2_X1 U1041 ( .A(G122), .B(G113), .Z(n1140) );
XNOR2_X1 U1042 ( .A(n1331), .B(KEYINPUT0), .ZN(n1142) );
XOR2_X1 U1043 ( .A(n1138), .B(n1141), .Z(n1329) );
NAND2_X1 U1044 ( .A1(KEYINPUT5), .A2(n1284), .ZN(n1141) );
INV_X1 U1045 ( .A(n1136), .ZN(n1138) );
XOR2_X1 U1046 ( .A(n1265), .B(n1332), .Z(n1136) );
XOR2_X1 U1047 ( .A(G107), .B(G104), .Z(n1332) );
NAND3_X1 U1048 ( .A1(n1333), .A2(n1334), .A3(KEYINPUT24), .ZN(n1327) );
NAND2_X1 U1049 ( .A1(n1335), .A2(n1209), .ZN(n1334) );
XOR2_X1 U1050 ( .A(KEYINPUT60), .B(n1336), .Z(n1333) );
NOR2_X1 U1051 ( .A1(n1335), .A2(n1209), .ZN(n1336) );
NAND2_X1 U1052 ( .A1(G224), .A2(n1055), .ZN(n1209) );
XOR2_X1 U1053 ( .A(n1337), .B(n1338), .Z(n1335) );
NOR2_X1 U1054 ( .A1(KEYINPUT32), .A2(n1205), .ZN(n1338) );
INV_X1 U1055 ( .A(n1175), .ZN(n1205) );
NOR2_X1 U1056 ( .A1(n1279), .A2(n1057), .ZN(n1098) );
XNOR2_X1 U1057 ( .A(n1339), .B(n1154), .ZN(n1057) );
NAND2_X1 U1058 ( .A1(G217), .A2(n1310), .ZN(n1154) );
NAND2_X1 U1059 ( .A1(G234), .A2(n1157), .ZN(n1310) );
NAND2_X1 U1060 ( .A1(n1152), .A2(n1157), .ZN(n1339) );
XNOR2_X1 U1061 ( .A(n1340), .B(n1341), .ZN(n1152) );
XNOR2_X1 U1062 ( .A(G137), .B(n1342), .ZN(n1341) );
NAND2_X1 U1063 ( .A1(n1343), .A2(KEYINPUT1), .ZN(n1342) );
XOR2_X1 U1064 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1065 ( .A(n1346), .B(n1347), .ZN(n1345) );
NOR2_X1 U1066 ( .A1(G110), .A2(KEYINPUT56), .ZN(n1347) );
NAND4_X1 U1067 ( .A1(KEYINPUT51), .A2(n1348), .A3(n1349), .A4(n1350), .ZN(n1346) );
NAND3_X1 U1068 ( .A1(n1123), .A2(n1351), .A3(G146), .ZN(n1350) );
NAND2_X1 U1069 ( .A1(n1352), .A2(n1353), .ZN(n1349) );
INV_X1 U1070 ( .A(G146), .ZN(n1353) );
NAND2_X1 U1071 ( .A1(n1354), .A2(n1351), .ZN(n1352) );
XOR2_X1 U1072 ( .A(KEYINPUT33), .B(n1123), .Z(n1354) );
OR2_X1 U1073 ( .A1(n1351), .A2(n1123), .ZN(n1348) );
XOR2_X1 U1074 ( .A(G140), .B(n1206), .Z(n1123) );
INV_X1 U1075 ( .A(n1337), .ZN(n1206) );
XNOR2_X1 U1076 ( .A(G125), .B(KEYINPUT34), .ZN(n1337) );
INV_X1 U1077 ( .A(KEYINPUT54), .ZN(n1351) );
XNOR2_X1 U1078 ( .A(G119), .B(n1355), .ZN(n1344) );
XOR2_X1 U1079 ( .A(KEYINPUT42), .B(G128), .Z(n1355) );
NAND2_X1 U1080 ( .A1(G221), .A2(n1304), .ZN(n1340) );
AND2_X1 U1081 ( .A1(n1356), .A2(n1055), .ZN(n1304) );
XOR2_X1 U1082 ( .A(KEYINPUT14), .B(G234), .Z(n1356) );
XOR2_X1 U1083 ( .A(n1066), .B(n1357), .Z(n1279) );
NOR2_X1 U1084 ( .A1(G472), .A2(KEYINPUT23), .ZN(n1357) );
NAND2_X1 U1085 ( .A1(n1358), .A2(n1157), .ZN(n1066) );
INV_X1 U1086 ( .A(G902), .ZN(n1157) );
XOR2_X1 U1087 ( .A(n1359), .B(n1360), .Z(n1358) );
XOR2_X1 U1088 ( .A(n1169), .B(n1176), .Z(n1360) );
XOR2_X1 U1089 ( .A(G113), .B(n1361), .Z(n1176) );
NOR2_X1 U1090 ( .A1(KEYINPUT47), .A2(n1331), .ZN(n1361) );
XNOR2_X1 U1091 ( .A(G116), .B(G119), .ZN(n1331) );
AND3_X1 U1092 ( .A1(n1289), .A2(n1055), .A3(G210), .ZN(n1169) );
INV_X1 U1093 ( .A(G953), .ZN(n1055) );
INV_X1 U1094 ( .A(G237), .ZN(n1289) );
XNOR2_X1 U1095 ( .A(n1362), .B(n1363), .ZN(n1359) );
NOR2_X1 U1096 ( .A1(KEYINPUT31), .A2(n1265), .ZN(n1363) );
INV_X1 U1097 ( .A(G101), .ZN(n1265) );
NOR2_X1 U1098 ( .A1(KEYINPUT38), .A2(n1364), .ZN(n1362) );
XOR2_X1 U1099 ( .A(n1179), .B(n1175), .Z(n1364) );
XOR2_X1 U1100 ( .A(n1263), .B(n1291), .Z(n1175) );
XOR2_X1 U1101 ( .A(G143), .B(G146), .Z(n1291) );
INV_X1 U1102 ( .A(G128), .ZN(n1263) );
NAND2_X1 U1103 ( .A1(n1365), .A2(n1366), .ZN(n1179) );
NAND2_X1 U1104 ( .A1(n1119), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1105 ( .A(KEYINPUT45), .B(n1368), .Z(n1365) );
NOR2_X1 U1106 ( .A1(n1119), .A2(n1367), .ZN(n1368) );
INV_X1 U1107 ( .A(G131), .ZN(n1367) );
XNOR2_X1 U1108 ( .A(G134), .B(G137), .ZN(n1119) );
INV_X1 U1109 ( .A(G110), .ZN(n1284) );
endmodule


