//Key = 1000110110100110100010100010110110001000111010101000011100100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332;

XOR2_X1 U729 ( .A(n1010), .B(n1011), .Z(G9) );
NAND3_X1 U730 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(G75) );
NAND2_X1 U731 ( .A1(G952), .A2(n1015), .ZN(n1014) );
NAND3_X1 U732 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NAND4_X1 U733 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1017) );
NAND2_X1 U734 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND3_X1 U735 ( .A1(n1025), .A2(n1026), .A3(KEYINPUT21), .ZN(n1024) );
NAND3_X1 U736 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1021) );
NAND2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
OR2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U739 ( .A1(n1025), .A2(n1034), .ZN(n1027) );
NAND2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U741 ( .A1(n1026), .A2(n1037), .ZN(n1036) );
INV_X1 U742 ( .A(KEYINPUT21), .ZN(n1037) );
NAND4_X1 U743 ( .A1(n1025), .A2(n1030), .A3(n1029), .A4(n1038), .ZN(n1016) );
NAND2_X1 U744 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U745 ( .A1(n1020), .A2(n1041), .ZN(n1040) );
NAND2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U747 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
INV_X1 U748 ( .A(KEYINPUT47), .ZN(n1045) );
NAND2_X1 U749 ( .A1(n1019), .A2(n1047), .ZN(n1039) );
NAND3_X1 U750 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NAND2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
XOR2_X1 U752 ( .A(n1053), .B(KEYINPUT30), .Z(n1051) );
NAND2_X1 U753 ( .A1(KEYINPUT47), .A2(n1020), .ZN(n1048) );
INV_X1 U754 ( .A(n1023), .ZN(n1029) );
XOR2_X1 U755 ( .A(n1054), .B(KEYINPUT54), .Z(n1023) );
NAND4_X1 U756 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1012) );
NOR4_X1 U757 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
XOR2_X1 U758 ( .A(KEYINPUT27), .B(n1046), .Z(n1062) );
XOR2_X1 U759 ( .A(KEYINPUT35), .B(n1063), .Z(n1061) );
XOR2_X1 U760 ( .A(n1064), .B(n1065), .Z(n1060) );
NOR2_X1 U761 ( .A1(KEYINPUT62), .A2(n1066), .ZN(n1065) );
NOR3_X1 U762 ( .A1(n1067), .A2(n1068), .A3(n1052), .ZN(n1057) );
INV_X1 U763 ( .A(n1069), .ZN(n1068) );
NOR2_X1 U764 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
XOR2_X1 U765 ( .A(KEYINPUT44), .B(G478), .Z(n1071) );
XOR2_X1 U766 ( .A(n1072), .B(n1073), .Z(n1056) );
NOR2_X1 U767 ( .A1(G475), .A2(KEYINPUT23), .ZN(n1073) );
XOR2_X1 U768 ( .A(n1074), .B(n1075), .Z(G72) );
NOR2_X1 U769 ( .A1(n1076), .A2(n1013), .ZN(n1075) );
XOR2_X1 U770 ( .A(n1077), .B(KEYINPUT14), .Z(n1076) );
NAND2_X1 U771 ( .A1(G900), .A2(G227), .ZN(n1077) );
NAND3_X1 U772 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1074) );
OR2_X1 U773 ( .A1(n1081), .A2(KEYINPUT58), .ZN(n1080) );
NAND3_X1 U774 ( .A1(KEYINPUT58), .A2(n1081), .A3(n1082), .ZN(n1079) );
AND2_X1 U775 ( .A1(n1013), .A2(n1083), .ZN(n1081) );
OR3_X1 U776 ( .A1(n1083), .A2(n1084), .A3(n1082), .ZN(n1078) );
XNOR2_X1 U777 ( .A(n1085), .B(n1086), .ZN(n1082) );
NOR2_X1 U778 ( .A1(KEYINPUT3), .A2(n1087), .ZN(n1086) );
XOR2_X1 U779 ( .A(n1088), .B(n1089), .Z(n1087) );
XOR2_X1 U780 ( .A(n1090), .B(n1091), .Z(n1089) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(n1088) );
NOR2_X1 U782 ( .A1(G134), .A2(KEYINPUT2), .ZN(n1093) );
NAND3_X1 U783 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1085) );
OR2_X1 U784 ( .A1(n1097), .A2(KEYINPUT13), .ZN(n1096) );
NAND3_X1 U785 ( .A1(KEYINPUT13), .A2(n1097), .A3(G125), .ZN(n1095) );
NAND2_X1 U786 ( .A1(n1098), .A2(n1099), .ZN(n1094) );
NAND2_X1 U787 ( .A1(KEYINPUT13), .A2(n1100), .ZN(n1098) );
XOR2_X1 U788 ( .A(KEYINPUT55), .B(G140), .Z(n1100) );
NOR2_X1 U789 ( .A1(n1013), .A2(G900), .ZN(n1084) );
NAND2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(G69) );
NAND2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U792 ( .A1(G953), .A2(n1105), .ZN(n1103) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1105) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
OR2_X1 U796 ( .A1(n1013), .A2(G224), .ZN(n1109) );
INV_X1 U797 ( .A(n1104), .ZN(n1106) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1104) );
NAND3_X1 U799 ( .A1(n1112), .A2(n1013), .A3(n1113), .ZN(n1111) );
XNOR2_X1 U800 ( .A(n1114), .B(n1115), .ZN(n1113) );
XOR2_X1 U801 ( .A(KEYINPUT60), .B(KEYINPUT11), .Z(n1115) );
XOR2_X1 U802 ( .A(n1116), .B(KEYINPUT61), .Z(n1110) );
NAND2_X1 U803 ( .A1(n1114), .A2(n1117), .ZN(n1116) );
XNOR2_X1 U804 ( .A(KEYINPUT6), .B(n1112), .ZN(n1117) );
AND2_X1 U805 ( .A1(n1118), .A2(n1108), .ZN(n1114) );
INV_X1 U806 ( .A(n1119), .ZN(n1108) );
XOR2_X1 U807 ( .A(n1120), .B(n1121), .Z(n1118) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND2_X1 U809 ( .A1(KEYINPUT31), .A2(n1124), .ZN(n1122) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XOR2_X1 U811 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U812 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n1125), .A2(n1131), .ZN(G63) );
XOR2_X1 U814 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U815 ( .A(n1134), .B(KEYINPUT63), .Z(n1133) );
NAND2_X1 U816 ( .A1(n1129), .A2(G478), .ZN(n1134) );
NOR2_X1 U817 ( .A1(n1125), .A2(n1135), .ZN(G60) );
XOR2_X1 U818 ( .A(n1136), .B(n1137), .Z(n1135) );
XNOR2_X1 U819 ( .A(n1138), .B(KEYINPUT9), .ZN(n1137) );
NAND3_X1 U820 ( .A1(n1129), .A2(G475), .A3(KEYINPUT36), .ZN(n1138) );
NAND2_X1 U821 ( .A1(n1139), .A2(n1140), .ZN(G6) );
NAND2_X1 U822 ( .A1(G104), .A2(n1141), .ZN(n1140) );
XOR2_X1 U823 ( .A(n1142), .B(KEYINPUT25), .Z(n1139) );
OR2_X1 U824 ( .A1(n1141), .A2(G104), .ZN(n1142) );
NAND2_X1 U825 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
XOR2_X1 U826 ( .A(n1145), .B(KEYINPUT53), .Z(n1143) );
NOR2_X1 U827 ( .A1(n1125), .A2(n1146), .ZN(G57) );
NOR3_X1 U828 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
NOR2_X1 U829 ( .A1(G101), .A2(n1150), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR3_X1 U831 ( .A1(n1153), .A2(n1154), .A3(n1152), .ZN(n1148) );
INV_X1 U832 ( .A(n1151), .ZN(n1154) );
AND2_X1 U833 ( .A1(n1152), .A2(n1155), .ZN(n1147) );
NOR2_X1 U834 ( .A1(KEYINPUT24), .A2(n1156), .ZN(n1152) );
XOR2_X1 U835 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U836 ( .A1(n1129), .A2(G472), .ZN(n1157) );
NOR2_X1 U837 ( .A1(n1125), .A2(n1159), .ZN(G54) );
XOR2_X1 U838 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U839 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U840 ( .A(n1164), .B(n1165), .Z(n1160) );
XNOR2_X1 U841 ( .A(n1166), .B(n1167), .ZN(n1165) );
NAND3_X1 U842 ( .A1(G902), .A2(G469), .A3(n1168), .ZN(n1167) );
XNOR2_X1 U843 ( .A(n1018), .B(KEYINPUT50), .ZN(n1168) );
NOR2_X1 U844 ( .A1(n1125), .A2(n1169), .ZN(G51) );
XOR2_X1 U845 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND3_X1 U846 ( .A1(n1129), .A2(n1064), .A3(KEYINPUT28), .ZN(n1171) );
NOR2_X1 U847 ( .A1(n1172), .A2(n1018), .ZN(n1129) );
NOR2_X1 U848 ( .A1(n1112), .A2(n1083), .ZN(n1018) );
NAND4_X1 U849 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1083) );
AND4_X1 U850 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NAND2_X1 U851 ( .A1(n1181), .A2(n1182), .ZN(n1175) );
NAND2_X1 U852 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND2_X1 U853 ( .A1(n1185), .A2(n1033), .ZN(n1184) );
NAND2_X1 U854 ( .A1(n1186), .A2(n1187), .ZN(n1183) );
NAND3_X1 U855 ( .A1(n1185), .A2(n1025), .A3(n1188), .ZN(n1173) );
XNOR2_X1 U856 ( .A(n1189), .B(KEYINPUT32), .ZN(n1188) );
NAND4_X1 U857 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1112) );
AND3_X1 U858 ( .A1(n1194), .A2(n1011), .A3(n1195), .ZN(n1193) );
NAND3_X1 U859 ( .A1(n1033), .A2(n1196), .A3(n1030), .ZN(n1011) );
NAND2_X1 U860 ( .A1(n1144), .A2(n1197), .ZN(n1192) );
NAND3_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1145), .ZN(n1197) );
NAND4_X1 U862 ( .A1(n1032), .A2(n1030), .A3(n1200), .A4(n1201), .ZN(n1145) );
NAND3_X1 U863 ( .A1(n1202), .A2(n1030), .A3(n1187), .ZN(n1190) );
NAND3_X1 U864 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1170) );
OR2_X1 U865 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U866 ( .A1(n1208), .A2(n1209), .ZN(n1204) );
INV_X1 U867 ( .A(KEYINPUT7), .ZN(n1209) );
NAND2_X1 U868 ( .A1(n1210), .A2(n1206), .ZN(n1208) );
XOR2_X1 U869 ( .A(n1211), .B(KEYINPUT42), .Z(n1210) );
NAND2_X1 U870 ( .A1(KEYINPUT7), .A2(n1212), .ZN(n1203) );
NAND2_X1 U871 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
OR2_X1 U872 ( .A1(n1207), .A2(KEYINPUT42), .ZN(n1214) );
NAND3_X1 U873 ( .A1(n1207), .A2(n1206), .A3(KEYINPUT42), .ZN(n1213) );
AND2_X1 U874 ( .A1(n1215), .A2(n1216), .ZN(n1125) );
XOR2_X1 U875 ( .A(KEYINPUT45), .B(G953), .Z(n1215) );
XNOR2_X1 U876 ( .A(G146), .B(n1174), .ZN(G48) );
NAND4_X1 U877 ( .A1(n1186), .A2(n1032), .A3(n1189), .A4(n1144), .ZN(n1174) );
XNOR2_X1 U878 ( .A(G143), .B(n1217), .ZN(G45) );
NAND3_X1 U879 ( .A1(n1186), .A2(n1187), .A3(n1218), .ZN(n1217) );
XOR2_X1 U880 ( .A(n1035), .B(KEYINPUT29), .Z(n1218) );
XOR2_X1 U881 ( .A(n1097), .B(n1180), .Z(G42) );
NAND3_X1 U882 ( .A1(n1032), .A2(n1026), .A3(n1185), .ZN(n1180) );
XOR2_X1 U883 ( .A(G137), .B(n1219), .Z(G39) );
NOR2_X1 U884 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XNOR2_X1 U885 ( .A(G134), .B(n1222), .ZN(G36) );
NAND4_X1 U886 ( .A1(n1186), .A2(n1181), .A3(n1033), .A4(n1223), .ZN(n1222) );
XOR2_X1 U887 ( .A(KEYINPUT43), .B(n1019), .Z(n1223) );
XOR2_X1 U888 ( .A(n1092), .B(n1179), .Z(G33) );
NAND3_X1 U889 ( .A1(n1032), .A2(n1181), .A3(n1185), .ZN(n1179) );
INV_X1 U890 ( .A(n1221), .ZN(n1185) );
NAND2_X1 U891 ( .A1(n1186), .A2(n1019), .ZN(n1221) );
AND2_X1 U892 ( .A1(n1044), .A2(n1224), .ZN(n1019) );
NOR2_X1 U893 ( .A1(n1225), .A2(n1050), .ZN(n1186) );
XNOR2_X1 U894 ( .A(n1200), .B(KEYINPUT17), .ZN(n1050) );
XNOR2_X1 U895 ( .A(G128), .B(n1178), .ZN(G30) );
NAND3_X1 U896 ( .A1(n1226), .A2(n1189), .A3(n1227), .ZN(n1178) );
AND3_X1 U897 ( .A1(n1033), .A2(n1200), .A3(n1144), .ZN(n1227) );
INV_X1 U898 ( .A(n1225), .ZN(n1226) );
NAND2_X1 U899 ( .A1(n1228), .A2(n1229), .ZN(G3) );
OR2_X1 U900 ( .A1(n1191), .A2(G101), .ZN(n1229) );
XOR2_X1 U901 ( .A(n1230), .B(KEYINPUT57), .Z(n1228) );
NAND2_X1 U902 ( .A1(G101), .A2(n1191), .ZN(n1230) );
NAND3_X1 U903 ( .A1(n1025), .A2(n1196), .A3(n1181), .ZN(n1191) );
XOR2_X1 U904 ( .A(n1099), .B(n1177), .Z(G27) );
NAND4_X1 U905 ( .A1(n1026), .A2(n1020), .A3(n1144), .A4(n1231), .ZN(n1177) );
NOR2_X1 U906 ( .A1(n1232), .A2(n1225), .ZN(n1231) );
NAND3_X1 U907 ( .A1(n1233), .A2(n1234), .A3(n1054), .ZN(n1225) );
NAND2_X1 U908 ( .A1(n1216), .A2(n1013), .ZN(n1234) );
INV_X1 U909 ( .A(G952), .ZN(n1216) );
NAND2_X1 U910 ( .A1(G953), .A2(n1235), .ZN(n1233) );
OR2_X1 U911 ( .A1(n1172), .A2(G900), .ZN(n1235) );
INV_X1 U912 ( .A(G125), .ZN(n1099) );
XNOR2_X1 U913 ( .A(G122), .B(n1236), .ZN(G24) );
NAND3_X1 U914 ( .A1(n1187), .A2(n1202), .A3(n1237), .ZN(n1236) );
XNOR2_X1 U915 ( .A(n1030), .B(KEYINPUT26), .ZN(n1237) );
NOR2_X1 U916 ( .A1(n1238), .A2(n1239), .ZN(n1030) );
INV_X1 U917 ( .A(n1055), .ZN(n1239) );
AND3_X1 U918 ( .A1(n1240), .A2(n1241), .A3(n1144), .ZN(n1187) );
OR2_X1 U919 ( .A1(n1033), .A2(KEYINPUT22), .ZN(n1241) );
NAND2_X1 U920 ( .A1(KEYINPUT22), .A2(n1242), .ZN(n1240) );
NAND2_X1 U921 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XOR2_X1 U922 ( .A(n1245), .B(n1246), .Z(G21) );
NAND3_X1 U923 ( .A1(n1144), .A2(n1247), .A3(KEYINPUT48), .ZN(n1246) );
XNOR2_X1 U924 ( .A(KEYINPUT37), .B(n1198), .ZN(n1247) );
OR2_X1 U925 ( .A1(n1220), .A2(n1248), .ZN(n1198) );
NAND2_X1 U926 ( .A1(n1025), .A2(n1189), .ZN(n1220) );
XNOR2_X1 U927 ( .A(G116), .B(n1194), .ZN(G18) );
NAND4_X1 U928 ( .A1(n1202), .A2(n1181), .A3(n1033), .A4(n1144), .ZN(n1194) );
NOR2_X1 U929 ( .A1(n1243), .A2(n1249), .ZN(n1033) );
XOR2_X1 U930 ( .A(G113), .B(n1250), .Z(G15) );
NOR2_X1 U931 ( .A1(n1251), .A2(n1042), .ZN(n1250) );
INV_X1 U932 ( .A(n1144), .ZN(n1042) );
XOR2_X1 U933 ( .A(n1199), .B(KEYINPUT52), .Z(n1251) );
NAND3_X1 U934 ( .A1(n1202), .A2(n1181), .A3(n1032), .ZN(n1199) );
INV_X1 U935 ( .A(n1232), .ZN(n1032) );
NAND2_X1 U936 ( .A1(n1252), .A2(n1249), .ZN(n1232) );
INV_X1 U937 ( .A(n1244), .ZN(n1249) );
XNOR2_X1 U938 ( .A(KEYINPUT22), .B(n1243), .ZN(n1252) );
INV_X1 U939 ( .A(n1035), .ZN(n1181) );
NAND2_X1 U940 ( .A1(n1055), .A2(n1238), .ZN(n1035) );
INV_X1 U941 ( .A(n1248), .ZN(n1202) );
NAND2_X1 U942 ( .A1(n1201), .A2(n1020), .ZN(n1248) );
NAND2_X1 U943 ( .A1(n1253), .A2(n1254), .ZN(n1020) );
OR3_X1 U944 ( .A1(n1059), .A2(n1052), .A3(KEYINPUT30), .ZN(n1254) );
INV_X1 U945 ( .A(n1053), .ZN(n1059) );
NAND2_X1 U946 ( .A1(KEYINPUT30), .A2(n1200), .ZN(n1253) );
XOR2_X1 U947 ( .A(n1195), .B(n1255), .Z(G12) );
XOR2_X1 U948 ( .A(KEYINPUT16), .B(G110), .Z(n1255) );
NAND3_X1 U949 ( .A1(n1196), .A2(n1026), .A3(n1025), .ZN(n1195) );
NOR2_X1 U950 ( .A1(n1244), .A2(n1243), .ZN(n1025) );
XOR2_X1 U951 ( .A(n1072), .B(G475), .Z(n1243) );
NOR2_X1 U952 ( .A1(n1136), .A2(G902), .ZN(n1072) );
XNOR2_X1 U953 ( .A(n1256), .B(n1257), .ZN(n1136) );
XOR2_X1 U954 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U955 ( .A(G122), .B(G104), .Z(n1259) );
XOR2_X1 U956 ( .A(G131), .B(G125), .Z(n1258) );
XNOR2_X1 U957 ( .A(n1260), .B(n1261), .ZN(n1256) );
XOR2_X1 U958 ( .A(n1262), .B(n1263), .Z(n1261) );
NOR2_X1 U959 ( .A1(G140), .A2(KEYINPUT15), .ZN(n1263) );
AND3_X1 U960 ( .A1(G214), .A2(n1013), .A3(n1264), .ZN(n1262) );
NAND2_X1 U961 ( .A1(n1265), .A2(n1069), .ZN(n1244) );
NAND2_X1 U962 ( .A1(n1070), .A2(n1266), .ZN(n1069) );
OR2_X1 U963 ( .A1(n1266), .A2(n1070), .ZN(n1265) );
NOR2_X1 U964 ( .A1(n1132), .A2(G902), .ZN(n1070) );
XOR2_X1 U965 ( .A(n1267), .B(n1268), .Z(n1132) );
XOR2_X1 U966 ( .A(G116), .B(n1269), .Z(n1268) );
XOR2_X1 U967 ( .A(KEYINPUT19), .B(G122), .Z(n1269) );
XOR2_X1 U968 ( .A(n1270), .B(n1271), .Z(n1267) );
XOR2_X1 U969 ( .A(n1010), .B(n1272), .Z(n1271) );
NAND2_X1 U970 ( .A1(KEYINPUT41), .A2(n1273), .ZN(n1272) );
XOR2_X1 U971 ( .A(G128), .B(n1274), .Z(n1273) );
XOR2_X1 U972 ( .A(G143), .B(G134), .Z(n1274) );
INV_X1 U973 ( .A(G107), .ZN(n1010) );
NAND2_X1 U974 ( .A1(n1275), .A2(G217), .ZN(n1270) );
INV_X1 U975 ( .A(G478), .ZN(n1266) );
NAND2_X1 U976 ( .A1(n1276), .A2(n1277), .ZN(n1026) );
OR3_X1 U977 ( .A1(n1055), .A2(n1238), .A3(KEYINPUT18), .ZN(n1277) );
INV_X1 U978 ( .A(n1278), .ZN(n1238) );
NAND2_X1 U979 ( .A1(KEYINPUT18), .A2(n1189), .ZN(n1276) );
NOR2_X1 U980 ( .A1(n1055), .A2(n1278), .ZN(n1189) );
XNOR2_X1 U981 ( .A(n1063), .B(KEYINPUT33), .ZN(n1278) );
XOR2_X1 U982 ( .A(G472), .B(n1279), .Z(n1063) );
NOR2_X1 U983 ( .A1(n1280), .A2(G902), .ZN(n1279) );
NOR2_X1 U984 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U985 ( .A(n1283), .B(KEYINPUT8), .Z(n1282) );
NAND2_X1 U986 ( .A1(n1158), .A2(n1284), .ZN(n1283) );
OR2_X1 U987 ( .A1(n1285), .A2(n1155), .ZN(n1284) );
NOR3_X1 U988 ( .A1(n1158), .A2(n1285), .A3(n1155), .ZN(n1281) );
NOR2_X1 U989 ( .A1(n1153), .A2(n1151), .ZN(n1155) );
AND2_X1 U990 ( .A1(n1286), .A2(n1153), .ZN(n1285) );
XOR2_X1 U991 ( .A(n1151), .B(KEYINPUT1), .Z(n1286) );
NAND3_X1 U992 ( .A1(n1264), .A2(n1013), .A3(G210), .ZN(n1151) );
XNOR2_X1 U993 ( .A(n1287), .B(n1288), .ZN(n1158) );
XOR2_X1 U994 ( .A(KEYINPUT39), .B(n1289), .Z(n1288) );
NOR2_X1 U995 ( .A1(KEYINPUT59), .A2(n1290), .ZN(n1289) );
XOR2_X1 U996 ( .A(G116), .B(n1245), .Z(n1290) );
XOR2_X1 U997 ( .A(n1163), .B(n1260), .Z(n1287) );
XNOR2_X1 U998 ( .A(G113), .B(n1291), .ZN(n1260) );
XOR2_X1 U999 ( .A(n1292), .B(n1293), .Z(n1163) );
XOR2_X1 U1000 ( .A(n1294), .B(n1130), .Z(n1055) );
AND2_X1 U1001 ( .A1(G217), .A2(n1295), .ZN(n1130) );
NAND2_X1 U1002 ( .A1(n1128), .A2(n1172), .ZN(n1294) );
XNOR2_X1 U1003 ( .A(n1296), .B(n1297), .ZN(n1128) );
XOR2_X1 U1004 ( .A(n1292), .B(n1298), .Z(n1297) );
XOR2_X1 U1005 ( .A(n1299), .B(n1300), .Z(n1298) );
NOR2_X1 U1006 ( .A1(KEYINPUT51), .A2(n1301), .ZN(n1300) );
XOR2_X1 U1007 ( .A(KEYINPUT10), .B(G110), .Z(n1301) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1275), .ZN(n1299) );
AND2_X1 U1009 ( .A1(G234), .A2(n1013), .ZN(n1275) );
XNOR2_X1 U1010 ( .A(G128), .B(n1091), .ZN(n1292) );
XOR2_X1 U1011 ( .A(n1302), .B(n1303), .Z(n1296) );
XOR2_X1 U1012 ( .A(G125), .B(G119), .Z(n1303) );
XOR2_X1 U1013 ( .A(G146), .B(n1097), .Z(n1302) );
INV_X1 U1014 ( .A(G140), .ZN(n1097) );
AND3_X1 U1015 ( .A1(n1200), .A2(n1201), .A3(n1144), .ZN(n1196) );
NOR2_X1 U1016 ( .A1(n1044), .A2(n1046), .ZN(n1144) );
INV_X1 U1017 ( .A(n1224), .ZN(n1046) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1304), .ZN(n1224) );
XNOR2_X1 U1019 ( .A(n1305), .B(n1064), .ZN(n1044) );
AND2_X1 U1020 ( .A1(G210), .A2(n1304), .ZN(n1064) );
NAND2_X1 U1021 ( .A1(n1264), .A2(n1172), .ZN(n1304) );
INV_X1 U1022 ( .A(G237), .ZN(n1264) );
NAND2_X1 U1023 ( .A1(KEYINPUT0), .A2(n1066), .ZN(n1305) );
NAND2_X1 U1024 ( .A1(n1306), .A2(n1172), .ZN(n1066) );
XOR2_X1 U1025 ( .A(n1307), .B(n1207), .Z(n1306) );
INV_X1 U1026 ( .A(n1211), .ZN(n1207) );
XOR2_X1 U1027 ( .A(n1308), .B(n1309), .Z(n1211) );
INV_X1 U1028 ( .A(n1123), .ZN(n1309) );
XOR2_X1 U1029 ( .A(n1310), .B(G113), .Z(n1123) );
NAND2_X1 U1030 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND2_X1 U1031 ( .A1(G116), .A2(n1245), .ZN(n1312) );
XOR2_X1 U1032 ( .A(KEYINPUT46), .B(n1313), .Z(n1311) );
NOR2_X1 U1033 ( .A1(G116), .A2(n1245), .ZN(n1313) );
INV_X1 U1034 ( .A(G119), .ZN(n1245) );
XOR2_X1 U1035 ( .A(n1314), .B(n1124), .Z(n1308) );
XNOR2_X1 U1036 ( .A(n1164), .B(n1315), .ZN(n1124) );
XOR2_X1 U1037 ( .A(KEYINPUT5), .B(KEYINPUT40), .Z(n1315) );
NAND2_X1 U1038 ( .A1(KEYINPUT20), .A2(n1120), .ZN(n1314) );
XOR2_X1 U1039 ( .A(G110), .B(G122), .Z(n1120) );
NAND2_X1 U1040 ( .A1(KEYINPUT4), .A2(n1206), .ZN(n1307) );
XNOR2_X1 U1041 ( .A(n1316), .B(n1317), .ZN(n1206) );
XOR2_X1 U1042 ( .A(G128), .B(G125), .Z(n1317) );
XNOR2_X1 U1043 ( .A(n1318), .B(n1291), .ZN(n1316) );
NAND2_X1 U1044 ( .A1(G224), .A2(n1013), .ZN(n1318) );
AND2_X1 U1045 ( .A1(n1319), .A2(n1054), .ZN(n1201) );
NAND2_X1 U1046 ( .A1(G237), .A2(G234), .ZN(n1054) );
NAND2_X1 U1047 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U1048 ( .A1(G902), .A2(n1119), .ZN(n1321) );
NOR2_X1 U1049 ( .A1(n1013), .A2(G898), .ZN(n1119) );
NAND2_X1 U1050 ( .A1(G952), .A2(n1013), .ZN(n1320) );
NOR2_X1 U1051 ( .A1(n1053), .A2(n1052), .ZN(n1200) );
AND2_X1 U1052 ( .A1(n1322), .A2(G221), .ZN(n1052) );
XOR2_X1 U1053 ( .A(n1295), .B(KEYINPUT12), .Z(n1322) );
NAND2_X1 U1054 ( .A1(G234), .A2(n1172), .ZN(n1295) );
XOR2_X1 U1055 ( .A(n1323), .B(G469), .Z(n1053) );
NAND2_X1 U1056 ( .A1(n1324), .A2(n1172), .ZN(n1323) );
INV_X1 U1057 ( .A(G902), .ZN(n1172) );
XOR2_X1 U1058 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1059 ( .A(n1162), .B(n1091), .Z(n1326) );
XOR2_X1 U1060 ( .A(G137), .B(KEYINPUT49), .Z(n1091) );
XOR2_X1 U1061 ( .A(n1327), .B(n1328), .Z(n1162) );
XOR2_X1 U1062 ( .A(G140), .B(G110), .Z(n1328) );
NAND2_X1 U1063 ( .A1(G227), .A2(n1013), .ZN(n1327) );
INV_X1 U1064 ( .A(G953), .ZN(n1013) );
XNOR2_X1 U1065 ( .A(n1293), .B(n1329), .ZN(n1325) );
NOR2_X1 U1066 ( .A1(KEYINPUT34), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1067 ( .A(n1164), .B(n1090), .Z(n1330) );
XOR2_X1 U1068 ( .A(G128), .B(n1166), .Z(n1090) );
NOR2_X1 U1069 ( .A1(KEYINPUT38), .A2(n1291), .ZN(n1166) );
XNOR2_X1 U1070 ( .A(G143), .B(G146), .ZN(n1291) );
XOR2_X1 U1071 ( .A(n1153), .B(n1331), .Z(n1164) );
XOR2_X1 U1072 ( .A(G107), .B(G104), .Z(n1331) );
INV_X1 U1073 ( .A(G101), .ZN(n1153) );
XOR2_X1 U1074 ( .A(G134), .B(n1332), .Z(n1293) );
NOR2_X1 U1075 ( .A1(KEYINPUT56), .A2(n1092), .ZN(n1332) );
INV_X1 U1076 ( .A(G131), .ZN(n1092) );
endmodule


