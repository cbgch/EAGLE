//Key = 1010110010010110101101110000101011000010000111000100010100100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330;

XOR2_X1 U739 ( .A(n1022), .B(n1023), .Z(G9) );
XOR2_X1 U740 ( .A(KEYINPUT29), .B(G107), .Z(n1023) );
NOR2_X1 U741 ( .A1(KEYINPUT3), .A2(n1024), .ZN(n1022) );
NOR2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR4_X1 U743 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
XOR2_X1 U744 ( .A(n1031), .B(KEYINPUT57), .Z(n1029) );
NAND2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U746 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND3_X1 U747 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1032) );
NAND3_X1 U748 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1038) );
NAND3_X1 U749 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NAND3_X1 U750 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1041) );
XNOR2_X1 U751 ( .A(n1045), .B(KEYINPUT63), .ZN(n1048) );
NAND3_X1 U752 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1040) );
NAND4_X1 U753 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1027) );
NAND3_X1 U754 ( .A1(n1056), .A2(n1057), .A3(n1037), .ZN(n1053) );
NAND2_X1 U755 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
INV_X1 U756 ( .A(n1039), .ZN(n1059) );
NAND3_X1 U757 ( .A1(n1051), .A2(n1060), .A3(KEYINPUT56), .ZN(n1058) );
NAND3_X1 U758 ( .A1(n1061), .A2(n1062), .A3(n1039), .ZN(n1056) );
NAND3_X1 U759 ( .A1(n1060), .A2(n1063), .A3(n1051), .ZN(n1062) );
INV_X1 U760 ( .A(KEYINPUT56), .ZN(n1063) );
NAND2_X1 U761 ( .A1(n1045), .A2(n1064), .ZN(n1061) );
NAND2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U764 ( .A1(n1069), .A2(n1047), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1035), .A2(n1070), .ZN(n1052) );
AND3_X1 U766 ( .A1(n1051), .A2(n1045), .A3(n1039), .ZN(n1035) );
NOR2_X1 U767 ( .A1(KEYINPUT48), .A2(n1071), .ZN(n1039) );
AND2_X1 U768 ( .A1(n1068), .A2(n1047), .ZN(n1051) );
NOR3_X1 U769 ( .A1(n1072), .A2(G953), .A3(G952), .ZN(n1025) );
INV_X1 U770 ( .A(n1054), .ZN(n1072) );
NAND4_X1 U771 ( .A1(n1049), .A2(n1037), .A3(n1073), .A4(n1074), .ZN(n1054) );
NOR4_X1 U772 ( .A1(n1050), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1074) );
XNOR2_X1 U773 ( .A(n1078), .B(KEYINPUT55), .ZN(n1076) );
XNOR2_X1 U774 ( .A(n1079), .B(n1080), .ZN(n1075) );
NAND2_X1 U775 ( .A1(KEYINPUT19), .A2(n1081), .ZN(n1079) );
XNOR2_X1 U776 ( .A(n1082), .B(KEYINPUT37), .ZN(n1073) );
XOR2_X1 U777 ( .A(n1083), .B(n1084), .Z(G72) );
NAND2_X1 U778 ( .A1(G953), .A2(n1085), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1086), .A2(G227), .ZN(n1085) );
XNOR2_X1 U780 ( .A(G900), .B(KEYINPUT22), .ZN(n1086) );
NAND2_X1 U781 ( .A1(KEYINPUT38), .A2(n1087), .ZN(n1083) );
XOR2_X1 U782 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U783 ( .A1(n1055), .A2(n1030), .ZN(n1089) );
NAND3_X1 U784 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1088) );
XOR2_X1 U785 ( .A(n1093), .B(KEYINPUT15), .Z(n1092) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
OR2_X1 U787 ( .A1(n1095), .A2(n1094), .ZN(n1091) );
AND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
OR2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U790 ( .A(n1100), .B(KEYINPUT10), .Z(n1096) );
NAND2_X1 U791 ( .A1(n1101), .A2(n1098), .ZN(n1100) );
XOR2_X1 U792 ( .A(n1102), .B(n1103), .Z(n1098) );
INV_X1 U793 ( .A(G134), .ZN(n1103) );
XNOR2_X1 U794 ( .A(KEYINPUT40), .B(n1104), .ZN(n1101) );
XNOR2_X1 U795 ( .A(n1105), .B(G125), .ZN(n1095) );
NAND2_X1 U796 ( .A1(KEYINPUT2), .A2(n1106), .ZN(n1105) );
XOR2_X1 U797 ( .A(n1107), .B(n1108), .Z(G69) );
XOR2_X1 U798 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U799 ( .A1(n1111), .A2(n1055), .ZN(n1110) );
AND2_X1 U800 ( .A1(G224), .A2(G898), .ZN(n1111) );
NAND2_X1 U801 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
NAND2_X1 U802 ( .A1(n1114), .A2(G953), .ZN(n1113) );
XOR2_X1 U803 ( .A(n1115), .B(n1116), .Z(n1112) );
NAND2_X1 U804 ( .A1(n1055), .A2(n1028), .ZN(n1107) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(G66) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
XOR2_X1 U808 ( .A(KEYINPUT46), .B(n1123), .Z(n1122) );
NOR2_X1 U809 ( .A1(n1117), .A2(n1124), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1125), .B(n1126), .ZN(n1124) );
NAND2_X1 U811 ( .A1(n1121), .A2(G478), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1117), .A2(n1127), .ZN(G60) );
XOR2_X1 U813 ( .A(n1128), .B(n1129), .Z(n1127) );
AND2_X1 U814 ( .A1(G475), .A2(n1121), .ZN(n1129) );
NAND2_X1 U815 ( .A1(KEYINPUT0), .A2(n1130), .ZN(n1128) );
INV_X1 U816 ( .A(n1131), .ZN(n1130) );
XNOR2_X1 U817 ( .A(G104), .B(n1132), .ZN(G6) );
NOR3_X1 U818 ( .A1(n1117), .A2(n1133), .A3(n1134), .ZN(G57) );
NOR2_X1 U819 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U820 ( .A(n1137), .B(KEYINPUT50), .Z(n1136) );
NOR2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
XOR2_X1 U822 ( .A(n1137), .B(KEYINPUT30), .Z(n1139) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(n1137) );
XOR2_X1 U824 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U825 ( .A1(KEYINPUT51), .A2(n1144), .ZN(n1142) );
XOR2_X1 U826 ( .A(n1145), .B(n1146), .Z(n1140) );
NOR2_X1 U827 ( .A1(n1080), .A2(n1147), .ZN(n1146) );
NAND2_X1 U828 ( .A1(KEYINPUT58), .A2(n1148), .ZN(n1145) );
NOR2_X1 U829 ( .A1(n1117), .A2(n1149), .ZN(G54) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U831 ( .A(n1152), .B(n1153), .Z(n1151) );
AND2_X1 U832 ( .A1(G469), .A2(n1121), .ZN(n1153) );
NOR2_X1 U833 ( .A1(KEYINPUT24), .A2(n1154), .ZN(n1152) );
XNOR2_X1 U834 ( .A(n1155), .B(n1099), .ZN(n1154) );
NOR2_X1 U835 ( .A1(n1117), .A2(n1156), .ZN(G51) );
XOR2_X1 U836 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U837 ( .A1(KEYINPUT33), .A2(n1159), .ZN(n1158) );
NAND2_X1 U838 ( .A1(n1121), .A2(G210), .ZN(n1157) );
INV_X1 U839 ( .A(n1147), .ZN(n1121) );
NAND2_X1 U840 ( .A1(G902), .A2(n1160), .ZN(n1147) );
OR2_X1 U841 ( .A1(n1028), .A2(n1030), .ZN(n1160) );
NAND4_X1 U842 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1030) );
AND4_X1 U843 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NAND2_X1 U844 ( .A1(n1046), .A2(n1169), .ZN(n1163) );
NAND2_X1 U845 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NAND2_X1 U846 ( .A1(n1172), .A2(n1067), .ZN(n1170) );
NAND4_X1 U847 ( .A1(n1173), .A2(n1069), .A3(n1174), .A4(n1175), .ZN(n1161) );
XOR2_X1 U848 ( .A(KEYINPUT1), .B(n1070), .Z(n1174) );
NAND4_X1 U849 ( .A1(n1132), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1028) );
AND4_X1 U850 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1024), .ZN(n1178) );
NAND3_X1 U851 ( .A1(n1046), .A2(n1182), .A3(n1070), .ZN(n1024) );
OR2_X1 U852 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
NOR3_X1 U853 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1177) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1188) );
NOR3_X1 U856 ( .A1(n1192), .A2(n1044), .A3(n1193), .ZN(n1191) );
AND3_X1 U857 ( .A1(n1194), .A2(n1067), .A3(n1069), .ZN(n1190) );
AND3_X1 U858 ( .A1(n1195), .A2(n1184), .A3(n1196), .ZN(n1194) );
INV_X1 U859 ( .A(KEYINPUT23), .ZN(n1184) );
NOR4_X1 U860 ( .A1(n1037), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1186) );
INV_X1 U861 ( .A(KEYINPUT35), .ZN(n1199) );
NAND2_X1 U862 ( .A1(n1082), .A2(n1077), .ZN(n1197) );
NOR2_X1 U863 ( .A1(KEYINPUT35), .A2(n1200), .ZN(n1185) );
NAND3_X1 U864 ( .A1(n1070), .A2(n1182), .A3(n1069), .ZN(n1132) );
NOR2_X1 U865 ( .A1(n1055), .A2(G952), .ZN(n1117) );
XNOR2_X1 U866 ( .A(G146), .B(n1201), .ZN(G48) );
NAND4_X1 U867 ( .A1(n1202), .A2(n1173), .A3(n1069), .A4(n1070), .ZN(n1201) );
XOR2_X1 U868 ( .A(n1175), .B(KEYINPUT52), .Z(n1202) );
XNOR2_X1 U869 ( .A(G143), .B(n1162), .ZN(G45) );
NAND4_X1 U870 ( .A1(n1070), .A2(n1060), .A3(n1067), .A4(n1203), .ZN(n1162) );
AND3_X1 U871 ( .A1(n1082), .A2(n1175), .A3(n1077), .ZN(n1203) );
XNOR2_X1 U872 ( .A(G140), .B(n1168), .ZN(G42) );
NAND2_X1 U873 ( .A1(n1172), .A2(n1204), .ZN(n1168) );
NAND2_X1 U874 ( .A1(n1205), .A2(n1206), .ZN(G39) );
NAND2_X1 U875 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U876 ( .A1(G137), .A2(n1209), .ZN(n1205) );
NAND2_X1 U877 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U878 ( .A1(KEYINPUT60), .A2(n1212), .ZN(n1211) );
OR2_X1 U879 ( .A1(n1207), .A2(KEYINPUT60), .ZN(n1210) );
AND2_X1 U880 ( .A1(KEYINPUT8), .A2(n1212), .ZN(n1207) );
INV_X1 U881 ( .A(n1167), .ZN(n1212) );
NAND3_X1 U882 ( .A1(n1043), .A2(n1213), .A3(n1172), .ZN(n1167) );
XNOR2_X1 U883 ( .A(G134), .B(n1214), .ZN(G36) );
NAND3_X1 U884 ( .A1(n1046), .A2(n1215), .A3(n1172), .ZN(n1214) );
XOR2_X1 U885 ( .A(KEYINPUT27), .B(n1067), .Z(n1215) );
XNOR2_X1 U886 ( .A(G131), .B(n1166), .ZN(G33) );
NAND3_X1 U887 ( .A1(n1069), .A2(n1067), .A3(n1172), .ZN(n1166) );
AND3_X1 U888 ( .A1(n1070), .A2(n1175), .A3(n1045), .ZN(n1172) );
AND2_X1 U889 ( .A1(n1049), .A2(n1216), .ZN(n1045) );
INV_X1 U890 ( .A(n1217), .ZN(n1049) );
XOR2_X1 U891 ( .A(n1218), .B(n1219), .Z(G30) );
NAND2_X1 U892 ( .A1(KEYINPUT49), .A2(G128), .ZN(n1219) );
NAND2_X1 U893 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
INV_X1 U894 ( .A(n1171), .ZN(n1221) );
NAND3_X1 U895 ( .A1(n1070), .A2(n1175), .A3(n1173), .ZN(n1171) );
AND3_X1 U896 ( .A1(n1078), .A2(n1213), .A3(n1060), .ZN(n1173) );
XNOR2_X1 U897 ( .A(n1046), .B(KEYINPUT16), .ZN(n1220) );
XNOR2_X1 U898 ( .A(G101), .B(n1176), .ZN(G3) );
NAND4_X1 U899 ( .A1(n1067), .A2(n1068), .A3(n1070), .A4(n1222), .ZN(n1176) );
XNOR2_X1 U900 ( .A(G125), .B(n1165), .ZN(G27) );
NAND4_X1 U901 ( .A1(n1204), .A2(n1037), .A3(n1060), .A4(n1175), .ZN(n1165) );
NAND2_X1 U902 ( .A1(n1223), .A2(n1224), .ZN(n1175) );
OR3_X1 U903 ( .A1(n1225), .A2(n1071), .A3(n1090), .ZN(n1224) );
NAND2_X1 U904 ( .A1(n1226), .A2(G953), .ZN(n1090) );
XNOR2_X1 U905 ( .A(G900), .B(KEYINPUT62), .ZN(n1226) );
INV_X1 U906 ( .A(n1227), .ZN(n1071) );
AND3_X1 U907 ( .A1(n1044), .A2(n1078), .A3(n1069), .ZN(n1204) );
XNOR2_X1 U908 ( .A(G122), .B(n1200), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1037), .A2(n1182), .A3(n1082), .A4(n1077), .ZN(n1200) );
INV_X1 U910 ( .A(n1198), .ZN(n1182) );
NAND2_X1 U911 ( .A1(n1222), .A2(n1047), .ZN(n1198) );
NOR2_X1 U912 ( .A1(n1213), .A2(n1078), .ZN(n1047) );
XOR2_X1 U913 ( .A(n1228), .B(n1229), .Z(G21) );
XOR2_X1 U914 ( .A(KEYINPUT41), .B(G119), .Z(n1229) );
NOR4_X1 U915 ( .A1(n1230), .A2(n1231), .A3(n1189), .A4(n1192), .ZN(n1228) );
NAND2_X1 U916 ( .A1(n1213), .A2(n1196), .ZN(n1231) );
XNOR2_X1 U917 ( .A(n1060), .B(KEYINPUT47), .ZN(n1230) );
XNOR2_X1 U918 ( .A(G116), .B(n1180), .ZN(G18) );
NAND4_X1 U919 ( .A1(n1067), .A2(n1037), .A3(n1046), .A4(n1222), .ZN(n1180) );
NOR2_X1 U920 ( .A1(n1077), .A2(n1232), .ZN(n1046) );
XNOR2_X1 U921 ( .A(G113), .B(n1183), .ZN(G15) );
NAND4_X1 U922 ( .A1(n1069), .A2(n1067), .A3(n1037), .A4(n1222), .ZN(n1183) );
INV_X1 U923 ( .A(n1189), .ZN(n1037) );
NAND2_X1 U924 ( .A1(n1034), .A2(n1233), .ZN(n1189) );
NOR2_X1 U925 ( .A1(n1078), .A2(n1044), .ZN(n1067) );
AND2_X1 U926 ( .A1(n1232), .A2(n1077), .ZN(n1069) );
INV_X1 U927 ( .A(n1082), .ZN(n1232) );
XNOR2_X1 U928 ( .A(G110), .B(n1179), .ZN(G12) );
NAND4_X1 U929 ( .A1(n1043), .A2(n1070), .A3(n1222), .A4(n1044), .ZN(n1179) );
INV_X1 U930 ( .A(n1213), .ZN(n1044) );
NAND2_X1 U931 ( .A1(n1234), .A2(n1235), .ZN(n1213) );
NAND2_X1 U932 ( .A1(n1236), .A2(n1080), .ZN(n1235) );
XOR2_X1 U933 ( .A(KEYINPUT28), .B(n1237), .Z(n1234) );
NOR2_X1 U934 ( .A1(n1236), .A2(n1080), .ZN(n1237) );
INV_X1 U935 ( .A(G472), .ZN(n1080) );
INV_X1 U936 ( .A(n1081), .ZN(n1236) );
NAND2_X1 U937 ( .A1(n1238), .A2(n1225), .ZN(n1081) );
XOR2_X1 U938 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U939 ( .A(n1241), .B(n1148), .Z(n1240) );
XNOR2_X1 U940 ( .A(n1242), .B(n1243), .ZN(n1148) );
NOR2_X1 U941 ( .A1(KEYINPUT54), .A2(n1135), .ZN(n1241) );
INV_X1 U942 ( .A(n1138), .ZN(n1135) );
XOR2_X1 U943 ( .A(n1244), .B(n1245), .Z(n1138) );
INV_X1 U944 ( .A(G101), .ZN(n1245) );
NAND3_X1 U945 ( .A1(n1246), .A2(n1055), .A3(G210), .ZN(n1244) );
XNOR2_X1 U946 ( .A(n1143), .B(n1144), .ZN(n1239) );
XNOR2_X1 U947 ( .A(n1247), .B(G113), .ZN(n1144) );
NAND2_X1 U948 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U949 ( .A1(G119), .A2(n1250), .ZN(n1249) );
XOR2_X1 U950 ( .A(KEYINPUT43), .B(n1251), .Z(n1248) );
NOR2_X1 U951 ( .A1(G119), .A2(n1250), .ZN(n1251) );
INV_X1 U952 ( .A(n1193), .ZN(n1222) );
NAND2_X1 U953 ( .A1(n1060), .A2(n1196), .ZN(n1193) );
NAND2_X1 U954 ( .A1(n1223), .A2(n1252), .ZN(n1196) );
NAND4_X1 U955 ( .A1(n1114), .A2(G953), .A3(G902), .A4(n1227), .ZN(n1252) );
XNOR2_X1 U956 ( .A(G898), .B(KEYINPUT20), .ZN(n1114) );
NAND3_X1 U957 ( .A1(n1227), .A2(n1055), .A3(G952), .ZN(n1223) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1227) );
INV_X1 U959 ( .A(n1195), .ZN(n1060) );
NAND2_X1 U960 ( .A1(n1216), .A2(n1217), .ZN(n1195) );
NAND2_X1 U961 ( .A1(n1253), .A2(n1254), .ZN(n1217) );
NAND2_X1 U962 ( .A1(G210), .A2(n1255), .ZN(n1254) );
NAND2_X1 U963 ( .A1(n1225), .A2(n1256), .ZN(n1255) );
OR2_X1 U964 ( .A1(n1246), .A2(n1257), .ZN(n1256) );
NAND3_X1 U965 ( .A1(n1258), .A2(n1225), .A3(n1257), .ZN(n1253) );
XOR2_X1 U966 ( .A(n1159), .B(KEYINPUT5), .Z(n1257) );
XOR2_X1 U967 ( .A(n1259), .B(n1260), .Z(n1159) );
XOR2_X1 U968 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U969 ( .A(KEYINPUT4), .B(n1263), .ZN(n1262) );
NOR2_X1 U970 ( .A1(KEYINPUT12), .A2(n1115), .ZN(n1263) );
XNOR2_X1 U971 ( .A(G110), .B(n1264), .ZN(n1115) );
NAND2_X1 U972 ( .A1(G224), .A2(n1055), .ZN(n1261) );
XNOR2_X1 U973 ( .A(n1116), .B(n1265), .ZN(n1259) );
XNOR2_X1 U974 ( .A(n1266), .B(n1242), .ZN(n1265) );
XNOR2_X1 U975 ( .A(n1267), .B(n1268), .ZN(n1116) );
XNOR2_X1 U976 ( .A(n1269), .B(n1270), .ZN(n1268) );
INV_X1 U977 ( .A(n1271), .ZN(n1270) );
NOR2_X1 U978 ( .A1(G119), .A2(KEYINPUT34), .ZN(n1269) );
XNOR2_X1 U979 ( .A(G104), .B(n1272), .ZN(n1267) );
XNOR2_X1 U980 ( .A(n1250), .B(G113), .ZN(n1272) );
INV_X1 U981 ( .A(G116), .ZN(n1250) );
NAND2_X1 U982 ( .A1(G210), .A2(G237), .ZN(n1258) );
XNOR2_X1 U983 ( .A(n1050), .B(KEYINPUT59), .ZN(n1216) );
AND2_X1 U984 ( .A1(G214), .A2(n1273), .ZN(n1050) );
NAND2_X1 U985 ( .A1(n1225), .A2(n1246), .ZN(n1273) );
NOR2_X1 U986 ( .A1(n1034), .A2(n1036), .ZN(n1070) );
INV_X1 U987 ( .A(n1233), .ZN(n1036) );
NAND2_X1 U988 ( .A1(n1274), .A2(n1275), .ZN(n1233) );
XNOR2_X1 U989 ( .A(G221), .B(KEYINPUT14), .ZN(n1274) );
XOR2_X1 U990 ( .A(n1276), .B(G469), .Z(n1034) );
NAND2_X1 U991 ( .A1(n1277), .A2(n1225), .ZN(n1276) );
XOR2_X1 U992 ( .A(n1150), .B(n1278), .Z(n1277) );
NOR2_X1 U993 ( .A1(KEYINPUT39), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U994 ( .A(n1280), .B(n1281), .ZN(n1279) );
INV_X1 U995 ( .A(n1155), .ZN(n1281) );
XOR2_X1 U996 ( .A(n1271), .B(n1282), .Z(n1155) );
NOR2_X1 U997 ( .A1(G104), .A2(KEYINPUT17), .ZN(n1282) );
XOR2_X1 U998 ( .A(G101), .B(G107), .Z(n1271) );
NAND2_X1 U999 ( .A1(KEYINPUT45), .A2(n1104), .ZN(n1280) );
INV_X1 U1000 ( .A(n1099), .ZN(n1104) );
XNOR2_X1 U1001 ( .A(n1283), .B(G128), .ZN(n1099) );
NAND2_X1 U1002 ( .A1(n1284), .A2(KEYINPUT32), .ZN(n1283) );
XNOR2_X1 U1003 ( .A(G143), .B(n1243), .ZN(n1284) );
XNOR2_X1 U1004 ( .A(n1143), .B(n1285), .ZN(n1150) );
XOR2_X1 U1005 ( .A(n1286), .B(n1287), .Z(n1285) );
AND2_X1 U1006 ( .A1(n1055), .A2(G227), .ZN(n1286) );
XNOR2_X1 U1007 ( .A(n1102), .B(n1288), .ZN(n1143) );
NOR2_X1 U1008 ( .A1(G134), .A2(KEYINPUT42), .ZN(n1288) );
XNOR2_X1 U1009 ( .A(G131), .B(n1289), .ZN(n1102) );
XNOR2_X1 U1010 ( .A(KEYINPUT61), .B(n1208), .ZN(n1289) );
INV_X1 U1011 ( .A(G137), .ZN(n1208) );
INV_X1 U1012 ( .A(n1192), .ZN(n1043) );
NAND2_X1 U1013 ( .A1(n1068), .A2(n1078), .ZN(n1192) );
XNOR2_X1 U1014 ( .A(n1290), .B(n1123), .ZN(n1078) );
AND2_X1 U1015 ( .A1(G217), .A2(n1275), .ZN(n1123) );
NAND2_X1 U1016 ( .A1(G234), .A2(n1225), .ZN(n1275) );
NAND2_X1 U1017 ( .A1(n1120), .A2(n1225), .ZN(n1290) );
INV_X1 U1018 ( .A(G902), .ZN(n1225) );
XNOR2_X1 U1019 ( .A(n1291), .B(n1292), .ZN(n1120) );
XOR2_X1 U1020 ( .A(n1266), .B(n1293), .Z(n1292) );
XOR2_X1 U1021 ( .A(n1294), .B(n1287), .Z(n1293) );
XNOR2_X1 U1022 ( .A(G110), .B(n1106), .ZN(n1287) );
INV_X1 U1023 ( .A(G140), .ZN(n1106) );
NOR2_X1 U1024 ( .A1(G137), .A2(KEYINPUT31), .ZN(n1294) );
XOR2_X1 U1025 ( .A(G125), .B(n1243), .Z(n1266) );
XOR2_X1 U1026 ( .A(n1295), .B(n1296), .Z(n1291) );
XOR2_X1 U1027 ( .A(KEYINPUT7), .B(G128), .Z(n1296) );
XOR2_X1 U1028 ( .A(n1297), .B(G119), .Z(n1295) );
NAND2_X1 U1029 ( .A1(n1298), .A2(G221), .ZN(n1297) );
NOR2_X1 U1030 ( .A1(n1082), .A2(n1077), .ZN(n1068) );
XOR2_X1 U1031 ( .A(G475), .B(n1299), .Z(n1077) );
NOR2_X1 U1032 ( .A1(G902), .A2(n1131), .ZN(n1299) );
NAND3_X1 U1033 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1131) );
NAND2_X1 U1034 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U1035 ( .A1(KEYINPUT11), .A2(n1305), .ZN(n1304) );
XOR2_X1 U1036 ( .A(n1306), .B(n1307), .Z(n1303) );
NAND4_X1 U1037 ( .A1(n1308), .A2(n1305), .A3(KEYINPUT11), .A4(n1309), .ZN(n1301) );
XNOR2_X1 U1038 ( .A(n1307), .B(n1306), .ZN(n1308) );
XOR2_X1 U1039 ( .A(n1310), .B(n1311), .Z(n1306) );
NOR2_X1 U1040 ( .A1(KEYINPUT25), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1041 ( .A(n1243), .B(n1313), .Z(n1312) );
XOR2_X1 U1042 ( .A(KEYINPUT7), .B(KEYINPUT18), .Z(n1313) );
XOR2_X1 U1043 ( .A(G146), .B(KEYINPUT44), .Z(n1243) );
XOR2_X1 U1044 ( .A(n1314), .B(G125), .Z(n1310) );
NAND3_X1 U1045 ( .A1(n1246), .A2(n1055), .A3(n1315), .ZN(n1314) );
XNOR2_X1 U1046 ( .A(G214), .B(KEYINPUT13), .ZN(n1315) );
INV_X1 U1047 ( .A(G237), .ZN(n1246) );
XNOR2_X1 U1048 ( .A(n1316), .B(n1317), .ZN(n1307) );
XOR2_X1 U1049 ( .A(KEYINPUT6), .B(G143), .Z(n1317) );
XNOR2_X1 U1050 ( .A(G131), .B(G140), .ZN(n1316) );
OR2_X1 U1051 ( .A1(n1309), .A2(n1305), .ZN(n1300) );
XNOR2_X1 U1052 ( .A(n1318), .B(G104), .ZN(n1305) );
NAND2_X1 U1053 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U1054 ( .A1(G113), .A2(n1264), .ZN(n1320) );
XOR2_X1 U1055 ( .A(KEYINPUT21), .B(n1321), .Z(n1319) );
NOR2_X1 U1056 ( .A1(G113), .A2(n1264), .ZN(n1321) );
INV_X1 U1057 ( .A(KEYINPUT36), .ZN(n1309) );
XOR2_X1 U1058 ( .A(G478), .B(n1322), .Z(n1082) );
NOR2_X1 U1059 ( .A1(G902), .A2(n1126), .ZN(n1322) );
XNOR2_X1 U1060 ( .A(n1323), .B(n1324), .ZN(n1126) );
XNOR2_X1 U1061 ( .A(n1325), .B(n1242), .ZN(n1324) );
XNOR2_X1 U1062 ( .A(G128), .B(G143), .ZN(n1242) );
NOR2_X1 U1063 ( .A1(n1326), .A2(KEYINPUT26), .ZN(n1325) );
AND2_X1 U1064 ( .A1(n1298), .A2(G217), .ZN(n1326) );
AND2_X1 U1065 ( .A1(G234), .A2(n1055), .ZN(n1298) );
INV_X1 U1066 ( .A(G953), .ZN(n1055) );
XOR2_X1 U1067 ( .A(n1327), .B(n1328), .Z(n1323) );
NOR2_X1 U1068 ( .A1(KEYINPUT9), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1069 ( .A(G107), .B(n1330), .Z(n1329) );
XNOR2_X1 U1070 ( .A(n1264), .B(G116), .ZN(n1330) );
INV_X1 U1071 ( .A(G122), .ZN(n1264) );
XNOR2_X1 U1072 ( .A(G134), .B(KEYINPUT53), .ZN(n1327) );
endmodule


