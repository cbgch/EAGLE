//Key = 0110101011110001110000001111010010111010100011101101110110100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;

XOR2_X1 U734 ( .A(n1006), .B(n1007), .Z(G9) );
NOR2_X1 U735 ( .A1(KEYINPUT5), .A2(n1008), .ZN(n1007) );
INV_X1 U736 ( .A(G107), .ZN(n1008) );
NOR2_X1 U737 ( .A1(n1009), .A2(n1010), .ZN(G75) );
NOR4_X1 U738 ( .A1(G953), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1010) );
NOR2_X1 U739 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR2_X1 U740 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR3_X1 U741 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NOR3_X1 U742 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1019) );
NOR2_X1 U743 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
XOR2_X1 U744 ( .A(KEYINPUT58), .B(n1026), .Z(n1025) );
NOR3_X1 U745 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1022) );
NOR2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1021) );
NOR2_X1 U747 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
XOR2_X1 U748 ( .A(n1034), .B(KEYINPUT55), .Z(n1033) );
NAND2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR3_X1 U750 ( .A1(n1031), .A2(n1037), .A3(n1029), .ZN(n1016) );
INV_X1 U751 ( .A(n1026), .ZN(n1029) );
NOR3_X1 U752 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NOR2_X1 U753 ( .A1(n1041), .A2(n1020), .ZN(n1040) );
NOR2_X1 U754 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
AND2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1038) );
NOR3_X1 U756 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1009) );
AND4_X1 U757 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1011) );
NOR4_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1035), .A4(n1052), .ZN(n1049) );
INV_X1 U759 ( .A(n1053), .ZN(n1052) );
NAND3_X1 U760 ( .A1(n1054), .A2(n1028), .A3(n1055), .ZN(n1050) );
NOR3_X1 U761 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1048) );
NOR2_X1 U762 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
INV_X1 U763 ( .A(n1061), .ZN(n1057) );
NAND2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(G72) );
NAND3_X1 U765 ( .A1(n1064), .A2(n1065), .A3(G953), .ZN(n1063) );
XOR2_X1 U766 ( .A(n1066), .B(KEYINPUT30), .Z(n1062) );
NAND3_X1 U767 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1065), .ZN(n1069) );
OR3_X1 U769 ( .A1(n1065), .A2(n1070), .A3(G953), .ZN(n1068) );
NAND2_X1 U770 ( .A1(G953), .A2(n1071), .ZN(n1067) );
OR2_X1 U771 ( .A1(n1065), .A2(n1064), .ZN(n1071) );
NAND2_X1 U772 ( .A1(G900), .A2(G227), .ZN(n1064) );
NAND2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(n1065) );
NAND2_X1 U774 ( .A1(G953), .A2(n1074), .ZN(n1073) );
XOR2_X1 U775 ( .A(n1075), .B(KEYINPUT8), .Z(n1072) );
NAND2_X1 U776 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U777 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U778 ( .A(KEYINPUT52), .B(n1080), .Z(n1076) );
NOR2_X1 U779 ( .A1(n1078), .A2(n1079), .ZN(n1080) );
XOR2_X1 U780 ( .A(n1081), .B(G140), .Z(n1079) );
NAND2_X1 U781 ( .A1(KEYINPUT34), .A2(n1082), .ZN(n1081) );
XOR2_X1 U782 ( .A(n1083), .B(n1084), .Z(G69) );
XOR2_X1 U783 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U784 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U785 ( .A1(G953), .A2(n1089), .ZN(n1088) );
XOR2_X1 U786 ( .A(n1090), .B(n1091), .Z(n1087) );
XNOR2_X1 U787 ( .A(n1092), .B(n1093), .ZN(n1091) );
XOR2_X1 U788 ( .A(n1094), .B(n1095), .Z(n1090) );
XOR2_X1 U789 ( .A(G107), .B(n1096), .Z(n1095) );
NAND2_X1 U790 ( .A1(n1097), .A2(KEYINPUT24), .ZN(n1094) );
XNOR2_X1 U791 ( .A(G122), .B(n1098), .ZN(n1097) );
NAND2_X1 U792 ( .A1(G953), .A2(n1099), .ZN(n1085) );
NAND2_X1 U793 ( .A1(n1100), .A2(G898), .ZN(n1099) );
XOR2_X1 U794 ( .A(n1101), .B(KEYINPUT2), .Z(n1100) );
NOR2_X1 U795 ( .A1(n1102), .A2(G953), .ZN(n1083) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1104), .ZN(G66) );
XOR2_X1 U797 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U798 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U799 ( .A1(n1103), .A2(n1109), .ZN(G63) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U801 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U802 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U803 ( .A1(n1107), .A2(G478), .ZN(n1112) );
NOR2_X1 U804 ( .A1(n1114), .A2(n1115), .ZN(n1110) );
INV_X1 U805 ( .A(KEYINPUT33), .ZN(n1115) );
NOR2_X1 U806 ( .A1(n1103), .A2(n1116), .ZN(G60) );
XOR2_X1 U807 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U808 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U809 ( .A(KEYINPUT50), .B(KEYINPUT15), .ZN(n1120) );
NAND3_X1 U810 ( .A1(n1121), .A2(n1122), .A3(G475), .ZN(n1117) );
OR2_X1 U811 ( .A1(n1107), .A2(KEYINPUT18), .ZN(n1122) );
NAND2_X1 U812 ( .A1(KEYINPUT18), .A2(n1123), .ZN(n1121) );
NAND2_X1 U813 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
INV_X1 U814 ( .A(n1013), .ZN(n1124) );
XOR2_X1 U815 ( .A(n1126), .B(n1127), .Z(G6) );
XOR2_X1 U816 ( .A(KEYINPUT56), .B(G104), .Z(n1127) );
NOR2_X1 U817 ( .A1(n1103), .A2(n1128), .ZN(G57) );
XNOR2_X1 U818 ( .A(n1129), .B(n1130), .ZN(n1128) );
XOR2_X1 U819 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR3_X1 U820 ( .A1(n1133), .A2(KEYINPUT22), .A3(n1134), .ZN(n1131) );
INV_X1 U821 ( .A(G472), .ZN(n1134) );
NOR2_X1 U822 ( .A1(n1103), .A2(n1135), .ZN(G54) );
XOR2_X1 U823 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U825 ( .A(n1140), .B(KEYINPUT36), .Z(n1139) );
NAND2_X1 U826 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U827 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U828 ( .A1(KEYINPUT29), .A2(n1145), .ZN(n1144) );
NAND2_X1 U829 ( .A1(KEYINPUT48), .A2(n1146), .ZN(n1145) );
NAND2_X1 U830 ( .A1(n1147), .A2(n1148), .ZN(n1141) );
NAND2_X1 U831 ( .A1(KEYINPUT48), .A2(n1149), .ZN(n1148) );
NAND2_X1 U832 ( .A1(KEYINPUT29), .A2(n1150), .ZN(n1149) );
INV_X1 U833 ( .A(n1143), .ZN(n1150) );
XNOR2_X1 U834 ( .A(n1151), .B(KEYINPUT19), .ZN(n1143) );
INV_X1 U835 ( .A(n1146), .ZN(n1147) );
NAND2_X1 U836 ( .A1(KEYINPUT49), .A2(n1152), .ZN(n1138) );
NAND2_X1 U837 ( .A1(n1107), .A2(G469), .ZN(n1152) );
XOR2_X1 U838 ( .A(n1078), .B(n1153), .Z(n1136) );
XOR2_X1 U839 ( .A(n1154), .B(n1155), .Z(n1078) );
NOR2_X1 U840 ( .A1(n1103), .A2(n1156), .ZN(G51) );
XOR2_X1 U841 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U842 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND3_X1 U843 ( .A1(n1107), .A2(G210), .A3(n1161), .ZN(n1159) );
XOR2_X1 U844 ( .A(n1162), .B(KEYINPUT3), .Z(n1161) );
INV_X1 U845 ( .A(n1133), .ZN(n1107) );
NAND2_X1 U846 ( .A1(n1125), .A2(n1013), .ZN(n1133) );
NAND2_X1 U847 ( .A1(n1102), .A2(n1070), .ZN(n1013) );
AND4_X1 U848 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1070) );
AND4_X1 U849 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR2_X1 U850 ( .A1(n1171), .A2(n1172), .ZN(n1165) );
NOR2_X1 U851 ( .A1(n1173), .A2(n1031), .ZN(n1172) );
NOR2_X1 U852 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U853 ( .A(KEYINPUT59), .B(n1176), .Z(n1175) );
NAND2_X1 U854 ( .A1(n1177), .A2(n1178), .ZN(n1164) );
INV_X1 U855 ( .A(KEYINPUT39), .ZN(n1178) );
NAND4_X1 U856 ( .A1(n1179), .A2(n1024), .A3(n1180), .A4(KEYINPUT39), .ZN(n1163) );
AND4_X1 U857 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1102) );
NOR4_X1 U858 ( .A1(n1185), .A2(n1006), .A3(n1186), .A4(n1187), .ZN(n1184) );
INV_X1 U859 ( .A(n1188), .ZN(n1187) );
AND3_X1 U860 ( .A1(n1189), .A2(n1190), .A3(n1042), .ZN(n1006) );
NOR2_X1 U861 ( .A1(n1191), .A2(n1192), .ZN(n1185) );
NOR2_X1 U862 ( .A1(n1193), .A2(n1039), .ZN(n1191) );
AND3_X1 U863 ( .A1(KEYINPUT14), .A2(n1020), .A3(n1043), .ZN(n1193) );
INV_X1 U864 ( .A(n1189), .ZN(n1020) );
NOR2_X1 U865 ( .A1(n1194), .A2(n1195), .ZN(n1183) );
NOR2_X1 U866 ( .A1(KEYINPUT14), .A2(n1126), .ZN(n1195) );
NAND3_X1 U867 ( .A1(n1189), .A2(n1190), .A3(n1043), .ZN(n1126) );
INV_X1 U868 ( .A(n1196), .ZN(n1194) );
XOR2_X1 U869 ( .A(G902), .B(KEYINPUT47), .Z(n1125) );
XOR2_X1 U870 ( .A(KEYINPUT45), .B(n1197), .Z(n1157) );
NOR2_X1 U871 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR2_X1 U872 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NOR2_X1 U873 ( .A1(G953), .A2(n1101), .ZN(n1200) );
NOR3_X1 U874 ( .A1(n1202), .A2(G953), .A3(n1101), .ZN(n1198) );
INV_X1 U875 ( .A(G224), .ZN(n1101) );
XNOR2_X1 U876 ( .A(KEYINPUT37), .B(n1201), .ZN(n1202) );
NOR2_X1 U877 ( .A1(n1203), .A2(G952), .ZN(n1103) );
XOR2_X1 U878 ( .A(n1204), .B(n1168), .Z(G48) );
NAND3_X1 U879 ( .A1(n1043), .A2(n1205), .A3(n1206), .ZN(n1168) );
XOR2_X1 U880 ( .A(G143), .B(n1177), .Z(G45) );
AND3_X1 U881 ( .A1(n1179), .A2(n1205), .A3(n1180), .ZN(n1177) );
XNOR2_X1 U882 ( .A(G140), .B(n1170), .ZN(G42) );
NAND3_X1 U883 ( .A1(n1207), .A2(n1032), .A3(n1208), .ZN(n1170) );
XOR2_X1 U884 ( .A(n1209), .B(n1210), .Z(G39) );
NAND2_X1 U885 ( .A1(n1176), .A2(n1207), .ZN(n1210) );
AND2_X1 U886 ( .A1(n1206), .A2(n1044), .ZN(n1176) );
XNOR2_X1 U887 ( .A(G134), .B(n1167), .ZN(G36) );
NAND3_X1 U888 ( .A1(n1180), .A2(n1042), .A3(n1207), .ZN(n1167) );
INV_X1 U889 ( .A(n1031), .ZN(n1207) );
XOR2_X1 U890 ( .A(G131), .B(n1211), .Z(G33) );
NOR2_X1 U891 ( .A1(n1031), .A2(n1212), .ZN(n1211) );
XOR2_X1 U892 ( .A(KEYINPUT4), .B(n1174), .Z(n1212) );
AND2_X1 U893 ( .A1(n1180), .A2(n1043), .ZN(n1174) );
AND3_X1 U894 ( .A1(n1032), .A2(n1213), .A3(n1045), .ZN(n1180) );
NAND2_X1 U895 ( .A1(n1214), .A2(n1028), .ZN(n1031) );
INV_X1 U896 ( .A(n1027), .ZN(n1214) );
XNOR2_X1 U897 ( .A(G128), .B(n1215), .ZN(G30) );
NAND2_X1 U898 ( .A1(KEYINPUT1), .A2(n1171), .ZN(n1215) );
AND3_X1 U899 ( .A1(n1042), .A2(n1205), .A3(n1206), .ZN(n1171) );
AND4_X1 U900 ( .A1(n1032), .A2(n1216), .A3(n1213), .A4(n1217), .ZN(n1206) );
XOR2_X1 U901 ( .A(n1218), .B(n1196), .Z(G3) );
NAND3_X1 U902 ( .A1(n1044), .A2(n1190), .A3(n1045), .ZN(n1196) );
XOR2_X1 U903 ( .A(n1082), .B(n1169), .Z(G27) );
NAND3_X1 U904 ( .A1(n1026), .A2(n1205), .A3(n1208), .ZN(n1169) );
AND4_X1 U905 ( .A1(n1219), .A2(n1043), .A3(n1213), .A4(n1217), .ZN(n1208) );
NAND2_X1 U906 ( .A1(n1015), .A2(n1220), .ZN(n1213) );
NAND4_X1 U907 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1074), .ZN(n1220) );
INV_X1 U908 ( .A(G900), .ZN(n1074) );
XNOR2_X1 U909 ( .A(G122), .B(n1181), .ZN(G24) );
NAND3_X1 U910 ( .A1(n1222), .A2(n1189), .A3(n1179), .ZN(n1181) );
NOR2_X1 U911 ( .A1(n1046), .A2(n1223), .ZN(n1179) );
NOR2_X1 U912 ( .A1(n1217), .A2(n1216), .ZN(n1189) );
XOR2_X1 U913 ( .A(n1224), .B(n1182), .Z(G21) );
NAND4_X1 U914 ( .A1(n1222), .A2(n1044), .A3(n1216), .A4(n1217), .ZN(n1182) );
INV_X1 U915 ( .A(n1219), .ZN(n1216) );
XOR2_X1 U916 ( .A(n1225), .B(n1188), .Z(G18) );
NAND3_X1 U917 ( .A1(n1222), .A2(n1042), .A3(n1045), .ZN(n1188) );
NOR2_X1 U918 ( .A1(n1056), .A2(n1046), .ZN(n1042) );
XOR2_X1 U919 ( .A(G113), .B(n1186), .Z(G15) );
AND3_X1 U920 ( .A1(n1222), .A2(n1043), .A3(n1045), .ZN(n1186) );
NOR2_X1 U921 ( .A1(n1217), .A2(n1219), .ZN(n1045) );
AND2_X1 U922 ( .A1(n1226), .A2(n1046), .ZN(n1043) );
XOR2_X1 U923 ( .A(n1223), .B(KEYINPUT51), .Z(n1226) );
AND3_X1 U924 ( .A1(n1205), .A2(n1227), .A3(n1026), .ZN(n1222) );
NOR2_X1 U925 ( .A1(n1228), .A2(n1035), .ZN(n1026) );
XNOR2_X1 U926 ( .A(G110), .B(n1229), .ZN(G12) );
NAND3_X1 U927 ( .A1(n1039), .A2(n1190), .A3(KEYINPUT11), .ZN(n1229) );
INV_X1 U928 ( .A(n1192), .ZN(n1190) );
NAND3_X1 U929 ( .A1(n1205), .A2(n1227), .A3(n1032), .ZN(n1192) );
NOR2_X1 U930 ( .A1(n1036), .A2(n1035), .ZN(n1032) );
AND2_X1 U931 ( .A1(G221), .A2(n1230), .ZN(n1035) );
INV_X1 U932 ( .A(n1228), .ZN(n1036) );
NAND2_X1 U933 ( .A1(n1053), .A2(n1231), .ZN(n1228) );
NAND2_X1 U934 ( .A1(G469), .A2(n1232), .ZN(n1231) );
XOR2_X1 U935 ( .A(KEYINPUT46), .B(n1059), .Z(n1232) );
NAND2_X1 U936 ( .A1(n1059), .A2(n1060), .ZN(n1053) );
INV_X1 U937 ( .A(G469), .ZN(n1060) );
AND2_X1 U938 ( .A1(n1233), .A2(n1234), .ZN(n1059) );
XOR2_X1 U939 ( .A(n1235), .B(n1236), .Z(n1233) );
XOR2_X1 U940 ( .A(n1155), .B(n1151), .Z(n1236) );
XOR2_X1 U941 ( .A(G110), .B(G140), .Z(n1151) );
XNOR2_X1 U942 ( .A(n1237), .B(n1238), .ZN(n1235) );
NOR2_X1 U943 ( .A1(KEYINPUT60), .A2(n1239), .ZN(n1238) );
XOR2_X1 U944 ( .A(n1146), .B(KEYINPUT7), .Z(n1239) );
NAND2_X1 U945 ( .A1(G227), .A2(n1203), .ZN(n1146) );
NAND2_X1 U946 ( .A1(KEYINPUT62), .A2(n1240), .ZN(n1237) );
XNOR2_X1 U947 ( .A(n1153), .B(n1241), .ZN(n1240) );
XOR2_X1 U948 ( .A(n1154), .B(KEYINPUT61), .Z(n1241) );
NAND3_X1 U949 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1154) );
OR2_X1 U950 ( .A1(n1245), .A2(KEYINPUT53), .ZN(n1244) );
NAND3_X1 U951 ( .A1(KEYINPUT53), .A2(n1246), .A3(n1247), .ZN(n1243) );
INV_X1 U952 ( .A(n1248), .ZN(n1246) );
NAND2_X1 U953 ( .A1(G128), .A2(n1248), .ZN(n1242) );
NAND2_X1 U954 ( .A1(KEYINPUT25), .A2(n1245), .ZN(n1248) );
XOR2_X1 U955 ( .A(G143), .B(n1249), .Z(n1245) );
XOR2_X1 U956 ( .A(KEYINPUT63), .B(G146), .Z(n1249) );
XNOR2_X1 U957 ( .A(n1250), .B(n1251), .ZN(n1153) );
XOR2_X1 U958 ( .A(G104), .B(G101), .Z(n1251) );
NAND2_X1 U959 ( .A1(KEYINPUT38), .A2(n1252), .ZN(n1250) );
XOR2_X1 U960 ( .A(KEYINPUT0), .B(G107), .Z(n1252) );
NAND2_X1 U961 ( .A1(n1015), .A2(n1253), .ZN(n1227) );
NAND4_X1 U962 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1089), .ZN(n1253) );
INV_X1 U963 ( .A(G898), .ZN(n1089) );
NAND3_X1 U964 ( .A1(n1221), .A2(n1203), .A3(G952), .ZN(n1015) );
NAND2_X1 U965 ( .A1(G237), .A2(G234), .ZN(n1221) );
INV_X1 U966 ( .A(n1024), .ZN(n1205) );
NAND2_X1 U967 ( .A1(n1254), .A2(n1027), .ZN(n1024) );
NAND2_X1 U968 ( .A1(n1255), .A2(n1055), .ZN(n1027) );
NAND3_X1 U969 ( .A1(n1256), .A2(n1162), .A3(G210), .ZN(n1055) );
NAND2_X1 U970 ( .A1(n1257), .A2(n1234), .ZN(n1256) );
XOR2_X1 U971 ( .A(n1054), .B(KEYINPUT31), .Z(n1255) );
NAND3_X1 U972 ( .A1(n1258), .A2(n1234), .A3(n1257), .ZN(n1054) );
XOR2_X1 U973 ( .A(n1259), .B(n1260), .Z(n1257) );
INV_X1 U974 ( .A(n1160), .ZN(n1260) );
XOR2_X1 U975 ( .A(n1261), .B(n1262), .Z(n1160) );
XOR2_X1 U976 ( .A(n1263), .B(n1098), .Z(n1262) );
XOR2_X1 U977 ( .A(G110), .B(KEYINPUT26), .Z(n1098) );
XOR2_X1 U978 ( .A(n1264), .B(n1265), .Z(n1261) );
NOR2_X1 U979 ( .A1(KEYINPUT54), .A2(n1266), .ZN(n1265) );
XOR2_X1 U980 ( .A(G113), .B(n1092), .Z(n1266) );
XNOR2_X1 U981 ( .A(n1225), .B(n1267), .ZN(n1092) );
XOR2_X1 U982 ( .A(KEYINPUT57), .B(G119), .Z(n1267) );
XOR2_X1 U983 ( .A(n1218), .B(n1096), .Z(n1264) );
NOR2_X1 U984 ( .A1(KEYINPUT21), .A2(G104), .ZN(n1096) );
INV_X1 U985 ( .A(G101), .ZN(n1218) );
XNOR2_X1 U986 ( .A(n1268), .B(n1201), .ZN(n1259) );
XNOR2_X1 U987 ( .A(G125), .B(n1269), .ZN(n1201) );
NAND3_X1 U988 ( .A1(G224), .A2(n1203), .A3(KEYINPUT9), .ZN(n1268) );
NAND2_X1 U989 ( .A1(G210), .A2(n1162), .ZN(n1258) );
XNOR2_X1 U990 ( .A(KEYINPUT35), .B(n1028), .ZN(n1254) );
NAND2_X1 U991 ( .A1(G214), .A2(n1162), .ZN(n1028) );
NAND2_X1 U992 ( .A1(n1270), .A2(n1271), .ZN(n1162) );
INV_X1 U993 ( .A(G237), .ZN(n1271) );
AND3_X1 U994 ( .A1(n1219), .A2(n1217), .A3(n1044), .ZN(n1039) );
INV_X1 U995 ( .A(n1018), .ZN(n1044) );
NAND2_X1 U996 ( .A1(n1046), .A2(n1272), .ZN(n1018) );
XOR2_X1 U997 ( .A(KEYINPUT27), .B(n1056), .Z(n1272) );
INV_X1 U998 ( .A(n1223), .ZN(n1056) );
XOR2_X1 U999 ( .A(n1273), .B(G475), .Z(n1223) );
OR2_X1 U1000 ( .A1(n1119), .A2(G902), .ZN(n1273) );
XOR2_X1 U1001 ( .A(n1274), .B(n1275), .Z(n1119) );
XOR2_X1 U1002 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U1003 ( .A(G122), .B(G113), .Z(n1277) );
XOR2_X1 U1004 ( .A(G143), .B(G131), .Z(n1276) );
XOR2_X1 U1005 ( .A(n1278), .B(n1279), .Z(n1274) );
XOR2_X1 U1006 ( .A(n1280), .B(G104), .Z(n1278) );
NAND3_X1 U1007 ( .A1(G214), .A2(n1281), .A3(KEYINPUT44), .ZN(n1280) );
XOR2_X1 U1008 ( .A(n1282), .B(G478), .Z(n1046) );
NAND2_X1 U1009 ( .A1(n1114), .A2(n1234), .ZN(n1282) );
XNOR2_X1 U1010 ( .A(n1283), .B(n1284), .ZN(n1114) );
XOR2_X1 U1011 ( .A(n1285), .B(n1286), .Z(n1284) );
NAND2_X1 U1012 ( .A1(n1287), .A2(KEYINPUT10), .ZN(n1285) );
XOR2_X1 U1013 ( .A(n1288), .B(n1263), .Z(n1287) );
XOR2_X1 U1014 ( .A(G107), .B(G122), .Z(n1263) );
NAND2_X1 U1015 ( .A1(KEYINPUT32), .A2(n1225), .ZN(n1288) );
XNOR2_X1 U1016 ( .A(G134), .B(n1289), .ZN(n1283) );
AND4_X1 U1017 ( .A1(n1290), .A2(n1203), .A3(G217), .A4(G234), .ZN(n1289) );
INV_X1 U1018 ( .A(KEYINPUT20), .ZN(n1290) );
NAND3_X1 U1019 ( .A1(n1291), .A2(n1292), .A3(n1061), .ZN(n1217) );
NAND3_X1 U1020 ( .A1(n1293), .A2(n1234), .A3(n1105), .ZN(n1061) );
NAND2_X1 U1021 ( .A1(KEYINPUT28), .A2(n1293), .ZN(n1292) );
NAND2_X1 U1022 ( .A1(n1051), .A2(n1294), .ZN(n1291) );
INV_X1 U1023 ( .A(KEYINPUT28), .ZN(n1294) );
AND2_X1 U1024 ( .A1(n1108), .A2(n1295), .ZN(n1051) );
NAND2_X1 U1025 ( .A1(n1105), .A2(n1234), .ZN(n1295) );
NAND2_X1 U1026 ( .A1(n1296), .A2(n1297), .ZN(n1105) );
NAND3_X1 U1027 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1297) );
XNOR2_X1 U1028 ( .A(n1301), .B(n1302), .ZN(n1300) );
NAND2_X1 U1029 ( .A1(n1303), .A2(n1304), .ZN(n1296) );
NAND2_X1 U1030 ( .A1(n1298), .A2(n1299), .ZN(n1304) );
NAND2_X1 U1031 ( .A1(n1305), .A2(n1279), .ZN(n1299) );
INV_X1 U1032 ( .A(n1306), .ZN(n1279) );
XNOR2_X1 U1033 ( .A(n1307), .B(n1308), .ZN(n1305) );
XNOR2_X1 U1034 ( .A(KEYINPUT16), .B(n1309), .ZN(n1298) );
NAND2_X1 U1035 ( .A1(n1310), .A2(n1306), .ZN(n1309) );
XOR2_X1 U1036 ( .A(n1082), .B(n1311), .Z(n1306) );
XOR2_X1 U1037 ( .A(G146), .B(G140), .Z(n1311) );
INV_X1 U1038 ( .A(G125), .ZN(n1082) );
XOR2_X1 U1039 ( .A(n1307), .B(n1308), .Z(n1310) );
XOR2_X1 U1040 ( .A(G110), .B(G119), .Z(n1308) );
NAND2_X1 U1041 ( .A1(KEYINPUT6), .A2(n1247), .ZN(n1307) );
INV_X1 U1042 ( .A(G128), .ZN(n1247) );
XOR2_X1 U1043 ( .A(n1301), .B(n1302), .Z(n1303) );
NAND2_X1 U1044 ( .A1(KEYINPUT17), .A2(n1209), .ZN(n1302) );
INV_X1 U1045 ( .A(G137), .ZN(n1209) );
NAND3_X1 U1046 ( .A1(G234), .A2(n1203), .A3(G221), .ZN(n1301) );
INV_X1 U1047 ( .A(G953), .ZN(n1203) );
INV_X1 U1048 ( .A(n1293), .ZN(n1108) );
NAND2_X1 U1049 ( .A1(G217), .A2(n1230), .ZN(n1293) );
NAND2_X1 U1050 ( .A1(n1270), .A2(G234), .ZN(n1230) );
XOR2_X1 U1051 ( .A(n1234), .B(KEYINPUT43), .Z(n1270) );
XOR2_X1 U1052 ( .A(n1047), .B(KEYINPUT13), .Z(n1219) );
XOR2_X1 U1053 ( .A(n1312), .B(G472), .Z(n1047) );
NAND2_X1 U1054 ( .A1(n1313), .A2(n1234), .ZN(n1312) );
INV_X1 U1055 ( .A(G902), .ZN(n1234) );
XNOR2_X1 U1056 ( .A(n1132), .B(n1314), .ZN(n1313) );
NOR2_X1 U1057 ( .A1(KEYINPUT23), .A2(n1129), .ZN(n1314) );
XNOR2_X1 U1058 ( .A(n1155), .B(n1269), .ZN(n1129) );
XNOR2_X1 U1059 ( .A(n1286), .B(n1315), .ZN(n1269) );
NOR2_X1 U1060 ( .A1(KEYINPUT12), .A2(n1204), .ZN(n1315) );
INV_X1 U1061 ( .A(G146), .ZN(n1204) );
XNOR2_X1 U1062 ( .A(G128), .B(G143), .ZN(n1286) );
XNOR2_X1 U1063 ( .A(n1316), .B(n1317), .ZN(n1155) );
XOR2_X1 U1064 ( .A(KEYINPUT40), .B(G137), .Z(n1317) );
XNOR2_X1 U1065 ( .A(G131), .B(G134), .ZN(n1316) );
XNOR2_X1 U1066 ( .A(n1318), .B(n1319), .ZN(n1132) );
NOR2_X1 U1067 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NOR2_X1 U1068 ( .A1(n1224), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1069 ( .A(n1225), .B(KEYINPUT41), .Z(n1322) );
INV_X1 U1070 ( .A(G116), .ZN(n1225) );
INV_X1 U1071 ( .A(G119), .ZN(n1224) );
NOR2_X1 U1072 ( .A1(G119), .A2(n1323), .ZN(n1320) );
XOR2_X1 U1073 ( .A(KEYINPUT42), .B(G116), .Z(n1323) );
XOR2_X1 U1074 ( .A(n1324), .B(n1093), .Z(n1318) );
XOR2_X1 U1075 ( .A(G101), .B(G113), .Z(n1093) );
NAND2_X1 U1076 ( .A1(G210), .A2(n1281), .ZN(n1324) );
NOR2_X1 U1077 ( .A1(G953), .A2(G237), .ZN(n1281) );
endmodule


