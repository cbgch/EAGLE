//Key = 0100001001100001101010101111011011001101000110011010101111101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201;

XNOR2_X1 U661 ( .A(G107), .B(n911), .ZN(G9) );
NOR2_X1 U662 ( .A1(n912), .A2(n913), .ZN(G75) );
NOR4_X1 U663 ( .A1(G953), .A2(n914), .A3(n915), .A4(n916), .ZN(n913) );
NOR2_X1 U664 ( .A1(n917), .A2(n918), .ZN(n915) );
NOR2_X1 U665 ( .A1(n919), .A2(n920), .ZN(n917) );
NOR2_X1 U666 ( .A1(n921), .A2(n922), .ZN(n920) );
NOR2_X1 U667 ( .A1(n923), .A2(n924), .ZN(n921) );
NOR2_X1 U668 ( .A1(n925), .A2(n926), .ZN(n924) );
NOR2_X1 U669 ( .A1(n927), .A2(n928), .ZN(n925) );
NOR2_X1 U670 ( .A1(n929), .A2(n930), .ZN(n928) );
XNOR2_X1 U671 ( .A(n931), .B(n932), .ZN(n929) );
NOR3_X1 U672 ( .A1(n933), .A2(KEYINPUT60), .A3(n934), .ZN(n927) );
NOR3_X1 U673 ( .A1(n930), .A2(n935), .A3(n936), .ZN(n923) );
NOR3_X1 U674 ( .A1(n926), .A2(n937), .A3(n936), .ZN(n919) );
NOR3_X1 U675 ( .A1(n938), .A2(n939), .A3(n940), .ZN(n937) );
NOR2_X1 U676 ( .A1(n941), .A2(n942), .ZN(n940) );
XNOR2_X1 U677 ( .A(KEYINPUT15), .B(n930), .ZN(n942) );
NOR3_X1 U678 ( .A1(n943), .A2(n944), .A3(n930), .ZN(n939) );
XNOR2_X1 U679 ( .A(KEYINPUT42), .B(n945), .ZN(n943) );
NOR2_X1 U680 ( .A1(n946), .A2(n922), .ZN(n938) );
NOR2_X1 U681 ( .A1(n947), .A2(n948), .ZN(n946) );
NOR2_X1 U682 ( .A1(n949), .A2(n950), .ZN(n948) );
AND2_X1 U683 ( .A1(n951), .A2(KEYINPUT60), .ZN(n947) );
NOR3_X1 U684 ( .A1(n914), .A2(G953), .A3(G952), .ZN(n912) );
AND4_X1 U685 ( .A1(n952), .A2(n945), .A3(n953), .A4(n954), .ZN(n914) );
NOR4_X1 U686 ( .A1(n955), .A2(n956), .A3(n957), .A4(n958), .ZN(n954) );
XOR2_X1 U687 ( .A(n959), .B(KEYINPUT11), .Z(n957) );
NAND2_X1 U688 ( .A1(n960), .A2(n961), .ZN(n959) );
XOR2_X1 U689 ( .A(n962), .B(KEYINPUT4), .Z(n960) );
XNOR2_X1 U690 ( .A(n932), .B(KEYINPUT3), .ZN(n956) );
INV_X1 U691 ( .A(n944), .ZN(n955) );
XOR2_X1 U692 ( .A(n963), .B(n964), .Z(G72) );
NOR2_X1 U693 ( .A1(n965), .A2(n966), .ZN(n964) );
AND2_X1 U694 ( .A1(G227), .A2(G900), .ZN(n965) );
NAND2_X1 U695 ( .A1(n967), .A2(n968), .ZN(n963) );
NAND2_X1 U696 ( .A1(n969), .A2(n966), .ZN(n968) );
XNOR2_X1 U697 ( .A(n970), .B(n971), .ZN(n969) );
OR3_X1 U698 ( .A1(n972), .A2(n971), .A3(n966), .ZN(n967) );
XNOR2_X1 U699 ( .A(n973), .B(n974), .ZN(n971) );
XOR2_X1 U700 ( .A(n975), .B(n976), .Z(n974) );
NAND2_X1 U701 ( .A1(KEYINPUT54), .A2(n977), .ZN(n975) );
XOR2_X1 U702 ( .A(n978), .B(n979), .Z(G69) );
XOR2_X1 U703 ( .A(n980), .B(n981), .Z(n979) );
NAND2_X1 U704 ( .A1(n966), .A2(n982), .ZN(n981) );
NAND2_X1 U705 ( .A1(n983), .A2(n984), .ZN(n980) );
NAND2_X1 U706 ( .A1(G953), .A2(n985), .ZN(n984) );
NOR2_X1 U707 ( .A1(n986), .A2(n966), .ZN(n978) );
NOR2_X1 U708 ( .A1(n987), .A2(n988), .ZN(n986) );
NOR2_X1 U709 ( .A1(n989), .A2(n990), .ZN(G66) );
XOR2_X1 U710 ( .A(n991), .B(n992), .Z(n990) );
NAND2_X1 U711 ( .A1(n993), .A2(G217), .ZN(n991) );
NOR2_X1 U712 ( .A1(n989), .A2(n994), .ZN(G63) );
XNOR2_X1 U713 ( .A(n995), .B(n996), .ZN(n994) );
NAND2_X1 U714 ( .A1(n993), .A2(G478), .ZN(n995) );
NOR3_X1 U715 ( .A1(n997), .A2(n998), .A3(n999), .ZN(G60) );
AND2_X1 U716 ( .A1(KEYINPUT36), .A2(n989), .ZN(n999) );
NOR3_X1 U717 ( .A1(KEYINPUT36), .A2(G953), .A3(G952), .ZN(n998) );
XOR2_X1 U718 ( .A(n1000), .B(n1001), .Z(n997) );
NAND2_X1 U719 ( .A1(n993), .A2(G475), .ZN(n1000) );
NOR2_X1 U720 ( .A1(n1002), .A2(n1003), .ZN(n993) );
XNOR2_X1 U721 ( .A(n1004), .B(n1005), .ZN(G6) );
NOR2_X1 U722 ( .A1(n989), .A2(n1006), .ZN(G57) );
XOR2_X1 U723 ( .A(n1007), .B(n1008), .Z(n1006) );
XOR2_X1 U724 ( .A(n1009), .B(n1010), .Z(n1008) );
XOR2_X1 U725 ( .A(KEYINPUT1), .B(n1011), .Z(n1010) );
NOR3_X1 U726 ( .A1(n1012), .A2(n1013), .A3(n1002), .ZN(n1011) );
XNOR2_X1 U727 ( .A(KEYINPUT41), .B(n916), .ZN(n1012) );
XOR2_X1 U728 ( .A(KEYINPUT49), .B(KEYINPUT35), .Z(n1009) );
XOR2_X1 U729 ( .A(n1014), .B(n1015), .Z(n1007) );
XNOR2_X1 U730 ( .A(n1016), .B(n1017), .ZN(n1015) );
XNOR2_X1 U731 ( .A(n1018), .B(n1019), .ZN(n1014) );
NOR2_X1 U732 ( .A1(n989), .A2(n1020), .ZN(G54) );
XOR2_X1 U733 ( .A(n1021), .B(n1022), .Z(n1020) );
XOR2_X1 U734 ( .A(n1023), .B(n1024), .Z(n1022) );
NAND2_X1 U735 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NAND2_X1 U736 ( .A1(n1018), .A2(n1027), .ZN(n1026) );
XOR2_X1 U737 ( .A(KEYINPUT29), .B(n1028), .Z(n1025) );
NOR2_X1 U738 ( .A1(n1018), .A2(n1027), .ZN(n1028) );
NAND3_X1 U739 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1027) );
NAND2_X1 U740 ( .A1(KEYINPUT40), .A2(n1032), .ZN(n1031) );
OR3_X1 U741 ( .A1(n1032), .A2(KEYINPUT40), .A3(n976), .ZN(n1030) );
NAND2_X1 U742 ( .A1(n976), .A2(n1033), .ZN(n1029) );
NAND2_X1 U743 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
INV_X1 U744 ( .A(KEYINPUT40), .ZN(n1035) );
XNOR2_X1 U745 ( .A(KEYINPUT34), .B(n1032), .ZN(n1034) );
XOR2_X1 U746 ( .A(n1036), .B(KEYINPUT14), .Z(n1021) );
NAND3_X1 U747 ( .A1(G902), .A2(n1037), .A3(G469), .ZN(n1036) );
XNOR2_X1 U748 ( .A(KEYINPUT37), .B(n916), .ZN(n1037) );
NOR2_X1 U749 ( .A1(n989), .A2(n1038), .ZN(G51) );
XOR2_X1 U750 ( .A(n1039), .B(n1040), .Z(n1038) );
NAND4_X1 U751 ( .A1(n1041), .A2(G210), .A3(n916), .A4(n1042), .ZN(n1040) );
INV_X1 U752 ( .A(n1003), .ZN(n916) );
NOR2_X1 U753 ( .A1(n970), .A2(n982), .ZN(n1003) );
NAND4_X1 U754 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n982) );
AND3_X1 U755 ( .A1(n1047), .A2(n911), .A3(n1048), .ZN(n1046) );
NAND2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n911) );
NAND2_X1 U757 ( .A1(n1005), .A2(n1051), .ZN(n1045) );
INV_X1 U758 ( .A(KEYINPUT28), .ZN(n1051) );
AND2_X1 U759 ( .A1(n1052), .A2(n1050), .ZN(n1005) );
NOR4_X1 U760 ( .A1(n936), .A2(n933), .A3(n941), .A4(n1053), .ZN(n1050) );
NAND2_X1 U761 ( .A1(n951), .A2(n1054), .ZN(n1043) );
NAND3_X1 U762 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
XNOR2_X1 U763 ( .A(KEYINPUT39), .B(n1058), .ZN(n1057) );
NAND3_X1 U764 ( .A1(n1059), .A2(n1060), .A3(n934), .ZN(n1055) );
NAND2_X1 U765 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND3_X1 U766 ( .A1(n941), .A2(n1052), .A3(KEYINPUT28), .ZN(n1062) );
INV_X1 U767 ( .A(n1063), .ZN(n941) );
OR3_X1 U768 ( .A1(n922), .A2(n1064), .A3(n1065), .ZN(n1061) );
NAND4_X1 U769 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n970) );
NOR4_X1 U770 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
NAND2_X1 U771 ( .A1(n1074), .A2(n951), .ZN(n1068) );
OR3_X1 U772 ( .A1(n930), .A2(n935), .A3(n1075), .ZN(n1066) );
NOR2_X1 U773 ( .A1(n1052), .A2(n1049), .ZN(n935) );
XNOR2_X1 U774 ( .A(G902), .B(KEYINPUT27), .ZN(n1041) );
NAND2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1039) );
NAND2_X1 U776 ( .A1(n1078), .A2(n983), .ZN(n1077) );
XOR2_X1 U777 ( .A(n1079), .B(KEYINPUT21), .Z(n1076) );
NAND2_X1 U778 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U779 ( .A(n1078), .B(KEYINPUT6), .Z(n1080) );
XNOR2_X1 U780 ( .A(n1082), .B(KEYINPUT33), .ZN(n1078) );
NOR2_X1 U781 ( .A1(n966), .A2(G952), .ZN(n989) );
XNOR2_X1 U782 ( .A(G146), .B(n1067), .ZN(G48) );
NAND3_X1 U783 ( .A1(n1052), .A2(n951), .A3(n1083), .ZN(n1067) );
XOR2_X1 U784 ( .A(G143), .B(n1073), .Z(G45) );
NOR4_X1 U785 ( .A1(n1065), .A2(n1075), .A3(n933), .A4(n1064), .ZN(n1073) );
XOR2_X1 U786 ( .A(G140), .B(n1072), .Z(G42) );
AND3_X1 U787 ( .A1(n953), .A2(n1063), .A3(n1084), .ZN(n1072) );
XOR2_X1 U788 ( .A(G137), .B(n1071), .Z(G39) );
AND3_X1 U789 ( .A1(n1085), .A2(n953), .A3(n1083), .ZN(n1071) );
XOR2_X1 U790 ( .A(n1086), .B(n1087), .Z(G36) );
NOR4_X1 U791 ( .A1(KEYINPUT0), .A2(n1088), .A3(n930), .A4(n1075), .ZN(n1087) );
XNOR2_X1 U792 ( .A(G134), .B(KEYINPUT63), .ZN(n1086) );
XOR2_X1 U793 ( .A(G131), .B(n1089), .Z(G33) );
NOR3_X1 U794 ( .A1(n1075), .A2(n1090), .A3(n1091), .ZN(n1089) );
INV_X1 U795 ( .A(n1052), .ZN(n1091) );
XNOR2_X1 U796 ( .A(n953), .B(KEYINPUT51), .ZN(n1090) );
INV_X1 U797 ( .A(n930), .ZN(n953) );
NAND2_X1 U798 ( .A1(n1092), .A2(n950), .ZN(n930) );
INV_X1 U799 ( .A(n949), .ZN(n1092) );
NAND4_X1 U800 ( .A1(n1093), .A2(n931), .A3(n1063), .A4(n1094), .ZN(n1075) );
XOR2_X1 U801 ( .A(G128), .B(n1095), .Z(G30) );
NOR2_X1 U802 ( .A1(n933), .A2(n1096), .ZN(n1095) );
XOR2_X1 U803 ( .A(KEYINPUT24), .B(n1074), .Z(n1096) );
AND2_X1 U804 ( .A1(n1083), .A2(n1049), .ZN(n1074) );
AND4_X1 U805 ( .A1(n1093), .A2(n1063), .A3(n1094), .A4(n1097), .ZN(n1083) );
XNOR2_X1 U806 ( .A(G101), .B(n1044), .ZN(G3) );
NAND3_X1 U807 ( .A1(n1085), .A2(n1063), .A3(n1098), .ZN(n1044) );
INV_X1 U808 ( .A(n926), .ZN(n1085) );
XOR2_X1 U809 ( .A(G125), .B(n1070), .Z(G27) );
AND3_X1 U810 ( .A1(n951), .A2(n1099), .A3(n1084), .ZN(n1070) );
AND4_X1 U811 ( .A1(n1052), .A2(n932), .A3(n1094), .A4(n1097), .ZN(n1084) );
NAND2_X1 U812 ( .A1(n918), .A2(n1100), .ZN(n1094) );
NAND4_X1 U813 ( .A1(G953), .A2(G902), .A3(n1101), .A4(n972), .ZN(n1100) );
INV_X1 U814 ( .A(G900), .ZN(n972) );
INV_X1 U815 ( .A(n933), .ZN(n951) );
XOR2_X1 U816 ( .A(n1102), .B(n1103), .Z(G24) );
NAND2_X1 U817 ( .A1(KEYINPUT50), .A2(G122), .ZN(n1103) );
NAND4_X1 U818 ( .A1(n1104), .A2(n1105), .A3(n1099), .A4(n1106), .ZN(n1102) );
NOR3_X1 U819 ( .A1(n1065), .A2(n933), .A3(n936), .ZN(n1106) );
INV_X1 U820 ( .A(n934), .ZN(n936) );
NOR2_X1 U821 ( .A1(n1097), .A2(n1093), .ZN(n934) );
XNOR2_X1 U822 ( .A(KEYINPUT18), .B(n1060), .ZN(n1104) );
XOR2_X1 U823 ( .A(G119), .B(n1107), .Z(G21) );
NOR2_X1 U824 ( .A1(n1108), .A2(n933), .ZN(n1107) );
XOR2_X1 U825 ( .A(n1056), .B(KEYINPUT7), .Z(n1108) );
NAND3_X1 U826 ( .A1(n1093), .A2(n1099), .A3(n1109), .ZN(n1056) );
INV_X1 U827 ( .A(n932), .ZN(n1093) );
XNOR2_X1 U828 ( .A(G116), .B(n1047), .ZN(G18) );
NAND3_X1 U829 ( .A1(n1049), .A2(n1099), .A3(n1098), .ZN(n1047) );
INV_X1 U830 ( .A(n1088), .ZN(n1049) );
NAND2_X1 U831 ( .A1(n952), .A2(n1105), .ZN(n1088) );
XNOR2_X1 U832 ( .A(G113), .B(n1048), .ZN(G15) );
NAND3_X1 U833 ( .A1(n1052), .A2(n1099), .A3(n1098), .ZN(n1048) );
NOR4_X1 U834 ( .A1(n932), .A2(n933), .A3(n1097), .A4(n1053), .ZN(n1098) );
NOR2_X1 U835 ( .A1(n1105), .A2(n1065), .ZN(n1052) );
XNOR2_X1 U836 ( .A(n952), .B(KEYINPUT9), .ZN(n1065) );
XOR2_X1 U837 ( .A(n1110), .B(n1111), .Z(G12) );
NOR3_X1 U838 ( .A1(n1058), .A2(KEYINPUT12), .A3(n933), .ZN(n1111) );
NAND2_X1 U839 ( .A1(n949), .A2(n950), .ZN(n933) );
NAND2_X1 U840 ( .A1(G214), .A2(n1112), .ZN(n950) );
XNOR2_X1 U841 ( .A(KEYINPUT57), .B(n1042), .ZN(n1112) );
INV_X1 U842 ( .A(n1113), .ZN(n1042) );
XNOR2_X1 U843 ( .A(n1114), .B(n1115), .ZN(n949) );
NOR2_X1 U844 ( .A1(n1113), .A2(n1116), .ZN(n1115) );
XOR2_X1 U845 ( .A(KEYINPUT52), .B(G210), .Z(n1116) );
NOR2_X1 U846 ( .A1(G237), .A2(G902), .ZN(n1113) );
NAND2_X1 U847 ( .A1(n1117), .A2(n1002), .ZN(n1114) );
XNOR2_X1 U848 ( .A(n983), .B(n1082), .ZN(n1117) );
XNOR2_X1 U849 ( .A(n1118), .B(n1019), .ZN(n1082) );
XNOR2_X1 U850 ( .A(G125), .B(n1119), .ZN(n1118) );
NOR2_X1 U851 ( .A1(G953), .A2(n988), .ZN(n1119) );
INV_X1 U852 ( .A(G224), .ZN(n988) );
INV_X1 U853 ( .A(n1081), .ZN(n983) );
XNOR2_X1 U854 ( .A(n1120), .B(n1121), .ZN(n1081) );
XOR2_X1 U855 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U856 ( .A(G104), .B(n1124), .ZN(n1123) );
NOR2_X1 U857 ( .A1(G110), .A2(KEYINPUT17), .ZN(n1124) );
XOR2_X1 U858 ( .A(n1125), .B(n1126), .Z(n1120) );
NAND2_X1 U859 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NAND3_X1 U860 ( .A1(G113), .A2(n1129), .A3(n1130), .ZN(n1128) );
OR2_X1 U861 ( .A1(n1130), .A2(n1016), .ZN(n1127) );
INV_X1 U862 ( .A(KEYINPUT25), .ZN(n1130) );
NAND3_X1 U863 ( .A1(n1063), .A2(n932), .A3(n1109), .ZN(n1058) );
NOR3_X1 U864 ( .A1(n931), .A2(n1053), .A3(n926), .ZN(n1109) );
NAND2_X1 U865 ( .A1(n1064), .A2(n952), .ZN(n926) );
XOR2_X1 U866 ( .A(n1131), .B(G475), .Z(n952) );
NAND2_X1 U867 ( .A1(n1001), .A2(n1002), .ZN(n1131) );
XOR2_X1 U868 ( .A(n1132), .B(n1133), .Z(n1001) );
XOR2_X1 U869 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND2_X1 U870 ( .A1(KEYINPUT20), .A2(n1136), .ZN(n1135) );
NAND2_X1 U871 ( .A1(G214), .A2(n1137), .ZN(n1134) );
XOR2_X1 U872 ( .A(n1138), .B(n1139), .Z(n1132) );
XOR2_X1 U873 ( .A(G143), .B(G131), .Z(n1139) );
NAND3_X1 U874 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1138) );
OR2_X1 U875 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND3_X1 U876 ( .A1(n1144), .A2(n1143), .A3(G104), .ZN(n1141) );
NAND2_X1 U877 ( .A1(n1145), .A2(n1004), .ZN(n1140) );
INV_X1 U878 ( .A(G104), .ZN(n1004) );
NAND2_X1 U879 ( .A1(n1146), .A2(n1143), .ZN(n1145) );
INV_X1 U880 ( .A(KEYINPUT53), .ZN(n1143) );
XNOR2_X1 U881 ( .A(n1144), .B(KEYINPUT10), .ZN(n1146) );
XOR2_X1 U882 ( .A(G113), .B(n1126), .Z(n1144) );
INV_X1 U883 ( .A(n1105), .ZN(n1064) );
XOR2_X1 U884 ( .A(n958), .B(KEYINPUT46), .Z(n1105) );
XNOR2_X1 U885 ( .A(n1147), .B(G478), .ZN(n958) );
NAND2_X1 U886 ( .A1(n1148), .A2(n1002), .ZN(n1147) );
XNOR2_X1 U887 ( .A(KEYINPUT43), .B(n1149), .ZN(n1148) );
INV_X1 U888 ( .A(n996), .ZN(n1149) );
XNOR2_X1 U889 ( .A(n1150), .B(n1151), .ZN(n996) );
XOR2_X1 U890 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U891 ( .A(G116), .B(G107), .Z(n1153) );
XOR2_X1 U892 ( .A(KEYINPUT30), .B(G134), .Z(n1152) );
XOR2_X1 U893 ( .A(n1154), .B(n1126), .Z(n1150) );
XOR2_X1 U894 ( .A(G122), .B(KEYINPUT19), .Z(n1126) );
XOR2_X1 U895 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U896 ( .A1(G217), .A2(n1157), .ZN(n1155) );
INV_X1 U897 ( .A(n1060), .ZN(n1053) );
NAND2_X1 U898 ( .A1(n1158), .A2(n918), .ZN(n1060) );
NAND3_X1 U899 ( .A1(n1101), .A2(n966), .A3(G952), .ZN(n918) );
NAND4_X1 U900 ( .A1(G953), .A2(G902), .A3(n985), .A4(n1101), .ZN(n1158) );
NAND2_X1 U901 ( .A1(G237), .A2(n1159), .ZN(n1101) );
XNOR2_X1 U902 ( .A(KEYINPUT61), .B(n987), .ZN(n985) );
INV_X1 U903 ( .A(G898), .ZN(n987) );
INV_X1 U904 ( .A(n1097), .ZN(n931) );
NAND2_X1 U905 ( .A1(n961), .A2(n962), .ZN(n1097) );
NAND2_X1 U906 ( .A1(G217), .A2(n1160), .ZN(n962) );
NAND2_X1 U907 ( .A1(n1161), .A2(n1002), .ZN(n1160) );
NAND2_X1 U908 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U909 ( .A(KEYINPUT56), .B(n992), .Z(n1163) );
NAND3_X1 U910 ( .A1(n1164), .A2(n1002), .A3(n1165), .ZN(n961) );
XNOR2_X1 U911 ( .A(n992), .B(KEYINPUT56), .ZN(n1165) );
XNOR2_X1 U912 ( .A(n1166), .B(n1167), .ZN(n992) );
XOR2_X1 U913 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U914 ( .A(G128), .B(G119), .Z(n1169) );
XOR2_X1 U915 ( .A(KEYINPUT8), .B(G137), .Z(n1168) );
XNOR2_X1 U916 ( .A(n1170), .B(n1136), .ZN(n1166) );
XOR2_X1 U917 ( .A(n973), .B(n1171), .Z(n1136) );
XNOR2_X1 U918 ( .A(G125), .B(G140), .ZN(n973) );
XOR2_X1 U919 ( .A(n1172), .B(G110), .Z(n1170) );
NAND2_X1 U920 ( .A1(G221), .A2(n1157), .ZN(n1172) );
AND2_X1 U921 ( .A1(G234), .A2(n966), .ZN(n1157) );
NAND2_X1 U922 ( .A1(n1162), .A2(G217), .ZN(n1164) );
INV_X1 U923 ( .A(n1159), .ZN(n1162) );
XNOR2_X1 U924 ( .A(n1173), .B(n1174), .ZN(n932) );
XNOR2_X1 U925 ( .A(KEYINPUT22), .B(n1013), .ZN(n1174) );
INV_X1 U926 ( .A(G472), .ZN(n1013) );
NAND2_X1 U927 ( .A1(n1175), .A2(n1002), .ZN(n1173) );
XOR2_X1 U928 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U929 ( .A(n1178), .B(n1019), .ZN(n1177) );
NAND2_X1 U930 ( .A1(KEYINPUT55), .A2(n1018), .ZN(n1178) );
XOR2_X1 U931 ( .A(n1179), .B(n1180), .Z(n1176) );
XOR2_X1 U932 ( .A(KEYINPUT59), .B(n1181), .Z(n1180) );
NOR2_X1 U933 ( .A1(KEYINPUT38), .A2(n1017), .ZN(n1181) );
XNOR2_X1 U934 ( .A(n1182), .B(G101), .ZN(n1017) );
NAND2_X1 U935 ( .A1(G210), .A2(n1137), .ZN(n1182) );
NOR2_X1 U936 ( .A1(G953), .A2(G237), .ZN(n1137) );
NOR2_X1 U937 ( .A1(KEYINPUT31), .A2(n1016), .ZN(n1179) );
XNOR2_X1 U938 ( .A(G113), .B(n1129), .ZN(n1016) );
XOR2_X1 U939 ( .A(G116), .B(G119), .Z(n1129) );
NAND2_X1 U940 ( .A1(n1183), .A2(n1184), .ZN(n1063) );
OR3_X1 U941 ( .A1(n1185), .A2(n945), .A3(KEYINPUT13), .ZN(n1184) );
NAND2_X1 U942 ( .A1(KEYINPUT13), .A2(n1099), .ZN(n1183) );
INV_X1 U943 ( .A(n922), .ZN(n1099) );
NAND2_X1 U944 ( .A1(n945), .A2(n1186), .ZN(n922) );
INV_X1 U945 ( .A(n1185), .ZN(n1186) );
XOR2_X1 U946 ( .A(n944), .B(KEYINPUT44), .Z(n1185) );
NAND2_X1 U947 ( .A1(G221), .A2(n1187), .ZN(n944) );
NAND2_X1 U948 ( .A1(n1159), .A2(n1002), .ZN(n1187) );
XOR2_X1 U949 ( .A(G234), .B(KEYINPUT23), .Z(n1159) );
XOR2_X1 U950 ( .A(n1188), .B(G469), .Z(n945) );
NAND2_X1 U951 ( .A1(n1189), .A2(n1002), .ZN(n1188) );
INV_X1 U952 ( .A(G902), .ZN(n1002) );
XNOR2_X1 U953 ( .A(n1190), .B(n1191), .ZN(n1189) );
XOR2_X1 U954 ( .A(n1192), .B(n1024), .Z(n1191) );
XOR2_X1 U955 ( .A(n1193), .B(n1194), .Z(n1024) );
XOR2_X1 U956 ( .A(G140), .B(G110), .Z(n1194) );
NAND2_X1 U957 ( .A1(G227), .A2(n966), .ZN(n1193) );
INV_X1 U958 ( .A(G953), .ZN(n966) );
NAND2_X1 U959 ( .A1(n1195), .A2(n1196), .ZN(n1192) );
XOR2_X1 U960 ( .A(n976), .B(n1197), .Z(n1196) );
XOR2_X1 U961 ( .A(n1032), .B(KEYINPUT16), .Z(n1197) );
XOR2_X1 U962 ( .A(n1122), .B(n1198), .Z(n1032) );
NOR2_X1 U963 ( .A1(KEYINPUT5), .A2(n1199), .ZN(n1198) );
XNOR2_X1 U964 ( .A(G104), .B(KEYINPUT47), .ZN(n1199) );
XNOR2_X1 U965 ( .A(G101), .B(G107), .ZN(n1122) );
XOR2_X1 U966 ( .A(n1200), .B(n1019), .Z(n976) );
XOR2_X1 U967 ( .A(n1156), .B(n1171), .Z(n1019) );
XOR2_X1 U968 ( .A(G146), .B(KEYINPUT45), .Z(n1171) );
XOR2_X1 U969 ( .A(G128), .B(G143), .Z(n1156) );
XNOR2_X1 U970 ( .A(KEYINPUT26), .B(KEYINPUT2), .ZN(n1200) );
XNOR2_X1 U971 ( .A(KEYINPUT62), .B(KEYINPUT58), .ZN(n1195) );
INV_X1 U972 ( .A(n1018), .ZN(n1190) );
XNOR2_X1 U973 ( .A(n977), .B(KEYINPUT48), .ZN(n1018) );
XNOR2_X1 U974 ( .A(G131), .B(n1201), .ZN(n977) );
XOR2_X1 U975 ( .A(G137), .B(G134), .Z(n1201) );
XNOR2_X1 U976 ( .A(G110), .B(KEYINPUT32), .ZN(n1110) );
endmodule


