//Key = 0100010001111111101010111100100001110001101000011001101000001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359;

XOR2_X1 U745 ( .A(n1035), .B(n1036), .Z(G9) );
NAND4_X1 U746 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(G75) );
INV_X1 U747 ( .A(n1041), .ZN(n1040) );
NAND4_X1 U748 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1039) );
NOR3_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NOR2_X1 U750 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
NAND3_X1 U752 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1046) );
NOR3_X1 U753 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1044) );
XOR2_X1 U754 ( .A(n1059), .B(KEYINPUT22), .Z(n1057) );
NAND2_X1 U755 ( .A1(n1052), .A2(n1051), .ZN(n1059) );
XOR2_X1 U756 ( .A(KEYINPUT62), .B(n1060), .Z(n1052) );
XNOR2_X1 U757 ( .A(n1061), .B(G472), .ZN(n1043) );
XOR2_X1 U758 ( .A(n1062), .B(n1063), .Z(n1042) );
NAND2_X1 U759 ( .A1(G952), .A2(n1064), .ZN(n1038) );
NAND3_X1 U760 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND2_X1 U762 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND4_X1 U763 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1055), .ZN(n1071) );
NAND2_X1 U764 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U765 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U766 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U767 ( .A1(n1081), .A2(n1082), .ZN(n1075) );
NAND2_X1 U768 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
OR2_X1 U769 ( .A1(n1053), .A2(n1085), .ZN(n1084) );
NAND3_X1 U770 ( .A1(n1077), .A2(n1086), .A3(n1081), .ZN(n1070) );
NAND2_X1 U771 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U772 ( .A1(n1089), .A2(n1090), .A3(n1073), .ZN(n1088) );
OR2_X1 U773 ( .A1(n1055), .A2(n1072), .ZN(n1090) );
NAND3_X1 U774 ( .A1(n1091), .A2(n1092), .A3(n1055), .ZN(n1089) );
INV_X1 U775 ( .A(n1093), .ZN(n1092) );
NAND2_X1 U776 ( .A1(n1094), .A2(n1056), .ZN(n1091) );
NAND2_X1 U777 ( .A1(n1072), .A2(n1095), .ZN(n1087) );
INV_X1 U778 ( .A(n1096), .ZN(n1068) );
NAND2_X1 U779 ( .A1(KEYINPUT17), .A2(n1097), .ZN(n1065) );
OR2_X1 U780 ( .A1(n1097), .A2(KEYINPUT17), .ZN(n1037) );
XOR2_X1 U781 ( .A(n1098), .B(n1099), .Z(G72) );
XOR2_X1 U782 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U783 ( .A1(n1102), .A2(n1097), .ZN(n1101) );
NOR2_X1 U784 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
NAND2_X1 U786 ( .A1(G953), .A2(n1104), .ZN(n1106) );
XOR2_X1 U787 ( .A(n1107), .B(n1108), .Z(n1105) );
XNOR2_X1 U788 ( .A(n1109), .B(n1110), .ZN(n1108) );
XOR2_X1 U789 ( .A(n1111), .B(n1112), .Z(n1107) );
NOR2_X1 U790 ( .A1(KEYINPUT21), .A2(n1113), .ZN(n1112) );
XOR2_X1 U791 ( .A(n1114), .B(G137), .Z(n1113) );
INV_X1 U792 ( .A(G134), .ZN(n1114) );
NAND2_X1 U793 ( .A1(n1097), .A2(n1115), .ZN(n1098) );
NAND2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U795 ( .A(n1118), .B(n1119), .Z(G69) );
NOR2_X1 U796 ( .A1(n1120), .A2(G953), .ZN(n1119) );
NAND2_X1 U797 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
NAND2_X1 U798 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
INV_X1 U799 ( .A(n1125), .ZN(n1123) );
NAND2_X1 U800 ( .A1(n1126), .A2(n1125), .ZN(n1121) );
NAND2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1127) );
NOR2_X1 U803 ( .A1(KEYINPUT58), .A2(n1131), .ZN(n1129) );
XOR2_X1 U804 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U805 ( .A1(n1128), .A2(n1124), .ZN(n1126) );
NAND2_X1 U806 ( .A1(G953), .A2(n1134), .ZN(n1124) );
INV_X1 U807 ( .A(n1135), .ZN(n1128) );
NOR2_X1 U808 ( .A1(n1041), .A2(n1136), .ZN(G66) );
XOR2_X1 U809 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U810 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NOR2_X1 U811 ( .A1(n1041), .A2(n1141), .ZN(G63) );
NOR3_X1 U812 ( .A1(n1060), .A2(n1142), .A3(n1143), .ZN(n1141) );
NOR3_X1 U813 ( .A1(n1144), .A2(n1145), .A3(n1140), .ZN(n1143) );
NOR2_X1 U814 ( .A1(n1146), .A2(n1147), .ZN(n1142) );
NOR2_X1 U815 ( .A1(n1067), .A2(n1145), .ZN(n1146) );
INV_X1 U816 ( .A(G478), .ZN(n1145) );
INV_X1 U817 ( .A(n1148), .ZN(n1067) );
NOR2_X1 U818 ( .A1(n1041), .A2(n1149), .ZN(G60) );
XOR2_X1 U819 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR3_X1 U820 ( .A1(n1140), .A2(KEYINPUT59), .A3(n1050), .ZN(n1150) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(G6) );
NOR2_X1 U822 ( .A1(G104), .A2(KEYINPUT50), .ZN(n1153) );
NOR3_X1 U823 ( .A1(n1041), .A2(n1154), .A3(n1155), .ZN(G57) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U825 ( .A(n1158), .B(n1159), .Z(n1156) );
NOR2_X1 U826 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
INV_X1 U827 ( .A(KEYINPUT33), .ZN(n1161) );
NOR2_X1 U828 ( .A1(n1162), .A2(n1163), .ZN(n1154) );
XOR2_X1 U829 ( .A(n1164), .B(n1159), .Z(n1163) );
XNOR2_X1 U830 ( .A(n1165), .B(n1166), .ZN(n1159) );
XOR2_X1 U831 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND3_X1 U832 ( .A1(G472), .A2(n1148), .A3(n1169), .ZN(n1168) );
XOR2_X1 U833 ( .A(n1170), .B(KEYINPUT51), .Z(n1169) );
NAND2_X1 U834 ( .A1(KEYINPUT16), .A2(n1171), .ZN(n1165) );
AND2_X1 U835 ( .A1(n1160), .A2(KEYINPUT33), .ZN(n1164) );
XOR2_X1 U836 ( .A(n1172), .B(n1173), .Z(n1160) );
XNOR2_X1 U837 ( .A(KEYINPUT6), .B(n1174), .ZN(n1172) );
NOR2_X1 U838 ( .A1(KEYINPUT38), .A2(n1175), .ZN(n1174) );
INV_X1 U839 ( .A(n1157), .ZN(n1162) );
NOR2_X1 U840 ( .A1(n1041), .A2(n1176), .ZN(G54) );
XOR2_X1 U841 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U842 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U843 ( .A1(G140), .A2(KEYINPUT29), .ZN(n1180) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1140), .ZN(n1179) );
XOR2_X1 U845 ( .A(n1182), .B(n1183), .Z(n1177) );
NOR2_X1 U846 ( .A1(KEYINPUT2), .A2(n1184), .ZN(n1183) );
XOR2_X1 U847 ( .A(n1109), .B(n1185), .Z(n1184) );
XNOR2_X1 U848 ( .A(n1186), .B(n1187), .ZN(n1185) );
NOR2_X1 U849 ( .A1(KEYINPUT36), .A2(n1175), .ZN(n1187) );
NAND2_X1 U850 ( .A1(KEYINPUT48), .A2(n1188), .ZN(n1186) );
XOR2_X1 U851 ( .A(n1189), .B(n1190), .Z(n1182) );
NOR2_X1 U852 ( .A1(n1041), .A2(n1191), .ZN(G51) );
XOR2_X1 U853 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U854 ( .A(n1194), .B(n1195), .Z(n1192) );
NOR2_X1 U855 ( .A1(n1196), .A2(n1140), .ZN(n1195) );
NAND2_X1 U856 ( .A1(G902), .A2(n1148), .ZN(n1140) );
NAND3_X1 U857 ( .A1(n1116), .A2(n1197), .A3(n1120), .ZN(n1148) );
AND4_X1 U858 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1120) );
AND4_X1 U859 ( .A1(n1202), .A2(n1203), .A3(n1152), .A4(n1204), .ZN(n1201) );
NAND4_X1 U860 ( .A1(n1095), .A2(n1205), .A3(n1077), .A4(n1206), .ZN(n1204) );
NAND3_X1 U861 ( .A1(n1207), .A2(n1072), .A3(n1208), .ZN(n1152) );
NOR2_X1 U862 ( .A1(n1209), .A2(n1210), .ZN(n1200) );
INV_X1 U863 ( .A(n1036), .ZN(n1210) );
NAND3_X1 U864 ( .A1(n1205), .A2(n1072), .A3(n1207), .ZN(n1036) );
XNOR2_X1 U865 ( .A(KEYINPUT39), .B(n1117), .ZN(n1197) );
AND4_X1 U866 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1116) );
NOR4_X1 U867 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NAND2_X1 U868 ( .A1(n1219), .A2(n1220), .ZN(n1213) );
NOR2_X1 U869 ( .A1(n1097), .A2(G952), .ZN(n1041) );
XOR2_X1 U870 ( .A(n1221), .B(n1211), .Z(G48) );
NAND2_X1 U871 ( .A1(n1222), .A2(n1208), .ZN(n1211) );
XOR2_X1 U872 ( .A(n1223), .B(n1224), .Z(G45) );
XOR2_X1 U873 ( .A(KEYINPUT12), .B(G143), .Z(n1224) );
NAND2_X1 U874 ( .A1(n1225), .A2(n1219), .ZN(n1223) );
AND3_X1 U875 ( .A1(n1093), .A2(n1226), .A3(n1227), .ZN(n1219) );
XOR2_X1 U876 ( .A(n1083), .B(KEYINPUT47), .Z(n1225) );
XNOR2_X1 U877 ( .A(G140), .B(n1212), .ZN(G42) );
NAND4_X1 U878 ( .A1(n1228), .A2(n1208), .A3(n1094), .A4(n1056), .ZN(n1212) );
XOR2_X1 U879 ( .A(G137), .B(n1218), .Z(G39) );
AND4_X1 U880 ( .A1(n1228), .A2(n1081), .A3(n1056), .A4(n1229), .ZN(n1218) );
XOR2_X1 U881 ( .A(G134), .B(n1217), .Z(G36) );
AND3_X1 U882 ( .A1(n1093), .A2(n1205), .A3(n1228), .ZN(n1217) );
XOR2_X1 U883 ( .A(G131), .B(n1216), .Z(G33) );
AND3_X1 U884 ( .A1(n1208), .A2(n1093), .A3(n1228), .ZN(n1216) );
AND4_X1 U885 ( .A1(n1220), .A2(n1073), .A3(n1226), .A4(n1055), .ZN(n1228) );
XOR2_X1 U886 ( .A(n1230), .B(n1117), .Z(G30) );
NAND2_X1 U887 ( .A1(n1222), .A2(n1205), .ZN(n1117) );
AND3_X1 U888 ( .A1(n1220), .A2(n1229), .A3(n1231), .ZN(n1222) );
XOR2_X1 U889 ( .A(n1203), .B(n1232), .Z(G3) );
XOR2_X1 U890 ( .A(n1171), .B(KEYINPUT0), .Z(n1232) );
NAND3_X1 U891 ( .A1(n1081), .A2(n1207), .A3(n1093), .ZN(n1203) );
XOR2_X1 U892 ( .A(G125), .B(n1215), .Z(G27) );
AND4_X1 U893 ( .A1(n1231), .A2(n1208), .A3(n1094), .A4(n1077), .ZN(n1215) );
AND3_X1 U894 ( .A1(n1056), .A2(n1226), .A3(n1095), .ZN(n1231) );
NAND2_X1 U895 ( .A1(n1233), .A2(n1096), .ZN(n1226) );
XOR2_X1 U896 ( .A(n1234), .B(KEYINPUT57), .Z(n1233) );
NAND4_X1 U897 ( .A1(G902), .A2(G953), .A3(n1235), .A4(n1104), .ZN(n1234) );
INV_X1 U898 ( .A(G900), .ZN(n1104) );
XOR2_X1 U899 ( .A(n1236), .B(n1202), .Z(G24) );
NAND4_X1 U900 ( .A1(n1227), .A2(n1077), .A3(n1072), .A4(n1237), .ZN(n1202) );
NOR2_X1 U901 ( .A1(n1229), .A2(n1056), .ZN(n1072) );
AND3_X1 U902 ( .A1(n1238), .A2(n1239), .A3(n1095), .ZN(n1227) );
XOR2_X1 U903 ( .A(n1240), .B(n1241), .Z(G21) );
NAND2_X1 U904 ( .A1(KEYINPUT9), .A2(n1209), .ZN(n1241) );
AND4_X1 U905 ( .A1(n1077), .A2(n1095), .A3(n1081), .A4(n1242), .ZN(n1209) );
AND3_X1 U906 ( .A1(n1056), .A2(n1237), .A3(n1229), .ZN(n1242) );
INV_X1 U907 ( .A(n1094), .ZN(n1229) );
XOR2_X1 U908 ( .A(G116), .B(n1243), .Z(G18) );
NOR4_X1 U909 ( .A1(n1244), .A2(n1080), .A3(n1245), .A4(n1246), .ZN(n1243) );
XOR2_X1 U910 ( .A(KEYINPUT63), .B(n1095), .Z(n1246) );
INV_X1 U911 ( .A(n1205), .ZN(n1080) );
NOR2_X1 U912 ( .A1(n1239), .A2(n1247), .ZN(n1205) );
XNOR2_X1 U913 ( .A(n1077), .B(KEYINPUT46), .ZN(n1244) );
XOR2_X1 U914 ( .A(n1132), .B(n1198), .Z(G15) );
NAND4_X1 U915 ( .A1(n1208), .A2(n1206), .A3(n1077), .A4(n1248), .ZN(n1198) );
NOR2_X1 U916 ( .A1(n1085), .A2(n1249), .ZN(n1077) );
INV_X1 U917 ( .A(n1053), .ZN(n1249) );
INV_X1 U918 ( .A(n1245), .ZN(n1206) );
NAND2_X1 U919 ( .A1(n1093), .A2(n1237), .ZN(n1245) );
NOR2_X1 U920 ( .A1(n1056), .A2(n1094), .ZN(n1093) );
INV_X1 U921 ( .A(n1079), .ZN(n1208) );
NAND2_X1 U922 ( .A1(n1247), .A2(n1239), .ZN(n1079) );
NAND2_X1 U923 ( .A1(n1250), .A2(n1251), .ZN(G12) );
NAND2_X1 U924 ( .A1(n1252), .A2(n1189), .ZN(n1251) );
XOR2_X1 U925 ( .A(KEYINPUT60), .B(n1253), .Z(n1250) );
NOR2_X1 U926 ( .A1(n1252), .A2(n1189), .ZN(n1253) );
INV_X1 U927 ( .A(n1199), .ZN(n1252) );
NAND4_X1 U928 ( .A1(n1081), .A2(n1207), .A3(n1094), .A4(n1056), .ZN(n1199) );
XOR2_X1 U929 ( .A(n1254), .B(n1139), .Z(n1056) );
NAND2_X1 U930 ( .A1(G217), .A2(n1255), .ZN(n1139) );
OR2_X1 U931 ( .A1(n1138), .A2(G902), .ZN(n1254) );
XNOR2_X1 U932 ( .A(n1256), .B(n1257), .ZN(n1138) );
XOR2_X1 U933 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U934 ( .A(n1260), .B(n1261), .Z(n1259) );
AND3_X1 U935 ( .A1(G221), .A2(n1097), .A3(G234), .ZN(n1261) );
NAND2_X1 U936 ( .A1(KEYINPUT35), .A2(n1262), .ZN(n1260) );
XOR2_X1 U937 ( .A(n1111), .B(n1263), .Z(n1262) );
NAND2_X1 U938 ( .A1(KEYINPUT25), .A2(G140), .ZN(n1263) );
INV_X1 U939 ( .A(G125), .ZN(n1111) );
NAND2_X1 U940 ( .A1(KEYINPUT24), .A2(n1240), .ZN(n1258) );
INV_X1 U941 ( .A(G119), .ZN(n1240) );
XOR2_X1 U942 ( .A(n1264), .B(n1265), .Z(n1256) );
XOR2_X1 U943 ( .A(G146), .B(G137), .Z(n1265) );
XOR2_X1 U944 ( .A(n1230), .B(G110), .Z(n1264) );
INV_X1 U945 ( .A(G128), .ZN(n1230) );
XOR2_X1 U946 ( .A(n1266), .B(G472), .Z(n1094) );
NAND2_X1 U947 ( .A1(KEYINPUT54), .A2(n1061), .ZN(n1266) );
AND3_X1 U948 ( .A1(n1267), .A2(n1268), .A3(n1170), .ZN(n1061) );
OR2_X1 U949 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND2_X1 U950 ( .A1(n1271), .A2(n1270), .ZN(n1267) );
XNOR2_X1 U951 ( .A(n1167), .B(G101), .ZN(n1270) );
NAND2_X1 U952 ( .A1(n1272), .A2(G210), .ZN(n1167) );
XOR2_X1 U953 ( .A(KEYINPUT4), .B(n1269), .Z(n1271) );
XNOR2_X1 U954 ( .A(n1273), .B(n1274), .ZN(n1269) );
XOR2_X1 U955 ( .A(n1157), .B(n1173), .Z(n1274) );
XOR2_X1 U956 ( .A(n1275), .B(n1276), .Z(n1157) );
NOR2_X1 U957 ( .A1(KEYINPUT37), .A2(n1133), .ZN(n1276) );
XOR2_X1 U958 ( .A(n1132), .B(KEYINPUT23), .Z(n1275) );
XNOR2_X1 U959 ( .A(n1175), .B(KEYINPUT45), .ZN(n1273) );
AND3_X1 U960 ( .A1(n1248), .A2(n1237), .A3(n1220), .ZN(n1207) );
INV_X1 U961 ( .A(n1083), .ZN(n1220) );
NAND2_X1 U962 ( .A1(n1085), .A2(n1053), .ZN(n1083) );
NAND2_X1 U963 ( .A1(G221), .A2(n1255), .ZN(n1053) );
NAND2_X1 U964 ( .A1(G234), .A2(n1170), .ZN(n1255) );
XOR2_X1 U965 ( .A(n1058), .B(KEYINPUT3), .Z(n1085) );
XNOR2_X1 U966 ( .A(n1181), .B(n1277), .ZN(n1058) );
NOR2_X1 U967 ( .A1(G902), .A2(n1278), .ZN(n1277) );
XOR2_X1 U968 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U969 ( .A(n1190), .B(n1281), .Z(n1280) );
NOR3_X1 U970 ( .A1(n1282), .A2(KEYINPUT26), .A3(n1283), .ZN(n1281) );
NOR2_X1 U971 ( .A1(n1284), .A2(n1175), .ZN(n1283) );
XOR2_X1 U972 ( .A(n1285), .B(KEYINPUT34), .Z(n1282) );
NAND2_X1 U973 ( .A1(n1284), .A2(n1175), .ZN(n1285) );
XNOR2_X1 U974 ( .A(n1286), .B(n1287), .ZN(n1175) );
XOR2_X1 U975 ( .A(G134), .B(G131), .Z(n1287) );
NAND2_X1 U976 ( .A1(KEYINPUT52), .A2(n1288), .ZN(n1286) );
XOR2_X1 U977 ( .A(KEYINPUT42), .B(G137), .Z(n1288) );
XOR2_X1 U978 ( .A(n1188), .B(n1289), .Z(n1284) );
NOR2_X1 U979 ( .A1(KEYINPUT19), .A2(n1109), .ZN(n1289) );
XNOR2_X1 U980 ( .A(n1290), .B(G128), .ZN(n1109) );
NAND3_X1 U981 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1290) );
NAND2_X1 U982 ( .A1(KEYINPUT53), .A2(G143), .ZN(n1293) );
NAND3_X1 U983 ( .A1(n1294), .A2(n1295), .A3(G146), .ZN(n1292) );
INV_X1 U984 ( .A(G143), .ZN(n1294) );
NAND2_X1 U985 ( .A1(n1296), .A2(n1221), .ZN(n1291) );
INV_X1 U986 ( .A(G146), .ZN(n1221) );
NAND2_X1 U987 ( .A1(n1297), .A2(n1295), .ZN(n1296) );
INV_X1 U988 ( .A(KEYINPUT53), .ZN(n1295) );
XOR2_X1 U989 ( .A(KEYINPUT18), .B(G143), .Z(n1297) );
NAND3_X1 U990 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1188) );
NAND2_X1 U991 ( .A1(n1301), .A2(n1171), .ZN(n1300) );
INV_X1 U992 ( .A(G101), .ZN(n1171) );
NAND2_X1 U993 ( .A1(n1302), .A2(n1303), .ZN(n1299) );
INV_X1 U994 ( .A(KEYINPUT5), .ZN(n1303) );
NAND2_X1 U995 ( .A1(G101), .A2(n1304), .ZN(n1302) );
XOR2_X1 U996 ( .A(KEYINPUT28), .B(n1301), .Z(n1304) );
INV_X1 U997 ( .A(n1305), .ZN(n1301) );
NAND2_X1 U998 ( .A1(KEYINPUT5), .A2(n1306), .ZN(n1298) );
NAND2_X1 U999 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
OR2_X1 U1000 ( .A1(n1305), .A2(KEYINPUT28), .ZN(n1308) );
NAND3_X1 U1001 ( .A1(G101), .A2(n1305), .A3(KEYINPUT28), .ZN(n1307) );
XOR2_X1 U1002 ( .A(n1309), .B(G107), .Z(n1305) );
NAND2_X1 U1003 ( .A1(KEYINPUT13), .A2(n1310), .ZN(n1309) );
INV_X1 U1004 ( .A(G104), .ZN(n1310) );
NOR2_X1 U1005 ( .A1(n1103), .A2(G953), .ZN(n1190) );
INV_X1 U1006 ( .A(G227), .ZN(n1103) );
NAND2_X1 U1007 ( .A1(n1311), .A2(KEYINPUT40), .ZN(n1279) );
XOR2_X1 U1008 ( .A(n1189), .B(n1312), .Z(n1311) );
XOR2_X1 U1009 ( .A(KEYINPUT11), .B(G140), .Z(n1312) );
INV_X1 U1010 ( .A(G469), .ZN(n1181) );
NAND2_X1 U1011 ( .A1(n1096), .A2(n1313), .ZN(n1237) );
NAND3_X1 U1012 ( .A1(n1135), .A2(n1235), .A3(G902), .ZN(n1313) );
NOR2_X1 U1013 ( .A1(G898), .A2(n1097), .ZN(n1135) );
NAND3_X1 U1014 ( .A1(n1235), .A2(n1097), .A3(G952), .ZN(n1096) );
NAND2_X1 U1015 ( .A1(G237), .A2(G234), .ZN(n1235) );
XOR2_X1 U1016 ( .A(n1095), .B(KEYINPUT7), .Z(n1248) );
NOR2_X1 U1017 ( .A1(n1073), .A2(n1314), .ZN(n1095) );
INV_X1 U1018 ( .A(n1055), .ZN(n1314) );
NAND2_X1 U1019 ( .A1(G214), .A2(n1315), .ZN(n1055) );
XNOR2_X1 U1020 ( .A(n1062), .B(n1316), .ZN(n1073) );
NOR2_X1 U1021 ( .A1(n1063), .A2(KEYINPUT41), .ZN(n1316) );
INV_X1 U1022 ( .A(n1196), .ZN(n1063) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1315), .ZN(n1196) );
NAND2_X1 U1024 ( .A1(n1317), .A2(n1170), .ZN(n1315) );
XNOR2_X1 U1025 ( .A(G237), .B(KEYINPUT49), .ZN(n1317) );
NAND2_X1 U1026 ( .A1(n1318), .A2(n1170), .ZN(n1062) );
INV_X1 U1027 ( .A(G902), .ZN(n1170) );
XOR2_X1 U1028 ( .A(n1319), .B(n1194), .Z(n1318) );
XNOR2_X1 U1029 ( .A(n1130), .B(n1320), .ZN(n1194) );
NOR2_X1 U1030 ( .A1(KEYINPUT44), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1031 ( .A(n1133), .B(G113), .Z(n1321) );
XNOR2_X1 U1032 ( .A(G116), .B(n1322), .ZN(n1133) );
XOR2_X1 U1033 ( .A(KEYINPUT27), .B(G119), .Z(n1322) );
XNOR2_X1 U1034 ( .A(n1323), .B(n1324), .ZN(n1130) );
XOR2_X1 U1035 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1036 ( .A(G107), .B(G101), .Z(n1326) );
NOR2_X1 U1037 ( .A1(G104), .A2(KEYINPUT56), .ZN(n1325) );
XOR2_X1 U1038 ( .A(n1189), .B(n1327), .Z(n1323) );
XOR2_X1 U1039 ( .A(KEYINPUT14), .B(G122), .Z(n1327) );
INV_X1 U1040 ( .A(G110), .ZN(n1189) );
NAND2_X1 U1041 ( .A1(KEYINPUT1), .A2(n1193), .ZN(n1319) );
XNOR2_X1 U1042 ( .A(n1173), .B(n1328), .ZN(n1193) );
XOR2_X1 U1043 ( .A(G125), .B(n1329), .Z(n1328) );
NOR2_X1 U1044 ( .A1(G953), .A2(n1134), .ZN(n1329) );
INV_X1 U1045 ( .A(G224), .ZN(n1134) );
XNOR2_X1 U1046 ( .A(G128), .B(n1330), .ZN(n1173) );
NOR2_X1 U1047 ( .A1(n1238), .A2(n1239), .ZN(n1081) );
NAND2_X1 U1048 ( .A1(n1331), .A2(n1332), .ZN(n1239) );
OR2_X1 U1049 ( .A1(n1050), .A2(n1049), .ZN(n1332) );
XOR2_X1 U1050 ( .A(n1054), .B(KEYINPUT8), .Z(n1331) );
NAND2_X1 U1051 ( .A1(n1049), .A2(n1050), .ZN(n1054) );
INV_X1 U1052 ( .A(G475), .ZN(n1050) );
NOR2_X1 U1053 ( .A1(n1151), .A2(G902), .ZN(n1049) );
XNOR2_X1 U1054 ( .A(n1333), .B(n1334), .ZN(n1151) );
NOR2_X1 U1055 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NOR2_X1 U1056 ( .A1(G122), .A2(n1337), .ZN(n1336) );
NOR2_X1 U1057 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NOR2_X1 U1058 ( .A1(KEYINPUT31), .A2(G113), .ZN(n1338) );
NOR2_X1 U1059 ( .A1(n1340), .A2(n1132), .ZN(n1335) );
INV_X1 U1060 ( .A(G113), .ZN(n1132) );
NOR2_X1 U1061 ( .A1(n1341), .A2(KEYINPUT31), .ZN(n1340) );
NOR2_X1 U1062 ( .A1(n1236), .A2(n1339), .ZN(n1341) );
INV_X1 U1063 ( .A(KEYINPUT20), .ZN(n1339) );
XOR2_X1 U1064 ( .A(n1342), .B(G104), .Z(n1333) );
NAND2_X1 U1065 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XOR2_X1 U1066 ( .A(n1345), .B(n1346), .Z(n1344) );
XNOR2_X1 U1067 ( .A(n1110), .B(n1330), .ZN(n1346) );
XOR2_X1 U1068 ( .A(G146), .B(G143), .Z(n1330) );
XOR2_X1 U1069 ( .A(G131), .B(G140), .Z(n1110) );
XOR2_X1 U1070 ( .A(n1347), .B(n1348), .Z(n1345) );
NOR2_X1 U1071 ( .A1(KEYINPUT32), .A2(G125), .ZN(n1348) );
NAND2_X1 U1072 ( .A1(n1272), .A2(G214), .ZN(n1347) );
NOR2_X1 U1073 ( .A1(G953), .A2(G237), .ZN(n1272) );
XNOR2_X1 U1074 ( .A(KEYINPUT15), .B(KEYINPUT10), .ZN(n1343) );
INV_X1 U1075 ( .A(n1247), .ZN(n1238) );
XNOR2_X1 U1076 ( .A(n1060), .B(n1051), .ZN(n1247) );
XOR2_X1 U1077 ( .A(G478), .B(KEYINPUT55), .Z(n1051) );
NOR2_X1 U1078 ( .A1(n1147), .A2(G902), .ZN(n1060) );
INV_X1 U1079 ( .A(n1144), .ZN(n1147) );
XOR2_X1 U1080 ( .A(n1349), .B(n1350), .Z(n1144) );
XOR2_X1 U1081 ( .A(n1351), .B(n1352), .Z(n1350) );
XOR2_X1 U1082 ( .A(G134), .B(G128), .Z(n1352) );
XOR2_X1 U1083 ( .A(KEYINPUT61), .B(G143), .Z(n1351) );
XOR2_X1 U1084 ( .A(n1353), .B(n1354), .Z(n1349) );
XOR2_X1 U1085 ( .A(n1035), .B(n1355), .Z(n1354) );
NAND2_X1 U1086 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1087 ( .A1(n1358), .A2(n1236), .ZN(n1357) );
XOR2_X1 U1088 ( .A(n1359), .B(KEYINPUT30), .Z(n1356) );
OR2_X1 U1089 ( .A1(n1358), .A2(n1236), .ZN(n1359) );
INV_X1 U1090 ( .A(G122), .ZN(n1236) );
XOR2_X1 U1091 ( .A(G116), .B(KEYINPUT43), .Z(n1358) );
INV_X1 U1092 ( .A(G107), .ZN(n1035) );
NAND3_X1 U1093 ( .A1(G234), .A2(n1097), .A3(G217), .ZN(n1353) );
INV_X1 U1094 ( .A(G953), .ZN(n1097) );
endmodule


