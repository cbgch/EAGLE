//Key = 1001110010110111111011100101000000011000000001010000010011110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367;

NAND2_X1 U747 ( .A1(n1036), .A2(n1037), .ZN(G9) );
NAND2_X1 U748 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XOR2_X1 U749 ( .A(KEYINPUT14), .B(n1040), .Z(n1036) );
NOR2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1040) );
INV_X1 U751 ( .A(n1041), .ZN(n1038) );
NOR2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
XOR2_X1 U754 ( .A(KEYINPUT31), .B(n1048), .Z(n1045) );
NOR3_X1 U755 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND4_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1044) );
NAND4_X1 U757 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1054) );
NAND2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U761 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1060) );
NAND2_X1 U763 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1053) );
NAND2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U767 ( .A1(n1058), .A2(n1078), .ZN(n1077) );
NAND2_X1 U768 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U769 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U770 ( .A1(n1057), .A2(n1083), .ZN(n1076) );
INV_X1 U771 ( .A(n1049), .ZN(n1074) );
NAND3_X1 U772 ( .A1(n1062), .A2(n1068), .A3(n1056), .ZN(n1049) );
INV_X1 U773 ( .A(n1084), .ZN(n1056) );
XOR2_X1 U774 ( .A(KEYINPUT12), .B(n1085), .Z(n1052) );
NOR3_X1 U775 ( .A1(n1047), .A2(G952), .A3(n1086), .ZN(n1042) );
INV_X1 U776 ( .A(n1055), .ZN(n1086) );
NAND4_X1 U777 ( .A1(n1087), .A2(n1068), .A3(n1088), .A4(n1089), .ZN(n1055) );
NOR4_X1 U778 ( .A1(n1081), .A2(n1072), .A3(n1090), .A4(n1091), .ZN(n1089) );
XNOR2_X1 U779 ( .A(n1092), .B(KEYINPUT53), .ZN(n1090) );
INV_X1 U780 ( .A(n1093), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1088) );
XNOR2_X1 U782 ( .A(G478), .B(n1096), .ZN(n1087) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(G72) );
OR3_X1 U784 ( .A1(n1099), .A2(KEYINPUT42), .A3(n1100), .ZN(n1098) );
NAND3_X1 U785 ( .A1(n1101), .A2(n1102), .A3(n1100), .ZN(n1097) );
XOR2_X1 U786 ( .A(n1103), .B(n1104), .Z(n1100) );
NAND2_X1 U787 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XOR2_X1 U789 ( .A(n1109), .B(n1110), .Z(n1105) );
XNOR2_X1 U790 ( .A(n1111), .B(n1112), .ZN(n1110) );
NAND2_X1 U791 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NAND2_X1 U792 ( .A1(G140), .A2(n1115), .ZN(n1114) );
XOR2_X1 U793 ( .A(n1116), .B(KEYINPUT49), .Z(n1113) );
OR2_X1 U794 ( .A1(n1115), .A2(G140), .ZN(n1116) );
XOR2_X1 U795 ( .A(G131), .B(n1117), .Z(n1109) );
XNOR2_X1 U796 ( .A(n1118), .B(G134), .ZN(n1117) );
NAND3_X1 U797 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1103) );
XNOR2_X1 U798 ( .A(KEYINPUT35), .B(n1122), .ZN(n1121) );
OR2_X1 U799 ( .A1(n1123), .A2(KEYINPUT21), .ZN(n1120) );
NAND2_X1 U800 ( .A1(KEYINPUT21), .A2(n1085), .ZN(n1119) );
NAND2_X1 U801 ( .A1(KEYINPUT32), .A2(n1099), .ZN(n1102) );
OR3_X1 U802 ( .A1(KEYINPUT32), .A2(KEYINPUT42), .A3(n1099), .ZN(n1101) );
NAND2_X1 U803 ( .A1(G953), .A2(n1124), .ZN(n1099) );
NAND2_X1 U804 ( .A1(G900), .A2(G227), .ZN(n1124) );
XOR2_X1 U805 ( .A(n1125), .B(n1126), .Z(G69) );
XOR2_X1 U806 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND3_X1 U807 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
XOR2_X1 U808 ( .A(KEYINPUT5), .B(n1132), .Z(n1131) );
NOR2_X1 U809 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XNOR2_X1 U810 ( .A(n1135), .B(KEYINPUT11), .ZN(n1134) );
INV_X1 U811 ( .A(n1136), .ZN(n1130) );
NAND3_X1 U812 ( .A1(n1137), .A2(n1122), .A3(KEYINPUT47), .ZN(n1127) );
XNOR2_X1 U813 ( .A(KEYINPUT45), .B(n1046), .ZN(n1137) );
NOR2_X1 U814 ( .A1(n1138), .A2(n1122), .ZN(n1125) );
AND2_X1 U815 ( .A1(G224), .A2(G898), .ZN(n1138) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U818 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NOR2_X1 U819 ( .A1(n1139), .A2(n1145), .ZN(G63) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U821 ( .A1(n1148), .A2(G478), .ZN(n1147) );
NAND2_X1 U822 ( .A1(KEYINPUT58), .A2(n1149), .ZN(n1146) );
NOR2_X1 U823 ( .A1(n1139), .A2(n1150), .ZN(G60) );
XNOR2_X1 U824 ( .A(n1151), .B(n1152), .ZN(n1150) );
AND2_X1 U825 ( .A1(G475), .A2(n1148), .ZN(n1152) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(G6) );
NAND2_X1 U827 ( .A1(KEYINPUT17), .A2(G104), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(G57) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U830 ( .A(n1159), .B(n1160), .ZN(n1158) );
XOR2_X1 U831 ( .A(n1161), .B(n1162), .Z(n1157) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1162) );
AND2_X1 U833 ( .A1(G472), .A2(n1148), .ZN(n1164) );
NOR2_X1 U834 ( .A1(KEYINPUT62), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U835 ( .A(n1166), .B(KEYINPUT54), .ZN(n1165) );
NAND2_X1 U836 ( .A1(n1167), .A2(n1168), .ZN(n1161) );
NAND3_X1 U837 ( .A1(G210), .A2(n1169), .A3(G101), .ZN(n1168) );
XOR2_X1 U838 ( .A(n1170), .B(KEYINPUT23), .Z(n1167) );
NOR2_X1 U839 ( .A1(G952), .A2(n1171), .ZN(n1155) );
XNOR2_X1 U840 ( .A(G953), .B(KEYINPUT46), .ZN(n1171) );
NOR2_X1 U841 ( .A1(n1139), .A2(n1172), .ZN(G54) );
XOR2_X1 U842 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U843 ( .A1(n1148), .A2(G469), .ZN(n1174) );
INV_X1 U844 ( .A(n1144), .ZN(n1148) );
NAND2_X1 U845 ( .A1(n1175), .A2(KEYINPUT18), .ZN(n1173) );
XOR2_X1 U846 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U847 ( .A(n1178), .B(n1179), .ZN(n1177) );
XNOR2_X1 U848 ( .A(n1180), .B(n1181), .ZN(n1176) );
NAND2_X1 U849 ( .A1(KEYINPUT57), .A2(n1182), .ZN(n1180) );
NOR2_X1 U850 ( .A1(n1139), .A2(n1183), .ZN(G51) );
XOR2_X1 U851 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U852 ( .A1(n1095), .A2(n1144), .ZN(n1185) );
NAND2_X1 U853 ( .A1(G902), .A2(n1186), .ZN(n1144) );
NAND2_X1 U854 ( .A1(n1187), .A2(n1085), .ZN(n1186) );
AND4_X1 U855 ( .A1(n1188), .A2(n1189), .A3(n1123), .A4(n1190), .ZN(n1085) );
AND4_X1 U856 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190) );
NAND3_X1 U857 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1123) );
XNOR2_X1 U858 ( .A(n1198), .B(KEYINPUT56), .ZN(n1197) );
NAND2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1189) );
XNOR2_X1 U860 ( .A(KEYINPUT9), .B(n1201), .ZN(n1200) );
INV_X1 U861 ( .A(n1202), .ZN(n1199) );
NAND2_X1 U862 ( .A1(n1203), .A2(n1204), .ZN(n1188) );
NAND2_X1 U863 ( .A1(n1205), .A2(n1202), .ZN(n1204) );
NAND2_X1 U864 ( .A1(n1206), .A2(n1062), .ZN(n1205) );
INV_X1 U865 ( .A(n1046), .ZN(n1187) );
NAND4_X1 U866 ( .A1(n1207), .A2(n1041), .A3(n1208), .A4(n1209), .ZN(n1046) );
AND3_X1 U867 ( .A1(n1210), .A2(n1211), .A3(n1153), .ZN(n1209) );
NAND3_X1 U868 ( .A1(n1068), .A2(n1212), .A3(n1203), .ZN(n1153) );
OR2_X1 U869 ( .A1(n1213), .A2(n1064), .ZN(n1210) );
NOR2_X1 U870 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
AND2_X1 U871 ( .A1(n1212), .A2(n1058), .ZN(n1215) );
NOR2_X1 U872 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NOR2_X1 U873 ( .A1(n1083), .A2(n1203), .ZN(n1216) );
NAND3_X1 U874 ( .A1(n1212), .A2(n1083), .A3(n1068), .ZN(n1041) );
XOR2_X1 U875 ( .A(n1218), .B(n1219), .Z(n1184) );
NOR2_X1 U876 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NOR2_X1 U877 ( .A1(n1122), .A2(G952), .ZN(n1139) );
XNOR2_X1 U878 ( .A(n1222), .B(n1223), .ZN(G48) );
NOR2_X1 U879 ( .A1(n1051), .A2(n1202), .ZN(n1223) );
XNOR2_X1 U880 ( .A(G143), .B(n1194), .ZN(G45) );
NAND4_X1 U881 ( .A1(n1224), .A2(n1206), .A3(n1225), .A4(n1226), .ZN(n1194) );
XNOR2_X1 U882 ( .A(KEYINPUT50), .B(n1227), .ZN(n1226) );
XNOR2_X1 U883 ( .A(G140), .B(n1192), .ZN(G42) );
NAND3_X1 U884 ( .A1(n1062), .A2(n1198), .A3(n1228), .ZN(n1192) );
XNOR2_X1 U885 ( .A(G137), .B(n1229), .ZN(G39) );
NAND3_X1 U886 ( .A1(n1195), .A2(n1198), .A3(n1230), .ZN(n1229) );
XNOR2_X1 U887 ( .A(n1196), .B(KEYINPUT10), .ZN(n1230) );
AND3_X1 U888 ( .A1(n1058), .A2(n1231), .A3(n1062), .ZN(n1195) );
XNOR2_X1 U889 ( .A(G134), .B(n1191), .ZN(G36) );
NAND3_X1 U890 ( .A1(n1062), .A2(n1083), .A3(n1206), .ZN(n1191) );
INV_X1 U891 ( .A(n1232), .ZN(n1206) );
XOR2_X1 U892 ( .A(G131), .B(n1233), .Z(G33) );
NOR4_X1 U893 ( .A1(KEYINPUT6), .A2(n1234), .A3(n1051), .A4(n1232), .ZN(n1233) );
NAND3_X1 U894 ( .A1(n1198), .A2(n1231), .A3(n1235), .ZN(n1232) );
INV_X1 U895 ( .A(n1203), .ZN(n1051) );
XNOR2_X1 U896 ( .A(n1062), .B(KEYINPUT44), .ZN(n1234) );
AND2_X1 U897 ( .A1(n1073), .A2(n1236), .ZN(n1062) );
XOR2_X1 U898 ( .A(G128), .B(n1237), .Z(G30) );
NOR2_X1 U899 ( .A1(n1201), .A2(n1202), .ZN(n1237) );
NAND4_X1 U900 ( .A1(n1196), .A2(n1225), .A3(n1198), .A4(n1231), .ZN(n1202) );
NAND2_X1 U901 ( .A1(n1238), .A2(n1239), .ZN(G3) );
NAND2_X1 U902 ( .A1(G101), .A2(n1240), .ZN(n1239) );
XOR2_X1 U903 ( .A(KEYINPUT25), .B(n1241), .Z(n1238) );
NOR2_X1 U904 ( .A1(G101), .A2(n1240), .ZN(n1241) );
NAND3_X1 U905 ( .A1(n1058), .A2(n1212), .A3(n1235), .ZN(n1240) );
XNOR2_X1 U906 ( .A(G125), .B(n1193), .ZN(G27) );
NAND3_X1 U907 ( .A1(n1057), .A2(n1225), .A3(n1228), .ZN(n1193) );
AND4_X1 U908 ( .A1(n1066), .A2(n1203), .A3(n1231), .A4(n1067), .ZN(n1228) );
NAND2_X1 U909 ( .A1(n1084), .A2(n1242), .ZN(n1231) );
NAND4_X1 U910 ( .A1(G902), .A2(n1107), .A3(n1243), .A4(n1108), .ZN(n1242) );
INV_X1 U911 ( .A(G900), .ZN(n1108) );
XNOR2_X1 U912 ( .A(G122), .B(n1211), .ZN(G24) );
NAND4_X1 U913 ( .A1(n1244), .A2(n1068), .A3(n1245), .A4(n1246), .ZN(n1211) );
NAND2_X1 U914 ( .A1(KEYINPUT50), .A2(n1201), .ZN(n1246) );
NAND2_X1 U915 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
INV_X1 U916 ( .A(KEYINPUT50), .ZN(n1248) );
NAND2_X1 U917 ( .A1(n1224), .A2(n1092), .ZN(n1247) );
AND2_X1 U918 ( .A1(n1249), .A2(n1250), .ZN(n1068) );
XNOR2_X1 U919 ( .A(G119), .B(n1208), .ZN(G21) );
NAND3_X1 U920 ( .A1(n1196), .A2(n1058), .A3(n1244), .ZN(n1208) );
AND2_X1 U921 ( .A1(n1251), .A2(n1067), .ZN(n1196) );
XNOR2_X1 U922 ( .A(G116), .B(n1252), .ZN(G18) );
NAND4_X1 U923 ( .A1(n1235), .A2(n1083), .A3(n1253), .A4(n1254), .ZN(n1252) );
OR2_X1 U924 ( .A1(n1244), .A2(KEYINPUT2), .ZN(n1254) );
NAND2_X1 U925 ( .A1(KEYINPUT2), .A2(n1255), .ZN(n1253) );
NAND2_X1 U926 ( .A1(n1256), .A2(n1070), .ZN(n1255) );
INV_X1 U927 ( .A(n1225), .ZN(n1070) );
INV_X1 U928 ( .A(n1201), .ZN(n1083) );
NAND2_X1 U929 ( .A1(n1224), .A2(n1227), .ZN(n1201) );
XNOR2_X1 U930 ( .A(n1257), .B(n1258), .ZN(G15) );
NAND2_X1 U931 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND4_X1 U932 ( .A1(n1261), .A2(n1244), .A3(n1235), .A4(n1262), .ZN(n1260) );
INV_X1 U933 ( .A(KEYINPUT30), .ZN(n1262) );
INV_X1 U934 ( .A(n1217), .ZN(n1244) );
NAND2_X1 U935 ( .A1(n1256), .A2(n1225), .ZN(n1217) );
NAND3_X1 U936 ( .A1(n1225), .A2(n1263), .A3(KEYINPUT30), .ZN(n1259) );
NAND3_X1 U937 ( .A1(n1235), .A2(n1256), .A3(n1261), .ZN(n1263) );
XNOR2_X1 U938 ( .A(n1203), .B(KEYINPUT8), .ZN(n1261) );
NOR2_X1 U939 ( .A1(n1227), .A2(n1224), .ZN(n1203) );
INV_X1 U940 ( .A(n1092), .ZN(n1227) );
AND2_X1 U941 ( .A1(n1057), .A2(n1264), .ZN(n1256) );
INV_X1 U942 ( .A(n1050), .ZN(n1057) );
NAND2_X1 U943 ( .A1(n1082), .A2(n1093), .ZN(n1050) );
INV_X1 U944 ( .A(n1064), .ZN(n1235) );
NAND2_X1 U945 ( .A1(n1251), .A2(n1249), .ZN(n1064) );
INV_X1 U946 ( .A(n1067), .ZN(n1249) );
XOR2_X1 U947 ( .A(n1250), .B(KEYINPUT27), .Z(n1251) );
XNOR2_X1 U948 ( .A(G110), .B(n1207), .ZN(G12) );
NAND4_X1 U949 ( .A1(n1066), .A2(n1058), .A3(n1212), .A4(n1067), .ZN(n1207) );
NAND3_X1 U950 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1067) );
NAND2_X1 U951 ( .A1(G902), .A2(G217), .ZN(n1267) );
OR3_X1 U952 ( .A1(n1142), .A2(G902), .A3(n1268), .ZN(n1266) );
NAND2_X1 U953 ( .A1(n1142), .A2(n1268), .ZN(n1265) );
NOR2_X1 U954 ( .A1(n1143), .A2(G234), .ZN(n1268) );
INV_X1 U955 ( .A(G217), .ZN(n1143) );
XNOR2_X1 U956 ( .A(n1269), .B(n1270), .ZN(n1142) );
XOR2_X1 U957 ( .A(n1271), .B(n1272), .Z(n1270) );
XNOR2_X1 U958 ( .A(n1273), .B(n1274), .ZN(n1272) );
NOR2_X1 U959 ( .A1(KEYINPUT48), .A2(n1222), .ZN(n1274) );
INV_X1 U960 ( .A(G146), .ZN(n1222) );
NAND2_X1 U961 ( .A1(KEYINPUT13), .A2(n1118), .ZN(n1273) );
XOR2_X1 U962 ( .A(n1275), .B(n1276), .Z(n1269) );
XOR2_X1 U963 ( .A(G128), .B(G119), .Z(n1276) );
XNOR2_X1 U964 ( .A(n1277), .B(n1278), .ZN(n1275) );
NAND2_X1 U965 ( .A1(G221), .A2(n1279), .ZN(n1277) );
AND3_X1 U966 ( .A1(n1198), .A2(n1264), .A3(n1225), .ZN(n1212) );
NOR2_X1 U967 ( .A1(n1073), .A2(n1072), .ZN(n1225) );
INV_X1 U968 ( .A(n1236), .ZN(n1072) );
NAND2_X1 U969 ( .A1(G214), .A2(n1280), .ZN(n1236) );
XNOR2_X1 U970 ( .A(n1095), .B(n1281), .ZN(n1073) );
NOR2_X1 U971 ( .A1(n1094), .A2(KEYINPUT1), .ZN(n1281) );
AND2_X1 U972 ( .A1(n1282), .A2(n1283), .ZN(n1094) );
XOR2_X1 U973 ( .A(n1284), .B(n1285), .Z(n1282) );
NOR4_X1 U974 ( .A1(n1286), .A2(n1287), .A3(KEYINPUT37), .A4(n1220), .ZN(n1285) );
NOR3_X1 U975 ( .A1(n1115), .A2(n1288), .A3(n1112), .ZN(n1220) );
AND2_X1 U976 ( .A1(n1289), .A2(n1221), .ZN(n1287) );
NAND2_X1 U977 ( .A1(n1290), .A2(n1291), .ZN(n1221) );
NAND2_X1 U978 ( .A1(n1292), .A2(n1115), .ZN(n1291) );
XNOR2_X1 U979 ( .A(n1288), .B(n1159), .ZN(n1292) );
NAND3_X1 U980 ( .A1(n1288), .A2(n1112), .A3(G125), .ZN(n1290) );
INV_X1 U981 ( .A(n1293), .ZN(n1288) );
NOR2_X1 U982 ( .A1(n1294), .A2(n1289), .ZN(n1286) );
INV_X1 U983 ( .A(KEYINPUT40), .ZN(n1289) );
XNOR2_X1 U984 ( .A(n1293), .B(n1295), .ZN(n1294) );
NOR2_X1 U985 ( .A1(G125), .A2(n1159), .ZN(n1295) );
NAND2_X1 U986 ( .A1(G224), .A2(n1122), .ZN(n1293) );
XOR2_X1 U987 ( .A(n1218), .B(KEYINPUT15), .Z(n1284) );
NAND2_X1 U988 ( .A1(n1129), .A2(n1296), .ZN(n1218) );
OR2_X1 U989 ( .A1(n1135), .A2(n1133), .ZN(n1296) );
NAND2_X1 U990 ( .A1(n1133), .A2(n1135), .ZN(n1129) );
XNOR2_X1 U991 ( .A(n1297), .B(n1298), .ZN(n1135) );
XNOR2_X1 U992 ( .A(n1039), .B(G104), .ZN(n1298) );
XNOR2_X1 U993 ( .A(n1299), .B(n1300), .ZN(n1297) );
XNOR2_X1 U994 ( .A(G110), .B(G122), .ZN(n1133) );
NAND2_X1 U995 ( .A1(G210), .A2(n1280), .ZN(n1095) );
NAND2_X1 U996 ( .A1(n1301), .A2(n1283), .ZN(n1280) );
INV_X1 U997 ( .A(G237), .ZN(n1301) );
NAND2_X1 U998 ( .A1(n1084), .A2(n1302), .ZN(n1264) );
NAND3_X1 U999 ( .A1(G902), .A2(n1243), .A3(n1136), .ZN(n1302) );
NOR2_X1 U1000 ( .A1(n1303), .A2(G898), .ZN(n1136) );
INV_X1 U1001 ( .A(n1107), .ZN(n1303) );
XNOR2_X1 U1002 ( .A(n1122), .B(KEYINPUT28), .ZN(n1107) );
NAND3_X1 U1003 ( .A1(n1304), .A2(n1243), .A3(G952), .ZN(n1084) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1243) );
INV_X1 U1005 ( .A(n1047), .ZN(n1304) );
XOR2_X1 U1006 ( .A(G953), .B(KEYINPUT63), .Z(n1047) );
INV_X1 U1007 ( .A(n1079), .ZN(n1198) );
NAND2_X1 U1008 ( .A1(n1305), .A2(n1093), .ZN(n1079) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1306), .ZN(n1093) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1283), .ZN(n1306) );
XOR2_X1 U1011 ( .A(KEYINPUT59), .B(n1082), .Z(n1305) );
XOR2_X1 U1012 ( .A(n1091), .B(KEYINPUT3), .Z(n1082) );
XNOR2_X1 U1013 ( .A(n1307), .B(G469), .ZN(n1091) );
NAND2_X1 U1014 ( .A1(n1283), .A2(n1308), .ZN(n1307) );
NAND2_X1 U1015 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND2_X1 U1016 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XNOR2_X1 U1017 ( .A(KEYINPUT22), .B(n1313), .ZN(n1312) );
XNOR2_X1 U1018 ( .A(n1181), .B(n1182), .ZN(n1311) );
XOR2_X1 U1019 ( .A(n1314), .B(KEYINPUT19), .Z(n1309) );
NAND2_X1 U1020 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U1021 ( .A(n1313), .B(KEYINPUT22), .Z(n1316) );
NAND3_X1 U1022 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(n1313) );
OR2_X1 U1023 ( .A1(n1320), .A2(n1178), .ZN(n1319) );
NAND3_X1 U1024 ( .A1(n1178), .A2(n1320), .A3(n1166), .ZN(n1318) );
NAND2_X1 U1025 ( .A1(n1179), .A2(n1321), .ZN(n1317) );
NAND2_X1 U1026 ( .A1(n1322), .A2(n1320), .ZN(n1321) );
INV_X1 U1027 ( .A(KEYINPUT52), .ZN(n1320) );
XNOR2_X1 U1028 ( .A(n1178), .B(KEYINPUT16), .ZN(n1322) );
XOR2_X1 U1029 ( .A(n1112), .B(n1323), .Z(n1178) );
XNOR2_X1 U1030 ( .A(n1300), .B(n1324), .ZN(n1323) );
NOR4_X1 U1031 ( .A1(n1325), .A2(n1326), .A3(KEYINPUT24), .A4(n1327), .ZN(n1324) );
AND2_X1 U1032 ( .A1(n1328), .A2(G104), .ZN(n1327) );
NOR2_X1 U1033 ( .A1(n1329), .A2(n1039), .ZN(n1326) );
NOR2_X1 U1034 ( .A1(G104), .A2(KEYINPUT34), .ZN(n1329) );
NOR4_X1 U1035 ( .A1(G107), .A2(n1328), .A3(KEYINPUT34), .A4(G104), .ZN(n1325) );
INV_X1 U1036 ( .A(KEYINPUT4), .ZN(n1328) );
XOR2_X1 U1037 ( .A(n1181), .B(n1182), .Z(n1315) );
XNOR2_X1 U1038 ( .A(n1278), .B(G140), .ZN(n1182) );
INV_X1 U1039 ( .A(G110), .ZN(n1278) );
NAND2_X1 U1040 ( .A1(G227), .A2(n1122), .ZN(n1181) );
NOR2_X1 U1041 ( .A1(n1092), .A2(n1224), .ZN(n1058) );
XOR2_X1 U1042 ( .A(n1330), .B(n1331), .Z(n1224) );
XOR2_X1 U1043 ( .A(KEYINPUT55), .B(n1096), .Z(n1331) );
NOR2_X1 U1044 ( .A1(n1149), .A2(G902), .ZN(n1096) );
XNOR2_X1 U1045 ( .A(n1332), .B(n1333), .ZN(n1149) );
XOR2_X1 U1046 ( .A(G128), .B(n1334), .Z(n1333) );
XNOR2_X1 U1047 ( .A(n1335), .B(G134), .ZN(n1334) );
INV_X1 U1048 ( .A(G143), .ZN(n1335) );
XOR2_X1 U1049 ( .A(n1336), .B(n1337), .Z(n1332) );
NOR2_X1 U1050 ( .A1(KEYINPUT41), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1051 ( .A(n1039), .B(n1339), .ZN(n1338) );
XOR2_X1 U1052 ( .A(G122), .B(G116), .Z(n1339) );
INV_X1 U1053 ( .A(G107), .ZN(n1039) );
NAND2_X1 U1054 ( .A1(n1279), .A2(G217), .ZN(n1336) );
AND2_X1 U1055 ( .A1(G234), .A2(n1122), .ZN(n1279) );
INV_X1 U1056 ( .A(G953), .ZN(n1122) );
NAND2_X1 U1057 ( .A1(KEYINPUT20), .A2(n1340), .ZN(n1330) );
INV_X1 U1058 ( .A(G478), .ZN(n1340) );
XNOR2_X1 U1059 ( .A(n1341), .B(G475), .ZN(n1092) );
NAND2_X1 U1060 ( .A1(n1151), .A2(n1283), .ZN(n1341) );
XNOR2_X1 U1061 ( .A(n1342), .B(n1343), .ZN(n1151) );
XNOR2_X1 U1062 ( .A(n1344), .B(n1345), .ZN(n1343) );
XNOR2_X1 U1063 ( .A(n1346), .B(n1347), .ZN(n1345) );
NOR2_X1 U1064 ( .A1(KEYINPUT26), .A2(n1258), .ZN(n1347) );
INV_X1 U1065 ( .A(G113), .ZN(n1258) );
NOR2_X1 U1066 ( .A1(KEYINPUT33), .A2(n1348), .ZN(n1346) );
XOR2_X1 U1067 ( .A(KEYINPUT36), .B(n1271), .Z(n1348) );
XNOR2_X1 U1068 ( .A(G140), .B(n1115), .ZN(n1271) );
INV_X1 U1069 ( .A(G125), .ZN(n1115) );
XOR2_X1 U1070 ( .A(n1349), .B(n1350), .Z(n1342) );
XOR2_X1 U1071 ( .A(G131), .B(G122), .Z(n1350) );
XOR2_X1 U1072 ( .A(n1351), .B(G104), .Z(n1349) );
NAND2_X1 U1073 ( .A1(G214), .A2(n1169), .ZN(n1351) );
XOR2_X1 U1074 ( .A(n1250), .B(KEYINPUT38), .Z(n1066) );
XOR2_X1 U1075 ( .A(n1352), .B(G472), .Z(n1250) );
NAND2_X1 U1076 ( .A1(n1353), .A2(n1283), .ZN(n1352) );
INV_X1 U1077 ( .A(G902), .ZN(n1283) );
XNOR2_X1 U1078 ( .A(n1160), .B(n1354), .ZN(n1353) );
XOR2_X1 U1079 ( .A(n1355), .B(n1356), .Z(n1354) );
NOR2_X1 U1080 ( .A1(KEYINPUT39), .A2(n1357), .ZN(n1356) );
XNOR2_X1 U1081 ( .A(n1358), .B(n1112), .ZN(n1357) );
INV_X1 U1082 ( .A(n1159), .ZN(n1112) );
XNOR2_X1 U1083 ( .A(G128), .B(n1344), .ZN(n1159) );
XOR2_X1 U1084 ( .A(G143), .B(G146), .Z(n1344) );
NAND2_X1 U1085 ( .A1(KEYINPUT0), .A2(n1179), .ZN(n1358) );
INV_X1 U1086 ( .A(n1166), .ZN(n1179) );
XOR2_X1 U1087 ( .A(G131), .B(n1359), .Z(n1166) );
NOR2_X1 U1088 ( .A1(KEYINPUT43), .A2(n1360), .ZN(n1359) );
XNOR2_X1 U1089 ( .A(n1118), .B(n1361), .ZN(n1360) );
NOR2_X1 U1090 ( .A1(G134), .A2(KEYINPUT51), .ZN(n1361) );
INV_X1 U1091 ( .A(G137), .ZN(n1118) );
NAND2_X1 U1092 ( .A1(n1362), .A2(n1170), .ZN(n1355) );
NAND2_X1 U1093 ( .A1(n1300), .A2(n1363), .ZN(n1170) );
NAND2_X1 U1094 ( .A1(G210), .A2(n1169), .ZN(n1363) );
INV_X1 U1095 ( .A(G101), .ZN(n1300) );
XOR2_X1 U1096 ( .A(n1364), .B(KEYINPUT29), .Z(n1362) );
NAND3_X1 U1097 ( .A1(G210), .A2(n1169), .A3(n1365), .ZN(n1364) );
XNOR2_X1 U1098 ( .A(G101), .B(KEYINPUT61), .ZN(n1365) );
NOR2_X1 U1099 ( .A1(G237), .A2(G953), .ZN(n1169) );
XNOR2_X1 U1100 ( .A(n1299), .B(n1366), .ZN(n1160) );
XOR2_X1 U1101 ( .A(KEYINPUT7), .B(KEYINPUT60), .Z(n1366) );
XNOR2_X1 U1102 ( .A(G113), .B(n1367), .ZN(n1299) );
XOR2_X1 U1103 ( .A(G119), .B(G116), .Z(n1367) );
endmodule


