//Key = 1000001010111101111101010111101001000000100101101110101111101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302;

XNOR2_X1 U717 ( .A(G107), .B(n988), .ZN(G9) );
NAND3_X1 U718 ( .A1(n989), .A2(n990), .A3(n991), .ZN(G75) );
NAND2_X1 U719 ( .A1(G952), .A2(n992), .ZN(n991) );
NAND2_X1 U720 ( .A1(n993), .A2(n994), .ZN(n992) );
NAND2_X1 U721 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U722 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND3_X1 U723 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NAND2_X1 U724 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NAND3_X1 U725 ( .A1(n1004), .A2(n1005), .A3(KEYINPUT32), .ZN(n1002) );
NAND3_X1 U726 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n999) );
NAND2_X1 U727 ( .A1(n1005), .A2(n1009), .ZN(n1007) );
NAND2_X1 U728 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
OR2_X1 U729 ( .A1(n1012), .A2(KEYINPUT32), .ZN(n1011) );
NAND2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1006) );
NAND2_X1 U731 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U732 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND3_X1 U733 ( .A1(n1005), .A2(n1019), .A3(n1013), .ZN(n997) );
NAND2_X1 U734 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U735 ( .A1(n1001), .A2(n1022), .ZN(n1021) );
NAND2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U737 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U738 ( .A1(n1008), .A2(n1027), .ZN(n1020) );
NAND2_X1 U739 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U740 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
XNOR2_X1 U741 ( .A(KEYINPUT54), .B(n1032), .ZN(n995) );
NAND4_X1 U742 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n989) );
NOR4_X1 U743 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
NOR2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(n1037) );
NOR2_X1 U745 ( .A1(n1003), .A2(n1043), .ZN(n1035) );
XOR2_X1 U746 ( .A(n1044), .B(n1045), .Z(n1043) );
XOR2_X1 U747 ( .A(KEYINPUT11), .B(G475), .Z(n1045) );
NOR2_X1 U748 ( .A1(KEYINPUT62), .A2(n1046), .ZN(n1044) );
NAND2_X1 U749 ( .A1(n1047), .A2(n1048), .ZN(n1034) );
INV_X1 U750 ( .A(KEYINPUT12), .ZN(n1048) );
NAND2_X1 U751 ( .A1(n1049), .A2(n1042), .ZN(n1047) );
XNOR2_X1 U752 ( .A(n1041), .B(KEYINPUT30), .ZN(n1049) );
NAND2_X1 U753 ( .A1(KEYINPUT12), .A2(n1050), .ZN(n1033) );
NAND2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
OR2_X1 U755 ( .A1(n1041), .A2(KEYINPUT30), .ZN(n1052) );
NAND3_X1 U756 ( .A1(n1041), .A2(n1042), .A3(KEYINPUT30), .ZN(n1051) );
XOR2_X1 U757 ( .A(n1053), .B(n1054), .Z(G72) );
NOR2_X1 U758 ( .A1(n1055), .A2(n990), .ZN(n1054) );
AND2_X1 U759 ( .A1(G227), .A2(G900), .ZN(n1055) );
NAND2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NAND3_X1 U761 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NAND2_X1 U762 ( .A1(G953), .A2(n1061), .ZN(n1059) );
XNOR2_X1 U763 ( .A(KEYINPUT41), .B(n1062), .ZN(n1058) );
NAND3_X1 U764 ( .A1(n1062), .A2(n990), .A3(n1063), .ZN(n1056) );
INV_X1 U765 ( .A(n1060), .ZN(n1063) );
XOR2_X1 U766 ( .A(n1064), .B(n1065), .Z(n1060) );
XOR2_X1 U767 ( .A(n1066), .B(n1067), .Z(n1065) );
NAND2_X1 U768 ( .A1(KEYINPUT61), .A2(n1068), .ZN(n1067) );
XOR2_X1 U769 ( .A(n1069), .B(n1070), .Z(n1068) );
XOR2_X1 U770 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U771 ( .A1(KEYINPUT40), .A2(n1073), .ZN(n1071) );
NAND2_X1 U772 ( .A1(KEYINPUT43), .A2(n1074), .ZN(n1064) );
XOR2_X1 U773 ( .A(n1075), .B(n1076), .Z(G69) );
XOR2_X1 U774 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U776 ( .A1(G953), .A2(n1081), .ZN(n1080) );
XNOR2_X1 U777 ( .A(n1082), .B(n1083), .ZN(n1079) );
NAND2_X1 U778 ( .A1(KEYINPUT25), .A2(n1084), .ZN(n1082) );
NAND2_X1 U779 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U780 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U781 ( .A(n1089), .B(KEYINPUT9), .Z(n1085) );
OR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(n1089) );
NAND2_X1 U783 ( .A1(G953), .A2(n1090), .ZN(n1077) );
NAND2_X1 U784 ( .A1(n1091), .A2(G224), .ZN(n1090) );
XOR2_X1 U785 ( .A(n1081), .B(KEYINPUT48), .Z(n1091) );
AND2_X1 U786 ( .A1(n1092), .A2(n990), .ZN(n1075) );
NOR2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(G66) );
XOR2_X1 U788 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U789 ( .A1(n1042), .A2(n1097), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1093), .A2(n1098), .ZN(G63) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U792 ( .A1(KEYINPUT59), .A2(n1101), .ZN(n1099) );
NOR3_X1 U793 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
INV_X1 U794 ( .A(G478), .ZN(n1103) );
XOR2_X1 U795 ( .A(KEYINPUT22), .B(n993), .Z(n1102) );
NOR3_X1 U796 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(G60) );
AND2_X1 U797 ( .A1(KEYINPUT50), .A2(n1093), .ZN(n1107) );
NOR3_X1 U798 ( .A1(KEYINPUT50), .A2(G953), .A3(G952), .ZN(n1106) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(n1105) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1097), .ZN(n1108) );
INV_X1 U801 ( .A(G475), .ZN(n1110) );
XOR2_X1 U802 ( .A(n1111), .B(n1112), .Z(G6) );
NOR2_X1 U803 ( .A1(n1093), .A2(n1113), .ZN(G57) );
NOR3_X1 U804 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U806 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
XOR2_X1 U807 ( .A(KEYINPUT37), .B(n1121), .Z(n1120) );
NOR3_X1 U808 ( .A1(n1122), .A2(n1121), .A3(n1119), .ZN(n1115) );
INV_X1 U809 ( .A(n1118), .ZN(n1122) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1118) );
XOR2_X1 U811 ( .A(KEYINPUT60), .B(n1125), .Z(n1124) );
NOR3_X1 U812 ( .A1(KEYINPUT39), .A2(n1126), .A3(n1127), .ZN(n1125) );
AND2_X1 U813 ( .A1(n1128), .A2(KEYINPUT28), .ZN(n1127) );
NOR2_X1 U814 ( .A1(KEYINPUT28), .A2(n1129), .ZN(n1126) );
AND2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U816 ( .A(n1132), .B(n1133), .ZN(n1123) );
NOR2_X1 U817 ( .A1(n1134), .A2(n1097), .ZN(n1133) );
INV_X1 U818 ( .A(G472), .ZN(n1134) );
AND2_X1 U819 ( .A1(n1119), .A2(n1121), .ZN(n1114) );
INV_X1 U820 ( .A(KEYINPUT0), .ZN(n1119) );
NOR2_X1 U821 ( .A1(n1093), .A2(n1135), .ZN(G54) );
XOR2_X1 U822 ( .A(n1136), .B(n1137), .Z(n1135) );
XNOR2_X1 U823 ( .A(n1138), .B(n1139), .ZN(n1137) );
XOR2_X1 U824 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U825 ( .A1(n1142), .A2(n1097), .ZN(n1141) );
INV_X1 U826 ( .A(G469), .ZN(n1142) );
NAND2_X1 U827 ( .A1(KEYINPUT56), .A2(n1074), .ZN(n1140) );
XOR2_X1 U828 ( .A(n1143), .B(n1144), .Z(n1136) );
XOR2_X1 U829 ( .A(G110), .B(n1145), .Z(n1144) );
NOR2_X1 U830 ( .A1(KEYINPUT4), .A2(n1146), .ZN(n1145) );
NAND2_X1 U831 ( .A1(KEYINPUT49), .A2(n1131), .ZN(n1143) );
NOR2_X1 U832 ( .A1(n1093), .A2(n1147), .ZN(G51) );
XOR2_X1 U833 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR3_X1 U834 ( .A1(n1150), .A2(n1151), .A3(n1097), .ZN(n1149) );
OR2_X1 U835 ( .A1(n1104), .A2(n993), .ZN(n1097) );
NOR2_X1 U836 ( .A1(n1092), .A2(n1062), .ZN(n993) );
NAND2_X1 U837 ( .A1(n1152), .A2(n1153), .ZN(n1062) );
AND4_X1 U838 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NOR4_X1 U839 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1152) );
NOR3_X1 U840 ( .A1(n1162), .A2(n1028), .A3(n1012), .ZN(n1161) );
INV_X1 U841 ( .A(n1163), .ZN(n1160) );
NAND4_X1 U842 ( .A1(n988), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1092) );
NOR4_X1 U843 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR2_X1 U844 ( .A1(n1023), .A2(n1171), .ZN(n1170) );
NOR3_X1 U845 ( .A1(n1172), .A2(n1031), .A3(n1173), .ZN(n1169) );
INV_X1 U846 ( .A(n1112), .ZN(n1168) );
NAND3_X1 U847 ( .A1(n1174), .A2(n1175), .A3(n1004), .ZN(n1112) );
NOR2_X1 U848 ( .A1(n1176), .A2(n1177), .ZN(n1165) );
NAND3_X1 U849 ( .A1(n1178), .A2(n1175), .A3(n1174), .ZN(n988) );
XNOR2_X1 U850 ( .A(n1179), .B(KEYINPUT55), .ZN(n1104) );
XOR2_X1 U851 ( .A(KEYINPUT3), .B(n1180), .Z(n1150) );
NOR2_X1 U852 ( .A1(KEYINPUT2), .A2(n1181), .ZN(n1148) );
XNOR2_X1 U853 ( .A(n1182), .B(n1183), .ZN(n1181) );
XOR2_X1 U854 ( .A(n1184), .B(n1185), .Z(n1182) );
NOR2_X1 U855 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
XOR2_X1 U856 ( .A(KEYINPUT38), .B(n1188), .Z(n1187) );
NOR2_X1 U857 ( .A1(n1066), .A2(n1130), .ZN(n1188) );
AND2_X1 U858 ( .A1(n1066), .A2(n1130), .ZN(n1186) );
NAND2_X1 U859 ( .A1(KEYINPUT45), .A2(n1189), .ZN(n1184) );
NOR2_X1 U860 ( .A1(n990), .A2(G952), .ZN(n1093) );
XOR2_X1 U861 ( .A(n1190), .B(n1163), .Z(G48) );
NAND4_X1 U862 ( .A1(n1191), .A2(n1192), .A3(n1004), .A4(n1038), .ZN(n1163) );
XOR2_X1 U863 ( .A(G143), .B(n1159), .Z(G45) );
AND4_X1 U864 ( .A1(n1193), .A2(n1194), .A3(n1191), .A4(n1195), .ZN(n1159) );
NOR3_X1 U865 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1195) );
XOR2_X1 U866 ( .A(n1199), .B(n1200), .Z(G42) );
XOR2_X1 U867 ( .A(KEYINPUT23), .B(G140), .Z(n1200) );
NAND2_X1 U868 ( .A1(KEYINPUT17), .A2(n1158), .ZN(n1199) );
NOR4_X1 U869 ( .A1(n1162), .A2(n1012), .A3(n1038), .A4(n1175), .ZN(n1158) );
INV_X1 U870 ( .A(n1201), .ZN(n1162) );
XOR2_X1 U871 ( .A(n1157), .B(n1202), .Z(G39) );
NAND2_X1 U872 ( .A1(KEYINPUT33), .A2(G137), .ZN(n1202) );
NAND3_X1 U873 ( .A1(n1203), .A2(n1038), .A3(n1201), .ZN(n1157) );
XNOR2_X1 U874 ( .A(G134), .B(n1156), .ZN(G36) );
NAND3_X1 U875 ( .A1(n1193), .A2(n1178), .A3(n1201), .ZN(n1156) );
XOR2_X1 U876 ( .A(n1204), .B(n1205), .Z(G33) );
NAND4_X1 U877 ( .A1(KEYINPUT57), .A2(n1201), .A3(n1004), .A4(n1193), .ZN(n1205) );
NOR3_X1 U878 ( .A1(n1003), .A2(n1197), .A3(n1015), .ZN(n1201) );
INV_X1 U879 ( .A(n1191), .ZN(n1015) );
XNOR2_X1 U880 ( .A(n1206), .B(KEYINPUT26), .ZN(n1191) );
INV_X1 U881 ( .A(n1008), .ZN(n1003) );
NOR2_X1 U882 ( .A1(n1207), .A2(n1025), .ZN(n1008) );
XOR2_X1 U883 ( .A(n1208), .B(n1155), .Z(G30) );
NAND4_X1 U884 ( .A1(n1192), .A2(n1178), .A3(n1206), .A4(n1038), .ZN(n1155) );
INV_X1 U885 ( .A(n1010), .ZN(n1178) );
XOR2_X1 U886 ( .A(G101), .B(n1209), .Z(G3) );
NOR2_X1 U887 ( .A1(n1023), .A2(n1210), .ZN(n1209) );
XNOR2_X1 U888 ( .A(KEYINPUT58), .B(n1171), .ZN(n1210) );
NAND4_X1 U889 ( .A1(n1193), .A2(n1013), .A3(n1206), .A4(n1211), .ZN(n1171) );
INV_X1 U890 ( .A(n1028), .ZN(n1193) );
XOR2_X1 U891 ( .A(n1066), .B(n1154), .Z(G27) );
NAND4_X1 U892 ( .A1(n1192), .A2(n1004), .A3(n1031), .A4(n1005), .ZN(n1154) );
INV_X1 U893 ( .A(n1012), .ZN(n1004) );
NOR3_X1 U894 ( .A1(n1023), .A2(n1197), .A3(n1175), .ZN(n1192) );
AND2_X1 U895 ( .A1(n1212), .A2(n1213), .ZN(n1197) );
NAND2_X1 U896 ( .A1(n1214), .A2(n1061), .ZN(n1213) );
INV_X1 U897 ( .A(G900), .ZN(n1061) );
INV_X1 U898 ( .A(G125), .ZN(n1066) );
XNOR2_X1 U899 ( .A(G122), .B(n1164), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1215), .A2(n1001), .A3(n1040), .A4(n1216), .ZN(n1164) );
NOR2_X1 U901 ( .A1(n1038), .A2(n1030), .ZN(n1001) );
INV_X1 U902 ( .A(n1173), .ZN(n1215) );
XNOR2_X1 U903 ( .A(G119), .B(n1217), .ZN(G21) );
NAND3_X1 U904 ( .A1(n1218), .A2(n1203), .A3(n1219), .ZN(n1217) );
AND3_X1 U905 ( .A1(n1005), .A2(n1211), .A3(n1038), .ZN(n1219) );
XOR2_X1 U906 ( .A(n1023), .B(KEYINPUT6), .Z(n1218) );
INV_X1 U907 ( .A(n1194), .ZN(n1023) );
XOR2_X1 U908 ( .A(G116), .B(n1167), .Z(G18) );
NOR3_X1 U909 ( .A1(n1173), .A2(n1010), .A3(n1028), .ZN(n1167) );
NAND2_X1 U910 ( .A1(n1198), .A2(n1040), .ZN(n1010) );
XOR2_X1 U911 ( .A(G113), .B(n1177), .Z(G15) );
NOR3_X1 U912 ( .A1(n1028), .A2(n1173), .A3(n1012), .ZN(n1177) );
NAND2_X1 U913 ( .A1(n1196), .A2(n1216), .ZN(n1012) );
NAND3_X1 U914 ( .A1(n1194), .A2(n1211), .A3(n1005), .ZN(n1173) );
INV_X1 U915 ( .A(n1039), .ZN(n1005) );
NAND2_X1 U916 ( .A1(n1018), .A2(n1220), .ZN(n1039) );
NAND2_X1 U917 ( .A1(n1038), .A2(n1175), .ZN(n1028) );
INV_X1 U918 ( .A(n1030), .ZN(n1175) );
INV_X1 U919 ( .A(n1031), .ZN(n1038) );
XOR2_X1 U920 ( .A(G110), .B(n1176), .Z(G12) );
AND2_X1 U921 ( .A1(n1203), .A2(n1174), .ZN(n1176) );
AND4_X1 U922 ( .A1(n1194), .A2(n1206), .A3(n1031), .A4(n1211), .ZN(n1174) );
NAND2_X1 U923 ( .A1(n1212), .A2(n1221), .ZN(n1211) );
NAND2_X1 U924 ( .A1(n1214), .A2(n1081), .ZN(n1221) );
INV_X1 U925 ( .A(G898), .ZN(n1081) );
AND3_X1 U926 ( .A1(G902), .A2(n1032), .A3(G953), .ZN(n1214) );
NAND3_X1 U927 ( .A1(n1032), .A2(n990), .A3(G952), .ZN(n1212) );
NAND2_X1 U928 ( .A1(G237), .A2(G234), .ZN(n1032) );
XOR2_X1 U929 ( .A(n1222), .B(G472), .Z(n1031) );
NAND2_X1 U930 ( .A1(n1223), .A2(n1179), .ZN(n1222) );
XOR2_X1 U931 ( .A(n1224), .B(n1128), .Z(n1223) );
XNOR2_X1 U932 ( .A(n1130), .B(n1131), .ZN(n1128) );
XNOR2_X1 U933 ( .A(n1121), .B(n1132), .ZN(n1224) );
XNOR2_X1 U934 ( .A(n1225), .B(G113), .ZN(n1132) );
NAND2_X1 U935 ( .A1(KEYINPUT8), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U936 ( .A(n1227), .B(G101), .ZN(n1121) );
NAND2_X1 U937 ( .A1(n1228), .A2(G210), .ZN(n1227) );
NOR2_X1 U938 ( .A1(n1018), .A2(n1017), .ZN(n1206) );
INV_X1 U939 ( .A(n1220), .ZN(n1017) );
NAND2_X1 U940 ( .A1(G221), .A2(n1229), .ZN(n1220) );
XOR2_X1 U941 ( .A(n1230), .B(G469), .Z(n1018) );
NAND2_X1 U942 ( .A1(n1231), .A2(n1179), .ZN(n1230) );
XOR2_X1 U943 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U944 ( .A(n1234), .B(n1131), .ZN(n1233) );
XNOR2_X1 U945 ( .A(n1073), .B(n1235), .ZN(n1131) );
INV_X1 U946 ( .A(n1072), .ZN(n1235) );
XNOR2_X1 U947 ( .A(G134), .B(G137), .ZN(n1072) );
XOR2_X1 U948 ( .A(n1204), .B(KEYINPUT34), .Z(n1073) );
NAND2_X1 U949 ( .A1(KEYINPUT18), .A2(n1236), .ZN(n1234) );
XOR2_X1 U950 ( .A(n1146), .B(n1237), .Z(n1232) );
NOR2_X1 U951 ( .A1(KEYINPUT5), .A2(n1138), .ZN(n1237) );
XOR2_X1 U952 ( .A(n1069), .B(n1238), .Z(n1138) );
XNOR2_X1 U953 ( .A(n1239), .B(n1240), .ZN(n1238) );
NAND2_X1 U954 ( .A1(KEYINPUT46), .A2(n1111), .ZN(n1239) );
XNOR2_X1 U955 ( .A(n1241), .B(n1242), .ZN(n1069) );
NAND2_X1 U956 ( .A1(KEYINPUT10), .A2(n1243), .ZN(n1241) );
XOR2_X1 U957 ( .A(KEYINPUT63), .B(G146), .Z(n1243) );
NAND2_X1 U958 ( .A1(G227), .A2(n990), .ZN(n1146) );
NOR2_X1 U959 ( .A1(n1026), .A2(n1025), .ZN(n1194) );
NOR2_X1 U960 ( .A1(n1244), .A2(n1180), .ZN(n1025) );
INV_X1 U961 ( .A(G214), .ZN(n1244) );
INV_X1 U962 ( .A(n1207), .ZN(n1026) );
XNOR2_X1 U963 ( .A(n1245), .B(n1246), .ZN(n1207) );
NOR2_X1 U964 ( .A1(n1180), .A2(n1151), .ZN(n1246) );
INV_X1 U965 ( .A(G210), .ZN(n1151) );
NOR2_X1 U966 ( .A1(G237), .A2(G902), .ZN(n1180) );
NAND2_X1 U967 ( .A1(n1247), .A2(n1179), .ZN(n1245) );
XOR2_X1 U968 ( .A(KEYINPUT44), .B(n1248), .Z(n1247) );
NOR2_X1 U969 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XOR2_X1 U970 ( .A(n1251), .B(KEYINPUT21), .Z(n1250) );
NAND2_X1 U971 ( .A1(n1183), .A2(n1252), .ZN(n1251) );
NOR2_X1 U972 ( .A1(n1183), .A2(n1252), .ZN(n1249) );
XNOR2_X1 U973 ( .A(n1253), .B(n1254), .ZN(n1252) );
XOR2_X1 U974 ( .A(KEYINPUT1), .B(G125), .Z(n1254) );
XOR2_X1 U975 ( .A(n1130), .B(n1189), .Z(n1253) );
AND2_X1 U976 ( .A1(G224), .A2(n990), .ZN(n1189) );
NAND2_X1 U977 ( .A1(n1255), .A2(n1256), .ZN(n1130) );
NAND2_X1 U978 ( .A1(G146), .A2(n1257), .ZN(n1256) );
NAND2_X1 U979 ( .A1(n1258), .A2(n1190), .ZN(n1255) );
INV_X1 U980 ( .A(G146), .ZN(n1190) );
XOR2_X1 U981 ( .A(KEYINPUT29), .B(n1242), .Z(n1258) );
XOR2_X1 U982 ( .A(n1259), .B(n1083), .Z(n1183) );
XOR2_X1 U983 ( .A(G110), .B(G122), .Z(n1083) );
NAND3_X1 U984 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1259) );
NAND2_X1 U985 ( .A1(KEYINPUT35), .A2(n1263), .ZN(n1262) );
OR3_X1 U986 ( .A1(n1263), .A2(KEYINPUT35), .A3(n1087), .ZN(n1261) );
NAND2_X1 U987 ( .A1(n1087), .A2(n1264), .ZN(n1260) );
NAND2_X1 U988 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
INV_X1 U989 ( .A(KEYINPUT35), .ZN(n1266) );
XNOR2_X1 U990 ( .A(KEYINPUT20), .B(n1263), .ZN(n1265) );
XNOR2_X1 U991 ( .A(n1088), .B(KEYINPUT13), .ZN(n1263) );
XOR2_X1 U992 ( .A(n1226), .B(G113), .Z(n1088) );
XOR2_X1 U993 ( .A(G116), .B(n1267), .Z(n1226) );
XOR2_X1 U994 ( .A(KEYINPUT7), .B(G119), .Z(n1267) );
XNOR2_X1 U995 ( .A(n1111), .B(n1240), .ZN(n1087) );
XOR2_X1 U996 ( .A(G101), .B(G107), .Z(n1240) );
INV_X1 U997 ( .A(n1172), .ZN(n1203) );
NAND2_X1 U998 ( .A1(n1013), .A2(n1030), .ZN(n1172) );
XOR2_X1 U999 ( .A(n1042), .B(n1268), .Z(n1030) );
NOR2_X1 U1000 ( .A1(n1041), .A2(KEYINPUT36), .ZN(n1268) );
NOR2_X1 U1001 ( .A1(n1095), .A2(G902), .ZN(n1041) );
XOR2_X1 U1002 ( .A(n1269), .B(n1270), .Z(n1095) );
XOR2_X1 U1003 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U1004 ( .A(KEYINPUT47), .B(KEYINPUT14), .Z(n1272) );
NOR2_X1 U1005 ( .A1(KEYINPUT51), .A2(n1273), .ZN(n1271) );
XOR2_X1 U1006 ( .A(G119), .B(n1274), .Z(n1273) );
XOR2_X1 U1007 ( .A(KEYINPUT19), .B(G128), .Z(n1274) );
XOR2_X1 U1008 ( .A(n1275), .B(n1276), .Z(n1269) );
XNOR2_X1 U1009 ( .A(n1277), .B(n1236), .ZN(n1275) );
XOR2_X1 U1010 ( .A(G110), .B(n1074), .Z(n1236) );
INV_X1 U1011 ( .A(G140), .ZN(n1074) );
NAND2_X1 U1012 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
OR2_X1 U1013 ( .A1(n1280), .A2(KEYINPUT27), .ZN(n1279) );
XOR2_X1 U1014 ( .A(n1281), .B(n1282), .Z(n1278) );
AND2_X1 U1015 ( .A1(G221), .A2(n1283), .ZN(n1282) );
NAND2_X1 U1016 ( .A1(KEYINPUT27), .A2(n1280), .ZN(n1281) );
XOR2_X1 U1017 ( .A(G137), .B(KEYINPUT52), .Z(n1280) );
NAND2_X1 U1018 ( .A1(G217), .A2(n1229), .ZN(n1042) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1179), .ZN(n1229) );
NOR2_X1 U1020 ( .A1(n1040), .A2(n1216), .ZN(n1013) );
INV_X1 U1021 ( .A(n1198), .ZN(n1216) );
XOR2_X1 U1022 ( .A(n1284), .B(G475), .Z(n1198) );
NAND2_X1 U1023 ( .A1(KEYINPUT16), .A2(n1046), .ZN(n1284) );
NOR2_X1 U1024 ( .A1(n1109), .A2(G902), .ZN(n1046) );
XNOR2_X1 U1025 ( .A(n1285), .B(n1286), .ZN(n1109) );
XOR2_X1 U1026 ( .A(G122), .B(G113), .Z(n1286) );
XOR2_X1 U1027 ( .A(n1111), .B(n1287), .Z(n1285) );
NOR2_X1 U1028 ( .A1(KEYINPUT31), .A2(n1288), .ZN(n1287) );
XOR2_X1 U1029 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U1030 ( .A(G143), .B(n1291), .Z(n1290) );
NOR2_X1 U1031 ( .A1(KEYINPUT42), .A2(n1204), .ZN(n1291) );
INV_X1 U1032 ( .A(G131), .ZN(n1204) );
XOR2_X1 U1033 ( .A(n1292), .B(n1293), .Z(n1289) );
NOR2_X1 U1034 ( .A1(KEYINPUT24), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1035 ( .A(n1276), .B(n1295), .Z(n1294) );
XOR2_X1 U1036 ( .A(KEYINPUT53), .B(G140), .Z(n1295) );
XOR2_X1 U1037 ( .A(G146), .B(G125), .Z(n1276) );
NAND2_X1 U1038 ( .A1(n1228), .A2(G214), .ZN(n1292) );
NOR2_X1 U1039 ( .A1(G953), .A2(G237), .ZN(n1228) );
INV_X1 U1040 ( .A(G104), .ZN(n1111) );
INV_X1 U1041 ( .A(n1196), .ZN(n1040) );
XOR2_X1 U1042 ( .A(n1296), .B(G478), .Z(n1196) );
NAND2_X1 U1043 ( .A1(n1100), .A2(n1179), .ZN(n1296) );
INV_X1 U1044 ( .A(G902), .ZN(n1179) );
XNOR2_X1 U1045 ( .A(n1297), .B(n1298), .ZN(n1100) );
XOR2_X1 U1046 ( .A(n1299), .B(n1300), .Z(n1298) );
XOR2_X1 U1047 ( .A(n1301), .B(G107), .Z(n1300) );
NAND2_X1 U1048 ( .A1(G217), .A2(n1283), .ZN(n1301) );
AND2_X1 U1049 ( .A1(G234), .A2(n990), .ZN(n1283) );
INV_X1 U1050 ( .A(G953), .ZN(n990) );
NAND2_X1 U1051 ( .A1(KEYINPUT15), .A2(n1242), .ZN(n1299) );
INV_X1 U1052 ( .A(n1257), .ZN(n1242) );
XOR2_X1 U1053 ( .A(n1208), .B(G143), .Z(n1257) );
INV_X1 U1054 ( .A(G128), .ZN(n1208) );
XNOR2_X1 U1055 ( .A(G116), .B(n1302), .ZN(n1297) );
XOR2_X1 U1056 ( .A(G134), .B(G122), .Z(n1302) );
endmodule


