//Key = 1110111100100100001001101100100001001010000000001010010010010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424;

XOR2_X1 U794 ( .A(G107), .B(n1094), .Z(G9) );
NOR2_X1 U795 ( .A1(n1095), .A2(n1096), .ZN(G75) );
NOR4_X1 U796 ( .A1(n1097), .A2(n1098), .A3(G953), .A4(n1099), .ZN(n1096) );
NOR4_X1 U797 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1098) );
NOR2_X1 U798 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
NOR2_X1 U799 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U800 ( .A(n1108), .B(KEYINPUT11), .ZN(n1106) );
NOR4_X1 U801 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1104) );
INV_X1 U802 ( .A(n1113), .ZN(n1110) );
NAND3_X1 U803 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1097) );
NAND3_X1 U804 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1115) );
NAND2_X1 U805 ( .A1(n1120), .A2(n1103), .ZN(n1118) );
OR4_X1 U806 ( .A1(n1101), .A2(n1121), .A3(n1111), .A4(KEYINPUT53), .ZN(n1120) );
NAND3_X1 U807 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1117) );
INV_X1 U808 ( .A(n1103), .ZN(n1124) );
NAND3_X1 U809 ( .A1(n1108), .A2(n1125), .A3(n1126), .ZN(n1123) );
NAND2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NAND2_X1 U811 ( .A1(KEYINPUT53), .A2(n1129), .ZN(n1128) );
NAND2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1122) );
NAND2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U814 ( .A1(n1108), .A2(n1134), .ZN(n1133) );
NAND2_X1 U815 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND3_X1 U816 ( .A1(n1137), .A2(n1138), .A3(KEYINPUT36), .ZN(n1136) );
NAND2_X1 U817 ( .A1(n1126), .A2(n1139), .ZN(n1132) );
NAND3_X1 U818 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
OR2_X1 U819 ( .A1(n1111), .A2(KEYINPUT36), .ZN(n1142) );
NOR3_X1 U820 ( .A1(n1099), .A2(G953), .A3(G952), .ZN(n1095) );
AND4_X1 U821 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1099) );
NOR4_X1 U822 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
NOR2_X1 U823 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XNOR2_X1 U824 ( .A(G472), .B(KEYINPUT46), .ZN(n1152) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1149) );
INV_X1 U826 ( .A(n1155), .ZN(n1154) );
XOR2_X1 U827 ( .A(n1156), .B(KEYINPUT48), .Z(n1153) );
XNOR2_X1 U828 ( .A(n1157), .B(n1158), .ZN(n1145) );
XNOR2_X1 U829 ( .A(KEYINPUT30), .B(n1159), .ZN(n1158) );
XOR2_X1 U830 ( .A(KEYINPUT29), .B(n1160), .Z(n1144) );
AND4_X1 U831 ( .A1(n1161), .A2(n1162), .A3(n1112), .A4(n1126), .ZN(n1160) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(G72) );
XOR2_X1 U833 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U834 ( .A1(n1114), .A2(G953), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1165) );
XOR2_X1 U836 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U837 ( .A(G131), .B(n1171), .ZN(n1170) );
XNOR2_X1 U838 ( .A(KEYINPUT18), .B(KEYINPUT16), .ZN(n1171) );
XOR2_X1 U839 ( .A(n1172), .B(n1173), .Z(n1169) );
XOR2_X1 U840 ( .A(n1174), .B(n1175), .Z(n1172) );
NAND2_X1 U841 ( .A1(n1176), .A2(KEYINPUT25), .ZN(n1174) );
XNOR2_X1 U842 ( .A(n1177), .B(n1178), .ZN(n1176) );
NAND2_X1 U843 ( .A1(KEYINPUT1), .A2(G140), .ZN(n1177) );
NOR2_X1 U844 ( .A1(n1179), .A2(n1180), .ZN(n1163) );
AND2_X1 U845 ( .A1(G227), .A2(G900), .ZN(n1179) );
XOR2_X1 U846 ( .A(n1181), .B(n1182), .Z(G69) );
NOR2_X1 U847 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U848 ( .A(n1185), .B(KEYINPUT10), .Z(n1184) );
NAND3_X1 U849 ( .A1(n1186), .A2(n1180), .A3(n1187), .ZN(n1185) );
NOR2_X1 U850 ( .A1(n1188), .A2(n1187), .ZN(n1183) );
NAND2_X1 U851 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
NAND2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U853 ( .A(n1193), .B(n1194), .Z(n1189) );
NOR2_X1 U854 ( .A1(KEYINPUT34), .A2(n1195), .ZN(n1193) );
NOR2_X1 U855 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U856 ( .A(n1198), .B(KEYINPUT28), .Z(n1197) );
NAND2_X1 U857 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NOR2_X1 U858 ( .A1(n1199), .A2(n1200), .ZN(n1196) );
XNOR2_X1 U859 ( .A(n1201), .B(KEYINPUT50), .ZN(n1199) );
NOR2_X1 U860 ( .A1(G953), .A2(n1116), .ZN(n1188) );
NAND2_X1 U861 ( .A1(G953), .A2(n1202), .ZN(n1181) );
NAND2_X1 U862 ( .A1(G224), .A2(G898), .ZN(n1202) );
NOR2_X1 U863 ( .A1(n1203), .A2(n1204), .ZN(G66) );
NOR2_X1 U864 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U865 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U866 ( .A1(n1156), .A2(n1209), .ZN(n1208) );
NOR2_X1 U867 ( .A1(KEYINPUT42), .A2(n1210), .ZN(n1207) );
AND2_X1 U868 ( .A1(n1210), .A2(KEYINPUT42), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1203), .A2(n1211), .ZN(G63) );
XNOR2_X1 U870 ( .A(n1212), .B(n1213), .ZN(n1211) );
NOR2_X1 U871 ( .A1(n1214), .A2(n1209), .ZN(n1213) );
NOR2_X1 U872 ( .A1(n1203), .A2(n1215), .ZN(G60) );
NOR3_X1 U873 ( .A1(n1157), .A2(n1216), .A3(n1217), .ZN(n1215) );
NOR3_X1 U874 ( .A1(n1218), .A2(n1159), .A3(n1209), .ZN(n1217) );
INV_X1 U875 ( .A(G475), .ZN(n1159) );
NOR2_X1 U876 ( .A1(n1219), .A2(n1220), .ZN(n1216) );
AND2_X1 U877 ( .A1(n1221), .A2(G475), .ZN(n1219) );
XNOR2_X1 U878 ( .A(n1222), .B(n1223), .ZN(G6) );
NOR3_X1 U879 ( .A1(n1224), .A2(n1127), .A3(n1225), .ZN(n1223) );
XNOR2_X1 U880 ( .A(KEYINPUT62), .B(n1107), .ZN(n1225) );
NAND3_X1 U881 ( .A1(n1226), .A2(n1227), .A3(n1108), .ZN(n1224) );
NOR2_X1 U882 ( .A1(n1203), .A2(n1228), .ZN(G57) );
XOR2_X1 U883 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U884 ( .A(n1231), .B(n1232), .Z(n1230) );
NAND2_X1 U885 ( .A1(KEYINPUT2), .A2(n1233), .ZN(n1231) );
XNOR2_X1 U886 ( .A(n1234), .B(n1235), .ZN(n1233) );
NOR2_X1 U887 ( .A1(n1236), .A2(KEYINPUT20), .ZN(n1235) );
XOR2_X1 U888 ( .A(n1237), .B(n1238), .Z(n1229) );
NOR2_X1 U889 ( .A1(n1239), .A2(n1209), .ZN(n1238) );
NOR2_X1 U890 ( .A1(KEYINPUT32), .A2(n1240), .ZN(n1237) );
NOR2_X1 U891 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U892 ( .A(n1243), .B(KEYINPUT61), .Z(n1242) );
INV_X1 U893 ( .A(n1244), .ZN(n1241) );
NOR2_X1 U894 ( .A1(n1203), .A2(n1245), .ZN(G54) );
XOR2_X1 U895 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U896 ( .A(G110), .B(n1248), .Z(n1247) );
NOR2_X1 U897 ( .A1(n1249), .A2(n1209), .ZN(n1248) );
XOR2_X1 U898 ( .A(n1250), .B(n1251), .Z(n1246) );
NAND2_X1 U899 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
NAND2_X1 U900 ( .A1(n1201), .A2(n1254), .ZN(n1253) );
NAND2_X1 U901 ( .A1(n1255), .A2(n1256), .ZN(n1252) );
XNOR2_X1 U902 ( .A(KEYINPUT45), .B(n1254), .ZN(n1255) );
NOR2_X1 U903 ( .A1(n1203), .A2(n1257), .ZN(G51) );
XOR2_X1 U904 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U905 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U906 ( .A1(n1262), .A2(n1209), .ZN(n1261) );
NAND2_X1 U907 ( .A1(G902), .A2(n1221), .ZN(n1209) );
NAND2_X1 U908 ( .A1(n1116), .A2(n1263), .ZN(n1221) );
XOR2_X1 U909 ( .A(KEYINPUT60), .B(n1114), .Z(n1263) );
AND4_X1 U910 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1114) );
NOR4_X1 U911 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1267) );
AND2_X1 U912 ( .A1(n1272), .A2(n1273), .ZN(n1266) );
NAND4_X1 U913 ( .A1(n1274), .A2(n1275), .A3(n1126), .A4(n1276), .ZN(n1265) );
NOR2_X1 U914 ( .A1(n1141), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U915 ( .A(KEYINPUT0), .B(n1107), .ZN(n1277) );
INV_X1 U916 ( .A(n1278), .ZN(n1141) );
XNOR2_X1 U917 ( .A(KEYINPUT23), .B(n1127), .ZN(n1274) );
NAND2_X1 U918 ( .A1(n1119), .A2(n1279), .ZN(n1264) );
XOR2_X1 U919 ( .A(KEYINPUT35), .B(n1280), .Z(n1279) );
INV_X1 U920 ( .A(n1186), .ZN(n1116) );
NAND4_X1 U921 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1186) );
NOR4_X1 U922 ( .A1(n1285), .A2(n1286), .A3(n1287), .A4(n1094), .ZN(n1284) );
AND3_X1 U923 ( .A1(n1129), .A2(n1108), .A3(n1288), .ZN(n1094) );
NOR2_X1 U924 ( .A1(n1289), .A2(n1290), .ZN(n1283) );
NAND4_X1 U925 ( .A1(n1291), .A2(n1129), .A3(n1292), .A4(n1293), .ZN(n1282) );
NAND2_X1 U926 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
INV_X1 U927 ( .A(KEYINPUT8), .ZN(n1295) );
NAND2_X1 U928 ( .A1(KEYINPUT8), .A2(n1296), .ZN(n1292) );
NAND3_X1 U929 ( .A1(n1126), .A2(n1297), .A3(n1298), .ZN(n1296) );
NAND3_X1 U930 ( .A1(n1288), .A2(n1108), .A3(n1299), .ZN(n1281) );
INV_X1 U931 ( .A(n1111), .ZN(n1108) );
INV_X1 U932 ( .A(G210), .ZN(n1262) );
NOR2_X1 U933 ( .A1(KEYINPUT40), .A2(n1300), .ZN(n1260) );
XNOR2_X1 U934 ( .A(n1301), .B(n1302), .ZN(n1300) );
NOR2_X1 U935 ( .A1(n1180), .A2(G952), .ZN(n1203) );
XNOR2_X1 U936 ( .A(G146), .B(n1273), .ZN(G48) );
NAND3_X1 U937 ( .A1(n1299), .A2(n1297), .A3(n1303), .ZN(n1273) );
NAND2_X1 U938 ( .A1(n1304), .A2(n1305), .ZN(G45) );
NAND2_X1 U939 ( .A1(G143), .A2(n1272), .ZN(n1305) );
XOR2_X1 U940 ( .A(KEYINPUT33), .B(n1306), .Z(n1304) );
NOR2_X1 U941 ( .A1(G143), .A2(n1272), .ZN(n1306) );
NAND4_X1 U942 ( .A1(n1307), .A2(n1275), .A3(n1297), .A4(n1308), .ZN(n1272) );
NOR3_X1 U943 ( .A1(n1140), .A2(n1135), .A3(n1309), .ZN(n1308) );
XNOR2_X1 U944 ( .A(n1310), .B(n1271), .ZN(G42) );
AND3_X1 U945 ( .A1(n1299), .A2(n1278), .A3(n1311), .ZN(n1271) );
XNOR2_X1 U946 ( .A(G137), .B(n1312), .ZN(G39) );
NAND3_X1 U947 ( .A1(n1280), .A2(n1119), .A3(KEYINPUT59), .ZN(n1312) );
AND2_X1 U948 ( .A1(n1303), .A2(n1130), .ZN(n1280) );
XOR2_X1 U949 ( .A(G134), .B(n1270), .Z(G36) );
AND3_X1 U950 ( .A1(n1291), .A2(n1129), .A3(n1311), .ZN(n1270) );
XNOR2_X1 U951 ( .A(n1313), .B(n1269), .ZN(G33) );
AND3_X1 U952 ( .A1(n1299), .A2(n1291), .A3(n1311), .ZN(n1269) );
AND3_X1 U953 ( .A1(n1226), .A2(n1275), .A3(n1119), .ZN(n1311) );
AND3_X1 U954 ( .A1(n1112), .A2(n1162), .A3(n1113), .ZN(n1119) );
XOR2_X1 U955 ( .A(G128), .B(n1268), .Z(G30) );
AND3_X1 U956 ( .A1(n1129), .A2(n1297), .A3(n1303), .ZN(n1268) );
NOR4_X1 U957 ( .A1(n1135), .A2(n1314), .A3(n1315), .A4(n1316), .ZN(n1303) );
XNOR2_X1 U958 ( .A(n1317), .B(n1287), .ZN(G3) );
AND3_X1 U959 ( .A1(n1130), .A2(n1288), .A3(n1291), .ZN(n1287) );
INV_X1 U960 ( .A(n1140), .ZN(n1291) );
XNOR2_X1 U961 ( .A(G125), .B(n1318), .ZN(G27) );
NAND4_X1 U962 ( .A1(n1299), .A2(n1126), .A3(n1319), .A4(n1297), .ZN(n1318) );
NOR2_X1 U963 ( .A1(n1314), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U964 ( .A(n1278), .B(KEYINPUT37), .ZN(n1320) );
INV_X1 U965 ( .A(n1275), .ZN(n1314) );
NAND2_X1 U966 ( .A1(n1103), .A2(n1321), .ZN(n1275) );
NAND3_X1 U967 ( .A1(G902), .A2(n1322), .A3(n1167), .ZN(n1321) );
NOR2_X1 U968 ( .A1(n1323), .A2(G900), .ZN(n1167) );
XOR2_X1 U969 ( .A(G122), .B(n1290), .Z(G24) );
NOR4_X1 U970 ( .A1(n1309), .A2(n1294), .A3(n1111), .A4(n1143), .ZN(n1290) );
NAND2_X1 U971 ( .A1(n1316), .A2(n1315), .ZN(n1111) );
XNOR2_X1 U972 ( .A(n1324), .B(n1289), .ZN(G21) );
NOR4_X1 U973 ( .A1(n1294), .A2(n1102), .A3(n1315), .A4(n1316), .ZN(n1289) );
INV_X1 U974 ( .A(n1130), .ZN(n1102) );
XOR2_X1 U975 ( .A(G116), .B(n1325), .Z(G18) );
NOR4_X1 U976 ( .A1(KEYINPUT27), .A2(n1121), .A3(n1140), .A4(n1294), .ZN(n1325) );
INV_X1 U977 ( .A(n1129), .ZN(n1121) );
NOR2_X1 U978 ( .A1(n1326), .A2(n1143), .ZN(n1129) );
INV_X1 U979 ( .A(n1307), .ZN(n1143) );
XOR2_X1 U980 ( .A(n1327), .B(n1286), .Z(G15) );
NOR3_X1 U981 ( .A1(n1294), .A2(n1140), .A3(n1127), .ZN(n1286) );
INV_X1 U982 ( .A(n1299), .ZN(n1127) );
NOR2_X1 U983 ( .A1(n1309), .A2(n1307), .ZN(n1299) );
NAND2_X1 U984 ( .A1(n1315), .A2(n1328), .ZN(n1140) );
XOR2_X1 U985 ( .A(KEYINPUT7), .B(n1316), .Z(n1328) );
NAND3_X1 U986 ( .A1(n1297), .A2(n1227), .A3(n1126), .ZN(n1294) );
INV_X1 U987 ( .A(n1101), .ZN(n1126) );
NAND2_X1 U988 ( .A1(n1137), .A2(n1329), .ZN(n1101) );
INV_X1 U989 ( .A(n1107), .ZN(n1297) );
NAND2_X1 U990 ( .A1(KEYINPUT5), .A2(n1330), .ZN(n1327) );
XOR2_X1 U991 ( .A(G110), .B(n1285), .Z(G12) );
AND3_X1 U992 ( .A1(n1278), .A2(n1288), .A3(n1130), .ZN(n1285) );
NOR2_X1 U993 ( .A1(n1307), .A2(n1326), .ZN(n1130) );
INV_X1 U994 ( .A(n1309), .ZN(n1326) );
XOR2_X1 U995 ( .A(G475), .B(n1331), .Z(n1309) );
NOR2_X1 U996 ( .A1(n1157), .A2(KEYINPUT17), .ZN(n1331) );
NOR2_X1 U997 ( .A1(n1220), .A2(G902), .ZN(n1157) );
INV_X1 U998 ( .A(n1218), .ZN(n1220) );
XNOR2_X1 U999 ( .A(n1332), .B(n1333), .ZN(n1218) );
XNOR2_X1 U1000 ( .A(n1334), .B(n1335), .ZN(n1333) );
NOR2_X1 U1001 ( .A1(KEYINPUT54), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1002 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1003 ( .A(n1339), .B(n1340), .Z(n1338) );
AND3_X1 U1004 ( .A1(n1341), .A2(G214), .A3(n1342), .ZN(n1339) );
XOR2_X1 U1005 ( .A(n1343), .B(n1344), .Z(n1337) );
XNOR2_X1 U1006 ( .A(n1313), .B(G125), .ZN(n1344) );
INV_X1 U1007 ( .A(G131), .ZN(n1313) );
NAND2_X1 U1008 ( .A1(KEYINPUT63), .A2(n1345), .ZN(n1343) );
NAND2_X1 U1009 ( .A1(KEYINPUT22), .A2(n1222), .ZN(n1334) );
XNOR2_X1 U1010 ( .A(G113), .B(G122), .ZN(n1332) );
XOR2_X1 U1011 ( .A(n1346), .B(n1214), .Z(n1307) );
INV_X1 U1012 ( .A(G478), .ZN(n1214) );
NAND2_X1 U1013 ( .A1(n1212), .A2(n1347), .ZN(n1346) );
XNOR2_X1 U1014 ( .A(n1348), .B(n1349), .ZN(n1212) );
XNOR2_X1 U1015 ( .A(n1350), .B(n1351), .ZN(n1349) );
XOR2_X1 U1016 ( .A(n1352), .B(n1353), .Z(n1351) );
AND3_X1 U1017 ( .A1(G217), .A2(G234), .A3(n1342), .ZN(n1353) );
NAND2_X1 U1018 ( .A1(KEYINPUT38), .A2(G128), .ZN(n1352) );
XOR2_X1 U1019 ( .A(n1354), .B(n1355), .Z(n1348) );
XNOR2_X1 U1020 ( .A(n1356), .B(G122), .ZN(n1355) );
INV_X1 U1021 ( .A(G143), .ZN(n1356) );
XNOR2_X1 U1022 ( .A(G107), .B(G116), .ZN(n1354) );
NOR3_X1 U1023 ( .A1(n1107), .A2(n1298), .A3(n1135), .ZN(n1288) );
INV_X1 U1024 ( .A(n1226), .ZN(n1135) );
NOR2_X1 U1025 ( .A1(n1137), .A2(n1138), .ZN(n1226) );
INV_X1 U1026 ( .A(n1329), .ZN(n1138) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1357), .ZN(n1329) );
XNOR2_X1 U1028 ( .A(n1358), .B(n1249), .ZN(n1137) );
INV_X1 U1029 ( .A(G469), .ZN(n1249) );
NAND2_X1 U1030 ( .A1(n1359), .A2(n1347), .ZN(n1358) );
XOR2_X1 U1031 ( .A(n1360), .B(n1361), .Z(n1359) );
XNOR2_X1 U1032 ( .A(n1254), .B(n1251), .ZN(n1361) );
XOR2_X1 U1033 ( .A(G140), .B(n1362), .Z(n1251) );
AND2_X1 U1034 ( .A1(n1342), .A2(G227), .ZN(n1362) );
XOR2_X1 U1035 ( .A(n1234), .B(n1173), .Z(n1254) );
XNOR2_X1 U1036 ( .A(n1363), .B(n1364), .ZN(n1173) );
NOR2_X1 U1037 ( .A1(G146), .A2(KEYINPUT15), .ZN(n1364) );
XNOR2_X1 U1038 ( .A(G143), .B(G128), .ZN(n1363) );
XNOR2_X1 U1039 ( .A(n1365), .B(n1256), .ZN(n1360) );
INV_X1 U1040 ( .A(n1201), .ZN(n1256) );
NOR2_X1 U1041 ( .A1(G110), .A2(KEYINPUT47), .ZN(n1365) );
INV_X1 U1042 ( .A(n1227), .ZN(n1298) );
NAND2_X1 U1043 ( .A1(n1103), .A2(n1366), .ZN(n1227) );
NAND4_X1 U1044 ( .A1(G902), .A2(n1191), .A3(n1192), .A4(n1322), .ZN(n1366) );
INV_X1 U1045 ( .A(n1323), .ZN(n1192) );
XOR2_X1 U1046 ( .A(n1180), .B(KEYINPUT31), .Z(n1323) );
XOR2_X1 U1047 ( .A(KEYINPUT21), .B(G898), .Z(n1191) );
NAND3_X1 U1048 ( .A1(n1322), .A2(n1180), .A3(G952), .ZN(n1103) );
INV_X1 U1049 ( .A(G953), .ZN(n1180) );
NAND2_X1 U1050 ( .A1(G237), .A2(G234), .ZN(n1322) );
NAND2_X1 U1051 ( .A1(n1112), .A2(n1367), .ZN(n1107) );
NAND2_X1 U1052 ( .A1(n1113), .A2(n1162), .ZN(n1367) );
INV_X1 U1053 ( .A(n1109), .ZN(n1162) );
NOR2_X1 U1054 ( .A1(n1368), .A2(n1369), .ZN(n1109) );
AND2_X1 U1055 ( .A1(G210), .A2(n1370), .ZN(n1369) );
XNOR2_X1 U1056 ( .A(n1371), .B(KEYINPUT6), .ZN(n1113) );
NAND2_X1 U1057 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
NAND2_X1 U1058 ( .A1(KEYINPUT49), .A2(n1368), .ZN(n1373) );
NAND2_X1 U1059 ( .A1(n1161), .A2(n1374), .ZN(n1372) );
INV_X1 U1060 ( .A(KEYINPUT49), .ZN(n1374) );
NAND3_X1 U1061 ( .A1(n1370), .A2(n1368), .A3(G210), .ZN(n1161) );
NAND2_X1 U1062 ( .A1(n1375), .A2(n1347), .ZN(n1368) );
XOR2_X1 U1063 ( .A(n1376), .B(n1377), .Z(n1375) );
NOR2_X1 U1064 ( .A1(KEYINPUT14), .A2(n1258), .ZN(n1377) );
XOR2_X1 U1065 ( .A(n1378), .B(n1200), .Z(n1258) );
XNOR2_X1 U1066 ( .A(n1379), .B(G113), .ZN(n1200) );
NAND2_X1 U1067 ( .A1(n1380), .A2(KEYINPUT4), .ZN(n1379) );
XNOR2_X1 U1068 ( .A(G116), .B(n1381), .ZN(n1380) );
NOR2_X1 U1069 ( .A1(G119), .A2(KEYINPUT12), .ZN(n1381) );
XNOR2_X1 U1070 ( .A(n1201), .B(n1194), .ZN(n1378) );
XOR2_X1 U1071 ( .A(G110), .B(n1382), .Z(n1194) );
XOR2_X1 U1072 ( .A(KEYINPUT41), .B(G122), .Z(n1382) );
XOR2_X1 U1073 ( .A(G101), .B(n1383), .Z(n1201) );
XNOR2_X1 U1074 ( .A(G107), .B(n1222), .ZN(n1383) );
INV_X1 U1075 ( .A(G104), .ZN(n1222) );
NAND2_X1 U1076 ( .A1(n1384), .A2(n1385), .ZN(n1376) );
NAND3_X1 U1077 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n1385) );
OR2_X1 U1078 ( .A1(n1389), .A2(n1302), .ZN(n1387) );
NAND3_X1 U1079 ( .A1(G125), .A2(n1390), .A3(n1389), .ZN(n1386) );
XOR2_X1 U1080 ( .A(n1391), .B(KEYINPUT57), .Z(n1384) );
NAND3_X1 U1081 ( .A1(n1392), .A2(n1393), .A3(n1301), .ZN(n1391) );
INV_X1 U1082 ( .A(n1388), .ZN(n1301) );
NAND2_X1 U1083 ( .A1(G224), .A2(n1342), .ZN(n1388) );
NAND2_X1 U1084 ( .A1(n1394), .A2(n1389), .ZN(n1393) );
INV_X1 U1085 ( .A(KEYINPUT24), .ZN(n1389) );
NAND2_X1 U1086 ( .A1(G125), .A2(n1390), .ZN(n1394) );
NAND2_X1 U1087 ( .A1(KEYINPUT24), .A2(n1302), .ZN(n1392) );
XNOR2_X1 U1088 ( .A(n1236), .B(n1178), .ZN(n1302) );
INV_X1 U1089 ( .A(G125), .ZN(n1178) );
INV_X1 U1090 ( .A(n1390), .ZN(n1236) );
NAND2_X1 U1091 ( .A1(G214), .A2(n1370), .ZN(n1112) );
NAND2_X1 U1092 ( .A1(n1395), .A2(n1347), .ZN(n1370) );
XNOR2_X1 U1093 ( .A(G237), .B(KEYINPUT55), .ZN(n1395) );
NOR2_X1 U1094 ( .A1(n1396), .A2(n1315), .ZN(n1278) );
NOR2_X1 U1095 ( .A1(n1397), .A2(n1148), .ZN(n1315) );
NOR2_X1 U1096 ( .A1(n1156), .A2(n1155), .ZN(n1148) );
AND2_X1 U1097 ( .A1(n1155), .A2(n1156), .ZN(n1397) );
NAND2_X1 U1098 ( .A1(G217), .A2(n1357), .ZN(n1156) );
NAND2_X1 U1099 ( .A1(G234), .A2(n1347), .ZN(n1357) );
NOR2_X1 U1100 ( .A1(n1210), .A2(G902), .ZN(n1155) );
XOR2_X1 U1101 ( .A(n1398), .B(n1399), .Z(n1210) );
XOR2_X1 U1102 ( .A(n1400), .B(n1401), .Z(n1399) );
XNOR2_X1 U1103 ( .A(n1402), .B(n1403), .ZN(n1401) );
NOR2_X1 U1104 ( .A1(KEYINPUT52), .A2(n1324), .ZN(n1403) );
INV_X1 U1105 ( .A(G119), .ZN(n1324) );
NAND2_X1 U1106 ( .A1(KEYINPUT56), .A2(n1404), .ZN(n1402) );
XOR2_X1 U1107 ( .A(n1405), .B(n1345), .Z(n1404) );
XNOR2_X1 U1108 ( .A(n1310), .B(KEYINPUT13), .ZN(n1345) );
INV_X1 U1109 ( .A(G140), .ZN(n1310) );
NOR2_X1 U1110 ( .A1(G125), .A2(KEYINPUT58), .ZN(n1405) );
AND3_X1 U1111 ( .A1(n1342), .A2(G234), .A3(G221), .ZN(n1400) );
XOR2_X1 U1112 ( .A(n1406), .B(n1407), .Z(n1398) );
XOR2_X1 U1113 ( .A(G128), .B(G110), .Z(n1407) );
XNOR2_X1 U1114 ( .A(G137), .B(G146), .ZN(n1406) );
INV_X1 U1115 ( .A(n1316), .ZN(n1396) );
NOR2_X1 U1116 ( .A1(n1408), .A2(n1147), .ZN(n1316) );
NOR2_X1 U1117 ( .A1(n1409), .A2(G472), .ZN(n1147) );
NOR2_X1 U1118 ( .A1(n1239), .A2(n1151), .ZN(n1408) );
INV_X1 U1119 ( .A(n1409), .ZN(n1151) );
NAND2_X1 U1120 ( .A1(n1410), .A2(n1347), .ZN(n1409) );
INV_X1 U1121 ( .A(G902), .ZN(n1347) );
XOR2_X1 U1122 ( .A(n1411), .B(n1412), .Z(n1410) );
XOR2_X1 U1123 ( .A(n1413), .B(n1232), .Z(n1412) );
XOR2_X1 U1124 ( .A(n1414), .B(n1415), .Z(n1232) );
XNOR2_X1 U1125 ( .A(n1330), .B(n1416), .ZN(n1415) );
NOR2_X1 U1126 ( .A1(G119), .A2(KEYINPUT43), .ZN(n1416) );
INV_X1 U1127 ( .A(G113), .ZN(n1330) );
XNOR2_X1 U1128 ( .A(G116), .B(KEYINPUT39), .ZN(n1414) );
NAND2_X1 U1129 ( .A1(n1243), .A2(n1244), .ZN(n1413) );
NAND4_X1 U1130 ( .A1(n1341), .A2(G210), .A3(n1342), .A4(G101), .ZN(n1244) );
NAND2_X1 U1131 ( .A1(n1317), .A2(n1417), .ZN(n1243) );
NAND3_X1 U1132 ( .A1(n1342), .A2(G210), .A3(n1341), .ZN(n1417) );
XNOR2_X1 U1133 ( .A(G237), .B(KEYINPUT3), .ZN(n1341) );
XNOR2_X1 U1134 ( .A(G953), .B(KEYINPUT44), .ZN(n1342) );
INV_X1 U1135 ( .A(G101), .ZN(n1317) );
XNOR2_X1 U1136 ( .A(n1418), .B(n1390), .ZN(n1411) );
NAND2_X1 U1137 ( .A1(n1419), .A2(n1420), .ZN(n1390) );
NAND2_X1 U1138 ( .A1(G128), .A2(n1340), .ZN(n1420) );
XOR2_X1 U1139 ( .A(n1421), .B(KEYINPUT26), .Z(n1419) );
OR2_X1 U1140 ( .A1(n1340), .A2(G128), .ZN(n1421) );
XOR2_X1 U1141 ( .A(G143), .B(G146), .Z(n1340) );
XOR2_X1 U1142 ( .A(n1234), .B(KEYINPUT19), .Z(n1418) );
NAND2_X1 U1143 ( .A1(n1422), .A2(n1423), .ZN(n1234) );
NAND2_X1 U1144 ( .A1(G131), .A2(n1175), .ZN(n1423) );
XOR2_X1 U1145 ( .A(n1424), .B(KEYINPUT51), .Z(n1422) );
OR2_X1 U1146 ( .A1(n1175), .A2(G131), .ZN(n1424) );
XOR2_X1 U1147 ( .A(G137), .B(n1350), .Z(n1175) );
XOR2_X1 U1148 ( .A(G134), .B(KEYINPUT9), .Z(n1350) );
INV_X1 U1149 ( .A(G472), .ZN(n1239) );
endmodule


