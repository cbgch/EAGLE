//Key = 1111000001011010111010000000110110110110010010111011000001000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376;

XOR2_X1 U756 ( .A(n1047), .B(G107), .Z(G9) );
NAND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
OR2_X1 U758 ( .A1(n1050), .A2(KEYINPUT26), .ZN(n1049) );
NAND3_X1 U759 ( .A1(n1051), .A2(n1052), .A3(KEYINPUT26), .ZN(n1048) );
NAND4_X1 U760 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NOR2_X1 U761 ( .A1(n1057), .A2(n1058), .ZN(G75) );
NOR4_X1 U762 ( .A1(G953), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1058) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR4_X1 U767 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
NOR3_X1 U768 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1071) );
NOR2_X1 U769 ( .A1(n1054), .A2(n1077), .ZN(n1070) );
NOR3_X1 U770 ( .A1(n1078), .A2(n1074), .A3(n1079), .ZN(n1068) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U772 ( .A1(n1082), .A2(n1073), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1072), .ZN(n1080) );
NOR2_X1 U774 ( .A1(n1084), .A2(n1055), .ZN(n1083) );
NOR2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR4_X1 U776 ( .A1(n1078), .A2(n1087), .A3(n1072), .A4(n1073), .ZN(n1064) );
INV_X1 U777 ( .A(n1088), .ZN(n1073) );
INV_X1 U778 ( .A(n1089), .ZN(n1072) );
INV_X1 U779 ( .A(n1054), .ZN(n1078) );
NOR3_X1 U780 ( .A1(n1059), .A2(G953), .A3(G952), .ZN(n1057) );
AND4_X1 U781 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1059) );
NOR3_X1 U782 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
XOR2_X1 U783 ( .A(n1097), .B(n1098), .Z(n1096) );
XNOR2_X1 U784 ( .A(KEYINPUT9), .B(n1099), .ZN(n1098) );
XOR2_X1 U785 ( .A(n1100), .B(n1101), .Z(n1095) );
NOR2_X1 U786 ( .A1(n1102), .A2(KEYINPUT24), .ZN(n1101) );
NAND3_X1 U787 ( .A1(n1077), .A2(n1103), .A3(n1086), .ZN(n1094) );
NOR3_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1092) );
NOR3_X1 U789 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
INV_X1 U790 ( .A(KEYINPUT3), .ZN(n1107) );
NOR2_X1 U791 ( .A1(KEYINPUT3), .A2(G475), .ZN(n1105) );
XOR2_X1 U792 ( .A(KEYINPUT51), .B(n1110), .Z(n1104) );
NOR2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
AND2_X1 U794 ( .A1(n1113), .A2(G478), .ZN(n1111) );
XOR2_X1 U795 ( .A(KEYINPUT35), .B(n1114), .Z(n1091) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(G72) );
NOR2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U798 ( .A(n1119), .B(KEYINPUT14), .Z(n1118) );
NAND3_X1 U799 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
NOR3_X1 U800 ( .A1(n1120), .A2(n1123), .A3(n1122), .ZN(n1117) );
XOR2_X1 U801 ( .A(n1124), .B(n1125), .Z(n1122) );
XOR2_X1 U802 ( .A(KEYINPUT1), .B(n1126), .Z(n1125) );
XOR2_X1 U803 ( .A(KEYINPUT53), .B(KEYINPUT44), .Z(n1126) );
XOR2_X1 U804 ( .A(n1127), .B(n1128), .Z(n1124) );
XOR2_X1 U805 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U806 ( .A1(G900), .A2(n1121), .ZN(n1123) );
NAND2_X1 U807 ( .A1(G953), .A2(n1131), .ZN(n1115) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1131) );
NAND2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(G69) );
NAND2_X1 U810 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND4_X1 U811 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1134) );
NOR2_X1 U812 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
OR2_X1 U813 ( .A1(n1121), .A2(G224), .ZN(n1138) );
NAND2_X1 U814 ( .A1(n1142), .A2(n1143), .ZN(n1132) );
NAND2_X1 U815 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND4_X1 U816 ( .A1(n1146), .A2(n1136), .A3(n1147), .A4(n1121), .ZN(n1145) );
INV_X1 U817 ( .A(n1140), .ZN(n1146) );
NAND2_X1 U818 ( .A1(G953), .A2(G224), .ZN(n1144) );
INV_X1 U819 ( .A(n1135), .ZN(n1142) );
NAND2_X1 U820 ( .A1(n1148), .A2(n1137), .ZN(n1135) );
INV_X1 U821 ( .A(n1149), .ZN(n1137) );
XOR2_X1 U822 ( .A(n1150), .B(n1151), .Z(n1148) );
NOR2_X1 U823 ( .A1(KEYINPUT30), .A2(n1152), .ZN(n1151) );
NOR3_X1 U824 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1150) );
NOR2_X1 U825 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR3_X1 U826 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1156) );
AND2_X1 U827 ( .A1(n1161), .A2(KEYINPUT27), .ZN(n1160) );
NOR2_X1 U828 ( .A1(KEYINPUT27), .A2(n1162), .ZN(n1159) );
NOR2_X1 U829 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U830 ( .A1(KEYINPUT52), .A2(n1165), .ZN(n1163) );
NOR2_X1 U831 ( .A1(KEYINPUT49), .A2(n1166), .ZN(n1158) );
NOR4_X1 U832 ( .A1(n1167), .A2(n1164), .A3(KEYINPUT52), .A4(KEYINPUT49), .ZN(n1154) );
NOR2_X1 U833 ( .A1(n1168), .A2(n1166), .ZN(n1153) );
INV_X1 U834 ( .A(KEYINPUT52), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1169), .A2(n1164), .ZN(n1168) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1167), .ZN(n1169) );
INV_X1 U837 ( .A(KEYINPUT49), .ZN(n1165) );
NOR3_X1 U838 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(G66) );
AND3_X1 U839 ( .A1(KEYINPUT5), .A2(G953), .A3(G952), .ZN(n1172) );
NOR2_X1 U840 ( .A1(KEYINPUT5), .A2(n1173), .ZN(n1171) );
INV_X1 U841 ( .A(n1174), .ZN(n1173) );
XOR2_X1 U842 ( .A(n1175), .B(n1176), .Z(n1170) );
NOR2_X1 U843 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U844 ( .A1(KEYINPUT16), .A2(n1179), .ZN(n1175) );
INV_X1 U845 ( .A(n1180), .ZN(n1179) );
NOR2_X1 U846 ( .A1(n1174), .A2(n1181), .ZN(G63) );
XOR2_X1 U847 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND2_X1 U848 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
XOR2_X1 U849 ( .A(KEYINPUT6), .B(G478), .Z(n1185) );
NOR3_X1 U850 ( .A1(n1174), .A2(n1186), .A3(n1187), .ZN(G60) );
NOR3_X1 U851 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
NOR2_X1 U852 ( .A1(KEYINPUT34), .A2(n1191), .ZN(n1190) );
NOR2_X1 U853 ( .A1(n1192), .A2(n1193), .ZN(n1186) );
NOR2_X1 U854 ( .A1(n1191), .A2(n1194), .ZN(n1192) );
INV_X1 U855 ( .A(KEYINPUT34), .ZN(n1194) );
XNOR2_X1 U856 ( .A(n1189), .B(KEYINPUT12), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1178), .A2(n1109), .ZN(n1189) );
XOR2_X1 U858 ( .A(n1195), .B(n1196), .Z(G6) );
XOR2_X1 U859 ( .A(KEYINPUT7), .B(G104), .Z(n1196) );
NOR2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
NOR2_X1 U861 ( .A1(n1174), .A2(n1199), .ZN(G57) );
XOR2_X1 U862 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U863 ( .A(n1202), .B(n1203), .Z(n1201) );
XOR2_X1 U864 ( .A(n1204), .B(KEYINPUT10), .Z(n1203) );
NAND2_X1 U865 ( .A1(n1184), .A2(G472), .ZN(n1202) );
XNOR2_X1 U866 ( .A(n1205), .B(n1206), .ZN(n1200) );
NOR2_X1 U867 ( .A1(n1207), .A2(n1208), .ZN(G54) );
XOR2_X1 U868 ( .A(KEYINPUT60), .B(n1174), .Z(n1208) );
XOR2_X1 U869 ( .A(n1209), .B(n1210), .Z(n1207) );
NAND2_X1 U870 ( .A1(n1184), .A2(G469), .ZN(n1210) );
NAND2_X1 U871 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
NAND2_X1 U872 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U873 ( .A(n1215), .B(KEYINPUT40), .Z(n1211) );
OR2_X1 U874 ( .A1(n1213), .A2(n1214), .ZN(n1215) );
XNOR2_X1 U875 ( .A(n1216), .B(n1217), .ZN(n1213) );
XOR2_X1 U876 ( .A(n1218), .B(n1219), .Z(n1217) );
XNOR2_X1 U877 ( .A(n1129), .B(KEYINPUT0), .ZN(n1216) );
NOR2_X1 U878 ( .A1(n1174), .A2(n1220), .ZN(G51) );
XOR2_X1 U879 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U880 ( .A(n1223), .B(n1224), .Z(n1222) );
NOR2_X1 U881 ( .A1(KEYINPUT4), .A2(n1225), .ZN(n1223) );
XNOR2_X1 U882 ( .A(G125), .B(n1226), .ZN(n1221) );
NAND2_X1 U883 ( .A1(n1184), .A2(n1102), .ZN(n1226) );
INV_X1 U884 ( .A(n1178), .ZN(n1184) );
NAND2_X1 U885 ( .A1(G902), .A2(n1061), .ZN(n1178) );
NAND4_X1 U886 ( .A1(n1227), .A2(n1147), .A3(n1228), .A4(n1229), .ZN(n1061) );
XNOR2_X1 U887 ( .A(KEYINPUT33), .B(n1140), .ZN(n1229) );
NAND3_X1 U888 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1140) );
OR2_X1 U889 ( .A1(n1233), .A2(n1082), .ZN(n1232) );
INV_X1 U890 ( .A(n1120), .ZN(n1228) );
NAND4_X1 U891 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1120) );
NOR3_X1 U892 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1237) );
NOR3_X1 U893 ( .A1(n1241), .A2(n1242), .A3(n1087), .ZN(n1240) );
NOR2_X1 U894 ( .A1(n1243), .A2(n1244), .ZN(n1238) );
NOR2_X1 U895 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
AND2_X1 U896 ( .A1(n1075), .A2(n1247), .ZN(n1246) );
NOR2_X1 U897 ( .A1(n1082), .A2(n1248), .ZN(n1245) );
NOR2_X1 U898 ( .A1(n1247), .A2(n1053), .ZN(n1082) );
INV_X1 U899 ( .A(n1249), .ZN(n1234) );
INV_X1 U900 ( .A(n1141), .ZN(n1147) );
NAND3_X1 U901 ( .A1(n1250), .A2(n1050), .A3(n1251), .ZN(n1141) );
NAND3_X1 U902 ( .A1(n1247), .A2(n1252), .A3(n1253), .ZN(n1251) );
XNOR2_X1 U903 ( .A(n1054), .B(KEYINPUT17), .ZN(n1253) );
OR2_X1 U904 ( .A1(n1197), .A2(n1242), .ZN(n1050) );
NAND2_X1 U905 ( .A1(n1252), .A2(n1054), .ZN(n1197) );
XOR2_X1 U906 ( .A(n1136), .B(KEYINPUT45), .Z(n1227) );
NOR2_X1 U907 ( .A1(n1121), .A2(G952), .ZN(n1174) );
XNOR2_X1 U908 ( .A(n1254), .B(n1249), .ZN(G48) );
NOR3_X1 U909 ( .A1(n1198), .A2(n1087), .A3(n1241), .ZN(n1249) );
XOR2_X1 U910 ( .A(n1239), .B(n1255), .Z(G45) );
NOR2_X1 U911 ( .A1(KEYINPUT55), .A2(n1256), .ZN(n1255) );
AND4_X1 U912 ( .A1(n1051), .A2(n1055), .A3(n1076), .A4(n1257), .ZN(n1239) );
NOR3_X1 U913 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1257) );
XNOR2_X1 U914 ( .A(G140), .B(n1261), .ZN(G42) );
NAND4_X1 U915 ( .A1(KEYINPUT63), .A2(n1262), .A3(n1247), .A4(n1075), .ZN(n1261) );
XNOR2_X1 U916 ( .A(G137), .B(n1235), .ZN(G39) );
NAND4_X1 U917 ( .A1(n1262), .A2(n1089), .A3(n1263), .A4(n1264), .ZN(n1235) );
NAND2_X1 U918 ( .A1(n1265), .A2(n1266), .ZN(G36) );
NAND2_X1 U919 ( .A1(G134), .A2(n1267), .ZN(n1266) );
XOR2_X1 U920 ( .A(KEYINPUT57), .B(n1268), .Z(n1265) );
NOR2_X1 U921 ( .A1(G134), .A2(n1267), .ZN(n1268) );
NAND3_X1 U922 ( .A1(n1053), .A2(n1269), .A3(n1262), .ZN(n1267) );
XNOR2_X1 U923 ( .A(KEYINPUT36), .B(n1248), .ZN(n1269) );
XOR2_X1 U924 ( .A(G131), .B(n1270), .Z(G33) );
NOR3_X1 U925 ( .A1(n1248), .A2(n1271), .A3(n1244), .ZN(n1270) );
INV_X1 U926 ( .A(n1262), .ZN(n1244) );
NOR4_X1 U927 ( .A1(n1067), .A2(n1272), .A3(n1258), .A4(n1074), .ZN(n1262) );
INV_X1 U928 ( .A(n1077), .ZN(n1074) );
XNOR2_X1 U929 ( .A(n1247), .B(KEYINPUT39), .ZN(n1271) );
XOR2_X1 U930 ( .A(G128), .B(n1273), .Z(G30) );
NOR3_X1 U931 ( .A1(n1241), .A2(n1274), .A3(n1242), .ZN(n1273) );
XNOR2_X1 U932 ( .A(n1051), .B(KEYINPUT43), .ZN(n1274) );
NAND4_X1 U933 ( .A1(n1055), .A2(n1263), .A3(n1275), .A4(n1264), .ZN(n1241) );
XNOR2_X1 U934 ( .A(G101), .B(n1136), .ZN(G3) );
NAND3_X1 U935 ( .A1(n1089), .A2(n1252), .A3(n1076), .ZN(n1136) );
XNOR2_X1 U936 ( .A(G125), .B(n1236), .ZN(G27) );
NAND4_X1 U937 ( .A1(n1088), .A2(n1247), .A3(n1276), .A4(n1075), .ZN(n1236) );
NOR2_X1 U938 ( .A1(n1258), .A2(n1087), .ZN(n1276) );
INV_X1 U939 ( .A(n1275), .ZN(n1258) );
NAND2_X1 U940 ( .A1(n1063), .A2(n1277), .ZN(n1275) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1278), .A4(n1279), .ZN(n1277) );
INV_X1 U942 ( .A(G900), .ZN(n1279) );
NAND2_X1 U943 ( .A1(n1280), .A2(n1281), .ZN(G24) );
NAND2_X1 U944 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
XOR2_X1 U945 ( .A(KEYINPUT37), .B(n1284), .Z(n1280) );
NOR2_X1 U946 ( .A1(n1282), .A2(n1283), .ZN(n1284) );
INV_X1 U947 ( .A(n1230), .ZN(n1282) );
NAND4_X1 U948 ( .A1(n1285), .A2(n1054), .A3(n1286), .A4(n1287), .ZN(n1230) );
NOR2_X1 U949 ( .A1(n1264), .A2(n1263), .ZN(n1054) );
XNOR2_X1 U950 ( .A(G119), .B(n1231), .ZN(G21) );
NAND4_X1 U951 ( .A1(n1285), .A2(n1089), .A3(n1263), .A4(n1264), .ZN(n1231) );
XNOR2_X1 U952 ( .A(G116), .B(n1288), .ZN(G18) );
NOR2_X1 U953 ( .A1(n1289), .A2(KEYINPUT19), .ZN(n1288) );
NOR2_X1 U954 ( .A1(n1242), .A2(n1233), .ZN(n1289) );
INV_X1 U955 ( .A(n1053), .ZN(n1242) );
NOR2_X1 U956 ( .A1(n1286), .A2(n1259), .ZN(n1053) );
INV_X1 U957 ( .A(n1287), .ZN(n1259) );
XNOR2_X1 U958 ( .A(G113), .B(n1290), .ZN(G15) );
NOR2_X1 U959 ( .A1(n1291), .A2(KEYINPUT59), .ZN(n1290) );
NOR2_X1 U960 ( .A1(n1198), .A2(n1233), .ZN(n1291) );
NAND2_X1 U961 ( .A1(n1285), .A2(n1076), .ZN(n1233) );
INV_X1 U962 ( .A(n1248), .ZN(n1076) );
NAND2_X1 U963 ( .A1(n1090), .A2(n1263), .ZN(n1248) );
AND3_X1 U964 ( .A1(n1051), .A2(n1056), .A3(n1088), .ZN(n1285) );
NOR2_X1 U965 ( .A1(n1085), .A2(n1292), .ZN(n1088) );
INV_X1 U966 ( .A(n1086), .ZN(n1292) );
INV_X1 U967 ( .A(n1247), .ZN(n1198) );
NOR2_X1 U968 ( .A1(n1287), .A2(n1260), .ZN(n1247) );
INV_X1 U969 ( .A(n1286), .ZN(n1260) );
XNOR2_X1 U970 ( .A(G110), .B(n1250), .ZN(G12) );
NAND3_X1 U971 ( .A1(n1075), .A2(n1252), .A3(n1089), .ZN(n1250) );
NOR2_X1 U972 ( .A1(n1287), .A2(n1286), .ZN(n1089) );
NAND2_X1 U973 ( .A1(n1103), .A2(n1293), .ZN(n1286) );
OR2_X1 U974 ( .A1(n1109), .A2(n1108), .ZN(n1293) );
NAND2_X1 U975 ( .A1(n1108), .A2(n1109), .ZN(n1103) );
INV_X1 U976 ( .A(G475), .ZN(n1109) );
NOR2_X1 U977 ( .A1(n1193), .A2(G902), .ZN(n1108) );
INV_X1 U978 ( .A(n1188), .ZN(n1193) );
XNOR2_X1 U979 ( .A(n1294), .B(n1295), .ZN(n1188) );
XNOR2_X1 U980 ( .A(n1296), .B(n1297), .ZN(n1295) );
NOR2_X1 U981 ( .A1(G104), .A2(KEYINPUT61), .ZN(n1297) );
NAND2_X1 U982 ( .A1(KEYINPUT41), .A2(n1254), .ZN(n1296) );
XOR2_X1 U983 ( .A(n1298), .B(n1299), .Z(n1294) );
XOR2_X1 U984 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U985 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U986 ( .A(n1304), .B(n1305), .ZN(n1302) );
INV_X1 U987 ( .A(G113), .ZN(n1305) );
NAND2_X1 U988 ( .A1(n1306), .A2(G214), .ZN(n1304) );
XNOR2_X1 U989 ( .A(G131), .B(n1307), .ZN(n1300) );
XNOR2_X1 U990 ( .A(KEYINPUT15), .B(n1256), .ZN(n1307) );
NAND2_X1 U991 ( .A1(KEYINPUT2), .A2(G122), .ZN(n1298) );
NAND3_X1 U992 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1287) );
INV_X1 U993 ( .A(n1112), .ZN(n1310) );
NOR2_X1 U994 ( .A1(n1113), .A2(G478), .ZN(n1112) );
OR2_X1 U995 ( .A1(G478), .A2(KEYINPUT11), .ZN(n1309) );
NAND3_X1 U996 ( .A1(G478), .A2(n1113), .A3(KEYINPUT11), .ZN(n1308) );
NAND2_X1 U997 ( .A1(n1183), .A2(n1311), .ZN(n1113) );
XOR2_X1 U998 ( .A(n1312), .B(n1313), .Z(n1183) );
XOR2_X1 U999 ( .A(n1314), .B(n1315), .Z(n1313) );
NAND2_X1 U1000 ( .A1(KEYINPUT50), .A2(n1316), .ZN(n1315) );
NAND2_X1 U1001 ( .A1(n1317), .A2(n1318), .ZN(n1314) );
NAND2_X1 U1002 ( .A1(G134), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1003 ( .A(KEYINPUT38), .B(n1320), .Z(n1317) );
NOR2_X1 U1004 ( .A1(G134), .A2(n1319), .ZN(n1320) );
NAND2_X1 U1005 ( .A1(n1321), .A2(n1322), .ZN(n1319) );
NAND2_X1 U1006 ( .A1(G128), .A2(n1256), .ZN(n1322) );
XOR2_X1 U1007 ( .A(KEYINPUT29), .B(n1323), .Z(n1321) );
NOR2_X1 U1008 ( .A1(G128), .A2(n1256), .ZN(n1323) );
INV_X1 U1009 ( .A(G143), .ZN(n1256) );
XOR2_X1 U1010 ( .A(n1324), .B(n1325), .Z(n1312) );
NOR4_X1 U1011 ( .A1(KEYINPUT25), .A2(G953), .A3(n1326), .A4(n1177), .ZN(n1325) );
XNOR2_X1 U1012 ( .A(G107), .B(G122), .ZN(n1324) );
AND3_X1 U1013 ( .A1(n1055), .A2(n1056), .A3(n1051), .ZN(n1252) );
INV_X1 U1014 ( .A(n1087), .ZN(n1051) );
NAND2_X1 U1015 ( .A1(n1067), .A2(n1077), .ZN(n1087) );
NAND2_X1 U1016 ( .A1(G214), .A2(n1327), .ZN(n1077) );
NAND2_X1 U1017 ( .A1(n1328), .A2(n1329), .ZN(n1067) );
OR2_X1 U1018 ( .A1(n1100), .A2(n1102), .ZN(n1329) );
XOR2_X1 U1019 ( .A(n1330), .B(KEYINPUT22), .Z(n1328) );
NAND2_X1 U1020 ( .A1(n1102), .A2(n1100), .ZN(n1330) );
NAND2_X1 U1021 ( .A1(n1331), .A2(n1311), .ZN(n1100) );
XOR2_X1 U1022 ( .A(n1224), .B(n1332), .Z(n1331) );
XOR2_X1 U1023 ( .A(G125), .B(n1225), .Z(n1332) );
XNOR2_X1 U1024 ( .A(n1333), .B(n1334), .ZN(n1225) );
XNOR2_X1 U1025 ( .A(n1335), .B(n1336), .ZN(n1224) );
XNOR2_X1 U1026 ( .A(n1161), .B(n1152), .ZN(n1336) );
XNOR2_X1 U1027 ( .A(G110), .B(n1283), .ZN(n1152) );
INV_X1 U1028 ( .A(G122), .ZN(n1283) );
XOR2_X1 U1029 ( .A(n1337), .B(n1338), .Z(n1335) );
NOR2_X1 U1030 ( .A1(KEYINPUT42), .A2(n1157), .ZN(n1338) );
INV_X1 U1031 ( .A(n1167), .ZN(n1157) );
XOR2_X1 U1032 ( .A(G113), .B(n1339), .Z(n1167) );
NOR2_X1 U1033 ( .A1(KEYINPUT62), .A2(n1340), .ZN(n1339) );
NAND2_X1 U1034 ( .A1(G224), .A2(n1121), .ZN(n1337) );
AND2_X1 U1035 ( .A1(G210), .A2(n1327), .ZN(n1102) );
NAND2_X1 U1036 ( .A1(n1341), .A2(n1311), .ZN(n1327) );
INV_X1 U1037 ( .A(G237), .ZN(n1341) );
NAND2_X1 U1038 ( .A1(n1063), .A2(n1342), .ZN(n1056) );
NAND3_X1 U1039 ( .A1(G902), .A2(n1278), .A3(n1149), .ZN(n1342) );
NOR2_X1 U1040 ( .A1(G898), .A2(n1121), .ZN(n1149) );
NAND3_X1 U1041 ( .A1(n1278), .A2(n1121), .A3(G952), .ZN(n1063) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1278) );
INV_X1 U1043 ( .A(n1272), .ZN(n1055) );
NAND2_X1 U1044 ( .A1(n1085), .A2(n1086), .ZN(n1272) );
NAND2_X1 U1045 ( .A1(G221), .A2(n1343), .ZN(n1086) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1311), .ZN(n1343) );
XNOR2_X1 U1047 ( .A(n1344), .B(n1097), .ZN(n1085) );
NAND2_X1 U1048 ( .A1(n1345), .A2(n1311), .ZN(n1097) );
XOR2_X1 U1049 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1050 ( .A(n1348), .B(n1214), .Z(n1347) );
XNOR2_X1 U1051 ( .A(n1349), .B(n1350), .ZN(n1214) );
XOR2_X1 U1052 ( .A(G140), .B(G110), .Z(n1350) );
NAND2_X1 U1053 ( .A1(G227), .A2(n1121), .ZN(n1349) );
INV_X1 U1054 ( .A(G953), .ZN(n1121) );
XNOR2_X1 U1055 ( .A(n1351), .B(n1352), .ZN(n1346) );
INV_X1 U1056 ( .A(G137), .ZN(n1352) );
NAND2_X1 U1057 ( .A1(KEYINPUT31), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1058 ( .A(n1354), .B(n1218), .Z(n1353) );
XNOR2_X1 U1059 ( .A(n1161), .B(KEYINPUT20), .ZN(n1218) );
INV_X1 U1060 ( .A(n1164), .ZN(n1161) );
XOR2_X1 U1061 ( .A(n1355), .B(n1206), .Z(n1164) );
INV_X1 U1062 ( .A(n1356), .ZN(n1206) );
XNOR2_X1 U1063 ( .A(G104), .B(G107), .ZN(n1355) );
NOR2_X1 U1064 ( .A1(KEYINPUT13), .A2(n1357), .ZN(n1354) );
XOR2_X1 U1065 ( .A(n1129), .B(n1334), .Z(n1357) );
NOR2_X1 U1066 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1129) );
NAND2_X1 U1067 ( .A1(KEYINPUT47), .A2(n1099), .ZN(n1344) );
INV_X1 U1068 ( .A(G469), .ZN(n1099) );
NOR2_X1 U1069 ( .A1(n1263), .A2(n1090), .ZN(n1075) );
INV_X1 U1070 ( .A(n1264), .ZN(n1090) );
NAND3_X1 U1071 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1264) );
NAND2_X1 U1072 ( .A1(n1361), .A2(n1180), .ZN(n1360) );
OR3_X1 U1073 ( .A1(n1180), .A2(n1361), .A3(G902), .ZN(n1359) );
NOR2_X1 U1074 ( .A1(n1177), .A2(G234), .ZN(n1361) );
INV_X1 U1075 ( .A(G217), .ZN(n1177) );
XNOR2_X1 U1076 ( .A(n1362), .B(n1363), .ZN(n1180) );
XOR2_X1 U1077 ( .A(n1364), .B(n1365), .Z(n1363) );
NOR2_X1 U1078 ( .A1(G110), .A2(KEYINPUT58), .ZN(n1365) );
NOR3_X1 U1079 ( .A1(n1366), .A2(G953), .A3(n1326), .ZN(n1364) );
XNOR2_X1 U1080 ( .A(G234), .B(KEYINPUT8), .ZN(n1326) );
INV_X1 U1081 ( .A(G221), .ZN(n1366) );
XOR2_X1 U1082 ( .A(n1127), .B(n1367), .Z(n1362) );
XOR2_X1 U1083 ( .A(n1368), .B(n1303), .Z(n1127) );
XOR2_X1 U1084 ( .A(G140), .B(G125), .Z(n1303) );
NAND2_X1 U1085 ( .A1(G902), .A2(G217), .ZN(n1358) );
XOR2_X1 U1086 ( .A(n1114), .B(KEYINPUT21), .Z(n1263) );
XNOR2_X1 U1087 ( .A(n1369), .B(G472), .ZN(n1114) );
NAND2_X1 U1088 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XNOR2_X1 U1089 ( .A(KEYINPUT32), .B(n1311), .ZN(n1371) );
INV_X1 U1090 ( .A(G902), .ZN(n1311) );
XNOR2_X1 U1091 ( .A(n1356), .B(n1372), .ZN(n1370) );
XNOR2_X1 U1092 ( .A(n1373), .B(n1374), .ZN(n1372) );
NOR2_X1 U1093 ( .A1(KEYINPUT23), .A2(n1204), .ZN(n1374) );
NAND2_X1 U1094 ( .A1(n1306), .A2(G210), .ZN(n1204) );
NOR2_X1 U1095 ( .A1(G953), .A2(G237), .ZN(n1306) );
NAND2_X1 U1096 ( .A1(KEYINPUT46), .A2(n1205), .ZN(n1373) );
XOR2_X1 U1097 ( .A(n1375), .B(n1376), .Z(n1205) );
XNOR2_X1 U1098 ( .A(G113), .B(n1333), .ZN(n1376) );
NAND2_X1 U1099 ( .A1(KEYINPUT18), .A2(G143), .ZN(n1333) );
XNOR2_X1 U1100 ( .A(n1219), .B(n1340), .ZN(n1375) );
XNOR2_X1 U1101 ( .A(n1316), .B(n1367), .ZN(n1340) );
XOR2_X1 U1102 ( .A(G119), .B(KEYINPUT54), .Z(n1367) );
INV_X1 U1103 ( .A(G116), .ZN(n1316) );
XNOR2_X1 U1104 ( .A(n1368), .B(n1348), .ZN(n1219) );
XOR2_X1 U1105 ( .A(n1130), .B(KEYINPUT28), .Z(n1348) );
XOR2_X1 U1106 ( .A(G131), .B(G134), .Z(n1130) );
XNOR2_X1 U1107 ( .A(G137), .B(n1334), .ZN(n1368) );
XNOR2_X1 U1108 ( .A(n1254), .B(G128), .ZN(n1334) );
INV_X1 U1109 ( .A(G146), .ZN(n1254) );
XOR2_X1 U1110 ( .A(G101), .B(KEYINPUT48), .Z(n1356) );
endmodule


