//Key = 1001100111011100111011011010010110001010101011000011011000110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346;

NAND3_X1 U737 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(G9) );
OR2_X1 U738 ( .A1(G107), .A2(KEYINPUT40), .ZN(n1025) );
NAND3_X1 U739 ( .A1(KEYINPUT40), .A2(G107), .A3(n1026), .ZN(n1024) );
NAND2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(n1023) );
NAND2_X1 U741 ( .A1(n1029), .A2(KEYINPUT40), .ZN(n1028) );
XNOR2_X1 U742 ( .A(G107), .B(KEYINPUT8), .ZN(n1029) );
NOR2_X1 U743 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR3_X1 U744 ( .A1(n1032), .A2(G953), .A3(G952), .ZN(n1031) );
NOR4_X1 U745 ( .A1(n1033), .A2(n1034), .A3(G953), .A4(n1032), .ZN(n1030) );
AND4_X1 U746 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1032) );
NOR3_X1 U747 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
XOR2_X1 U748 ( .A(n1042), .B(KEYINPUT32), .Z(n1041) );
NAND3_X1 U749 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1039) );
NOR3_X1 U750 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1037) );
AND3_X1 U751 ( .A1(KEYINPUT42), .A2(n1049), .A3(G475), .ZN(n1048) );
NOR2_X1 U752 ( .A1(KEYINPUT42), .A2(n1049), .ZN(n1047) );
XOR2_X1 U753 ( .A(n1050), .B(n1051), .Z(n1046) );
XOR2_X1 U754 ( .A(n1052), .B(KEYINPUT27), .Z(n1051) );
NAND2_X1 U755 ( .A1(KEYINPUT7), .A2(n1053), .ZN(n1050) );
INV_X1 U756 ( .A(n1054), .ZN(n1053) );
NOR4_X1 U757 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1034) );
NOR3_X1 U758 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1056) );
AND3_X1 U759 ( .A1(n1062), .A2(n1063), .A3(KEYINPUT56), .ZN(n1061) );
INV_X1 U760 ( .A(n1064), .ZN(n1063) );
NOR2_X1 U761 ( .A1(n1065), .A2(n1062), .ZN(n1060) );
NOR3_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
AND2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U764 ( .A1(n1071), .A2(n1072), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U766 ( .A1(KEYINPUT56), .A2(n1064), .ZN(n1066) );
AND2_X1 U767 ( .A1(n1075), .A2(KEYINPUT61), .ZN(n1059) );
NAND3_X1 U768 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1033) );
NAND2_X1 U769 ( .A1(n1075), .A2(n1079), .ZN(n1077) );
NAND2_X1 U770 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND3_X1 U771 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1055), .A2(n1057), .ZN(n1083) );
NAND3_X1 U773 ( .A1(n1085), .A2(n1086), .A3(n1045), .ZN(n1082) );
NAND4_X1 U774 ( .A1(n1040), .A2(n1042), .A3(n1043), .A4(n1087), .ZN(n1085) );
INV_X1 U775 ( .A(KEYINPUT61), .ZN(n1087) );
INV_X1 U776 ( .A(n1088), .ZN(n1040) );
NAND2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1080) );
NOR3_X1 U778 ( .A1(n1091), .A2(n1072), .A3(n1062), .ZN(n1075) );
INV_X1 U779 ( .A(n1036), .ZN(n1072) );
XOR2_X1 U780 ( .A(n1092), .B(n1093), .Z(G72) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U782 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U783 ( .A1(G953), .A2(n1098), .ZN(n1097) );
XOR2_X1 U784 ( .A(n1099), .B(n1100), .Z(n1096) );
XOR2_X1 U785 ( .A(n1101), .B(n1102), .Z(n1100) );
NAND2_X1 U786 ( .A1(KEYINPUT29), .A2(n1103), .ZN(n1102) );
NAND3_X1 U787 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1101) );
NAND2_X1 U788 ( .A1(KEYINPUT30), .A2(n1107), .ZN(n1105) );
NAND2_X1 U789 ( .A1(n1108), .A2(n1109), .ZN(n1104) );
INV_X1 U790 ( .A(KEYINPUT30), .ZN(n1109) );
XOR2_X1 U791 ( .A(n1110), .B(G131), .Z(n1099) );
NAND2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1094) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1112) );
XNOR2_X1 U794 ( .A(KEYINPUT22), .B(n1113), .ZN(n1111) );
NOR2_X1 U795 ( .A1(n1076), .A2(G953), .ZN(n1092) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(G69) );
XOR2_X1 U797 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U799 ( .A1(G953), .A2(n1120), .ZN(n1119) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(n1118) );
NAND2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NAND2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
INV_X1 U803 ( .A(KEYINPUT35), .ZN(n1126) );
XOR2_X1 U804 ( .A(G113), .B(n1127), .Z(n1125) );
NAND3_X1 U805 ( .A1(n1128), .A2(n1129), .A3(KEYINPUT35), .ZN(n1123) );
XOR2_X1 U806 ( .A(G113), .B(n1130), .Z(n1128) );
NAND2_X1 U807 ( .A1(G953), .A2(n1131), .ZN(n1116) );
NAND2_X1 U808 ( .A1(n1132), .A2(G898), .ZN(n1131) );
XNOR2_X1 U809 ( .A(G224), .B(KEYINPUT4), .ZN(n1132) );
NOR2_X1 U810 ( .A1(n1078), .A2(G953), .ZN(n1114) );
NOR2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XNOR2_X1 U812 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR2_X1 U813 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR4_X1 U814 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(G63) );
AND2_X1 U815 ( .A1(KEYINPUT45), .A2(n1133), .ZN(n1142) );
NOR3_X1 U816 ( .A1(KEYINPUT45), .A2(G953), .A3(G952), .ZN(n1141) );
NOR4_X1 U817 ( .A1(n1143), .A2(n1138), .A3(KEYINPUT48), .A4(n1144), .ZN(n1140) );
NOR2_X1 U818 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
NOR3_X1 U819 ( .A1(n1138), .A2(n1147), .A3(n1144), .ZN(n1146) );
NOR2_X1 U820 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
INV_X1 U821 ( .A(KEYINPUT48), .ZN(n1149) );
INV_X1 U822 ( .A(n1143), .ZN(n1145) );
NAND2_X1 U823 ( .A1(KEYINPUT23), .A2(n1148), .ZN(n1143) );
NOR2_X1 U824 ( .A1(n1133), .A2(n1150), .ZN(G60) );
XOR2_X1 U825 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U826 ( .A1(KEYINPUT25), .A2(n1153), .ZN(n1152) );
OR2_X1 U827 ( .A1(n1138), .A2(n1154), .ZN(n1151) );
XNOR2_X1 U828 ( .A(G104), .B(n1155), .ZN(G6) );
NOR2_X1 U829 ( .A1(n1156), .A2(n1157), .ZN(G57) );
XOR2_X1 U830 ( .A(n1158), .B(KEYINPUT63), .Z(n1157) );
NAND2_X1 U831 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NAND2_X1 U832 ( .A1(n1133), .A2(n1161), .ZN(n1160) );
OR3_X1 U833 ( .A1(G952), .A2(G953), .A3(n1161), .ZN(n1159) );
INV_X1 U834 ( .A(KEYINPUT52), .ZN(n1161) );
XNOR2_X1 U835 ( .A(n1162), .B(n1163), .ZN(n1156) );
NOR2_X1 U836 ( .A1(n1164), .A2(n1138), .ZN(n1163) );
NOR2_X1 U837 ( .A1(n1133), .A2(n1165), .ZN(G54) );
XOR2_X1 U838 ( .A(n1166), .B(n1167), .Z(n1165) );
XNOR2_X1 U839 ( .A(n1168), .B(KEYINPUT3), .ZN(n1167) );
NAND2_X1 U840 ( .A1(n1169), .A2(KEYINPUT13), .ZN(n1168) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U842 ( .A(KEYINPUT26), .B(n1172), .ZN(n1171) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1138), .ZN(n1166) );
NOR2_X1 U844 ( .A1(n1133), .A2(n1174), .ZN(G51) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U846 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR2_X1 U847 ( .A1(G125), .A2(KEYINPUT6), .ZN(n1178) );
NOR2_X1 U848 ( .A1(n1054), .A2(n1138), .ZN(n1177) );
NAND2_X1 U849 ( .A1(G902), .A2(n1179), .ZN(n1138) );
NAND2_X1 U850 ( .A1(n1078), .A2(n1076), .ZN(n1179) );
AND2_X1 U851 ( .A1(n1180), .A2(n1181), .ZN(n1076) );
AND4_X1 U852 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
AND4_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1180) );
AND4_X1 U854 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1078) );
NOR4_X1 U855 ( .A1(n1027), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1193) );
INV_X1 U856 ( .A(n1026), .ZN(n1027) );
NAND3_X1 U857 ( .A1(n1073), .A2(n1036), .A3(n1197), .ZN(n1026) );
NOR2_X1 U858 ( .A1(n1198), .A2(n1199), .ZN(n1192) );
INV_X1 U859 ( .A(n1155), .ZN(n1199) );
NAND3_X1 U860 ( .A1(n1197), .A2(n1036), .A3(n1074), .ZN(n1155) );
NOR3_X1 U861 ( .A1(n1064), .A2(n1200), .A3(n1201), .ZN(n1198) );
NOR2_X1 U862 ( .A1(KEYINPUT36), .A2(n1202), .ZN(n1201) );
NOR2_X1 U863 ( .A1(n1090), .A2(n1203), .ZN(n1202) );
AND2_X1 U864 ( .A1(n1204), .A2(KEYINPUT36), .ZN(n1200) );
NOR2_X1 U865 ( .A1(n1113), .A2(G952), .ZN(n1133) );
NAND2_X1 U866 ( .A1(n1205), .A2(n1206), .ZN(G48) );
NAND2_X1 U867 ( .A1(n1207), .A2(n1189), .ZN(n1206) );
NAND2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U869 ( .A1(KEYINPUT43), .A2(KEYINPUT18), .ZN(n1209) );
NAND3_X1 U870 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1205) );
INV_X1 U871 ( .A(KEYINPUT43), .ZN(n1212) );
OR2_X1 U872 ( .A1(G146), .A2(KEYINPUT18), .ZN(n1211) );
NAND2_X1 U873 ( .A1(KEYINPUT18), .A2(n1213), .ZN(n1210) );
OR2_X1 U874 ( .A1(n1189), .A2(G146), .ZN(n1213) );
NAND4_X1 U875 ( .A1(n1214), .A2(n1074), .A3(n1215), .A4(n1216), .ZN(n1189) );
XNOR2_X1 U876 ( .A(G143), .B(n1188), .ZN(G45) );
NAND4_X1 U877 ( .A1(n1090), .A2(n1215), .A3(n1069), .A4(n1217), .ZN(n1188) );
NOR3_X1 U878 ( .A1(n1035), .A2(n1218), .A3(n1219), .ZN(n1217) );
XNOR2_X1 U879 ( .A(n1220), .B(n1172), .ZN(G42) );
NAND2_X1 U880 ( .A1(KEYINPUT20), .A2(n1187), .ZN(n1220) );
NAND4_X1 U881 ( .A1(n1221), .A2(n1074), .A3(n1222), .A4(n1223), .ZN(n1187) );
XNOR2_X1 U882 ( .A(G137), .B(n1224), .ZN(G39) );
NAND2_X1 U883 ( .A1(KEYINPUT21), .A2(n1225), .ZN(n1224) );
INV_X1 U884 ( .A(n1186), .ZN(n1225) );
NAND2_X1 U885 ( .A1(n1221), .A2(n1226), .ZN(n1186) );
XOR2_X1 U886 ( .A(G134), .B(n1227), .Z(G36) );
NOR2_X1 U887 ( .A1(KEYINPUT2), .A2(n1185), .ZN(n1227) );
NAND3_X1 U888 ( .A1(n1069), .A2(n1073), .A3(n1221), .ZN(n1185) );
XOR2_X1 U889 ( .A(G131), .B(n1228), .Z(G33) );
NOR2_X1 U890 ( .A1(KEYINPUT57), .A2(n1184), .ZN(n1228) );
NAND3_X1 U891 ( .A1(n1074), .A2(n1069), .A3(n1221), .ZN(n1184) );
NOR4_X1 U892 ( .A1(n1058), .A2(n1086), .A3(n1055), .A4(n1219), .ZN(n1221) );
XNOR2_X1 U893 ( .A(G128), .B(n1183), .ZN(G30) );
NAND4_X1 U894 ( .A1(n1214), .A2(n1073), .A3(n1229), .A4(n1216), .ZN(n1183) );
XNOR2_X1 U895 ( .A(G101), .B(n1190), .ZN(G3) );
NAND3_X1 U896 ( .A1(n1069), .A2(n1197), .A3(n1070), .ZN(n1190) );
XNOR2_X1 U897 ( .A(G125), .B(n1182), .ZN(G27) );
NAND4_X1 U898 ( .A1(n1214), .A2(n1074), .A3(n1222), .A4(n1089), .ZN(n1182) );
NOR3_X1 U899 ( .A1(n1230), .A2(n1219), .A3(n1231), .ZN(n1214) );
AND2_X1 U900 ( .A1(n1232), .A2(n1062), .ZN(n1219) );
XOR2_X1 U901 ( .A(n1233), .B(KEYINPUT62), .Z(n1232) );
NAND4_X1 U902 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1098), .ZN(n1233) );
INV_X1 U903 ( .A(G900), .ZN(n1098) );
XNOR2_X1 U904 ( .A(G122), .B(n1191), .ZN(G24) );
NAND4_X1 U905 ( .A1(n1235), .A2(n1036), .A3(n1236), .A4(n1237), .ZN(n1191) );
NOR2_X1 U906 ( .A1(n1223), .A2(n1216), .ZN(n1036) );
XNOR2_X1 U907 ( .A(n1196), .B(n1238), .ZN(G21) );
NAND2_X1 U908 ( .A1(KEYINPUT54), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U909 ( .A(KEYINPUT5), .B(n1240), .ZN(n1239) );
AND2_X1 U910 ( .A1(n1226), .A2(n1235), .ZN(n1196) );
NOR3_X1 U911 ( .A1(n1222), .A2(n1230), .A3(n1091), .ZN(n1226) );
INV_X1 U912 ( .A(n1070), .ZN(n1091) );
INV_X1 U913 ( .A(n1223), .ZN(n1230) );
XOR2_X1 U914 ( .A(G116), .B(n1195), .Z(G18) );
AND3_X1 U915 ( .A1(n1069), .A2(n1073), .A3(n1235), .ZN(n1195) );
NOR2_X1 U916 ( .A1(n1237), .A2(n1035), .ZN(n1073) );
INV_X1 U917 ( .A(n1236), .ZN(n1035) );
XOR2_X1 U918 ( .A(G113), .B(n1194), .Z(G15) );
AND3_X1 U919 ( .A1(n1074), .A2(n1069), .A3(n1235), .ZN(n1194) );
AND3_X1 U920 ( .A1(n1090), .A2(n1241), .A3(n1089), .ZN(n1235) );
INV_X1 U921 ( .A(n1057), .ZN(n1089) );
NAND3_X1 U922 ( .A1(n1088), .A2(n1043), .A3(n1042), .ZN(n1057) );
NOR2_X1 U923 ( .A1(n1223), .A2(n1222), .ZN(n1069) );
NOR2_X1 U924 ( .A1(n1236), .A2(n1218), .ZN(n1074) );
INV_X1 U925 ( .A(n1237), .ZN(n1218) );
XOR2_X1 U926 ( .A(G110), .B(n1242), .Z(G12) );
NOR3_X1 U927 ( .A1(n1064), .A2(KEYINPUT15), .A3(n1204), .ZN(n1242) );
INV_X1 U928 ( .A(n1197), .ZN(n1204) );
NOR2_X1 U929 ( .A1(n1231), .A2(n1203), .ZN(n1197) );
NAND2_X1 U930 ( .A1(n1229), .A2(n1241), .ZN(n1203) );
NAND2_X1 U931 ( .A1(n1062), .A2(n1243), .ZN(n1241) );
NAND4_X1 U932 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1120), .ZN(n1243) );
INV_X1 U933 ( .A(G898), .ZN(n1120) );
NAND3_X1 U934 ( .A1(n1234), .A2(n1113), .A3(G952), .ZN(n1062) );
NAND2_X1 U935 ( .A1(G234), .A2(G237), .ZN(n1234) );
XNOR2_X1 U936 ( .A(n1215), .B(KEYINPUT59), .ZN(n1229) );
INV_X1 U937 ( .A(n1086), .ZN(n1215) );
NAND2_X1 U938 ( .A1(n1088), .A2(n1244), .ZN(n1086) );
NAND2_X1 U939 ( .A1(n1042), .A2(n1043), .ZN(n1244) );
NAND3_X1 U940 ( .A1(n1173), .A2(n1245), .A3(n1246), .ZN(n1043) );
INV_X1 U941 ( .A(G469), .ZN(n1173) );
NAND2_X1 U942 ( .A1(G469), .A2(n1247), .ZN(n1042) );
NAND2_X1 U943 ( .A1(n1246), .A2(n1245), .ZN(n1247) );
XOR2_X1 U944 ( .A(n1170), .B(n1248), .Z(n1246) );
XNOR2_X1 U945 ( .A(n1249), .B(KEYINPUT33), .ZN(n1248) );
NAND2_X1 U946 ( .A1(KEYINPUT58), .A2(n1250), .ZN(n1249) );
XNOR2_X1 U947 ( .A(KEYINPUT17), .B(n1172), .ZN(n1250) );
XOR2_X1 U948 ( .A(n1251), .B(n1252), .Z(n1170) );
XOR2_X1 U949 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U950 ( .A(n1255), .B(n1256), .ZN(n1254) );
AND2_X1 U951 ( .A1(n1113), .A2(G227), .ZN(n1256) );
XOR2_X1 U952 ( .A(n1257), .B(n1258), .Z(n1251) );
XOR2_X1 U953 ( .A(KEYINPUT49), .B(G110), .Z(n1258) );
XNOR2_X1 U954 ( .A(n1110), .B(n1259), .ZN(n1257) );
NAND2_X1 U955 ( .A1(n1260), .A2(n1261), .ZN(n1110) );
NAND2_X1 U956 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XOR2_X1 U957 ( .A(KEYINPUT51), .B(n1264), .Z(n1260) );
NOR2_X1 U958 ( .A1(n1262), .A2(n1263), .ZN(n1264) );
XNOR2_X1 U959 ( .A(G143), .B(G146), .ZN(n1262) );
NAND2_X1 U960 ( .A1(G221), .A2(n1265), .ZN(n1088) );
INV_X1 U961 ( .A(n1090), .ZN(n1231) );
NOR2_X1 U962 ( .A1(n1084), .A2(n1055), .ZN(n1090) );
INV_X1 U963 ( .A(n1045), .ZN(n1055) );
NAND2_X1 U964 ( .A1(G214), .A2(n1266), .ZN(n1045) );
INV_X1 U965 ( .A(n1058), .ZN(n1084) );
XOR2_X1 U966 ( .A(n1267), .B(n1054), .Z(n1058) );
NAND2_X1 U967 ( .A1(G210), .A2(n1266), .ZN(n1054) );
NAND2_X1 U968 ( .A1(n1268), .A2(n1245), .ZN(n1266) );
XNOR2_X1 U969 ( .A(G237), .B(KEYINPUT37), .ZN(n1268) );
XOR2_X1 U970 ( .A(n1052), .B(KEYINPUT34), .Z(n1267) );
NAND2_X1 U971 ( .A1(n1269), .A2(n1245), .ZN(n1052) );
XNOR2_X1 U972 ( .A(n1175), .B(n1270), .ZN(n1269) );
XNOR2_X1 U973 ( .A(KEYINPUT24), .B(n1107), .ZN(n1270) );
XNOR2_X1 U974 ( .A(n1271), .B(n1272), .ZN(n1175) );
XOR2_X1 U975 ( .A(n1273), .B(n1274), .Z(n1272) );
NOR2_X1 U976 ( .A1(KEYINPUT60), .A2(n1122), .ZN(n1274) );
XNOR2_X1 U977 ( .A(G110), .B(G122), .ZN(n1122) );
AND2_X1 U978 ( .A1(n1113), .A2(G224), .ZN(n1273) );
XOR2_X1 U979 ( .A(n1275), .B(n1127), .Z(n1271) );
XOR2_X1 U980 ( .A(n1130), .B(n1129), .Z(n1127) );
XNOR2_X1 U981 ( .A(n1253), .B(n1276), .ZN(n1129) );
NOR2_X1 U982 ( .A1(KEYINPUT10), .A2(n1259), .ZN(n1276) );
INV_X1 U983 ( .A(G107), .ZN(n1259) );
XNOR2_X1 U984 ( .A(G101), .B(G104), .ZN(n1253) );
XNOR2_X1 U985 ( .A(G119), .B(n1277), .ZN(n1130) );
NAND3_X1 U986 ( .A1(n1222), .A2(n1223), .A3(n1070), .ZN(n1064) );
NOR2_X1 U987 ( .A1(n1236), .A2(n1237), .ZN(n1070) );
NAND2_X1 U988 ( .A1(n1278), .A2(n1044), .ZN(n1237) );
NAND2_X1 U989 ( .A1(n1279), .A2(n1154), .ZN(n1044) );
INV_X1 U990 ( .A(G475), .ZN(n1154) );
NAND2_X1 U991 ( .A1(G475), .A2(n1049), .ZN(n1278) );
INV_X1 U992 ( .A(n1279), .ZN(n1049) );
NOR2_X1 U993 ( .A1(n1153), .A2(G902), .ZN(n1279) );
XNOR2_X1 U994 ( .A(n1280), .B(n1281), .ZN(n1153) );
XOR2_X1 U995 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U996 ( .A(n1284), .B(n1285), .ZN(n1283) );
NAND2_X1 U997 ( .A1(KEYINPUT12), .A2(n1286), .ZN(n1285) );
INV_X1 U998 ( .A(G104), .ZN(n1286) );
NAND4_X1 U999 ( .A1(KEYINPUT0), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n1284) );
NAND3_X1 U1000 ( .A1(KEYINPUT38), .A2(n1290), .A3(n1208), .ZN(n1289) );
INV_X1 U1001 ( .A(n1291), .ZN(n1290) );
NAND2_X1 U1002 ( .A1(G146), .A2(n1291), .ZN(n1288) );
NAND2_X1 U1003 ( .A1(KEYINPUT11), .A2(n1292), .ZN(n1291) );
OR2_X1 U1004 ( .A1(n1292), .A2(KEYINPUT38), .ZN(n1287) );
NAND3_X1 U1005 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1292) );
XNOR2_X1 U1006 ( .A(n1108), .B(KEYINPUT55), .ZN(n1295) );
OR3_X1 U1007 ( .A1(G125), .A2(G140), .A3(KEYINPUT44), .ZN(n1294) );
NAND2_X1 U1008 ( .A1(n1296), .A2(KEYINPUT44), .ZN(n1293) );
XNOR2_X1 U1009 ( .A(G113), .B(n1297), .ZN(n1282) );
NOR2_X1 U1010 ( .A1(n1298), .A2(KEYINPUT19), .ZN(n1297) );
NOR2_X1 U1011 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
INV_X1 U1012 ( .A(G214), .ZN(n1299) );
XOR2_X1 U1013 ( .A(n1301), .B(n1302), .Z(n1280) );
XNOR2_X1 U1014 ( .A(KEYINPUT41), .B(n1303), .ZN(n1302) );
XNOR2_X1 U1015 ( .A(G122), .B(G131), .ZN(n1301) );
XOR2_X1 U1016 ( .A(n1304), .B(n1144), .Z(n1236) );
INV_X1 U1017 ( .A(G478), .ZN(n1144) );
NAND2_X1 U1018 ( .A1(n1245), .A2(n1148), .ZN(n1304) );
NAND2_X1 U1019 ( .A1(n1305), .A2(n1306), .ZN(n1148) );
NAND4_X1 U1020 ( .A1(G217), .A2(G234), .A3(n1307), .A4(n1113), .ZN(n1306) );
NAND2_X1 U1021 ( .A1(n1308), .A2(n1309), .ZN(n1305) );
NAND3_X1 U1022 ( .A1(G234), .A2(n1113), .A3(G217), .ZN(n1309) );
XNOR2_X1 U1023 ( .A(n1307), .B(KEYINPUT14), .ZN(n1308) );
XNOR2_X1 U1024 ( .A(n1310), .B(n1311), .ZN(n1307) );
XNOR2_X1 U1025 ( .A(G107), .B(n1312), .ZN(n1311) );
NAND2_X1 U1026 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND2_X1 U1027 ( .A1(n1315), .A2(n1303), .ZN(n1314) );
XOR2_X1 U1028 ( .A(KEYINPUT16), .B(n1316), .Z(n1313) );
NOR2_X1 U1029 ( .A1(n1315), .A2(n1303), .ZN(n1316) );
XNOR2_X1 U1030 ( .A(G116), .B(n1317), .ZN(n1310) );
XOR2_X1 U1031 ( .A(G134), .B(G122), .Z(n1317) );
XOR2_X1 U1032 ( .A(n1318), .B(n1137), .Z(n1223) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1265), .ZN(n1137) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1245), .ZN(n1265) );
NAND2_X1 U1035 ( .A1(n1135), .A2(n1245), .ZN(n1318) );
XNOR2_X1 U1036 ( .A(n1319), .B(n1320), .ZN(n1135) );
XOR2_X1 U1037 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1038 ( .A(n1323), .B(n1324), .Z(n1322) );
NAND2_X1 U1039 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1040 ( .A1(G119), .A2(n1263), .ZN(n1326) );
XOR2_X1 U1041 ( .A(n1327), .B(KEYINPUT1), .Z(n1325) );
NAND2_X1 U1042 ( .A1(n1315), .A2(n1240), .ZN(n1327) );
INV_X1 U1043 ( .A(G119), .ZN(n1240) );
NAND2_X1 U1044 ( .A1(n1328), .A2(n1106), .ZN(n1323) );
INV_X1 U1045 ( .A(n1296), .ZN(n1106) );
NOR2_X1 U1046 ( .A1(n1172), .A2(G125), .ZN(n1296) );
XOR2_X1 U1047 ( .A(KEYINPUT46), .B(n1329), .Z(n1328) );
NOR2_X1 U1048 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
AND2_X1 U1049 ( .A1(KEYINPUT9), .A2(n1108), .ZN(n1331) );
NOR2_X1 U1050 ( .A1(n1107), .A2(G140), .ZN(n1108) );
INV_X1 U1051 ( .A(G125), .ZN(n1107) );
NOR2_X1 U1052 ( .A1(KEYINPUT9), .A2(n1172), .ZN(n1330) );
INV_X1 U1053 ( .A(G140), .ZN(n1172) );
AND3_X1 U1054 ( .A1(G221), .A2(n1113), .A3(G234), .ZN(n1321) );
INV_X1 U1055 ( .A(G953), .ZN(n1113) );
XOR2_X1 U1056 ( .A(n1332), .B(n1333), .Z(n1319) );
XNOR2_X1 U1057 ( .A(KEYINPUT28), .B(n1208), .ZN(n1333) );
XNOR2_X1 U1058 ( .A(G137), .B(G110), .ZN(n1332) );
INV_X1 U1059 ( .A(n1216), .ZN(n1222) );
XOR2_X1 U1060 ( .A(n1334), .B(n1164), .Z(n1216) );
INV_X1 U1061 ( .A(G472), .ZN(n1164) );
NAND2_X1 U1062 ( .A1(n1162), .A2(n1245), .ZN(n1334) );
INV_X1 U1063 ( .A(G902), .ZN(n1245) );
XNOR2_X1 U1064 ( .A(n1335), .B(n1336), .ZN(n1162) );
XOR2_X1 U1065 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1066 ( .A(G101), .B(n1339), .Z(n1338) );
NOR2_X1 U1067 ( .A1(KEYINPUT47), .A2(n1340), .ZN(n1339) );
XNOR2_X1 U1068 ( .A(G119), .B(n1341), .ZN(n1340) );
NAND2_X1 U1069 ( .A1(KEYINPUT31), .A2(n1277), .ZN(n1341) );
XNOR2_X1 U1070 ( .A(G116), .B(KEYINPUT39), .ZN(n1277) );
NOR2_X1 U1071 ( .A1(n1342), .A2(n1300), .ZN(n1337) );
OR2_X1 U1072 ( .A1(G953), .A2(G237), .ZN(n1300) );
INV_X1 U1073 ( .A(G210), .ZN(n1342) );
XNOR2_X1 U1074 ( .A(n1275), .B(n1343), .ZN(n1335) );
INV_X1 U1075 ( .A(n1255), .ZN(n1343) );
XNOR2_X1 U1076 ( .A(G131), .B(n1103), .ZN(n1255) );
XNOR2_X1 U1077 ( .A(G134), .B(G137), .ZN(n1103) );
XOR2_X1 U1078 ( .A(n1344), .B(n1345), .Z(n1275) );
XNOR2_X1 U1079 ( .A(n1303), .B(G113), .ZN(n1345) );
INV_X1 U1080 ( .A(G143), .ZN(n1303) );
XNOR2_X1 U1081 ( .A(n1346), .B(n1315), .ZN(n1344) );
INV_X1 U1082 ( .A(n1263), .ZN(n1315) );
XOR2_X1 U1083 ( .A(G128), .B(KEYINPUT53), .Z(n1263) );
NAND2_X1 U1084 ( .A1(KEYINPUT50), .A2(n1208), .ZN(n1346) );
INV_X1 U1085 ( .A(G146), .ZN(n1208) );
endmodule


