//Key = 0100000100101100000000001011101101111110000000101110101010000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;

XNOR2_X1 U794 ( .A(G107), .B(n1103), .ZN(G9) );
NAND2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U796 ( .A(n1106), .B(KEYINPUT50), .Z(n1104) );
NOR2_X1 U797 ( .A1(n1107), .A2(n1108), .ZN(G75) );
NOR4_X1 U798 ( .A1(G953), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NOR2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR3_X1 U801 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
NOR3_X1 U802 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1117) );
NOR3_X1 U803 ( .A1(n1122), .A2(KEYINPUT56), .A3(n1123), .ZN(n1121) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1120) );
NOR3_X1 U805 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1124) );
AND2_X1 U806 ( .A1(n1129), .A2(KEYINPUT22), .ZN(n1128) );
NOR3_X1 U807 ( .A1(KEYINPUT22), .A2(n1130), .A3(n1131), .ZN(n1127) );
AND2_X1 U808 ( .A1(n1132), .A2(KEYINPUT56), .ZN(n1126) );
NOR2_X1 U809 ( .A1(n1133), .A2(n1134), .ZN(n1119) );
NOR2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR3_X1 U811 ( .A1(n1125), .A2(n1137), .A3(n1134), .ZN(n1114) );
NOR2_X1 U812 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U813 ( .A1(n1140), .A2(n1118), .ZN(n1139) );
NOR2_X1 U814 ( .A1(n1141), .A2(n1105), .ZN(n1140) );
NOR2_X1 U815 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1144), .A2(n1116), .ZN(n1138) );
INV_X1 U817 ( .A(n1145), .ZN(n1116) );
NOR2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
NOR3_X1 U819 ( .A1(n1109), .A2(G953), .A3(G952), .ZN(n1107) );
AND3_X1 U820 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1109) );
NOR4_X1 U821 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
INV_X1 U822 ( .A(n1155), .ZN(n1152) );
NAND3_X1 U823 ( .A1(n1156), .A2(n1157), .A3(n1131), .ZN(n1151) );
NOR3_X1 U824 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1149) );
XOR2_X1 U825 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U826 ( .A1(KEYINPUT11), .A2(n1163), .ZN(n1162) );
XNOR2_X1 U827 ( .A(G478), .B(KEYINPUT33), .ZN(n1163) );
NOR2_X1 U828 ( .A1(n1164), .A2(n1165), .ZN(n1159) );
NOR3_X1 U829 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1148) );
NOR3_X1 U830 ( .A1(n1169), .A2(KEYINPUT60), .A3(n1170), .ZN(n1168) );
AND2_X1 U831 ( .A1(n1169), .A2(KEYINPUT60), .ZN(n1167) );
XOR2_X1 U832 ( .A(n1171), .B(n1172), .Z(n1166) );
NOR3_X1 U833 ( .A1(n1173), .A2(KEYINPUT47), .A3(G902), .ZN(n1172) );
XOR2_X1 U834 ( .A(n1174), .B(n1175), .Z(G72) );
NOR2_X1 U835 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
AND2_X1 U836 ( .A1(G227), .A2(G900), .ZN(n1176) );
NAND2_X1 U837 ( .A1(n1178), .A2(n1179), .ZN(n1174) );
NAND2_X1 U838 ( .A1(n1180), .A2(n1177), .ZN(n1179) );
XOR2_X1 U839 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND3_X1 U840 ( .A1(n1182), .A2(G900), .A3(G953), .ZN(n1178) );
AND2_X1 U841 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND2_X1 U842 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U843 ( .A(n1187), .B(n1188), .Z(n1185) );
NAND2_X1 U844 ( .A1(n1189), .A2(n1190), .ZN(n1183) );
XOR2_X1 U845 ( .A(G125), .B(n1188), .Z(n1190) );
NOR2_X1 U846 ( .A1(KEYINPUT9), .A2(n1191), .ZN(n1188) );
XNOR2_X1 U847 ( .A(KEYINPUT29), .B(n1186), .ZN(n1189) );
XOR2_X1 U848 ( .A(n1192), .B(n1193), .Z(n1186) );
NOR2_X1 U849 ( .A1(KEYINPUT8), .A2(n1194), .ZN(n1193) );
XOR2_X1 U850 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U851 ( .A1(KEYINPUT43), .A2(n1197), .ZN(n1195) );
NAND2_X1 U852 ( .A1(n1198), .A2(n1199), .ZN(G69) );
NAND3_X1 U853 ( .A1(G953), .A2(n1200), .A3(n1201), .ZN(n1199) );
XOR2_X1 U854 ( .A(KEYINPUT30), .B(n1202), .Z(n1198) );
NOR2_X1 U855 ( .A1(n1203), .A2(n1201), .ZN(n1202) );
XOR2_X1 U856 ( .A(n1204), .B(n1205), .Z(n1201) );
NOR2_X1 U857 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U858 ( .A1(G898), .A2(n1177), .ZN(n1206) );
NAND2_X1 U859 ( .A1(n1177), .A2(n1208), .ZN(n1204) );
AND2_X1 U860 ( .A1(n1200), .A2(G953), .ZN(n1203) );
NAND2_X1 U861 ( .A1(G898), .A2(G224), .ZN(n1200) );
NOR2_X1 U862 ( .A1(n1209), .A2(n1210), .ZN(G66) );
XOR2_X1 U863 ( .A(n1211), .B(n1212), .Z(n1210) );
NAND2_X1 U864 ( .A1(n1213), .A2(n1164), .ZN(n1211) );
NOR2_X1 U865 ( .A1(n1209), .A2(n1214), .ZN(G63) );
NOR3_X1 U866 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
AND3_X1 U867 ( .A1(n1218), .A2(G478), .A3(n1213), .ZN(n1217) );
NOR2_X1 U868 ( .A1(n1219), .A2(n1218), .ZN(n1216) );
AND2_X1 U869 ( .A1(n1111), .A2(G478), .ZN(n1219) );
NOR2_X1 U870 ( .A1(n1209), .A2(n1220), .ZN(G60) );
XOR2_X1 U871 ( .A(n1221), .B(n1222), .Z(n1220) );
NAND2_X1 U872 ( .A1(n1213), .A2(G475), .ZN(n1221) );
XOR2_X1 U873 ( .A(n1223), .B(n1224), .Z(G6) );
NAND2_X1 U874 ( .A1(KEYINPUT37), .A2(G104), .ZN(n1224) );
NAND4_X1 U875 ( .A1(n1136), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
XOR2_X1 U876 ( .A(KEYINPUT20), .B(n1105), .Z(n1227) );
NOR2_X1 U877 ( .A1(n1209), .A2(n1228), .ZN(G57) );
XOR2_X1 U878 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U879 ( .A(n1231), .B(n1232), .Z(n1230) );
NAND2_X1 U880 ( .A1(n1233), .A2(KEYINPUT46), .ZN(n1232) );
XOR2_X1 U881 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND2_X1 U882 ( .A1(n1213), .A2(G472), .ZN(n1234) );
NOR2_X1 U883 ( .A1(KEYINPUT58), .A2(n1236), .ZN(n1229) );
NOR2_X1 U884 ( .A1(n1209), .A2(n1237), .ZN(G54) );
XOR2_X1 U885 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U886 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR2_X1 U887 ( .A1(n1242), .A2(n1243), .ZN(n1238) );
XOR2_X1 U888 ( .A(KEYINPUT0), .B(n1244), .Z(n1243) );
NOR2_X1 U889 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
INV_X1 U890 ( .A(n1247), .ZN(n1245) );
NOR2_X1 U891 ( .A1(n1248), .A2(n1247), .ZN(n1242) );
NAND3_X1 U892 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1247) );
OR2_X1 U893 ( .A1(n1252), .A2(KEYINPUT27), .ZN(n1251) );
NAND3_X1 U894 ( .A1(KEYINPUT27), .A2(n1252), .A3(n1253), .ZN(n1250) );
INV_X1 U895 ( .A(n1254), .ZN(n1253) );
NAND2_X1 U896 ( .A1(n1255), .A2(n1254), .ZN(n1249) );
NAND2_X1 U897 ( .A1(n1256), .A2(KEYINPUT27), .ZN(n1255) );
XNOR2_X1 U898 ( .A(n1252), .B(KEYINPUT31), .ZN(n1256) );
XNOR2_X1 U899 ( .A(n1257), .B(KEYINPUT32), .ZN(n1252) );
XNOR2_X1 U900 ( .A(n1246), .B(KEYINPUT4), .ZN(n1248) );
XNOR2_X1 U901 ( .A(n1258), .B(n1259), .ZN(n1246) );
NAND2_X1 U902 ( .A1(n1260), .A2(KEYINPUT38), .ZN(n1258) );
XOR2_X1 U903 ( .A(n1192), .B(n1261), .Z(n1260) );
NOR3_X1 U904 ( .A1(n1262), .A2(n1209), .A3(n1263), .ZN(G51) );
NOR3_X1 U905 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
XOR2_X1 U906 ( .A(n1267), .B(n1268), .Z(n1264) );
NAND2_X1 U907 ( .A1(KEYINPUT28), .A2(n1269), .ZN(n1268) );
INV_X1 U908 ( .A(n1270), .ZN(n1269) );
NOR2_X1 U909 ( .A1(n1177), .A2(G952), .ZN(n1209) );
NOR2_X1 U910 ( .A1(n1271), .A2(n1272), .ZN(n1262) );
XOR2_X1 U911 ( .A(n1267), .B(n1273), .Z(n1272) );
NAND2_X1 U912 ( .A1(KEYINPUT28), .A2(n1270), .ZN(n1273) );
NAND2_X1 U913 ( .A1(n1274), .A2(n1275), .ZN(n1270) );
NAND2_X1 U914 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
OR2_X1 U915 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
XOR2_X1 U916 ( .A(KEYINPUT12), .B(n1280), .Z(n1274) );
NOR3_X1 U917 ( .A1(n1277), .A2(n1278), .A3(n1279), .ZN(n1280) );
NAND2_X1 U918 ( .A1(n1213), .A2(n1171), .ZN(n1267) );
INV_X1 U919 ( .A(n1241), .ZN(n1213) );
NAND2_X1 U920 ( .A1(G902), .A2(n1111), .ZN(n1241) );
NAND3_X1 U921 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1111) );
INV_X1 U922 ( .A(n1208), .ZN(n1283) );
NAND4_X1 U923 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1208) );
NOR3_X1 U924 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1287) );
INV_X1 U925 ( .A(n1291), .ZN(n1290) );
AND3_X1 U926 ( .A1(n1136), .A2(n1292), .A3(n1147), .ZN(n1288) );
OR2_X1 U927 ( .A1(n1293), .A2(KEYINPUT25), .ZN(n1286) );
NAND2_X1 U928 ( .A1(n1105), .A2(n1294), .ZN(n1285) );
NAND4_X1 U929 ( .A1(n1295), .A2(n1296), .A3(n1297), .A4(n1298), .ZN(n1294) );
NAND2_X1 U930 ( .A1(n1226), .A2(n1299), .ZN(n1298) );
NAND2_X1 U931 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND3_X1 U932 ( .A1(n1146), .A2(n1125), .A3(KEYINPUT40), .ZN(n1301) );
INV_X1 U933 ( .A(n1122), .ZN(n1125) );
NAND2_X1 U934 ( .A1(n1136), .A2(n1225), .ZN(n1300) );
OR2_X1 U935 ( .A1(n1106), .A2(KEYINPUT23), .ZN(n1297) );
OR2_X1 U936 ( .A1(n1302), .A2(KEYINPUT40), .ZN(n1296) );
XOR2_X1 U937 ( .A(n1303), .B(KEYINPUT53), .Z(n1295) );
NAND2_X1 U938 ( .A1(n1304), .A2(n1305), .ZN(n1284) );
NAND2_X1 U939 ( .A1(n1306), .A2(n1307), .ZN(n1304) );
NAND4_X1 U940 ( .A1(n1122), .A2(n1129), .A3(KEYINPUT25), .A4(n1308), .ZN(n1307) );
NOR3_X1 U941 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1308) );
NAND2_X1 U942 ( .A1(KEYINPUT23), .A2(n1312), .ZN(n1306) );
INV_X1 U943 ( .A(n1106), .ZN(n1312) );
NAND3_X1 U944 ( .A1(n1225), .A2(n1226), .A3(n1135), .ZN(n1106) );
INV_X1 U945 ( .A(n1118), .ZN(n1225) );
NAND2_X1 U946 ( .A1(n1181), .A2(n1313), .ZN(n1282) );
INV_X1 U947 ( .A(KEYINPUT42), .ZN(n1313) );
NAND4_X1 U948 ( .A1(n1314), .A2(n1315), .A3(n1316), .A4(n1317), .ZN(n1181) );
NOR4_X1 U949 ( .A1(n1318), .A2(n1319), .A3(n1320), .A4(n1321), .ZN(n1317) );
NOR2_X1 U950 ( .A1(n1322), .A2(n1323), .ZN(n1316) );
NAND2_X1 U951 ( .A1(n1324), .A2(n1105), .ZN(n1314) );
NAND2_X1 U952 ( .A1(KEYINPUT42), .A2(n1325), .ZN(n1281) );
NOR2_X1 U953 ( .A1(n1266), .A2(n1265), .ZN(n1271) );
INV_X1 U954 ( .A(KEYINPUT10), .ZN(n1265) );
INV_X1 U955 ( .A(n1207), .ZN(n1266) );
XOR2_X1 U956 ( .A(G146), .B(n1319), .Z(G48) );
AND3_X1 U957 ( .A1(n1136), .A2(n1105), .A3(n1326), .ZN(n1319) );
XOR2_X1 U958 ( .A(G143), .B(n1327), .Z(G45) );
NOR2_X1 U959 ( .A1(n1305), .A2(n1328), .ZN(n1327) );
XOR2_X1 U960 ( .A(KEYINPUT1), .B(n1324), .Z(n1328) );
AND3_X1 U961 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1324) );
XOR2_X1 U962 ( .A(n1191), .B(n1315), .Z(G42) );
NAND3_X1 U963 ( .A1(n1145), .A2(n1132), .A3(n1332), .ZN(n1315) );
XOR2_X1 U964 ( .A(G137), .B(n1318), .Z(G39) );
AND3_X1 U965 ( .A1(n1326), .A2(n1122), .A3(n1145), .ZN(n1318) );
XOR2_X1 U966 ( .A(G134), .B(n1323), .Z(G36) );
AND3_X1 U967 ( .A1(n1145), .A2(n1135), .A3(n1331), .ZN(n1323) );
XOR2_X1 U968 ( .A(G131), .B(n1322), .Z(G33) );
AND3_X1 U969 ( .A1(n1145), .A2(n1136), .A3(n1331), .ZN(n1322) );
AND3_X1 U970 ( .A1(n1132), .A2(n1333), .A3(n1147), .ZN(n1331) );
NOR2_X1 U971 ( .A1(n1143), .A2(n1153), .ZN(n1145) );
INV_X1 U972 ( .A(n1142), .ZN(n1153) );
NAND2_X1 U973 ( .A1(n1334), .A2(n1335), .ZN(G30) );
NAND2_X1 U974 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U975 ( .A(KEYINPUT39), .B(n1320), .Z(n1336) );
INV_X1 U976 ( .A(n1325), .ZN(n1320) );
NAND2_X1 U977 ( .A1(G128), .A2(n1338), .ZN(n1334) );
XOR2_X1 U978 ( .A(n1325), .B(KEYINPUT16), .Z(n1338) );
NAND3_X1 U979 ( .A1(n1105), .A2(n1135), .A3(n1326), .ZN(n1325) );
AND4_X1 U980 ( .A1(n1132), .A2(n1158), .A3(n1333), .A4(n1339), .ZN(n1326) );
INV_X1 U981 ( .A(n1123), .ZN(n1132) );
XOR2_X1 U982 ( .A(n1231), .B(n1291), .Z(G3) );
NAND4_X1 U983 ( .A1(n1122), .A2(n1147), .A3(n1105), .A4(n1226), .ZN(n1291) );
XOR2_X1 U984 ( .A(G125), .B(n1321), .Z(G27) );
AND3_X1 U985 ( .A1(n1129), .A2(n1105), .A3(n1332), .ZN(n1321) );
AND3_X1 U986 ( .A1(n1136), .A2(n1333), .A3(n1146), .ZN(n1332) );
NAND2_X1 U987 ( .A1(n1113), .A2(n1340), .ZN(n1333) );
NAND4_X1 U988 ( .A1(G953), .A2(G902), .A3(n1341), .A4(n1342), .ZN(n1340) );
INV_X1 U989 ( .A(G900), .ZN(n1342) );
INV_X1 U990 ( .A(n1134), .ZN(n1129) );
NAND2_X1 U991 ( .A1(n1343), .A2(n1344), .ZN(G24) );
OR2_X1 U992 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XOR2_X1 U993 ( .A(n1347), .B(KEYINPUT3), .Z(n1343) );
NAND2_X1 U994 ( .A1(n1346), .A2(n1348), .ZN(n1347) );
XOR2_X1 U995 ( .A(KEYINPUT7), .B(G122), .Z(n1348) );
NOR2_X1 U996 ( .A1(n1303), .A2(n1305), .ZN(n1346) );
NAND4_X1 U997 ( .A1(n1329), .A2(n1330), .A3(n1349), .A4(n1350), .ZN(n1303) );
NOR2_X1 U998 ( .A1(n1118), .A2(n1134), .ZN(n1350) );
NAND2_X1 U999 ( .A1(n1310), .A2(n1309), .ZN(n1118) );
XOR2_X1 U1000 ( .A(n1293), .B(n1351), .Z(G21) );
XNOR2_X1 U1001 ( .A(G119), .B(KEYINPUT21), .ZN(n1351) );
NAND4_X1 U1002 ( .A1(n1122), .A2(n1292), .A3(n1158), .A4(n1339), .ZN(n1293) );
XOR2_X1 U1003 ( .A(n1289), .B(n1352), .Z(G18) );
NOR2_X1 U1004 ( .A1(KEYINPUT6), .A2(n1353), .ZN(n1352) );
INV_X1 U1005 ( .A(G116), .ZN(n1353) );
AND3_X1 U1006 ( .A1(n1292), .A2(n1135), .A3(n1147), .ZN(n1289) );
AND2_X1 U1007 ( .A1(n1354), .A2(n1330), .ZN(n1135) );
XOR2_X1 U1008 ( .A(n1355), .B(n1356), .Z(G15) );
NAND3_X1 U1009 ( .A1(n1136), .A2(n1292), .A3(n1357), .ZN(n1356) );
XNOR2_X1 U1010 ( .A(n1147), .B(KEYINPUT54), .ZN(n1357) );
NOR2_X1 U1011 ( .A1(n1339), .A2(n1309), .ZN(n1147) );
NOR3_X1 U1012 ( .A1(n1305), .A2(n1311), .A3(n1134), .ZN(n1292) );
NAND2_X1 U1013 ( .A1(n1358), .A2(n1131), .ZN(n1134) );
INV_X1 U1014 ( .A(n1130), .ZN(n1358) );
NOR2_X1 U1015 ( .A1(n1330), .A2(n1354), .ZN(n1136) );
NAND2_X1 U1016 ( .A1(n1359), .A2(n1360), .ZN(G12) );
NAND3_X1 U1017 ( .A1(n1361), .A2(n1362), .A3(n1105), .ZN(n1360) );
XOR2_X1 U1018 ( .A(n1363), .B(KEYINPUT19), .Z(n1359) );
NAND2_X1 U1019 ( .A1(G110), .A2(n1364), .ZN(n1363) );
NAND2_X1 U1020 ( .A1(n1105), .A2(n1361), .ZN(n1364) );
XNOR2_X1 U1021 ( .A(n1302), .B(KEYINPUT17), .ZN(n1361) );
NAND3_X1 U1022 ( .A1(n1122), .A2(n1226), .A3(n1146), .ZN(n1302) );
NOR2_X1 U1023 ( .A1(n1158), .A2(n1310), .ZN(n1146) );
INV_X1 U1024 ( .A(n1339), .ZN(n1310) );
NAND2_X1 U1025 ( .A1(n1365), .A2(n1156), .ZN(n1339) );
NAND2_X1 U1026 ( .A1(n1164), .A2(n1165), .ZN(n1156) );
NAND2_X1 U1027 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
INV_X1 U1028 ( .A(n1165), .ZN(n1367) );
NAND2_X1 U1029 ( .A1(n1212), .A2(n1368), .ZN(n1165) );
XNOR2_X1 U1030 ( .A(n1369), .B(n1370), .ZN(n1212) );
XOR2_X1 U1031 ( .A(G119), .B(n1371), .Z(n1370) );
XOR2_X1 U1032 ( .A(G137), .B(G128), .Z(n1371) );
XOR2_X1 U1033 ( .A(n1372), .B(n1373), .Z(n1369) );
INV_X1 U1034 ( .A(n1374), .ZN(n1373) );
XOR2_X1 U1035 ( .A(n1257), .B(n1375), .Z(n1372) );
AND3_X1 U1036 ( .A1(G221), .A2(n1177), .A3(G234), .ZN(n1375) );
XNOR2_X1 U1037 ( .A(n1164), .B(KEYINPUT5), .ZN(n1366) );
AND2_X1 U1038 ( .A1(G217), .A2(n1376), .ZN(n1164) );
INV_X1 U1039 ( .A(n1309), .ZN(n1158) );
XOR2_X1 U1040 ( .A(n1377), .B(G472), .Z(n1309) );
NAND2_X1 U1041 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
XNOR2_X1 U1042 ( .A(n1380), .B(n1235), .ZN(n1379) );
XNOR2_X1 U1043 ( .A(n1381), .B(n1382), .ZN(n1235) );
XOR2_X1 U1044 ( .A(n1383), .B(n1384), .Z(n1382) );
XOR2_X1 U1045 ( .A(n1259), .B(n1355), .Z(n1381) );
INV_X1 U1046 ( .A(G113), .ZN(n1355) );
NAND2_X1 U1047 ( .A1(n1385), .A2(n1386), .ZN(n1380) );
NAND2_X1 U1048 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
XOR2_X1 U1049 ( .A(KEYINPUT45), .B(G101), .Z(n1388) );
INV_X1 U1050 ( .A(n1236), .ZN(n1387) );
XOR2_X1 U1051 ( .A(n1389), .B(KEYINPUT57), .Z(n1385) );
NAND2_X1 U1052 ( .A1(n1231), .A2(n1236), .ZN(n1389) );
NAND3_X1 U1053 ( .A1(n1390), .A2(n1177), .A3(G210), .ZN(n1236) );
INV_X1 U1054 ( .A(G101), .ZN(n1231) );
XOR2_X1 U1055 ( .A(KEYINPUT36), .B(G902), .Z(n1378) );
NOR2_X1 U1056 ( .A1(n1123), .A2(n1311), .ZN(n1226) );
INV_X1 U1057 ( .A(n1349), .ZN(n1311) );
NAND2_X1 U1058 ( .A1(n1113), .A2(n1391), .ZN(n1349) );
NAND4_X1 U1059 ( .A1(G953), .A2(G902), .A3(n1341), .A4(n1392), .ZN(n1391) );
INV_X1 U1060 ( .A(G898), .ZN(n1392) );
NAND3_X1 U1061 ( .A1(n1341), .A2(n1177), .A3(G952), .ZN(n1113) );
NAND2_X1 U1062 ( .A1(G237), .A2(G234), .ZN(n1341) );
NAND2_X1 U1063 ( .A1(n1130), .A2(n1131), .ZN(n1123) );
NAND2_X1 U1064 ( .A1(G221), .A2(n1376), .ZN(n1131) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1393), .ZN(n1376) );
NAND2_X1 U1066 ( .A1(n1394), .A2(n1155), .ZN(n1130) );
NAND2_X1 U1067 ( .A1(G469), .A2(n1395), .ZN(n1155) );
NAND2_X1 U1068 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
XNOR2_X1 U1069 ( .A(KEYINPUT13), .B(n1157), .ZN(n1394) );
NAND3_X1 U1070 ( .A1(n1397), .A2(n1240), .A3(n1396), .ZN(n1157) );
XOR2_X1 U1071 ( .A(n1368), .B(KEYINPUT44), .Z(n1396) );
INV_X1 U1072 ( .A(G469), .ZN(n1240) );
XOR2_X1 U1073 ( .A(n1398), .B(n1399), .Z(n1397) );
XOR2_X1 U1074 ( .A(n1257), .B(n1192), .Z(n1399) );
NAND2_X1 U1075 ( .A1(n1400), .A2(n1401), .ZN(n1192) );
NAND2_X1 U1076 ( .A1(n1402), .A2(G146), .ZN(n1401) );
NAND2_X1 U1077 ( .A1(n1403), .A2(n1404), .ZN(n1400) );
XNOR2_X1 U1078 ( .A(n1402), .B(KEYINPUT61), .ZN(n1403) );
XOR2_X1 U1079 ( .A(n1191), .B(n1405), .Z(n1257) );
XOR2_X1 U1080 ( .A(n1406), .B(n1259), .Z(n1398) );
XNOR2_X1 U1081 ( .A(n1197), .B(n1196), .ZN(n1259) );
XOR2_X1 U1082 ( .A(G131), .B(G134), .Z(n1196) );
INV_X1 U1083 ( .A(G137), .ZN(n1197) );
XOR2_X1 U1084 ( .A(n1254), .B(n1407), .Z(n1406) );
NOR2_X1 U1085 ( .A1(KEYINPUT63), .A2(n1261), .ZN(n1407) );
NAND2_X1 U1086 ( .A1(G227), .A2(n1177), .ZN(n1254) );
NOR2_X1 U1087 ( .A1(n1330), .A2(n1329), .ZN(n1122) );
INV_X1 U1088 ( .A(n1354), .ZN(n1329) );
NOR2_X1 U1089 ( .A1(n1154), .A2(n1408), .ZN(n1354) );
NOR2_X1 U1090 ( .A1(n1169), .A2(n1170), .ZN(n1408) );
INV_X1 U1091 ( .A(n1409), .ZN(n1170) );
INV_X1 U1092 ( .A(G475), .ZN(n1169) );
NOR2_X1 U1093 ( .A1(n1409), .A2(G475), .ZN(n1154) );
NAND2_X1 U1094 ( .A1(n1222), .A2(n1368), .ZN(n1409) );
XOR2_X1 U1095 ( .A(n1410), .B(n1411), .Z(n1222) );
XOR2_X1 U1096 ( .A(n1412), .B(n1374), .Z(n1411) );
XOR2_X1 U1097 ( .A(n1187), .B(n1413), .Z(n1374) );
XOR2_X1 U1098 ( .A(KEYINPUT26), .B(G146), .Z(n1413) );
NAND2_X1 U1099 ( .A1(KEYINPUT62), .A2(n1191), .ZN(n1412) );
INV_X1 U1100 ( .A(G140), .ZN(n1191) );
XOR2_X1 U1101 ( .A(n1414), .B(n1415), .Z(n1410) );
NOR2_X1 U1102 ( .A1(n1416), .A2(n1417), .ZN(n1415) );
XOR2_X1 U1103 ( .A(n1418), .B(KEYINPUT34), .Z(n1417) );
NAND2_X1 U1104 ( .A1(G104), .A2(n1419), .ZN(n1418) );
XOR2_X1 U1105 ( .A(KEYINPUT14), .B(n1420), .Z(n1419) );
NOR2_X1 U1106 ( .A1(G104), .A2(n1420), .ZN(n1416) );
XOR2_X1 U1107 ( .A(G113), .B(G122), .Z(n1420) );
XOR2_X1 U1108 ( .A(n1421), .B(n1422), .Z(n1414) );
NOR2_X1 U1109 ( .A1(KEYINPUT59), .A2(n1423), .ZN(n1422) );
XOR2_X1 U1110 ( .A(G143), .B(n1424), .Z(n1423) );
AND3_X1 U1111 ( .A1(G214), .A2(n1177), .A3(n1390), .ZN(n1424) );
INV_X1 U1112 ( .A(G131), .ZN(n1421) );
NAND2_X1 U1113 ( .A1(n1425), .A2(n1426), .ZN(n1330) );
NAND2_X1 U1114 ( .A1(G478), .A2(n1161), .ZN(n1426) );
XOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1427), .Z(n1425) );
NOR2_X1 U1116 ( .A1(G478), .A2(n1161), .ZN(n1427) );
INV_X1 U1117 ( .A(n1215), .ZN(n1161) );
NOR2_X1 U1118 ( .A1(n1218), .A2(G902), .ZN(n1215) );
XOR2_X1 U1119 ( .A(n1428), .B(n1429), .Z(n1218) );
XOR2_X1 U1120 ( .A(G116), .B(n1430), .Z(n1429) );
XOR2_X1 U1121 ( .A(G134), .B(G122), .Z(n1430) );
XOR2_X1 U1122 ( .A(n1431), .B(n1432), .Z(n1428) );
AND3_X1 U1123 ( .A1(G234), .A2(n1177), .A3(G217), .ZN(n1432) );
XNOR2_X1 U1124 ( .A(G107), .B(n1433), .ZN(n1431) );
NOR2_X1 U1125 ( .A1(KEYINPUT15), .A2(n1434), .ZN(n1433) );
XOR2_X1 U1126 ( .A(G143), .B(n1435), .Z(n1434) );
NOR2_X1 U1127 ( .A1(G128), .A2(KEYINPUT18), .ZN(n1435) );
INV_X1 U1128 ( .A(n1305), .ZN(n1105) );
NAND2_X1 U1129 ( .A1(n1436), .A2(n1143), .ZN(n1305) );
XNOR2_X1 U1130 ( .A(n1437), .B(n1171), .ZN(n1143) );
AND2_X1 U1131 ( .A1(G210), .A2(n1438), .ZN(n1171) );
NAND3_X1 U1132 ( .A1(n1439), .A2(n1368), .A3(KEYINPUT35), .ZN(n1437) );
INV_X1 U1133 ( .A(G902), .ZN(n1368) );
INV_X1 U1134 ( .A(n1173), .ZN(n1439) );
XOR2_X1 U1135 ( .A(n1207), .B(n1440), .Z(n1173) );
XOR2_X1 U1136 ( .A(n1441), .B(n1442), .Z(n1440) );
NOR2_X1 U1137 ( .A1(KEYINPUT2), .A2(n1277), .ZN(n1442) );
NAND2_X1 U1138 ( .A1(G224), .A2(n1177), .ZN(n1277) );
INV_X1 U1139 ( .A(G953), .ZN(n1177) );
NOR3_X1 U1140 ( .A1(n1278), .A2(n1443), .A3(n1444), .ZN(n1441) );
AND2_X1 U1141 ( .A1(KEYINPUT24), .A2(n1279), .ZN(n1444) );
NOR2_X1 U1142 ( .A1(n1187), .A2(n1383), .ZN(n1279) );
NOR2_X1 U1143 ( .A1(KEYINPUT24), .A2(G125), .ZN(n1443) );
AND2_X1 U1144 ( .A1(n1383), .A2(n1187), .ZN(n1278) );
INV_X1 U1145 ( .A(G125), .ZN(n1187) );
XNOR2_X1 U1146 ( .A(n1404), .B(n1402), .ZN(n1383) );
XNOR2_X1 U1147 ( .A(n1337), .B(G143), .ZN(n1402) );
INV_X1 U1148 ( .A(G128), .ZN(n1337) );
INV_X1 U1149 ( .A(G146), .ZN(n1404) );
XOR2_X1 U1150 ( .A(n1445), .B(n1446), .Z(n1207) );
XOR2_X1 U1151 ( .A(n1345), .B(n1447), .Z(n1446) );
NAND2_X1 U1152 ( .A1(n1448), .A2(n1449), .ZN(n1447) );
NAND2_X1 U1153 ( .A1(G113), .A2(n1384), .ZN(n1449) );
XOR2_X1 U1154 ( .A(n1450), .B(KEYINPUT41), .Z(n1448) );
OR2_X1 U1155 ( .A1(n1384), .A2(G113), .ZN(n1450) );
XOR2_X1 U1156 ( .A(G116), .B(G119), .Z(n1384) );
INV_X1 U1157 ( .A(G122), .ZN(n1345) );
XOR2_X1 U1158 ( .A(n1405), .B(n1261), .Z(n1445) );
XOR2_X1 U1159 ( .A(n1451), .B(n1452), .Z(n1261) );
XOR2_X1 U1160 ( .A(G104), .B(G101), .Z(n1452) );
XNOR2_X1 U1161 ( .A(G107), .B(KEYINPUT55), .ZN(n1451) );
XNOR2_X1 U1162 ( .A(n1362), .B(KEYINPUT49), .ZN(n1405) );
INV_X1 U1163 ( .A(G110), .ZN(n1362) );
XOR2_X1 U1164 ( .A(n1142), .B(KEYINPUT51), .Z(n1436) );
NAND2_X1 U1165 ( .A1(G214), .A2(n1438), .ZN(n1142) );
NAND2_X1 U1166 ( .A1(n1393), .A2(n1390), .ZN(n1438) );
INV_X1 U1167 ( .A(G237), .ZN(n1390) );
XOR2_X1 U1168 ( .A(G902), .B(KEYINPUT48), .Z(n1393) );
endmodule


