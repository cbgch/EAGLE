//Key = 1001000001100011010000001000011000001100100001010001001100110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373;

XNOR2_X1 U755 ( .A(G107), .B(n1037), .ZN(G9) );
NOR2_X1 U756 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR4_X1 U757 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NOR3_X1 U758 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NOR2_X1 U759 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U760 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U761 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U762 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
INV_X1 U763 ( .A(n1055), .ZN(n1054) );
XNOR2_X1 U764 ( .A(n1056), .B(KEYINPUT11), .ZN(n1053) );
NOR2_X1 U765 ( .A1(n1057), .A2(n1058), .ZN(n1051) );
NOR2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U768 ( .A1(KEYINPUT4), .A2(n1063), .ZN(n1059) );
NOR3_X1 U769 ( .A1(n1064), .A2(n1065), .A3(n1058), .ZN(n1047) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U772 ( .A1(KEYINPUT25), .A2(n1070), .ZN(n1066) );
NOR3_X1 U773 ( .A1(n1071), .A2(n1072), .A3(n1064), .ZN(n1042) );
NOR4_X1 U774 ( .A1(n1070), .A2(n1058), .A3(n1046), .A4(n1044), .ZN(n1072) );
INV_X1 U775 ( .A(n1073), .ZN(n1046) );
INV_X1 U776 ( .A(KEYINPUT25), .ZN(n1071) );
NAND4_X1 U777 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1040) );
NAND4_X1 U778 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1075) );
NOR2_X1 U779 ( .A1(n1082), .A2(n1050), .ZN(n1080) );
XNOR2_X1 U780 ( .A(n1073), .B(KEYINPUT56), .ZN(n1082) );
XNOR2_X1 U781 ( .A(n1056), .B(KEYINPUT58), .ZN(n1078) );
NAND4_X1 U782 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1074) );
NAND2_X1 U783 ( .A1(n1087), .A2(n1044), .ZN(n1086) );
NAND3_X1 U784 ( .A1(n1073), .A2(n1088), .A3(KEYINPUT4), .ZN(n1087) );
NAND2_X1 U785 ( .A1(n1079), .A2(n1089), .ZN(n1085) );
NAND2_X1 U786 ( .A1(n1056), .A2(n1090), .ZN(n1089) );
OR2_X1 U787 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
INV_X1 U788 ( .A(n1064), .ZN(n1056) );
INV_X1 U789 ( .A(n1044), .ZN(n1079) );
NOR3_X1 U790 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1038) );
INV_X1 U791 ( .A(n1076), .ZN(n1093) );
NAND4_X1 U792 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1076) );
NOR3_X1 U793 ( .A1(n1098), .A2(n1061), .A3(n1099), .ZN(n1097) );
XNOR2_X1 U794 ( .A(n1100), .B(n1101), .ZN(n1099) );
NAND3_X1 U795 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1098) );
XNOR2_X1 U796 ( .A(n1105), .B(n1106), .ZN(n1104) );
OR3_X1 U797 ( .A1(n1107), .A2(KEYINPUT43), .A3(n1108), .ZN(n1103) );
NAND2_X1 U798 ( .A1(n1109), .A2(n1108), .ZN(n1102) );
NAND2_X1 U799 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
INV_X1 U800 ( .A(KEYINPUT43), .ZN(n1111) );
XNOR2_X1 U801 ( .A(n1107), .B(KEYINPUT20), .ZN(n1110) );
NOR3_X1 U802 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1096) );
XOR2_X1 U803 ( .A(n1115), .B(KEYINPUT3), .Z(n1112) );
NAND2_X1 U804 ( .A1(KEYINPUT43), .A2(n1107), .ZN(n1095) );
XOR2_X1 U805 ( .A(n1116), .B(n1117), .Z(G72) );
NOR2_X1 U806 ( .A1(n1118), .A2(n1077), .ZN(n1117) );
AND2_X1 U807 ( .A1(G227), .A2(G900), .ZN(n1118) );
NAND2_X1 U808 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
NAND2_X1 U809 ( .A1(n1121), .A2(n1077), .ZN(n1120) );
XNOR2_X1 U810 ( .A(n1122), .B(n1123), .ZN(n1121) );
NOR3_X1 U811 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
XOR2_X1 U812 ( .A(n1127), .B(KEYINPUT60), .Z(n1126) );
NAND2_X1 U813 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U814 ( .A(n1130), .B(KEYINPUT31), .Z(n1128) );
NAND3_X1 U815 ( .A1(G900), .A2(n1122), .A3(G953), .ZN(n1119) );
XOR2_X1 U816 ( .A(n1131), .B(n1132), .Z(n1122) );
NOR2_X1 U817 ( .A1(KEYINPUT12), .A2(n1133), .ZN(n1132) );
XOR2_X1 U818 ( .A(n1134), .B(n1135), .Z(n1133) );
XNOR2_X1 U819 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR2_X1 U820 ( .A1(KEYINPUT53), .A2(n1138), .ZN(n1137) );
INV_X1 U821 ( .A(n1139), .ZN(n1138) );
XNOR2_X1 U822 ( .A(G131), .B(KEYINPUT27), .ZN(n1134) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(G69) );
NOR3_X1 U824 ( .A1(n1077), .A2(KEYINPUT52), .A3(n1142), .ZN(n1141) );
AND2_X1 U825 ( .A1(G224), .A2(G898), .ZN(n1142) );
NAND2_X1 U826 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
NAND2_X1 U827 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND3_X1 U828 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1143) );
NAND2_X1 U829 ( .A1(G953), .A2(n1150), .ZN(n1148) );
XOR2_X1 U830 ( .A(KEYINPUT14), .B(n1145), .Z(n1147) );
AND2_X1 U831 ( .A1(n1151), .A2(n1077), .ZN(n1145) );
NAND2_X1 U832 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XNOR2_X1 U833 ( .A(KEYINPUT36), .B(n1154), .ZN(n1153) );
NOR2_X1 U834 ( .A1(n1155), .A2(n1156), .ZN(G66) );
NOR3_X1 U835 ( .A1(n1100), .A2(n1157), .A3(n1158), .ZN(n1156) );
NOR3_X1 U836 ( .A1(n1159), .A2(n1101), .A3(n1160), .ZN(n1158) );
NOR2_X1 U837 ( .A1(n1161), .A2(n1162), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1163), .A2(n1101), .ZN(n1161) );
NOR2_X1 U839 ( .A1(n1155), .A2(n1164), .ZN(G63) );
XNOR2_X1 U840 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U841 ( .A1(n1167), .A2(n1160), .ZN(n1166) );
NOR2_X1 U842 ( .A1(n1155), .A2(n1168), .ZN(G60) );
NOR3_X1 U843 ( .A1(n1107), .A2(n1169), .A3(n1170), .ZN(n1168) );
NOR3_X1 U844 ( .A1(n1171), .A2(n1108), .A3(n1160), .ZN(n1170) );
NOR2_X1 U845 ( .A1(n1172), .A2(n1173), .ZN(n1169) );
NOR2_X1 U846 ( .A1(n1163), .A2(n1108), .ZN(n1172) );
INV_X1 U847 ( .A(n1041), .ZN(n1163) );
XOR2_X1 U848 ( .A(n1174), .B(n1175), .Z(G6) );
XOR2_X1 U849 ( .A(KEYINPUT45), .B(G104), .Z(n1175) );
NAND4_X1 U850 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1174) );
NOR2_X1 U851 ( .A1(n1058), .A2(n1180), .ZN(n1179) );
XNOR2_X1 U852 ( .A(KEYINPUT8), .B(n1063), .ZN(n1176) );
INV_X1 U853 ( .A(n1088), .ZN(n1063) );
NOR2_X1 U854 ( .A1(n1155), .A2(n1181), .ZN(G57) );
XOR2_X1 U855 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U856 ( .A(n1184), .B(n1185), .ZN(n1183) );
XNOR2_X1 U857 ( .A(n1186), .B(n1187), .ZN(n1182) );
NOR2_X1 U858 ( .A1(n1188), .A2(n1160), .ZN(n1187) );
NOR2_X1 U859 ( .A1(n1155), .A2(n1189), .ZN(G54) );
XOR2_X1 U860 ( .A(n1190), .B(n1191), .Z(n1189) );
XOR2_X1 U861 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U862 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U863 ( .A1(n1106), .A2(n1160), .ZN(n1195) );
INV_X1 U864 ( .A(G469), .ZN(n1106) );
NOR3_X1 U865 ( .A1(n1196), .A2(KEYINPUT57), .A3(n1197), .ZN(n1194) );
XOR2_X1 U866 ( .A(n1198), .B(KEYINPUT40), .Z(n1196) );
NAND2_X1 U867 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XNOR2_X1 U868 ( .A(G110), .B(KEYINPUT15), .ZN(n1199) );
XOR2_X1 U869 ( .A(n1201), .B(n1202), .Z(n1190) );
XNOR2_X1 U870 ( .A(n1186), .B(n1203), .ZN(n1202) );
XNOR2_X1 U871 ( .A(KEYINPUT61), .B(n1204), .ZN(n1201) );
NOR2_X1 U872 ( .A1(KEYINPUT23), .A2(n1205), .ZN(n1204) );
XNOR2_X1 U873 ( .A(n1139), .B(KEYINPUT21), .ZN(n1205) );
NOR2_X1 U874 ( .A1(n1155), .A2(n1206), .ZN(G51) );
XOR2_X1 U875 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U876 ( .A1(n1209), .A2(n1160), .ZN(n1208) );
NAND2_X1 U877 ( .A1(G902), .A2(n1041), .ZN(n1160) );
NAND4_X1 U878 ( .A1(n1210), .A2(n1152), .A3(n1211), .A4(n1212), .ZN(n1041) );
AND3_X1 U879 ( .A1(n1129), .A2(n1154), .A3(n1130), .ZN(n1212) );
NOR3_X1 U880 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1129) );
XNOR2_X1 U881 ( .A(n1125), .B(KEYINPUT35), .ZN(n1211) );
AND4_X1 U882 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1152) );
AND4_X1 U883 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1037), .ZN(n1219) );
NAND3_X1 U884 ( .A1(n1092), .A2(n1084), .A3(n1223), .ZN(n1037) );
NAND2_X1 U885 ( .A1(n1088), .A2(n1224), .ZN(n1218) );
XOR2_X1 U886 ( .A(KEYINPUT16), .B(n1225), .Z(n1224) );
NAND3_X1 U887 ( .A1(n1223), .A2(n1084), .A3(n1091), .ZN(n1216) );
INV_X1 U888 ( .A(n1124), .ZN(n1210) );
NAND3_X1 U889 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1124) );
NAND3_X1 U890 ( .A1(n1091), .A2(n1081), .A3(n1229), .ZN(n1228) );
NOR2_X1 U891 ( .A1(n1230), .A2(n1231), .ZN(n1207) );
XOR2_X1 U892 ( .A(n1232), .B(KEYINPUT9), .Z(n1231) );
NAND2_X1 U893 ( .A1(n1233), .A2(n1149), .ZN(n1232) );
NOR2_X1 U894 ( .A1(n1149), .A2(n1233), .ZN(n1230) );
XOR2_X1 U895 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND2_X1 U896 ( .A1(KEYINPUT59), .A2(n1236), .ZN(n1235) );
XOR2_X1 U897 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U898 ( .A(n1239), .B(KEYINPUT18), .ZN(n1238) );
INV_X1 U899 ( .A(n1146), .ZN(n1149) );
NOR2_X1 U900 ( .A1(n1077), .A2(G952), .ZN(n1155) );
XOR2_X1 U901 ( .A(G146), .B(n1215), .Z(G48) );
AND2_X1 U902 ( .A1(n1240), .A2(n1091), .ZN(n1215) );
XNOR2_X1 U903 ( .A(G143), .B(n1130), .ZN(G45) );
NAND4_X1 U904 ( .A1(n1088), .A2(n1178), .A3(n1081), .A4(n1241), .ZN(n1130) );
NOR3_X1 U905 ( .A1(n1094), .A2(n1242), .A3(n1243), .ZN(n1241) );
XNOR2_X1 U906 ( .A(n1200), .B(n1213), .ZN(G42) );
AND3_X1 U907 ( .A1(n1091), .A2(n1055), .A3(n1229), .ZN(n1213) );
XNOR2_X1 U908 ( .A(n1244), .B(n1214), .ZN(G39) );
AND3_X1 U909 ( .A1(n1073), .A2(n1245), .A3(n1229), .ZN(n1214) );
XNOR2_X1 U910 ( .A(G134), .B(n1226), .ZN(G36) );
NAND3_X1 U911 ( .A1(n1081), .A2(n1092), .A3(n1229), .ZN(n1226) );
XNOR2_X1 U912 ( .A(G131), .B(n1246), .ZN(G33) );
NAND4_X1 U913 ( .A1(n1247), .A2(n1229), .A3(n1091), .A4(n1081), .ZN(n1246) );
NOR3_X1 U914 ( .A1(n1070), .A2(n1242), .A3(n1064), .ZN(n1229) );
NAND2_X1 U915 ( .A1(n1248), .A2(n1249), .ZN(n1064) );
XNOR2_X1 U916 ( .A(n1113), .B(KEYINPUT1), .ZN(n1248) );
INV_X1 U917 ( .A(n1250), .ZN(n1242) );
INV_X1 U918 ( .A(n1178), .ZN(n1070) );
XNOR2_X1 U919 ( .A(KEYINPUT22), .B(KEYINPUT2), .ZN(n1247) );
XOR2_X1 U920 ( .A(G128), .B(n1125), .Z(G30) );
AND2_X1 U921 ( .A1(n1240), .A2(n1092), .ZN(n1125) );
AND4_X1 U922 ( .A1(n1245), .A2(n1088), .A3(n1178), .A4(n1250), .ZN(n1240) );
XNOR2_X1 U923 ( .A(G101), .B(n1217), .ZN(G3) );
NAND3_X1 U924 ( .A1(n1073), .A2(n1223), .A3(n1081), .ZN(n1217) );
NAND3_X1 U925 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(G27) );
OR2_X1 U926 ( .A1(G125), .A2(KEYINPUT30), .ZN(n1253) );
NAND3_X1 U927 ( .A1(KEYINPUT30), .A2(G125), .A3(n1227), .ZN(n1252) );
NAND2_X1 U928 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
NAND2_X1 U929 ( .A1(KEYINPUT30), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U930 ( .A(KEYINPUT6), .B(n1257), .ZN(n1256) );
INV_X1 U931 ( .A(n1227), .ZN(n1254) );
NAND4_X1 U932 ( .A1(n1055), .A2(n1250), .A3(n1088), .A4(n1258), .ZN(n1227) );
NOR2_X1 U933 ( .A1(n1050), .A2(n1180), .ZN(n1258) );
INV_X1 U934 ( .A(n1091), .ZN(n1180) );
INV_X1 U935 ( .A(n1083), .ZN(n1050) );
NAND2_X1 U936 ( .A1(n1044), .A2(n1259), .ZN(n1250) );
NAND4_X1 U937 ( .A1(n1260), .A2(G953), .A3(n1261), .A4(n1262), .ZN(n1259) );
INV_X1 U938 ( .A(G900), .ZN(n1262) );
XNOR2_X1 U939 ( .A(G902), .B(KEYINPUT17), .ZN(n1260) );
XNOR2_X1 U940 ( .A(G122), .B(n1222), .ZN(G24) );
NAND4_X1 U941 ( .A1(n1263), .A2(n1084), .A3(n1264), .A4(n1265), .ZN(n1222) );
INV_X1 U942 ( .A(n1058), .ZN(n1084) );
NAND2_X1 U943 ( .A1(n1115), .A2(n1266), .ZN(n1058) );
XNOR2_X1 U944 ( .A(G119), .B(n1154), .ZN(G21) );
NAND3_X1 U945 ( .A1(n1263), .A2(n1245), .A3(n1073), .ZN(n1154) );
XOR2_X1 U946 ( .A(n1267), .B(n1268), .Z(G18) );
NAND2_X1 U947 ( .A1(n1225), .A2(n1088), .ZN(n1268) );
AND4_X1 U948 ( .A1(n1081), .A2(n1083), .A3(n1092), .A4(n1177), .ZN(n1225) );
NOR2_X1 U949 ( .A1(n1265), .A2(n1094), .ZN(n1092) );
INV_X1 U950 ( .A(n1264), .ZN(n1094) );
NAND2_X1 U951 ( .A1(KEYINPUT10), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U952 ( .A(KEYINPUT46), .B(n1270), .ZN(n1269) );
XNOR2_X1 U953 ( .A(G113), .B(n1221), .ZN(G15) );
NAND3_X1 U954 ( .A1(n1081), .A2(n1263), .A3(n1091), .ZN(n1221) );
NOR2_X1 U955 ( .A1(n1264), .A2(n1243), .ZN(n1091) );
AND3_X1 U956 ( .A1(n1088), .A2(n1177), .A3(n1083), .ZN(n1263) );
NOR2_X1 U957 ( .A1(n1068), .A2(n1114), .ZN(n1083) );
NOR2_X1 U958 ( .A1(n1271), .A2(n1115), .ZN(n1081) );
XNOR2_X1 U959 ( .A(G110), .B(n1220), .ZN(G12) );
NAND3_X1 U960 ( .A1(n1223), .A2(n1055), .A3(n1073), .ZN(n1220) );
NOR2_X1 U961 ( .A1(n1264), .A2(n1265), .ZN(n1073) );
INV_X1 U962 ( .A(n1243), .ZN(n1265) );
XOR2_X1 U963 ( .A(n1107), .B(n1108), .Z(n1243) );
INV_X1 U964 ( .A(G475), .ZN(n1108) );
NOR2_X1 U965 ( .A1(n1173), .A2(G902), .ZN(n1107) );
INV_X1 U966 ( .A(n1171), .ZN(n1173) );
XNOR2_X1 U967 ( .A(n1272), .B(n1273), .ZN(n1171) );
XOR2_X1 U968 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U969 ( .A(n1276), .B(n1131), .Z(n1275) );
XOR2_X1 U970 ( .A(G125), .B(G140), .Z(n1131) );
NAND2_X1 U971 ( .A1(n1277), .A2(G214), .ZN(n1276) );
XOR2_X1 U972 ( .A(n1278), .B(G104), .Z(n1274) );
NAND2_X1 U973 ( .A1(KEYINPUT47), .A2(n1279), .ZN(n1278) );
XOR2_X1 U974 ( .A(G122), .B(G113), .Z(n1279) );
XOR2_X1 U975 ( .A(n1280), .B(n1281), .Z(n1272) );
XOR2_X1 U976 ( .A(G143), .B(G131), .Z(n1281) );
XNOR2_X1 U977 ( .A(G146), .B(KEYINPUT39), .ZN(n1280) );
XOR2_X1 U978 ( .A(n1282), .B(n1167), .Z(n1264) );
INV_X1 U979 ( .A(G478), .ZN(n1167) );
NAND2_X1 U980 ( .A1(n1165), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U981 ( .A(n1284), .B(n1285), .ZN(n1165) );
XOR2_X1 U982 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U983 ( .A(G128), .B(G122), .Z(n1287) );
XOR2_X1 U984 ( .A(G143), .B(G134), .Z(n1286) );
XOR2_X1 U985 ( .A(n1288), .B(n1289), .Z(n1284) );
XNOR2_X1 U986 ( .A(n1270), .B(G107), .ZN(n1289) );
NAND2_X1 U987 ( .A1(G217), .A2(n1290), .ZN(n1288) );
NAND2_X1 U988 ( .A1(n1291), .A2(n1292), .ZN(n1055) );
NAND3_X1 U989 ( .A1(n1115), .A2(n1271), .A3(n1293), .ZN(n1292) );
INV_X1 U990 ( .A(KEYINPUT50), .ZN(n1293) );
INV_X1 U991 ( .A(n1266), .ZN(n1271) );
NAND2_X1 U992 ( .A1(KEYINPUT50), .A2(n1245), .ZN(n1291) );
NOR2_X1 U993 ( .A1(n1266), .A2(n1115), .ZN(n1245) );
XNOR2_X1 U994 ( .A(n1294), .B(n1188), .ZN(n1115) );
INV_X1 U995 ( .A(G472), .ZN(n1188) );
NAND2_X1 U996 ( .A1(n1295), .A2(n1283), .ZN(n1294) );
XNOR2_X1 U997 ( .A(n1296), .B(n1297), .ZN(n1295) );
XNOR2_X1 U998 ( .A(n1298), .B(KEYINPUT62), .ZN(n1297) );
NAND2_X1 U999 ( .A1(KEYINPUT55), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U1000 ( .A(n1186), .B(n1300), .ZN(n1299) );
NAND2_X1 U1001 ( .A1(KEYINPUT54), .A2(n1185), .ZN(n1300) );
INV_X1 U1002 ( .A(n1239), .ZN(n1185) );
INV_X1 U1003 ( .A(n1301), .ZN(n1186) );
INV_X1 U1004 ( .A(n1184), .ZN(n1296) );
XNOR2_X1 U1005 ( .A(n1302), .B(n1303), .ZN(n1184) );
XNOR2_X1 U1006 ( .A(n1270), .B(n1304), .ZN(n1303) );
XOR2_X1 U1007 ( .A(KEYINPUT37), .B(G119), .Z(n1304) );
XOR2_X1 U1008 ( .A(n1305), .B(n1306), .Z(n1302) );
XOR2_X1 U1009 ( .A(n1307), .B(G101), .Z(n1305) );
NAND2_X1 U1010 ( .A1(n1277), .A2(G210), .ZN(n1307) );
NOR2_X1 U1011 ( .A1(G953), .A2(G237), .ZN(n1277) );
XOR2_X1 U1012 ( .A(n1100), .B(n1308), .Z(n1266) );
NOR2_X1 U1013 ( .A1(n1309), .A2(KEYINPUT7), .ZN(n1308) );
INV_X1 U1014 ( .A(n1101), .ZN(n1309) );
NAND2_X1 U1015 ( .A1(G217), .A2(n1310), .ZN(n1101) );
NOR2_X1 U1016 ( .A1(n1162), .A2(G902), .ZN(n1100) );
INV_X1 U1017 ( .A(n1159), .ZN(n1162) );
NAND2_X1 U1018 ( .A1(n1311), .A2(n1312), .ZN(n1159) );
NAND2_X1 U1019 ( .A1(n1313), .A2(n1244), .ZN(n1312) );
NAND2_X1 U1020 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND2_X1 U1021 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
INV_X1 U1022 ( .A(n1318), .ZN(n1316) );
NAND2_X1 U1023 ( .A1(n1318), .A2(n1319), .ZN(n1314) );
XNOR2_X1 U1024 ( .A(n1320), .B(KEYINPUT48), .ZN(n1318) );
NAND2_X1 U1025 ( .A1(G137), .A2(n1321), .ZN(n1311) );
NAND2_X1 U1026 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NAND2_X1 U1027 ( .A1(n1324), .A2(n1317), .ZN(n1323) );
NAND2_X1 U1028 ( .A1(n1319), .A2(n1325), .ZN(n1322) );
INV_X1 U1029 ( .A(n1324), .ZN(n1325) );
XNOR2_X1 U1030 ( .A(n1320), .B(KEYINPUT44), .ZN(n1324) );
NAND2_X1 U1031 ( .A1(n1290), .A2(G221), .ZN(n1320) );
AND2_X1 U1032 ( .A1(G234), .A2(n1077), .ZN(n1290) );
XOR2_X1 U1033 ( .A(n1317), .B(KEYINPUT51), .Z(n1319) );
XOR2_X1 U1034 ( .A(n1326), .B(n1327), .Z(n1317) );
XOR2_X1 U1035 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U1036 ( .A(KEYINPUT41), .B(n1330), .ZN(n1326) );
NOR2_X1 U1037 ( .A1(KEYINPUT34), .A2(n1331), .ZN(n1330) );
XNOR2_X1 U1038 ( .A(n1200), .B(n1332), .ZN(n1331) );
NOR2_X1 U1039 ( .A1(KEYINPUT33), .A2(n1257), .ZN(n1332) );
INV_X1 U1040 ( .A(G125), .ZN(n1257) );
AND3_X1 U1041 ( .A1(n1178), .A2(n1177), .A3(n1088), .ZN(n1223) );
NOR2_X1 U1042 ( .A1(n1249), .A2(n1113), .ZN(n1088) );
INV_X1 U1043 ( .A(n1062), .ZN(n1113) );
NAND2_X1 U1044 ( .A1(G214), .A2(n1333), .ZN(n1062) );
INV_X1 U1045 ( .A(n1061), .ZN(n1249) );
XOR2_X1 U1046 ( .A(n1334), .B(n1209), .Z(n1061) );
NAND2_X1 U1047 ( .A1(G210), .A2(n1333), .ZN(n1209) );
NAND2_X1 U1048 ( .A1(n1335), .A2(n1283), .ZN(n1333) );
INV_X1 U1049 ( .A(G237), .ZN(n1335) );
NAND2_X1 U1050 ( .A1(n1336), .A2(n1283), .ZN(n1334) );
XNOR2_X1 U1051 ( .A(n1146), .B(n1337), .ZN(n1336) );
XNOR2_X1 U1052 ( .A(n1338), .B(n1234), .ZN(n1337) );
NAND2_X1 U1053 ( .A1(G224), .A2(n1077), .ZN(n1234) );
NAND2_X1 U1054 ( .A1(n1339), .A2(KEYINPUT24), .ZN(n1338) );
XOR2_X1 U1055 ( .A(n1237), .B(n1340), .Z(n1339) );
NOR2_X1 U1056 ( .A1(KEYINPUT42), .A2(n1239), .ZN(n1340) );
XOR2_X1 U1057 ( .A(n1139), .B(KEYINPUT26), .Z(n1239) );
XNOR2_X1 U1058 ( .A(G125), .B(KEYINPUT28), .ZN(n1237) );
XNOR2_X1 U1059 ( .A(n1341), .B(n1342), .ZN(n1146) );
XOR2_X1 U1060 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1061 ( .A(G122), .B(G101), .Z(n1344) );
NOR2_X1 U1062 ( .A1(KEYINPUT13), .A2(n1345), .ZN(n1343) );
XOR2_X1 U1063 ( .A(n1346), .B(n1306), .Z(n1341) );
XOR2_X1 U1064 ( .A(G113), .B(KEYINPUT63), .Z(n1306) );
NAND2_X1 U1065 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NAND2_X1 U1066 ( .A1(n1349), .A2(n1270), .ZN(n1348) );
INV_X1 U1067 ( .A(G116), .ZN(n1270) );
XOR2_X1 U1068 ( .A(KEYINPUT49), .B(n1329), .Z(n1349) );
NAND2_X1 U1069 ( .A1(n1350), .A2(G116), .ZN(n1347) );
XOR2_X1 U1070 ( .A(KEYINPUT29), .B(n1329), .Z(n1350) );
XOR2_X1 U1071 ( .A(G119), .B(G110), .Z(n1329) );
NAND2_X1 U1072 ( .A1(n1044), .A2(n1351), .ZN(n1177) );
NAND4_X1 U1073 ( .A1(G953), .A2(G902), .A3(n1261), .A4(n1150), .ZN(n1351) );
INV_X1 U1074 ( .A(G898), .ZN(n1150) );
NAND3_X1 U1075 ( .A1(n1261), .A2(n1077), .A3(G952), .ZN(n1044) );
NAND2_X1 U1076 ( .A1(G237), .A2(G234), .ZN(n1261) );
NOR2_X1 U1077 ( .A1(n1352), .A2(n1114), .ZN(n1178) );
INV_X1 U1078 ( .A(n1069), .ZN(n1114) );
NAND2_X1 U1079 ( .A1(G221), .A2(n1310), .ZN(n1069) );
NAND2_X1 U1080 ( .A1(G234), .A2(n1283), .ZN(n1310) );
INV_X1 U1081 ( .A(n1068), .ZN(n1352) );
XOR2_X1 U1082 ( .A(G469), .B(n1353), .Z(n1068) );
NOR2_X1 U1083 ( .A1(KEYINPUT19), .A2(n1105), .ZN(n1353) );
NAND3_X1 U1084 ( .A1(n1354), .A2(n1355), .A3(n1283), .ZN(n1105) );
INV_X1 U1085 ( .A(G902), .ZN(n1283) );
NAND2_X1 U1086 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
INV_X1 U1087 ( .A(KEYINPUT32), .ZN(n1357) );
XOR2_X1 U1088 ( .A(n1358), .B(n1359), .Z(n1356) );
NAND2_X1 U1089 ( .A1(KEYINPUT0), .A2(n1360), .ZN(n1359) );
NAND3_X1 U1090 ( .A1(n1361), .A2(n1358), .A3(KEYINPUT32), .ZN(n1354) );
NAND3_X1 U1091 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1358) );
NAND2_X1 U1092 ( .A1(n1197), .A2(n1365), .ZN(n1364) );
NOR2_X1 U1093 ( .A1(n1200), .A2(G110), .ZN(n1197) );
NAND3_X1 U1094 ( .A1(n1203), .A2(G110), .A3(G140), .ZN(n1363) );
INV_X1 U1095 ( .A(n1365), .ZN(n1203) );
NAND2_X1 U1096 ( .A1(n1366), .A2(n1200), .ZN(n1362) );
INV_X1 U1097 ( .A(G140), .ZN(n1200) );
XNOR2_X1 U1098 ( .A(G110), .B(n1365), .ZN(n1366) );
NAND2_X1 U1099 ( .A1(G227), .A2(n1077), .ZN(n1365) );
INV_X1 U1100 ( .A(G953), .ZN(n1077) );
INV_X1 U1101 ( .A(n1360), .ZN(n1361) );
XOR2_X1 U1102 ( .A(n1367), .B(n1301), .Z(n1360) );
NAND2_X1 U1103 ( .A1(n1368), .A2(n1369), .ZN(n1301) );
NAND2_X1 U1104 ( .A1(G131), .A2(n1136), .ZN(n1369) );
XOR2_X1 U1105 ( .A(n1370), .B(KEYINPUT38), .Z(n1368) );
OR2_X1 U1106 ( .A1(n1136), .A2(G131), .ZN(n1370) );
XNOR2_X1 U1107 ( .A(G134), .B(n1244), .ZN(n1136) );
INV_X1 U1108 ( .A(G137), .ZN(n1244) );
NAND2_X1 U1109 ( .A1(n1371), .A2(n1372), .ZN(n1367) );
OR2_X1 U1110 ( .A1(n1192), .A2(n1139), .ZN(n1372) );
XOR2_X1 U1111 ( .A(n1373), .B(KEYINPUT5), .Z(n1371) );
NAND2_X1 U1112 ( .A1(n1192), .A2(n1139), .ZN(n1373) );
XOR2_X1 U1113 ( .A(G143), .B(n1328), .Z(n1139) );
XOR2_X1 U1114 ( .A(G128), .B(G146), .Z(n1328) );
XNOR2_X1 U1115 ( .A(G101), .B(n1345), .ZN(n1192) );
XNOR2_X1 U1116 ( .A(G104), .B(G107), .ZN(n1345) );
endmodule


