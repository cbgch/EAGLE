//Key = 1010000000101101101000011100010000101011000001010000010011101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;

XNOR2_X1 U737 ( .A(G107), .B(n1029), .ZN(G9) );
NOR2_X1 U738 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NAND3_X1 U740 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1032) );
NAND4_X1 U741 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1038) );
NAND2_X1 U742 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U743 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1043) );
NAND3_X1 U744 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1041) );
NAND4_X1 U745 ( .A1(KEYINPUT33), .A2(n1045), .A3(n1051), .A4(n1052), .ZN(n1049) );
NAND2_X1 U746 ( .A1(n1047), .A2(n1053), .ZN(n1048) );
NAND2_X1 U747 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND3_X1 U748 ( .A1(n1056), .A2(n1045), .A3(n1057), .ZN(n1055) );
NAND2_X1 U749 ( .A1(n1046), .A2(n1058), .ZN(n1054) );
NAND2_X1 U750 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U751 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND4_X1 U752 ( .A1(n1063), .A2(n1047), .A3(n1045), .A4(n1050), .ZN(n1036) );
NOR2_X1 U753 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U754 ( .A1(n1039), .A2(n1066), .ZN(n1065) );
NOR2_X1 U755 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U756 ( .A1(n1069), .A2(n1052), .ZN(n1064) );
NAND3_X1 U757 ( .A1(n1070), .A2(n1071), .A3(n1047), .ZN(n1052) );
OR3_X1 U758 ( .A1(n1067), .A2(KEYINPUT33), .A3(n1072), .ZN(n1071) );
NAND2_X1 U759 ( .A1(n1046), .A2(n1073), .ZN(n1070) );
NAND2_X1 U760 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XNOR2_X1 U761 ( .A(n1076), .B(KEYINPUT51), .ZN(n1074) );
NOR3_X1 U762 ( .A1(n1035), .A2(G952), .A3(n1077), .ZN(n1030) );
INV_X1 U763 ( .A(n1037), .ZN(n1077) );
NAND4_X1 U764 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1037) );
NOR4_X1 U765 ( .A1(n1044), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1081) );
XNOR2_X1 U766 ( .A(KEYINPUT54), .B(n1085), .ZN(n1084) );
NOR3_X1 U767 ( .A1(n1086), .A2(n1057), .A3(n1062), .ZN(n1080) );
NAND2_X1 U768 ( .A1(G472), .A2(n1087), .ZN(n1079) );
XNOR2_X1 U769 ( .A(KEYINPUT39), .B(n1056), .ZN(n1078) );
XOR2_X1 U770 ( .A(n1088), .B(n1089), .Z(G72) );
NOR2_X1 U771 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U772 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
XOR2_X1 U773 ( .A(KEYINPUT56), .B(G900), .Z(n1093) );
INV_X1 U774 ( .A(G227), .ZN(n1092) );
NAND2_X1 U775 ( .A1(n1094), .A2(n1095), .ZN(n1088) );
OR2_X1 U776 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U777 ( .A(n1098), .B(KEYINPUT40), .Z(n1094) );
NAND2_X1 U778 ( .A1(n1097), .A2(n1096), .ZN(n1098) );
NAND2_X1 U779 ( .A1(n1099), .A2(n1100), .ZN(n1096) );
NAND2_X1 U780 ( .A1(G953), .A2(n1101), .ZN(n1100) );
XOR2_X1 U781 ( .A(n1102), .B(n1103), .Z(n1099) );
XOR2_X1 U782 ( .A(KEYINPUT22), .B(n1104), .Z(n1103) );
XNOR2_X1 U783 ( .A(n1105), .B(n1106), .ZN(n1102) );
AND2_X1 U784 ( .A1(n1091), .A2(n1033), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1107), .B(n1108), .Z(G69) );
NOR2_X1 U786 ( .A1(n1109), .A2(n1091), .ZN(n1108) );
AND2_X1 U787 ( .A1(G224), .A2(G898), .ZN(n1109) );
NAND2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NAND3_X1 U789 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NAND2_X1 U790 ( .A1(n1115), .A2(n1116), .ZN(n1110) );
NAND2_X1 U791 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U792 ( .A1(KEYINPUT28), .A2(n1112), .ZN(n1118) );
NAND2_X1 U793 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
INV_X1 U794 ( .A(KEYINPUT28), .ZN(n1120) );
NAND2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1119) );
INV_X1 U796 ( .A(KEYINPUT62), .ZN(n1113) );
AND3_X1 U797 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1112) );
XOR2_X1 U798 ( .A(KEYINPUT47), .B(n1124), .Z(n1123) );
NOR2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
AND2_X1 U800 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NAND3_X1 U801 ( .A1(n1128), .A2(n1127), .A3(n1126), .ZN(n1122) );
NAND2_X1 U802 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XNOR2_X1 U803 ( .A(n1131), .B(KEYINPUT26), .ZN(n1129) );
NAND2_X1 U804 ( .A1(G953), .A2(n1132), .ZN(n1121) );
INV_X1 U805 ( .A(n1114), .ZN(n1115) );
NAND2_X1 U806 ( .A1(n1091), .A2(n1034), .ZN(n1114) );
NOR2_X1 U807 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U808 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U809 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U810 ( .A1(n1133), .A2(n1139), .ZN(G63) );
XOR2_X1 U811 ( .A(n1140), .B(n1141), .Z(n1139) );
AND2_X1 U812 ( .A1(G478), .A2(n1142), .ZN(n1140) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1143), .ZN(G60) );
XNOR2_X1 U814 ( .A(n1144), .B(n1145), .ZN(n1143) );
AND2_X1 U815 ( .A1(G475), .A2(n1142), .ZN(n1145) );
XNOR2_X1 U816 ( .A(n1146), .B(n1147), .ZN(G6) );
NAND2_X1 U817 ( .A1(KEYINPUT58), .A2(G104), .ZN(n1147) );
NOR2_X1 U818 ( .A1(n1133), .A2(n1148), .ZN(G57) );
XOR2_X1 U819 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U820 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U821 ( .A1(G472), .A2(n1142), .ZN(n1152) );
NOR2_X1 U822 ( .A1(KEYINPUT30), .A2(n1153), .ZN(n1151) );
XOR2_X1 U823 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U824 ( .A1(KEYINPUT7), .A2(n1156), .ZN(n1154) );
NOR2_X1 U825 ( .A1(n1133), .A2(n1157), .ZN(G54) );
XOR2_X1 U826 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U827 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND2_X1 U828 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
INV_X1 U829 ( .A(n1164), .ZN(n1163) );
XNOR2_X1 U830 ( .A(n1165), .B(KEYINPUT21), .ZN(n1162) );
NAND2_X1 U831 ( .A1(n1166), .A2(n1164), .ZN(n1160) );
XNOR2_X1 U832 ( .A(KEYINPUT52), .B(n1167), .ZN(n1166) );
INV_X1 U833 ( .A(n1165), .ZN(n1167) );
XOR2_X1 U834 ( .A(G110), .B(n1168), .Z(n1165) );
AND2_X1 U835 ( .A1(G469), .A2(n1142), .ZN(n1168) );
NOR2_X1 U836 ( .A1(n1133), .A2(n1169), .ZN(G51) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U838 ( .A(n1172), .B(n1156), .ZN(n1171) );
NAND3_X1 U839 ( .A1(KEYINPUT2), .A2(n1142), .A3(n1173), .ZN(n1172) );
NOR2_X1 U840 ( .A1(KEYINPUT20), .A2(n1174), .ZN(n1173) );
INV_X1 U841 ( .A(n1138), .ZN(n1142) );
NAND2_X1 U842 ( .A1(G902), .A2(n1175), .ZN(n1138) );
OR2_X1 U843 ( .A1(n1033), .A2(n1034), .ZN(n1175) );
NAND4_X1 U844 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1034) );
AND4_X1 U845 ( .A1(n1180), .A2(n1029), .A3(n1181), .A4(n1182), .ZN(n1179) );
NAND3_X1 U846 ( .A1(n1183), .A2(n1184), .A3(n1076), .ZN(n1029) );
NOR2_X1 U847 ( .A1(n1146), .A2(n1185), .ZN(n1178) );
NOR4_X1 U848 ( .A1(n1186), .A2(n1187), .A3(n1067), .A4(n1188), .ZN(n1185) );
NOR2_X1 U849 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
INV_X1 U850 ( .A(KEYINPUT46), .ZN(n1190) );
NOR2_X1 U851 ( .A1(n1051), .A2(n1191), .ZN(n1189) );
NOR2_X1 U852 ( .A1(KEYINPUT46), .A2(n1192), .ZN(n1186) );
NOR3_X1 U853 ( .A1(n1193), .A2(n1194), .A3(n1075), .ZN(n1146) );
NAND4_X1 U854 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1033) );
AND4_X1 U855 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NOR2_X1 U856 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
NOR2_X1 U857 ( .A1(n1068), .A2(n1205), .ZN(n1204) );
NOR2_X1 U858 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
NOR2_X1 U859 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
NOR2_X1 U860 ( .A1(n1072), .A2(n1210), .ZN(n1209) );
NOR2_X1 U861 ( .A1(n1067), .A2(n1211), .ZN(n1208) );
XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n1068), .ZN(n1211) );
NAND4_X1 U863 ( .A1(n1212), .A2(n1075), .A3(n1213), .A4(n1214), .ZN(n1196) );
INV_X1 U864 ( .A(KEYINPUT24), .ZN(n1214) );
NAND2_X1 U865 ( .A1(n1215), .A2(KEYINPUT24), .ZN(n1195) );
XOR2_X1 U866 ( .A(n1216), .B(n1217), .Z(n1170) );
XNOR2_X1 U867 ( .A(n1218), .B(n1219), .ZN(n1217) );
NAND2_X1 U868 ( .A1(KEYINPUT53), .A2(n1220), .ZN(n1216) );
NOR2_X1 U869 ( .A1(n1091), .A2(G952), .ZN(n1133) );
INV_X1 U870 ( .A(G953), .ZN(n1091) );
XNOR2_X1 U871 ( .A(n1202), .B(n1221), .ZN(G48) );
NOR2_X1 U872 ( .A1(KEYINPUT3), .A2(n1222), .ZN(n1221) );
INV_X1 U873 ( .A(G146), .ZN(n1222) );
OR3_X1 U874 ( .A1(n1075), .A2(n1072), .A3(n1207), .ZN(n1202) );
XNOR2_X1 U875 ( .A(G143), .B(n1201), .ZN(G45) );
NAND3_X1 U876 ( .A1(n1223), .A2(n1051), .A3(n1224), .ZN(n1201) );
AND3_X1 U877 ( .A1(n1225), .A2(n1212), .A3(n1082), .ZN(n1224) );
XOR2_X1 U878 ( .A(G140), .B(n1226), .Z(G42) );
NOR2_X1 U879 ( .A1(n1227), .A2(n1068), .ZN(n1226) );
XOR2_X1 U880 ( .A(n1205), .B(KEYINPUT11), .Z(n1227) );
NAND4_X1 U881 ( .A1(n1228), .A2(n1184), .A3(n1212), .A4(n1044), .ZN(n1205) );
XOR2_X1 U882 ( .A(G137), .B(n1229), .Z(G39) );
NOR3_X1 U883 ( .A1(n1207), .A2(n1067), .A3(n1068), .ZN(n1229) );
INV_X1 U884 ( .A(n1040), .ZN(n1067) );
XNOR2_X1 U885 ( .A(G134), .B(n1200), .ZN(G36) );
NAND2_X1 U886 ( .A1(n1230), .A2(n1076), .ZN(n1200) );
XNOR2_X1 U887 ( .A(G131), .B(n1199), .ZN(G33) );
NAND2_X1 U888 ( .A1(n1228), .A2(n1230), .ZN(n1199) );
NOR3_X1 U889 ( .A1(n1068), .A2(n1231), .A3(n1188), .ZN(n1230) );
INV_X1 U890 ( .A(n1046), .ZN(n1068) );
NOR2_X1 U891 ( .A1(n1232), .A2(n1057), .ZN(n1046) );
XNOR2_X1 U892 ( .A(n1233), .B(n1234), .ZN(G30) );
NOR3_X1 U893 ( .A1(n1235), .A2(n1210), .A3(n1207), .ZN(n1234) );
OR4_X1 U894 ( .A1(n1059), .A2(n1231), .A3(n1039), .A4(n1050), .ZN(n1207) );
INV_X1 U895 ( .A(n1212), .ZN(n1231) );
INV_X1 U896 ( .A(n1076), .ZN(n1210) );
XNOR2_X1 U897 ( .A(KEYINPUT25), .B(n1072), .ZN(n1235) );
XOR2_X1 U898 ( .A(G101), .B(n1236), .Z(G3) );
NOR2_X1 U899 ( .A1(n1188), .A2(n1237), .ZN(n1236) );
INV_X1 U900 ( .A(n1223), .ZN(n1188) );
NOR3_X1 U901 ( .A1(n1044), .A2(n1039), .A3(n1059), .ZN(n1223) );
XNOR2_X1 U902 ( .A(n1219), .B(n1215), .ZN(G27) );
AND3_X1 U903 ( .A1(n1228), .A2(n1212), .A3(n1213), .ZN(n1215) );
NOR4_X1 U904 ( .A1(n1238), .A2(n1069), .A3(n1072), .A4(n1050), .ZN(n1213) );
NAND2_X1 U905 ( .A1(n1239), .A2(n1240), .ZN(n1212) );
NAND3_X1 U906 ( .A1(G902), .A2(n1101), .A3(n1241), .ZN(n1240) );
XOR2_X1 U907 ( .A(KEYINPUT29), .B(G900), .Z(n1101) );
XNOR2_X1 U908 ( .A(G122), .B(n1176), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1225), .A2(n1082), .A3(n1039), .A4(n1242), .ZN(n1176) );
NOR2_X1 U910 ( .A1(n1193), .A2(n1238), .ZN(n1242) );
NAND2_X1 U911 ( .A1(n1243), .A2(n1244), .ZN(G21) );
NAND2_X1 U912 ( .A1(G119), .A2(n1177), .ZN(n1244) );
XOR2_X1 U913 ( .A(n1245), .B(KEYINPUT4), .Z(n1243) );
OR2_X1 U914 ( .A1(n1177), .A2(G119), .ZN(n1245) );
OR4_X1 U915 ( .A1(n1237), .A2(n1238), .A3(n1039), .A4(n1050), .ZN(n1177) );
XNOR2_X1 U916 ( .A(G116), .B(n1180), .ZN(G18) );
NAND4_X1 U917 ( .A1(n1045), .A2(n1076), .A3(n1183), .A4(n1069), .ZN(n1180) );
XNOR2_X1 U918 ( .A(G113), .B(n1182), .ZN(G15) );
NAND4_X1 U919 ( .A1(n1045), .A2(n1228), .A3(n1183), .A4(n1069), .ZN(n1182) );
INV_X1 U920 ( .A(n1193), .ZN(n1183) );
NAND2_X1 U921 ( .A1(n1192), .A2(n1050), .ZN(n1193) );
INV_X1 U922 ( .A(n1075), .ZN(n1228) );
NAND2_X1 U923 ( .A1(n1246), .A2(n1082), .ZN(n1075) );
XNOR2_X1 U924 ( .A(KEYINPUT27), .B(n1225), .ZN(n1246) );
INV_X1 U925 ( .A(n1238), .ZN(n1045) );
NAND2_X1 U926 ( .A1(n1247), .A2(n1061), .ZN(n1238) );
INV_X1 U927 ( .A(n1083), .ZN(n1061) );
XNOR2_X1 U928 ( .A(G110), .B(n1181), .ZN(G12) );
OR3_X1 U929 ( .A1(n1194), .A2(n1050), .A3(n1237), .ZN(n1181) );
NAND2_X1 U930 ( .A1(n1192), .A2(n1040), .ZN(n1237) );
NAND2_X1 U931 ( .A1(n1248), .A2(n1249), .ZN(n1040) );
OR3_X1 U932 ( .A1(n1082), .A2(n1225), .A3(KEYINPUT27), .ZN(n1249) );
NAND2_X1 U933 ( .A1(KEYINPUT27), .A2(n1076), .ZN(n1248) );
NOR2_X1 U934 ( .A1(n1082), .A2(n1085), .ZN(n1076) );
INV_X1 U935 ( .A(n1225), .ZN(n1085) );
XNOR2_X1 U936 ( .A(n1250), .B(G478), .ZN(n1225) );
OR2_X1 U937 ( .A1(n1141), .A2(G902), .ZN(n1250) );
XNOR2_X1 U938 ( .A(n1251), .B(n1252), .ZN(n1141) );
XNOR2_X1 U939 ( .A(n1253), .B(n1254), .ZN(n1252) );
NOR3_X1 U940 ( .A1(n1137), .A2(KEYINPUT55), .A3(n1255), .ZN(n1254) );
NAND2_X1 U941 ( .A1(n1256), .A2(KEYINPUT16), .ZN(n1253) );
XNOR2_X1 U942 ( .A(G128), .B(G143), .ZN(n1256) );
XOR2_X1 U943 ( .A(n1257), .B(n1258), .Z(n1251) );
XOR2_X1 U944 ( .A(KEYINPUT35), .B(G134), .Z(n1258) );
NAND2_X1 U945 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND2_X1 U946 ( .A1(G107), .A2(n1261), .ZN(n1260) );
XOR2_X1 U947 ( .A(KEYINPUT60), .B(n1262), .Z(n1259) );
NOR2_X1 U948 ( .A1(G107), .A2(n1261), .ZN(n1262) );
XNOR2_X1 U949 ( .A(n1263), .B(G116), .ZN(n1261) );
XNOR2_X1 U950 ( .A(n1264), .B(G475), .ZN(n1082) );
NAND2_X1 U951 ( .A1(n1144), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U952 ( .A(n1266), .B(n1267), .ZN(n1144) );
XOR2_X1 U953 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U954 ( .A(G104), .B(n1270), .Z(n1269) );
NOR2_X1 U955 ( .A1(KEYINPUT31), .A2(n1271), .ZN(n1270) );
XNOR2_X1 U956 ( .A(G143), .B(n1272), .ZN(n1271) );
NAND3_X1 U957 ( .A1(n1273), .A2(n1274), .A3(G214), .ZN(n1272) );
XOR2_X1 U958 ( .A(KEYINPUT17), .B(n1275), .Z(n1273) );
XNOR2_X1 U959 ( .A(KEYINPUT43), .B(n1276), .ZN(n1268) );
INV_X1 U960 ( .A(G131), .ZN(n1276) );
XOR2_X1 U961 ( .A(n1277), .B(n1278), .Z(n1266) );
XNOR2_X1 U962 ( .A(n1279), .B(n1280), .ZN(n1278) );
NOR2_X1 U963 ( .A1(KEYINPUT37), .A2(n1105), .ZN(n1280) );
NAND2_X1 U964 ( .A1(KEYINPUT13), .A2(n1281), .ZN(n1279) );
XNOR2_X1 U965 ( .A(n1263), .B(G113), .ZN(n1281) );
NOR2_X1 U966 ( .A1(n1072), .A2(n1191), .ZN(n1192) );
AND2_X1 U967 ( .A1(n1282), .A2(n1239), .ZN(n1191) );
INV_X1 U968 ( .A(n1047), .ZN(n1239) );
NOR3_X1 U969 ( .A1(n1035), .A2(n1283), .A3(n1284), .ZN(n1047) );
INV_X1 U970 ( .A(G952), .ZN(n1284) );
AND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n1283) );
XOR2_X1 U972 ( .A(G953), .B(KEYINPUT63), .Z(n1035) );
NAND3_X1 U973 ( .A1(n1285), .A2(n1132), .A3(n1241), .ZN(n1282) );
AND2_X1 U974 ( .A1(G953), .A2(n1286), .ZN(n1241) );
NAND2_X1 U975 ( .A1(G237), .A2(G234), .ZN(n1286) );
INV_X1 U976 ( .A(G898), .ZN(n1132) );
XNOR2_X1 U977 ( .A(KEYINPUT9), .B(n1265), .ZN(n1285) );
INV_X1 U978 ( .A(n1051), .ZN(n1072) );
NOR2_X1 U979 ( .A1(n1056), .A2(n1057), .ZN(n1051) );
NOR2_X1 U980 ( .A1(n1287), .A2(n1288), .ZN(n1057) );
INV_X1 U981 ( .A(G214), .ZN(n1287) );
INV_X1 U982 ( .A(n1232), .ZN(n1056) );
XNOR2_X1 U983 ( .A(n1289), .B(n1290), .ZN(n1232) );
NOR2_X1 U984 ( .A1(n1288), .A2(n1174), .ZN(n1290) );
INV_X1 U985 ( .A(G210), .ZN(n1174) );
NOR2_X1 U986 ( .A1(G902), .A2(G237), .ZN(n1288) );
NAND2_X1 U987 ( .A1(n1291), .A2(n1265), .ZN(n1289) );
XOR2_X1 U988 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U989 ( .A(n1220), .B(KEYINPUT50), .ZN(n1293) );
AND2_X1 U990 ( .A1(n1294), .A2(n1295), .ZN(n1220) );
NAND3_X1 U991 ( .A1(n1296), .A2(n1127), .A3(n1126), .ZN(n1295) );
NAND2_X1 U992 ( .A1(n1297), .A2(n1131), .ZN(n1127) );
NAND2_X1 U993 ( .A1(n1298), .A2(n1130), .ZN(n1296) );
INV_X1 U994 ( .A(n1131), .ZN(n1298) );
NAND2_X1 U995 ( .A1(n1299), .A2(n1300), .ZN(n1294) );
XNOR2_X1 U996 ( .A(n1131), .B(n1297), .ZN(n1300) );
INV_X1 U997 ( .A(n1130), .ZN(n1297) );
XOR2_X1 U998 ( .A(n1301), .B(n1302), .Z(n1130) );
NOR2_X1 U999 ( .A1(KEYINPUT19), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1000 ( .A(n1304), .B(G101), .Z(n1131) );
XNOR2_X1 U1001 ( .A(n1126), .B(KEYINPUT6), .ZN(n1299) );
XNOR2_X1 U1002 ( .A(n1305), .B(G110), .ZN(n1126) );
NAND2_X1 U1003 ( .A1(n1306), .A2(n1263), .ZN(n1305) );
INV_X1 U1004 ( .A(G122), .ZN(n1263) );
XNOR2_X1 U1005 ( .A(KEYINPUT10), .B(KEYINPUT0), .ZN(n1306) );
NAND2_X1 U1006 ( .A1(n1307), .A2(n1308), .ZN(n1292) );
OR2_X1 U1007 ( .A1(n1218), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1008 ( .A(n1310), .B(KEYINPUT1), .Z(n1307) );
NAND2_X1 U1009 ( .A1(n1309), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U1010 ( .A(KEYINPUT36), .B(n1218), .ZN(n1311) );
NAND2_X1 U1011 ( .A1(G224), .A2(n1275), .ZN(n1218) );
XOR2_X1 U1012 ( .A(n1156), .B(n1312), .Z(n1309) );
NOR2_X1 U1013 ( .A1(KEYINPUT42), .A2(n1219), .ZN(n1312) );
INV_X1 U1014 ( .A(n1044), .ZN(n1050) );
NAND3_X1 U1015 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1044) );
NAND2_X1 U1016 ( .A1(n1316), .A2(n1135), .ZN(n1315) );
OR3_X1 U1017 ( .A1(n1135), .A2(n1316), .A3(G902), .ZN(n1314) );
NOR2_X1 U1018 ( .A1(n1137), .A2(G234), .ZN(n1316) );
INV_X1 U1019 ( .A(G217), .ZN(n1137) );
XOR2_X1 U1020 ( .A(n1317), .B(G137), .Z(n1135) );
XOR2_X1 U1021 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1022 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1023 ( .A(KEYINPUT23), .B(G119), .Z(n1321) );
XOR2_X1 U1024 ( .A(KEYINPUT38), .B(KEYINPUT32), .Z(n1320) );
XOR2_X1 U1025 ( .A(n1322), .B(n1323), .Z(n1318) );
XOR2_X1 U1026 ( .A(G110), .B(n1324), .Z(n1323) );
NOR2_X1 U1027 ( .A1(n1255), .A2(n1325), .ZN(n1324) );
INV_X1 U1028 ( .A(G221), .ZN(n1325) );
NAND2_X1 U1029 ( .A1(G234), .A2(n1275), .ZN(n1255) );
XNOR2_X1 U1030 ( .A(n1326), .B(n1105), .ZN(n1322) );
XNOR2_X1 U1031 ( .A(G140), .B(n1219), .ZN(n1105) );
INV_X1 U1032 ( .A(G125), .ZN(n1219) );
NAND2_X1 U1033 ( .A1(G902), .A2(G217), .ZN(n1313) );
INV_X1 U1034 ( .A(n1184), .ZN(n1194) );
NOR2_X1 U1035 ( .A1(n1059), .A2(n1069), .ZN(n1184) );
INV_X1 U1036 ( .A(n1039), .ZN(n1069) );
NOR2_X1 U1037 ( .A1(n1086), .A2(n1327), .ZN(n1039) );
AND2_X1 U1038 ( .A1(n1328), .A2(n1087), .ZN(n1327) );
XOR2_X1 U1039 ( .A(KEYINPUT59), .B(G472), .Z(n1328) );
NOR2_X1 U1040 ( .A1(n1087), .A2(G472), .ZN(n1086) );
NAND2_X1 U1041 ( .A1(n1329), .A2(n1265), .ZN(n1087) );
XOR2_X1 U1042 ( .A(n1330), .B(n1149), .Z(n1329) );
XOR2_X1 U1043 ( .A(n1331), .B(n1332), .Z(n1149) );
XNOR2_X1 U1044 ( .A(n1303), .B(G101), .ZN(n1332) );
INV_X1 U1045 ( .A(G113), .ZN(n1303) );
XOR2_X1 U1046 ( .A(n1333), .B(n1301), .Z(n1331) );
XOR2_X1 U1047 ( .A(G116), .B(G119), .Z(n1301) );
NAND3_X1 U1048 ( .A1(n1275), .A2(n1274), .A3(G210), .ZN(n1333) );
INV_X1 U1049 ( .A(G237), .ZN(n1274) );
NAND2_X1 U1050 ( .A1(n1334), .A2(n1335), .ZN(n1330) );
NAND2_X1 U1051 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
INV_X1 U1052 ( .A(n1156), .ZN(n1337) );
XOR2_X1 U1053 ( .A(KEYINPUT15), .B(n1155), .Z(n1336) );
XOR2_X1 U1054 ( .A(n1338), .B(KEYINPUT61), .Z(n1334) );
NAND2_X1 U1055 ( .A1(n1339), .A2(n1156), .ZN(n1338) );
XOR2_X1 U1056 ( .A(n1340), .B(n1233), .Z(n1156) );
INV_X1 U1057 ( .A(G128), .ZN(n1233) );
NAND2_X1 U1058 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1059 ( .A1(KEYINPUT45), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1060 ( .A(G143), .B(n1277), .Z(n1343) );
NAND3_X1 U1061 ( .A1(G143), .A2(n1277), .A3(n1344), .ZN(n1341) );
INV_X1 U1062 ( .A(KEYINPUT45), .ZN(n1344) );
XNOR2_X1 U1063 ( .A(n1155), .B(KEYINPUT57), .ZN(n1339) );
NAND2_X1 U1064 ( .A1(n1247), .A2(n1083), .ZN(n1059) );
XNOR2_X1 U1065 ( .A(n1345), .B(G469), .ZN(n1083) );
NAND2_X1 U1066 ( .A1(n1346), .A2(n1265), .ZN(n1345) );
XOR2_X1 U1067 ( .A(n1347), .B(n1159), .Z(n1346) );
XOR2_X1 U1068 ( .A(n1348), .B(n1349), .Z(n1159) );
XNOR2_X1 U1069 ( .A(G140), .B(KEYINPUT41), .ZN(n1349) );
XNOR2_X1 U1070 ( .A(n1155), .B(n1350), .ZN(n1348) );
AND2_X1 U1071 ( .A1(n1275), .A2(G227), .ZN(n1350) );
XOR2_X1 U1072 ( .A(G953), .B(KEYINPUT12), .Z(n1275) );
XOR2_X1 U1073 ( .A(n1104), .B(KEYINPUT44), .Z(n1155) );
XOR2_X1 U1074 ( .A(G131), .B(n1351), .Z(n1104) );
XOR2_X1 U1075 ( .A(G137), .B(G134), .Z(n1351) );
XNOR2_X1 U1076 ( .A(n1164), .B(n1352), .ZN(n1347) );
NOR2_X1 U1077 ( .A1(G110), .A2(KEYINPUT5), .ZN(n1352) );
XNOR2_X1 U1078 ( .A(n1353), .B(n1304), .ZN(n1164) );
XOR2_X1 U1079 ( .A(G104), .B(n1354), .Z(n1304) );
XOR2_X1 U1080 ( .A(KEYINPUT18), .B(G107), .Z(n1354) );
XNOR2_X1 U1081 ( .A(n1106), .B(n1355), .ZN(n1353) );
NOR2_X1 U1082 ( .A1(G101), .A2(KEYINPUT14), .ZN(n1355) );
XNOR2_X1 U1083 ( .A(n1356), .B(n1326), .ZN(n1106) );
XNOR2_X1 U1084 ( .A(G128), .B(n1277), .ZN(n1326) );
XNOR2_X1 U1085 ( .A(G146), .B(KEYINPUT48), .ZN(n1277) );
XNOR2_X1 U1086 ( .A(G143), .B(KEYINPUT49), .ZN(n1356) );
XNOR2_X1 U1087 ( .A(KEYINPUT8), .B(n1062), .ZN(n1247) );
AND2_X1 U1088 ( .A1(G221), .A2(n1357), .ZN(n1062) );
NAND2_X1 U1089 ( .A1(G234), .A2(n1265), .ZN(n1357) );
INV_X1 U1090 ( .A(G902), .ZN(n1265) );
endmodule


