//Key = 1100101010101100001000110111101010100100111100111000000001000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
n1434, n1435, n1436;

XOR2_X1 U806 ( .A(G107), .B(n1094), .Z(G9) );
NOR2_X1 U807 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U808 ( .A1(n1097), .A2(n1098), .ZN(G75) );
NOR4_X1 U809 ( .A1(n1099), .A2(n1100), .A3(G953), .A4(n1101), .ZN(n1098) );
NOR2_X1 U810 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U811 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR2_X1 U812 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U813 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR3_X1 U814 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NOR2_X1 U815 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U816 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
AND3_X1 U817 ( .A1(n1117), .A2(n1115), .A3(n1116), .ZN(n1108) );
AND3_X1 U818 ( .A1(n1118), .A2(n1115), .A3(n1119), .ZN(n1104) );
NAND3_X1 U819 ( .A1(n1120), .A2(G952), .A3(n1121), .ZN(n1099) );
XOR2_X1 U820 ( .A(n1122), .B(KEYINPUT3), .Z(n1121) );
NAND3_X1 U821 ( .A1(n1116), .A2(n1123), .A3(n1124), .ZN(n1122) );
INV_X1 U822 ( .A(n1103), .ZN(n1124) );
NAND2_X1 U823 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND3_X1 U824 ( .A1(n1115), .A2(n1127), .A3(n1128), .ZN(n1126) );
NAND2_X1 U825 ( .A1(n1119), .A2(n1129), .ZN(n1125) );
NAND2_X1 U826 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U827 ( .A1(n1132), .A2(n1128), .ZN(n1131) );
NAND3_X1 U828 ( .A1(n1133), .A2(n1134), .A3(n1115), .ZN(n1130) );
OR2_X1 U829 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U830 ( .A1(n1135), .A2(n1137), .ZN(n1133) );
NAND2_X1 U831 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U832 ( .A1(n1140), .A2(KEYINPUT55), .ZN(n1135) );
NOR3_X1 U833 ( .A1(n1141), .A2(G953), .A3(n1101), .ZN(n1097) );
AND4_X1 U834 ( .A1(n1119), .A2(n1142), .A3(n1128), .A4(n1143), .ZN(n1101) );
NOR3_X1 U835 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1143) );
XNOR2_X1 U836 ( .A(G469), .B(n1147), .ZN(n1146) );
NAND2_X1 U837 ( .A1(KEYINPUT25), .A2(n1148), .ZN(n1147) );
XNOR2_X1 U838 ( .A(G472), .B(n1149), .ZN(n1145) );
XOR2_X1 U839 ( .A(KEYINPUT17), .B(n1150), .Z(n1144) );
NOR2_X1 U840 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
INV_X1 U841 ( .A(n1107), .ZN(n1128) );
NAND2_X1 U842 ( .A1(n1151), .A2(n1152), .ZN(n1142) );
XNOR2_X1 U843 ( .A(n1153), .B(KEYINPUT14), .ZN(n1152) );
XOR2_X1 U844 ( .A(KEYINPUT49), .B(G952), .Z(n1141) );
XOR2_X1 U845 ( .A(n1154), .B(n1155), .Z(G72) );
NOR2_X1 U846 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR2_X1 U847 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
INV_X1 U848 ( .A(n1160), .ZN(n1158) );
NOR3_X1 U849 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1156) );
XNOR2_X1 U850 ( .A(KEYINPUT50), .B(n1159), .ZN(n1162) );
NAND2_X1 U851 ( .A1(n1163), .A2(n1164), .ZN(n1159) );
NAND2_X1 U852 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U853 ( .A(KEYINPUT36), .B(n1167), .Z(n1166) );
NOR2_X1 U854 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U855 ( .A(KEYINPUT59), .B(n1170), .Z(n1169) );
INV_X1 U856 ( .A(n1171), .ZN(n1165) );
XNOR2_X1 U857 ( .A(n1172), .B(n1173), .ZN(n1160) );
XOR2_X1 U858 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U859 ( .A(n1176), .B(n1177), .ZN(n1172) );
NAND2_X1 U860 ( .A1(KEYINPUT0), .A2(n1178), .ZN(n1176) );
NAND2_X1 U861 ( .A1(G953), .A2(n1179), .ZN(n1154) );
NAND2_X1 U862 ( .A1(G227), .A2(n1180), .ZN(n1179) );
XOR2_X1 U863 ( .A(KEYINPUT58), .B(G900), .Z(n1180) );
XOR2_X1 U864 ( .A(n1181), .B(n1182), .Z(G69) );
XOR2_X1 U865 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U866 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XNOR2_X1 U867 ( .A(G953), .B(KEYINPUT12), .ZN(n1186) );
NOR2_X1 U868 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NAND2_X1 U869 ( .A1(n1189), .A2(n1190), .ZN(n1183) );
NAND2_X1 U870 ( .A1(G953), .A2(n1191), .ZN(n1190) );
XOR2_X1 U871 ( .A(n1192), .B(n1193), .Z(n1189) );
XNOR2_X1 U872 ( .A(n1194), .B(n1195), .ZN(n1193) );
NOR2_X1 U873 ( .A1(KEYINPUT38), .A2(n1196), .ZN(n1195) );
NAND2_X1 U874 ( .A1(KEYINPUT40), .A2(n1197), .ZN(n1194) );
NAND2_X1 U875 ( .A1(G953), .A2(n1198), .ZN(n1181) );
XOR2_X1 U876 ( .A(KEYINPUT18), .B(n1199), .Z(n1198) );
NOR2_X1 U877 ( .A1(n1200), .A2(n1191), .ZN(n1199) );
NOR2_X1 U878 ( .A1(n1201), .A2(n1202), .ZN(G66) );
NOR3_X1 U879 ( .A1(n1153), .A2(n1203), .A3(n1204), .ZN(n1202) );
AND3_X1 U880 ( .A1(n1205), .A2(n1151), .A3(n1206), .ZN(n1204) );
NOR2_X1 U881 ( .A1(n1207), .A2(n1205), .ZN(n1203) );
NOR2_X1 U882 ( .A1(n1120), .A2(n1208), .ZN(n1207) );
NOR2_X1 U883 ( .A1(n1201), .A2(n1209), .ZN(G63) );
XNOR2_X1 U884 ( .A(n1210), .B(n1211), .ZN(n1209) );
AND2_X1 U885 ( .A1(G478), .A2(n1206), .ZN(n1211) );
NOR2_X1 U886 ( .A1(n1201), .A2(n1212), .ZN(G60) );
XNOR2_X1 U887 ( .A(n1213), .B(n1214), .ZN(n1212) );
AND2_X1 U888 ( .A1(G475), .A2(n1206), .ZN(n1214) );
XNOR2_X1 U889 ( .A(G104), .B(n1215), .ZN(G6) );
NOR2_X1 U890 ( .A1(n1201), .A2(n1216), .ZN(G57) );
XOR2_X1 U891 ( .A(n1217), .B(n1218), .Z(n1216) );
XNOR2_X1 U892 ( .A(n1219), .B(n1220), .ZN(n1218) );
XOR2_X1 U893 ( .A(n1221), .B(KEYINPUT56), .Z(n1217) );
NAND2_X1 U894 ( .A1(n1206), .A2(G472), .ZN(n1221) );
NOR2_X1 U895 ( .A1(n1201), .A2(n1222), .ZN(G54) );
XOR2_X1 U896 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U897 ( .A(n1225), .B(n1226), .Z(n1224) );
NOR2_X1 U898 ( .A1(KEYINPUT52), .A2(n1227), .ZN(n1225) );
XOR2_X1 U899 ( .A(n1228), .B(n1229), .Z(n1223) );
NOR3_X1 U900 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1229) );
NOR2_X1 U901 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NOR3_X1 U902 ( .A1(G140), .A2(KEYINPUT15), .A3(n1235), .ZN(n1231) );
INV_X1 U903 ( .A(n1233), .ZN(n1235) );
NOR2_X1 U904 ( .A1(G110), .A2(KEYINPUT24), .ZN(n1233) );
AND2_X1 U905 ( .A1(G110), .A2(KEYINPUT15), .ZN(n1230) );
XOR2_X1 U906 ( .A(n1236), .B(n1237), .Z(n1228) );
NOR2_X1 U907 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NOR2_X1 U908 ( .A1(n1201), .A2(n1240), .ZN(G51) );
XNOR2_X1 U909 ( .A(n1241), .B(n1242), .ZN(n1240) );
XNOR2_X1 U910 ( .A(n1243), .B(n1244), .ZN(n1242) );
NOR4_X1 U911 ( .A1(n1245), .A2(n1246), .A3(KEYINPUT11), .A4(n1247), .ZN(n1244) );
INV_X1 U912 ( .A(G210), .ZN(n1247) );
NOR2_X1 U913 ( .A1(KEYINPUT30), .A2(n1248), .ZN(n1246) );
AND2_X1 U914 ( .A1(G902), .A2(n1120), .ZN(n1248) );
AND2_X1 U915 ( .A1(n1239), .A2(KEYINPUT30), .ZN(n1245) );
INV_X1 U916 ( .A(n1206), .ZN(n1239) );
NOR2_X1 U917 ( .A1(n1249), .A2(n1120), .ZN(n1206) );
NOR3_X1 U918 ( .A1(n1188), .A2(n1168), .A3(n1250), .ZN(n1120) );
OR3_X1 U919 ( .A1(n1171), .A2(n1170), .A3(n1251), .ZN(n1250) );
XNOR2_X1 U920 ( .A(n1187), .B(KEYINPUT23), .ZN(n1251) );
INV_X1 U921 ( .A(n1252), .ZN(n1187) );
AND4_X1 U922 ( .A1(n1253), .A2(n1119), .A3(n1254), .A4(n1255), .ZN(n1170) );
OR2_X1 U923 ( .A1(n1256), .A2(KEYINPUT33), .ZN(n1255) );
NAND2_X1 U924 ( .A1(KEYINPUT33), .A2(n1257), .ZN(n1254) );
NAND4_X1 U925 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1171) );
NAND2_X1 U926 ( .A1(n1262), .A2(n1256), .ZN(n1259) );
NAND2_X1 U927 ( .A1(n1263), .A2(n1264), .ZN(n1168) );
NAND2_X1 U928 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U929 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND3_X1 U930 ( .A1(n1269), .A2(n1270), .A3(n1113), .ZN(n1268) );
NAND2_X1 U931 ( .A1(n1117), .A2(n1253), .ZN(n1267) );
NAND4_X1 U932 ( .A1(n1271), .A2(n1215), .A3(n1272), .A4(n1273), .ZN(n1188) );
AND4_X1 U933 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1273) );
NAND2_X1 U934 ( .A1(n1278), .A2(n1279), .ZN(n1272) );
XOR2_X1 U935 ( .A(n1095), .B(KEYINPUT4), .Z(n1278) );
NAND3_X1 U936 ( .A1(n1115), .A2(n1127), .A3(n1280), .ZN(n1095) );
AND3_X1 U937 ( .A1(n1114), .A2(n1281), .A3(n1282), .ZN(n1280) );
NAND3_X1 U938 ( .A1(n1283), .A2(n1115), .A3(n1117), .ZN(n1215) );
NAND3_X1 U939 ( .A1(n1119), .A2(n1284), .A3(n1285), .ZN(n1271) );
XNOR2_X1 U940 ( .A(KEYINPUT53), .B(n1286), .ZN(n1284) );
NOR2_X1 U941 ( .A1(n1163), .A2(G952), .ZN(n1201) );
XNOR2_X1 U942 ( .A(G146), .B(n1287), .ZN(G48) );
NAND4_X1 U943 ( .A1(KEYINPUT63), .A2(n1265), .A3(n1117), .A4(n1253), .ZN(n1287) );
XNOR2_X1 U944 ( .A(G143), .B(n1288), .ZN(G45) );
NAND3_X1 U945 ( .A1(KEYINPUT22), .A2(n1265), .A3(n1289), .ZN(n1288) );
AND3_X1 U946 ( .A1(n1113), .A2(n1270), .A3(n1269), .ZN(n1289) );
XNOR2_X1 U947 ( .A(G140), .B(n1263), .ZN(G42) );
NAND2_X1 U948 ( .A1(n1256), .A2(n1290), .ZN(n1263) );
XOR2_X1 U949 ( .A(G137), .B(n1291), .Z(G39) );
NOR4_X1 U950 ( .A1(KEYINPUT7), .A2(n1110), .A3(n1286), .A4(n1292), .ZN(n1291) );
XNOR2_X1 U951 ( .A(G134), .B(n1293), .ZN(G36) );
NAND3_X1 U952 ( .A1(n1294), .A2(n1295), .A3(n1262), .ZN(n1293) );
OR2_X1 U953 ( .A1(n1256), .A2(KEYINPUT51), .ZN(n1295) );
NAND2_X1 U954 ( .A1(KEYINPUT51), .A2(n1257), .ZN(n1294) );
NAND2_X1 U955 ( .A1(n1296), .A2(n1297), .ZN(n1257) );
INV_X1 U956 ( .A(n1298), .ZN(n1296) );
XNOR2_X1 U957 ( .A(G131), .B(n1260), .ZN(G33) );
NAND3_X1 U958 ( .A1(n1113), .A2(n1117), .A3(n1256), .ZN(n1260) );
INV_X1 U959 ( .A(n1292), .ZN(n1256) );
NAND2_X1 U960 ( .A1(n1297), .A2(n1298), .ZN(n1292) );
NOR2_X1 U961 ( .A1(n1107), .A2(n1116), .ZN(n1297) );
NAND2_X1 U962 ( .A1(n1136), .A2(n1281), .ZN(n1107) );
AND2_X1 U963 ( .A1(n1139), .A2(n1299), .ZN(n1136) );
NAND3_X1 U964 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(G30) );
NAND2_X1 U965 ( .A1(n1261), .A2(n1303), .ZN(n1302) );
OR3_X1 U966 ( .A1(n1303), .A2(n1261), .A3(G128), .ZN(n1301) );
INV_X1 U967 ( .A(KEYINPUT13), .ZN(n1303) );
NAND2_X1 U968 ( .A1(G128), .A2(n1304), .ZN(n1300) );
NAND2_X1 U969 ( .A1(KEYINPUT13), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U970 ( .A(KEYINPUT16), .B(n1261), .ZN(n1305) );
NAND3_X1 U971 ( .A1(n1253), .A2(n1127), .A3(n1265), .ZN(n1261) );
AND2_X1 U972 ( .A1(n1306), .A2(n1298), .ZN(n1265) );
XNOR2_X1 U973 ( .A(G101), .B(n1277), .ZN(G3) );
NAND3_X1 U974 ( .A1(n1283), .A2(n1119), .A3(n1113), .ZN(n1277) );
XNOR2_X1 U975 ( .A(G125), .B(n1307), .ZN(G27) );
NOR2_X1 U976 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NOR2_X1 U977 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND4_X1 U978 ( .A1(n1118), .A2(n1132), .A3(n1312), .A4(n1298), .ZN(n1311) );
INV_X1 U979 ( .A(KEYINPUT20), .ZN(n1310) );
NOR2_X1 U980 ( .A1(KEYINPUT20), .A2(n1258), .ZN(n1308) );
NAND3_X1 U981 ( .A1(n1118), .A2(n1298), .A3(n1290), .ZN(n1258) );
AND2_X1 U982 ( .A1(n1117), .A2(n1132), .ZN(n1290) );
NAND2_X1 U983 ( .A1(n1103), .A2(n1313), .ZN(n1298) );
NAND3_X1 U984 ( .A1(G902), .A2(n1314), .A3(n1161), .ZN(n1313) );
NOR2_X1 U985 ( .A1(n1163), .A2(G900), .ZN(n1161) );
XNOR2_X1 U986 ( .A(G122), .B(n1276), .ZN(G24) );
NAND4_X1 U987 ( .A1(n1269), .A2(n1285), .A3(n1115), .A4(n1270), .ZN(n1276) );
NOR2_X1 U988 ( .A1(n1315), .A2(n1316), .ZN(n1115) );
XNOR2_X1 U989 ( .A(G119), .B(n1317), .ZN(G21) );
NAND4_X1 U990 ( .A1(n1318), .A2(n1118), .A3(n1253), .A4(n1119), .ZN(n1317) );
INV_X1 U991 ( .A(n1286), .ZN(n1253) );
NAND2_X1 U992 ( .A1(n1316), .A2(n1315), .ZN(n1286) );
INV_X1 U993 ( .A(n1319), .ZN(n1315) );
XOR2_X1 U994 ( .A(n1282), .B(KEYINPUT5), .Z(n1318) );
XNOR2_X1 U995 ( .A(G116), .B(n1252), .ZN(G18) );
NAND2_X1 U996 ( .A1(n1262), .A2(n1285), .ZN(n1252) );
AND2_X1 U997 ( .A1(n1113), .A2(n1127), .ZN(n1262) );
AND2_X1 U998 ( .A1(n1320), .A2(n1270), .ZN(n1127) );
XNOR2_X1 U999 ( .A(G113), .B(n1275), .ZN(G15) );
NAND3_X1 U1000 ( .A1(n1285), .A2(n1117), .A3(n1113), .ZN(n1275) );
NOR2_X1 U1001 ( .A1(n1319), .A2(n1316), .ZN(n1113) );
INV_X1 U1002 ( .A(n1312), .ZN(n1117) );
NAND2_X1 U1003 ( .A1(n1269), .A2(n1321), .ZN(n1312) );
XOR2_X1 U1004 ( .A(n1320), .B(KEYINPUT26), .Z(n1269) );
AND2_X1 U1005 ( .A1(n1118), .A2(n1282), .ZN(n1285) );
NOR3_X1 U1006 ( .A1(n1096), .A2(n1140), .A3(n1114), .ZN(n1118) );
INV_X1 U1007 ( .A(n1116), .ZN(n1114) );
NAND3_X1 U1008 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(G12) );
NAND2_X1 U1009 ( .A1(G110), .A2(n1274), .ZN(n1324) );
NAND2_X1 U1010 ( .A1(KEYINPUT60), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1011 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
XNOR2_X1 U1012 ( .A(KEYINPUT2), .B(n1274), .ZN(n1326) );
NAND2_X1 U1013 ( .A1(n1328), .A2(n1329), .ZN(n1322) );
INV_X1 U1014 ( .A(KEYINPUT60), .ZN(n1329) );
NAND2_X1 U1015 ( .A1(n1330), .A2(n1331), .ZN(n1328) );
NAND2_X1 U1016 ( .A1(KEYINPUT2), .A2(n1274), .ZN(n1331) );
OR3_X1 U1017 ( .A1(G110), .A2(KEYINPUT2), .A3(n1274), .ZN(n1330) );
NAND3_X1 U1018 ( .A1(n1132), .A2(n1119), .A3(n1283), .ZN(n1274) );
AND2_X1 U1019 ( .A1(n1306), .A2(n1282), .ZN(n1283) );
NAND2_X1 U1020 ( .A1(n1103), .A2(n1332), .ZN(n1282) );
NAND4_X1 U1021 ( .A1(G953), .A2(G902), .A3(n1314), .A4(n1191), .ZN(n1332) );
INV_X1 U1022 ( .A(G898), .ZN(n1191) );
NAND3_X1 U1023 ( .A1(n1314), .A2(n1163), .A3(G952), .ZN(n1103) );
NAND2_X1 U1024 ( .A1(G234), .A2(G237), .ZN(n1314) );
NOR3_X1 U1025 ( .A1(n1116), .A2(n1140), .A3(n1096), .ZN(n1306) );
INV_X1 U1026 ( .A(n1279), .ZN(n1096) );
NOR2_X1 U1027 ( .A1(n1139), .A2(n1138), .ZN(n1279) );
INV_X1 U1028 ( .A(n1299), .ZN(n1138) );
NAND2_X1 U1029 ( .A1(G214), .A2(n1333), .ZN(n1299) );
XOR2_X1 U1030 ( .A(n1334), .B(n1335), .Z(n1139) );
AND2_X1 U1031 ( .A1(n1333), .A2(G210), .ZN(n1335) );
NAND2_X1 U1032 ( .A1(n1336), .A2(n1249), .ZN(n1333) );
XNOR2_X1 U1033 ( .A(G237), .B(KEYINPUT31), .ZN(n1336) );
NAND3_X1 U1034 ( .A1(n1337), .A2(n1338), .A3(n1249), .ZN(n1334) );
NAND2_X1 U1035 ( .A1(G125), .A2(n1241), .ZN(n1338) );
NAND2_X1 U1036 ( .A1(n1339), .A2(n1243), .ZN(n1337) );
XNOR2_X1 U1037 ( .A(KEYINPUT28), .B(n1340), .ZN(n1339) );
INV_X1 U1038 ( .A(n1241), .ZN(n1340) );
XNOR2_X1 U1039 ( .A(n1341), .B(n1342), .ZN(n1241) );
XOR2_X1 U1040 ( .A(n1197), .B(n1196), .Z(n1342) );
NAND2_X1 U1041 ( .A1(n1343), .A2(n1344), .ZN(n1196) );
NAND2_X1 U1042 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1043 ( .A1(n1347), .A2(G116), .ZN(n1343) );
XOR2_X1 U1044 ( .A(n1345), .B(KEYINPUT61), .Z(n1347) );
XNOR2_X1 U1045 ( .A(G113), .B(G119), .ZN(n1345) );
XNOR2_X1 U1046 ( .A(G122), .B(G110), .ZN(n1197) );
XOR2_X1 U1047 ( .A(n1348), .B(n1349), .Z(n1341) );
XOR2_X1 U1048 ( .A(n1350), .B(n1351), .Z(n1348) );
NOR2_X1 U1049 ( .A1(G953), .A2(n1200), .ZN(n1351) );
INV_X1 U1050 ( .A(G224), .ZN(n1200) );
NAND2_X1 U1051 ( .A1(KEYINPUT37), .A2(n1192), .ZN(n1350) );
INV_X1 U1052 ( .A(n1281), .ZN(n1140) );
NAND2_X1 U1053 ( .A1(G221), .A2(n1352), .ZN(n1281) );
XOR2_X1 U1054 ( .A(n1148), .B(n1238), .Z(n1116) );
INV_X1 U1055 ( .A(G469), .ZN(n1238) );
AND2_X1 U1056 ( .A1(n1353), .A2(n1249), .ZN(n1148) );
XOR2_X1 U1057 ( .A(n1227), .B(n1354), .Z(n1353) );
XNOR2_X1 U1058 ( .A(n1355), .B(n1226), .ZN(n1354) );
XOR2_X1 U1059 ( .A(G131), .B(n1356), .Z(n1226) );
NAND2_X1 U1060 ( .A1(n1357), .A2(n1358), .ZN(n1355) );
NAND2_X1 U1061 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
XOR2_X1 U1062 ( .A(n1361), .B(KEYINPUT62), .Z(n1357) );
OR2_X1 U1063 ( .A1(n1360), .A2(n1359), .ZN(n1361) );
XOR2_X1 U1064 ( .A(n1362), .B(G140), .Z(n1359) );
NAND2_X1 U1065 ( .A1(KEYINPUT27), .A2(n1327), .ZN(n1362) );
XNOR2_X1 U1066 ( .A(n1236), .B(KEYINPUT41), .ZN(n1360) );
NAND2_X1 U1067 ( .A1(G227), .A2(n1163), .ZN(n1236) );
XOR2_X1 U1068 ( .A(n1178), .B(n1192), .Z(n1227) );
XOR2_X1 U1069 ( .A(n1363), .B(n1364), .Z(n1192) );
XOR2_X1 U1070 ( .A(KEYINPUT6), .B(G107), .Z(n1364) );
XNOR2_X1 U1071 ( .A(G101), .B(G104), .ZN(n1363) );
AND2_X1 U1072 ( .A1(n1365), .A2(n1366), .ZN(n1178) );
NAND2_X1 U1073 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
XOR2_X1 U1074 ( .A(KEYINPUT46), .B(n1369), .Z(n1365) );
NOR2_X1 U1075 ( .A1(n1370), .A2(n1368), .ZN(n1369) );
XNOR2_X1 U1076 ( .A(KEYINPUT47), .B(n1367), .ZN(n1370) );
NAND2_X1 U1077 ( .A1(n1371), .A2(n1372), .ZN(n1367) );
NAND2_X1 U1078 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XNOR2_X1 U1079 ( .A(G143), .B(KEYINPUT44), .ZN(n1373) );
NAND2_X1 U1080 ( .A1(G146), .A2(n1375), .ZN(n1371) );
XNOR2_X1 U1081 ( .A(G143), .B(KEYINPUT42), .ZN(n1375) );
INV_X1 U1082 ( .A(n1110), .ZN(n1119) );
NAND2_X1 U1083 ( .A1(n1321), .A2(n1320), .ZN(n1110) );
XOR2_X1 U1084 ( .A(n1376), .B(G475), .Z(n1320) );
NAND2_X1 U1085 ( .A1(n1213), .A2(n1249), .ZN(n1376) );
XNOR2_X1 U1086 ( .A(n1377), .B(n1378), .ZN(n1213) );
XOR2_X1 U1087 ( .A(n1379), .B(n1380), .Z(n1378) );
XOR2_X1 U1088 ( .A(n1381), .B(n1382), .Z(n1380) );
AND3_X1 U1089 ( .A1(G214), .A2(n1163), .A3(n1383), .ZN(n1382) );
NAND2_X1 U1090 ( .A1(KEYINPUT57), .A2(n1384), .ZN(n1381) );
INV_X1 U1091 ( .A(G104), .ZN(n1384) );
XNOR2_X1 U1092 ( .A(G122), .B(KEYINPUT34), .ZN(n1379) );
XNOR2_X1 U1093 ( .A(n1175), .B(n1385), .ZN(n1377) );
XOR2_X1 U1094 ( .A(n1386), .B(n1387), .Z(n1385) );
XNOR2_X1 U1095 ( .A(G125), .B(n1234), .ZN(n1175) );
INV_X1 U1096 ( .A(n1270), .ZN(n1321) );
XNOR2_X1 U1097 ( .A(n1388), .B(G478), .ZN(n1270) );
NAND2_X1 U1098 ( .A1(n1249), .A2(n1210), .ZN(n1388) );
NAND2_X1 U1099 ( .A1(n1389), .A2(n1390), .ZN(n1210) );
NAND4_X1 U1100 ( .A1(n1391), .A2(G217), .A3(G234), .A4(n1392), .ZN(n1390) );
XOR2_X1 U1101 ( .A(n1393), .B(KEYINPUT9), .Z(n1389) );
NAND2_X1 U1102 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
NAND3_X1 U1103 ( .A1(G217), .A2(G234), .A3(n1391), .ZN(n1395) );
XNOR2_X1 U1104 ( .A(G953), .B(KEYINPUT35), .ZN(n1391) );
INV_X1 U1105 ( .A(n1392), .ZN(n1394) );
XNOR2_X1 U1106 ( .A(n1396), .B(n1397), .ZN(n1392) );
XNOR2_X1 U1107 ( .A(G107), .B(n1398), .ZN(n1397) );
NAND2_X1 U1108 ( .A1(n1399), .A2(KEYINPUT43), .ZN(n1398) );
XNOR2_X1 U1109 ( .A(G128), .B(n1400), .ZN(n1399) );
XOR2_X1 U1110 ( .A(G143), .B(G134), .Z(n1400) );
XNOR2_X1 U1111 ( .A(G122), .B(G116), .ZN(n1396) );
AND2_X1 U1112 ( .A1(n1316), .A2(n1319), .ZN(n1132) );
NAND2_X1 U1113 ( .A1(n1401), .A2(n1402), .ZN(n1319) );
NAND2_X1 U1114 ( .A1(KEYINPUT48), .A2(n1403), .ZN(n1402) );
XOR2_X1 U1115 ( .A(n1149), .B(G472), .Z(n1403) );
NAND3_X1 U1116 ( .A1(G472), .A2(n1149), .A3(n1404), .ZN(n1401) );
INV_X1 U1117 ( .A(KEYINPUT48), .ZN(n1404) );
NAND2_X1 U1118 ( .A1(n1405), .A2(n1249), .ZN(n1149) );
XNOR2_X1 U1119 ( .A(n1406), .B(n1407), .ZN(n1405) );
INV_X1 U1120 ( .A(n1219), .ZN(n1407) );
XNOR2_X1 U1121 ( .A(n1408), .B(G101), .ZN(n1219) );
NAND3_X1 U1122 ( .A1(n1383), .A2(n1163), .A3(G210), .ZN(n1408) );
INV_X1 U1123 ( .A(G237), .ZN(n1383) );
NAND2_X1 U1124 ( .A1(KEYINPUT10), .A2(n1220), .ZN(n1406) );
XOR2_X1 U1125 ( .A(n1409), .B(n1410), .Z(n1220) );
XOR2_X1 U1126 ( .A(n1411), .B(n1356), .Z(n1410) );
XNOR2_X1 U1127 ( .A(n1412), .B(KEYINPUT32), .ZN(n1356) );
NAND3_X1 U1128 ( .A1(n1413), .A2(n1414), .A3(KEYINPUT8), .ZN(n1412) );
OR2_X1 U1129 ( .A1(n1174), .A2(KEYINPUT19), .ZN(n1414) );
XOR2_X1 U1130 ( .A(G134), .B(G137), .Z(n1174) );
NAND3_X1 U1131 ( .A1(G134), .A2(n1415), .A3(KEYINPUT19), .ZN(n1413) );
INV_X1 U1132 ( .A(G137), .ZN(n1415) );
NOR2_X1 U1133 ( .A1(n1416), .A2(n1417), .ZN(n1411) );
XOR2_X1 U1134 ( .A(KEYINPUT21), .B(n1418), .Z(n1417) );
NOR2_X1 U1135 ( .A1(G116), .A2(n1419), .ZN(n1418) );
NOR2_X1 U1136 ( .A1(G119), .A2(n1346), .ZN(n1416) );
INV_X1 U1137 ( .A(G116), .ZN(n1346) );
XNOR2_X1 U1138 ( .A(n1349), .B(n1387), .ZN(n1409) );
XNOR2_X1 U1139 ( .A(G113), .B(n1177), .ZN(n1387) );
INV_X1 U1140 ( .A(G131), .ZN(n1177) );
XOR2_X1 U1141 ( .A(G128), .B(n1386), .Z(n1349) );
XNOR2_X1 U1142 ( .A(G143), .B(n1374), .ZN(n1386) );
XNOR2_X1 U1143 ( .A(n1153), .B(n1420), .ZN(n1316) );
NOR2_X1 U1144 ( .A1(n1151), .A2(KEYINPUT39), .ZN(n1420) );
INV_X1 U1145 ( .A(n1208), .ZN(n1151) );
NAND2_X1 U1146 ( .A1(G217), .A2(n1352), .ZN(n1208) );
NAND2_X1 U1147 ( .A1(G234), .A2(n1249), .ZN(n1352) );
INV_X1 U1148 ( .A(G902), .ZN(n1249) );
NOR2_X1 U1149 ( .A1(n1205), .A2(G902), .ZN(n1153) );
XOR2_X1 U1150 ( .A(n1421), .B(n1422), .Z(n1205) );
XNOR2_X1 U1151 ( .A(n1243), .B(n1423), .ZN(n1422) );
XNOR2_X1 U1152 ( .A(n1374), .B(G137), .ZN(n1423) );
INV_X1 U1153 ( .A(G146), .ZN(n1374) );
INV_X1 U1154 ( .A(G125), .ZN(n1243) );
XOR2_X1 U1155 ( .A(n1424), .B(n1425), .Z(n1421) );
XOR2_X1 U1156 ( .A(n1426), .B(n1427), .Z(n1425) );
NAND2_X1 U1157 ( .A1(KEYINPUT1), .A2(n1234), .ZN(n1427) );
INV_X1 U1158 ( .A(G140), .ZN(n1234) );
NAND3_X1 U1159 ( .A1(n1428), .A2(n1429), .A3(n1430), .ZN(n1426) );
NAND2_X1 U1160 ( .A1(KEYINPUT54), .A2(n1431), .ZN(n1430) );
NAND3_X1 U1161 ( .A1(n1432), .A2(n1433), .A3(n1327), .ZN(n1429) );
INV_X1 U1162 ( .A(KEYINPUT54), .ZN(n1433) );
OR2_X1 U1163 ( .A1(n1327), .A2(n1432), .ZN(n1428) );
NOR2_X1 U1164 ( .A1(n1431), .A2(KEYINPUT29), .ZN(n1432) );
AND2_X1 U1165 ( .A1(n1434), .A2(n1435), .ZN(n1431) );
NAND2_X1 U1166 ( .A1(G128), .A2(n1419), .ZN(n1435) );
INV_X1 U1167 ( .A(G119), .ZN(n1419) );
XOR2_X1 U1168 ( .A(n1436), .B(KEYINPUT45), .Z(n1434) );
NAND2_X1 U1169 ( .A1(G119), .A2(n1368), .ZN(n1436) );
INV_X1 U1170 ( .A(G128), .ZN(n1368) );
INV_X1 U1171 ( .A(G110), .ZN(n1327) );
NAND3_X1 U1172 ( .A1(G234), .A2(n1163), .A3(G221), .ZN(n1424) );
INV_X1 U1173 ( .A(G953), .ZN(n1163) );
endmodule


