//Key = 0100110011011010111101101111110001110011011000011001100101111110


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
n2308, n2309, n2310;

OR2_X1 U1295 ( .A1(n2310), .A2(n1739), .ZN(U280) );
OR2_X1 U1296 ( .A1(n1878), .A2(STATO_REG_0__SCAN_IN), .ZN(n1738) );
INV_X2 U1297 ( .A(n1738), .ZN(n1739) );
INV_X2 U1298 ( .A(U280), .ZN(n1740) );
XOR2_X1 U1299 ( .A(n1741), .B(KEYINPUT55), .Z(U375) );
NAND2_X1 U1300 ( .A1(n1742), .A2(n1743), .ZN(U344) );
NAND2_X1 U1301 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1744), .ZN(n1743) );
NAND2_X1 U1302 ( .A1(n1745), .A2(DATA_IN_7_), .ZN(n1742) );
NAND2_X1 U1303 ( .A1(n1746), .A2(n1747), .ZN(U343) );
NAND2_X1 U1304 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1744), .ZN(n1747) );
NAND2_X1 U1305 ( .A1(n1745), .A2(DATA_IN_6_), .ZN(n1746) );
NAND2_X1 U1306 ( .A1(n1748), .A2(n1749), .ZN(U342) );
NAND2_X1 U1307 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1744), .ZN(n1749) );
NAND2_X1 U1308 ( .A1(n1745), .A2(DATA_IN_5_), .ZN(n1748) );
NAND2_X1 U1309 ( .A1(n1750), .A2(n1751), .ZN(U341) );
NAND2_X1 U1310 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1744), .ZN(n1751) );
NAND2_X1 U1311 ( .A1(n1745), .A2(DATA_IN_4_), .ZN(n1750) );
NAND2_X1 U1312 ( .A1(n1752), .A2(n1753), .ZN(U340) );
NAND2_X1 U1313 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1744), .ZN(n1753) );
NAND2_X1 U1314 ( .A1(n1745), .A2(DATA_IN_3_), .ZN(n1752) );
NAND2_X1 U1315 ( .A1(n1754), .A2(n1755), .ZN(U339) );
NAND2_X1 U1316 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1744), .ZN(n1755) );
NAND2_X1 U1317 ( .A1(n1745), .A2(DATA_IN_2_), .ZN(n1754) );
NAND2_X1 U1318 ( .A1(n1756), .A2(n1757), .ZN(U338) );
NAND2_X1 U1319 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1744), .ZN(n1757) );
NAND2_X1 U1320 ( .A1(n1745), .A2(DATA_IN_1_), .ZN(n1756) );
NAND2_X1 U1321 ( .A1(n1758), .A2(n1759), .ZN(U337) );
NAND2_X1 U1322 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1744), .ZN(n1759) );
NAND2_X1 U1323 ( .A1(n1745), .A2(n1760), .ZN(n1758) );
XNOR2_X1 U1324 ( .A(DATA_IN_0_), .B(KEYINPUT57), .ZN(n1760) );
INV_X1 U1325 ( .A(n1744), .ZN(n1745) );
NAND2_X1 U1326 ( .A1(n1741), .A2(n1761), .ZN(n1744) );
NAND3_X1 U1327 ( .A1(n1762), .A2(n1763), .A3(n1764), .ZN(n1761) );
NAND2_X1 U1328 ( .A1(n1765), .A2(n1766), .ZN(U336) );
NAND2_X1 U1329 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1767), .ZN(n1766) );
NAND2_X1 U1330 ( .A1(n1768), .A2(DATA_IN_7_), .ZN(n1765) );
NAND2_X1 U1331 ( .A1(n1769), .A2(n1770), .ZN(U335) );
NAND2_X1 U1332 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1767), .ZN(n1770) );
NAND2_X1 U1333 ( .A1(n1768), .A2(DATA_IN_6_), .ZN(n1769) );
NAND2_X1 U1334 ( .A1(n1771), .A2(n1772), .ZN(U334) );
NAND2_X1 U1335 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1767), .ZN(n1772) );
NAND2_X1 U1336 ( .A1(n1768), .A2(DATA_IN_5_), .ZN(n1771) );
NAND2_X1 U1337 ( .A1(n1773), .A2(n1774), .ZN(U333) );
NAND2_X1 U1338 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1767), .ZN(n1774) );
NAND2_X1 U1339 ( .A1(n1768), .A2(DATA_IN_4_), .ZN(n1773) );
NAND2_X1 U1340 ( .A1(n1775), .A2(n1776), .ZN(U332) );
NAND2_X1 U1341 ( .A1(DATA_IN_3_), .A2(n1777), .ZN(n1776) );
XNOR2_X1 U1342 ( .A(KEYINPUT46), .B(n1767), .ZN(n1777) );
NAND2_X1 U1343 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1767), .ZN(n1775) );
NAND2_X1 U1344 ( .A1(n1778), .A2(n1779), .ZN(U331) );
NAND2_X1 U1345 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1767), .ZN(n1779) );
NAND2_X1 U1346 ( .A1(n1768), .A2(DATA_IN_2_), .ZN(n1778) );
NAND2_X1 U1347 ( .A1(n1780), .A2(n1781), .ZN(U330) );
NAND2_X1 U1348 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1782), .ZN(n1781) );
XNOR2_X1 U1349 ( .A(KEYINPUT22), .B(n1767), .ZN(n1782) );
NAND2_X1 U1350 ( .A1(n1768), .A2(DATA_IN_1_), .ZN(n1780) );
NAND2_X1 U1351 ( .A1(n1783), .A2(n1784), .ZN(U329) );
NAND2_X1 U1352 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1767), .ZN(n1784) );
NAND2_X1 U1353 ( .A1(n1768), .A2(DATA_IN_0_), .ZN(n1783) );
INV_X1 U1354 ( .A(n1767), .ZN(n1768) );
NAND2_X1 U1355 ( .A1(n1741), .A2(n1785), .ZN(n1767) );
NAND2_X1 U1356 ( .A1(n1786), .A2(n1763), .ZN(n1785) );
NAND3_X1 U1357 ( .A1(n1764), .A2(n1762), .A3(n1787), .ZN(n1786) );
NAND2_X1 U1358 ( .A1(n1788), .A2(n1789), .ZN(n1787) );
NAND3_X1 U1359 ( .A1(n1790), .A2(n1791), .A3(n1792), .ZN(n1789) );
NAND2_X1 U1360 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1793), .ZN(n1792) );
NAND3_X1 U1361 ( .A1(n1794), .A2(n1795), .A3(n1796), .ZN(n1791) );
NAND2_X1 U1362 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1797), .ZN(n1796) );
NAND3_X1 U1363 ( .A1(n1798), .A2(n1799), .A3(n1800), .ZN(n1795) );
NAND2_X1 U1364 ( .A1(DATA_IN_5_), .A2(n1801), .ZN(n1800) );
NAND3_X1 U1365 ( .A1(n1802), .A2(n1803), .A3(n1804), .ZN(n1799) );
NAND2_X1 U1366 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1805), .ZN(n1804) );
NAND3_X1 U1367 ( .A1(n1806), .A2(n1807), .A3(n1808), .ZN(n1803) );
NAND2_X1 U1368 ( .A1(DATA_IN_3_), .A2(n1809), .ZN(n1808) );
NAND3_X1 U1369 ( .A1(n1810), .A2(n1811), .A3(n1812), .ZN(n1807) );
NAND2_X1 U1370 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1813), .ZN(n1812) );
NAND3_X1 U1371 ( .A1(n1814), .A2(n1815), .A3(n1816), .ZN(n1811) );
XNOR2_X1 U1372 ( .A(KEYINPUT25), .B(n1817), .ZN(n1816) );
NAND2_X1 U1373 ( .A1(DATA_IN_1_), .A2(n1818), .ZN(n1815) );
XOR2_X1 U1374 ( .A(RMIN_REG_0__SCAN_IN), .B(KEYINPUT31), .Z(n1814) );
NAND2_X1 U1375 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1819), .ZN(n1810) );
NAND2_X1 U1376 ( .A1(DATA_IN_2_), .A2(n1820), .ZN(n1806) );
NAND2_X1 U1377 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1821), .ZN(n1802) );
XNOR2_X1 U1378 ( .A(DATA_IN_3_), .B(n1822), .ZN(n1821) );
XNOR2_X1 U1379 ( .A(KEYINPUT40), .B(KEYINPUT35), .ZN(n1822) );
NAND2_X1 U1380 ( .A1(DATA_IN_4_), .A2(n1823), .ZN(n1798) );
NAND2_X1 U1381 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1824), .ZN(n1794) );
NAND2_X1 U1382 ( .A1(DATA_IN_6_), .A2(n1825), .ZN(n1790) );
XNOR2_X1 U1383 ( .A(n1826), .B(KEYINPUT16), .ZN(n1825) );
NAND2_X1 U1384 ( .A1(DATA_IN_7_), .A2(n1827), .ZN(n1788) );
NAND3_X1 U1385 ( .A1(n1828), .A2(n1829), .A3(n1830), .ZN(n1762) );
NAND2_X1 U1386 ( .A1(DATA_IN_7_), .A2(n1831), .ZN(n1830) );
NAND3_X1 U1387 ( .A1(n1832), .A2(n1833), .A3(n1834), .ZN(n1829) );
NAND2_X1 U1388 ( .A1(DATA_IN_6_), .A2(n1835), .ZN(n1834) );
NAND3_X1 U1389 ( .A1(n1836), .A2(n1837), .A3(n1838), .ZN(n1833) );
NAND2_X1 U1390 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1824), .ZN(n1838) );
NAND3_X1 U1391 ( .A1(n1839), .A2(n1840), .A3(n1841), .ZN(n1837) );
XOR2_X1 U1392 ( .A(KEYINPUT5), .B(n1842), .Z(n1841) );
NOR2_X1 U1393 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1843), .ZN(n1842) );
XNOR2_X1 U1394 ( .A(DATA_IN_4_), .B(KEYINPUT6), .ZN(n1843) );
NAND3_X1 U1395 ( .A1(n1844), .A2(n1845), .A3(n1846), .ZN(n1840) );
NAND2_X1 U1396 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1847), .ZN(n1846) );
NAND3_X1 U1397 ( .A1(n1848), .A2(n1849), .A3(n1850), .ZN(n1845) );
NAND2_X1 U1398 ( .A1(DATA_IN_2_), .A2(n1851), .ZN(n1850) );
NAND3_X1 U1399 ( .A1(DATA_IN_0_), .A2(n1852), .A3(n1853), .ZN(n1849) );
XNOR2_X1 U1400 ( .A(RMAX_REG_0__SCAN_IN), .B(KEYINPUT53), .ZN(n1853) );
NAND2_X1 U1401 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1819), .ZN(n1852) );
NAND2_X1 U1402 ( .A1(DATA_IN_1_), .A2(n1854), .ZN(n1848) );
XNOR2_X1 U1403 ( .A(n1855), .B(KEYINPUT38), .ZN(n1854) );
NAND2_X1 U1404 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1813), .ZN(n1844) );
NAND2_X1 U1405 ( .A1(DATA_IN_3_), .A2(n1856), .ZN(n1839) );
NAND2_X1 U1406 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1805), .ZN(n1836) );
INV_X1 U1407 ( .A(DATA_IN_4_), .ZN(n1805) );
NAND2_X1 U1408 ( .A1(DATA_IN_5_), .A2(n1857), .ZN(n1832) );
NAND2_X1 U1409 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1797), .ZN(n1828) );
INV_X1 U1410 ( .A(DATA_IN_6_), .ZN(n1797) );
NAND2_X1 U1411 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1793), .ZN(n1764) );
INV_X1 U1412 ( .A(DATA_IN_7_), .ZN(n1793) );
NAND2_X1 U1413 ( .A1(n1858), .A2(n1859), .ZN(U328) );
NAND2_X1 U1414 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1860), .ZN(n1859) );
NAND2_X1 U1415 ( .A1(n1861), .A2(DATA_IN_7_), .ZN(n1858) );
NAND2_X1 U1416 ( .A1(n1862), .A2(n1863), .ZN(U327) );
NAND2_X1 U1417 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1860), .ZN(n1863) );
NAND2_X1 U1418 ( .A1(n1861), .A2(DATA_IN_6_), .ZN(n1862) );
NAND2_X1 U1419 ( .A1(n1864), .A2(n1865), .ZN(U326) );
NAND2_X1 U1420 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1860), .ZN(n1865) );
NAND2_X1 U1421 ( .A1(n1861), .A2(DATA_IN_5_), .ZN(n1864) );
NAND2_X1 U1422 ( .A1(n1866), .A2(n1867), .ZN(U325) );
NAND2_X1 U1423 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1860), .ZN(n1867) );
NAND2_X1 U1424 ( .A1(n1861), .A2(DATA_IN_4_), .ZN(n1866) );
NAND2_X1 U1425 ( .A1(n1868), .A2(n1869), .ZN(U324) );
NAND2_X1 U1426 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1860), .ZN(n1869) );
NAND2_X1 U1427 ( .A1(n1861), .A2(DATA_IN_3_), .ZN(n1868) );
NAND2_X1 U1428 ( .A1(n1870), .A2(n1871), .ZN(U323) );
NAND2_X1 U1429 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1860), .ZN(n1871) );
NAND2_X1 U1430 ( .A1(n1861), .A2(DATA_IN_2_), .ZN(n1870) );
NAND2_X1 U1431 ( .A1(n1872), .A2(n1873), .ZN(U322) );
NAND2_X1 U1432 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1860), .ZN(n1873) );
NAND2_X1 U1433 ( .A1(n1861), .A2(DATA_IN_1_), .ZN(n1872) );
INV_X1 U1434 ( .A(n1874), .ZN(n1861) );
NAND2_X1 U1435 ( .A1(n1875), .A2(n1876), .ZN(U321) );
NAND2_X1 U1436 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1860), .ZN(n1876) );
NAND2_X1 U1437 ( .A1(n1741), .A2(n1877), .ZN(n1860) );
NAND2_X1 U1438 ( .A1(n1878), .A2(n1763), .ZN(n1741) );
XOR2_X1 U1439 ( .A(KEYINPUT8), .B(n1879), .Z(n1875) );
NOR2_X1 U1440 ( .A1(n1817), .A2(n1874), .ZN(n1879) );
NAND2_X1 U1441 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1877), .ZN(n1874) );
NAND2_X1 U1442 ( .A1(n1880), .A2(n1763), .ZN(n1877) );
NAND2_X1 U1443 ( .A1(n1881), .A2(n1882), .ZN(U320) );
NAND2_X1 U1444 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1740), .ZN(n1882) );
NAND2_X1 U1445 ( .A1(n1739), .A2(DATA_IN_7_), .ZN(n1881) );
NAND2_X1 U1446 ( .A1(n1883), .A2(n1884), .ZN(U319) );
NAND2_X1 U1447 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1740), .ZN(n1884) );
NAND2_X1 U1448 ( .A1(n1739), .A2(DATA_IN_6_), .ZN(n1883) );
NAND2_X1 U1449 ( .A1(n1885), .A2(n1886), .ZN(U318) );
NAND2_X1 U1450 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1740), .ZN(n1886) );
NAND2_X1 U1451 ( .A1(n1739), .A2(DATA_IN_5_), .ZN(n1885) );
NAND2_X1 U1452 ( .A1(n1887), .A2(n1888), .ZN(U317) );
NAND2_X1 U1453 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1740), .ZN(n1888) );
NAND2_X1 U1454 ( .A1(n1739), .A2(DATA_IN_4_), .ZN(n1887) );
NAND2_X1 U1455 ( .A1(n1889), .A2(n1890), .ZN(U316) );
NAND2_X1 U1456 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1740), .ZN(n1890) );
NAND2_X1 U1457 ( .A1(n1739), .A2(DATA_IN_3_), .ZN(n1889) );
NAND2_X1 U1458 ( .A1(n1891), .A2(n1892), .ZN(U315) );
NAND2_X1 U1459 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1740), .ZN(n1892) );
NAND2_X1 U1460 ( .A1(n1739), .A2(DATA_IN_2_), .ZN(n1891) );
NAND2_X1 U1461 ( .A1(n1893), .A2(n1894), .ZN(U314) );
NAND2_X1 U1462 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1740), .ZN(n1894) );
NAND2_X1 U1463 ( .A1(n1739), .A2(DATA_IN_1_), .ZN(n1893) );
NAND2_X1 U1464 ( .A1(n1895), .A2(n1896), .ZN(U313) );
NAND2_X1 U1465 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1740), .ZN(n1896) );
NAND2_X1 U1466 ( .A1(n1739), .A2(DATA_IN_0_), .ZN(n1895) );
NAND2_X1 U1467 ( .A1(n1897), .A2(n1898), .ZN(U312) );
NAND2_X1 U1468 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1740), .ZN(n1898) );
NAND2_X1 U1469 ( .A1(n1739), .A2(REG1_REG_7__SCAN_IN), .ZN(n1897) );
NAND2_X1 U1470 ( .A1(n1899), .A2(n1900), .ZN(U311) );
NAND2_X1 U1471 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1740), .ZN(n1900) );
NAND2_X1 U1472 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1739), .ZN(n1899) );
NAND2_X1 U1473 ( .A1(n1901), .A2(n1902), .ZN(U310) );
NAND2_X1 U1474 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1740), .ZN(n1902) );
NAND2_X1 U1475 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1739), .ZN(n1901) );
NAND2_X1 U1476 ( .A1(n1903), .A2(n1904), .ZN(U309) );
NAND2_X1 U1477 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1740), .ZN(n1904) );
NAND2_X1 U1478 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1739), .ZN(n1903) );
NAND2_X1 U1479 ( .A1(n1905), .A2(n1906), .ZN(U308) );
NAND2_X1 U1480 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1740), .ZN(n1906) );
NAND2_X1 U1481 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1739), .ZN(n1905) );
NAND2_X1 U1482 ( .A1(n1907), .A2(n1908), .ZN(U307) );
NAND2_X1 U1483 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1740), .ZN(n1908) );
NAND2_X1 U1484 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1739), .ZN(n1907) );
NAND2_X1 U1485 ( .A1(n1909), .A2(n1910), .ZN(U306) );
NAND2_X1 U1486 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1740), .ZN(n1910) );
NAND2_X1 U1487 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1739), .ZN(n1909) );
NAND2_X1 U1488 ( .A1(n1911), .A2(n1912), .ZN(U305) );
NAND2_X1 U1489 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1740), .ZN(n1912) );
NAND2_X1 U1490 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1739), .ZN(n1911) );
NAND2_X1 U1491 ( .A1(n1913), .A2(n1914), .ZN(U304) );
NAND2_X1 U1492 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1740), .ZN(n1914) );
NAND2_X1 U1493 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1739), .ZN(n1913) );
NAND2_X1 U1494 ( .A1(n1915), .A2(n1916), .ZN(U303) );
NAND2_X1 U1495 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1739), .ZN(n1916) );
XOR2_X1 U1496 ( .A(n1917), .B(KEYINPUT50), .Z(n1915) );
NAND2_X1 U1497 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1740), .ZN(n1917) );
NAND2_X1 U1498 ( .A1(n1918), .A2(n1919), .ZN(U302) );
NAND2_X1 U1499 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1740), .ZN(n1919) );
NAND2_X1 U1500 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1739), .ZN(n1918) );
NAND2_X1 U1501 ( .A1(n1920), .A2(n1921), .ZN(U301) );
NAND2_X1 U1502 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1922), .ZN(n1921) );
XNOR2_X1 U1503 ( .A(KEYINPUT54), .B(U280), .ZN(n1922) );
NAND2_X1 U1504 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1739), .ZN(n1920) );
NAND2_X1 U1505 ( .A1(n1923), .A2(n1924), .ZN(U300) );
NAND2_X1 U1506 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1740), .ZN(n1924) );
NAND2_X1 U1507 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1739), .ZN(n1923) );
NAND2_X1 U1508 ( .A1(n1925), .A2(n1926), .ZN(U299) );
NAND2_X1 U1509 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1740), .ZN(n1926) );
NAND2_X1 U1510 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1739), .ZN(n1925) );
NAND2_X1 U1511 ( .A1(n1927), .A2(n1928), .ZN(U298) );
NAND2_X1 U1512 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1740), .ZN(n1928) );
NAND2_X1 U1513 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1739), .ZN(n1927) );
NAND2_X1 U1514 ( .A1(n1929), .A2(n1930), .ZN(U297) );
NAND2_X1 U1515 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1740), .ZN(n1930) );
NAND2_X1 U1516 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1739), .ZN(n1929) );
NAND2_X1 U1517 ( .A1(n1931), .A2(n1932), .ZN(U296) );
NAND2_X1 U1518 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1740), .ZN(n1932) );
NAND2_X1 U1519 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1739), .ZN(n1931) );
NAND2_X1 U1520 ( .A1(n1933), .A2(n1934), .ZN(U295) );
NAND2_X1 U1521 ( .A1(n1935), .A2(n1740), .ZN(n1934) );
XNOR2_X1 U1522 ( .A(REG4_REG_6__SCAN_IN), .B(KEYINPUT47), .ZN(n1935) );
NAND2_X1 U1523 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1739), .ZN(n1933) );
NAND2_X1 U1524 ( .A1(n1936), .A2(n1937), .ZN(U294) );
NAND2_X1 U1525 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1740), .ZN(n1937) );
NAND2_X1 U1526 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1739), .ZN(n1936) );
NAND2_X1 U1527 ( .A1(n1938), .A2(n1939), .ZN(U293) );
NAND2_X1 U1528 ( .A1(n1940), .A2(REG4_REG_4__SCAN_IN), .ZN(n1939) );
XNOR2_X1 U1529 ( .A(n1740), .B(KEYINPUT24), .ZN(n1940) );
NAND2_X1 U1530 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1739), .ZN(n1938) );
NAND2_X1 U1531 ( .A1(n1941), .A2(n1942), .ZN(U292) );
NAND2_X1 U1532 ( .A1(n1739), .A2(n1943), .ZN(n1942) );
XOR2_X1 U1533 ( .A(REG3_REG_3__SCAN_IN), .B(KEYINPUT30), .Z(n1943) );
NAND2_X1 U1534 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1740), .ZN(n1941) );
NAND2_X1 U1535 ( .A1(n1944), .A2(n1945), .ZN(U291) );
NAND2_X1 U1536 ( .A1(n1946), .A2(n1739), .ZN(n1945) );
XNOR2_X1 U1537 ( .A(REG3_REG_2__SCAN_IN), .B(KEYINPUT52), .ZN(n1946) );
NAND2_X1 U1538 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1740), .ZN(n1944) );
NAND2_X1 U1539 ( .A1(n1947), .A2(n1948), .ZN(U290) );
NAND2_X1 U1540 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1740), .ZN(n1948) );
NAND2_X1 U1541 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1739), .ZN(n1947) );
NAND2_X1 U1542 ( .A1(n1949), .A2(n1950), .ZN(U289) );
NAND2_X1 U1543 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1740), .ZN(n1950) );
NAND2_X1 U1544 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1739), .ZN(n1949) );
NAND2_X1 U1545 ( .A1(n1951), .A2(n1952), .ZN(U288) );
NAND2_X1 U1546 ( .A1(n1953), .A2(REG4_REG_7__SCAN_IN), .ZN(n1952) );
XOR2_X1 U1547 ( .A(n1954), .B(KEYINPUT62), .Z(n1951) );
NAND3_X1 U1548 ( .A1(n1955), .A2(n1956), .A3(n1957), .ZN(n1954) );
NAND2_X1 U1549 ( .A1(n1958), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1956) );
NAND2_X1 U1550 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1740), .ZN(n1955) );
NAND4_X1 U1551 ( .A1(n1959), .A2(n1960), .A3(n1957), .A4(n1961), .ZN(U287));
NOR3_X1 U1552 ( .A1(n1962), .A2(n1963), .A3(n1964), .ZN(n1961) );
NOR3_X1 U1553 ( .A1(n1965), .A2(n1966), .A3(n1967), .ZN(n1964) );
NOR2_X1 U1554 ( .A1(n1968), .A2(n1969), .ZN(n1967) );
INV_X1 U1555 ( .A(KEYINPUT4), .ZN(n1969) );
NOR2_X1 U1556 ( .A1(n1970), .A2(n1971), .ZN(n1968) );
NOR2_X1 U1557 ( .A1(KEYINPUT4), .A2(n1971), .ZN(n1966) );
NOR4_X1 U1558 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .ZN(n1963));
AND2_X1 U1559 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1958), .ZN(n1962) );
AND2_X1 U1560 ( .A1(n1976), .A2(n1977), .ZN(n1957) );
NAND3_X1 U1561 ( .A1(n1970), .A2(n1971), .A3(n1978), .ZN(n1977) );
NAND3_X1 U1562 ( .A1(n1979), .A2(n1980), .A3(n1972), .ZN(n1976) );
AND2_X1 U1563 ( .A1(n1981), .A2(n1982), .ZN(n1972) );
XNOR2_X1 U1564 ( .A(KEYINPUT37), .B(n1983), .ZN(n1982) );
XNOR2_X1 U1565 ( .A(n1984), .B(KEYINPUT43), .ZN(n1981) );
OR2_X1 U1566 ( .A1(n1974), .A2(n1973), .ZN(n1980) );
NAND2_X1 U1567 ( .A1(n1953), .A2(REG4_REG_6__SCAN_IN), .ZN(n1960) );
NAND2_X1 U1568 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1740), .ZN(n1959) );
NAND4_X1 U1569 ( .A1(n1985), .A2(n1986), .A3(n1987), .A4(n1988), .ZN(U286));
NOR3_X1 U1570 ( .A1(n1989), .A2(n1990), .A3(n1991), .ZN(n1988) );
AND2_X1 U1571 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1958), .ZN(n1991) );
NOR2_X1 U1572 ( .A1(U280), .A2(n1992), .ZN(n1990) );
XOR2_X1 U1573 ( .A(KEYINPUT29), .B(DATA_OUT_REG_5__SCAN_IN), .Z(n1992) );
NOR2_X1 U1574 ( .A1(n1993), .A2(n1994), .ZN(n1989) );
NAND2_X1 U1575 ( .A1(n1979), .A2(n1995), .ZN(n1987) );
XNOR2_X1 U1576 ( .A(n1996), .B(n1973), .ZN(n1995) );
XNOR2_X1 U1577 ( .A(n1984), .B(n1997), .ZN(n1973) );
NOR2_X1 U1578 ( .A1(KEYINPUT43), .A2(n1983), .ZN(n1997) );
NAND3_X1 U1579 ( .A1(n1998), .A2(n1999), .A3(n2000), .ZN(n1986) );
XOR2_X1 U1580 ( .A(n1971), .B(KEYINPUT49), .Z(n2000) );
NAND2_X1 U1581 ( .A1(n2001), .A2(n2002), .ZN(n1971) );
XOR2_X1 U1582 ( .A(KEYINPUT28), .B(n2003), .Z(n2002) );
NAND2_X1 U1583 ( .A1(n2003), .A2(n2004), .ZN(n1999) );
INV_X1 U1584 ( .A(n2001), .ZN(n2004) );
NOR2_X1 U1585 ( .A1(n2005), .A2(n1970), .ZN(n2003) );
NOR2_X1 U1586 ( .A1(n2006), .A2(n1984), .ZN(n1970) );
AND2_X1 U1587 ( .A1(n1984), .A2(n2006), .ZN(n2005) );
XNOR2_X1 U1588 ( .A(n1978), .B(KEYINPUT21), .ZN(n1998) );
NAND2_X1 U1589 ( .A1(n1984), .A2(n2007), .ZN(n1985) );
XNOR2_X1 U1590 ( .A(KEYINPUT32), .B(n2008), .ZN(n2007) );
AND2_X1 U1591 ( .A1(n2009), .A2(n2010), .ZN(n1984) );
NAND4_X1 U1592 ( .A1(n2011), .A2(n2012), .A3(n2013), .A4(n2014), .ZN(n2010));
NAND2_X1 U1593 ( .A1(n2015), .A2(n2016), .ZN(n2014) );
XNOR2_X1 U1594 ( .A(n2017), .B(DATA_IN_6_), .ZN(n2015) );
NAND2_X1 U1595 ( .A1(n2018), .A2(RESTART), .ZN(n2013) );
XNOR2_X1 U1596 ( .A(n1826), .B(RMAX_REG_6__SCAN_IN), .ZN(n2018) );
NAND2_X1 U1597 ( .A1(n2019), .A2(n2020), .ZN(n2012) );
XNOR2_X1 U1598 ( .A(KEYINPUT11), .B(n2021), .ZN(n2011) );
NAND4_X1 U1599 ( .A1(n2022), .A2(n2020), .A3(n2023), .A4(n2024), .ZN(n2009));
NAND2_X1 U1600 ( .A1(n2025), .A2(n2016), .ZN(n2024) );
XNOR2_X1 U1601 ( .A(REG4_REG_6__SCAN_IN), .B(DATA_IN_6_), .ZN(n2025) );
NAND2_X1 U1602 ( .A1(n2026), .A2(RESTART), .ZN(n2023) );
XNOR2_X1 U1603 ( .A(RMAX_REG_6__SCAN_IN), .B(RMIN_REG_6__SCAN_IN), .ZN(n2026) );
NAND2_X1 U1604 ( .A1(n2021), .A2(n2027), .ZN(n2022) );
NAND4_X1 U1605 ( .A1(n2028), .A2(n2029), .A3(n2030), .A4(n2031), .ZN(U285));
NOR3_X1 U1606 ( .A1(n2032), .A2(n2033), .A3(n2034), .ZN(n2031) );
NOR3_X1 U1607 ( .A1(n1965), .A2(n2035), .A3(n2001), .ZN(n2034) );
NOR2_X1 U1608 ( .A1(n2036), .A2(n2037), .ZN(n2001) );
AND2_X1 U1609 ( .A1(n2038), .A2(n2006), .ZN(n2037) );
AND3_X1 U1610 ( .A1(n2038), .A2(n2036), .A3(n2006), .ZN(n2035) );
NAND3_X1 U1611 ( .A1(n2039), .A2(n2040), .A3(n2041), .ZN(n2006) );
NAND2_X1 U1612 ( .A1(n2042), .A2(n2043), .ZN(n2036) );
NAND2_X1 U1613 ( .A1(n2044), .A2(n2045), .ZN(n2038) );
NAND2_X1 U1614 ( .A1(n2041), .A2(n2040), .ZN(n2045) );
NOR3_X1 U1615 ( .A1(n1975), .A2(n1996), .A3(n2046), .ZN(n2033) );
NOR3_X1 U1616 ( .A1(n2047), .A2(n2048), .A3(n2049), .ZN(n2046) );
INV_X1 U1617 ( .A(n1983), .ZN(n2049) );
NAND2_X1 U1618 ( .A1(n2039), .A2(n2050), .ZN(n1983) );
XOR2_X1 U1619 ( .A(KEYINPUT36), .B(n2051), .Z(n2050) );
NOR2_X1 U1620 ( .A1(n2051), .A2(n2039), .ZN(n2047) );
INV_X1 U1621 ( .A(n1974), .ZN(n1996) );
NAND2_X1 U1622 ( .A1(n2052), .A2(n2048), .ZN(n1974) );
XNOR2_X1 U1623 ( .A(n2051), .B(n2053), .ZN(n2052) );
NOR2_X1 U1624 ( .A1(KEYINPUT36), .A2(n2044), .ZN(n2053) );
NOR2_X1 U1625 ( .A1(n2039), .A2(n2008), .ZN(n2032) );
INV_X1 U1626 ( .A(n2044), .ZN(n2039) );
NAND2_X1 U1627 ( .A1(n2054), .A2(n2055), .ZN(n2044) );
NAND2_X1 U1628 ( .A1(n2019), .A2(n2056), .ZN(n2055) );
NAND2_X1 U1629 ( .A1(n2021), .A2(n2020), .ZN(n2056) );
INV_X1 U1630 ( .A(n2027), .ZN(n2019) );
NAND4_X1 U1631 ( .A1(n2057), .A2(n2058), .A3(n2020), .A4(n2027), .ZN(n2054));
NAND2_X1 U1632 ( .A1(n2059), .A2(n2060), .ZN(n2027) );
NAND2_X1 U1633 ( .A1(n2061), .A2(n2062), .ZN(n2060) );
NAND2_X1 U1634 ( .A1(n2063), .A2(n2064), .ZN(n2062) );
OR2_X1 U1635 ( .A1(n2064), .A2(n2063), .ZN(n2059) );
NAND3_X1 U1636 ( .A1(n2065), .A2(n2066), .A3(n2067), .ZN(n2020) );
NAND2_X1 U1637 ( .A1(REG4_REG_5__SCAN_IN), .A2(n2016), .ZN(n2066) );
NAND2_X1 U1638 ( .A1(RESTART), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2065) );
OR2_X1 U1639 ( .A1(n2068), .A2(KEYINPUT17), .ZN(n2058) );
NAND2_X1 U1640 ( .A1(n2069), .A2(KEYINPUT17), .ZN(n2057) );
INV_X1 U1641 ( .A(n2021), .ZN(n2069) );
NAND3_X1 U1642 ( .A1(n2070), .A2(n2071), .A3(n2068), .ZN(n2021) );
INV_X1 U1643 ( .A(n2067), .ZN(n2068) );
NAND2_X1 U1644 ( .A1(n2072), .A2(n2073), .ZN(n2067) );
NAND2_X1 U1645 ( .A1(RESTART), .A2(n1857), .ZN(n2073) );
NAND2_X1 U1646 ( .A1(n1824), .A2(n2016), .ZN(n2072) );
INV_X1 U1647 ( .A(DATA_IN_5_), .ZN(n1824) );
NAND2_X1 U1648 ( .A1(RESTART), .A2(n1801), .ZN(n2071) );
NAND2_X1 U1649 ( .A1(n1993), .A2(n2016), .ZN(n2070) );
NAND2_X1 U1650 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1740), .ZN(n2030) );
NAND2_X1 U1651 ( .A1(n1958), .A2(RLAST_REG_4__SCAN_IN), .ZN(n2029) );
NAND2_X1 U1652 ( .A1(n1953), .A2(REG4_REG_4__SCAN_IN), .ZN(n2028) );
NAND4_X1 U1653 ( .A1(n2074), .A2(n2075), .A3(n2076), .A4(n2077), .ZN(U284));
NOR3_X1 U1654 ( .A1(n2078), .A2(n2079), .A3(n2080), .ZN(n2077) );
NOR2_X1 U1655 ( .A1(n2081), .A2(n1965), .ZN(n2080) );
XNOR2_X1 U1656 ( .A(n2042), .B(n2043), .ZN(n2081) );
XNOR2_X1 U1657 ( .A(n2082), .B(n2083), .ZN(n2043) );
NOR2_X1 U1658 ( .A1(KEYINPUT63), .A2(n2040), .ZN(n2083) );
NOR3_X1 U1659 ( .A1(n1975), .A2(n2048), .A3(n2084), .ZN(n2079) );
XOR2_X1 U1660 ( .A(n2085), .B(KEYINPUT26), .Z(n2084) );
NAND2_X1 U1661 ( .A1(n2086), .A2(n2087), .ZN(n2085) );
NOR2_X1 U1662 ( .A1(n2088), .A2(n2086), .ZN(n2048) );
NOR2_X1 U1663 ( .A1(n2089), .A2(n2051), .ZN(n2086) );
AND2_X1 U1664 ( .A1(n2090), .A2(n2040), .ZN(n2051) );
NOR2_X1 U1665 ( .A1(n2040), .A2(n2090), .ZN(n2089) );
XNOR2_X1 U1666 ( .A(n2087), .B(KEYINPUT34), .ZN(n2088) );
NOR2_X1 U1667 ( .A1(n2040), .A2(n2008), .ZN(n2078) );
XOR2_X1 U1668 ( .A(n2061), .B(n2091), .Z(n2040) );
NOR2_X1 U1669 ( .A1(n2092), .A2(n2093), .ZN(n2091) );
NOR2_X1 U1670 ( .A1(n2094), .A2(n2095), .ZN(n2093) );
NOR2_X1 U1671 ( .A1(KEYINPUT44), .A2(n2064), .ZN(n2094) );
NOR2_X1 U1672 ( .A1(n2063), .A2(n2064), .ZN(n2092) );
NAND2_X1 U1673 ( .A1(n2096), .A2(n2097), .ZN(n2064) );
NAND2_X1 U1674 ( .A1(RESTART), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2097) );
XOR2_X1 U1675 ( .A(n2098), .B(KEYINPUT7), .Z(n2096) );
NAND2_X1 U1676 ( .A1(n2099), .A2(n2016), .ZN(n2098) );
XNOR2_X1 U1677 ( .A(REG4_REG_4__SCAN_IN), .B(KEYINPUT9), .ZN(n2099) );
INV_X1 U1678 ( .A(n2095), .ZN(n2063) );
NAND2_X1 U1679 ( .A1(n2100), .A2(n2101), .ZN(n2095) );
NAND2_X1 U1680 ( .A1(n2102), .A2(n2103), .ZN(n2101) );
OR2_X1 U1681 ( .A1(n2104), .A2(n2105), .ZN(n2102) );
NAND2_X1 U1682 ( .A1(n2104), .A2(n2105), .ZN(n2100) );
AND2_X1 U1683 ( .A1(n2106), .A2(n2107), .ZN(n2061) );
NAND2_X1 U1684 ( .A1(DATA_IN_4_), .A2(n2016), .ZN(n2107) );
NAND2_X1 U1685 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2106) );
NAND2_X1 U1686 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1740), .ZN(n2076) );
NAND2_X1 U1687 ( .A1(n1958), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2075) );
NAND2_X1 U1688 ( .A1(n1953), .A2(REG4_REG_3__SCAN_IN), .ZN(n2074) );
NAND4_X1 U1689 ( .A1(n2108), .A2(n2109), .A3(n2110), .A4(n2111), .ZN(U283));
NOR3_X1 U1690 ( .A1(n2112), .A2(n2113), .A3(n2114), .ZN(n2111) );
NOR3_X1 U1691 ( .A1(n1975), .A2(n2115), .A3(n2116), .ZN(n2114) );
XOR2_X1 U1692 ( .A(n2087), .B(KEYINPUT41), .Z(n2116) );
NAND3_X1 U1693 ( .A1(n2117), .A2(n2118), .A3(n2119), .ZN(n2087) );
NAND2_X1 U1694 ( .A1(n2120), .A2(n2121), .ZN(n2117) );
INV_X1 U1695 ( .A(n2090), .ZN(n2121) );
NAND2_X1 U1696 ( .A1(n2122), .A2(n2123), .ZN(n2120) );
NOR3_X1 U1697 ( .A1(n2124), .A2(n2090), .A3(n2125), .ZN(n2115) );
NOR2_X1 U1698 ( .A1(n2126), .A2(n2127), .ZN(n2125) );
NOR2_X1 U1699 ( .A1(n2122), .A2(n2123), .ZN(n2090) );
AND2_X1 U1700 ( .A1(n2118), .A2(n2119), .ZN(n2124) );
NOR3_X1 U1701 ( .A1(n1965), .A2(n2042), .A3(n2128), .ZN(n2113) );
NOR2_X1 U1702 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
NOR2_X1 U1703 ( .A1(n2131), .A2(n2132), .ZN(n2129) );
AND3_X1 U1704 ( .A1(n2133), .A2(n2134), .A3(n2130), .ZN(n2042) );
NAND2_X1 U1705 ( .A1(n2082), .A2(n2135), .ZN(n2130) );
NAND2_X1 U1706 ( .A1(n2136), .A2(n2122), .ZN(n2135) );
INV_X1 U1707 ( .A(n2041), .ZN(n2082) );
NOR2_X1 U1708 ( .A1(n2122), .A2(n2136), .ZN(n2041) );
INV_X1 U1709 ( .A(n2137), .ZN(n2136) );
NOR2_X1 U1710 ( .A1(n2127), .A2(n2008), .ZN(n2112) );
INV_X1 U1711 ( .A(n2122), .ZN(n2127) );
XOR2_X1 U1712 ( .A(n2138), .B(n2105), .Z(n2122) );
NAND2_X1 U1713 ( .A1(n2139), .A2(n2140), .ZN(n2105) );
NAND2_X1 U1714 ( .A1(RESTART), .A2(n1809), .ZN(n2140) );
NAND2_X1 U1715 ( .A1(n2141), .A2(n2016), .ZN(n2139) );
NAND2_X1 U1716 ( .A1(n2142), .A2(n2143), .ZN(n2138) );
NAND2_X1 U1717 ( .A1(n2144), .A2(n2145), .ZN(n2143) );
NAND2_X1 U1718 ( .A1(KEYINPUT39), .A2(n2104), .ZN(n2145) );
INV_X1 U1719 ( .A(n2103), .ZN(n2144) );
NAND2_X1 U1720 ( .A1(n2104), .A2(n2103), .ZN(n2142) );
NAND2_X1 U1721 ( .A1(n2146), .A2(n2147), .ZN(n2103) );
NAND2_X1 U1722 ( .A1(n2148), .A2(n2149), .ZN(n2147) );
OR2_X1 U1723 ( .A1(n2150), .A2(n2151), .ZN(n2148) );
NAND2_X1 U1724 ( .A1(n2151), .A2(n2150), .ZN(n2146) );
NAND2_X1 U1725 ( .A1(n2152), .A2(n2153), .ZN(n2104) );
NAND2_X1 U1726 ( .A1(RESTART), .A2(n1856), .ZN(n2153) );
NAND2_X1 U1727 ( .A1(n1847), .A2(n2016), .ZN(n2152) );
NAND2_X1 U1728 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1740), .ZN(n2110) );
NAND2_X1 U1729 ( .A1(n1958), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2109) );
NAND2_X1 U1730 ( .A1(n1953), .A2(REG4_REG_2__SCAN_IN), .ZN(n2108) );
INV_X1 U1731 ( .A(n1994), .ZN(n1953) );
NAND4_X1 U1732 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(U282));
NOR3_X1 U1733 ( .A1(n2158), .A2(n2159), .A3(n2160), .ZN(n2157) );
NOR2_X1 U1734 ( .A1(n1975), .A2(n2161), .ZN(n2160) );
XNOR2_X1 U1735 ( .A(n2119), .B(n2118), .ZN(n2161) );
NAND2_X1 U1736 ( .A1(n2123), .A2(n2162), .ZN(n2118) );
INV_X1 U1737 ( .A(n2126), .ZN(n2123) );
INV_X1 U1738 ( .A(n2163), .ZN(n2119) );
NOR2_X1 U1739 ( .A1(n1994), .A2(n2164), .ZN(n2159) );
XNOR2_X1 U1740 ( .A(n2165), .B(KEYINPUT48), .ZN(n2164) );
NOR3_X1 U1741 ( .A1(n1965), .A2(n2166), .A3(n2167), .ZN(n2158) );
NOR3_X1 U1742 ( .A1(n2132), .A2(n2131), .A3(n2168), .ZN(n2167) );
NOR2_X1 U1743 ( .A1(KEYINPUT1), .A2(n2169), .ZN(n2168) );
INV_X1 U1744 ( .A(n2133), .ZN(n2132) );
NOR2_X1 U1745 ( .A1(n2170), .A2(n2133), .ZN(n2166) );
NAND2_X1 U1746 ( .A1(n2171), .A2(n2162), .ZN(n2133) );
NAND2_X1 U1747 ( .A1(n2172), .A2(n2173), .ZN(n2162) );
XNOR2_X1 U1748 ( .A(KEYINPUT56), .B(n2137), .ZN(n2171) );
NAND2_X1 U1749 ( .A1(n2174), .A2(n2175), .ZN(n2137) );
OR4_X1 U1750 ( .A1(n2172), .A2(n2176), .A3(n2177), .A4(KEYINPUT27), .ZN(n2175) );
NAND2_X1 U1751 ( .A1(KEYINPUT27), .A2(n2126), .ZN(n2174) );
NOR2_X1 U1752 ( .A1(n2173), .A2(n2172), .ZN(n2126) );
NOR2_X1 U1753 ( .A1(n2169), .A2(n2178), .ZN(n2170) );
INV_X1 U1754 ( .A(KEYINPUT1), .ZN(n2178) );
XNOR2_X1 U1755 ( .A(n2134), .B(KEYINPUT15), .ZN(n2169) );
INV_X1 U1756 ( .A(n1978), .ZN(n1965) );
XOR2_X1 U1757 ( .A(KEYINPUT18), .B(n2179), .Z(n2156) );
AND2_X1 U1758 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1958), .ZN(n2179) );
NAND2_X1 U1759 ( .A1(n2180), .A2(n2172), .ZN(n2155) );
XNOR2_X1 U1760 ( .A(n2150), .B(n2181), .ZN(n2172) );
XOR2_X1 U1761 ( .A(n2149), .B(n2151), .Z(n2181) );
NAND2_X1 U1762 ( .A1(n2182), .A2(n2183), .ZN(n2151) );
NAND2_X1 U1763 ( .A1(RESTART), .A2(n1820), .ZN(n2183) );
NAND2_X1 U1764 ( .A1(n2184), .A2(n2016), .ZN(n2182) );
NAND2_X1 U1765 ( .A1(n2185), .A2(n2186), .ZN(n2149) );
NAND2_X1 U1766 ( .A1(n2187), .A2(n2188), .ZN(n2186) );
NAND2_X1 U1767 ( .A1(n2189), .A2(n2190), .ZN(n2188) );
NAND2_X1 U1768 ( .A1(n2191), .A2(n2192), .ZN(n2185) );
NAND2_X1 U1769 ( .A1(n2193), .A2(n2194), .ZN(n2150) );
NAND2_X1 U1770 ( .A1(RESTART), .A2(n1851), .ZN(n2194) );
NAND2_X1 U1771 ( .A1(n1813), .A2(n2016), .ZN(n2193) );
INV_X1 U1772 ( .A(n2008), .ZN(n2180) );
NAND2_X1 U1773 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1740), .ZN(n2154) );
NAND4_X1 U1774 ( .A1(n2195), .A2(n2196), .A3(n2197), .A4(n2198), .ZN(U281));
NOR3_X1 U1775 ( .A1(n2199), .A2(n2200), .A3(n2201), .ZN(n2198) );
NOR2_X1 U1776 ( .A1(n2177), .A2(n2008), .ZN(n2201) );
NAND4_X1 U1777 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2202), .A3(n2203), .A4(U280), .ZN(n2008) );
NAND2_X1 U1778 ( .A1(n2204), .A2(n2205), .ZN(n2202) );
NAND2_X1 U1779 ( .A1(n2206), .A2(n2207), .ZN(n2205) );
XNOR2_X1 U1780 ( .A(KEYINPUT12), .B(n2208), .ZN(n2207) );
XNOR2_X1 U1781 ( .A(RESTART), .B(KEYINPUT45), .ZN(n2204) );
INV_X1 U1782 ( .A(n2209), .ZN(n2177) );
NOR2_X1 U1783 ( .A1(n2210), .A2(n2211), .ZN(n2200) );
INV_X1 U1784 ( .A(RLAST_REG_0__SCAN_IN), .ZN(n2211) );
XNOR2_X1 U1785 ( .A(n1958), .B(KEYINPUT0), .ZN(n2210) );
AND2_X1 U1786 ( .A1(n2212), .A2(n1880), .ZN(n1958) );
INV_X1 U1787 ( .A(ENABLE), .ZN(n1880) );
NOR2_X1 U1788 ( .A1(n2213), .A2(n1994), .ZN(n2199) );
NAND3_X1 U1789 ( .A1(AVERAGE), .A2(n2212), .A3(ENABLE), .ZN(n1994) );
NAND2_X1 U1790 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1740), .ZN(n2197) );
NAND2_X1 U1791 ( .A1(n2131), .A2(n1978), .ZN(n2196) );
NOR3_X1 U1792 ( .A1(n1878), .A2(n1740), .A3(n2203), .ZN(n1978) );
NAND3_X1 U1793 ( .A1(n2214), .A2(n2215), .A3(RESTART), .ZN(n2203) );
NAND3_X1 U1794 ( .A1(n2216), .A2(n2217), .A3(n2218), .ZN(n2215) );
NAND2_X1 U1795 ( .A1(n2219), .A2(n1835), .ZN(n2218) );
NAND2_X1 U1796 ( .A1(n2220), .A2(n1826), .ZN(n2217) );
INV_X1 U1797 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1826) );
OR2_X1 U1798 ( .A1(n2219), .A2(n1835), .ZN(n2220) );
INV_X1 U1799 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1835) );
NAND2_X1 U1800 ( .A1(n2221), .A2(n2222), .ZN(n2219) );
NAND2_X1 U1801 ( .A1(n2223), .A2(n1801), .ZN(n2222) );
INV_X1 U1802 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1801) );
NAND2_X1 U1803 ( .A1(n2224), .A2(n2225), .ZN(n2223) );
XNOR2_X1 U1804 ( .A(n1857), .B(KEYINPUT2), .ZN(n2224) );
INV_X1 U1805 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1857) );
OR2_X1 U1806 ( .A1(n2225), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2221) );
NAND2_X1 U1807 ( .A1(n2226), .A2(n2227), .ZN(n2225) );
NAND3_X1 U1808 ( .A1(n2228), .A2(n2229), .A3(n2230), .ZN(n2227) );
NAND2_X1 U1809 ( .A1(n2231), .A2(n1823), .ZN(n2230) );
NAND3_X1 U1810 ( .A1(n2232), .A2(n2233), .A3(n2234), .ZN(n2229) );
NAND2_X1 U1811 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2234) );
NAND3_X1 U1812 ( .A1(n2235), .A2(n2236), .A3(n2237), .ZN(n2233) );
NAND2_X1 U1813 ( .A1(n1851), .A2(n1820), .ZN(n2237) );
INV_X1 U1814 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1820) );
INV_X1 U1815 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1851) );
NAND2_X1 U1816 ( .A1(n2238), .A2(n1855), .ZN(n2236) );
NAND2_X1 U1817 ( .A1(n2239), .A2(n2240), .ZN(n2238) );
XNOR2_X1 U1818 ( .A(n1818), .B(KEYINPUT20), .ZN(n2240) );
INV_X1 U1819 ( .A(n2241), .ZN(n2239) );
NAND2_X1 U1820 ( .A1(n2241), .A2(n1818), .ZN(n2235) );
NAND2_X1 U1821 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2241) );
NAND2_X1 U1822 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2232) );
NAND2_X1 U1823 ( .A1(n1856), .A2(n1809), .ZN(n2228) );
INV_X1 U1824 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1809) );
INV_X1 U1825 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1856) );
XOR2_X1 U1826 ( .A(KEYINPUT14), .B(n2242), .Z(n2226) );
NOR2_X1 U1827 ( .A1(n2231), .A2(n1823), .ZN(n2242) );
INV_X1 U1828 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1823) );
INV_X1 U1829 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n2231) );
NAND2_X1 U1830 ( .A1(n2243), .A2(RMIN_REG_7__SCAN_IN), .ZN(n2216) );
XNOR2_X1 U1831 ( .A(RMAX_REG_7__SCAN_IN), .B(KEYINPUT59), .ZN(n2243) );
NAND2_X1 U1832 ( .A1(n1831), .A2(n1827), .ZN(n2214) );
INV_X1 U1833 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1827) );
INV_X1 U1834 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1831) );
INV_X1 U1835 ( .A(n2134), .ZN(n2131) );
NAND2_X1 U1836 ( .A1(n2173), .A2(n2244), .ZN(n2134) );
NAND2_X1 U1837 ( .A1(n2176), .A2(n2209), .ZN(n2244) );
NAND2_X1 U1838 ( .A1(n1979), .A2(n2163), .ZN(n2195) );
NAND3_X1 U1839 ( .A1(n2245), .A2(n2246), .A3(n2247), .ZN(n2163) );
XOR2_X1 U1840 ( .A(n2248), .B(KEYINPUT58), .Z(n2247) );
NAND2_X1 U1841 ( .A1(n2249), .A2(n2250), .ZN(n2248) );
OR2_X1 U1842 ( .A1(n2173), .A2(KEYINPUT60), .ZN(n2250) );
INV_X1 U1843 ( .A(n2251), .ZN(n2173) );
NAND3_X1 U1844 ( .A1(n2209), .A2(n2252), .A3(KEYINPUT60), .ZN(n2249) );
OR3_X1 U1845 ( .A1(n2252), .A2(n2209), .A3(KEYINPUT23), .ZN(n2246) );
NAND2_X1 U1846 ( .A1(KEYINPUT23), .A2(n2251), .ZN(n2245) );
NOR2_X1 U1847 ( .A1(n2209), .A2(n2176), .ZN(n2251) );
INV_X1 U1848 ( .A(n2252), .ZN(n2176) );
NAND3_X1 U1849 ( .A1(n2253), .A2(n2254), .A3(n2255), .ZN(n2252) );
NAND2_X1 U1850 ( .A1(n2256), .A2(n2257), .ZN(n2255) );
NAND2_X1 U1851 ( .A1(KEYINPUT33), .A2(n2258), .ZN(n2257) );
INV_X1 U1852 ( .A(n2259), .ZN(n2258) );
NAND3_X1 U1853 ( .A1(KEYINPUT33), .A2(n2189), .A3(n2260), .ZN(n2254) );
INV_X1 U1854 ( .A(KEYINPUT3), .ZN(n2260) );
NAND2_X1 U1855 ( .A1(KEYINPUT3), .A2(n2259), .ZN(n2253) );
NAND2_X1 U1856 ( .A1(n2261), .A2(n2262), .ZN(n2209) );
NAND2_X1 U1857 ( .A1(n2191), .A2(n2263), .ZN(n2262) );
XOR2_X1 U1858 ( .A(n2264), .B(KEYINPUT10), .Z(n2263) );
NAND3_X1 U1859 ( .A1(n2265), .A2(n2266), .A3(n2267), .ZN(n2264) );
OR2_X1 U1860 ( .A1(n2268), .A2(KEYINPUT19), .ZN(n2267) );
NAND3_X1 U1861 ( .A1(KEYINPUT19), .A2(n2268), .A3(n2192), .ZN(n2266) );
INV_X1 U1862 ( .A(n2189), .ZN(n2192) );
NAND2_X1 U1863 ( .A1(n2189), .A2(n2269), .ZN(n2265) );
NAND2_X1 U1864 ( .A1(KEYINPUT19), .A2(n2270), .ZN(n2269) );
XNOR2_X1 U1865 ( .A(n2268), .B(KEYINPUT61), .ZN(n2270) );
NAND2_X1 U1866 ( .A1(n2271), .A2(n2190), .ZN(n2261) );
INV_X1 U1867 ( .A(n2191), .ZN(n2190) );
NAND2_X1 U1868 ( .A1(n2272), .A2(n2273), .ZN(n2191) );
NAND2_X1 U1869 ( .A1(RESTART), .A2(n1855), .ZN(n2273) );
INV_X1 U1870 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1855) );
NAND2_X1 U1871 ( .A1(n1819), .A2(n2016), .ZN(n2272) );
INV_X1 U1872 ( .A(DATA_IN_1_), .ZN(n1819) );
XNOR2_X1 U1873 ( .A(n2268), .B(n2189), .ZN(n2271) );
NOR2_X1 U1874 ( .A1(n2259), .A2(n2256), .ZN(n2189) );
AND2_X1 U1875 ( .A1(n2274), .A2(n2275), .ZN(n2256) );
NAND2_X1 U1876 ( .A1(REG4_REG_0__SCAN_IN), .A2(n2016), .ZN(n2275) );
NAND2_X1 U1877 ( .A1(RESTART), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2274) );
NAND2_X1 U1878 ( .A1(n2276), .A2(n2277), .ZN(n2259) );
OR2_X1 U1879 ( .A1(n2016), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2277) );
NAND2_X1 U1880 ( .A1(n1817), .A2(n2016), .ZN(n2276) );
INV_X1 U1881 ( .A(n2187), .ZN(n2268) );
NAND2_X1 U1882 ( .A1(n2278), .A2(n2279), .ZN(n2187) );
NAND2_X1 U1883 ( .A1(RESTART), .A2(n1818), .ZN(n2279) );
INV_X1 U1884 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1818) );
NAND2_X1 U1885 ( .A1(n2165), .A2(n2016), .ZN(n2278) );
INV_X1 U1886 ( .A(RESTART), .ZN(n2016) );
INV_X1 U1887 ( .A(n1975), .ZN(n1979) );
NAND3_X1 U1888 ( .A1(n2206), .A2(n2212), .A3(n2280), .ZN(n1975) );
XOR2_X1 U1889 ( .A(n2208), .B(KEYINPUT12), .Z(n2280) );
NAND2_X1 U1890 ( .A1(n2281), .A2(n2282), .ZN(n2208) );
NAND2_X1 U1891 ( .A1(n2283), .A2(n2284), .ZN(n2282) );
INV_X1 U1892 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2284) );
NAND2_X1 U1893 ( .A1(DATA_IN_7_), .A2(n2285), .ZN(n2283) );
OR2_X1 U1894 ( .A1(n2285), .A2(DATA_IN_7_), .ZN(n2281) );
NAND2_X1 U1895 ( .A1(n2286), .A2(n2287), .ZN(n2285) );
NAND2_X1 U1896 ( .A1(n2288), .A2(n2017), .ZN(n2287) );
INV_X1 U1897 ( .A(REG4_REG_6__SCAN_IN), .ZN(n2017) );
NAND2_X1 U1898 ( .A1(n2289), .A2(DATA_IN_6_), .ZN(n2288) );
XOR2_X1 U1899 ( .A(KEYINPUT51), .B(n2290), .Z(n2286) );
NOR2_X1 U1900 ( .A1(n2289), .A2(DATA_IN_6_), .ZN(n2290) );
AND2_X1 U1901 ( .A1(n2291), .A2(n2292), .ZN(n2289) );
NAND2_X1 U1902 ( .A1(n1993), .A2(n2293), .ZN(n2292) );
NAND2_X1 U1903 ( .A1(DATA_IN_5_), .A2(n2294), .ZN(n2293) );
INV_X1 U1904 ( .A(REG4_REG_5__SCAN_IN), .ZN(n1993) );
OR2_X1 U1905 ( .A1(n2294), .A2(DATA_IN_5_), .ZN(n2291) );
NAND2_X1 U1906 ( .A1(n2295), .A2(n2296), .ZN(n2294) );
NAND2_X1 U1907 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2296) );
NAND3_X1 U1908 ( .A1(n2297), .A2(n2298), .A3(n2299), .ZN(n2295) );
OR2_X1 U1909 ( .A1(DATA_IN_4_), .A2(REG4_REG_4__SCAN_IN), .ZN(n2299) );
NAND3_X1 U1910 ( .A1(n2300), .A2(n2301), .A3(n2302), .ZN(n2298) );
XOR2_X1 U1911 ( .A(n2303), .B(KEYINPUT13), .Z(n2302) );
NAND3_X1 U1912 ( .A1(n2304), .A2(n2305), .A3(n2306), .ZN(n2303) );
NAND2_X1 U1913 ( .A1(n1813), .A2(n2184), .ZN(n2306) );
INV_X1 U1914 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2184) );
INV_X1 U1915 ( .A(DATA_IN_2_), .ZN(n1813) );
NAND2_X1 U1916 ( .A1(n2307), .A2(n2165), .ZN(n2305) );
INV_X1 U1917 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2165) );
NAND2_X1 U1918 ( .A1(n2308), .A2(DATA_IN_1_), .ZN(n2307) );
OR2_X1 U1919 ( .A1(n2308), .A2(DATA_IN_1_), .ZN(n2304) );
NOR2_X1 U1920 ( .A1(n2213), .A2(n1817), .ZN(n2308) );
INV_X1 U1921 ( .A(DATA_IN_0_), .ZN(n1817) );
INV_X1 U1922 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2213) );
NAND2_X1 U1923 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2301) );
NAND2_X1 U1924 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2300) );
NAND2_X1 U1925 ( .A1(n1847), .A2(n2141), .ZN(n2297) );
INV_X1 U1926 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2141) );
INV_X1 U1927 ( .A(DATA_IN_3_), .ZN(n1847) );
NOR3_X1 U1928 ( .A1(n1740), .A2(RESTART), .A3(n1878), .ZN(n2212) );
AND2_X1 U1929 ( .A1(ENABLE), .A2(n2309), .ZN(n2206) );
XOR2_X1 U1930 ( .A(KEYINPUT42), .B(AVERAGE), .Z(n2309) );
INV_X1 U1931 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1878) );
NOR2_X1 U1932 ( .A1(n1763), .A2(STATO_REG_1__SCAN_IN), .ZN(n2310) );
INV_X1 U1933 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1763) );
endmodule


