//Key = 0000101001000111101000010010100100111101001110111110100100100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346;

XOR2_X1 U739 ( .A(n1027), .B(n1028), .Z(G9) );
NOR2_X1 U740 ( .A1(KEYINPUT56), .A2(n1029), .ZN(n1028) );
NOR3_X1 U741 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
XNOR2_X1 U742 ( .A(n1033), .B(KEYINPUT24), .ZN(n1031) );
XNOR2_X1 U743 ( .A(G107), .B(KEYINPUT51), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR4_X1 U745 ( .A1(G953), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR3_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NOR3_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1044) );
NOR2_X1 U750 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U751 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U752 ( .A1(n1053), .A2(n1054), .ZN(n1047) );
XNOR2_X1 U753 ( .A(n1055), .B(KEYINPUT10), .ZN(n1053) );
NOR2_X1 U754 ( .A1(n1056), .A2(n1030), .ZN(n1046) );
NOR3_X1 U755 ( .A1(n1050), .A2(n1057), .A3(n1030), .ZN(n1041) );
NOR2_X1 U756 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U757 ( .A1(n1060), .A2(n1045), .ZN(n1059) );
NOR2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
XNOR2_X1 U759 ( .A(n1063), .B(KEYINPUT28), .ZN(n1062) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NOR2_X1 U761 ( .A1(n1066), .A2(n1043), .ZN(n1058) );
NOR2_X1 U762 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
AND2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR3_X1 U764 ( .A1(n1036), .A2(G953), .A3(G952), .ZN(n1034) );
AND4_X1 U765 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1036) );
NOR4_X1 U766 ( .A1(n1075), .A2(n1070), .A3(n1076), .A4(n1077), .ZN(n1074) );
AND2_X1 U767 ( .A1(n1078), .A2(G478), .ZN(n1077) );
NOR2_X1 U768 ( .A1(n1079), .A2(n1030), .ZN(n1073) );
XNOR2_X1 U769 ( .A(n1080), .B(n1081), .ZN(n1079) );
NOR2_X1 U770 ( .A1(G475), .A2(KEYINPUT22), .ZN(n1081) );
XNOR2_X1 U771 ( .A(n1082), .B(n1083), .ZN(n1072) );
NAND2_X1 U772 ( .A1(KEYINPUT35), .A2(G469), .ZN(n1082) );
XOR2_X1 U773 ( .A(n1084), .B(n1085), .Z(n1071) );
NAND3_X1 U774 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(G72) );
OR2_X1 U775 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(n1087) );
INV_X1 U777 ( .A(KEYINPUT42), .ZN(n1092) );
NAND2_X1 U778 ( .A1(n1093), .A2(n1090), .ZN(n1091) );
XNOR2_X1 U779 ( .A(KEYINPUT46), .B(n1089), .ZN(n1093) );
NAND2_X1 U780 ( .A1(KEYINPUT42), .A2(n1094), .ZN(n1086) );
NAND2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
OR2_X1 U782 ( .A1(n1089), .A2(KEYINPUT46), .ZN(n1096) );
NAND3_X1 U783 ( .A1(n1090), .A2(n1089), .A3(KEYINPUT46), .ZN(n1095) );
NAND2_X1 U784 ( .A1(G953), .A2(n1097), .ZN(n1089) );
NAND2_X1 U785 ( .A1(G900), .A2(G227), .ZN(n1097) );
NAND2_X1 U786 ( .A1(n1098), .A2(n1099), .ZN(n1090) );
NAND3_X1 U787 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
NAND2_X1 U788 ( .A1(G953), .A2(n1103), .ZN(n1101) );
OR2_X1 U789 ( .A1(n1100), .A2(n1102), .ZN(n1098) );
NAND2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(n1100) );
XNOR2_X1 U793 ( .A(n1110), .B(n1111), .ZN(n1109) );
XNOR2_X1 U794 ( .A(n1112), .B(G137), .ZN(n1111) );
XOR2_X1 U795 ( .A(n1113), .B(n1114), .Z(n1108) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1113) );
NOR2_X1 U797 ( .A1(KEYINPUT5), .A2(G125), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1117), .A2(n1118), .ZN(G69) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U800 ( .A(KEYINPUT47), .B(n1121), .Z(n1117) );
NOR2_X1 U801 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XNOR2_X1 U802 ( .A(KEYINPUT52), .B(n1119), .ZN(n1123) );
NAND2_X1 U803 ( .A1(n1124), .A2(n1125), .ZN(n1119) );
OR2_X1 U804 ( .A1(n1104), .A2(G224), .ZN(n1125) );
NOR2_X1 U805 ( .A1(n1126), .A2(n1127), .ZN(n1122) );
INV_X1 U806 ( .A(n1120), .ZN(n1127) );
NAND2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(n1120) );
NOR2_X1 U808 ( .A1(n1129), .A2(n1128), .ZN(n1126) );
AND2_X1 U809 ( .A1(n1130), .A2(n1124), .ZN(n1128) );
INV_X1 U810 ( .A(n1131), .ZN(n1124) );
XOR2_X1 U811 ( .A(KEYINPUT54), .B(n1132), .Z(n1130) );
NOR2_X1 U812 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U813 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1139), .ZN(G63) );
XNOR2_X1 U816 ( .A(n1140), .B(n1141), .ZN(n1139) );
AND2_X1 U817 ( .A1(G478), .A2(n1142), .ZN(n1141) );
NOR2_X1 U818 ( .A1(n1133), .A2(n1143), .ZN(G60) );
NOR3_X1 U819 ( .A1(n1080), .A2(n1144), .A3(n1145), .ZN(n1143) );
AND3_X1 U820 ( .A1(n1146), .A2(G475), .A3(n1142), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1147), .A2(n1146), .ZN(n1144) );
AND2_X1 U822 ( .A1(n1038), .A2(G475), .ZN(n1147) );
XOR2_X1 U823 ( .A(n1148), .B(n1149), .Z(G6) );
XNOR2_X1 U824 ( .A(G104), .B(KEYINPUT14), .ZN(n1148) );
NOR2_X1 U825 ( .A1(n1133), .A2(n1150), .ZN(G57) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U827 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U829 ( .A1(KEYINPUT60), .A2(n1157), .ZN(n1156) );
AND2_X1 U830 ( .A1(G472), .A2(n1142), .ZN(n1155) );
NOR2_X1 U831 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
NOR3_X1 U832 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1159) );
INV_X1 U833 ( .A(KEYINPUT40), .ZN(n1160) );
NOR2_X1 U834 ( .A1(KEYINPUT40), .A2(n1163), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1151) );
XNOR2_X1 U836 ( .A(G101), .B(KEYINPUT19), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(G54) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1167) );
XNOR2_X1 U839 ( .A(n1170), .B(n1171), .ZN(n1169) );
XNOR2_X1 U840 ( .A(n1172), .B(n1173), .ZN(n1168) );
NAND3_X1 U841 ( .A1(n1142), .A2(G469), .A3(KEYINPUT43), .ZN(n1172) );
INV_X1 U842 ( .A(n1138), .ZN(n1142) );
XNOR2_X1 U843 ( .A(n1133), .B(KEYINPUT31), .ZN(n1166) );
NOR2_X1 U844 ( .A1(n1133), .A2(n1174), .ZN(G51) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U846 ( .A(n1177), .B(n1178), .ZN(n1176) );
NOR3_X1 U847 ( .A1(n1138), .A2(KEYINPUT38), .A3(n1085), .ZN(n1178) );
NAND2_X1 U848 ( .A1(G902), .A2(n1038), .ZN(n1138) );
NAND3_X1 U849 ( .A1(n1129), .A2(n1106), .A3(n1179), .ZN(n1038) );
XNOR2_X1 U850 ( .A(n1107), .B(KEYINPUT39), .ZN(n1179) );
AND4_X1 U851 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1107) );
NAND3_X1 U852 ( .A1(n1033), .A2(n1184), .A3(n1185), .ZN(n1181) );
NAND2_X1 U853 ( .A1(n1186), .A2(n1187), .ZN(n1184) );
NAND3_X1 U854 ( .A1(n1063), .A2(n1188), .A3(KEYINPUT53), .ZN(n1187) );
NAND2_X1 U855 ( .A1(n1189), .A2(n1052), .ZN(n1186) );
OR2_X1 U856 ( .A1(n1190), .A2(KEYINPUT53), .ZN(n1180) );
AND4_X1 U857 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1106) );
AND4_X1 U858 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1129) );
NOR4_X1 U859 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1149), .ZN(n1198) );
NOR3_X1 U860 ( .A1(n1030), .A2(n1032), .A3(n1054), .ZN(n1149) );
NOR2_X1 U861 ( .A1(n1202), .A2(n1203), .ZN(n1197) );
NOR3_X1 U862 ( .A1(n1030), .A2(n1056), .A3(n1032), .ZN(n1203) );
INV_X1 U863 ( .A(n1055), .ZN(n1030) );
NAND4_X1 U864 ( .A1(n1204), .A2(n1052), .A3(n1205), .A4(n1206), .ZN(n1196) );
OR2_X1 U865 ( .A1(n1207), .A2(KEYINPUT27), .ZN(n1206) );
NAND2_X1 U866 ( .A1(KEYINPUT27), .A2(n1208), .ZN(n1205) );
NAND2_X1 U867 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
INV_X1 U868 ( .A(n1068), .ZN(n1210) );
NOR2_X1 U869 ( .A1(n1104), .A2(G952), .ZN(n1133) );
XNOR2_X1 U870 ( .A(G146), .B(n1191), .ZN(G48) );
NAND2_X1 U871 ( .A1(n1211), .A2(n1212), .ZN(n1191) );
NAND2_X1 U872 ( .A1(n1213), .A2(n1214), .ZN(G45) );
NAND2_X1 U873 ( .A1(G143), .A2(n1192), .ZN(n1214) );
XOR2_X1 U874 ( .A(KEYINPUT13), .B(n1215), .Z(n1213) );
NOR2_X1 U875 ( .A1(G143), .A2(n1192), .ZN(n1215) );
NAND4_X1 U876 ( .A1(n1216), .A2(n1063), .A3(n1217), .A4(n1218), .ZN(n1192) );
XNOR2_X1 U877 ( .A(G140), .B(n1193), .ZN(G42) );
NAND4_X1 U878 ( .A1(n1185), .A2(n1189), .A3(n1051), .A4(n1212), .ZN(n1193) );
XNOR2_X1 U879 ( .A(G137), .B(n1194), .ZN(G39) );
NAND4_X1 U880 ( .A1(n1185), .A2(n1189), .A3(n1204), .A4(n1219), .ZN(n1194) );
XOR2_X1 U881 ( .A(G134), .B(n1220), .Z(G36) );
NOR2_X1 U882 ( .A1(n1221), .A2(n1043), .ZN(n1220) );
INV_X1 U883 ( .A(n1189), .ZN(n1043) );
XOR2_X1 U884 ( .A(n1222), .B(KEYINPUT21), .Z(n1221) );
NAND2_X1 U885 ( .A1(n1216), .A2(n1033), .ZN(n1222) );
NAND2_X1 U886 ( .A1(n1223), .A2(n1224), .ZN(G33) );
NAND2_X1 U887 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
INV_X1 U888 ( .A(G131), .ZN(n1226) );
XNOR2_X1 U889 ( .A(KEYINPUT59), .B(n1182), .ZN(n1225) );
NAND2_X1 U890 ( .A1(n1227), .A2(G131), .ZN(n1223) );
XNOR2_X1 U891 ( .A(KEYINPUT4), .B(n1182), .ZN(n1227) );
NAND3_X1 U892 ( .A1(n1189), .A2(n1212), .A3(n1216), .ZN(n1182) );
AND2_X1 U893 ( .A1(n1185), .A2(n1052), .ZN(n1216) );
NOR2_X1 U894 ( .A1(n1064), .A2(n1076), .ZN(n1189) );
INV_X1 U895 ( .A(n1065), .ZN(n1076) );
XNOR2_X1 U896 ( .A(G128), .B(n1190), .ZN(G30) );
NAND2_X1 U897 ( .A1(n1211), .A2(n1033), .ZN(n1190) );
AND3_X1 U898 ( .A1(n1219), .A2(n1063), .A3(n1185), .ZN(n1211) );
AND2_X1 U899 ( .A1(n1068), .A2(n1228), .ZN(n1185) );
NAND2_X1 U900 ( .A1(n1040), .A2(n1229), .ZN(n1228) );
XOR2_X1 U901 ( .A(n1230), .B(n1231), .Z(G3) );
XNOR2_X1 U902 ( .A(KEYINPUT6), .B(n1232), .ZN(n1231) );
NAND4_X1 U903 ( .A1(KEYINPUT18), .A2(n1204), .A3(n1052), .A4(n1207), .ZN(n1230) );
XNOR2_X1 U904 ( .A(G125), .B(n1183), .ZN(G27) );
NAND4_X1 U905 ( .A1(n1051), .A2(n1212), .A3(n1233), .A4(n1234), .ZN(n1183) );
NOR2_X1 U906 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
AND2_X1 U907 ( .A1(n1040), .A2(n1229), .ZN(n1235) );
NAND4_X1 U908 ( .A1(G953), .A2(n1237), .A3(n1238), .A4(n1103), .ZN(n1229) );
INV_X1 U909 ( .A(G900), .ZN(n1103) );
XNOR2_X1 U910 ( .A(KEYINPUT30), .B(n1239), .ZN(n1237) );
XNOR2_X1 U911 ( .A(n1201), .B(n1240), .ZN(G24) );
NAND2_X1 U912 ( .A1(KEYINPUT49), .A2(G122), .ZN(n1240) );
AND4_X1 U913 ( .A1(n1241), .A2(n1055), .A3(n1217), .A4(n1218), .ZN(n1201) );
NOR2_X1 U914 ( .A1(n1242), .A2(n1243), .ZN(n1055) );
XOR2_X1 U915 ( .A(G119), .B(n1200), .Z(G21) );
AND3_X1 U916 ( .A1(n1219), .A2(n1241), .A3(n1204), .ZN(n1200) );
INV_X1 U917 ( .A(n1188), .ZN(n1219) );
NAND2_X1 U918 ( .A1(n1243), .A2(n1242), .ZN(n1188) );
NAND2_X1 U919 ( .A1(n1244), .A2(n1245), .ZN(G18) );
NAND2_X1 U920 ( .A1(n1199), .A2(n1246), .ZN(n1245) );
XOR2_X1 U921 ( .A(KEYINPUT9), .B(n1247), .Z(n1244) );
NOR2_X1 U922 ( .A1(n1199), .A2(n1246), .ZN(n1247) );
AND3_X1 U923 ( .A1(n1241), .A2(n1033), .A3(n1052), .ZN(n1199) );
INV_X1 U924 ( .A(n1056), .ZN(n1033) );
NAND2_X1 U925 ( .A1(n1248), .A2(n1218), .ZN(n1056) );
AND3_X1 U926 ( .A1(n1063), .A2(n1249), .A3(n1234), .ZN(n1241) );
INV_X1 U927 ( .A(n1236), .ZN(n1063) );
XOR2_X1 U928 ( .A(G113), .B(n1202), .Z(G15) );
AND4_X1 U929 ( .A1(n1212), .A2(n1052), .A3(n1234), .A4(n1209), .ZN(n1202) );
INV_X1 U930 ( .A(n1045), .ZN(n1234) );
NAND2_X1 U931 ( .A1(n1069), .A2(n1250), .ZN(n1045) );
AND2_X1 U932 ( .A1(n1251), .A2(n1242), .ZN(n1052) );
INV_X1 U933 ( .A(n1054), .ZN(n1212) );
NAND2_X1 U934 ( .A1(n1252), .A2(n1217), .ZN(n1054) );
INV_X1 U935 ( .A(n1248), .ZN(n1217) );
XNOR2_X1 U936 ( .A(G110), .B(n1195), .ZN(G12) );
NAND3_X1 U937 ( .A1(n1204), .A2(n1207), .A3(n1051), .ZN(n1195) );
NOR2_X1 U938 ( .A1(n1242), .A2(n1251), .ZN(n1051) );
INV_X1 U939 ( .A(n1243), .ZN(n1251) );
XOR2_X1 U940 ( .A(n1253), .B(n1137), .Z(n1243) );
NAND2_X1 U941 ( .A1(G217), .A2(n1254), .ZN(n1137) );
OR2_X1 U942 ( .A1(n1136), .A2(G902), .ZN(n1253) );
XNOR2_X1 U943 ( .A(n1255), .B(n1256), .ZN(n1136) );
XOR2_X1 U944 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U945 ( .A(n1110), .B(G119), .ZN(n1258) );
XOR2_X1 U946 ( .A(KEYINPUT34), .B(G146), .Z(n1257) );
XOR2_X1 U947 ( .A(n1259), .B(n1260), .Z(n1255) );
XOR2_X1 U948 ( .A(n1261), .B(n1262), .Z(n1260) );
NAND2_X1 U949 ( .A1(G221), .A2(n1263), .ZN(n1262) );
NAND2_X1 U950 ( .A1(KEYINPUT36), .A2(n1264), .ZN(n1261) );
XNOR2_X1 U951 ( .A(n1265), .B(n1266), .ZN(n1259) );
NAND3_X1 U952 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1265) );
NAND2_X1 U953 ( .A1(KEYINPUT12), .A2(G140), .ZN(n1269) );
NAND3_X1 U954 ( .A1(n1112), .A2(n1270), .A3(G125), .ZN(n1268) );
NAND2_X1 U955 ( .A1(n1271), .A2(n1177), .ZN(n1267) );
NAND2_X1 U956 ( .A1(n1272), .A2(n1270), .ZN(n1271) );
INV_X1 U957 ( .A(KEYINPUT12), .ZN(n1270) );
XNOR2_X1 U958 ( .A(G140), .B(KEYINPUT61), .ZN(n1272) );
XNOR2_X1 U959 ( .A(n1273), .B(G472), .ZN(n1242) );
NAND2_X1 U960 ( .A1(n1274), .A2(n1239), .ZN(n1273) );
XOR2_X1 U961 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U962 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U963 ( .A(KEYINPUT0), .B(n1232), .ZN(n1278) );
NOR2_X1 U964 ( .A1(KEYINPUT57), .A2(n1164), .ZN(n1277) );
NAND3_X1 U965 ( .A1(n1279), .A2(n1104), .A3(G210), .ZN(n1164) );
XNOR2_X1 U966 ( .A(KEYINPUT37), .B(n1280), .ZN(n1279) );
XOR2_X1 U967 ( .A(n1163), .B(n1157), .Z(n1275) );
XNOR2_X1 U968 ( .A(n1281), .B(KEYINPUT20), .ZN(n1157) );
XNOR2_X1 U969 ( .A(n1161), .B(n1162), .ZN(n1163) );
INV_X1 U970 ( .A(n1032), .ZN(n1207) );
NAND2_X1 U971 ( .A1(n1068), .A2(n1209), .ZN(n1032) );
AND2_X1 U972 ( .A1(n1282), .A2(n1249), .ZN(n1209) );
NAND2_X1 U973 ( .A1(n1040), .A2(n1283), .ZN(n1249) );
NAND3_X1 U974 ( .A1(n1131), .A2(n1238), .A3(G902), .ZN(n1283) );
NOR2_X1 U975 ( .A1(G898), .A2(n1104), .ZN(n1131) );
NAND3_X1 U976 ( .A1(n1238), .A2(n1104), .A3(G952), .ZN(n1040) );
NAND2_X1 U977 ( .A1(G234), .A2(G237), .ZN(n1238) );
XNOR2_X1 U978 ( .A(KEYINPUT25), .B(n1236), .ZN(n1282) );
NAND2_X1 U979 ( .A1(n1064), .A2(n1065), .ZN(n1236) );
NAND2_X1 U980 ( .A1(G214), .A2(n1284), .ZN(n1065) );
XOR2_X1 U981 ( .A(n1085), .B(n1285), .Z(n1064) );
NOR2_X1 U982 ( .A1(n1084), .A2(KEYINPUT3), .ZN(n1285) );
AND2_X1 U983 ( .A1(n1286), .A2(n1239), .ZN(n1084) );
XOR2_X1 U984 ( .A(n1175), .B(n1287), .Z(n1286) );
NOR2_X1 U985 ( .A1(G125), .A2(KEYINPUT11), .ZN(n1287) );
XOR2_X1 U986 ( .A(n1288), .B(n1289), .Z(n1175) );
XOR2_X1 U987 ( .A(n1290), .B(n1162), .Z(n1289) );
XOR2_X1 U988 ( .A(n1291), .B(n1292), .Z(n1162) );
XNOR2_X1 U989 ( .A(G143), .B(n1110), .ZN(n1292) );
INV_X1 U990 ( .A(G128), .ZN(n1110) );
NAND2_X1 U991 ( .A1(KEYINPUT50), .A2(G146), .ZN(n1291) );
NAND2_X1 U992 ( .A1(G224), .A2(n1104), .ZN(n1290) );
NAND2_X1 U993 ( .A1(n1293), .A2(n1294), .ZN(n1288) );
NAND2_X1 U994 ( .A1(n1132), .A2(n1295), .ZN(n1294) );
INV_X1 U995 ( .A(KEYINPUT2), .ZN(n1295) );
XNOR2_X1 U996 ( .A(n1296), .B(n1297), .ZN(n1132) );
XOR2_X1 U997 ( .A(n1298), .B(n1281), .Z(n1297) );
NAND2_X1 U998 ( .A1(KEYINPUT2), .A2(n1299), .ZN(n1293) );
XOR2_X1 U999 ( .A(n1300), .B(n1298), .Z(n1299) );
XNOR2_X1 U1000 ( .A(n1266), .B(n1301), .ZN(n1298) );
INV_X1 U1001 ( .A(G110), .ZN(n1266) );
NAND2_X1 U1002 ( .A1(n1296), .A2(n1281), .ZN(n1300) );
XOR2_X1 U1003 ( .A(G113), .B(n1302), .Z(n1281) );
XNOR2_X1 U1004 ( .A(G119), .B(n1246), .ZN(n1302) );
XNOR2_X1 U1005 ( .A(n1303), .B(n1232), .ZN(n1296) );
NAND2_X1 U1006 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U1007 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1008 ( .A(KEYINPUT58), .B(n1308), .Z(n1304) );
NOR2_X1 U1009 ( .A1(n1306), .A2(n1307), .ZN(n1308) );
XOR2_X1 U1010 ( .A(KEYINPUT62), .B(G107), .Z(n1307) );
NAND2_X1 U1011 ( .A1(G210), .A2(n1284), .ZN(n1085) );
NAND2_X1 U1012 ( .A1(n1280), .A2(n1239), .ZN(n1284) );
INV_X1 U1013 ( .A(G237), .ZN(n1280) );
NOR2_X1 U1014 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
INV_X1 U1015 ( .A(n1250), .ZN(n1070) );
NAND2_X1 U1016 ( .A1(G221), .A2(n1254), .ZN(n1250) );
NAND2_X1 U1017 ( .A1(G234), .A2(n1239), .ZN(n1254) );
XNOR2_X1 U1018 ( .A(n1083), .B(n1309), .ZN(n1069) );
XOR2_X1 U1019 ( .A(KEYINPUT44), .B(G469), .Z(n1309) );
NAND2_X1 U1020 ( .A1(n1310), .A2(n1239), .ZN(n1083) );
XNOR2_X1 U1021 ( .A(n1311), .B(n1312), .ZN(n1310) );
INV_X1 U1022 ( .A(n1173), .ZN(n1312) );
XNOR2_X1 U1023 ( .A(n1313), .B(n1314), .ZN(n1173) );
XOR2_X1 U1024 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1025 ( .A(n1115), .B(KEYINPUT45), .Z(n1316) );
NAND2_X1 U1026 ( .A1(KEYINPUT23), .A2(n1317), .ZN(n1115) );
NAND2_X1 U1027 ( .A1(KEYINPUT15), .A2(n1232), .ZN(n1315) );
INV_X1 U1028 ( .A(G101), .ZN(n1232) );
XNOR2_X1 U1029 ( .A(n1318), .B(n1306), .ZN(n1313) );
XNOR2_X1 U1030 ( .A(G104), .B(KEYINPUT29), .ZN(n1306) );
XOR2_X1 U1031 ( .A(n1319), .B(n1320), .Z(n1318) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1104), .ZN(n1319) );
XNOR2_X1 U1033 ( .A(n1321), .B(n1322), .ZN(n1311) );
NOR2_X1 U1034 ( .A1(KEYINPUT32), .A2(n1161), .ZN(n1322) );
INV_X1 U1035 ( .A(n1171), .ZN(n1161) );
NAND2_X1 U1036 ( .A1(n1323), .A2(n1324), .ZN(n1171) );
NAND2_X1 U1037 ( .A1(n1114), .A2(n1264), .ZN(n1324) );
INV_X1 U1038 ( .A(G137), .ZN(n1264) );
NAND2_X1 U1039 ( .A1(n1325), .A2(G137), .ZN(n1323) );
XOR2_X1 U1040 ( .A(KEYINPUT26), .B(n1114), .Z(n1325) );
XOR2_X1 U1041 ( .A(G134), .B(G131), .Z(n1114) );
NOR2_X1 U1042 ( .A1(KEYINPUT1), .A2(n1170), .ZN(n1321) );
XNOR2_X1 U1043 ( .A(G110), .B(n1112), .ZN(n1170) );
INV_X1 U1044 ( .A(n1050), .ZN(n1204) );
NAND2_X1 U1045 ( .A1(n1252), .A2(n1248), .ZN(n1050) );
XNOR2_X1 U1046 ( .A(n1080), .B(G475), .ZN(n1248) );
NOR2_X1 U1047 ( .A1(n1146), .A2(G902), .ZN(n1080) );
XNOR2_X1 U1048 ( .A(n1326), .B(n1327), .ZN(n1146) );
XNOR2_X1 U1049 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U1050 ( .A1(G104), .A2(KEYINPUT33), .ZN(n1329) );
NAND2_X1 U1051 ( .A1(KEYINPUT48), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1052 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1053 ( .A(n1317), .B(n1333), .ZN(n1332) );
XNOR2_X1 U1054 ( .A(n1177), .B(n1334), .ZN(n1333) );
NOR4_X1 U1055 ( .A1(KEYINPUT41), .A2(G953), .A3(G237), .A4(n1335), .ZN(n1334) );
INV_X1 U1056 ( .A(G214), .ZN(n1335) );
INV_X1 U1057 ( .A(G125), .ZN(n1177) );
XNOR2_X1 U1058 ( .A(G143), .B(G146), .ZN(n1317) );
XOR2_X1 U1059 ( .A(n1336), .B(n1337), .Z(n1331) );
XNOR2_X1 U1060 ( .A(n1112), .B(G131), .ZN(n1337) );
INV_X1 U1061 ( .A(G140), .ZN(n1112) );
XOR2_X1 U1062 ( .A(KEYINPUT63), .B(KEYINPUT17), .Z(n1336) );
XNOR2_X1 U1063 ( .A(G113), .B(n1338), .ZN(n1326) );
NOR2_X1 U1064 ( .A1(KEYINPUT7), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1065 ( .A(n1218), .B(KEYINPUT16), .Z(n1252) );
NAND2_X1 U1066 ( .A1(n1340), .A2(n1341), .ZN(n1218) );
NAND2_X1 U1067 ( .A1(G478), .A2(n1078), .ZN(n1341) );
XOR2_X1 U1068 ( .A(KEYINPUT55), .B(n1075), .Z(n1340) );
NOR2_X1 U1069 ( .A1(n1078), .A2(G478), .ZN(n1075) );
NAND2_X1 U1070 ( .A1(n1140), .A2(n1239), .ZN(n1078) );
INV_X1 U1071 ( .A(G902), .ZN(n1239) );
XNOR2_X1 U1072 ( .A(n1342), .B(n1343), .ZN(n1140) );
XNOR2_X1 U1073 ( .A(n1246), .B(n1344), .ZN(n1343) );
XOR2_X1 U1074 ( .A(G143), .B(G134), .Z(n1344) );
INV_X1 U1075 ( .A(G116), .ZN(n1246) );
XNOR2_X1 U1076 ( .A(n1345), .B(n1339), .ZN(n1342) );
INV_X1 U1077 ( .A(n1301), .ZN(n1339) );
XOR2_X1 U1078 ( .A(G122), .B(KEYINPUT8), .Z(n1301) );
XOR2_X1 U1079 ( .A(n1346), .B(n1320), .Z(n1345) );
XOR2_X1 U1080 ( .A(G107), .B(G128), .Z(n1320) );
NAND2_X1 U1081 ( .A1(n1263), .A2(G217), .ZN(n1346) );
AND2_X1 U1082 ( .A1(G234), .A2(n1104), .ZN(n1263) );
INV_X1 U1083 ( .A(G953), .ZN(n1104) );
endmodule


