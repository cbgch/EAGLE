//Key = 1101110011111000101001101110111010100010000001011110111001101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291;

XOR2_X1 U706 ( .A(n985), .B(n986), .Z(G9) );
XOR2_X1 U707 ( .A(KEYINPUT63), .B(G107), .Z(n986) );
NAND3_X1 U708 ( .A1(n987), .A2(n988), .A3(n989), .ZN(G75) );
NAND2_X1 U709 ( .A1(G952), .A2(n990), .ZN(n989) );
NAND3_X1 U710 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n990) );
NAND2_X1 U711 ( .A1(n994), .A2(n995), .ZN(n992) );
NAND2_X1 U712 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND3_X1 U713 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
NAND2_X1 U714 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NAND2_X1 U715 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U716 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U717 ( .A1(n1007), .A2(n1008), .ZN(n1001) );
NAND2_X1 U718 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U719 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND3_X1 U720 ( .A1(n1007), .A2(n1013), .A3(n1003), .ZN(n996) );
NAND2_X1 U721 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U722 ( .A1(n998), .A2(n1016), .ZN(n1015) );
NAND2_X1 U723 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U724 ( .A1(n1000), .A2(n1019), .ZN(n1014) );
NAND2_X1 U725 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U726 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
XNOR2_X1 U727 ( .A(KEYINPUT29), .B(n1024), .ZN(n994) );
NAND4_X1 U728 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n987) );
NOR4_X1 U729 ( .A1(n1011), .A2(n1022), .A3(n1029), .A4(n1030), .ZN(n1028) );
XOR2_X1 U730 ( .A(n1031), .B(n1032), .Z(n1030) );
NOR2_X1 U731 ( .A1(G472), .A2(n1033), .ZN(n1032) );
XOR2_X1 U732 ( .A(KEYINPUT2), .B(KEYINPUT19), .Z(n1033) );
XOR2_X1 U733 ( .A(n1034), .B(n1035), .Z(n1029) );
NOR2_X1 U734 ( .A1(n1036), .A2(KEYINPUT41), .ZN(n1035) );
NOR2_X1 U735 ( .A1(n1037), .A2(n1038), .ZN(n1027) );
XOR2_X1 U736 ( .A(G469), .B(n1039), .Z(n1038) );
NOR2_X1 U737 ( .A1(KEYINPUT14), .A2(n1040), .ZN(n1039) );
XOR2_X1 U738 ( .A(n1023), .B(KEYINPUT34), .Z(n1037) );
XOR2_X1 U739 ( .A(n1041), .B(n1042), .Z(n1026) );
XOR2_X1 U740 ( .A(n1043), .B(n1044), .Z(n1025) );
XOR2_X1 U741 ( .A(n1045), .B(n1046), .Z(G72) );
XOR2_X1 U742 ( .A(n1047), .B(n1048), .Z(n1046) );
NAND2_X1 U743 ( .A1(G953), .A2(n1049), .ZN(n1048) );
NAND2_X1 U744 ( .A1(G900), .A2(G227), .ZN(n1049) );
NAND3_X1 U745 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1047) );
NAND2_X1 U746 ( .A1(G953), .A2(n1053), .ZN(n1052) );
NAND2_X1 U747 ( .A1(n1054), .A2(n1055), .ZN(n1051) );
NAND2_X1 U748 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XOR2_X1 U749 ( .A(G140), .B(n1058), .Z(n1054) );
NAND3_X1 U750 ( .A1(n1056), .A2(n1057), .A3(n1059), .ZN(n1050) );
XOR2_X1 U751 ( .A(n1060), .B(n1058), .Z(n1059) );
NOR2_X1 U752 ( .A1(KEYINPUT59), .A2(n1061), .ZN(n1058) );
NAND2_X1 U753 ( .A1(n1062), .A2(n1063), .ZN(n1057) );
XOR2_X1 U754 ( .A(KEYINPUT56), .B(n1064), .Z(n1062) );
XNOR2_X1 U755 ( .A(KEYINPUT9), .B(n1065), .ZN(n1056) );
NAND2_X1 U756 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XOR2_X1 U757 ( .A(KEYINPUT11), .B(n1063), .Z(n1067) );
XNOR2_X1 U758 ( .A(n1064), .B(KEYINPUT56), .ZN(n1066) );
NOR2_X1 U759 ( .A1(n993), .A2(G953), .ZN(n1045) );
XOR2_X1 U760 ( .A(n1068), .B(n1069), .Z(G69) );
XOR2_X1 U761 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U762 ( .A1(n991), .A2(G953), .ZN(n1071) );
NOR2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
XNOR2_X1 U764 ( .A(n1074), .B(n1075), .ZN(n1073) );
XOR2_X1 U765 ( .A(n1076), .B(KEYINPUT15), .Z(n1075) );
NOR2_X1 U766 ( .A1(G898), .A2(n988), .ZN(n1072) );
NOR2_X1 U767 ( .A1(n1077), .A2(n988), .ZN(n1068) );
AND2_X1 U768 ( .A1(G224), .A2(G898), .ZN(n1077) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(G66) );
XOR2_X1 U770 ( .A(n1080), .B(n1081), .Z(n1079) );
XOR2_X1 U771 ( .A(KEYINPUT1), .B(n1082), .Z(n1081) );
NOR2_X1 U772 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U773 ( .A1(n1078), .A2(n1085), .ZN(G63) );
XOR2_X1 U774 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U775 ( .A1(n1044), .A2(n1084), .ZN(n1087) );
NOR2_X1 U776 ( .A1(n1078), .A2(n1088), .ZN(G60) );
XOR2_X1 U777 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U778 ( .A1(n1042), .A2(n1084), .ZN(n1089) );
INV_X1 U779 ( .A(G475), .ZN(n1042) );
NAND2_X1 U780 ( .A1(n1091), .A2(n1092), .ZN(G6) );
NAND3_X1 U781 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
XOR2_X1 U782 ( .A(KEYINPUT60), .B(G104), .Z(n1093) );
NAND2_X1 U783 ( .A1(n1096), .A2(n1097), .ZN(n1091) );
NAND2_X1 U784 ( .A1(n1095), .A2(n1094), .ZN(n1097) );
XOR2_X1 U785 ( .A(n1098), .B(KEYINPUT54), .Z(n1096) );
INV_X1 U786 ( .A(G104), .ZN(n1098) );
NOR2_X1 U787 ( .A1(n1078), .A2(n1099), .ZN(G57) );
XOR2_X1 U788 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U789 ( .A(KEYINPUT16), .B(n1102), .Z(n1101) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1084), .ZN(n1102) );
INV_X1 U791 ( .A(G472), .ZN(n1103) );
NOR2_X1 U792 ( .A1(n1078), .A2(n1104), .ZN(G54) );
XOR2_X1 U793 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XOR2_X1 U795 ( .A(n1109), .B(KEYINPUT49), .Z(n1108) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1110), .A2(n1112), .ZN(n1107) );
XOR2_X1 U798 ( .A(KEYINPUT35), .B(n1111), .Z(n1112) );
AND2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NAND2_X1 U800 ( .A1(n1115), .A2(G110), .ZN(n1114) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
XNOR2_X1 U802 ( .A(KEYINPUT36), .B(n1115), .ZN(n1116) );
XOR2_X1 U803 ( .A(n1118), .B(n1119), .Z(n1115) );
XOR2_X1 U804 ( .A(n1120), .B(n1121), .Z(n1110) );
NOR2_X1 U805 ( .A1(KEYINPUT17), .A2(n1122), .ZN(n1121) );
NOR2_X1 U806 ( .A1(n1084), .A2(n1123), .ZN(n1105) );
XOR2_X1 U807 ( .A(KEYINPUT45), .B(G469), .Z(n1123) );
NOR2_X1 U808 ( .A1(n1078), .A2(n1124), .ZN(G51) );
XOR2_X1 U809 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U811 ( .A(KEYINPUT44), .B(n1129), .Z(n1128) );
AND2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U813 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
XNOR2_X1 U814 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR2_X1 U815 ( .A1(n1084), .A2(n1134), .ZN(n1125) );
XOR2_X1 U816 ( .A(KEYINPUT24), .B(G210), .Z(n1134) );
NAND2_X1 U817 ( .A1(G902), .A2(n1135), .ZN(n1084) );
NAND2_X1 U818 ( .A1(n993), .A2(n991), .ZN(n1135) );
AND2_X1 U819 ( .A1(n1136), .A2(n1137), .ZN(n991) );
NOR4_X1 U820 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1137) );
NOR4_X1 U821 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
INV_X1 U822 ( .A(n1146), .ZN(n1144) );
NOR2_X1 U823 ( .A1(KEYINPUT28), .A2(n1147), .ZN(n1143) );
NOR2_X1 U824 ( .A1(n1020), .A2(n1148), .ZN(n1147) );
AND2_X1 U825 ( .A1(n1149), .A2(KEYINPUT28), .ZN(n1142) );
NOR4_X1 U826 ( .A1(n985), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1136) );
NOR3_X1 U827 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
NOR3_X1 U828 ( .A1(n1156), .A2(n1005), .A3(n1009), .ZN(n1151) );
NAND3_X1 U829 ( .A1(n1157), .A2(n1158), .A3(n1000), .ZN(n1156) );
INV_X1 U830 ( .A(n1154), .ZN(n1000) );
OR2_X1 U831 ( .A1(n1159), .A2(KEYINPUT51), .ZN(n1158) );
NAND2_X1 U832 ( .A1(KEYINPUT51), .A2(n1160), .ZN(n1157) );
NAND2_X1 U833 ( .A1(n1020), .A2(n1148), .ZN(n1160) );
NOR4_X1 U834 ( .A1(n1161), .A2(n1162), .A3(n1006), .A4(n1018), .ZN(n1150) );
NOR2_X1 U835 ( .A1(KEYINPUT48), .A2(n1163), .ZN(n1162) );
NOR2_X1 U836 ( .A1(n1003), .A2(n1149), .ZN(n1163) );
AND2_X1 U837 ( .A1(n1153), .A2(KEYINPUT48), .ZN(n1161) );
AND2_X1 U838 ( .A1(n1164), .A2(n1095), .ZN(n985) );
NOR3_X1 U839 ( .A1(n1009), .A2(n1149), .A3(n1154), .ZN(n1095) );
AND2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(n993) );
NOR4_X1 U841 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
AND4_X1 U842 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1165) );
NAND4_X1 U843 ( .A1(n1175), .A2(n1176), .A3(n1003), .A4(n1177), .ZN(n1173) );
XOR2_X1 U844 ( .A(KEYINPUT4), .B(n1017), .Z(n1177) );
NOR2_X1 U845 ( .A1(n988), .A2(G952), .ZN(n1078) );
NAND2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(G48) );
OR2_X1 U847 ( .A1(n1174), .A2(G146), .ZN(n1179) );
XOR2_X1 U848 ( .A(n1180), .B(KEYINPUT39), .Z(n1178) );
NAND2_X1 U849 ( .A1(G146), .A2(n1174), .ZN(n1180) );
NAND3_X1 U850 ( .A1(n1175), .A2(n1094), .A3(n1181), .ZN(n1174) );
XNOR2_X1 U851 ( .A(G143), .B(n1172), .ZN(G45) );
NAND4_X1 U852 ( .A1(n1146), .A2(n1182), .A3(n1175), .A4(n1183), .ZN(n1172) );
XOR2_X1 U853 ( .A(n1060), .B(n1171), .Z(G42) );
NAND4_X1 U854 ( .A1(n1184), .A2(n1176), .A3(n1185), .A4(n998), .ZN(n1171) );
XOR2_X1 U855 ( .A(G137), .B(n1170), .Z(G39) );
AND3_X1 U856 ( .A1(n1181), .A2(n998), .A3(n1007), .ZN(n1170) );
XOR2_X1 U857 ( .A(G134), .B(n1169), .Z(G36) );
AND4_X1 U858 ( .A1(n1146), .A2(n1164), .A3(n998), .A4(n1183), .ZN(n1169) );
XOR2_X1 U859 ( .A(G131), .B(n1168), .Z(G33) );
AND3_X1 U860 ( .A1(n1146), .A2(n998), .A3(n1176), .ZN(n1168) );
NAND2_X1 U861 ( .A1(n1186), .A2(n1187), .ZN(n998) );
OR2_X1 U862 ( .A1(n1020), .A2(KEYINPUT52), .ZN(n1187) );
NAND3_X1 U863 ( .A1(n1023), .A2(n1188), .A3(KEYINPUT52), .ZN(n1186) );
INV_X1 U864 ( .A(n1022), .ZN(n1188) );
XOR2_X1 U865 ( .A(G128), .B(n1167), .Z(G30) );
AND3_X1 U866 ( .A1(n1164), .A2(n1175), .A3(n1181), .ZN(n1167) );
NOR4_X1 U867 ( .A1(n1009), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1181) );
XNOR2_X1 U868 ( .A(G101), .B(n1192), .ZN(G3) );
NAND3_X1 U869 ( .A1(n1146), .A2(n1159), .A3(n1007), .ZN(n1192) );
INV_X1 U870 ( .A(n1145), .ZN(n1007) );
NOR2_X1 U871 ( .A1(n1018), .A2(n1009), .ZN(n1146) );
XOR2_X1 U872 ( .A(G125), .B(n1193), .Z(G27) );
NOR2_X1 U873 ( .A1(n1194), .A2(n1020), .ZN(n1193) );
INV_X1 U874 ( .A(n1175), .ZN(n1020) );
XOR2_X1 U875 ( .A(n1195), .B(KEYINPUT55), .Z(n1194) );
NAND3_X1 U876 ( .A1(n1184), .A2(n1176), .A3(n1003), .ZN(n1195) );
NOR2_X1 U877 ( .A1(n1005), .A2(n1191), .ZN(n1176) );
INV_X1 U878 ( .A(n1183), .ZN(n1191) );
NAND2_X1 U879 ( .A1(n1196), .A2(n1197), .ZN(n1183) );
NAND2_X1 U880 ( .A1(n1198), .A2(n1053), .ZN(n1197) );
INV_X1 U881 ( .A(G900), .ZN(n1053) );
XOR2_X1 U882 ( .A(G122), .B(n1199), .Z(G24) );
NOR4_X1 U883 ( .A1(KEYINPUT46), .A2(n1154), .A3(n1153), .A4(n1200), .ZN(n1199) );
XOR2_X1 U884 ( .A(KEYINPUT47), .B(n1182), .Z(n1200) );
NAND2_X1 U885 ( .A1(n1190), .A2(n1189), .ZN(n1154) );
XOR2_X1 U886 ( .A(G119), .B(n1140), .Z(G21) );
NOR4_X1 U887 ( .A1(n1153), .A2(n1145), .A3(n1189), .A4(n1190), .ZN(n1140) );
XOR2_X1 U888 ( .A(G116), .B(n1201), .Z(G18) );
NOR3_X1 U889 ( .A1(n1153), .A2(n1006), .A3(n1018), .ZN(n1201) );
INV_X1 U890 ( .A(n1164), .ZN(n1006) );
NOR2_X1 U891 ( .A1(n1202), .A2(n1203), .ZN(n1164) );
XOR2_X1 U892 ( .A(n1139), .B(n1204), .Z(G15) );
NOR2_X1 U893 ( .A1(KEYINPUT27), .A2(n1205), .ZN(n1204) );
NOR3_X1 U894 ( .A1(n1018), .A2(n1005), .A3(n1153), .ZN(n1139) );
NAND2_X1 U895 ( .A1(n1003), .A2(n1159), .ZN(n1153) );
INV_X1 U896 ( .A(n1149), .ZN(n1159) );
NOR2_X1 U897 ( .A1(n1206), .A2(n1011), .ZN(n1003) );
INV_X1 U898 ( .A(n1094), .ZN(n1005) );
NAND2_X1 U899 ( .A1(n1207), .A2(n1208), .ZN(n1094) );
OR2_X1 U900 ( .A1(n1155), .A2(KEYINPUT61), .ZN(n1208) );
INV_X1 U901 ( .A(n1182), .ZN(n1155) );
NOR2_X1 U902 ( .A1(n1202), .A2(n1209), .ZN(n1182) );
NAND3_X1 U903 ( .A1(n1203), .A2(n1202), .A3(KEYINPUT61), .ZN(n1207) );
INV_X1 U904 ( .A(n1209), .ZN(n1203) );
NAND2_X1 U905 ( .A1(n1189), .A2(n1210), .ZN(n1018) );
XOR2_X1 U906 ( .A(G110), .B(n1138), .Z(G12) );
NOR4_X1 U907 ( .A1(n1017), .A2(n1145), .A3(n1009), .A4(n1149), .ZN(n1138) );
NAND2_X1 U908 ( .A1(n1175), .A2(n1148), .ZN(n1149) );
NAND2_X1 U909 ( .A1(n1196), .A2(n1211), .ZN(n1148) );
NAND2_X1 U910 ( .A1(n1198), .A2(n1212), .ZN(n1211) );
INV_X1 U911 ( .A(G898), .ZN(n1212) );
AND3_X1 U912 ( .A1(G902), .A2(n1024), .A3(G953), .ZN(n1198) );
NAND3_X1 U913 ( .A1(n1024), .A2(n988), .A3(G952), .ZN(n1196) );
NAND2_X1 U914 ( .A1(n1213), .A2(G237), .ZN(n1024) );
XOR2_X1 U915 ( .A(n1214), .B(KEYINPUT25), .Z(n1213) );
NOR2_X1 U916 ( .A1(n1023), .A2(n1022), .ZN(n1175) );
NOR2_X1 U917 ( .A1(n1215), .A2(n1216), .ZN(n1022) );
XOR2_X1 U918 ( .A(G214), .B(KEYINPUT22), .Z(n1215) );
XOR2_X1 U919 ( .A(n1217), .B(n1218), .Z(n1023) );
NOR2_X1 U920 ( .A1(n1216), .A2(n1219), .ZN(n1218) );
NOR2_X1 U921 ( .A1(G902), .A2(G237), .ZN(n1216) );
NAND2_X1 U922 ( .A1(n1220), .A2(n1221), .ZN(n1217) );
XOR2_X1 U923 ( .A(n1222), .B(n1223), .Z(n1220) );
NOR2_X1 U924 ( .A1(KEYINPUT42), .A2(n1130), .ZN(n1223) );
XNOR2_X1 U925 ( .A(n1076), .B(n1224), .ZN(n1130) );
NOR2_X1 U926 ( .A1(KEYINPUT13), .A2(n1074), .ZN(n1224) );
XNOR2_X1 U927 ( .A(n1225), .B(G122), .ZN(n1074) );
NAND2_X1 U928 ( .A1(KEYINPUT12), .A2(G110), .ZN(n1225) );
XOR2_X1 U929 ( .A(n1226), .B(n1227), .Z(n1076) );
XOR2_X1 U930 ( .A(n1132), .B(n1228), .Z(n1222) );
NOR2_X1 U931 ( .A1(KEYINPUT6), .A2(n1133), .ZN(n1228) );
XOR2_X1 U932 ( .A(G125), .B(n1063), .Z(n1133) );
NAND2_X1 U933 ( .A1(G224), .A2(n988), .ZN(n1132) );
INV_X1 U934 ( .A(n1185), .ZN(n1009) );
NOR2_X1 U935 ( .A1(n1012), .A2(n1011), .ZN(n1185) );
NOR2_X1 U936 ( .A1(n1229), .A2(n1230), .ZN(n1011) );
INV_X1 U937 ( .A(n1206), .ZN(n1012) );
XNOR2_X1 U938 ( .A(n1040), .B(G469), .ZN(n1206) );
NAND2_X1 U939 ( .A1(n1231), .A2(n1221), .ZN(n1040) );
XOR2_X1 U940 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U941 ( .A(n1118), .B(n1234), .ZN(n1233) );
XOR2_X1 U942 ( .A(KEYINPUT40), .B(G110), .Z(n1234) );
NAND2_X1 U943 ( .A1(G227), .A2(n988), .ZN(n1118) );
XOR2_X1 U944 ( .A(n1235), .B(n1119), .Z(n1232) );
XOR2_X1 U945 ( .A(G140), .B(KEYINPUT23), .Z(n1119) );
XNOR2_X1 U946 ( .A(n1120), .B(n1122), .ZN(n1235) );
XOR2_X1 U947 ( .A(n1236), .B(n1227), .Z(n1122) );
XOR2_X1 U948 ( .A(G107), .B(n1237), .Z(n1227) );
NAND2_X1 U949 ( .A1(KEYINPUT21), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U950 ( .A(n1239), .B(KEYINPUT58), .ZN(n1120) );
NAND2_X1 U951 ( .A1(n1209), .A2(n1202), .ZN(n1145) );
XNOR2_X1 U952 ( .A(n1044), .B(n1240), .ZN(n1202) );
NOR2_X1 U953 ( .A1(n1043), .A2(KEYINPUT33), .ZN(n1240) );
AND2_X1 U954 ( .A1(n1241), .A2(n1221), .ZN(n1043) );
XOR2_X1 U955 ( .A(KEYINPUT62), .B(n1242), .Z(n1241) );
INV_X1 U956 ( .A(n1086), .ZN(n1242) );
XOR2_X1 U957 ( .A(n1243), .B(n1244), .Z(n1086) );
XOR2_X1 U958 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U959 ( .A(G107), .B(n1247), .Z(n1246) );
NOR3_X1 U960 ( .A1(n1214), .A2(G953), .A3(n1083), .ZN(n1247) );
INV_X1 U961 ( .A(G217), .ZN(n1083) );
XNOR2_X1 U962 ( .A(G116), .B(n1248), .ZN(n1243) );
XOR2_X1 U963 ( .A(G134), .B(G122), .Z(n1248) );
INV_X1 U964 ( .A(G478), .ZN(n1044) );
XOR2_X1 U965 ( .A(n1249), .B(G475), .Z(n1209) );
NAND2_X1 U966 ( .A1(KEYINPUT26), .A2(n1041), .ZN(n1249) );
NOR2_X1 U967 ( .A1(n1090), .A2(n1250), .ZN(n1041) );
INV_X1 U968 ( .A(n1221), .ZN(n1250) );
XNOR2_X1 U969 ( .A(n1251), .B(n1252), .ZN(n1090) );
XOR2_X1 U970 ( .A(G122), .B(n1253), .Z(n1252) );
XOR2_X1 U971 ( .A(G146), .B(G131), .Z(n1253) );
XOR2_X1 U972 ( .A(n1254), .B(n1255), .Z(n1251) );
XOR2_X1 U973 ( .A(n1205), .B(n1256), .Z(n1255) );
NAND3_X1 U974 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
OR2_X1 U975 ( .A1(n1060), .A2(n1260), .ZN(n1259) );
NAND3_X1 U976 ( .A1(n1260), .A2(n1060), .A3(KEYINPUT3), .ZN(n1258) );
INV_X1 U977 ( .A(G140), .ZN(n1060) );
NOR2_X1 U978 ( .A1(G125), .A2(KEYINPUT20), .ZN(n1260) );
OR2_X1 U979 ( .A1(n1061), .A2(KEYINPUT3), .ZN(n1257) );
INV_X1 U980 ( .A(G125), .ZN(n1061) );
NAND2_X1 U981 ( .A1(n1261), .A2(n1262), .ZN(n1254) );
NAND2_X1 U982 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XNOR2_X1 U983 ( .A(KEYINPUT38), .B(n1265), .ZN(n1263) );
NAND2_X1 U984 ( .A1(n1266), .A2(n1267), .ZN(n1261) );
XOR2_X1 U985 ( .A(n1265), .B(KEYINPUT53), .Z(n1267) );
NAND2_X1 U986 ( .A1(KEYINPUT18), .A2(n1237), .ZN(n1265) );
XOR2_X1 U987 ( .A(G104), .B(KEYINPUT50), .Z(n1237) );
INV_X1 U988 ( .A(n1264), .ZN(n1266) );
XOR2_X1 U989 ( .A(n1268), .B(G143), .Z(n1264) );
NAND3_X1 U990 ( .A1(n1269), .A2(n988), .A3(G214), .ZN(n1268) );
INV_X1 U991 ( .A(G953), .ZN(n988) );
INV_X1 U992 ( .A(n1184), .ZN(n1017) );
NOR2_X1 U993 ( .A1(n1210), .A2(n1189), .ZN(n1184) );
XOR2_X1 U994 ( .A(n1034), .B(n1036), .Z(n1189) );
AND2_X1 U995 ( .A1(G217), .A2(n1270), .ZN(n1036) );
XOR2_X1 U996 ( .A(KEYINPUT10), .B(n1230), .Z(n1270) );
NOR2_X1 U997 ( .A1(n1214), .A2(G902), .ZN(n1230) );
NAND2_X1 U998 ( .A1(n1080), .A2(n1221), .ZN(n1034) );
XNOR2_X1 U999 ( .A(n1271), .B(n1272), .ZN(n1080) );
NOR4_X1 U1000 ( .A1(KEYINPUT7), .A2(G953), .A3(n1214), .A4(n1229), .ZN(n1272) );
INV_X1 U1001 ( .A(G221), .ZN(n1229) );
INV_X1 U1002 ( .A(G234), .ZN(n1214) );
XOR2_X1 U1003 ( .A(n1273), .B(n1274), .Z(n1271) );
NOR2_X1 U1004 ( .A1(KEYINPUT31), .A2(n1275), .ZN(n1274) );
XOR2_X1 U1005 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U1006 ( .A(G140), .B(n1278), .Z(n1277) );
XOR2_X1 U1007 ( .A(KEYINPUT0), .B(G146), .Z(n1278) );
XOR2_X1 U1008 ( .A(n1279), .B(n1280), .Z(n1276) );
NOR2_X1 U1009 ( .A1(KEYINPUT43), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1010 ( .A(n1282), .B(n1283), .Z(n1281) );
INV_X1 U1011 ( .A(G128), .ZN(n1282) );
XOR2_X1 U1012 ( .A(n1117), .B(G125), .Z(n1279) );
INV_X1 U1013 ( .A(G110), .ZN(n1117) );
INV_X1 U1014 ( .A(G137), .ZN(n1273) );
INV_X1 U1015 ( .A(n1190), .ZN(n1210) );
XOR2_X1 U1016 ( .A(n1031), .B(G472), .Z(n1190) );
NAND2_X1 U1017 ( .A1(n1284), .A2(n1221), .ZN(n1031) );
XOR2_X1 U1018 ( .A(G902), .B(KEYINPUT8), .Z(n1221) );
XOR2_X1 U1019 ( .A(n1100), .B(KEYINPUT37), .Z(n1284) );
XOR2_X1 U1020 ( .A(n1285), .B(n1239), .Z(n1100) );
XOR2_X1 U1021 ( .A(n1064), .B(n1063), .Z(n1239) );
XOR2_X1 U1022 ( .A(G146), .B(n1245), .Z(n1063) );
XOR2_X1 U1023 ( .A(G128), .B(G143), .Z(n1245) );
XOR2_X1 U1024 ( .A(G131), .B(n1286), .Z(n1064) );
XOR2_X1 U1025 ( .A(G137), .B(G134), .Z(n1286) );
XOR2_X1 U1026 ( .A(n1226), .B(n1287), .Z(n1285) );
NOR3_X1 U1027 ( .A1(n1219), .A2(G953), .A3(n1288), .ZN(n1287) );
XOR2_X1 U1028 ( .A(n1269), .B(KEYINPUT57), .Z(n1288) );
INV_X1 U1029 ( .A(G237), .ZN(n1269) );
INV_X1 U1030 ( .A(G210), .ZN(n1219) );
XOR2_X1 U1031 ( .A(n1289), .B(n1290), .Z(n1226) );
XOR2_X1 U1032 ( .A(n1238), .B(n1283), .Z(n1290) );
XOR2_X1 U1033 ( .A(G119), .B(KEYINPUT30), .Z(n1283) );
XOR2_X1 U1034 ( .A(G101), .B(KEYINPUT5), .Z(n1238) );
XOR2_X1 U1035 ( .A(n1205), .B(n1291), .Z(n1289) );
XOR2_X1 U1036 ( .A(KEYINPUT32), .B(G116), .Z(n1291) );
INV_X1 U1037 ( .A(G113), .ZN(n1205) );
endmodule


