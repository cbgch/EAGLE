//Key = 0010101111010000111101101011100000000110101011100010011011111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;

XOR2_X1 U738 ( .A(n1013), .B(n1014), .Z(G9) );
NAND3_X1 U739 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND2_X1 U740 ( .A1(KEYINPUT58), .A2(G107), .ZN(n1013) );
NAND4_X1 U741 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(G75) );
NOR2_X1 U742 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR4_X1 U743 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
XOR2_X1 U744 ( .A(n1028), .B(KEYINPUT7), .Z(n1027) );
NAND2_X1 U745 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR2_X1 U746 ( .A1(G475), .A2(n1031), .ZN(n1026) );
NAND3_X1 U747 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1025) );
NAND2_X1 U748 ( .A1(G469), .A2(n1035), .ZN(n1034) );
NAND4_X1 U749 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1024) );
NOR2_X1 U750 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
XNOR2_X1 U751 ( .A(G472), .B(n1042), .ZN(n1041) );
XOR2_X1 U752 ( .A(KEYINPUT3), .B(n1043), .Z(n1040) );
NOR3_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
AND2_X1 U754 ( .A1(n1047), .A2(KEYINPUT0), .ZN(n1046) );
NOR3_X1 U755 ( .A1(KEYINPUT0), .A2(n1048), .A3(n1049), .ZN(n1045) );
AND2_X1 U756 ( .A1(n1049), .A2(n1048), .ZN(n1044) );
NAND2_X1 U757 ( .A1(KEYINPUT11), .A2(n1050), .ZN(n1049) );
XOR2_X1 U758 ( .A(KEYINPUT4), .B(n1051), .Z(n1037) );
NOR2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U760 ( .A1(G953), .A2(n1054), .ZN(n1019) );
NAND3_X1 U761 ( .A1(G952), .A2(n1055), .A3(n1056), .ZN(n1018) );
NAND2_X1 U762 ( .A1(n1054), .A2(n1057), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U764 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND3_X1 U765 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NAND3_X1 U766 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1063) );
NAND2_X1 U767 ( .A1(n1016), .A2(n1068), .ZN(n1067) );
OR2_X1 U768 ( .A1(n1069), .A2(n1015), .ZN(n1068) );
NAND2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
NAND2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U771 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
INV_X1 U772 ( .A(KEYINPUT20), .ZN(n1075) );
INV_X1 U773 ( .A(n1076), .ZN(n1072) );
NAND3_X1 U774 ( .A1(KEYINPUT20), .A2(n1074), .A3(n1077), .ZN(n1065) );
INV_X1 U775 ( .A(n1070), .ZN(n1077) );
NAND3_X1 U776 ( .A1(n1016), .A2(n1078), .A3(n1070), .ZN(n1060) );
NAND3_X1 U777 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NAND2_X1 U778 ( .A1(n1062), .A2(n1082), .ZN(n1081) );
NAND2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1038), .ZN(n1084) );
XOR2_X1 U781 ( .A(n1033), .B(KEYINPUT9), .Z(n1085) );
NAND3_X1 U782 ( .A1(n1064), .A2(n1086), .A3(n1087), .ZN(n1079) );
XOR2_X1 U783 ( .A(n1088), .B(KEYINPUT52), .Z(n1058) );
INV_X1 U784 ( .A(KEYINPUT39), .ZN(n1054) );
XOR2_X1 U785 ( .A(n1089), .B(n1090), .Z(G72) );
XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U788 ( .A(n1095), .B(n1096), .Z(n1094) );
XNOR2_X1 U789 ( .A(n1097), .B(n1098), .ZN(n1096) );
XNOR2_X1 U790 ( .A(n1099), .B(n1100), .ZN(n1095) );
XNOR2_X1 U791 ( .A(KEYINPUT63), .B(KEYINPUT32), .ZN(n1099) );
NOR2_X1 U792 ( .A1(G900), .A2(n1056), .ZN(n1093) );
NOR2_X1 U793 ( .A1(G953), .A2(n1101), .ZN(n1091) );
NOR2_X1 U794 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U795 ( .A(KEYINPUT1), .B(n1104), .Z(n1103) );
NOR2_X1 U796 ( .A1(n1105), .A2(n1056), .ZN(n1089) );
AND2_X1 U797 ( .A1(G227), .A2(G900), .ZN(n1105) );
XOR2_X1 U798 ( .A(n1106), .B(n1107), .Z(G69) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U800 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND2_X1 U801 ( .A1(n1111), .A2(G898), .ZN(n1110) );
XNOR2_X1 U802 ( .A(G224), .B(KEYINPUT60), .ZN(n1111) );
NAND2_X1 U803 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
OR2_X1 U804 ( .A1(n1056), .A2(G898), .ZN(n1113) );
XOR2_X1 U805 ( .A(n1114), .B(n1115), .Z(n1112) );
XOR2_X1 U806 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U807 ( .A1(KEYINPUT45), .A2(n1118), .ZN(n1116) );
AND2_X1 U808 ( .A1(n1119), .A2(n1056), .ZN(n1106) );
NOR2_X1 U809 ( .A1(n1022), .A2(n1120), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1048), .A2(n1121), .A3(n1122), .ZN(n1120) );
NOR4_X1 U811 ( .A1(n1123), .A2(n1124), .A3(KEYINPUT15), .A4(n1050), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
NOR3_X1 U813 ( .A1(n1050), .A2(KEYINPUT15), .A3(n1020), .ZN(n1125) );
NOR2_X1 U814 ( .A1(n1022), .A2(n1127), .ZN(G63) );
XOR2_X1 U815 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U816 ( .A1(n1130), .A2(n1124), .ZN(n1128) );
NOR2_X1 U817 ( .A1(n1022), .A2(n1131), .ZN(G60) );
NOR3_X1 U818 ( .A1(n1052), .A2(n1132), .A3(n1133), .ZN(n1131) );
NOR3_X1 U819 ( .A1(n1134), .A2(n1053), .A3(n1124), .ZN(n1133) );
NOR2_X1 U820 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1020), .A2(n1053), .ZN(n1135) );
INV_X1 U822 ( .A(G475), .ZN(n1053) );
XNOR2_X1 U823 ( .A(n1137), .B(n1138), .ZN(G6) );
XNOR2_X1 U824 ( .A(G104), .B(KEYINPUT62), .ZN(n1138) );
NOR2_X1 U825 ( .A1(n1139), .A2(n1140), .ZN(G57) );
XOR2_X1 U826 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U827 ( .A(KEYINPUT42), .B(n1143), .Z(n1142) );
NOR2_X1 U828 ( .A1(n1144), .A2(n1124), .ZN(n1143) );
XNOR2_X1 U829 ( .A(n1145), .B(n1146), .ZN(n1141) );
NOR2_X1 U830 ( .A1(KEYINPUT34), .A2(n1147), .ZN(n1146) );
NOR2_X1 U831 ( .A1(n1148), .A2(n1056), .ZN(n1139) );
XNOR2_X1 U832 ( .A(G952), .B(KEYINPUT16), .ZN(n1148) );
NOR2_X1 U833 ( .A1(n1022), .A2(n1149), .ZN(G54) );
XOR2_X1 U834 ( .A(n1150), .B(n1151), .Z(n1149) );
XNOR2_X1 U835 ( .A(n1152), .B(n1153), .ZN(n1151) );
NAND2_X1 U836 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND3_X1 U837 ( .A1(n1156), .A2(n1097), .A3(n1157), .ZN(n1155) );
INV_X1 U838 ( .A(KEYINPUT38), .ZN(n1157) );
NAND2_X1 U839 ( .A1(n1158), .A2(KEYINPUT38), .ZN(n1154) );
XOR2_X1 U840 ( .A(n1159), .B(n1160), .Z(n1150) );
NOR2_X1 U841 ( .A1(n1030), .A2(n1124), .ZN(n1160) );
INV_X1 U842 ( .A(G469), .ZN(n1030) );
NAND2_X1 U843 ( .A1(KEYINPUT50), .A2(n1161), .ZN(n1159) );
NOR2_X1 U844 ( .A1(n1022), .A2(n1162), .ZN(G51) );
XNOR2_X1 U845 ( .A(n1163), .B(n1164), .ZN(n1162) );
NOR2_X1 U846 ( .A1(n1165), .A2(n1124), .ZN(n1164) );
OR2_X1 U847 ( .A1(n1166), .A2(n1020), .ZN(n1124) );
NOR3_X1 U848 ( .A1(n1102), .A2(n1104), .A3(n1119), .ZN(n1020) );
NAND4_X1 U849 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1119) );
AND4_X1 U850 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1170) );
NOR2_X1 U851 ( .A1(n1137), .A2(n1175), .ZN(n1169) );
NOR4_X1 U852 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
INV_X1 U853 ( .A(n1016), .ZN(n1178) );
NOR2_X1 U854 ( .A1(KEYINPUT46), .A2(n1180), .ZN(n1177) );
NOR3_X1 U855 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1180) );
NOR2_X1 U856 ( .A1(n1017), .A2(n1184), .ZN(n1176) );
INV_X1 U857 ( .A(KEYINPUT46), .ZN(n1184) );
AND3_X1 U858 ( .A1(n1017), .A2(n1016), .A3(n1069), .ZN(n1137) );
NAND4_X1 U859 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1102) );
AND4_X1 U860 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188) );
NAND2_X1 U861 ( .A1(KEYINPUT19), .A2(n1193), .ZN(n1187) );
NAND3_X1 U862 ( .A1(n1194), .A2(n1015), .A3(n1195), .ZN(n1186) );
NAND2_X1 U863 ( .A1(n1196), .A2(n1197), .ZN(n1185) );
NAND2_X1 U864 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
OR3_X1 U865 ( .A1(n1064), .A2(KEYINPUT19), .A3(n1181), .ZN(n1199) );
NAND2_X1 U866 ( .A1(n1062), .A2(n1182), .ZN(n1198) );
NOR2_X1 U867 ( .A1(n1056), .A2(G952), .ZN(n1022) );
XOR2_X1 U868 ( .A(G146), .B(n1104), .Z(G48) );
AND3_X1 U869 ( .A1(n1069), .A2(n1182), .A3(n1200), .ZN(n1104) );
XNOR2_X1 U870 ( .A(G143), .B(n1192), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1074), .A2(n1201), .A3(n1194), .A4(n1202), .ZN(n1192) );
NOR3_X1 U872 ( .A1(n1083), .A2(n1036), .A3(n1203), .ZN(n1202) );
INV_X1 U873 ( .A(n1204), .ZN(n1036) );
XOR2_X1 U874 ( .A(G140), .B(n1193), .Z(G42) );
AND2_X1 U875 ( .A1(n1196), .A2(n1205), .ZN(n1193) );
AND3_X1 U876 ( .A1(n1076), .A2(n1069), .A3(n1194), .ZN(n1196) );
XOR2_X1 U877 ( .A(n1191), .B(n1206), .Z(G39) );
NAND2_X1 U878 ( .A1(KEYINPUT27), .A2(G137), .ZN(n1206) );
NAND3_X1 U879 ( .A1(n1200), .A2(n1070), .A3(n1064), .ZN(n1191) );
XOR2_X1 U880 ( .A(n1207), .B(G134), .Z(G36) );
NAND2_X1 U881 ( .A1(KEYINPUT2), .A2(n1208), .ZN(n1207) );
NAND3_X1 U882 ( .A1(n1195), .A2(n1015), .A3(n1209), .ZN(n1208) );
XNOR2_X1 U883 ( .A(n1194), .B(KEYINPUT26), .ZN(n1209) );
XNOR2_X1 U884 ( .A(G131), .B(n1190), .ZN(G33) );
NAND3_X1 U885 ( .A1(n1194), .A2(n1069), .A3(n1195), .ZN(n1190) );
AND2_X1 U886 ( .A1(n1205), .A2(n1074), .ZN(n1195) );
INV_X1 U887 ( .A(n1080), .ZN(n1205) );
NAND2_X1 U888 ( .A1(n1064), .A2(n1201), .ZN(n1080) );
AND2_X1 U889 ( .A1(n1210), .A2(n1038), .ZN(n1064) );
INV_X1 U890 ( .A(n1211), .ZN(n1038) );
XOR2_X1 U891 ( .A(n1033), .B(KEYINPUT35), .Z(n1210) );
NAND2_X1 U892 ( .A1(n1212), .A2(n1213), .ZN(G30) );
OR2_X1 U893 ( .A1(n1214), .A2(G128), .ZN(n1213) );
NAND2_X1 U894 ( .A1(G128), .A2(n1215), .ZN(n1212) );
NAND2_X1 U895 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U896 ( .A1(KEYINPUT29), .A2(n1218), .ZN(n1217) );
NAND2_X1 U897 ( .A1(n1214), .A2(n1219), .ZN(n1216) );
INV_X1 U898 ( .A(KEYINPUT29), .ZN(n1219) );
NAND2_X1 U899 ( .A1(KEYINPUT54), .A2(n1218), .ZN(n1214) );
INV_X1 U900 ( .A(n1189), .ZN(n1218) );
NAND3_X1 U901 ( .A1(n1015), .A2(n1182), .A3(n1200), .ZN(n1189) );
NOR4_X1 U902 ( .A1(n1220), .A2(n1221), .A3(n1181), .A4(n1222), .ZN(n1200) );
XOR2_X1 U903 ( .A(n1167), .B(n1223), .Z(G3) );
XNOR2_X1 U904 ( .A(KEYINPUT28), .B(n1224), .ZN(n1223) );
NAND3_X1 U905 ( .A1(n1074), .A2(n1017), .A3(n1070), .ZN(n1167) );
XNOR2_X1 U906 ( .A(G125), .B(n1225), .ZN(G27) );
NAND2_X1 U907 ( .A1(n1226), .A2(n1182), .ZN(n1225) );
INV_X1 U908 ( .A(n1083), .ZN(n1182) );
XOR2_X1 U909 ( .A(n1227), .B(KEYINPUT18), .Z(n1226) );
NAND4_X1 U910 ( .A1(n1194), .A2(n1076), .A3(n1062), .A4(n1228), .ZN(n1227) );
XOR2_X1 U911 ( .A(KEYINPUT48), .B(n1069), .Z(n1228) );
INV_X1 U912 ( .A(n1229), .ZN(n1062) );
INV_X1 U913 ( .A(n1221), .ZN(n1194) );
NAND2_X1 U914 ( .A1(n1230), .A2(n1231), .ZN(n1221) );
NAND2_X1 U915 ( .A1(G900), .A2(G953), .ZN(n1231) );
XNOR2_X1 U916 ( .A(G122), .B(n1168), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1232), .A2(n1016), .A3(n1233), .A4(n1204), .ZN(n1168) );
NOR2_X1 U918 ( .A1(n1234), .A2(n1235), .ZN(n1016) );
XNOR2_X1 U919 ( .A(G119), .B(n1174), .ZN(G21) );
NAND4_X1 U920 ( .A1(n1235), .A2(n1070), .A3(n1232), .A4(n1234), .ZN(n1174) );
XNOR2_X1 U921 ( .A(G116), .B(n1173), .ZN(G18) );
NAND3_X1 U922 ( .A1(n1232), .A2(n1015), .A3(n1074), .ZN(n1173) );
INV_X1 U923 ( .A(n1179), .ZN(n1015) );
NAND2_X1 U924 ( .A1(n1236), .A2(n1204), .ZN(n1179) );
XNOR2_X1 U925 ( .A(n1233), .B(KEYINPUT23), .ZN(n1236) );
XNOR2_X1 U926 ( .A(G113), .B(n1172), .ZN(G15) );
NAND3_X1 U927 ( .A1(n1074), .A2(n1232), .A3(n1069), .ZN(n1172) );
NOR2_X1 U928 ( .A1(n1204), .A2(n1203), .ZN(n1069) );
INV_X1 U929 ( .A(n1233), .ZN(n1203) );
NOR3_X1 U930 ( .A1(n1083), .A2(n1183), .A3(n1229), .ZN(n1232) );
NAND2_X1 U931 ( .A1(n1032), .A2(n1086), .ZN(n1229) );
NOR2_X1 U932 ( .A1(n1235), .A2(n1222), .ZN(n1074) );
INV_X1 U933 ( .A(n1234), .ZN(n1222) );
INV_X1 U934 ( .A(n1220), .ZN(n1235) );
XOR2_X1 U935 ( .A(n1171), .B(n1237), .Z(G12) );
NOR2_X1 U936 ( .A1(G110), .A2(KEYINPUT41), .ZN(n1237) );
NAND3_X1 U937 ( .A1(n1070), .A2(n1017), .A3(n1076), .ZN(n1171) );
NOR2_X1 U938 ( .A1(n1220), .A2(n1234), .ZN(n1076) );
XOR2_X1 U939 ( .A(n1238), .B(n1144), .Z(n1234) );
INV_X1 U940 ( .A(G472), .ZN(n1144) );
NAND2_X1 U941 ( .A1(KEYINPUT57), .A2(n1239), .ZN(n1238) );
INV_X1 U942 ( .A(n1042), .ZN(n1239) );
NAND2_X1 U943 ( .A1(n1240), .A2(n1166), .ZN(n1042) );
XNOR2_X1 U944 ( .A(n1147), .B(n1241), .ZN(n1240) );
INV_X1 U945 ( .A(n1145), .ZN(n1241) );
XNOR2_X1 U946 ( .A(n1242), .B(n1243), .ZN(n1145) );
XNOR2_X1 U947 ( .A(G113), .B(n1224), .ZN(n1243) );
XNOR2_X1 U948 ( .A(n1244), .B(n1245), .ZN(n1242) );
NOR2_X1 U949 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
INV_X1 U950 ( .A(G210), .ZN(n1246) );
XNOR2_X1 U951 ( .A(n1248), .B(n1249), .ZN(n1147) );
INV_X1 U952 ( .A(n1152), .ZN(n1249) );
XOR2_X1 U953 ( .A(n1048), .B(n1250), .Z(n1220) );
NOR2_X1 U954 ( .A1(n1047), .A2(KEYINPUT12), .ZN(n1250) );
INV_X1 U955 ( .A(n1050), .ZN(n1047) );
NAND2_X1 U956 ( .A1(G217), .A2(n1251), .ZN(n1050) );
NOR2_X1 U957 ( .A1(n1126), .A2(G902), .ZN(n1048) );
INV_X1 U958 ( .A(n1123), .ZN(n1126) );
XNOR2_X1 U959 ( .A(n1252), .B(n1253), .ZN(n1123) );
XOR2_X1 U960 ( .A(G137), .B(n1254), .Z(n1253) );
AND3_X1 U961 ( .A1(G221), .A2(n1056), .A3(G234), .ZN(n1254) );
NAND2_X1 U962 ( .A1(n1255), .A2(KEYINPUT37), .ZN(n1252) );
XOR2_X1 U963 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U964 ( .A(G110), .B(n1258), .Z(n1257) );
XOR2_X1 U965 ( .A(KEYINPUT33), .B(G119), .Z(n1258) );
XOR2_X1 U966 ( .A(n1259), .B(n1260), .Z(n1256) );
NOR3_X1 U967 ( .A1(n1083), .A2(n1183), .A3(n1181), .ZN(n1017) );
INV_X1 U968 ( .A(n1201), .ZN(n1181) );
NOR2_X1 U969 ( .A1(n1086), .A2(n1087), .ZN(n1201) );
INV_X1 U970 ( .A(n1032), .ZN(n1087) );
NAND2_X1 U971 ( .A1(G221), .A2(n1251), .ZN(n1032) );
NAND2_X1 U972 ( .A1(n1261), .A2(n1166), .ZN(n1251) );
NAND3_X1 U973 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1086) );
NAND2_X1 U974 ( .A1(G469), .A2(n1265), .ZN(n1264) );
OR3_X1 U975 ( .A1(n1265), .A2(G469), .A3(KEYINPUT43), .ZN(n1263) );
OR2_X1 U976 ( .A1(n1029), .A2(KEYINPUT55), .ZN(n1265) );
NAND2_X1 U977 ( .A1(KEYINPUT43), .A2(n1029), .ZN(n1262) );
INV_X1 U978 ( .A(n1035), .ZN(n1029) );
NAND2_X1 U979 ( .A1(n1266), .A2(n1166), .ZN(n1035) );
XOR2_X1 U980 ( .A(n1161), .B(n1267), .Z(n1266) );
XNOR2_X1 U981 ( .A(n1158), .B(n1152), .ZN(n1267) );
XOR2_X1 U982 ( .A(G131), .B(n1268), .Z(n1152) );
NOR2_X1 U983 ( .A1(KEYINPUT30), .A2(n1100), .ZN(n1268) );
XNOR2_X1 U984 ( .A(G134), .B(G137), .ZN(n1100) );
XOR2_X1 U985 ( .A(n1097), .B(n1156), .Z(n1158) );
AND3_X1 U986 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1156) );
NAND2_X1 U987 ( .A1(n1272), .A2(n1224), .ZN(n1271) );
OR3_X1 U988 ( .A1(n1224), .A2(G104), .A3(G107), .ZN(n1270) );
INV_X1 U989 ( .A(G101), .ZN(n1224) );
NAND2_X1 U990 ( .A1(n1273), .A2(G107), .ZN(n1269) );
XNOR2_X1 U991 ( .A(G101), .B(G104), .ZN(n1273) );
XNOR2_X1 U992 ( .A(n1248), .B(KEYINPUT49), .ZN(n1097) );
XOR2_X1 U993 ( .A(n1274), .B(n1275), .Z(n1161) );
XOR2_X1 U994 ( .A(G140), .B(G110), .Z(n1275) );
NAND2_X1 U995 ( .A1(G227), .A2(n1056), .ZN(n1274) );
NAND2_X1 U996 ( .A1(n1230), .A2(n1276), .ZN(n1183) );
NAND2_X1 U997 ( .A1(G898), .A2(G953), .ZN(n1276) );
AND3_X1 U998 ( .A1(n1277), .A2(n1278), .A3(n1088), .ZN(n1230) );
NAND2_X1 U999 ( .A1(n1261), .A2(n1279), .ZN(n1088) );
XNOR2_X1 U1000 ( .A(KEYINPUT36), .B(n1280), .ZN(n1279) );
XNOR2_X1 U1001 ( .A(G234), .B(KEYINPUT44), .ZN(n1261) );
OR2_X1 U1002 ( .A1(G952), .A2(G953), .ZN(n1278) );
NAND2_X1 U1003 ( .A1(n1281), .A2(G953), .ZN(n1277) );
XNOR2_X1 U1004 ( .A(KEYINPUT56), .B(n1166), .ZN(n1281) );
NAND2_X1 U1005 ( .A1(n1211), .A2(n1033), .ZN(n1083) );
NAND2_X1 U1006 ( .A1(G214), .A2(n1282), .ZN(n1033) );
XOR2_X1 U1007 ( .A(n1283), .B(n1165), .Z(n1211) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1282), .ZN(n1165) );
NAND2_X1 U1009 ( .A1(n1166), .A2(n1280), .ZN(n1282) );
NAND2_X1 U1010 ( .A1(n1163), .A2(n1166), .ZN(n1283) );
INV_X1 U1011 ( .A(G902), .ZN(n1166) );
XNOR2_X1 U1012 ( .A(n1284), .B(n1285), .ZN(n1163) );
XOR2_X1 U1013 ( .A(G125), .B(n1286), .Z(n1285) );
NOR2_X1 U1014 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U1015 ( .A(n1289), .B(KEYINPUT53), .Z(n1288) );
NAND2_X1 U1016 ( .A1(n1290), .A2(n1117), .ZN(n1289) );
NOR2_X1 U1017 ( .A1(n1117), .A2(n1290), .ZN(n1287) );
XNOR2_X1 U1018 ( .A(n1114), .B(n1118), .ZN(n1290) );
XNOR2_X1 U1019 ( .A(n1291), .B(G113), .ZN(n1118) );
NAND2_X1 U1020 ( .A1(KEYINPUT21), .A2(n1244), .ZN(n1291) );
XOR2_X1 U1021 ( .A(G116), .B(G119), .Z(n1244) );
XOR2_X1 U1022 ( .A(G101), .B(n1292), .Z(n1114) );
NOR2_X1 U1023 ( .A1(n1272), .A2(n1293), .ZN(n1292) );
XOR2_X1 U1024 ( .A(KEYINPUT25), .B(n1294), .Z(n1293) );
NOR2_X1 U1025 ( .A1(G104), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1026 ( .A(KEYINPUT6), .B(G107), .Z(n1295) );
NOR2_X1 U1027 ( .A1(n1296), .A2(G107), .ZN(n1272) );
XNOR2_X1 U1028 ( .A(G110), .B(G122), .ZN(n1117) );
XOR2_X1 U1029 ( .A(n1248), .B(n1297), .Z(n1284) );
AND2_X1 U1030 ( .A1(n1056), .A2(G224), .ZN(n1297) );
XNOR2_X1 U1031 ( .A(n1259), .B(n1298), .ZN(n1248) );
INV_X1 U1032 ( .A(G143), .ZN(n1298) );
XNOR2_X1 U1033 ( .A(G146), .B(n1299), .ZN(n1259) );
NOR2_X1 U1034 ( .A1(n1204), .A2(n1233), .ZN(n1070) );
XOR2_X1 U1035 ( .A(n1300), .B(n1031), .Z(n1233) );
INV_X1 U1036 ( .A(n1052), .ZN(n1031) );
NOR2_X1 U1037 ( .A1(n1136), .A2(G902), .ZN(n1052) );
INV_X1 U1038 ( .A(n1134), .ZN(n1136) );
XNOR2_X1 U1039 ( .A(n1301), .B(n1302), .ZN(n1134) );
XOR2_X1 U1040 ( .A(n1098), .B(n1303), .Z(n1302) );
XNOR2_X1 U1041 ( .A(n1304), .B(n1305), .ZN(n1303) );
NOR2_X1 U1042 ( .A1(KEYINPUT14), .A2(n1296), .ZN(n1305) );
INV_X1 U1043 ( .A(G104), .ZN(n1296) );
NAND2_X1 U1044 ( .A1(n1306), .A2(KEYINPUT22), .ZN(n1304) );
XNOR2_X1 U1045 ( .A(G146), .B(KEYINPUT61), .ZN(n1306) );
XOR2_X1 U1046 ( .A(G131), .B(n1260), .Z(n1098) );
XOR2_X1 U1047 ( .A(G125), .B(G140), .Z(n1260) );
XOR2_X1 U1048 ( .A(n1307), .B(n1308), .Z(n1301) );
XOR2_X1 U1049 ( .A(G113), .B(n1309), .Z(n1308) );
NOR2_X1 U1050 ( .A1(n1310), .A2(n1247), .ZN(n1309) );
NAND2_X1 U1051 ( .A1(n1311), .A2(n1056), .ZN(n1247) );
XNOR2_X1 U1052 ( .A(KEYINPUT59), .B(n1280), .ZN(n1311) );
INV_X1 U1053 ( .A(G237), .ZN(n1280) );
INV_X1 U1054 ( .A(G214), .ZN(n1310) );
XNOR2_X1 U1055 ( .A(G122), .B(G143), .ZN(n1307) );
NAND2_X1 U1056 ( .A1(KEYINPUT17), .A2(G475), .ZN(n1300) );
XOR2_X1 U1057 ( .A(n1312), .B(n1130), .Z(n1204) );
INV_X1 U1058 ( .A(G478), .ZN(n1130) );
OR2_X1 U1059 ( .A1(n1129), .A2(G902), .ZN(n1312) );
XNOR2_X1 U1060 ( .A(n1313), .B(n1314), .ZN(n1129) );
XOR2_X1 U1061 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1062 ( .A(n1317), .B(G107), .ZN(n1316) );
INV_X1 U1063 ( .A(G122), .ZN(n1317) );
NOR4_X1 U1064 ( .A1(KEYINPUT13), .A2(n1318), .A3(n1319), .A4(n1320), .ZN(n1315) );
XNOR2_X1 U1065 ( .A(KEYINPUT51), .B(n1056), .ZN(n1320) );
INV_X1 U1066 ( .A(G953), .ZN(n1056) );
INV_X1 U1067 ( .A(G217), .ZN(n1319) );
INV_X1 U1068 ( .A(G234), .ZN(n1318) );
XOR2_X1 U1069 ( .A(n1321), .B(n1322), .Z(n1313) );
NOR2_X1 U1070 ( .A1(G116), .A2(KEYINPUT10), .ZN(n1322) );
NAND2_X1 U1071 ( .A1(n1323), .A2(n1324), .ZN(n1321) );
NAND2_X1 U1072 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1073 ( .A(n1327), .B(KEYINPUT5), .Z(n1323) );
OR2_X1 U1074 ( .A1(n1326), .A2(n1325), .ZN(n1327) );
XOR2_X1 U1075 ( .A(G134), .B(KEYINPUT31), .Z(n1325) );
NAND2_X1 U1076 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
OR2_X1 U1077 ( .A1(n1330), .A2(G143), .ZN(n1329) );
XOR2_X1 U1078 ( .A(n1331), .B(KEYINPUT47), .Z(n1328) );
NAND2_X1 U1079 ( .A1(n1332), .A2(n1330), .ZN(n1331) );
XNOR2_X1 U1080 ( .A(n1299), .B(KEYINPUT8), .ZN(n1330) );
XOR2_X1 U1081 ( .A(G128), .B(KEYINPUT24), .Z(n1299) );
XNOR2_X1 U1082 ( .A(G143), .B(KEYINPUT40), .ZN(n1332) );
endmodule


