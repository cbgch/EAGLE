//Key = 1101110111101100110101010111111101111010001000110111000100101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;

XNOR2_X1 U766 ( .A(G107), .B(n1061), .ZN(G9) );
NOR2_X1 U767 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR4_X1 U768 ( .A1(G953), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1063) );
NOR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR3_X1 U771 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
NOR2_X1 U772 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR3_X1 U773 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NOR3_X1 U774 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NOR2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1077) );
NOR2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1074) );
NOR3_X1 U778 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1069) );
NOR3_X1 U779 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1088) );
AND3_X1 U780 ( .A1(n1071), .A2(n1093), .A3(KEYINPUT43), .ZN(n1092) );
NOR2_X1 U781 ( .A1(n1094), .A2(n1071), .ZN(n1091) );
NOR2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U784 ( .A1(KEYINPUT43), .A2(n1099), .ZN(n1095) );
NOR2_X1 U785 ( .A1(n1100), .A2(n1073), .ZN(n1090) );
INV_X1 U786 ( .A(n1101), .ZN(n1073) );
NOR2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
INV_X1 U788 ( .A(n1084), .ZN(n1087) );
NOR3_X1 U789 ( .A1(n1064), .A2(G953), .A3(G952), .ZN(n1062) );
AND4_X1 U790 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1064) );
NOR4_X1 U791 ( .A1(n1108), .A2(n1109), .A3(n1089), .A4(n1110), .ZN(n1107) );
XNOR2_X1 U792 ( .A(n1111), .B(n1112), .ZN(n1110) );
NOR2_X1 U793 ( .A1(KEYINPUT54), .A2(n1113), .ZN(n1112) );
XOR2_X1 U794 ( .A(n1114), .B(n1115), .Z(n1108) );
NAND2_X1 U795 ( .A1(KEYINPUT38), .A2(n1116), .ZN(n1114) );
NOR3_X1 U796 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1104) );
XNOR2_X1 U798 ( .A(n1122), .B(KEYINPUT51), .ZN(n1120) );
XOR2_X1 U799 ( .A(n1123), .B(n1124), .Z(G72) );
NOR2_X1 U800 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
AND2_X1 U801 ( .A1(G227), .A2(G900), .ZN(n1125) );
NAND3_X1 U802 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1123) );
OR2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND3_X1 U804 ( .A1(n1131), .A2(n1130), .A3(n1132), .ZN(n1128) );
NAND2_X1 U805 ( .A1(n1133), .A2(n1134), .ZN(n1127) );
NAND2_X1 U806 ( .A1(n1135), .A2(n1130), .ZN(n1134) );
INV_X1 U807 ( .A(KEYINPUT20), .ZN(n1130) );
XNOR2_X1 U808 ( .A(n1131), .B(KEYINPUT16), .ZN(n1135) );
NOR2_X1 U809 ( .A1(G953), .A2(n1136), .ZN(n1131) );
INV_X1 U810 ( .A(n1132), .ZN(n1133) );
NAND2_X1 U811 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
XOR2_X1 U812 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U813 ( .A(n1141), .B(n1142), .ZN(n1140) );
XOR2_X1 U814 ( .A(n1143), .B(n1144), .Z(n1139) );
NOR2_X1 U815 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U816 ( .A(G125), .B(KEYINPUT27), .ZN(n1143) );
XOR2_X1 U817 ( .A(KEYINPUT13), .B(n1147), .Z(n1137) );
XOR2_X1 U818 ( .A(n1148), .B(n1149), .Z(G69) );
XOR2_X1 U819 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U820 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XNOR2_X1 U821 ( .A(KEYINPUT62), .B(n1126), .ZN(n1153) );
NOR2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1150) );
NAND2_X1 U824 ( .A1(G953), .A2(n1155), .ZN(n1157) );
XNOR2_X1 U825 ( .A(n1158), .B(n1159), .ZN(n1156) );
INV_X1 U826 ( .A(n1160), .ZN(n1159) );
XOR2_X1 U827 ( .A(n1161), .B(KEYINPUT34), .Z(n1158) );
NAND3_X1 U828 ( .A1(n1162), .A2(n1126), .A3(KEYINPUT19), .ZN(n1148) );
NAND2_X1 U829 ( .A1(n1163), .A2(n1061), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1164), .A2(n1165), .ZN(G66) );
XOR2_X1 U831 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U832 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
AND2_X1 U833 ( .A1(KEYINPUT37), .A2(n1170), .ZN(n1169) );
NOR2_X1 U834 ( .A1(KEYINPUT15), .A2(n1170), .ZN(n1168) );
OR2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XNOR2_X1 U836 ( .A(n1173), .B(KEYINPUT63), .ZN(n1164) );
NOR2_X1 U837 ( .A1(n1173), .A2(n1174), .ZN(G63) );
XNOR2_X1 U838 ( .A(n1175), .B(n1176), .ZN(n1174) );
NOR2_X1 U839 ( .A1(n1177), .A2(n1171), .ZN(n1176) );
INV_X1 U840 ( .A(G478), .ZN(n1177) );
NOR2_X1 U841 ( .A1(n1173), .A2(n1178), .ZN(G60) );
XNOR2_X1 U842 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U843 ( .A1(n1181), .A2(n1171), .ZN(n1180) );
XNOR2_X1 U844 ( .A(G104), .B(n1182), .ZN(G6) );
NOR2_X1 U845 ( .A1(n1183), .A2(n1184), .ZN(G57) );
XNOR2_X1 U846 ( .A(n1173), .B(KEYINPUT35), .ZN(n1184) );
NOR2_X1 U847 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
XOR2_X1 U848 ( .A(KEYINPUT48), .B(n1187), .Z(n1186) );
NOR2_X1 U849 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XNOR2_X1 U850 ( .A(G101), .B(n1190), .ZN(n1189) );
INV_X1 U851 ( .A(n1191), .ZN(n1188) );
NOR2_X1 U852 ( .A1(n1192), .A2(n1191), .ZN(n1185) );
XNOR2_X1 U853 ( .A(n1193), .B(n1194), .ZN(n1191) );
NOR2_X1 U854 ( .A1(n1111), .A2(n1171), .ZN(n1194) );
NAND2_X1 U855 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
INV_X1 U856 ( .A(n1197), .ZN(n1196) );
XNOR2_X1 U857 ( .A(n1198), .B(G101), .ZN(n1192) );
NOR2_X1 U858 ( .A1(n1173), .A2(n1199), .ZN(G54) );
XOR2_X1 U859 ( .A(n1200), .B(n1201), .Z(n1199) );
XOR2_X1 U860 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U861 ( .A1(n1204), .A2(n1171), .ZN(n1203) );
XOR2_X1 U862 ( .A(n1205), .B(KEYINPUT9), .Z(n1200) );
NAND2_X1 U863 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U864 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U865 ( .A(n1210), .B(KEYINPUT40), .Z(n1206) );
OR2_X1 U866 ( .A1(n1208), .A2(n1209), .ZN(n1210) );
NAND2_X1 U867 ( .A1(n1211), .A2(n1212), .ZN(n1208) );
NAND2_X1 U868 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U869 ( .A(n1215), .B(KEYINPUT44), .Z(n1211) );
NAND2_X1 U870 ( .A1(n1142), .A2(n1216), .ZN(n1215) );
NOR3_X1 U871 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(G51) );
AND2_X1 U872 ( .A1(KEYINPUT42), .A2(n1173), .ZN(n1219) );
NOR2_X1 U873 ( .A1(n1126), .A2(G952), .ZN(n1173) );
NOR3_X1 U874 ( .A1(KEYINPUT42), .A2(G953), .A3(G952), .ZN(n1218) );
XOR2_X1 U875 ( .A(n1220), .B(n1221), .Z(n1217) );
XNOR2_X1 U876 ( .A(n1222), .B(n1223), .ZN(n1221) );
NOR2_X1 U877 ( .A1(KEYINPUT18), .A2(n1224), .ZN(n1222) );
XOR2_X1 U878 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U879 ( .A(n1227), .B(n1228), .ZN(n1226) );
NAND2_X1 U880 ( .A1(KEYINPUT3), .A2(n1229), .ZN(n1225) );
XNOR2_X1 U881 ( .A(n1160), .B(n1230), .ZN(n1220) );
NOR2_X1 U882 ( .A1(n1231), .A2(n1171), .ZN(n1230) );
NAND2_X1 U883 ( .A1(G902), .A2(n1066), .ZN(n1171) );
NAND3_X1 U884 ( .A1(n1136), .A2(n1163), .A3(n1232), .ZN(n1066) );
XOR2_X1 U885 ( .A(n1061), .B(KEYINPUT45), .Z(n1232) );
NAND3_X1 U886 ( .A1(n1101), .A2(n1102), .A3(n1233), .ZN(n1061) );
AND4_X1 U887 ( .A1(n1234), .A2(n1235), .A3(n1182), .A4(n1236), .ZN(n1163) );
AND4_X1 U888 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
NAND3_X1 U889 ( .A1(n1233), .A2(n1101), .A3(n1103), .ZN(n1182) );
AND4_X1 U890 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1136) );
AND4_X1 U891 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1244) );
NOR2_X1 U892 ( .A1(n1249), .A2(n1250), .ZN(n1243) );
NOR2_X1 U893 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NOR2_X1 U894 ( .A1(n1253), .A2(n1254), .ZN(n1251) );
XNOR2_X1 U895 ( .A(n1103), .B(KEYINPUT25), .ZN(n1254) );
NOR2_X1 U896 ( .A1(KEYINPUT6), .A2(n1255), .ZN(n1253) );
NOR4_X1 U897 ( .A1(n1080), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1249) );
INV_X1 U898 ( .A(KEYINPUT6), .ZN(n1257) );
XOR2_X1 U899 ( .A(G122), .B(n1258), .Z(n1160) );
NAND2_X1 U900 ( .A1(n1259), .A2(n1260), .ZN(G48) );
NAND2_X1 U901 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U902 ( .A(n1263), .B(n1264), .Z(n1259) );
NOR2_X1 U903 ( .A1(n1261), .A2(n1262), .ZN(n1264) );
INV_X1 U904 ( .A(KEYINPUT28), .ZN(n1262) );
OR2_X1 U905 ( .A1(n1252), .A2(n1265), .ZN(n1263) );
XNOR2_X1 U906 ( .A(G143), .B(n1241), .ZN(G45) );
NAND4_X1 U907 ( .A1(n1266), .A2(n1080), .A3(n1109), .A4(n1267), .ZN(n1241) );
XNOR2_X1 U908 ( .A(G140), .B(n1242), .ZN(G42) );
NAND3_X1 U909 ( .A1(n1268), .A2(n1076), .A3(n1084), .ZN(n1242) );
XOR2_X1 U910 ( .A(n1248), .B(n1269), .Z(G39) );
NAND2_X1 U911 ( .A1(G137), .A2(n1270), .ZN(n1269) );
XOR2_X1 U912 ( .A(KEYINPUT39), .B(KEYINPUT17), .Z(n1270) );
NAND3_X1 U913 ( .A1(n1271), .A2(n1084), .A3(n1272), .ZN(n1248) );
XNOR2_X1 U914 ( .A(G134), .B(n1247), .ZN(G36) );
NAND3_X1 U915 ( .A1(n1266), .A2(n1102), .A3(n1084), .ZN(n1247) );
XNOR2_X1 U916 ( .A(G131), .B(n1246), .ZN(G33) );
NAND3_X1 U917 ( .A1(n1266), .A2(n1103), .A3(n1084), .ZN(n1246) );
NOR2_X1 U918 ( .A1(n1082), .A2(n1117), .ZN(n1084) );
INV_X1 U919 ( .A(n1083), .ZN(n1117) );
NOR3_X1 U920 ( .A1(n1086), .A2(n1273), .A3(n1099), .ZN(n1266) );
INV_X1 U921 ( .A(n1093), .ZN(n1099) );
XOR2_X1 U922 ( .A(n1274), .B(n1275), .Z(G30) );
NOR2_X1 U923 ( .A1(n1255), .A2(n1252), .ZN(n1275) );
NAND2_X1 U924 ( .A1(n1271), .A2(n1080), .ZN(n1252) );
INV_X1 U925 ( .A(n1256), .ZN(n1271) );
NAND3_X1 U926 ( .A1(n1098), .A2(n1076), .A3(n1276), .ZN(n1256) );
NOR2_X1 U927 ( .A1(KEYINPUT41), .A2(n1277), .ZN(n1274) );
XOR2_X1 U928 ( .A(n1234), .B(n1278), .Z(G3) );
XNOR2_X1 U929 ( .A(KEYINPUT49), .B(n1279), .ZN(n1278) );
NAND3_X1 U930 ( .A1(n1093), .A2(n1233), .A3(n1272), .ZN(n1234) );
XNOR2_X1 U931 ( .A(G125), .B(n1245), .ZN(G27) );
NAND3_X1 U932 ( .A1(n1280), .A2(n1080), .A3(n1268), .ZN(n1245) );
AND3_X1 U933 ( .A1(n1281), .A2(n1276), .A3(n1103), .ZN(n1268) );
NOR3_X1 U934 ( .A1(n1079), .A2(n1097), .A3(n1273), .ZN(n1276) );
AND2_X1 U935 ( .A1(n1068), .A2(n1282), .ZN(n1273) );
NAND3_X1 U936 ( .A1(G902), .A2(n1283), .A3(n1147), .ZN(n1282) );
NOR2_X1 U937 ( .A1(n1126), .A2(G900), .ZN(n1147) );
INV_X1 U938 ( .A(n1085), .ZN(n1079) );
XNOR2_X1 U939 ( .A(n1284), .B(n1235), .ZN(G24) );
NAND4_X1 U940 ( .A1(n1285), .A2(n1101), .A3(n1109), .A4(n1267), .ZN(n1235) );
NOR2_X1 U941 ( .A1(n1286), .A2(n1098), .ZN(n1101) );
NAND2_X1 U942 ( .A1(KEYINPUT29), .A2(n1287), .ZN(n1284) );
INV_X1 U943 ( .A(G122), .ZN(n1287) );
XNOR2_X1 U944 ( .A(G119), .B(n1240), .ZN(G21) );
NAND4_X1 U945 ( .A1(n1285), .A2(n1272), .A3(n1098), .A4(n1286), .ZN(n1240) );
XOR2_X1 U946 ( .A(n1237), .B(n1288), .Z(G18) );
NAND2_X1 U947 ( .A1(KEYINPUT36), .A2(G116), .ZN(n1288) );
NAND3_X1 U948 ( .A1(n1093), .A2(n1102), .A3(n1285), .ZN(n1237) );
INV_X1 U949 ( .A(n1255), .ZN(n1102) );
NAND2_X1 U950 ( .A1(n1289), .A2(n1267), .ZN(n1255) );
XNOR2_X1 U951 ( .A(G113), .B(n1239), .ZN(G15) );
NAND3_X1 U952 ( .A1(n1093), .A2(n1103), .A3(n1285), .ZN(n1239) );
NOR2_X1 U953 ( .A1(n1089), .A2(n1290), .ZN(n1285) );
NAND2_X1 U954 ( .A1(n1280), .A2(n1085), .ZN(n1089) );
INV_X1 U955 ( .A(n1076), .ZN(n1280) );
INV_X1 U956 ( .A(n1265), .ZN(n1103) );
NAND2_X1 U957 ( .A1(n1291), .A2(n1109), .ZN(n1265) );
NOR2_X1 U958 ( .A1(n1286), .A2(n1281), .ZN(n1093) );
NAND3_X1 U959 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(G12) );
OR2_X1 U960 ( .A1(G110), .A2(KEYINPUT47), .ZN(n1294) );
NAND3_X1 U961 ( .A1(KEYINPUT47), .A2(G110), .A3(n1238), .ZN(n1293) );
NAND2_X1 U962 ( .A1(n1295), .A2(n1296), .ZN(n1292) );
NAND2_X1 U963 ( .A1(n1297), .A2(KEYINPUT47), .ZN(n1296) );
XNOR2_X1 U964 ( .A(G110), .B(KEYINPUT1), .ZN(n1297) );
INV_X1 U965 ( .A(n1238), .ZN(n1295) );
NAND4_X1 U966 ( .A1(n1272), .A2(n1233), .A3(n1281), .A4(n1286), .ZN(n1238) );
INV_X1 U967 ( .A(n1097), .ZN(n1286) );
NOR2_X1 U968 ( .A1(n1298), .A2(n1119), .ZN(n1097) );
NOR2_X1 U969 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
INV_X1 U970 ( .A(n1172), .ZN(n1122) );
AND2_X1 U971 ( .A1(n1299), .A2(n1121), .ZN(n1298) );
NAND2_X1 U972 ( .A1(n1166), .A2(n1300), .ZN(n1121) );
XOR2_X1 U973 ( .A(n1301), .B(n1302), .Z(n1166) );
XOR2_X1 U974 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U975 ( .A(n1305), .B(n1306), .ZN(n1304) );
NOR2_X1 U976 ( .A1(KEYINPUT14), .A2(n1141), .ZN(n1306) );
NAND3_X1 U977 ( .A1(n1307), .A2(G221), .A3(KEYINPUT30), .ZN(n1305) );
XOR2_X1 U978 ( .A(n1308), .B(n1309), .Z(n1301) );
XNOR2_X1 U979 ( .A(n1310), .B(G125), .ZN(n1309) );
XNOR2_X1 U980 ( .A(G119), .B(G110), .ZN(n1308) );
XNOR2_X1 U981 ( .A(KEYINPUT32), .B(n1172), .ZN(n1299) );
NAND2_X1 U982 ( .A1(G217), .A2(n1311), .ZN(n1172) );
INV_X1 U983 ( .A(n1098), .ZN(n1281) );
XOR2_X1 U984 ( .A(n1113), .B(n1111), .Z(n1098) );
INV_X1 U985 ( .A(G472), .ZN(n1111) );
NAND2_X1 U986 ( .A1(n1312), .A2(n1300), .ZN(n1113) );
XOR2_X1 U987 ( .A(n1313), .B(n1314), .Z(n1312) );
NOR2_X1 U988 ( .A1(n1197), .A2(n1315), .ZN(n1314) );
XOR2_X1 U989 ( .A(n1195), .B(KEYINPUT12), .Z(n1315) );
NAND2_X1 U990 ( .A1(n1316), .A2(n1317), .ZN(n1195) );
NOR2_X1 U991 ( .A1(n1317), .A2(n1316), .ZN(n1197) );
XOR2_X1 U992 ( .A(n1318), .B(KEYINPUT5), .Z(n1316) );
NAND2_X1 U993 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
NAND2_X1 U994 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U995 ( .A(n1323), .B(KEYINPUT33), .Z(n1321) );
XNOR2_X1 U996 ( .A(n1209), .B(n1229), .ZN(n1317) );
NAND2_X1 U997 ( .A1(n1324), .A2(n1325), .ZN(n1313) );
NAND2_X1 U998 ( .A1(n1198), .A2(n1326), .ZN(n1325) );
NAND2_X1 U999 ( .A1(KEYINPUT58), .A2(n1327), .ZN(n1326) );
NAND2_X1 U1000 ( .A1(n1279), .A2(n1328), .ZN(n1327) );
INV_X1 U1001 ( .A(G101), .ZN(n1279) );
INV_X1 U1002 ( .A(n1190), .ZN(n1198) );
NAND2_X1 U1003 ( .A1(G101), .A2(n1329), .ZN(n1324) );
NAND2_X1 U1004 ( .A1(n1328), .A2(n1330), .ZN(n1329) );
NAND2_X1 U1005 ( .A1(KEYINPUT58), .A2(n1190), .ZN(n1330) );
NAND2_X1 U1006 ( .A1(n1331), .A2(n1332), .ZN(n1190) );
XNOR2_X1 U1007 ( .A(KEYINPUT59), .B(n1231), .ZN(n1332) );
INV_X1 U1008 ( .A(G210), .ZN(n1231) );
INV_X1 U1009 ( .A(KEYINPUT56), .ZN(n1328) );
NOR2_X1 U1010 ( .A1(n1290), .A2(n1086), .ZN(n1233) );
NAND2_X1 U1011 ( .A1(n1076), .A2(n1085), .ZN(n1086) );
NAND2_X1 U1012 ( .A1(G221), .A2(n1311), .ZN(n1085) );
NAND2_X1 U1013 ( .A1(G234), .A2(n1300), .ZN(n1311) );
XOR2_X1 U1014 ( .A(n1333), .B(n1204), .Z(n1076) );
INV_X1 U1015 ( .A(G469), .ZN(n1204) );
NAND2_X1 U1016 ( .A1(n1334), .A2(n1300), .ZN(n1333) );
XOR2_X1 U1017 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U1018 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1019 ( .A(n1209), .B(KEYINPUT11), .Z(n1338) );
NAND3_X1 U1020 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1209) );
INV_X1 U1021 ( .A(n1145), .ZN(n1341) );
NOR3_X1 U1022 ( .A1(n1342), .A2(G137), .A3(n1343), .ZN(n1145) );
NAND2_X1 U1023 ( .A1(n1146), .A2(n1344), .ZN(n1340) );
INV_X1 U1024 ( .A(KEYINPUT57), .ZN(n1344) );
NAND2_X1 U1025 ( .A1(n1345), .A2(n1346), .ZN(n1146) );
NAND3_X1 U1026 ( .A1(n1342), .A2(n1343), .A3(n1310), .ZN(n1346) );
NAND2_X1 U1027 ( .A1(n1347), .A2(G137), .ZN(n1345) );
XNOR2_X1 U1028 ( .A(n1343), .B(G131), .ZN(n1347) );
NAND2_X1 U1029 ( .A1(n1348), .A2(KEYINPUT57), .ZN(n1339) );
XNOR2_X1 U1030 ( .A(n1342), .B(n1349), .ZN(n1348) );
NOR2_X1 U1031 ( .A1(G134), .A2(n1310), .ZN(n1349) );
INV_X1 U1032 ( .A(G137), .ZN(n1310) );
INV_X1 U1033 ( .A(G131), .ZN(n1342) );
NAND2_X1 U1034 ( .A1(KEYINPUT31), .A2(n1213), .ZN(n1337) );
INV_X1 U1035 ( .A(n1142), .ZN(n1213) );
XOR2_X1 U1036 ( .A(n1229), .B(KEYINPUT22), .Z(n1142) );
XNOR2_X1 U1037 ( .A(n1350), .B(n1214), .ZN(n1335) );
NAND3_X1 U1038 ( .A1(n1351), .A2(n1352), .A3(KEYINPUT50), .ZN(n1350) );
NAND2_X1 U1039 ( .A1(KEYINPUT46), .A2(n1202), .ZN(n1352) );
XOR2_X1 U1040 ( .A(n1353), .B(n1354), .Z(n1202) );
OR3_X1 U1041 ( .A1(n1353), .A2(n1354), .A3(KEYINPUT46), .ZN(n1351) );
XNOR2_X1 U1042 ( .A(G110), .B(n1355), .ZN(n1354) );
INV_X1 U1043 ( .A(n1141), .ZN(n1355) );
NAND2_X1 U1044 ( .A1(G227), .A2(n1126), .ZN(n1353) );
NAND2_X1 U1045 ( .A1(n1080), .A2(n1356), .ZN(n1290) );
NAND2_X1 U1046 ( .A1(n1068), .A2(n1357), .ZN(n1356) );
NAND4_X1 U1047 ( .A1(G953), .A2(G902), .A3(n1283), .A4(n1155), .ZN(n1357) );
INV_X1 U1048 ( .A(G898), .ZN(n1155) );
NAND3_X1 U1049 ( .A1(n1283), .A2(n1126), .A3(G952), .ZN(n1068) );
NAND2_X1 U1050 ( .A1(G237), .A2(G234), .ZN(n1283) );
AND2_X1 U1051 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1358), .ZN(n1083) );
NAND2_X1 U1053 ( .A1(n1359), .A2(n1360), .ZN(n1082) );
NAND2_X1 U1054 ( .A1(n1115), .A2(n1116), .ZN(n1360) );
XOR2_X1 U1055 ( .A(n1361), .B(KEYINPUT52), .Z(n1359) );
OR2_X1 U1056 ( .A1(n1116), .A2(n1115), .ZN(n1361) );
AND2_X1 U1057 ( .A1(n1362), .A2(G210), .ZN(n1115) );
XOR2_X1 U1058 ( .A(n1358), .B(KEYINPUT24), .Z(n1362) );
OR2_X1 U1059 ( .A1(G902), .A2(G237), .ZN(n1358) );
NAND2_X1 U1060 ( .A1(n1363), .A2(n1300), .ZN(n1116) );
XOR2_X1 U1061 ( .A(n1364), .B(n1365), .Z(n1363) );
XNOR2_X1 U1062 ( .A(n1229), .B(n1258), .ZN(n1365) );
XOR2_X1 U1063 ( .A(G110), .B(KEYINPUT26), .Z(n1258) );
XOR2_X1 U1064 ( .A(G143), .B(n1303), .Z(n1229) );
XNOR2_X1 U1065 ( .A(n1277), .B(G146), .ZN(n1303) );
XOR2_X1 U1066 ( .A(n1366), .B(n1367), .Z(n1364) );
XOR2_X1 U1067 ( .A(n1223), .B(n1228), .Z(n1366) );
NOR2_X1 U1068 ( .A1(n1154), .A2(G953), .ZN(n1228) );
INV_X1 U1069 ( .A(G224), .ZN(n1154) );
NAND2_X1 U1070 ( .A1(KEYINPUT23), .A2(n1161), .ZN(n1223) );
XNOR2_X1 U1071 ( .A(n1368), .B(n1214), .ZN(n1161) );
INV_X1 U1072 ( .A(n1216), .ZN(n1214) );
XOR2_X1 U1073 ( .A(G101), .B(n1369), .Z(n1216) );
XNOR2_X1 U1074 ( .A(n1370), .B(G104), .ZN(n1369) );
NAND2_X1 U1075 ( .A1(n1319), .A2(n1371), .ZN(n1368) );
NAND2_X1 U1076 ( .A1(n1372), .A2(n1322), .ZN(n1371) );
INV_X1 U1077 ( .A(G119), .ZN(n1322) );
XOR2_X1 U1078 ( .A(n1323), .B(KEYINPUT0), .Z(n1372) );
NAND2_X1 U1079 ( .A1(G119), .A2(n1323), .ZN(n1319) );
XNOR2_X1 U1080 ( .A(G113), .B(n1373), .ZN(n1323) );
XOR2_X1 U1081 ( .A(KEYINPUT61), .B(G116), .Z(n1373) );
INV_X1 U1082 ( .A(n1071), .ZN(n1272) );
NAND2_X1 U1083 ( .A1(n1289), .A2(n1291), .ZN(n1071) );
XNOR2_X1 U1084 ( .A(KEYINPUT2), .B(n1267), .ZN(n1291) );
NAND2_X1 U1085 ( .A1(n1374), .A2(n1105), .ZN(n1267) );
NAND2_X1 U1086 ( .A1(G478), .A2(n1375), .ZN(n1105) );
NAND2_X1 U1087 ( .A1(n1175), .A2(n1300), .ZN(n1375) );
XOR2_X1 U1088 ( .A(KEYINPUT10), .B(n1118), .Z(n1374) );
NOR3_X1 U1089 ( .A1(G478), .A2(G902), .A3(n1376), .ZN(n1118) );
INV_X1 U1090 ( .A(n1175), .ZN(n1376) );
XNOR2_X1 U1091 ( .A(n1377), .B(n1378), .ZN(n1175) );
AND2_X1 U1092 ( .A1(n1307), .A2(G217), .ZN(n1378) );
AND2_X1 U1093 ( .A1(G234), .A2(n1126), .ZN(n1307) );
INV_X1 U1094 ( .A(G953), .ZN(n1126) );
NAND2_X1 U1095 ( .A1(n1379), .A2(KEYINPUT4), .ZN(n1377) );
XOR2_X1 U1096 ( .A(n1380), .B(n1381), .Z(n1379) );
XOR2_X1 U1097 ( .A(n1382), .B(n1383), .Z(n1381) );
XNOR2_X1 U1098 ( .A(n1384), .B(n1385), .ZN(n1383) );
NAND2_X1 U1099 ( .A1(KEYINPUT60), .A2(n1386), .ZN(n1385) );
INV_X1 U1100 ( .A(G143), .ZN(n1386) );
NAND2_X1 U1101 ( .A1(KEYINPUT55), .A2(n1370), .ZN(n1384) );
INV_X1 U1102 ( .A(G107), .ZN(n1370) );
NAND2_X1 U1103 ( .A1(KEYINPUT21), .A2(n1343), .ZN(n1382) );
INV_X1 U1104 ( .A(G134), .ZN(n1343) );
XNOR2_X1 U1105 ( .A(G116), .B(n1387), .ZN(n1380) );
XNOR2_X1 U1106 ( .A(n1277), .B(G122), .ZN(n1387) );
INV_X1 U1107 ( .A(G128), .ZN(n1277) );
INV_X1 U1108 ( .A(n1109), .ZN(n1289) );
XOR2_X1 U1109 ( .A(n1388), .B(n1181), .Z(n1109) );
INV_X1 U1110 ( .A(G475), .ZN(n1181) );
NAND2_X1 U1111 ( .A1(n1179), .A2(n1300), .ZN(n1388) );
INV_X1 U1112 ( .A(G902), .ZN(n1300) );
XOR2_X1 U1113 ( .A(G104), .B(n1389), .Z(n1179) );
XOR2_X1 U1114 ( .A(n1390), .B(n1391), .Z(n1389) );
XOR2_X1 U1115 ( .A(n1392), .B(n1393), .Z(n1391) );
XOR2_X1 U1116 ( .A(n1394), .B(n1395), .Z(n1393) );
NAND2_X1 U1117 ( .A1(KEYINPUT8), .A2(n1396), .ZN(n1395) );
INV_X1 U1118 ( .A(G113), .ZN(n1396) );
NAND2_X1 U1119 ( .A1(n1331), .A2(G214), .ZN(n1394) );
NOR2_X1 U1120 ( .A1(G953), .A2(G237), .ZN(n1331) );
XNOR2_X1 U1121 ( .A(n1367), .B(n1141), .ZN(n1392) );
XOR2_X1 U1122 ( .A(G140), .B(KEYINPUT53), .Z(n1141) );
XNOR2_X1 U1123 ( .A(G122), .B(n1227), .ZN(n1367) );
INV_X1 U1124 ( .A(G125), .ZN(n1227) );
XOR2_X1 U1125 ( .A(n1397), .B(n1398), .Z(n1390) );
XNOR2_X1 U1126 ( .A(KEYINPUT7), .B(n1261), .ZN(n1398) );
INV_X1 U1127 ( .A(G146), .ZN(n1261) );
XNOR2_X1 U1128 ( .A(G143), .B(G131), .ZN(n1397) );
endmodule


