//Key = 0100000111110110011010110011001100011001100001111111011011000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;

XOR2_X1 U732 ( .A(G107), .B(n1008), .Z(G9) );
NOR2_X1 U733 ( .A1(n1009), .A2(n1010), .ZN(G75) );
XOR2_X1 U734 ( .A(n1011), .B(KEYINPUT30), .Z(n1010) );
OR3_X1 U735 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
NOR2_X1 U736 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
AND2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND4_X1 U738 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NAND2_X1 U739 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
OR2_X1 U741 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U742 ( .A1(n1029), .A2(n1030), .ZN(n1023) );
NAND2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND3_X1 U745 ( .A1(n1029), .A2(n1035), .A3(n1025), .ZN(n1017) );
NAND2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U747 ( .A1(n1038), .A2(n1039), .A3(n1019), .ZN(n1037) );
OR2_X1 U748 ( .A1(n1022), .A2(n1020), .ZN(n1039) );
NAND3_X1 U749 ( .A1(n1040), .A2(n1041), .A3(n1022), .ZN(n1038) );
NAND2_X1 U750 ( .A1(n1042), .A2(n1020), .ZN(n1036) );
NOR2_X1 U751 ( .A1(G952), .A2(n1012), .ZN(n1009) );
NAND2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1012) );
NAND4_X1 U753 ( .A1(n1045), .A2(n1025), .A3(n1046), .A4(n1047), .ZN(n1044) );
NOR3_X1 U754 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
XOR2_X1 U755 ( .A(n1051), .B(KEYINPUT40), .Z(n1049) );
NAND3_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1022), .ZN(n1048) );
NOR3_X1 U757 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1046) );
NOR3_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
INV_X1 U759 ( .A(KEYINPUT47), .ZN(n1057) );
NOR2_X1 U760 ( .A1(KEYINPUT47), .A2(G475), .ZN(n1055) );
XOR2_X1 U761 ( .A(n1060), .B(n1061), .Z(n1054) );
XOR2_X1 U762 ( .A(n1062), .B(n1063), .Z(n1045) );
NOR2_X1 U763 ( .A1(KEYINPUT6), .A2(n1064), .ZN(n1063) );
XOR2_X1 U764 ( .A(n1065), .B(n1066), .Z(G72) );
XOR2_X1 U765 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U766 ( .A1(n1069), .A2(n1043), .ZN(n1068) );
AND2_X1 U767 ( .A1(G227), .A2(G900), .ZN(n1069) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
NAND2_X1 U769 ( .A1(G953), .A2(n1072), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1073), .B(n1074), .Z(n1070) );
XOR2_X1 U771 ( .A(n1075), .B(n1076), .Z(n1074) );
XNOR2_X1 U772 ( .A(n1077), .B(n1078), .ZN(n1073) );
NAND2_X1 U773 ( .A1(KEYINPUT61), .A2(n1079), .ZN(n1078) );
NAND2_X1 U774 ( .A1(KEYINPUT9), .A2(n1080), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1043), .A2(n1081), .ZN(n1065) );
NAND2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(G69) );
NAND2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
OR2_X1 U779 ( .A1(n1043), .A2(G224), .ZN(n1087) );
NAND3_X1 U780 ( .A1(n1088), .A2(n1089), .A3(G953), .ZN(n1084) );
NAND2_X1 U781 ( .A1(G898), .A2(G224), .ZN(n1089) );
XOR2_X1 U782 ( .A(KEYINPUT20), .B(n1086), .Z(n1088) );
XNOR2_X1 U783 ( .A(n1090), .B(n1091), .ZN(n1086) );
NOR2_X1 U784 ( .A1(n1092), .A2(G953), .ZN(n1091) );
NAND3_X1 U785 ( .A1(KEYINPUT7), .A2(n1093), .A3(n1094), .ZN(n1090) );
XOR2_X1 U786 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U787 ( .A1(KEYINPUT17), .A2(n1097), .ZN(n1095) );
NAND2_X1 U788 ( .A1(G953), .A2(n1098), .ZN(n1093) );
NOR2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XNOR2_X1 U790 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U792 ( .A1(n1099), .A2(n1105), .ZN(G63) );
XOR2_X1 U793 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U794 ( .A1(n1108), .A2(n1104), .ZN(n1107) );
INV_X1 U795 ( .A(G478), .ZN(n1108) );
NOR2_X1 U796 ( .A1(n1099), .A2(n1109), .ZN(G60) );
XOR2_X1 U797 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U798 ( .A1(n1059), .A2(n1104), .ZN(n1111) );
XOR2_X1 U799 ( .A(G104), .B(n1112), .Z(G6) );
NOR2_X1 U800 ( .A1(n1099), .A2(n1113), .ZN(G57) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND3_X1 U802 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1114) );
OR2_X1 U803 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND3_X1 U804 ( .A1(n1121), .A2(n1119), .A3(n1122), .ZN(n1117) );
INV_X1 U805 ( .A(KEYINPUT15), .ZN(n1119) );
OR2_X1 U806 ( .A1(n1122), .A2(n1121), .ZN(n1116) );
AND2_X1 U807 ( .A1(KEYINPUT13), .A2(n1120), .ZN(n1121) );
NOR2_X1 U808 ( .A1(n1104), .A2(n1062), .ZN(n1120) );
INV_X1 U809 ( .A(G472), .ZN(n1062) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U811 ( .A(n1125), .B(n1079), .Z(n1123) );
NOR2_X1 U812 ( .A1(n1099), .A2(n1126), .ZN(G54) );
XOR2_X1 U813 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U814 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U815 ( .A(n1131), .B(n1079), .Z(n1130) );
NOR2_X1 U816 ( .A1(n1132), .A2(n1104), .ZN(n1131) );
INV_X1 U817 ( .A(G469), .ZN(n1132) );
XOR2_X1 U818 ( .A(n1133), .B(n1134), .Z(n1127) );
XOR2_X1 U819 ( .A(n1135), .B(KEYINPUT45), .Z(n1134) );
NAND4_X1 U820 ( .A1(KEYINPUT35), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1133) );
NAND3_X1 U821 ( .A1(KEYINPUT50), .A2(n1139), .A3(n1140), .ZN(n1138) );
OR2_X1 U822 ( .A1(n1140), .A2(n1139), .ZN(n1137) );
NOR2_X1 U823 ( .A1(G110), .A2(KEYINPUT59), .ZN(n1139) );
INV_X1 U824 ( .A(G140), .ZN(n1140) );
NAND2_X1 U825 ( .A1(G110), .A2(n1141), .ZN(n1136) );
INV_X1 U826 ( .A(KEYINPUT50), .ZN(n1141) );
NOR2_X1 U827 ( .A1(n1142), .A2(G952), .ZN(n1099) );
NOR2_X1 U828 ( .A1(n1143), .A2(n1144), .ZN(G51) );
XOR2_X1 U829 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U830 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U831 ( .A1(n1061), .A2(n1104), .ZN(n1148) );
NAND2_X1 U832 ( .A1(G902), .A2(n1014), .ZN(n1104) );
NAND3_X1 U833 ( .A1(n1082), .A2(n1149), .A3(n1092), .ZN(n1014) );
AND4_X1 U834 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1092) );
NOR4_X1 U835 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NOR2_X1 U836 ( .A1(n1008), .A2(n1112), .ZN(n1152) );
AND3_X1 U837 ( .A1(n1158), .A2(n1020), .A3(n1028), .ZN(n1112) );
AND3_X1 U838 ( .A1(n1020), .A2(n1027), .A3(n1158), .ZN(n1008) );
NAND2_X1 U839 ( .A1(n1159), .A2(n1042), .ZN(n1150) );
XNOR2_X1 U840 ( .A(KEYINPUT8), .B(n1083), .ZN(n1149) );
AND4_X1 U841 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1082) );
NOR4_X1 U842 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
INV_X1 U843 ( .A(n1168), .ZN(n1167) );
INV_X1 U844 ( .A(n1169), .ZN(n1166) );
NAND3_X1 U845 ( .A1(n1027), .A2(n1170), .A3(n1171), .ZN(n1162) );
NAND3_X1 U846 ( .A1(n1028), .A2(n1172), .A3(n1173), .ZN(n1160) );
NOR2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(n1147) );
NOR2_X1 U848 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NOR2_X1 U849 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
AND2_X1 U850 ( .A1(n1180), .A2(KEYINPUT56), .ZN(n1178) );
NOR2_X1 U851 ( .A1(n1181), .A2(n1180), .ZN(n1174) );
XNOR2_X1 U852 ( .A(n1182), .B(KEYINPUT18), .ZN(n1180) );
NOR2_X1 U853 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
INV_X1 U854 ( .A(KEYINPUT56), .ZN(n1184) );
NOR2_X1 U855 ( .A1(n1185), .A2(n1179), .ZN(n1183) );
INV_X1 U856 ( .A(KEYINPUT1), .ZN(n1179) );
NAND2_X1 U857 ( .A1(KEYINPUT26), .A2(n1186), .ZN(n1145) );
NOR2_X1 U858 ( .A1(n1187), .A2(n1142), .ZN(n1143) );
XOR2_X1 U859 ( .A(KEYINPUT53), .B(G953), .Z(n1142) );
XOR2_X1 U860 ( .A(KEYINPUT25), .B(G952), .Z(n1187) );
XOR2_X1 U861 ( .A(G146), .B(n1188), .Z(G48) );
NOR2_X1 U862 ( .A1(KEYINPUT2), .A2(n1161), .ZN(n1188) );
NAND3_X1 U863 ( .A1(n1028), .A2(n1170), .A3(n1171), .ZN(n1161) );
XOR2_X1 U864 ( .A(n1189), .B(n1168), .Z(G45) );
NAND4_X1 U865 ( .A1(n1190), .A2(n1042), .A3(n1172), .A4(n1191), .ZN(n1168) );
AND3_X1 U866 ( .A1(n1050), .A2(n1192), .A3(n1170), .ZN(n1191) );
XOR2_X1 U867 ( .A(G140), .B(n1165), .Z(G42) );
AND3_X1 U868 ( .A1(n1193), .A2(n1028), .A3(n1173), .ZN(n1165) );
XOR2_X1 U869 ( .A(G137), .B(n1164), .Z(G39) );
AND3_X1 U870 ( .A1(n1194), .A2(n1029), .A3(n1173), .ZN(n1164) );
XNOR2_X1 U871 ( .A(G134), .B(n1083), .ZN(G36) );
NAND3_X1 U872 ( .A1(n1172), .A2(n1027), .A3(n1173), .ZN(n1083) );
AND4_X1 U873 ( .A1(n1019), .A2(n1190), .A3(n1170), .A4(n1022), .ZN(n1173) );
XOR2_X1 U874 ( .A(n1080), .B(n1195), .Z(G33) );
NAND4_X1 U875 ( .A1(n1028), .A2(n1172), .A3(n1019), .A4(n1196), .ZN(n1195) );
NOR3_X1 U876 ( .A1(n1031), .A2(n1197), .A3(n1198), .ZN(n1196) );
XOR2_X1 U877 ( .A(n1170), .B(KEYINPUT23), .Z(n1198) );
INV_X1 U878 ( .A(n1190), .ZN(n1031) );
NAND2_X1 U879 ( .A1(n1199), .A2(n1200), .ZN(G30) );
NAND2_X1 U880 ( .A1(G128), .A2(n1201), .ZN(n1200) );
XOR2_X1 U881 ( .A(n1202), .B(KEYINPUT34), .Z(n1199) );
OR2_X1 U882 ( .A1(n1201), .A2(G128), .ZN(n1202) );
NAND3_X1 U883 ( .A1(n1171), .A2(n1027), .A3(n1203), .ZN(n1201) );
XOR2_X1 U884 ( .A(n1170), .B(KEYINPUT55), .Z(n1203) );
AND3_X1 U885 ( .A1(n1190), .A2(n1042), .A3(n1194), .ZN(n1171) );
XOR2_X1 U886 ( .A(G101), .B(n1157), .Z(G3) );
AND3_X1 U887 ( .A1(n1172), .A2(n1029), .A3(n1158), .ZN(n1157) );
AND3_X1 U888 ( .A1(n1042), .A2(n1204), .A3(n1190), .ZN(n1158) );
XOR2_X1 U889 ( .A(n1205), .B(n1169), .Z(G27) );
NAND4_X1 U890 ( .A1(n1042), .A2(n1170), .A3(n1025), .A4(n1206), .ZN(n1169) );
AND2_X1 U891 ( .A1(n1028), .A2(n1193), .ZN(n1206) );
NAND2_X1 U892 ( .A1(n1015), .A2(n1207), .ZN(n1170) );
NAND4_X1 U893 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1072), .ZN(n1207) );
INV_X1 U894 ( .A(G900), .ZN(n1072) );
XOR2_X1 U895 ( .A(n1209), .B(n1151), .Z(G24) );
NAND4_X1 U896 ( .A1(n1210), .A2(n1020), .A3(n1050), .A4(n1192), .ZN(n1151) );
NAND2_X1 U897 ( .A1(n1211), .A2(n1212), .ZN(n1020) );
OR2_X1 U898 ( .A1(n1041), .A2(KEYINPUT49), .ZN(n1212) );
NAND3_X1 U899 ( .A1(n1213), .A2(n1214), .A3(KEYINPUT49), .ZN(n1211) );
XOR2_X1 U900 ( .A(G119), .B(n1156), .Z(G21) );
AND3_X1 U901 ( .A1(n1210), .A2(n1029), .A3(n1194), .ZN(n1156) );
AND2_X1 U902 ( .A1(n1215), .A2(n1216), .ZN(n1194) );
XOR2_X1 U903 ( .A(G116), .B(n1155), .Z(G18) );
AND3_X1 U904 ( .A1(n1172), .A2(n1027), .A3(n1210), .ZN(n1155) );
NAND2_X1 U905 ( .A1(n1217), .A2(n1218), .ZN(n1027) );
NAND3_X1 U906 ( .A1(n1219), .A2(n1050), .A3(n1220), .ZN(n1218) );
INV_X1 U907 ( .A(KEYINPUT28), .ZN(n1220) );
NAND2_X1 U908 ( .A1(KEYINPUT28), .A2(n1029), .ZN(n1217) );
XOR2_X1 U909 ( .A(n1154), .B(n1221), .Z(G15) );
NOR2_X1 U910 ( .A1(KEYINPUT37), .A2(n1222), .ZN(n1221) );
AND3_X1 U911 ( .A1(n1028), .A2(n1172), .A3(n1210), .ZN(n1154) );
AND3_X1 U912 ( .A1(n1042), .A2(n1204), .A3(n1025), .ZN(n1210) );
NOR2_X1 U913 ( .A1(n1223), .A2(n1033), .ZN(n1025) );
INV_X1 U914 ( .A(n1034), .ZN(n1223) );
INV_X1 U915 ( .A(n1041), .ZN(n1172) );
NAND2_X1 U916 ( .A1(n1215), .A2(n1213), .ZN(n1041) );
XNOR2_X1 U917 ( .A(n1216), .B(KEYINPUT41), .ZN(n1213) );
INV_X1 U918 ( .A(n1214), .ZN(n1215) );
NOR2_X1 U919 ( .A1(n1050), .A2(n1219), .ZN(n1028) );
INV_X1 U920 ( .A(n1192), .ZN(n1219) );
XOR2_X1 U921 ( .A(n1224), .B(n1225), .Z(G12) );
XNOR2_X1 U922 ( .A(G110), .B(KEYINPUT63), .ZN(n1225) );
NAND2_X1 U923 ( .A1(n1226), .A2(n1042), .ZN(n1224) );
NOR2_X1 U924 ( .A1(n1019), .A2(n1197), .ZN(n1042) );
INV_X1 U925 ( .A(n1022), .ZN(n1197) );
NAND2_X1 U926 ( .A1(G214), .A2(n1227), .ZN(n1022) );
XOR2_X1 U927 ( .A(n1060), .B(n1228), .Z(n1019) );
NOR2_X1 U928 ( .A1(KEYINPUT16), .A2(n1061), .ZN(n1228) );
NAND2_X1 U929 ( .A1(G210), .A2(n1227), .ZN(n1061) );
NAND2_X1 U930 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
INV_X1 U931 ( .A(G237), .ZN(n1229) );
NAND2_X1 U932 ( .A1(n1231), .A2(n1230), .ZN(n1060) );
XOR2_X1 U933 ( .A(n1232), .B(n1233), .Z(n1231) );
NOR2_X1 U934 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NOR3_X1 U935 ( .A1(KEYINPUT27), .A2(n1079), .A3(n1205), .ZN(n1235) );
AND2_X1 U936 ( .A1(n1185), .A2(KEYINPUT27), .ZN(n1234) );
INV_X1 U937 ( .A(n1177), .ZN(n1185) );
XNOR2_X1 U938 ( .A(n1205), .B(n1079), .ZN(n1177) );
INV_X1 U939 ( .A(n1236), .ZN(n1079) );
INV_X1 U940 ( .A(G125), .ZN(n1205) );
XNOR2_X1 U941 ( .A(n1186), .B(n1182), .ZN(n1232) );
NAND2_X1 U942 ( .A1(G224), .A2(n1043), .ZN(n1182) );
NAND2_X1 U943 ( .A1(n1237), .A2(n1238), .ZN(n1186) );
NAND2_X1 U944 ( .A1(n1096), .A2(n1239), .ZN(n1238) );
XOR2_X1 U945 ( .A(n1240), .B(KEYINPUT32), .Z(n1237) );
OR2_X1 U946 ( .A1(n1239), .A2(n1096), .ZN(n1240) );
XNOR2_X1 U947 ( .A(n1241), .B(G110), .ZN(n1096) );
NAND2_X1 U948 ( .A1(KEYINPUT39), .A2(G122), .ZN(n1241) );
INV_X1 U949 ( .A(n1097), .ZN(n1239) );
XOR2_X1 U950 ( .A(n1242), .B(n1243), .Z(n1097) );
XOR2_X1 U951 ( .A(KEYINPUT60), .B(n1244), .Z(n1243) );
NOR2_X1 U952 ( .A1(KEYINPUT42), .A2(n1245), .ZN(n1244) );
XNOR2_X1 U953 ( .A(n1246), .B(n1247), .ZN(n1242) );
XNOR2_X1 U954 ( .A(n1159), .B(KEYINPUT11), .ZN(n1226) );
AND4_X1 U955 ( .A1(n1193), .A2(n1029), .A3(n1190), .A4(n1204), .ZN(n1159) );
NAND2_X1 U956 ( .A1(n1015), .A2(n1248), .ZN(n1204) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1208), .A4(n1098), .ZN(n1248) );
INV_X1 U958 ( .A(G898), .ZN(n1098) );
NAND3_X1 U959 ( .A1(n1208), .A2(n1043), .A3(G952), .ZN(n1015) );
NAND2_X1 U960 ( .A1(G237), .A2(G234), .ZN(n1208) );
NOR2_X1 U961 ( .A1(n1034), .A2(n1033), .ZN(n1190) );
AND2_X1 U962 ( .A1(G221), .A2(n1249), .ZN(n1033) );
XOR2_X1 U963 ( .A(n1250), .B(G469), .Z(n1034) );
NAND2_X1 U964 ( .A1(n1251), .A2(n1230), .ZN(n1250) );
XNOR2_X1 U965 ( .A(n1129), .B(n1252), .ZN(n1251) );
XOR2_X1 U966 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U967 ( .A1(KEYINPUT29), .A2(n1236), .ZN(n1254) );
NOR2_X1 U968 ( .A1(KEYINPUT24), .A2(n1255), .ZN(n1253) );
XNOR2_X1 U969 ( .A(n1135), .B(n1256), .ZN(n1255) );
XOR2_X1 U970 ( .A(G140), .B(G110), .Z(n1256) );
NAND2_X1 U971 ( .A1(G227), .A2(n1043), .ZN(n1135) );
XNOR2_X1 U972 ( .A(n1125), .B(n1247), .ZN(n1129) );
XNOR2_X1 U973 ( .A(n1257), .B(n1258), .ZN(n1247) );
XOR2_X1 U974 ( .A(KEYINPUT36), .B(G107), .Z(n1258) );
XOR2_X1 U975 ( .A(n1259), .B(G104), .Z(n1257) );
INV_X1 U976 ( .A(G101), .ZN(n1259) );
NOR2_X1 U977 ( .A1(n1192), .A2(n1050), .ZN(n1029) );
XOR2_X1 U978 ( .A(G478), .B(n1260), .Z(n1050) );
NOR2_X1 U979 ( .A1(G902), .A2(n1106), .ZN(n1260) );
XOR2_X1 U980 ( .A(n1261), .B(n1262), .Z(n1106) );
NOR2_X1 U981 ( .A1(KEYINPUT58), .A2(n1263), .ZN(n1262) );
XOR2_X1 U982 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U983 ( .A(G122), .B(n1266), .Z(n1265) );
XOR2_X1 U984 ( .A(KEYINPUT31), .B(G134), .Z(n1266) );
XOR2_X1 U985 ( .A(n1267), .B(n1268), .Z(n1264) );
XOR2_X1 U986 ( .A(G116), .B(G107), .Z(n1268) );
NAND3_X1 U987 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1267) );
OR2_X1 U988 ( .A1(n1272), .A2(KEYINPUT14), .ZN(n1271) );
NAND3_X1 U989 ( .A1(KEYINPUT14), .A2(n1272), .A3(G143), .ZN(n1270) );
NAND2_X1 U990 ( .A1(n1273), .A2(n1189), .ZN(n1269) );
INV_X1 U991 ( .A(G143), .ZN(n1189) );
NAND2_X1 U992 ( .A1(n1274), .A2(KEYINPUT14), .ZN(n1273) );
XOR2_X1 U993 ( .A(n1272), .B(KEYINPUT21), .Z(n1274) );
NAND2_X1 U994 ( .A1(G217), .A2(n1275), .ZN(n1261) );
NAND2_X1 U995 ( .A1(n1052), .A2(n1276), .ZN(n1192) );
OR2_X1 U996 ( .A1(n1059), .A2(n1058), .ZN(n1276) );
NAND2_X1 U997 ( .A1(n1058), .A2(n1059), .ZN(n1052) );
INV_X1 U998 ( .A(G475), .ZN(n1059) );
NOR2_X1 U999 ( .A1(n1110), .A2(G902), .ZN(n1058) );
XOR2_X1 U1000 ( .A(n1277), .B(n1278), .Z(n1110) );
XOR2_X1 U1001 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U1002 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR3_X1 U1003 ( .A1(n1283), .A2(KEYINPUT5), .A3(n1284), .ZN(n1282) );
NOR2_X1 U1004 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XNOR2_X1 U1005 ( .A(n1287), .B(KEYINPUT10), .ZN(n1286) );
NOR2_X1 U1006 ( .A1(n1288), .A2(n1287), .ZN(n1285) );
NOR2_X1 U1007 ( .A1(G104), .A2(n1289), .ZN(n1288) );
NOR2_X1 U1008 ( .A1(n1290), .A2(n1291), .ZN(n1283) );
INV_X1 U1009 ( .A(G104), .ZN(n1291) );
NOR2_X1 U1010 ( .A1(n1287), .A2(n1289), .ZN(n1290) );
INV_X1 U1011 ( .A(KEYINPUT51), .ZN(n1289) );
AND2_X1 U1012 ( .A1(n1292), .A2(n1293), .ZN(n1287) );
NAND2_X1 U1013 ( .A1(G122), .A2(n1222), .ZN(n1293) );
INV_X1 U1014 ( .A(G113), .ZN(n1222) );
XOR2_X1 U1015 ( .A(n1294), .B(KEYINPUT0), .Z(n1292) );
NAND2_X1 U1016 ( .A1(G113), .A2(n1209), .ZN(n1294) );
INV_X1 U1017 ( .A(G122), .ZN(n1209) );
NAND2_X1 U1018 ( .A1(n1295), .A2(G214), .ZN(n1281) );
NAND2_X1 U1019 ( .A1(KEYINPUT48), .A2(n1080), .ZN(n1279) );
XNOR2_X1 U1020 ( .A(n1296), .B(n1076), .ZN(n1277) );
INV_X1 U1021 ( .A(n1040), .ZN(n1193) );
NAND2_X1 U1022 ( .A1(n1214), .A2(n1216), .ZN(n1040) );
NAND2_X1 U1023 ( .A1(n1051), .A2(n1053), .ZN(n1216) );
NAND3_X1 U1024 ( .A1(n1103), .A2(n1230), .A3(n1101), .ZN(n1053) );
NAND2_X1 U1025 ( .A1(n1297), .A2(n1298), .ZN(n1051) );
NAND2_X1 U1026 ( .A1(n1101), .A2(n1230), .ZN(n1298) );
XNOR2_X1 U1027 ( .A(n1299), .B(n1300), .ZN(n1101) );
XOR2_X1 U1028 ( .A(n1301), .B(n1302), .Z(n1300) );
NOR2_X1 U1029 ( .A1(KEYINPUT3), .A2(n1303), .ZN(n1302) );
NOR2_X1 U1030 ( .A1(n1304), .A2(n1305), .ZN(n1301) );
XOR2_X1 U1031 ( .A(n1306), .B(KEYINPUT46), .Z(n1305) );
NAND2_X1 U1032 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XOR2_X1 U1033 ( .A(n1309), .B(KEYINPUT43), .Z(n1307) );
NOR2_X1 U1034 ( .A1(n1309), .A2(n1308), .ZN(n1304) );
XOR2_X1 U1035 ( .A(n1310), .B(n1311), .Z(n1308) );
NOR2_X1 U1036 ( .A1(KEYINPUT38), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1037 ( .A(KEYINPUT12), .B(G128), .Z(n1312) );
XOR2_X1 U1038 ( .A(n1245), .B(G110), .Z(n1310) );
INV_X1 U1039 ( .A(G119), .ZN(n1245) );
XNOR2_X1 U1040 ( .A(G146), .B(n1076), .ZN(n1309) );
XOR2_X1 U1041 ( .A(G125), .B(G140), .Z(n1076) );
NAND2_X1 U1042 ( .A1(n1275), .A2(G221), .ZN(n1299) );
AND2_X1 U1043 ( .A1(G234), .A2(n1043), .ZN(n1275) );
INV_X1 U1044 ( .A(G953), .ZN(n1043) );
INV_X1 U1045 ( .A(n1103), .ZN(n1297) );
NAND2_X1 U1046 ( .A1(G217), .A2(n1249), .ZN(n1103) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1230), .ZN(n1249) );
XOR2_X1 U1048 ( .A(n1064), .B(G472), .Z(n1214) );
NAND2_X1 U1049 ( .A1(n1313), .A2(n1230), .ZN(n1064) );
INV_X1 U1050 ( .A(G902), .ZN(n1230) );
XOR2_X1 U1051 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1052 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1053 ( .A(n1318), .B(KEYINPUT44), .ZN(n1317) );
NAND2_X1 U1054 ( .A1(KEYINPUT54), .A2(n1236), .ZN(n1318) );
XOR2_X1 U1055 ( .A(n1272), .B(n1296), .Z(n1236) );
XOR2_X1 U1056 ( .A(G146), .B(G143), .Z(n1296) );
INV_X1 U1057 ( .A(G128), .ZN(n1272) );
XOR2_X1 U1058 ( .A(KEYINPUT62), .B(KEYINPUT57), .Z(n1316) );
XOR2_X1 U1059 ( .A(n1125), .B(n1319), .Z(n1314) );
XOR2_X1 U1060 ( .A(n1320), .B(n1321), .Z(n1319) );
INV_X1 U1061 ( .A(n1115), .ZN(n1321) );
XOR2_X1 U1062 ( .A(n1322), .B(G101), .Z(n1115) );
NAND2_X1 U1063 ( .A1(n1295), .A2(G210), .ZN(n1322) );
NOR2_X1 U1064 ( .A1(G953), .A2(G237), .ZN(n1295) );
NOR2_X1 U1065 ( .A1(KEYINPUT33), .A2(n1124), .ZN(n1320) );
XNOR2_X1 U1066 ( .A(G119), .B(n1246), .ZN(n1124) );
XOR2_X1 U1067 ( .A(G116), .B(G113), .Z(n1246) );
XOR2_X1 U1068 ( .A(n1323), .B(n1324), .Z(n1125) );
XOR2_X1 U1069 ( .A(KEYINPUT52), .B(KEYINPUT19), .Z(n1324) );
XOR2_X1 U1070 ( .A(n1325), .B(n1326), .Z(n1323) );
INV_X1 U1071 ( .A(n1075), .ZN(n1326) );
XNOR2_X1 U1072 ( .A(G134), .B(n1303), .ZN(n1075) );
XOR2_X1 U1073 ( .A(G137), .B(KEYINPUT4), .Z(n1303) );
NAND2_X1 U1074 ( .A1(KEYINPUT22), .A2(n1080), .ZN(n1325) );
INV_X1 U1075 ( .A(G131), .ZN(n1080) );
endmodule


