//Key = 1110101100101111100110111110011100100100101110101100010101010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275;

XNOR2_X1 U707 ( .A(G107), .B(n972), .ZN(G9) );
NOR2_X1 U708 ( .A1(n973), .A2(n974), .ZN(G75) );
NOR4_X1 U709 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .ZN(n974) );
NAND4_X1 U710 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(n975) );
NAND2_X1 U711 ( .A1(n983), .A2(n984), .ZN(n980) );
NAND3_X1 U712 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n979) );
NAND2_X1 U713 ( .A1(n988), .A2(n989), .ZN(n986) );
XNOR2_X1 U714 ( .A(n983), .B(KEYINPUT39), .ZN(n989) );
AND4_X1 U715 ( .A1(n990), .A2(n991), .A3(n992), .A4(n993), .ZN(n983) );
NAND2_X1 U716 ( .A1(n994), .A2(n995), .ZN(n985) );
NAND2_X1 U717 ( .A1(n996), .A2(n997), .ZN(n994) );
NAND2_X1 U718 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND3_X1 U719 ( .A1(n993), .A2(n1000), .A3(n1001), .ZN(n998) );
INV_X1 U720 ( .A(KEYINPUT61), .ZN(n1000) );
NAND3_X1 U721 ( .A1(n1002), .A2(n1003), .A3(n990), .ZN(n996) );
INV_X1 U722 ( .A(n999), .ZN(n990) );
NAND3_X1 U723 ( .A1(n992), .A2(n1004), .A3(n991), .ZN(n1003) );
NAND2_X1 U724 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U725 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND2_X1 U726 ( .A1(n993), .A2(n1009), .ZN(n1002) );
NAND4_X1 U727 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1009) );
NAND3_X1 U728 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
XNOR2_X1 U729 ( .A(n991), .B(KEYINPUT43), .ZN(n1016) );
NAND2_X1 U730 ( .A1(KEYINPUT61), .A2(n1001), .ZN(n1012) );
NAND2_X1 U731 ( .A1(n992), .A2(n1017), .ZN(n1011) );
NAND2_X1 U732 ( .A1(n991), .A2(n1018), .ZN(n1010) );
NOR3_X1 U733 ( .A1(n1019), .A2(G953), .A3(G952), .ZN(n973) );
INV_X1 U734 ( .A(n981), .ZN(n1019) );
NAND4_X1 U735 ( .A1(n987), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n981) );
NOR3_X1 U736 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
XNOR2_X1 U737 ( .A(n1007), .B(KEYINPUT24), .ZN(n1025) );
XOR2_X1 U738 ( .A(n1026), .B(KEYINPUT29), .Z(n1024) );
OR2_X1 U739 ( .A1(n1027), .A2(G472), .ZN(n1026) );
NAND3_X1 U740 ( .A1(n995), .A2(n1028), .A3(n1029), .ZN(n1023) );
NAND2_X1 U741 ( .A1(G472), .A2(n1027), .ZN(n1029) );
NOR3_X1 U742 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1021) );
AND3_X1 U743 ( .A1(KEYINPUT23), .A2(n1033), .A3(G475), .ZN(n1032) );
NOR2_X1 U744 ( .A1(KEYINPUT23), .A2(G475), .ZN(n1031) );
XOR2_X1 U745 ( .A(n1034), .B(n1035), .Z(G72) );
XOR2_X1 U746 ( .A(n1036), .B(n1037), .Z(n1035) );
NAND2_X1 U747 ( .A1(G953), .A2(n1038), .ZN(n1037) );
NAND2_X1 U748 ( .A1(G900), .A2(G227), .ZN(n1038) );
NAND2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1036) );
NAND2_X1 U750 ( .A1(n1041), .A2(G953), .ZN(n1040) );
XOR2_X1 U751 ( .A(n1042), .B(n1043), .Z(n1039) );
XOR2_X1 U752 ( .A(n1044), .B(n1045), .Z(n1043) );
NOR2_X1 U753 ( .A1(KEYINPUT51), .A2(n1046), .ZN(n1045) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
XOR2_X1 U755 ( .A(n1049), .B(KEYINPUT10), .Z(n1048) );
INV_X1 U756 ( .A(n1050), .ZN(n1047) );
NAND2_X1 U757 ( .A1(KEYINPUT6), .A2(n1051), .ZN(n1042) );
AND2_X1 U758 ( .A1(n976), .A2(n982), .ZN(n1034) );
XOR2_X1 U759 ( .A(n1052), .B(n1053), .Z(G69) );
XOR2_X1 U760 ( .A(n1054), .B(n1055), .Z(n1053) );
NOR2_X1 U761 ( .A1(G953), .A2(n1056), .ZN(n1055) );
XOR2_X1 U762 ( .A(KEYINPUT38), .B(n1057), .Z(n1056) );
NOR2_X1 U763 ( .A1(n1058), .A2(n978), .ZN(n1057) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(n1054) );
XOR2_X1 U765 ( .A(KEYINPUT41), .B(n1061), .Z(n1060) );
NOR2_X1 U766 ( .A1(G898), .A2(n982), .ZN(n1061) );
XOR2_X1 U767 ( .A(n1062), .B(n1063), .Z(n1059) );
XNOR2_X1 U768 ( .A(n1064), .B(n1065), .ZN(n1063) );
XOR2_X1 U769 ( .A(n1066), .B(n1067), .Z(n1062) );
XNOR2_X1 U770 ( .A(KEYINPUT54), .B(KEYINPUT19), .ZN(n1066) );
NOR2_X1 U771 ( .A1(n1068), .A2(n982), .ZN(n1052) );
AND2_X1 U772 ( .A1(G224), .A2(G898), .ZN(n1068) );
NOR2_X1 U773 ( .A1(n1069), .A2(n1070), .ZN(G66) );
XOR2_X1 U774 ( .A(n1071), .B(n1072), .Z(n1070) );
NOR2_X1 U775 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U776 ( .A1(KEYINPUT31), .A2(n1075), .ZN(n1071) );
NOR2_X1 U777 ( .A1(n1069), .A2(n1076), .ZN(G63) );
XOR2_X1 U778 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND2_X1 U779 ( .A1(n1079), .A2(G478), .ZN(n1077) );
NOR2_X1 U780 ( .A1(n1069), .A2(n1080), .ZN(G60) );
XOR2_X1 U781 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U782 ( .A1(n1079), .A2(G475), .ZN(n1081) );
XOR2_X1 U783 ( .A(n1083), .B(G104), .Z(G6) );
NAND2_X1 U784 ( .A1(KEYINPUT53), .A2(n1084), .ZN(n1083) );
NOR2_X1 U785 ( .A1(n1069), .A2(n1085), .ZN(G57) );
XOR2_X1 U786 ( .A(n1086), .B(n1087), .Z(n1085) );
XOR2_X1 U787 ( .A(n1088), .B(n1089), .Z(n1086) );
NOR2_X1 U788 ( .A1(n1090), .A2(n1074), .ZN(n1089) );
NAND2_X1 U789 ( .A1(KEYINPUT0), .A2(n1091), .ZN(n1088) );
NOR2_X1 U790 ( .A1(n1069), .A2(n1092), .ZN(G54) );
XNOR2_X1 U791 ( .A(n1093), .B(n1094), .ZN(n1092) );
XOR2_X1 U792 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR3_X1 U793 ( .A1(n1097), .A2(KEYINPUT33), .A3(n1098), .ZN(n1096) );
NAND2_X1 U794 ( .A1(n1079), .A2(G469), .ZN(n1095) );
INV_X1 U795 ( .A(n1074), .ZN(n1079) );
NOR2_X1 U796 ( .A1(n1069), .A2(n1099), .ZN(G51) );
XOR2_X1 U797 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U798 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U799 ( .A(n1104), .B(n1105), .Z(n1100) );
NOR2_X1 U800 ( .A1(n1106), .A2(n1074), .ZN(n1105) );
NAND2_X1 U801 ( .A1(G902), .A2(n1107), .ZN(n1074) );
OR3_X1 U802 ( .A1(n978), .A2(n977), .A3(n976), .ZN(n1107) );
NAND4_X1 U803 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n976) );
NOR4_X1 U804 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1111) );
INV_X1 U805 ( .A(n1116), .ZN(n1115) );
AND2_X1 U806 ( .A1(n1117), .A2(n1118), .ZN(n1110) );
XNOR2_X1 U807 ( .A(n1058), .B(KEYINPUT13), .ZN(n977) );
NAND4_X1 U808 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n978) );
NOR4_X1 U809 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1122) );
INV_X1 U810 ( .A(n972), .ZN(n1126) );
NAND4_X1 U811 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n993), .ZN(n972) );
INV_X1 U812 ( .A(n1084), .ZN(n1125) );
NAND4_X1 U813 ( .A1(n1127), .A2(n993), .A3(n1129), .A4(n1017), .ZN(n1084) );
INV_X1 U814 ( .A(n1130), .ZN(n993) );
XNOR2_X1 U815 ( .A(n1131), .B(n1132), .ZN(n1104) );
AND2_X1 U816 ( .A1(G953), .A2(n1133), .ZN(n1069) );
XOR2_X1 U817 ( .A(KEYINPUT15), .B(G952), .Z(n1133) );
XNOR2_X1 U818 ( .A(G146), .B(n1134), .ZN(G48) );
NAND2_X1 U819 ( .A1(KEYINPUT44), .A2(n1114), .ZN(n1134) );
AND4_X1 U820 ( .A1(n1135), .A2(n1018), .A3(n1017), .A4(n1136), .ZN(n1114) );
XNOR2_X1 U821 ( .A(G143), .B(n1108), .ZN(G45) );
NAND4_X1 U822 ( .A1(n1018), .A2(n984), .A3(n1137), .A4(n1138), .ZN(n1108) );
AND3_X1 U823 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
XOR2_X1 U824 ( .A(G140), .B(n1142), .Z(G42) );
NOR2_X1 U825 ( .A1(KEYINPUT3), .A2(n1109), .ZN(n1142) );
NAND4_X1 U826 ( .A1(n1143), .A2(n1017), .A3(n1007), .A4(n1008), .ZN(n1109) );
XNOR2_X1 U827 ( .A(G137), .B(n1118), .ZN(G39) );
NAND4_X1 U828 ( .A1(n1143), .A2(n991), .A3(n1136), .A4(n1007), .ZN(n1118) );
XNOR2_X1 U829 ( .A(G134), .B(n1117), .ZN(G36) );
NAND3_X1 U830 ( .A1(n1137), .A2(n1128), .A3(n1143), .ZN(n1117) );
XNOR2_X1 U831 ( .A(n1113), .B(n1144), .ZN(G33) );
NAND2_X1 U832 ( .A1(KEYINPUT49), .A2(G131), .ZN(n1144) );
AND3_X1 U833 ( .A1(n1137), .A2(n1017), .A3(n1143), .ZN(n1113) );
AND4_X1 U834 ( .A1(n987), .A2(n1018), .A3(n1141), .A4(n995), .ZN(n1143) );
NAND2_X1 U835 ( .A1(n1145), .A2(n1146), .ZN(G30) );
NAND2_X1 U836 ( .A1(n1112), .A2(n1147), .ZN(n1146) );
XOR2_X1 U837 ( .A(KEYINPUT40), .B(n1148), .Z(n1145) );
NOR2_X1 U838 ( .A1(n1112), .A2(n1147), .ZN(n1148) );
AND4_X1 U839 ( .A1(n1135), .A2(n1128), .A3(n1129), .A4(n1136), .ZN(n1112) );
XNOR2_X1 U840 ( .A(G101), .B(n1121), .ZN(G3) );
NAND4_X1 U841 ( .A1(n1137), .A2(n991), .A3(n1129), .A4(n1127), .ZN(n1121) );
XNOR2_X1 U842 ( .A(G125), .B(n1116), .ZN(G27) );
NAND4_X1 U843 ( .A1(n1135), .A2(n992), .A3(n1017), .A4(n1008), .ZN(n1116) );
AND3_X1 U844 ( .A1(n1007), .A2(n1141), .A3(n984), .ZN(n1135) );
NAND2_X1 U845 ( .A1(n999), .A2(n1149), .ZN(n1141) );
NAND4_X1 U846 ( .A1(n1041), .A2(G953), .A3(G902), .A4(n1150), .ZN(n1149) );
XNOR2_X1 U847 ( .A(G900), .B(KEYINPUT35), .ZN(n1041) );
XNOR2_X1 U848 ( .A(G122), .B(n1119), .ZN(G24) );
NAND3_X1 U849 ( .A1(n992), .A2(n1127), .A3(n1151), .ZN(n1119) );
NOR3_X1 U850 ( .A1(n1130), .A2(n1152), .A3(n1020), .ZN(n1151) );
NAND2_X1 U851 ( .A1(n1153), .A2(n1008), .ZN(n1130) );
XOR2_X1 U852 ( .A(n1124), .B(n1154), .Z(G21) );
NOR2_X1 U853 ( .A1(KEYINPUT58), .A2(n1155), .ZN(n1154) );
AND3_X1 U854 ( .A1(n992), .A2(n1136), .A3(n1156), .ZN(n1124) );
XOR2_X1 U855 ( .A(G116), .B(n1058), .Z(G18) );
AND3_X1 U856 ( .A1(n1137), .A2(n1127), .A3(n1001), .ZN(n1058) );
AND2_X1 U857 ( .A1(n992), .A2(n1128), .ZN(n1001) );
NOR2_X1 U858 ( .A1(n1140), .A2(n1020), .ZN(n1128) );
INV_X1 U859 ( .A(n1139), .ZN(n1020) );
XNOR2_X1 U860 ( .A(n1157), .B(n1158), .ZN(G15) );
NOR2_X1 U861 ( .A1(KEYINPUT63), .A2(n1120), .ZN(n1158) );
NAND4_X1 U862 ( .A1(n1137), .A2(n992), .A3(n1127), .A4(n1017), .ZN(n1120) );
NAND2_X1 U863 ( .A1(n1159), .A2(n1160), .ZN(n1017) );
OR3_X1 U864 ( .A1(n1139), .A2(n1152), .A3(KEYINPUT56), .ZN(n1160) );
INV_X1 U865 ( .A(n1140), .ZN(n1152) );
NAND2_X1 U866 ( .A1(KEYINPUT56), .A2(n991), .ZN(n1159) );
INV_X1 U867 ( .A(n1030), .ZN(n992) );
NAND2_X1 U868 ( .A1(n1014), .A2(n1161), .ZN(n1030) );
INV_X1 U869 ( .A(n1005), .ZN(n1137) );
NAND2_X1 U870 ( .A1(n1136), .A2(n1153), .ZN(n1005) );
XNOR2_X1 U871 ( .A(n1162), .B(KEYINPUT1), .ZN(n1153) );
INV_X1 U872 ( .A(n1007), .ZN(n1162) );
XNOR2_X1 U873 ( .A(n1008), .B(KEYINPUT9), .ZN(n1136) );
XNOR2_X1 U874 ( .A(G110), .B(n1163), .ZN(G12) );
NAND2_X1 U875 ( .A1(KEYINPUT55), .A2(n1123), .ZN(n1163) );
AND3_X1 U876 ( .A1(n1129), .A2(n1008), .A3(n1156), .ZN(n1123) );
AND3_X1 U877 ( .A1(n1127), .A2(n1007), .A3(n991), .ZN(n1156) );
NOR2_X1 U878 ( .A1(n1139), .A2(n1140), .ZN(n991) );
NAND3_X1 U879 ( .A1(n1164), .A2(n1165), .A3(n1028), .ZN(n1140) );
NAND2_X1 U880 ( .A1(n1166), .A2(n1167), .ZN(n1028) );
OR3_X1 U881 ( .A1(n1167), .A2(n1166), .A3(KEYINPUT36), .ZN(n1165) );
INV_X1 U882 ( .A(n1033), .ZN(n1166) );
NAND2_X1 U883 ( .A1(n1082), .A2(n1168), .ZN(n1033) );
XOR2_X1 U884 ( .A(n1169), .B(n1170), .Z(n1082) );
XOR2_X1 U885 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U886 ( .A(G122), .B(n1157), .ZN(n1172) );
XOR2_X1 U887 ( .A(KEYINPUT5), .B(G131), .Z(n1171) );
XNOR2_X1 U888 ( .A(n1173), .B(n1174), .ZN(n1169) );
INV_X1 U889 ( .A(n1175), .ZN(n1174) );
XOR2_X1 U890 ( .A(n1176), .B(n1177), .Z(n1173) );
NOR2_X1 U891 ( .A1(G104), .A2(KEYINPUT8), .ZN(n1177) );
NAND2_X1 U892 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
NAND4_X1 U893 ( .A1(n1180), .A2(G214), .A3(n1181), .A4(n982), .ZN(n1179) );
NAND2_X1 U894 ( .A1(n1182), .A2(n1183), .ZN(n1178) );
NAND3_X1 U895 ( .A1(n1181), .A2(n982), .A3(G214), .ZN(n1183) );
XNOR2_X1 U896 ( .A(KEYINPUT28), .B(n1180), .ZN(n1182) );
XOR2_X1 U897 ( .A(n1184), .B(KEYINPUT22), .Z(n1180) );
NAND2_X1 U898 ( .A1(KEYINPUT36), .A2(n1167), .ZN(n1164) );
INV_X1 U899 ( .A(G475), .ZN(n1167) );
XNOR2_X1 U900 ( .A(n1185), .B(G478), .ZN(n1139) );
NAND2_X1 U901 ( .A1(n1078), .A2(n1168), .ZN(n1185) );
XOR2_X1 U902 ( .A(n1186), .B(n1187), .Z(n1078) );
XOR2_X1 U903 ( .A(n1188), .B(n1189), .Z(n1187) );
XNOR2_X1 U904 ( .A(n1190), .B(n1191), .ZN(n1189) );
NAND2_X1 U905 ( .A1(G217), .A2(n1192), .ZN(n1190) );
NAND2_X1 U906 ( .A1(KEYINPUT34), .A2(n1193), .ZN(n1188) );
INV_X1 U907 ( .A(G134), .ZN(n1193) );
XOR2_X1 U908 ( .A(n1194), .B(n1195), .Z(n1186) );
XNOR2_X1 U909 ( .A(n1184), .B(G128), .ZN(n1195) );
XNOR2_X1 U910 ( .A(G116), .B(G122), .ZN(n1194) );
XOR2_X1 U911 ( .A(n1196), .B(n1073), .Z(n1007) );
NAND2_X1 U912 ( .A1(G217), .A2(n1197), .ZN(n1073) );
NAND2_X1 U913 ( .A1(n1075), .A2(n1168), .ZN(n1196) );
XOR2_X1 U914 ( .A(n1198), .B(n1199), .Z(n1075) );
XOR2_X1 U915 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND2_X1 U916 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U917 ( .A(KEYINPUT2), .B(n1204), .ZN(n1203) );
XOR2_X1 U918 ( .A(KEYINPUT42), .B(KEYINPUT32), .Z(n1202) );
NAND2_X1 U919 ( .A1(KEYINPUT14), .A2(n1205), .ZN(n1200) );
XOR2_X1 U920 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U921 ( .A(n1175), .B(G110), .ZN(n1207) );
XOR2_X1 U922 ( .A(G146), .B(n1051), .Z(n1175) );
XNOR2_X1 U923 ( .A(n1131), .B(G140), .ZN(n1051) );
XNOR2_X1 U924 ( .A(G119), .B(G128), .ZN(n1206) );
NAND2_X1 U925 ( .A1(G221), .A2(n1192), .ZN(n1198) );
AND2_X1 U926 ( .A1(G234), .A2(n982), .ZN(n1192) );
AND2_X1 U927 ( .A1(n984), .A2(n1208), .ZN(n1127) );
NAND2_X1 U928 ( .A1(n999), .A2(n1209), .ZN(n1208) );
NAND4_X1 U929 ( .A1(G953), .A2(G902), .A3(n1150), .A4(n1210), .ZN(n1209) );
INV_X1 U930 ( .A(G898), .ZN(n1210) );
NAND3_X1 U931 ( .A1(n1150), .A2(n982), .A3(G952), .ZN(n999) );
NAND2_X1 U932 ( .A1(G237), .A2(G234), .ZN(n1150) );
NOR2_X1 U933 ( .A1(n987), .A2(n988), .ZN(n984) );
INV_X1 U934 ( .A(n995), .ZN(n988) );
NAND2_X1 U935 ( .A1(G214), .A2(n1211), .ZN(n995) );
XNOR2_X1 U936 ( .A(n1212), .B(n1106), .ZN(n987) );
NAND2_X1 U937 ( .A1(G210), .A2(n1211), .ZN(n1106) );
NAND2_X1 U938 ( .A1(n1181), .A2(n1168), .ZN(n1211) );
NAND2_X1 U939 ( .A1(n1213), .A2(n1168), .ZN(n1212) );
XOR2_X1 U940 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U941 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U942 ( .A(KEYINPUT60), .B(KEYINPUT30), .Z(n1217) );
NOR2_X1 U943 ( .A1(KEYINPUT17), .A2(n1132), .ZN(n1216) );
NAND2_X1 U944 ( .A1(G224), .A2(n982), .ZN(n1132) );
XOR2_X1 U945 ( .A(n1218), .B(n1103), .Z(n1214) );
XNOR2_X1 U946 ( .A(n1219), .B(n1067), .ZN(n1103) );
XNOR2_X1 U947 ( .A(n1220), .B(G122), .ZN(n1067) );
XNOR2_X1 U948 ( .A(KEYINPUT27), .B(n1221), .ZN(n1219) );
NOR2_X1 U949 ( .A1(KEYINPUT50), .A2(n1222), .ZN(n1221) );
XNOR2_X1 U950 ( .A(n1065), .B(n1223), .ZN(n1222) );
NOR2_X1 U951 ( .A1(KEYINPUT52), .A2(n1064), .ZN(n1223) );
XNOR2_X1 U952 ( .A(n1224), .B(n1225), .ZN(n1064) );
NAND2_X1 U953 ( .A1(KEYINPUT16), .A2(n1157), .ZN(n1224) );
INV_X1 U954 ( .A(G113), .ZN(n1157) );
XOR2_X1 U955 ( .A(G101), .B(n1226), .Z(n1065) );
XNOR2_X1 U956 ( .A(n1191), .B(G104), .ZN(n1226) );
NAND2_X1 U957 ( .A1(n1227), .A2(n1228), .ZN(n1218) );
NAND2_X1 U958 ( .A1(n1229), .A2(n1131), .ZN(n1228) );
INV_X1 U959 ( .A(G125), .ZN(n1131) );
XOR2_X1 U960 ( .A(KEYINPUT4), .B(n1102), .Z(n1229) );
NAND2_X1 U961 ( .A1(G125), .A2(n1230), .ZN(n1227) );
XNOR2_X1 U962 ( .A(n1102), .B(KEYINPUT59), .ZN(n1230) );
NAND3_X1 U963 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1008) );
OR2_X1 U964 ( .A1(n1090), .A2(n1234), .ZN(n1233) );
NAND3_X1 U965 ( .A1(n1234), .A2(n1090), .A3(KEYINPUT7), .ZN(n1232) );
INV_X1 U966 ( .A(G472), .ZN(n1090) );
NOR2_X1 U967 ( .A1(KEYINPUT21), .A2(n1235), .ZN(n1234) );
NAND2_X1 U968 ( .A1(n1235), .A2(n1236), .ZN(n1231) );
INV_X1 U969 ( .A(KEYINPUT7), .ZN(n1236) );
XOR2_X1 U970 ( .A(n1027), .B(KEYINPUT48), .Z(n1235) );
NAND2_X1 U971 ( .A1(n1237), .A2(n1168), .ZN(n1027) );
XOR2_X1 U972 ( .A(n1087), .B(n1238), .Z(n1237) );
XNOR2_X1 U973 ( .A(KEYINPUT25), .B(n1091), .ZN(n1238) );
XNOR2_X1 U974 ( .A(n1102), .B(n1239), .ZN(n1091) );
XNOR2_X1 U975 ( .A(n1240), .B(n1241), .ZN(n1102) );
NOR2_X1 U976 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U977 ( .A(n1244), .B(KEYINPUT37), .Z(n1243) );
NAND2_X1 U978 ( .A1(KEYINPUT46), .A2(n1147), .ZN(n1240) );
INV_X1 U979 ( .A(G128), .ZN(n1147) );
XOR2_X1 U980 ( .A(n1245), .B(n1246), .Z(n1087) );
XNOR2_X1 U981 ( .A(n1247), .B(n1248), .ZN(n1246) );
AND3_X1 U982 ( .A1(G210), .A2(n982), .A3(n1181), .ZN(n1248) );
INV_X1 U983 ( .A(G237), .ZN(n1181) );
XNOR2_X1 U984 ( .A(G113), .B(n1225), .ZN(n1245) );
XNOR2_X1 U985 ( .A(G116), .B(n1155), .ZN(n1225) );
INV_X1 U986 ( .A(G119), .ZN(n1155) );
XNOR2_X1 U987 ( .A(n1018), .B(KEYINPUT26), .ZN(n1129) );
NOR2_X1 U988 ( .A1(n1014), .A2(n1015), .ZN(n1018) );
INV_X1 U989 ( .A(n1161), .ZN(n1015) );
NAND2_X1 U990 ( .A1(G221), .A2(n1249), .ZN(n1161) );
XNOR2_X1 U991 ( .A(KEYINPUT20), .B(n1197), .ZN(n1249) );
NAND2_X1 U992 ( .A1(G234), .A2(n1168), .ZN(n1197) );
XOR2_X1 U993 ( .A(n1250), .B(G469), .Z(n1014) );
NAND2_X1 U994 ( .A1(n1251), .A2(n1168), .ZN(n1250) );
INV_X1 U995 ( .A(G902), .ZN(n1168) );
XOR2_X1 U996 ( .A(n1252), .B(n1253), .Z(n1251) );
NOR2_X1 U997 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
AND2_X1 U998 ( .A1(KEYINPUT11), .A2(n1098), .ZN(n1255) );
NOR3_X1 U999 ( .A1(KEYINPUT11), .A2(n1098), .A3(n1097), .ZN(n1254) );
AND2_X1 U1000 ( .A1(n1256), .A2(n1257), .ZN(n1097) );
NAND2_X1 U1001 ( .A1(G227), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U1002 ( .A(G140), .B(n1220), .ZN(n1256) );
INV_X1 U1003 ( .A(G110), .ZN(n1220) );
AND3_X1 U1004 ( .A1(G227), .A2(n1258), .A3(n1259), .ZN(n1098) );
XNOR2_X1 U1005 ( .A(G110), .B(G140), .ZN(n1259) );
XNOR2_X1 U1006 ( .A(KEYINPUT57), .B(n982), .ZN(n1258) );
INV_X1 U1007 ( .A(G953), .ZN(n982) );
NAND2_X1 U1008 ( .A1(n1260), .A2(n1261), .ZN(n1252) );
NAND2_X1 U1009 ( .A1(n1093), .A2(n1262), .ZN(n1261) );
XOR2_X1 U1010 ( .A(n1239), .B(n1263), .Z(n1093) );
OR3_X1 U1011 ( .A1(n1263), .A2(n1239), .A3(n1262), .ZN(n1260) );
INV_X1 U1012 ( .A(KEYINPUT47), .ZN(n1262) );
XNOR2_X1 U1013 ( .A(n1264), .B(KEYINPUT62), .ZN(n1239) );
NAND2_X1 U1014 ( .A1(n1049), .A2(n1050), .ZN(n1264) );
NAND2_X1 U1015 ( .A1(G131), .A2(n1265), .ZN(n1050) );
OR2_X1 U1016 ( .A1(n1265), .A2(G131), .ZN(n1049) );
XNOR2_X1 U1017 ( .A(G134), .B(n1204), .ZN(n1265) );
INV_X1 U1018 ( .A(G137), .ZN(n1204) );
XNOR2_X1 U1019 ( .A(n1266), .B(n1046), .ZN(n1263) );
XNOR2_X1 U1020 ( .A(n1267), .B(G128), .ZN(n1046) );
NAND2_X1 U1021 ( .A1(n1268), .A2(n1244), .ZN(n1267) );
NAND2_X1 U1022 ( .A1(n1269), .A2(n1270), .ZN(n1244) );
INV_X1 U1023 ( .A(G146), .ZN(n1270) );
XNOR2_X1 U1024 ( .A(KEYINPUT45), .B(n1184), .ZN(n1269) );
INV_X1 U1025 ( .A(G143), .ZN(n1184) );
XNOR2_X1 U1026 ( .A(n1242), .B(KEYINPUT18), .ZN(n1268) );
AND2_X1 U1027 ( .A1(n1271), .A2(G146), .ZN(n1242) );
XNOR2_X1 U1028 ( .A(KEYINPUT45), .B(G143), .ZN(n1271) );
XNOR2_X1 U1029 ( .A(n1272), .B(n1247), .ZN(n1266) );
INV_X1 U1030 ( .A(G101), .ZN(n1247) );
NAND2_X1 U1031 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U1032 ( .A1(G104), .A2(n1191), .ZN(n1274) );
XOR2_X1 U1033 ( .A(KEYINPUT12), .B(n1275), .Z(n1273) );
NOR2_X1 U1034 ( .A1(G104), .A2(n1191), .ZN(n1275) );
INV_X1 U1035 ( .A(G107), .ZN(n1191) );
endmodule


