//Key = 1111111100100010110011101101001100001100001100111101110011110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;

XOR2_X1 U745 ( .A(G107), .B(n1043), .Z(G9) );
NOR2_X1 U746 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U747 ( .A1(KEYINPUT50), .A2(n1046), .ZN(n1045) );
NOR2_X1 U748 ( .A1(KEYINPUT56), .A2(n1047), .ZN(n1044) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(G75) );
NOR4_X1 U750 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
NAND3_X1 U751 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1050) );
NAND2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U753 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND2_X1 U754 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U755 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U756 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND2_X1 U757 ( .A1(n1068), .A2(n1069), .ZN(n1063) );
NAND3_X1 U758 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U759 ( .A1(n1073), .A2(n1066), .ZN(n1072) );
XOR2_X1 U760 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U761 ( .A1(KEYINPUT12), .A2(n1076), .ZN(n1075) );
NAND3_X1 U762 ( .A1(n1065), .A2(n1077), .A3(KEYINPUT0), .ZN(n1070) );
NAND2_X1 U763 ( .A1(n1078), .A2(n1079), .ZN(n1059) );
INV_X1 U764 ( .A(KEYINPUT0), .ZN(n1079) );
NAND4_X1 U765 ( .A1(n1061), .A2(n1065), .A3(n1077), .A4(n1068), .ZN(n1078) );
NAND3_X1 U766 ( .A1(n1066), .A2(n1080), .A3(n1065), .ZN(n1054) );
NAND2_X1 U767 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U768 ( .A1(n1083), .A2(n1057), .A3(n1084), .ZN(n1082) );
XOR2_X1 U769 ( .A(n1085), .B(KEYINPUT57), .Z(n1084) );
NAND2_X1 U770 ( .A1(n1068), .A2(n1086), .ZN(n1081) );
NAND2_X1 U771 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U772 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
XOR2_X1 U773 ( .A(n1085), .B(KEYINPUT21), .Z(n1091) );
NAND2_X1 U774 ( .A1(n1061), .A2(n1092), .ZN(n1087) );
INV_X1 U775 ( .A(n1085), .ZN(n1061) );
NOR3_X1 U776 ( .A1(n1052), .A2(G952), .A3(n1093), .ZN(n1048) );
INV_X1 U777 ( .A(n1055), .ZN(n1093) );
NAND4_X1 U778 ( .A1(n1094), .A2(n1066), .A3(n1095), .A4(n1096), .ZN(n1055) );
NOR3_X1 U779 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
XNOR2_X1 U780 ( .A(n1100), .B(n1101), .ZN(n1095) );
NOR2_X1 U781 ( .A1(KEYINPUT54), .A2(n1102), .ZN(n1101) );
XOR2_X1 U782 ( .A(n1103), .B(G469), .Z(n1094) );
XOR2_X1 U783 ( .A(n1104), .B(n1105), .Z(G72) );
XOR2_X1 U784 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U785 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
AND2_X1 U786 ( .A1(G227), .A2(G900), .ZN(n1108) );
NOR2_X1 U787 ( .A1(n1110), .A2(n1111), .ZN(n1106) );
XOR2_X1 U788 ( .A(n1112), .B(KEYINPUT62), .Z(n1111) );
NAND2_X1 U789 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NAND3_X1 U790 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
XOR2_X1 U791 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U792 ( .A1(G125), .A2(KEYINPUT39), .ZN(n1118) );
NAND2_X1 U793 ( .A1(n1120), .A2(n1121), .ZN(n1113) );
NAND2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1121) );
INV_X1 U795 ( .A(KEYINPUT40), .ZN(n1116) );
INV_X1 U796 ( .A(G140), .ZN(n1115) );
XOR2_X1 U797 ( .A(n1122), .B(n1119), .Z(n1120) );
XNOR2_X1 U798 ( .A(n1123), .B(n1124), .ZN(n1119) );
XOR2_X1 U799 ( .A(KEYINPUT33), .B(G131), .Z(n1124) );
NOR2_X1 U800 ( .A1(KEYINPUT39), .A2(n1125), .ZN(n1122) );
NOR2_X1 U801 ( .A1(n1126), .A2(G953), .ZN(n1104) );
NAND3_X1 U802 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(G69) );
XOR2_X1 U803 ( .A(n1130), .B(KEYINPUT9), .Z(n1129) );
OR2_X1 U804 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U805 ( .A1(n1132), .A2(n1131), .ZN(n1128) );
NAND2_X1 U806 ( .A1(G953), .A2(n1133), .ZN(n1131) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1133) );
NOR2_X1 U808 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
XNOR2_X1 U809 ( .A(KEYINPUT42), .B(n1136), .ZN(n1135) );
NAND2_X1 U810 ( .A1(n1136), .A2(n1134), .ZN(n1127) );
NAND3_X1 U811 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U813 ( .A1(n1142), .A2(n1143), .ZN(n1138) );
XOR2_X1 U814 ( .A(n1144), .B(KEYINPUT46), .Z(n1142) );
NAND2_X1 U815 ( .A1(n1144), .A2(n1145), .ZN(n1137) );
NOR2_X1 U816 ( .A1(G953), .A2(n1146), .ZN(n1136) );
NOR2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(G66) );
NOR3_X1 U818 ( .A1(n1100), .A2(n1149), .A3(n1150), .ZN(n1148) );
NOR3_X1 U819 ( .A1(n1151), .A2(n1102), .A3(n1152), .ZN(n1150) );
INV_X1 U820 ( .A(n1153), .ZN(n1151) );
NOR2_X1 U821 ( .A1(n1154), .A2(n1153), .ZN(n1149) );
NOR2_X1 U822 ( .A1(n1155), .A2(n1102), .ZN(n1154) );
NOR2_X1 U823 ( .A1(n1053), .A2(n1051), .ZN(n1155) );
NOR2_X1 U824 ( .A1(n1147), .A2(n1156), .ZN(G63) );
XNOR2_X1 U825 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR2_X1 U826 ( .A1(n1159), .A2(n1152), .ZN(n1158) );
INV_X1 U827 ( .A(G478), .ZN(n1159) );
NOR2_X1 U828 ( .A1(n1147), .A2(n1160), .ZN(G60) );
XOR2_X1 U829 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U830 ( .A1(n1163), .A2(n1152), .ZN(n1161) );
INV_X1 U831 ( .A(G475), .ZN(n1163) );
XOR2_X1 U832 ( .A(G104), .B(n1164), .Z(G6) );
NOR2_X1 U833 ( .A1(n1147), .A2(n1165), .ZN(G57) );
XOR2_X1 U834 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U835 ( .A(G101), .B(n1168), .Z(n1167) );
NOR3_X1 U836 ( .A1(KEYINPUT35), .A2(n1169), .A3(n1170), .ZN(n1168) );
NOR2_X1 U837 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U838 ( .A(KEYINPUT37), .B(n1173), .Z(n1171) );
NOR2_X1 U839 ( .A1(n1173), .A2(n1174), .ZN(n1169) );
INV_X1 U840 ( .A(n1172), .ZN(n1174) );
XOR2_X1 U841 ( .A(n1175), .B(n1176), .Z(n1172) );
NOR2_X1 U842 ( .A1(KEYINPUT38), .A2(n1177), .ZN(n1176) );
NOR2_X1 U843 ( .A1(n1152), .A2(n1178), .ZN(n1173) );
NOR2_X1 U844 ( .A1(n1147), .A2(n1179), .ZN(G54) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U846 ( .A(n1182), .B(n1183), .ZN(n1181) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U848 ( .A1(n1186), .A2(n1152), .ZN(n1185) );
NOR2_X1 U849 ( .A1(KEYINPUT55), .A2(n1187), .ZN(n1184) );
XOR2_X1 U850 ( .A(n1188), .B(KEYINPUT58), .Z(n1187) );
XOR2_X1 U851 ( .A(n1123), .B(n1189), .Z(n1180) );
XOR2_X1 U852 ( .A(n1190), .B(n1191), .Z(n1123) );
NOR2_X1 U853 ( .A1(n1147), .A2(n1192), .ZN(G51) );
XOR2_X1 U854 ( .A(n1193), .B(n1194), .Z(n1192) );
XNOR2_X1 U855 ( .A(n1195), .B(n1196), .ZN(n1194) );
NOR2_X1 U856 ( .A1(n1197), .A2(n1152), .ZN(n1196) );
NAND2_X1 U857 ( .A1(G902), .A2(n1198), .ZN(n1152) );
NAND2_X1 U858 ( .A1(n1126), .A2(n1146), .ZN(n1198) );
INV_X1 U859 ( .A(n1053), .ZN(n1146) );
NAND2_X1 U860 ( .A1(n1199), .A2(n1200), .ZN(n1053) );
NOR4_X1 U861 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NOR4_X1 U862 ( .A1(n1164), .A2(n1046), .A3(n1205), .A4(n1206), .ZN(n1199) );
NOR2_X1 U863 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR4_X1 U864 ( .A1(n1209), .A2(n1071), .A3(n1210), .A4(n1211), .ZN(n1205) );
XOR2_X1 U865 ( .A(KEYINPUT43), .B(n1092), .Z(n1211) );
INV_X1 U866 ( .A(n1047), .ZN(n1046) );
NAND3_X1 U867 ( .A1(n1077), .A2(n1068), .A3(n1212), .ZN(n1047) );
AND3_X1 U868 ( .A1(n1212), .A2(n1068), .A3(n1213), .ZN(n1164) );
INV_X1 U869 ( .A(n1051), .ZN(n1126) );
NAND2_X1 U870 ( .A1(n1214), .A2(n1215), .ZN(n1051) );
NOR4_X1 U871 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
NOR4_X1 U872 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1214) );
NOR4_X1 U873 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1210), .ZN(n1223) );
NAND2_X1 U874 ( .A1(n1227), .A2(n1228), .ZN(n1193) );
NAND2_X1 U875 ( .A1(n1229), .A2(G125), .ZN(n1228) );
NAND2_X1 U876 ( .A1(n1230), .A2(n1125), .ZN(n1227) );
XOR2_X1 U877 ( .A(n1229), .B(n1231), .Z(n1230) );
XNOR2_X1 U878 ( .A(KEYINPUT60), .B(KEYINPUT34), .ZN(n1231) );
XOR2_X1 U879 ( .A(n1232), .B(n1233), .Z(n1229) );
NOR2_X1 U880 ( .A1(n1109), .A2(G952), .ZN(n1147) );
XOR2_X1 U881 ( .A(G146), .B(n1222), .Z(G48) );
AND3_X1 U882 ( .A1(n1213), .A2(n1234), .A3(n1235), .ZN(n1222) );
XOR2_X1 U883 ( .A(n1236), .B(n1237), .Z(G45) );
NAND2_X1 U884 ( .A1(KEYINPUT53), .A2(G143), .ZN(n1237) );
NAND4_X1 U885 ( .A1(n1238), .A2(n1235), .A3(n1239), .A4(n1240), .ZN(n1236) );
XOR2_X1 U886 ( .A(n1210), .B(KEYINPUT25), .Z(n1238) );
XOR2_X1 U887 ( .A(G140), .B(n1221), .Z(G42) );
AND3_X1 U888 ( .A1(n1083), .A2(n1213), .A3(n1241), .ZN(n1221) );
XOR2_X1 U889 ( .A(G137), .B(n1220), .Z(G39) );
AND3_X1 U890 ( .A1(n1066), .A2(n1234), .A3(n1241), .ZN(n1220) );
XOR2_X1 U891 ( .A(G134), .B(n1219), .Z(G36) );
AND3_X1 U892 ( .A1(n1067), .A2(n1077), .A3(n1241), .ZN(n1219) );
XOR2_X1 U893 ( .A(G131), .B(n1218), .Z(G33) );
AND3_X1 U894 ( .A1(n1067), .A2(n1213), .A3(n1241), .ZN(n1218) );
AND4_X1 U895 ( .A1(n1076), .A2(n1057), .A3(n1242), .A4(n1074), .ZN(n1241) );
INV_X1 U896 ( .A(n1097), .ZN(n1057) );
NAND2_X1 U897 ( .A1(n1089), .A2(n1243), .ZN(n1097) );
INV_X1 U898 ( .A(n1090), .ZN(n1243) );
NAND2_X1 U899 ( .A1(n1244), .A2(n1245), .ZN(G30) );
NAND2_X1 U900 ( .A1(n1217), .A2(n1246), .ZN(n1245) );
XOR2_X1 U901 ( .A(KEYINPUT22), .B(n1247), .Z(n1244) );
NOR2_X1 U902 ( .A1(n1217), .A2(n1246), .ZN(n1247) );
AND3_X1 U903 ( .A1(n1077), .A2(n1234), .A3(n1235), .ZN(n1217) );
INV_X1 U904 ( .A(n1226), .ZN(n1235) );
NAND4_X1 U905 ( .A1(n1076), .A2(n1092), .A3(n1242), .A4(n1074), .ZN(n1226) );
XOR2_X1 U906 ( .A(G101), .B(n1204), .Z(G3) );
AND3_X1 U907 ( .A1(n1066), .A2(n1212), .A3(n1067), .ZN(n1204) );
XOR2_X1 U908 ( .A(n1125), .B(n1248), .Z(G27) );
NAND2_X1 U909 ( .A1(KEYINPUT7), .A2(n1216), .ZN(n1248) );
AND4_X1 U910 ( .A1(n1083), .A2(n1249), .A3(n1092), .A4(n1242), .ZN(n1216) );
NAND2_X1 U911 ( .A1(n1085), .A2(n1250), .ZN(n1242) );
NAND3_X1 U912 ( .A1(G902), .A2(n1251), .A3(n1110), .ZN(n1250) );
NOR2_X1 U913 ( .A1(n1252), .A2(G900), .ZN(n1110) );
INV_X1 U914 ( .A(n1140), .ZN(n1252) );
INV_X1 U915 ( .A(n1071), .ZN(n1249) );
NAND2_X1 U916 ( .A1(n1065), .A2(n1213), .ZN(n1071) );
INV_X1 U917 ( .A(n1253), .ZN(n1213) );
XNOR2_X1 U918 ( .A(G122), .B(n1254), .ZN(G24) );
NAND2_X1 U919 ( .A1(n1255), .A2(n1092), .ZN(n1254) );
XOR2_X1 U920 ( .A(n1208), .B(KEYINPUT5), .Z(n1255) );
NAND3_X1 U921 ( .A1(n1065), .A2(n1068), .A3(n1256), .ZN(n1208) );
NOR3_X1 U922 ( .A1(n1225), .A2(n1209), .A3(n1224), .ZN(n1256) );
NOR2_X1 U923 ( .A1(n1099), .A2(n1257), .ZN(n1068) );
XOR2_X1 U924 ( .A(G119), .B(n1203), .Z(G21) );
AND3_X1 U925 ( .A1(n1066), .A2(n1234), .A3(n1258), .ZN(n1203) );
NAND2_X1 U926 ( .A1(n1259), .A2(n1260), .ZN(n1234) );
NAND3_X1 U927 ( .A1(n1257), .A2(n1099), .A3(n1261), .ZN(n1260) );
INV_X1 U928 ( .A(KEYINPUT45), .ZN(n1261) );
INV_X1 U929 ( .A(n1262), .ZN(n1257) );
NAND2_X1 U930 ( .A1(KEYINPUT45), .A2(n1083), .ZN(n1259) );
XOR2_X1 U931 ( .A(G116), .B(n1202), .Z(G18) );
AND3_X1 U932 ( .A1(n1067), .A2(n1077), .A3(n1258), .ZN(n1202) );
INV_X1 U933 ( .A(n1263), .ZN(n1258) );
NOR2_X1 U934 ( .A1(n1239), .A2(n1224), .ZN(n1077) );
XOR2_X1 U935 ( .A(n1264), .B(n1265), .Z(G15) );
NOR2_X1 U936 ( .A1(KEYINPUT15), .A2(n1266), .ZN(n1265) );
NOR3_X1 U937 ( .A1(n1267), .A2(n1253), .A3(n1263), .ZN(n1264) );
NAND3_X1 U938 ( .A1(n1092), .A2(n1268), .A3(n1065), .ZN(n1263) );
AND2_X1 U939 ( .A1(n1269), .A2(n1270), .ZN(n1065) );
XOR2_X1 U940 ( .A(n1074), .B(KEYINPUT19), .Z(n1269) );
NAND2_X1 U941 ( .A1(n1224), .A2(n1239), .ZN(n1253) );
XOR2_X1 U942 ( .A(KEYINPUT27), .B(n1067), .Z(n1267) );
INV_X1 U943 ( .A(n1210), .ZN(n1067) );
NAND2_X1 U944 ( .A1(n1262), .A2(n1271), .ZN(n1210) );
XOR2_X1 U945 ( .A(KEYINPUT45), .B(n1099), .Z(n1271) );
XNOR2_X1 U946 ( .A(n1201), .B(n1272), .ZN(G12) );
NAND2_X1 U947 ( .A1(KEYINPUT49), .A2(G110), .ZN(n1272) );
AND3_X1 U948 ( .A1(n1066), .A2(n1212), .A3(n1083), .ZN(n1201) );
NOR2_X1 U949 ( .A1(n1099), .A2(n1262), .ZN(n1083) );
XOR2_X1 U950 ( .A(n1100), .B(n1102), .Z(n1262) );
NAND2_X1 U951 ( .A1(G217), .A2(n1273), .ZN(n1102) );
NOR2_X1 U952 ( .A1(n1153), .A2(G902), .ZN(n1100) );
XOR2_X1 U953 ( .A(n1274), .B(n1275), .Z(n1153) );
XOR2_X1 U954 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U955 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR2_X1 U956 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U957 ( .A(n1282), .B(KEYINPUT52), .Z(n1281) );
NAND2_X1 U958 ( .A1(n1283), .A2(n1125), .ZN(n1282) );
NOR2_X1 U959 ( .A1(n1125), .A2(n1283), .ZN(n1280) );
XOR2_X1 U960 ( .A(KEYINPUT11), .B(G140), .Z(n1283) );
INV_X1 U961 ( .A(G125), .ZN(n1125) );
NAND3_X1 U962 ( .A1(n1284), .A2(G221), .A3(KEYINPUT20), .ZN(n1278) );
XNOR2_X1 U963 ( .A(G110), .B(n1285), .ZN(n1274) );
XOR2_X1 U964 ( .A(G137), .B(G119), .Z(n1285) );
XOR2_X1 U965 ( .A(n1286), .B(n1178), .Z(n1099) );
INV_X1 U966 ( .A(G472), .ZN(n1178) );
NAND2_X1 U967 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U968 ( .A(n1289), .B(n1290), .Z(n1287) );
XOR2_X1 U969 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U970 ( .A(KEYINPUT32), .B(G101), .Z(n1292) );
NOR2_X1 U971 ( .A1(n1166), .A2(KEYINPUT13), .ZN(n1291) );
AND2_X1 U972 ( .A1(n1293), .A2(G210), .ZN(n1166) );
XOR2_X1 U973 ( .A(n1175), .B(n1177), .Z(n1289) );
XOR2_X1 U974 ( .A(n1294), .B(n1233), .Z(n1177) );
XOR2_X1 U975 ( .A(n1295), .B(n1296), .Z(n1175) );
XNOR2_X1 U976 ( .A(KEYINPUT59), .B(n1297), .ZN(n1295) );
NOR2_X1 U977 ( .A1(G113), .A2(KEYINPUT8), .ZN(n1297) );
NOR4_X1 U978 ( .A1(n1270), .A2(n1207), .A3(n1209), .A4(n1098), .ZN(n1212) );
INV_X1 U979 ( .A(n1074), .ZN(n1098) );
NAND2_X1 U980 ( .A1(G221), .A2(n1273), .ZN(n1074) );
NAND2_X1 U981 ( .A1(G234), .A2(n1288), .ZN(n1273) );
INV_X1 U982 ( .A(n1268), .ZN(n1209) );
NAND2_X1 U983 ( .A1(n1085), .A2(n1298), .ZN(n1268) );
NAND4_X1 U984 ( .A1(n1299), .A2(n1140), .A3(n1251), .A4(n1141), .ZN(n1298) );
INV_X1 U985 ( .A(G898), .ZN(n1141) );
XOR2_X1 U986 ( .A(n1109), .B(KEYINPUT63), .Z(n1140) );
XOR2_X1 U987 ( .A(n1288), .B(KEYINPUT2), .Z(n1299) );
NAND3_X1 U988 ( .A1(n1300), .A2(n1251), .A3(G952), .ZN(n1085) );
NAND2_X1 U989 ( .A1(G237), .A2(G234), .ZN(n1251) );
INV_X1 U990 ( .A(n1052), .ZN(n1300) );
XOR2_X1 U991 ( .A(n1109), .B(KEYINPUT1), .Z(n1052) );
INV_X1 U992 ( .A(n1092), .ZN(n1207) );
NOR2_X1 U993 ( .A1(n1089), .A2(n1090), .ZN(n1092) );
AND2_X1 U994 ( .A1(G214), .A2(n1301), .ZN(n1090) );
XNOR2_X1 U995 ( .A(n1302), .B(n1197), .ZN(n1089) );
NAND2_X1 U996 ( .A1(G210), .A2(n1301), .ZN(n1197) );
NAND2_X1 U997 ( .A1(n1288), .A2(n1303), .ZN(n1301) );
INV_X1 U998 ( .A(G237), .ZN(n1303) );
NAND2_X1 U999 ( .A1(n1304), .A2(n1288), .ZN(n1302) );
XOR2_X1 U1000 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1001 ( .A(n1307), .B(n1232), .ZN(n1306) );
NAND2_X1 U1002 ( .A1(G224), .A2(n1109), .ZN(n1232) );
NAND2_X1 U1003 ( .A1(n1308), .A2(KEYINPUT4), .ZN(n1307) );
XNOR2_X1 U1004 ( .A(n1233), .B(n1309), .ZN(n1308) );
XOR2_X1 U1005 ( .A(KEYINPUT16), .B(G125), .Z(n1309) );
XNOR2_X1 U1006 ( .A(n1276), .B(n1310), .ZN(n1233) );
NOR2_X1 U1007 ( .A1(G143), .A2(KEYINPUT23), .ZN(n1310) );
XOR2_X1 U1008 ( .A(n1246), .B(n1311), .Z(n1276) );
INV_X1 U1009 ( .A(G128), .ZN(n1246) );
NAND2_X1 U1010 ( .A1(KEYINPUT24), .A2(n1195), .ZN(n1305) );
XNOR2_X1 U1011 ( .A(n1144), .B(n1145), .ZN(n1195) );
INV_X1 U1012 ( .A(n1143), .ZN(n1145) );
XOR2_X1 U1013 ( .A(n1312), .B(n1313), .Z(n1143) );
NOR2_X1 U1014 ( .A1(G101), .A2(KEYINPUT18), .ZN(n1313) );
XOR2_X1 U1015 ( .A(n1314), .B(n1315), .Z(n1312) );
NOR2_X1 U1016 ( .A1(KEYINPUT29), .A2(n1316), .ZN(n1315) );
INV_X1 U1017 ( .A(G104), .ZN(n1316) );
INV_X1 U1018 ( .A(G107), .ZN(n1314) );
XOR2_X1 U1019 ( .A(n1317), .B(n1318), .Z(n1144) );
XOR2_X1 U1020 ( .A(G110), .B(n1319), .Z(n1318) );
XOR2_X1 U1021 ( .A(KEYINPUT44), .B(G113), .Z(n1319) );
XOR2_X1 U1022 ( .A(n1320), .B(n1321), .Z(n1317) );
NOR2_X1 U1023 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NOR3_X1 U1024 ( .A1(KEYINPUT47), .A2(G119), .A3(n1324), .ZN(n1323) );
INV_X1 U1025 ( .A(G116), .ZN(n1324) );
NOR2_X1 U1026 ( .A1(n1296), .A2(n1325), .ZN(n1322) );
INV_X1 U1027 ( .A(KEYINPUT47), .ZN(n1325) );
XOR2_X1 U1028 ( .A(G116), .B(G119), .Z(n1296) );
INV_X1 U1029 ( .A(n1076), .ZN(n1270) );
XOR2_X1 U1030 ( .A(n1186), .B(n1326), .Z(n1076) );
NOR2_X1 U1031 ( .A1(KEYINPUT26), .A2(n1327), .ZN(n1326) );
XOR2_X1 U1032 ( .A(n1103), .B(KEYINPUT3), .Z(n1327) );
NAND2_X1 U1033 ( .A1(n1328), .A2(n1288), .ZN(n1103) );
XOR2_X1 U1034 ( .A(n1329), .B(n1189), .Z(n1328) );
XNOR2_X1 U1035 ( .A(n1330), .B(n1331), .ZN(n1189) );
XOR2_X1 U1036 ( .A(G140), .B(G110), .Z(n1331) );
NAND2_X1 U1037 ( .A1(G227), .A2(n1109), .ZN(n1330) );
NOR2_X1 U1038 ( .A1(n1332), .A2(n1333), .ZN(n1329) );
XOR2_X1 U1039 ( .A(n1334), .B(KEYINPUT51), .Z(n1333) );
NAND2_X1 U1040 ( .A1(n1335), .A2(n1294), .ZN(n1334) );
NOR2_X1 U1041 ( .A1(n1335), .A2(n1294), .ZN(n1332) );
XNOR2_X1 U1042 ( .A(n1182), .B(n1191), .ZN(n1294) );
XNOR2_X1 U1043 ( .A(G137), .B(n1336), .ZN(n1191) );
NAND2_X1 U1044 ( .A1(KEYINPUT10), .A2(G131), .ZN(n1182) );
XOR2_X1 U1045 ( .A(n1190), .B(n1337), .Z(n1335) );
INV_X1 U1046 ( .A(n1188), .ZN(n1337) );
XOR2_X1 U1047 ( .A(n1338), .B(n1339), .Z(n1188) );
XOR2_X1 U1048 ( .A(KEYINPUT61), .B(G107), .Z(n1339) );
XOR2_X1 U1049 ( .A(n1340), .B(G104), .Z(n1338) );
INV_X1 U1050 ( .A(G101), .ZN(n1340) );
XOR2_X1 U1051 ( .A(n1341), .B(G128), .Z(n1190) );
NAND2_X1 U1052 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1053 ( .A1(G143), .A2(n1311), .ZN(n1343) );
XOR2_X1 U1054 ( .A(KEYINPUT31), .B(n1344), .Z(n1342) );
NOR2_X1 U1055 ( .A1(G143), .A2(n1311), .ZN(n1344) );
INV_X1 U1056 ( .A(G469), .ZN(n1186) );
NOR2_X1 U1057 ( .A1(n1240), .A2(n1239), .ZN(n1066) );
INV_X1 U1058 ( .A(n1225), .ZN(n1239) );
XOR2_X1 U1059 ( .A(n1345), .B(G475), .Z(n1225) );
OR2_X1 U1060 ( .A1(n1162), .A2(G902), .ZN(n1345) );
XNOR2_X1 U1061 ( .A(n1346), .B(n1347), .ZN(n1162) );
XOR2_X1 U1062 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1063 ( .A(n1311), .B(n1350), .Z(n1349) );
XOR2_X1 U1064 ( .A(G146), .B(KEYINPUT6), .Z(n1311) );
XOR2_X1 U1065 ( .A(G104), .B(n1351), .Z(n1348) );
NOR2_X1 U1066 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1067 ( .A(n1354), .B(KEYINPUT14), .Z(n1353) );
NAND2_X1 U1068 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NOR2_X1 U1069 ( .A1(n1356), .A2(n1355), .ZN(n1352) );
XOR2_X1 U1070 ( .A(KEYINPUT30), .B(G131), .Z(n1355) );
XNOR2_X1 U1071 ( .A(n1357), .B(G143), .ZN(n1356) );
NAND2_X1 U1072 ( .A1(n1293), .A2(G214), .ZN(n1357) );
NOR2_X1 U1073 ( .A1(G953), .A2(G237), .ZN(n1293) );
XOR2_X1 U1074 ( .A(n1358), .B(n1359), .Z(n1346) );
XOR2_X1 U1075 ( .A(KEYINPUT28), .B(G140), .Z(n1359) );
XOR2_X1 U1076 ( .A(n1266), .B(G125), .Z(n1358) );
INV_X1 U1077 ( .A(G113), .ZN(n1266) );
INV_X1 U1078 ( .A(n1224), .ZN(n1240) );
XOR2_X1 U1079 ( .A(n1360), .B(G478), .Z(n1224) );
NAND2_X1 U1080 ( .A1(n1157), .A2(n1288), .ZN(n1360) );
INV_X1 U1081 ( .A(G902), .ZN(n1288) );
XNOR2_X1 U1082 ( .A(n1361), .B(n1362), .ZN(n1157) );
XOR2_X1 U1083 ( .A(n1363), .B(n1364), .Z(n1362) );
NAND2_X1 U1084 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NAND2_X1 U1085 ( .A1(n1367), .A2(n1336), .ZN(n1366) );
INV_X1 U1086 ( .A(G134), .ZN(n1336) );
XOR2_X1 U1087 ( .A(KEYINPUT41), .B(n1368), .Z(n1367) );
NAND2_X1 U1088 ( .A1(n1369), .A2(G134), .ZN(n1365) );
XOR2_X1 U1089 ( .A(KEYINPUT36), .B(n1368), .Z(n1369) );
XOR2_X1 U1090 ( .A(G128), .B(G143), .Z(n1368) );
NAND2_X1 U1091 ( .A1(KEYINPUT48), .A2(n1370), .ZN(n1363) );
XOR2_X1 U1092 ( .A(G116), .B(n1350), .Z(n1370) );
INV_X1 U1093 ( .A(n1320), .ZN(n1350) );
XNOR2_X1 U1094 ( .A(G122), .B(KEYINPUT17), .ZN(n1320) );
XOR2_X1 U1095 ( .A(n1371), .B(G107), .Z(n1361) );
NAND2_X1 U1096 ( .A1(G217), .A2(n1284), .ZN(n1371) );
AND2_X1 U1097 ( .A1(G234), .A2(n1109), .ZN(n1284) );
INV_X1 U1098 ( .A(G953), .ZN(n1109) );
endmodule


