//Key = 1001101001101101011011100000001110101011010000000000111010100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319;

XNOR2_X1 U732 ( .A(n1004), .B(n1005), .ZN(G9) );
NAND2_X1 U733 ( .A1(KEYINPUT22), .A2(n1006), .ZN(n1004) );
NOR2_X1 U734 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR3_X1 U735 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
XOR2_X1 U736 ( .A(KEYINPUT18), .B(G952), .Z(n1011) );
NAND3_X1 U737 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1009) );
NAND2_X1 U738 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U739 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND4_X1 U740 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NAND3_X1 U741 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
OR2_X1 U743 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND3_X1 U744 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1023) );
NAND4_X1 U745 ( .A1(n1032), .A2(n1026), .A3(n1033), .A4(n1034), .ZN(n1017) );
NAND2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U747 ( .A1(n1020), .A2(n1019), .ZN(n1036) );
NAND4_X1 U748 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1021), .ZN(n1033) );
NAND3_X1 U749 ( .A1(n1040), .A2(n1041), .A3(n1019), .ZN(n1038) );
NAND2_X1 U750 ( .A1(n1020), .A2(n1042), .ZN(n1037) );
INV_X1 U751 ( .A(n1043), .ZN(n1015) );
NOR3_X1 U752 ( .A1(n1044), .A2(G953), .A3(n1045), .ZN(n1007) );
INV_X1 U753 ( .A(n1012), .ZN(n1045) );
NAND4_X1 U754 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1012) );
NOR4_X1 U755 ( .A1(n1031), .A2(n1040), .A3(n1050), .A4(n1051), .ZN(n1049) );
XNOR2_X1 U756 ( .A(G469), .B(n1052), .ZN(n1050) );
NOR2_X1 U757 ( .A1(n1053), .A2(KEYINPUT63), .ZN(n1052) );
NOR2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1048) );
XNOR2_X1 U759 ( .A(G472), .B(n1056), .ZN(n1055) );
XNOR2_X1 U760 ( .A(n1057), .B(n1058), .ZN(n1054) );
XNOR2_X1 U761 ( .A(n1059), .B(n1060), .ZN(n1046) );
XNOR2_X1 U762 ( .A(n1061), .B(KEYINPUT48), .ZN(n1059) );
XOR2_X1 U763 ( .A(KEYINPUT45), .B(G952), .Z(n1044) );
XOR2_X1 U764 ( .A(n1062), .B(n1063), .Z(G72) );
XOR2_X1 U765 ( .A(n1064), .B(n1065), .Z(n1063) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1013), .ZN(n1065) );
AND2_X1 U767 ( .A1(G227), .A2(G900), .ZN(n1066) );
NAND2_X1 U768 ( .A1(n1067), .A2(n1068), .ZN(n1064) );
NAND2_X1 U769 ( .A1(G953), .A2(n1069), .ZN(n1068) );
XOR2_X1 U770 ( .A(n1070), .B(n1071), .Z(n1067) );
XOR2_X1 U771 ( .A(n1072), .B(n1073), .Z(n1071) );
XNOR2_X1 U772 ( .A(n1074), .B(n1075), .ZN(n1073) );
NOR2_X1 U773 ( .A1(G134), .A2(KEYINPUT44), .ZN(n1075) );
XOR2_X1 U774 ( .A(n1076), .B(n1077), .Z(n1070) );
XOR2_X1 U775 ( .A(KEYINPUT12), .B(G140), .Z(n1077) );
NOR2_X1 U776 ( .A1(G125), .A2(KEYINPUT14), .ZN(n1076) );
NAND2_X1 U777 ( .A1(n1013), .A2(n1078), .ZN(n1062) );
XOR2_X1 U778 ( .A(n1079), .B(n1080), .Z(G69) );
NOR2_X1 U779 ( .A1(n1081), .A2(n1013), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U781 ( .A1(n1084), .A2(KEYINPUT51), .A3(n1085), .ZN(n1079) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U783 ( .A(KEYINPUT57), .B(n1088), .ZN(n1087) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NOR2_X1 U785 ( .A1(G898), .A2(n1013), .ZN(n1089) );
NOR2_X1 U786 ( .A1(n1090), .A2(n1088), .ZN(n1084) );
NAND2_X1 U787 ( .A1(n1013), .A2(n1091), .ZN(n1088) );
XOR2_X1 U788 ( .A(n1092), .B(n1093), .Z(n1090) );
NOR2_X1 U789 ( .A1(n1094), .A2(n1095), .ZN(G66) );
XOR2_X1 U790 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U791 ( .A(KEYINPUT35), .B(n1098), .Z(n1097) );
NOR2_X1 U792 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR2_X1 U793 ( .A1(n1094), .A2(n1101), .ZN(G63) );
XNOR2_X1 U794 ( .A(n1102), .B(n1103), .ZN(n1101) );
AND2_X1 U795 ( .A1(G478), .A2(n1104), .ZN(n1102) );
NOR2_X1 U796 ( .A1(n1094), .A2(n1105), .ZN(G60) );
XNOR2_X1 U797 ( .A(n1106), .B(n1107), .ZN(n1105) );
AND2_X1 U798 ( .A1(G475), .A2(n1104), .ZN(n1107) );
XNOR2_X1 U799 ( .A(G104), .B(n1108), .ZN(G6) );
NOR3_X1 U800 ( .A1(n1109), .A2(n1094), .A3(n1110), .ZN(G57) );
NOR3_X1 U801 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1110) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(n1112) );
NOR2_X1 U803 ( .A1(G101), .A2(n1116), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1117), .A2(n1118), .ZN(n1109) );
XOR2_X1 U805 ( .A(n1114), .B(n1119), .Z(n1118) );
NOR2_X1 U806 ( .A1(n1120), .A2(n1116), .ZN(n1119) );
INV_X1 U807 ( .A(KEYINPUT9), .ZN(n1116) );
XNOR2_X1 U808 ( .A(n1121), .B(n1122), .ZN(n1114) );
NOR2_X1 U809 ( .A1(n1123), .A2(n1100), .ZN(n1122) );
NOR2_X1 U810 ( .A1(n1113), .A2(n1111), .ZN(n1117) );
INV_X1 U811 ( .A(KEYINPUT20), .ZN(n1111) );
NOR2_X1 U812 ( .A1(n1094), .A2(n1124), .ZN(G54) );
XOR2_X1 U813 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U814 ( .A(n1072), .B(n1127), .Z(n1126) );
XOR2_X1 U815 ( .A(n1128), .B(n1129), .Z(n1125) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U817 ( .A1(KEYINPUT46), .A2(n1132), .ZN(n1131) );
NAND2_X1 U818 ( .A1(KEYINPUT4), .A2(n1133), .ZN(n1130) );
XOR2_X1 U819 ( .A(KEYINPUT6), .B(n1134), .Z(n1133) );
NAND3_X1 U820 ( .A1(n1104), .A2(G469), .A3(KEYINPUT41), .ZN(n1128) );
INV_X1 U821 ( .A(n1100), .ZN(n1104) );
NOR2_X1 U822 ( .A1(n1094), .A2(n1135), .ZN(G51) );
XOR2_X1 U823 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U825 ( .A1(n1060), .A2(n1100), .ZN(n1139) );
NAND2_X1 U826 ( .A1(G902), .A2(n1010), .ZN(n1100) );
OR2_X1 U827 ( .A1(n1078), .A2(n1091), .ZN(n1010) );
NAND4_X1 U828 ( .A1(n1140), .A2(n1108), .A3(n1141), .A4(n1142), .ZN(n1091) );
NOR4_X1 U829 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1142) );
INV_X1 U830 ( .A(n1006), .ZN(n1144) );
NAND3_X1 U831 ( .A1(n1029), .A2(n1147), .A3(n1148), .ZN(n1006) );
NOR3_X1 U832 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1141) );
NOR3_X1 U833 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
INV_X1 U834 ( .A(KEYINPUT47), .ZN(n1152) );
NOR2_X1 U835 ( .A1(KEYINPUT47), .A2(n1155), .ZN(n1150) );
NOR2_X1 U836 ( .A1(n1156), .A2(n1157), .ZN(n1149) );
NAND3_X1 U837 ( .A1(n1148), .A2(n1147), .A3(n1028), .ZN(n1108) );
NAND2_X1 U838 ( .A1(n1026), .A2(n1158), .ZN(n1140) );
NAND2_X1 U839 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NAND4_X1 U840 ( .A1(n1154), .A2(n1157), .A3(n1019), .A4(n1161), .ZN(n1160) );
NOR2_X1 U841 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
INV_X1 U842 ( .A(KEYINPUT61), .ZN(n1157) );
NAND2_X1 U843 ( .A1(n1164), .A2(n1028), .ZN(n1159) );
NAND2_X1 U844 ( .A1(n1165), .A2(n1166), .ZN(n1078) );
NOR4_X1 U845 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
INV_X1 U846 ( .A(n1171), .ZN(n1169) );
NOR4_X1 U847 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1165) );
NOR3_X1 U848 ( .A1(n1163), .A2(n1154), .A3(n1176), .ZN(n1175) );
INV_X1 U849 ( .A(n1177), .ZN(n1174) );
INV_X1 U850 ( .A(n1178), .ZN(n1173) );
NOR2_X1 U851 ( .A1(n1179), .A2(n1180), .ZN(n1138) );
XOR2_X1 U852 ( .A(n1181), .B(KEYINPUT13), .Z(n1180) );
NAND2_X1 U853 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U854 ( .A1(n1183), .A2(n1182), .ZN(n1179) );
NOR2_X1 U855 ( .A1(n1013), .A2(G952), .ZN(n1094) );
XNOR2_X1 U856 ( .A(n1172), .B(n1184), .ZN(G48) );
NAND2_X1 U857 ( .A1(KEYINPUT30), .A2(G146), .ZN(n1184) );
AND3_X1 U858 ( .A1(n1028), .A2(n1185), .A3(n1186), .ZN(n1172) );
XOR2_X1 U859 ( .A(n1187), .B(n1188), .Z(G45) );
NAND2_X1 U860 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1188) );
NAND3_X1 U861 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1187) );
XNOR2_X1 U862 ( .A(KEYINPUT33), .B(n1154), .ZN(n1190) );
XOR2_X1 U863 ( .A(G140), .B(n1170), .Z(G42) );
AND3_X1 U864 ( .A1(n1192), .A2(n1148), .A3(n1020), .ZN(n1170) );
XNOR2_X1 U865 ( .A(G137), .B(n1171), .ZN(G39) );
NAND3_X1 U866 ( .A1(n1186), .A2(n1020), .A3(n1032), .ZN(n1171) );
XOR2_X1 U867 ( .A(G134), .B(n1168), .Z(G36) );
AND3_X1 U868 ( .A1(n1189), .A2(n1029), .A3(n1020), .ZN(n1168) );
NAND2_X1 U869 ( .A1(n1193), .A2(n1194), .ZN(G33) );
OR2_X1 U870 ( .A1(n1177), .A2(G131), .ZN(n1194) );
XOR2_X1 U871 ( .A(n1195), .B(KEYINPUT40), .Z(n1193) );
NAND2_X1 U872 ( .A1(G131), .A2(n1177), .ZN(n1195) );
NAND3_X1 U873 ( .A1(n1189), .A2(n1028), .A3(n1020), .ZN(n1177) );
NOR2_X1 U874 ( .A1(n1196), .A2(n1040), .ZN(n1020) );
INV_X1 U875 ( .A(n1176), .ZN(n1189) );
NAND4_X1 U876 ( .A1(n1035), .A2(n1148), .A3(n1019), .A4(n1197), .ZN(n1176) );
NAND2_X1 U877 ( .A1(n1198), .A2(n1199), .ZN(G30) );
OR2_X1 U878 ( .A1(n1178), .A2(G128), .ZN(n1199) );
XOR2_X1 U879 ( .A(n1200), .B(KEYINPUT16), .Z(n1198) );
NAND2_X1 U880 ( .A1(G128), .A2(n1178), .ZN(n1200) );
NAND3_X1 U881 ( .A1(n1029), .A2(n1185), .A3(n1186), .ZN(n1178) );
AND4_X1 U882 ( .A1(n1035), .A2(n1148), .A3(n1042), .A4(n1197), .ZN(n1186) );
NAND2_X1 U883 ( .A1(n1201), .A2(n1202), .ZN(G3) );
NAND2_X1 U884 ( .A1(G101), .A2(n1203), .ZN(n1202) );
NAND2_X1 U885 ( .A1(n1143), .A2(n1204), .ZN(n1203) );
NAND2_X1 U886 ( .A1(KEYINPUT5), .A2(KEYINPUT31), .ZN(n1204) );
NAND3_X1 U887 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1201) );
INV_X1 U888 ( .A(KEYINPUT5), .ZN(n1207) );
NAND2_X1 U889 ( .A1(n1143), .A2(n1208), .ZN(n1206) );
INV_X1 U890 ( .A(KEYINPUT31), .ZN(n1208) );
NAND2_X1 U891 ( .A1(KEYINPUT31), .A2(n1209), .ZN(n1205) );
NAND2_X1 U892 ( .A1(n1143), .A2(n1120), .ZN(n1209) );
NOR2_X1 U893 ( .A1(n1210), .A2(n1024), .ZN(n1143) );
INV_X1 U894 ( .A(n1164), .ZN(n1210) );
XNOR2_X1 U895 ( .A(n1183), .B(n1167), .ZN(G27) );
AND3_X1 U896 ( .A1(n1026), .A2(n1185), .A3(n1192), .ZN(n1167) );
AND4_X1 U897 ( .A1(n1028), .A2(n1042), .A3(n1021), .A4(n1197), .ZN(n1192) );
NAND2_X1 U898 ( .A1(n1043), .A2(n1211), .ZN(n1197) );
NAND2_X1 U899 ( .A1(n1212), .A2(n1069), .ZN(n1211) );
INV_X1 U900 ( .A(G900), .ZN(n1069) );
XNOR2_X1 U901 ( .A(G122), .B(n1156), .ZN(G24) );
NAND3_X1 U902 ( .A1(n1026), .A2(n1147), .A3(n1191), .ZN(n1156) );
INV_X1 U903 ( .A(n1163), .ZN(n1191) );
NAND2_X1 U904 ( .A1(n1213), .A2(n1051), .ZN(n1163) );
NOR2_X1 U905 ( .A1(n1162), .A2(n1039), .ZN(n1147) );
XOR2_X1 U906 ( .A(G119), .B(n1146), .Z(G21) );
AND4_X1 U907 ( .A1(n1214), .A2(n1032), .A3(n1185), .A4(n1042), .ZN(n1146) );
XOR2_X1 U908 ( .A(G116), .B(n1145), .Z(G18) );
AND3_X1 U909 ( .A1(n1026), .A2(n1029), .A3(n1164), .ZN(n1145) );
NOR3_X1 U910 ( .A1(n1039), .A2(n1215), .A3(n1021), .ZN(n1164) );
INV_X1 U911 ( .A(n1216), .ZN(n1215) );
NAND2_X1 U912 ( .A1(n1185), .A2(n1019), .ZN(n1039) );
NOR2_X1 U913 ( .A1(n1051), .A2(n1047), .ZN(n1029) );
NAND2_X1 U914 ( .A1(n1217), .A2(n1218), .ZN(G15) );
NAND2_X1 U915 ( .A1(G113), .A2(n1219), .ZN(n1218) );
XOR2_X1 U916 ( .A(KEYINPUT39), .B(n1220), .Z(n1217) );
NOR2_X1 U917 ( .A1(G113), .A2(n1219), .ZN(n1220) );
NAND4_X1 U918 ( .A1(n1214), .A2(n1028), .A3(n1019), .A4(n1221), .ZN(n1219) );
XNOR2_X1 U919 ( .A(KEYINPUT50), .B(n1154), .ZN(n1221) );
INV_X1 U920 ( .A(n1185), .ZN(n1154) );
AND2_X1 U921 ( .A1(n1222), .A2(n1051), .ZN(n1028) );
XOR2_X1 U922 ( .A(KEYINPUT28), .B(n1223), .Z(n1222) );
AND3_X1 U923 ( .A1(n1026), .A2(n1216), .A3(n1035), .ZN(n1214) );
INV_X1 U924 ( .A(n1021), .ZN(n1035) );
AND2_X1 U925 ( .A1(n1030), .A2(n1224), .ZN(n1026) );
XOR2_X1 U926 ( .A(KEYINPUT58), .B(n1031), .Z(n1224) );
XNOR2_X1 U927 ( .A(n1155), .B(n1225), .ZN(G12) );
NOR2_X1 U928 ( .A1(KEYINPUT11), .A2(n1226), .ZN(n1225) );
NAND2_X1 U929 ( .A1(n1153), .A2(n1185), .ZN(n1155) );
NOR2_X1 U930 ( .A1(n1041), .A2(n1040), .ZN(n1185) );
AND2_X1 U931 ( .A1(G214), .A2(n1227), .ZN(n1040) );
INV_X1 U932 ( .A(n1196), .ZN(n1041) );
NAND3_X1 U933 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1196) );
NAND2_X1 U934 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
OR3_X1 U935 ( .A1(n1232), .A2(n1231), .A3(n1233), .ZN(n1229) );
INV_X1 U936 ( .A(n1060), .ZN(n1231) );
NOR2_X1 U937 ( .A1(n1061), .A2(KEYINPUT60), .ZN(n1232) );
NAND2_X1 U938 ( .A1(n1234), .A2(n1233), .ZN(n1228) );
INV_X1 U939 ( .A(KEYINPUT62), .ZN(n1233) );
NAND2_X1 U940 ( .A1(n1061), .A2(n1060), .ZN(n1234) );
NAND2_X1 U941 ( .A1(G210), .A2(n1227), .ZN(n1060) );
NAND2_X1 U942 ( .A1(n1235), .A2(n1236), .ZN(n1227) );
XOR2_X1 U943 ( .A(KEYINPUT52), .B(G237), .Z(n1235) );
AND2_X1 U944 ( .A1(n1237), .A2(n1236), .ZN(n1061) );
XOR2_X1 U945 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U946 ( .A(n1182), .B(n1136), .Z(n1239) );
XNOR2_X1 U947 ( .A(n1092), .B(n1240), .ZN(n1136) );
XOR2_X1 U948 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U949 ( .A1(KEYINPUT19), .A2(n1093), .ZN(n1242) );
NOR2_X1 U950 ( .A1(G953), .A2(n1082), .ZN(n1241) );
INV_X1 U951 ( .A(G224), .ZN(n1082) );
XOR2_X1 U952 ( .A(n1243), .B(n1244), .Z(n1092) );
XNOR2_X1 U953 ( .A(n1226), .B(n1245), .ZN(n1244) );
XOR2_X1 U954 ( .A(KEYINPUT38), .B(G122), .Z(n1245) );
XNOR2_X1 U955 ( .A(G107), .B(n1246), .ZN(n1243) );
XNOR2_X1 U956 ( .A(G125), .B(KEYINPUT36), .ZN(n1238) );
NOR3_X1 U957 ( .A1(n1162), .A2(n1019), .A3(n1024), .ZN(n1153) );
NAND2_X1 U958 ( .A1(n1032), .A2(n1148), .ZN(n1024) );
NOR2_X1 U959 ( .A1(n1030), .A2(n1031), .ZN(n1148) );
AND2_X1 U960 ( .A1(n1247), .A2(G221), .ZN(n1031) );
XOR2_X1 U961 ( .A(n1248), .B(KEYINPUT49), .Z(n1247) );
XNOR2_X1 U962 ( .A(n1053), .B(G469), .ZN(n1030) );
AND2_X1 U963 ( .A1(n1249), .A2(n1236), .ZN(n1053) );
XOR2_X1 U964 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U965 ( .A(n1127), .B(n1132), .Z(n1251) );
XNOR2_X1 U966 ( .A(n1252), .B(n1253), .ZN(n1132) );
XNOR2_X1 U967 ( .A(G140), .B(n1226), .ZN(n1253) );
NAND2_X1 U968 ( .A1(G227), .A2(n1013), .ZN(n1252) );
NAND2_X1 U969 ( .A1(n1254), .A2(n1255), .ZN(n1127) );
NAND2_X1 U970 ( .A1(n1256), .A2(n1005), .ZN(n1255) );
INV_X1 U971 ( .A(G107), .ZN(n1005) );
XOR2_X1 U972 ( .A(KEYINPUT53), .B(n1246), .Z(n1256) );
NAND2_X1 U973 ( .A1(n1246), .A2(G107), .ZN(n1254) );
XOR2_X1 U974 ( .A(G104), .B(G101), .Z(n1246) );
XNOR2_X1 U975 ( .A(n1257), .B(n1258), .ZN(n1250) );
NOR2_X1 U976 ( .A1(KEYINPUT29), .A2(n1134), .ZN(n1258) );
NOR2_X1 U977 ( .A1(KEYINPUT1), .A2(n1072), .ZN(n1257) );
XOR2_X1 U978 ( .A(n1259), .B(KEYINPUT26), .Z(n1072) );
AND2_X1 U979 ( .A1(n1260), .A2(n1223), .ZN(n1032) );
XNOR2_X1 U980 ( .A(n1047), .B(KEYINPUT15), .ZN(n1223) );
INV_X1 U981 ( .A(n1213), .ZN(n1047) );
XNOR2_X1 U982 ( .A(n1261), .B(G478), .ZN(n1213) );
NAND2_X1 U983 ( .A1(n1262), .A2(n1103), .ZN(n1261) );
XOR2_X1 U984 ( .A(n1263), .B(n1264), .Z(n1103) );
XOR2_X1 U985 ( .A(n1265), .B(n1266), .Z(n1264) );
NAND2_X1 U986 ( .A1(G217), .A2(n1267), .ZN(n1266) );
NAND2_X1 U987 ( .A1(n1268), .A2(KEYINPUT17), .ZN(n1265) );
XNOR2_X1 U988 ( .A(G134), .B(n1269), .ZN(n1268) );
XNOR2_X1 U989 ( .A(G107), .B(n1270), .ZN(n1263) );
XOR2_X1 U990 ( .A(G122), .B(G116), .Z(n1270) );
XNOR2_X1 U991 ( .A(G902), .B(KEYINPUT27), .ZN(n1262) );
XOR2_X1 U992 ( .A(KEYINPUT32), .B(n1051), .Z(n1260) );
XNOR2_X1 U993 ( .A(n1271), .B(G475), .ZN(n1051) );
NAND2_X1 U994 ( .A1(n1106), .A2(n1236), .ZN(n1271) );
XNOR2_X1 U995 ( .A(n1272), .B(n1273), .ZN(n1106) );
XOR2_X1 U996 ( .A(n1274), .B(n1275), .Z(n1273) );
NOR2_X1 U997 ( .A1(KEYINPUT23), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U998 ( .A(G146), .B(n1277), .ZN(n1276) );
NOR2_X1 U999 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
AND2_X1 U1000 ( .A1(KEYINPUT7), .A2(n1280), .ZN(n1279) );
NOR2_X1 U1001 ( .A1(KEYINPUT24), .A2(n1280), .ZN(n1278) );
NOR2_X1 U1002 ( .A1(n1281), .A2(n1282), .ZN(n1274) );
XOR2_X1 U1003 ( .A(n1283), .B(KEYINPUT34), .Z(n1282) );
NAND2_X1 U1004 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U1005 ( .A(KEYINPUT59), .B(G131), .Z(n1285) );
NOR2_X1 U1006 ( .A1(G131), .A2(n1284), .ZN(n1281) );
XOR2_X1 U1007 ( .A(n1286), .B(G143), .Z(n1284) );
NAND2_X1 U1008 ( .A1(G214), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U1009 ( .A(G104), .B(n1288), .ZN(n1272) );
XOR2_X1 U1010 ( .A(G122), .B(G113), .Z(n1288) );
INV_X1 U1011 ( .A(n1042), .ZN(n1019) );
XOR2_X1 U1012 ( .A(n1289), .B(n1058), .Z(n1042) );
OR2_X1 U1013 ( .A1(n1290), .A2(n1096), .ZN(n1058) );
XNOR2_X1 U1014 ( .A(n1291), .B(n1292), .ZN(n1096) );
XOR2_X1 U1015 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U1016 ( .A(G128), .B(G119), .Z(n1294) );
XNOR2_X1 U1017 ( .A(KEYINPUT42), .B(n1295), .ZN(n1293) );
INV_X1 U1018 ( .A(G137), .ZN(n1295) );
XOR2_X1 U1019 ( .A(n1296), .B(n1297), .Z(n1291) );
XOR2_X1 U1020 ( .A(n1298), .B(n1299), .Z(n1297) );
NAND2_X1 U1021 ( .A1(KEYINPUT10), .A2(n1226), .ZN(n1299) );
INV_X1 U1022 ( .A(G110), .ZN(n1226) );
NAND3_X1 U1023 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1298) );
NAND2_X1 U1024 ( .A1(KEYINPUT8), .A2(G146), .ZN(n1302) );
OR3_X1 U1025 ( .A1(G146), .A2(KEYINPUT8), .A3(n1303), .ZN(n1301) );
NAND2_X1 U1026 ( .A1(n1303), .A2(n1304), .ZN(n1300) );
NAND2_X1 U1027 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
INV_X1 U1028 ( .A(KEYINPUT8), .ZN(n1306) );
XNOR2_X1 U1029 ( .A(G146), .B(KEYINPUT25), .ZN(n1305) );
INV_X1 U1030 ( .A(n1280), .ZN(n1303) );
XOR2_X1 U1031 ( .A(G140), .B(n1183), .Z(n1280) );
INV_X1 U1032 ( .A(G125), .ZN(n1183) );
NAND2_X1 U1033 ( .A1(n1267), .A2(G221), .ZN(n1296) );
AND2_X1 U1034 ( .A1(G234), .A2(n1013), .ZN(n1267) );
XNOR2_X1 U1035 ( .A(n1236), .B(KEYINPUT37), .ZN(n1290) );
NAND2_X1 U1036 ( .A1(KEYINPUT54), .A2(n1057), .ZN(n1289) );
INV_X1 U1037 ( .A(n1099), .ZN(n1057) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1248), .ZN(n1099) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1236), .ZN(n1248) );
NAND2_X1 U1040 ( .A1(n1021), .A2(n1216), .ZN(n1162) );
NAND2_X1 U1041 ( .A1(n1043), .A2(n1307), .ZN(n1216) );
NAND2_X1 U1042 ( .A1(n1212), .A2(n1083), .ZN(n1307) );
INV_X1 U1043 ( .A(G898), .ZN(n1083) );
AND3_X1 U1044 ( .A1(n1308), .A2(n1309), .A3(G953), .ZN(n1212) );
XNOR2_X1 U1045 ( .A(KEYINPUT43), .B(n1236), .ZN(n1308) );
NAND3_X1 U1046 ( .A1(n1309), .A2(n1013), .A3(G952), .ZN(n1043) );
INV_X1 U1047 ( .A(G953), .ZN(n1013) );
NAND2_X1 U1048 ( .A1(G237), .A2(G234), .ZN(n1309) );
XOR2_X1 U1049 ( .A(n1310), .B(n1056), .Z(n1021) );
NAND2_X1 U1050 ( .A1(n1311), .A2(n1236), .ZN(n1056) );
INV_X1 U1051 ( .A(G902), .ZN(n1236) );
XNOR2_X1 U1052 ( .A(n1312), .B(n1313), .ZN(n1311) );
INV_X1 U1053 ( .A(n1121), .ZN(n1313) );
XOR2_X1 U1054 ( .A(n1134), .B(n1314), .Z(n1121) );
XOR2_X1 U1055 ( .A(n1182), .B(n1093), .Z(n1314) );
XOR2_X1 U1056 ( .A(G113), .B(n1315), .Z(n1093) );
XOR2_X1 U1057 ( .A(G119), .B(G116), .Z(n1315) );
XNOR2_X1 U1058 ( .A(n1259), .B(KEYINPUT55), .ZN(n1182) );
XNOR2_X1 U1059 ( .A(G146), .B(n1269), .ZN(n1259) );
XOR2_X1 U1060 ( .A(G143), .B(G128), .Z(n1269) );
XNOR2_X1 U1061 ( .A(n1316), .B(n1074), .ZN(n1134) );
XOR2_X1 U1062 ( .A(G137), .B(G131), .Z(n1074) );
XNOR2_X1 U1063 ( .A(G134), .B(KEYINPUT0), .ZN(n1316) );
NAND3_X1 U1064 ( .A1(KEYINPUT21), .A2(n1317), .A3(n1318), .ZN(n1312) );
XOR2_X1 U1065 ( .A(n1319), .B(KEYINPUT2), .Z(n1318) );
OR2_X1 U1066 ( .A1(n1113), .A2(n1120), .ZN(n1319) );
NAND2_X1 U1067 ( .A1(n1113), .A2(n1120), .ZN(n1317) );
INV_X1 U1068 ( .A(G101), .ZN(n1120) );
NAND2_X1 U1069 ( .A1(G210), .A2(n1287), .ZN(n1113) );
NOR2_X1 U1070 ( .A1(G953), .A2(G237), .ZN(n1287) );
NAND2_X1 U1071 ( .A1(KEYINPUT3), .A2(n1123), .ZN(n1310) );
INV_X1 U1072 ( .A(G472), .ZN(n1123) );
endmodule


