//Key = 1000100100111000010111001011001100001000010010101110111010100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253;

XNOR2_X1 U694 ( .A(G107), .B(n954), .ZN(G9) );
NOR2_X1 U695 ( .A1(n955), .A2(n956), .ZN(G75) );
NOR4_X1 U696 ( .A1(G953), .A2(n957), .A3(n958), .A4(n959), .ZN(n956) );
NOR2_X1 U697 ( .A1(n960), .A2(n961), .ZN(n958) );
NOR2_X1 U698 ( .A1(n962), .A2(n963), .ZN(n960) );
NOR3_X1 U699 ( .A1(n964), .A2(n965), .A3(n966), .ZN(n963) );
NOR2_X1 U700 ( .A1(n967), .A2(n968), .ZN(n965) );
NOR2_X1 U701 ( .A1(n969), .A2(n970), .ZN(n968) );
NOR2_X1 U702 ( .A1(n971), .A2(n972), .ZN(n969) );
NOR2_X1 U703 ( .A1(n973), .A2(n974), .ZN(n972) );
XNOR2_X1 U704 ( .A(n975), .B(KEYINPUT60), .ZN(n973) );
NOR2_X1 U705 ( .A1(n976), .A2(n977), .ZN(n971) );
NOR2_X1 U706 ( .A1(n978), .A2(n979), .ZN(n976) );
NOR3_X1 U707 ( .A1(n977), .A2(n980), .A3(n981), .ZN(n967) );
NOR2_X1 U708 ( .A1(n982), .A2(n983), .ZN(n980) );
NOR3_X1 U709 ( .A1(n981), .A2(n984), .A3(n970), .ZN(n962) );
INV_X1 U710 ( .A(n985), .ZN(n970) );
NOR2_X1 U711 ( .A1(n986), .A2(n987), .ZN(n984) );
AND2_X1 U712 ( .A1(n988), .A2(n989), .ZN(n987) );
NOR3_X1 U713 ( .A1(n977), .A2(n990), .A3(n966), .ZN(n986) );
NOR2_X1 U714 ( .A1(n991), .A2(n992), .ZN(n990) );
AND2_X1 U715 ( .A1(n993), .A2(n994), .ZN(n991) );
INV_X1 U716 ( .A(n975), .ZN(n981) );
NOR3_X1 U717 ( .A1(n957), .A2(G953), .A3(G952), .ZN(n955) );
AND3_X1 U718 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n957) );
NOR3_X1 U719 ( .A1(n966), .A2(n998), .A3(n994), .ZN(n997) );
XOR2_X1 U720 ( .A(n999), .B(KEYINPUT53), .Z(n996) );
NAND4_X1 U721 ( .A1(n1000), .A2(n975), .A3(n1001), .A4(n1002), .ZN(n999) );
NAND2_X1 U722 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
XOR2_X1 U723 ( .A(KEYINPUT31), .B(n1005), .Z(n1001) );
NOR2_X1 U724 ( .A1(n1003), .A2(n1004), .ZN(n1005) );
XNOR2_X1 U725 ( .A(n1006), .B(n1007), .ZN(n995) );
NAND2_X1 U726 ( .A1(n1008), .A2(KEYINPUT7), .ZN(n1006) );
XNOR2_X1 U727 ( .A(G469), .B(KEYINPUT27), .ZN(n1008) );
XOR2_X1 U728 ( .A(n1009), .B(n1010), .Z(G72) );
XOR2_X1 U729 ( .A(n1011), .B(n1012), .Z(n1010) );
NOR3_X1 U730 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR2_X1 U731 ( .A1(G900), .A2(n1016), .ZN(n1015) );
NOR2_X1 U732 ( .A1(n1017), .A2(n1018), .ZN(n1014) );
XOR2_X1 U733 ( .A(n1019), .B(KEYINPUT21), .Z(n1013) );
NAND2_X1 U734 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
XOR2_X1 U735 ( .A(n1020), .B(n1021), .Z(n1018) );
NAND2_X1 U736 ( .A1(n1022), .A2(G953), .ZN(n1011) );
XOR2_X1 U737 ( .A(n1023), .B(KEYINPUT2), .Z(n1022) );
NAND2_X1 U738 ( .A1(G900), .A2(G227), .ZN(n1023) );
NAND2_X1 U739 ( .A1(n1016), .A2(n1024), .ZN(n1009) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(G69) );
NAND2_X1 U741 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XOR2_X1 U742 ( .A(KEYINPUT44), .B(n1029), .Z(n1025) );
NOR2_X1 U743 ( .A1(n1028), .A2(n1030), .ZN(n1029) );
XOR2_X1 U744 ( .A(KEYINPUT63), .B(n1027), .Z(n1030) );
XNOR2_X1 U745 ( .A(n1031), .B(n1032), .ZN(n1027) );
NOR2_X1 U746 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
XNOR2_X1 U747 ( .A(G953), .B(KEYINPUT24), .ZN(n1034) );
NOR2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
XOR2_X1 U749 ( .A(n1037), .B(KEYINPUT9), .Z(n1035) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1039), .ZN(n1031) );
NAND2_X1 U751 ( .A1(G953), .A2(n1040), .ZN(n1039) );
XOR2_X1 U752 ( .A(KEYINPUT57), .B(n1041), .Z(n1038) );
NAND2_X1 U753 ( .A1(G953), .A2(n1042), .ZN(n1028) );
NAND2_X1 U754 ( .A1(G898), .A2(G224), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1043), .A2(n1044), .ZN(G66) );
XOR2_X1 U756 ( .A(n1045), .B(n1046), .Z(n1044) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U758 ( .A1(n1043), .A2(n1049), .ZN(G63) );
XOR2_X1 U759 ( .A(n1050), .B(n1051), .Z(n1049) );
XNOR2_X1 U760 ( .A(KEYINPUT0), .B(n1052), .ZN(n1051) );
NAND2_X1 U761 ( .A1(n1047), .A2(G478), .ZN(n1050) );
NOR2_X1 U762 ( .A1(n1043), .A2(n1053), .ZN(G60) );
NOR2_X1 U763 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U764 ( .A(n1056), .B(n1057), .Z(n1055) );
NAND2_X1 U765 ( .A1(n1047), .A2(G475), .ZN(n1057) );
NAND2_X1 U766 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U767 ( .A1(n1058), .A2(n1059), .ZN(n1054) );
INV_X1 U768 ( .A(KEYINPUT47), .ZN(n1059) );
XNOR2_X1 U769 ( .A(G104), .B(n1060), .ZN(G6) );
NOR2_X1 U770 ( .A1(n1043), .A2(n1061), .ZN(G57) );
XOR2_X1 U771 ( .A(n1062), .B(n1063), .Z(n1061) );
NAND2_X1 U772 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U773 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XNOR2_X1 U774 ( .A(n1068), .B(KEYINPUT55), .ZN(n1067) );
XNOR2_X1 U775 ( .A(n1069), .B(n1070), .ZN(n1066) );
XOR2_X1 U776 ( .A(n1071), .B(KEYINPUT51), .Z(n1064) );
NAND2_X1 U777 ( .A1(n1068), .A2(n1072), .ZN(n1071) );
XNOR2_X1 U778 ( .A(n1070), .B(n1073), .ZN(n1072) );
NOR2_X1 U779 ( .A1(KEYINPUT25), .A2(n1074), .ZN(n1070) );
AND2_X1 U780 ( .A1(n1047), .A2(G472), .ZN(n1068) );
NOR2_X1 U781 ( .A1(n1043), .A2(n1075), .ZN(G54) );
XOR2_X1 U782 ( .A(n1076), .B(n1077), .Z(n1075) );
NAND2_X1 U783 ( .A1(n1047), .A2(G469), .ZN(n1077) );
NAND2_X1 U784 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NAND2_X1 U785 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U786 ( .A(KEYINPUT49), .B(n1082), .Z(n1078) );
NOR2_X1 U787 ( .A1(n1080), .A2(n1081), .ZN(n1082) );
XOR2_X1 U788 ( .A(n1083), .B(n1084), .Z(n1081) );
OR2_X1 U789 ( .A1(KEYINPUT37), .A2(n1020), .ZN(n1083) );
NOR2_X1 U790 ( .A1(n1043), .A2(n1085), .ZN(G51) );
XOR2_X1 U791 ( .A(n1086), .B(n1087), .Z(n1085) );
XNOR2_X1 U792 ( .A(n1088), .B(n1089), .ZN(n1087) );
NOR2_X1 U793 ( .A1(KEYINPUT38), .A2(n1090), .ZN(n1088) );
XOR2_X1 U794 ( .A(KEYINPUT10), .B(n1091), .Z(n1090) );
XOR2_X1 U795 ( .A(n1092), .B(n1041), .Z(n1086) );
NAND3_X1 U796 ( .A1(n1047), .A2(n1093), .A3(KEYINPUT54), .ZN(n1092) );
AND2_X1 U797 ( .A1(G902), .A2(n959), .ZN(n1047) );
OR3_X1 U798 ( .A1(n1037), .A2(n1024), .A3(n1036), .ZN(n959) );
NAND4_X1 U799 ( .A1(n1094), .A2(n1060), .A3(n1095), .A4(n954), .ZN(n1036) );
NAND3_X1 U800 ( .A1(n985), .A2(n1096), .A3(n978), .ZN(n954) );
NAND3_X1 U801 ( .A1(n985), .A2(n1096), .A3(n979), .ZN(n1060) );
NAND2_X1 U802 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
XNOR2_X1 U803 ( .A(KEYINPUT13), .B(n1099), .ZN(n1097) );
NAND4_X1 U804 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1024) );
AND4_X1 U805 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1103) );
NAND2_X1 U806 ( .A1(n1108), .A2(n1109), .ZN(n1102) );
NAND2_X1 U807 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U808 ( .A1(n979), .A2(n983), .ZN(n1110) );
NAND4_X1 U809 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1037) );
NOR2_X1 U810 ( .A1(n1016), .A2(G952), .ZN(n1043) );
XNOR2_X1 U811 ( .A(n1116), .B(n1100), .ZN(G48) );
NAND2_X1 U812 ( .A1(n1117), .A2(n979), .ZN(n1100) );
XNOR2_X1 U813 ( .A(G146), .B(KEYINPUT30), .ZN(n1116) );
XNOR2_X1 U814 ( .A(G143), .B(n1101), .ZN(G45) );
NAND3_X1 U815 ( .A1(n1118), .A2(n982), .A3(n1119), .ZN(n1101) );
AND3_X1 U816 ( .A1(n992), .A2(n1120), .A3(n1121), .ZN(n1119) );
XOR2_X1 U817 ( .A(G140), .B(n1122), .Z(G42) );
NOR3_X1 U818 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
XNOR2_X1 U819 ( .A(n979), .B(KEYINPUT22), .ZN(n1124) );
XNOR2_X1 U820 ( .A(G137), .B(n1126), .ZN(G39) );
NAND4_X1 U821 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
NOR3_X1 U822 ( .A1(n966), .A2(KEYINPUT32), .A3(n1131), .ZN(n1130) );
XOR2_X1 U823 ( .A(n1132), .B(KEYINPUT29), .Z(n1129) );
XNOR2_X1 U824 ( .A(G134), .B(n1105), .ZN(G36) );
NAND3_X1 U825 ( .A1(n982), .A2(n978), .A3(n1108), .ZN(n1105) );
XNOR2_X1 U826 ( .A(n1133), .B(n1104), .ZN(G33) );
NAND3_X1 U827 ( .A1(n982), .A2(n979), .A3(n1108), .ZN(n1104) );
INV_X1 U828 ( .A(n1123), .ZN(n1108) );
NAND4_X1 U829 ( .A1(n1127), .A2(n1134), .A3(n992), .A4(n1132), .ZN(n1123) );
INV_X1 U830 ( .A(n977), .ZN(n1127) );
XOR2_X1 U831 ( .A(n998), .B(KEYINPUT35), .Z(n977) );
NAND2_X1 U832 ( .A1(KEYINPUT46), .A2(n1135), .ZN(n1133) );
XOR2_X1 U833 ( .A(n1136), .B(G128), .Z(G30) );
NAND2_X1 U834 ( .A1(KEYINPUT17), .A2(n1107), .ZN(n1136) );
NAND2_X1 U835 ( .A1(n1117), .A2(n978), .ZN(n1107) );
AND4_X1 U836 ( .A1(n1118), .A2(n992), .A3(n1137), .A4(n1138), .ZN(n1117) );
XOR2_X1 U837 ( .A(G101), .B(n1139), .Z(G3) );
NOR2_X1 U838 ( .A1(n1140), .A2(n1099), .ZN(n1139) );
NAND4_X1 U839 ( .A1(n982), .A2(n975), .A3(n992), .A4(n1141), .ZN(n1099) );
XNOR2_X1 U840 ( .A(G125), .B(n1106), .ZN(G27) );
NAND4_X1 U841 ( .A1(n1118), .A2(n989), .A3(n979), .A4(n983), .ZN(n1106) );
INV_X1 U842 ( .A(n1142), .ZN(n979) );
AND2_X1 U843 ( .A1(n988), .A2(n1132), .ZN(n1118) );
NAND2_X1 U844 ( .A1(n961), .A2(n1143), .ZN(n1132) );
NAND4_X1 U845 ( .A1(G953), .A2(G902), .A3(n1144), .A4(n1145), .ZN(n1143) );
INV_X1 U846 ( .A(G900), .ZN(n1145) );
XNOR2_X1 U847 ( .A(G122), .B(n1112), .ZN(G24) );
NAND4_X1 U848 ( .A1(n1146), .A2(n985), .A3(n1121), .A4(n1120), .ZN(n1112) );
NOR2_X1 U849 ( .A1(n1138), .A2(n1137), .ZN(n985) );
XNOR2_X1 U850 ( .A(G119), .B(n1113), .ZN(G21) );
NAND2_X1 U851 ( .A1(n1128), .A2(n1146), .ZN(n1113) );
INV_X1 U852 ( .A(n1111), .ZN(n1128) );
NAND3_X1 U853 ( .A1(n1137), .A2(n1138), .A3(n975), .ZN(n1111) );
XOR2_X1 U854 ( .A(n1114), .B(n1147), .Z(G18) );
NAND2_X1 U855 ( .A1(KEYINPUT11), .A2(G116), .ZN(n1147) );
NAND3_X1 U856 ( .A1(n982), .A2(n978), .A3(n1146), .ZN(n1114) );
AND3_X1 U857 ( .A1(n988), .A2(n1141), .A3(n989), .ZN(n1146) );
NOR2_X1 U858 ( .A1(n1120), .A2(n1148), .ZN(n978) );
INV_X1 U859 ( .A(n1121), .ZN(n1148) );
XOR2_X1 U860 ( .A(n1115), .B(n1149), .Z(G15) );
NAND2_X1 U861 ( .A1(KEYINPUT12), .A2(G113), .ZN(n1149) );
NAND3_X1 U862 ( .A1(n989), .A2(n982), .A3(n1150), .ZN(n1115) );
NOR3_X1 U863 ( .A1(n1142), .A2(n1151), .A3(n1140), .ZN(n1150) );
NAND2_X1 U864 ( .A1(n1152), .A2(n1120), .ZN(n1142) );
XNOR2_X1 U865 ( .A(n1121), .B(KEYINPUT14), .ZN(n1152) );
NOR2_X1 U866 ( .A1(n1137), .A2(n1153), .ZN(n982) );
INV_X1 U867 ( .A(n964), .ZN(n989) );
NAND2_X1 U868 ( .A1(n1154), .A2(n1155), .ZN(n964) );
XOR2_X1 U869 ( .A(KEYINPUT34), .B(n993), .Z(n1154) );
XNOR2_X1 U870 ( .A(G110), .B(n1095), .ZN(G12) );
NAND3_X1 U871 ( .A1(n975), .A2(n1096), .A3(n983), .ZN(n1095) );
INV_X1 U872 ( .A(n1125), .ZN(n983) );
NAND2_X1 U873 ( .A1(n1153), .A2(n1137), .ZN(n1125) );
XNOR2_X1 U874 ( .A(n1000), .B(KEYINPUT28), .ZN(n1137) );
XOR2_X1 U875 ( .A(n1156), .B(n1048), .Z(n1000) );
AND2_X1 U876 ( .A1(G217), .A2(n1157), .ZN(n1048) );
NAND2_X1 U877 ( .A1(n1046), .A2(n1158), .ZN(n1156) );
XOR2_X1 U878 ( .A(n1159), .B(n1160), .Z(n1046) );
NOR2_X1 U879 ( .A1(KEYINPUT62), .A2(n1161), .ZN(n1160) );
XOR2_X1 U880 ( .A(n1162), .B(n1163), .Z(n1159) );
AND3_X1 U881 ( .A1(G221), .A2(n1016), .A3(n1164), .ZN(n1163) );
NAND2_X1 U882 ( .A1(n1165), .A2(KEYINPUT48), .ZN(n1162) );
XOR2_X1 U883 ( .A(n1166), .B(n1167), .Z(n1165) );
XNOR2_X1 U884 ( .A(G128), .B(n1168), .ZN(n1167) );
XNOR2_X1 U885 ( .A(KEYINPUT61), .B(KEYINPUT43), .ZN(n1168) );
XNOR2_X1 U886 ( .A(n1169), .B(n1170), .ZN(n1166) );
NOR2_X1 U887 ( .A1(KEYINPUT18), .A2(n1171), .ZN(n1170) );
XNOR2_X1 U888 ( .A(G146), .B(n1017), .ZN(n1171) );
INV_X1 U889 ( .A(n1138), .ZN(n1153) );
XOR2_X1 U890 ( .A(n1172), .B(n1004), .Z(n1138) );
INV_X1 U891 ( .A(G472), .ZN(n1004) );
NAND2_X1 U892 ( .A1(KEYINPUT20), .A2(n1003), .ZN(n1172) );
AND2_X1 U893 ( .A1(n1173), .A2(n1158), .ZN(n1003) );
XNOR2_X1 U894 ( .A(n1063), .B(n1174), .ZN(n1173) );
XOR2_X1 U895 ( .A(n1175), .B(n1074), .Z(n1174) );
AND2_X1 U896 ( .A1(n1176), .A2(n1177), .ZN(n1074) );
NAND2_X1 U897 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U898 ( .A(KEYINPUT19), .B(n1180), .Z(n1176) );
NOR2_X1 U899 ( .A1(n1179), .A2(n1178), .ZN(n1180) );
XOR2_X1 U900 ( .A(G116), .B(n1181), .Z(n1178) );
XOR2_X1 U901 ( .A(KEYINPUT41), .B(G119), .Z(n1181) );
NAND2_X1 U902 ( .A1(KEYINPUT52), .A2(n1073), .ZN(n1175) );
INV_X1 U903 ( .A(n1069), .ZN(n1073) );
XNOR2_X1 U904 ( .A(n1182), .B(n1020), .ZN(n1069) );
XNOR2_X1 U905 ( .A(n1183), .B(G101), .ZN(n1063) );
NAND2_X1 U906 ( .A1(G210), .A2(n1184), .ZN(n1183) );
NOR3_X1 U907 ( .A1(n1140), .A2(n1151), .A3(n1131), .ZN(n1096) );
INV_X1 U908 ( .A(n992), .ZN(n1131) );
NOR2_X1 U909 ( .A1(n993), .A2(n994), .ZN(n992) );
INV_X1 U910 ( .A(n1155), .ZN(n994) );
NAND2_X1 U911 ( .A1(G221), .A2(n1157), .ZN(n1155) );
NAND2_X1 U912 ( .A1(G234), .A2(n1158), .ZN(n1157) );
XNOR2_X1 U913 ( .A(n1007), .B(n1185), .ZN(n993) );
NOR2_X1 U914 ( .A1(G469), .A2(KEYINPUT15), .ZN(n1185) );
NAND2_X1 U915 ( .A1(n1186), .A2(n1187), .ZN(n1007) );
XOR2_X1 U916 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U917 ( .A(n1084), .B(n1020), .Z(n1189) );
XNOR2_X1 U918 ( .A(n1135), .B(n1190), .ZN(n1020) );
XNOR2_X1 U919 ( .A(n1161), .B(G134), .ZN(n1190) );
INV_X1 U920 ( .A(G137), .ZN(n1161) );
XOR2_X1 U921 ( .A(n1191), .B(n1192), .Z(n1084) );
XNOR2_X1 U922 ( .A(n1193), .B(KEYINPUT6), .ZN(n1192) );
NAND2_X1 U923 ( .A1(KEYINPUT36), .A2(G101), .ZN(n1193) );
XOR2_X1 U924 ( .A(n1194), .B(n1021), .Z(n1191) );
XNOR2_X1 U925 ( .A(n1195), .B(n1196), .ZN(n1021) );
XNOR2_X1 U926 ( .A(G128), .B(KEYINPUT50), .ZN(n1195) );
XNOR2_X1 U927 ( .A(n1080), .B(KEYINPUT3), .ZN(n1188) );
AND2_X1 U928 ( .A1(n1197), .A2(n1198), .ZN(n1080) );
NAND3_X1 U929 ( .A1(G227), .A2(n1016), .A3(n1199), .ZN(n1198) );
XNOR2_X1 U930 ( .A(G110), .B(G140), .ZN(n1199) );
NAND2_X1 U931 ( .A1(n1200), .A2(n1201), .ZN(n1197) );
NAND2_X1 U932 ( .A1(G227), .A2(n1016), .ZN(n1201) );
XOR2_X1 U933 ( .A(G140), .B(G110), .Z(n1200) );
XNOR2_X1 U934 ( .A(KEYINPUT4), .B(n1158), .ZN(n1186) );
INV_X1 U935 ( .A(n1141), .ZN(n1151) );
NAND2_X1 U936 ( .A1(n961), .A2(n1202), .ZN(n1141) );
NAND4_X1 U937 ( .A1(G953), .A2(G902), .A3(n1144), .A4(n1040), .ZN(n1202) );
INV_X1 U938 ( .A(G898), .ZN(n1040) );
NAND3_X1 U939 ( .A1(n1144), .A2(n1016), .A3(G952), .ZN(n961) );
NAND2_X1 U940 ( .A1(G237), .A2(G234), .ZN(n1144) );
INV_X1 U941 ( .A(n1098), .ZN(n1140) );
XOR2_X1 U942 ( .A(n988), .B(KEYINPUT5), .Z(n1098) );
NOR2_X1 U943 ( .A1(n1134), .A2(n998), .ZN(n988) );
INV_X1 U944 ( .A(n974), .ZN(n998) );
NAND2_X1 U945 ( .A1(G214), .A2(n1203), .ZN(n974) );
INV_X1 U946 ( .A(n966), .ZN(n1134) );
XNOR2_X1 U947 ( .A(n1204), .B(n1093), .ZN(n966) );
AND2_X1 U948 ( .A1(G210), .A2(n1203), .ZN(n1093) );
NAND2_X1 U949 ( .A1(n1205), .A2(n1158), .ZN(n1203) );
INV_X1 U950 ( .A(G237), .ZN(n1205) );
NAND3_X1 U951 ( .A1(n1206), .A2(n1158), .A3(n1207), .ZN(n1204) );
XOR2_X1 U952 ( .A(n1208), .B(KEYINPUT45), .Z(n1207) );
NAND2_X1 U953 ( .A1(n1209), .A2(n1041), .ZN(n1208) );
OR2_X1 U954 ( .A1(n1041), .A2(n1209), .ZN(n1206) );
XOR2_X1 U955 ( .A(n1091), .B(n1210), .Z(n1209) );
NOR2_X1 U956 ( .A1(KEYINPUT59), .A2(n1089), .ZN(n1210) );
NAND2_X1 U957 ( .A1(G224), .A2(n1016), .ZN(n1089) );
XNOR2_X1 U958 ( .A(n1182), .B(n1211), .ZN(n1091) );
XOR2_X1 U959 ( .A(KEYINPUT23), .B(G125), .Z(n1211) );
XOR2_X1 U960 ( .A(n1212), .B(n1213), .Z(n1182) );
NAND2_X1 U961 ( .A1(KEYINPUT56), .A2(n1214), .ZN(n1212) );
INV_X1 U962 ( .A(G146), .ZN(n1214) );
XNOR2_X1 U963 ( .A(n1215), .B(n1216), .ZN(n1041) );
XOR2_X1 U964 ( .A(G101), .B(n1217), .Z(n1216) );
XNOR2_X1 U965 ( .A(G116), .B(n1179), .ZN(n1217) );
XOR2_X1 U966 ( .A(n1194), .B(n1218), .Z(n1215) );
XOR2_X1 U967 ( .A(n1219), .B(n1169), .Z(n1218) );
XOR2_X1 U968 ( .A(G119), .B(G110), .Z(n1169) );
NOR2_X1 U969 ( .A1(G122), .A2(KEYINPUT1), .ZN(n1219) );
XNOR2_X1 U970 ( .A(G104), .B(G107), .ZN(n1194) );
NOR2_X1 U971 ( .A1(n1121), .A2(n1120), .ZN(n975) );
XNOR2_X1 U972 ( .A(n1220), .B(G475), .ZN(n1120) );
NAND2_X1 U973 ( .A1(n1058), .A2(n1158), .ZN(n1220) );
XNOR2_X1 U974 ( .A(n1221), .B(n1222), .ZN(n1058) );
XOR2_X1 U975 ( .A(n1223), .B(n1224), .Z(n1222) );
XNOR2_X1 U976 ( .A(G122), .B(n1179), .ZN(n1224) );
INV_X1 U977 ( .A(G113), .ZN(n1179) );
XNOR2_X1 U978 ( .A(KEYINPUT8), .B(n1135), .ZN(n1223) );
INV_X1 U979 ( .A(G131), .ZN(n1135) );
XOR2_X1 U980 ( .A(n1225), .B(n1226), .Z(n1221) );
XOR2_X1 U981 ( .A(n1196), .B(n1017), .Z(n1226) );
XOR2_X1 U982 ( .A(G125), .B(G140), .Z(n1017) );
XNOR2_X1 U983 ( .A(n1227), .B(G146), .ZN(n1196) );
INV_X1 U984 ( .A(G143), .ZN(n1227) );
XNOR2_X1 U985 ( .A(n1228), .B(n1229), .ZN(n1225) );
INV_X1 U986 ( .A(G104), .ZN(n1229) );
NAND2_X1 U987 ( .A1(G214), .A2(n1184), .ZN(n1228) );
NOR2_X1 U988 ( .A1(G953), .A2(G237), .ZN(n1184) );
XNOR2_X1 U989 ( .A(n1230), .B(G478), .ZN(n1121) );
NAND2_X1 U990 ( .A1(n1158), .A2(n1052), .ZN(n1230) );
NAND3_X1 U991 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1052) );
NAND2_X1 U992 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND3_X1 U993 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1235) );
NAND2_X1 U994 ( .A1(KEYINPUT33), .A2(n1239), .ZN(n1238) );
NAND2_X1 U995 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
INV_X1 U996 ( .A(KEYINPUT26), .ZN(n1241) );
NAND2_X1 U997 ( .A1(KEYINPUT26), .A2(n1242), .ZN(n1236) );
NAND2_X1 U998 ( .A1(n1240), .A2(n1243), .ZN(n1242) );
NAND2_X1 U999 ( .A1(KEYINPUT16), .A2(n1244), .ZN(n1243) );
NAND4_X1 U1000 ( .A1(n1245), .A2(n1239), .A3(n1240), .A4(n1244), .ZN(n1232) );
INV_X1 U1001 ( .A(KEYINPUT33), .ZN(n1244) );
INV_X1 U1002 ( .A(KEYINPUT16), .ZN(n1239) );
NAND2_X1 U1003 ( .A1(KEYINPUT33), .A2(n1246), .ZN(n1231) );
NAND2_X1 U1004 ( .A1(n1240), .A2(n1247), .ZN(n1246) );
NAND2_X1 U1005 ( .A1(KEYINPUT16), .A2(n1245), .ZN(n1247) );
INV_X1 U1006 ( .A(n1234), .ZN(n1245) );
XNOR2_X1 U1007 ( .A(n1248), .B(n1249), .ZN(n1234) );
XOR2_X1 U1008 ( .A(G107), .B(n1250), .Z(n1249) );
XOR2_X1 U1009 ( .A(G134), .B(G116), .Z(n1250) );
XNOR2_X1 U1010 ( .A(n1251), .B(n1252), .ZN(n1248) );
NOR2_X1 U1011 ( .A1(G122), .A2(KEYINPUT40), .ZN(n1252) );
NOR2_X1 U1012 ( .A1(KEYINPUT42), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U1013 ( .A(n1213), .B(KEYINPUT58), .ZN(n1253) );
XOR2_X1 U1014 ( .A(G143), .B(G128), .Z(n1213) );
AND3_X1 U1015 ( .A1(n1164), .A2(n1016), .A3(G217), .ZN(n1240) );
INV_X1 U1016 ( .A(G953), .ZN(n1016) );
XOR2_X1 U1017 ( .A(G234), .B(KEYINPUT39), .Z(n1164) );
INV_X1 U1018 ( .A(G902), .ZN(n1158) );
endmodule


