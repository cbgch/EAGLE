//Key = 1011001111110001011111000000111011100000011101001011011100111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377;

XNOR2_X1 U739 ( .A(n1034), .B(n1035), .ZN(G9) );
NOR2_X1 U740 ( .A1(n1036), .A2(n1037), .ZN(G75) );
NOR4_X1 U741 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1037) );
INV_X1 U742 ( .A(G952), .ZN(n1041) );
NOR2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U745 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U746 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
AND4_X1 U747 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(KEYINPUT7), .ZN(n1044) );
OR2_X1 U748 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U749 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U750 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U751 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U752 ( .A1(n1061), .A2(n1062), .ZN(n1053) );
NOR2_X1 U753 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U754 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
INV_X1 U755 ( .A(n1067), .ZN(n1039) );
NAND3_X1 U756 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1038) );
NAND3_X1 U757 ( .A1(n1052), .A2(n1071), .A3(n1072), .ZN(n1070) );
INV_X1 U758 ( .A(n1047), .ZN(n1072) );
NAND4_X1 U759 ( .A1(KEYINPUT7), .A2(n1073), .A3(n1074), .A4(n1050), .ZN(n1047) );
NAND2_X1 U760 ( .A1(n1075), .A2(n1076), .ZN(n1071) );
NAND2_X1 U761 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XNOR2_X1 U762 ( .A(n1079), .B(KEYINPUT8), .ZN(n1077) );
NOR3_X1 U763 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1036) );
NOR2_X1 U764 ( .A1(KEYINPUT23), .A2(n1083), .ZN(n1082) );
NOR2_X1 U765 ( .A1(G953), .A2(G952), .ZN(n1083) );
NOR2_X1 U766 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
INV_X1 U767 ( .A(KEYINPUT23), .ZN(n1085) );
INV_X1 U768 ( .A(n1068), .ZN(n1080) );
NAND4_X1 U769 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1068) );
NOR4_X1 U770 ( .A1(n1090), .A2(n1091), .A3(n1079), .A4(n1092), .ZN(n1089) );
NOR2_X1 U771 ( .A1(n1062), .A2(n1093), .ZN(n1088) );
NAND2_X1 U772 ( .A1(n1094), .A2(n1095), .ZN(n1087) );
XNOR2_X1 U773 ( .A(n1096), .B(KEYINPUT28), .ZN(n1094) );
XOR2_X1 U774 ( .A(KEYINPUT1), .B(n1097), .Z(n1086) );
NOR2_X1 U775 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U776 ( .A(KEYINPUT40), .B(n1100), .Z(n1099) );
AND2_X1 U777 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U778 ( .A(n1103), .B(n1104), .Z(G72) );
XOR2_X1 U779 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U780 ( .A1(n1069), .A2(n1107), .ZN(n1106) );
NAND2_X1 U781 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
XOR2_X1 U782 ( .A(n1110), .B(n1111), .Z(n1108) );
XNOR2_X1 U783 ( .A(n1112), .B(n1113), .ZN(n1111) );
XNOR2_X1 U784 ( .A(G134), .B(n1114), .ZN(n1110) );
NAND2_X1 U785 ( .A1(KEYINPUT21), .A2(G137), .ZN(n1114) );
NOR2_X1 U786 ( .A1(n1115), .A2(n1069), .ZN(n1103) );
AND2_X1 U787 ( .A1(G227), .A2(G900), .ZN(n1115) );
XOR2_X1 U788 ( .A(n1116), .B(n1117), .Z(G69) );
XOR2_X1 U789 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U790 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U791 ( .A1(G898), .A2(G224), .ZN(n1121) );
XNOR2_X1 U792 ( .A(KEYINPUT16), .B(n1069), .ZN(n1120) );
NAND2_X1 U793 ( .A1(n1122), .A2(n1123), .ZN(n1118) );
NAND2_X1 U794 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U795 ( .A(n1126), .B(n1127), .Z(n1122) );
XNOR2_X1 U796 ( .A(G122), .B(G110), .ZN(n1127) );
NAND4_X1 U797 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1126) );
NAND3_X1 U798 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
INV_X1 U799 ( .A(KEYINPUT25), .ZN(n1134) );
NAND2_X1 U800 ( .A1(KEYINPUT33), .A2(n1135), .ZN(n1133) );
NAND3_X1 U801 ( .A1(n1136), .A2(n1137), .A3(KEYINPUT25), .ZN(n1130) );
NAND2_X1 U802 ( .A1(n1135), .A2(n1138), .ZN(n1137) );
NAND3_X1 U803 ( .A1(n1139), .A2(n1135), .A3(n1140), .ZN(n1129) );
XNOR2_X1 U804 ( .A(n1138), .B(n1132), .ZN(n1139) );
INV_X1 U805 ( .A(KEYINPUT33), .ZN(n1138) );
OR2_X1 U806 ( .A1(n1135), .A2(n1140), .ZN(n1128) );
INV_X1 U807 ( .A(KEYINPUT5), .ZN(n1140) );
XNOR2_X1 U808 ( .A(G107), .B(n1141), .ZN(n1135) );
NOR2_X1 U809 ( .A1(n1142), .A2(G953), .ZN(n1116) );
NOR2_X1 U810 ( .A1(n1035), .A2(n1143), .ZN(n1142) );
NOR2_X1 U811 ( .A1(n1084), .A2(n1144), .ZN(G66) );
NOR3_X1 U812 ( .A1(n1102), .A2(n1145), .A3(n1146), .ZN(n1144) );
NOR2_X1 U813 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U814 ( .A1(n1067), .A2(n1101), .ZN(n1147) );
AND3_X1 U815 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1145) );
NOR2_X1 U816 ( .A1(n1084), .A2(n1151), .ZN(G63) );
XOR2_X1 U817 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U818 ( .A1(n1150), .A2(G478), .ZN(n1152) );
NOR2_X1 U819 ( .A1(n1084), .A2(n1154), .ZN(G60) );
XOR2_X1 U820 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U821 ( .A1(KEYINPUT49), .A2(n1157), .ZN(n1156) );
NAND2_X1 U822 ( .A1(n1150), .A2(G475), .ZN(n1155) );
XOR2_X1 U823 ( .A(G104), .B(n1158), .Z(G6) );
AND2_X1 U824 ( .A1(n1159), .A2(n1049), .ZN(n1158) );
NOR2_X1 U825 ( .A1(n1084), .A2(n1160), .ZN(G57) );
XNOR2_X1 U826 ( .A(n1161), .B(n1162), .ZN(n1160) );
NAND3_X1 U827 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1161) );
NAND2_X1 U828 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
OR3_X1 U829 ( .A1(n1167), .A2(n1166), .A3(KEYINPUT57), .ZN(n1164) );
NAND2_X1 U830 ( .A1(KEYINPUT3), .A2(n1168), .ZN(n1167) );
INV_X1 U831 ( .A(n1169), .ZN(n1168) );
NAND2_X1 U832 ( .A1(KEYINPUT57), .A2(n1169), .ZN(n1163) );
NAND2_X1 U833 ( .A1(n1150), .A2(G472), .ZN(n1169) );
NOR2_X1 U834 ( .A1(n1084), .A2(n1170), .ZN(G54) );
NOR3_X1 U835 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
NOR2_X1 U836 ( .A1(KEYINPUT58), .A2(n1174), .ZN(n1173) );
AND3_X1 U837 ( .A1(n1174), .A2(n1175), .A3(KEYINPUT58), .ZN(n1172) );
NOR2_X1 U838 ( .A1(n1176), .A2(n1175), .ZN(n1171) );
XNOR2_X1 U839 ( .A(n1177), .B(n1178), .ZN(n1175) );
XNOR2_X1 U840 ( .A(KEYINPUT10), .B(n1179), .ZN(n1178) );
XOR2_X1 U841 ( .A(n1180), .B(n1181), .Z(n1177) );
NAND2_X1 U842 ( .A1(KEYINPUT6), .A2(n1112), .ZN(n1180) );
NOR2_X1 U843 ( .A1(n1182), .A2(n1183), .ZN(n1176) );
INV_X1 U844 ( .A(KEYINPUT58), .ZN(n1183) );
XNOR2_X1 U845 ( .A(n1174), .B(KEYINPUT35), .ZN(n1182) );
AND2_X1 U846 ( .A1(n1150), .A2(G469), .ZN(n1174) );
NOR2_X1 U847 ( .A1(n1084), .A2(n1184), .ZN(G51) );
XOR2_X1 U848 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND2_X1 U849 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NAND2_X1 U850 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U851 ( .A(n1191), .B(KEYINPUT46), .Z(n1189) );
NAND2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(n1187) );
XOR2_X1 U853 ( .A(n1191), .B(KEYINPUT59), .Z(n1193) );
NAND2_X1 U854 ( .A1(n1150), .A2(n1194), .ZN(n1191) );
NOR2_X1 U855 ( .A1(n1195), .A2(n1067), .ZN(n1150) );
NOR3_X1 U856 ( .A1(n1143), .A2(n1196), .A3(n1107), .ZN(n1067) );
NAND2_X1 U857 ( .A1(n1197), .A2(n1198), .ZN(n1107) );
NOR4_X1 U858 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NOR4_X1 U859 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1197) );
INV_X1 U860 ( .A(n1207), .ZN(n1206) );
XNOR2_X1 U861 ( .A(KEYINPUT48), .B(n1035), .ZN(n1196) );
AND2_X1 U862 ( .A1(n1048), .A2(n1159), .ZN(n1035) );
NOR3_X1 U863 ( .A1(n1056), .A2(n1208), .A3(n1209), .ZN(n1159) );
NAND4_X1 U864 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1143) );
NOR4_X1 U865 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
AND2_X1 U866 ( .A1(n1218), .A2(KEYINPUT61), .ZN(n1217) );
NOR4_X1 U867 ( .A1(n1056), .A2(n1209), .A3(n1219), .A4(n1220), .ZN(n1216) );
XNOR2_X1 U868 ( .A(KEYINPUT41), .B(n1208), .ZN(n1220) );
INV_X1 U869 ( .A(n1074), .ZN(n1056) );
NOR2_X1 U870 ( .A1(n1221), .A2(n1222), .ZN(n1215) );
NOR2_X1 U871 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
XOR2_X1 U872 ( .A(KEYINPUT27), .B(n1225), .Z(n1224) );
XNOR2_X1 U873 ( .A(KEYINPUT44), .B(n1226), .ZN(n1223) );
NOR4_X1 U874 ( .A1(n1058), .A2(n1227), .A3(n1066), .A4(n1228), .ZN(n1214) );
OR2_X1 U875 ( .A1(n1075), .A2(KEYINPUT61), .ZN(n1227) );
NOR2_X1 U876 ( .A1(n1069), .A2(G952), .ZN(n1084) );
XNOR2_X1 U877 ( .A(n1229), .B(n1203), .ZN(G48) );
AND2_X1 U878 ( .A1(n1049), .A2(n1230), .ZN(n1203) );
XOR2_X1 U879 ( .A(n1231), .B(n1202), .Z(G45) );
AND3_X1 U880 ( .A1(n1232), .A2(n1064), .A3(n1233), .ZN(n1202) );
NOR3_X1 U881 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NOR2_X1 U882 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
INV_X1 U883 ( .A(KEYINPUT50), .ZN(n1238) );
NOR2_X1 U884 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
NOR2_X1 U885 ( .A1(KEYINPUT50), .A2(n1048), .ZN(n1235) );
NAND2_X1 U886 ( .A1(KEYINPUT20), .A2(n1241), .ZN(n1231) );
XNOR2_X1 U887 ( .A(G140), .B(n1242), .ZN(G42) );
NOR2_X1 U888 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NOR3_X1 U889 ( .A1(n1245), .A2(n1246), .A3(n1062), .ZN(n1244) );
INV_X1 U890 ( .A(KEYINPUT56), .ZN(n1245) );
NOR2_X1 U891 ( .A1(KEYINPUT56), .A2(n1207), .ZN(n1243) );
NAND2_X1 U892 ( .A1(n1246), .A2(n1073), .ZN(n1207) );
INV_X1 U893 ( .A(n1062), .ZN(n1073) );
AND2_X1 U894 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND3_X1 U895 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(G39) );
NAND2_X1 U896 ( .A1(G137), .A2(n1252), .ZN(n1251) );
NAND2_X1 U897 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
INV_X1 U898 ( .A(KEYINPUT4), .ZN(n1254) );
XNOR2_X1 U899 ( .A(n1205), .B(KEYINPUT15), .ZN(n1253) );
INV_X1 U900 ( .A(n1255), .ZN(n1205) );
OR3_X1 U901 ( .A1(n1255), .A2(G137), .A3(KEYINPUT4), .ZN(n1250) );
NAND2_X1 U902 ( .A1(KEYINPUT4), .A2(n1255), .ZN(n1249) );
NAND4_X1 U903 ( .A1(n1256), .A2(n1066), .A3(n1248), .A4(n1257), .ZN(n1255) );
NOR3_X1 U904 ( .A1(n1234), .A2(n1062), .A3(n1093), .ZN(n1257) );
XOR2_X1 U905 ( .A(n1201), .B(n1258), .Z(G36) );
NOR2_X1 U906 ( .A1(KEYINPUT38), .A2(n1259), .ZN(n1258) );
INV_X1 U907 ( .A(G134), .ZN(n1259) );
AND2_X1 U908 ( .A1(n1260), .A2(n1048), .ZN(n1201) );
XOR2_X1 U909 ( .A(G131), .B(n1200), .Z(G33) );
AND2_X1 U910 ( .A1(n1049), .A2(n1260), .ZN(n1200) );
NOR4_X1 U911 ( .A1(n1234), .A2(n1062), .A3(n1075), .A4(n1261), .ZN(n1260) );
NAND2_X1 U912 ( .A1(n1262), .A2(n1060), .ZN(n1062) );
INV_X1 U913 ( .A(n1059), .ZN(n1262) );
XOR2_X1 U914 ( .A(G128), .B(n1199), .Z(G30) );
AND2_X1 U915 ( .A1(n1230), .A2(n1048), .ZN(n1199) );
NOR4_X1 U916 ( .A1(n1234), .A2(n1209), .A3(n1065), .A4(n1263), .ZN(n1230) );
XNOR2_X1 U917 ( .A(G101), .B(n1212), .ZN(G3) );
NAND4_X1 U918 ( .A1(n1052), .A2(n1232), .A3(n1264), .A4(n1064), .ZN(n1212) );
XOR2_X1 U919 ( .A(G125), .B(n1204), .Z(G27) );
AND3_X1 U920 ( .A1(n1247), .A2(n1058), .A3(n1265), .ZN(n1204) );
NOR4_X1 U921 ( .A1(n1219), .A2(n1234), .A3(n1066), .A4(n1065), .ZN(n1247) );
INV_X1 U922 ( .A(n1256), .ZN(n1065) );
NAND2_X1 U923 ( .A1(n1266), .A2(n1050), .ZN(n1234) );
NAND2_X1 U924 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
OR2_X1 U925 ( .A1(n1109), .A2(n1195), .ZN(n1268) );
NAND2_X1 U926 ( .A1(n1269), .A2(n1124), .ZN(n1109) );
XOR2_X1 U927 ( .A(KEYINPUT55), .B(G900), .Z(n1269) );
XOR2_X1 U928 ( .A(n1270), .B(n1271), .Z(G24) );
NOR2_X1 U929 ( .A1(n1222), .A2(n1226), .ZN(n1271) );
NAND4_X1 U930 ( .A1(n1272), .A2(n1265), .A3(n1273), .A4(n1074), .ZN(n1226) );
NOR2_X1 U931 ( .A1(n1239), .A2(n1208), .ZN(n1273) );
INV_X1 U932 ( .A(n1043), .ZN(n1265) );
XNOR2_X1 U933 ( .A(KEYINPUT50), .B(n1274), .ZN(n1272) );
NAND2_X1 U934 ( .A1(KEYINPUT11), .A2(n1275), .ZN(n1270) );
XNOR2_X1 U935 ( .A(G119), .B(n1210), .ZN(G21) );
OR4_X1 U936 ( .A1(n1228), .A2(n1043), .A3(n1222), .A4(n1263), .ZN(n1210) );
XNOR2_X1 U937 ( .A(G116), .B(n1211), .ZN(G18) );
NAND3_X1 U938 ( .A1(n1048), .A2(n1058), .A3(n1276), .ZN(n1211) );
NOR2_X1 U939 ( .A1(n1274), .A2(n1239), .ZN(n1048) );
XNOR2_X1 U940 ( .A(G113), .B(n1277), .ZN(G15) );
NAND2_X1 U941 ( .A1(n1225), .A2(n1058), .ZN(n1277) );
INV_X1 U942 ( .A(n1222), .ZN(n1058) );
AND2_X1 U943 ( .A1(n1276), .A2(n1049), .ZN(n1225) );
INV_X1 U944 ( .A(n1219), .ZN(n1049) );
NAND2_X1 U945 ( .A1(n1239), .A2(n1274), .ZN(n1219) );
NOR3_X1 U946 ( .A1(n1208), .A2(n1261), .A3(n1043), .ZN(n1276) );
NAND2_X1 U947 ( .A1(n1078), .A2(n1278), .ZN(n1043) );
INV_X1 U948 ( .A(n1064), .ZN(n1261) );
NAND2_X1 U949 ( .A1(n1279), .A2(n1280), .ZN(n1064) );
OR3_X1 U950 ( .A1(n1256), .A2(n1263), .A3(KEYINPUT47), .ZN(n1280) );
NAND2_X1 U951 ( .A1(KEYINPUT47), .A2(n1074), .ZN(n1279) );
NOR2_X1 U952 ( .A1(n1066), .A2(n1256), .ZN(n1074) );
XOR2_X1 U953 ( .A(n1281), .B(n1218), .Z(G12) );
NOR3_X1 U954 ( .A1(n1209), .A2(n1066), .A3(n1228), .ZN(n1218) );
NAND3_X1 U955 ( .A1(n1264), .A2(n1256), .A3(n1052), .ZN(n1228) );
INV_X1 U956 ( .A(n1093), .ZN(n1052) );
NAND2_X1 U957 ( .A1(n1239), .A2(n1240), .ZN(n1093) );
INV_X1 U958 ( .A(n1274), .ZN(n1240) );
XNOR2_X1 U959 ( .A(n1282), .B(G475), .ZN(n1274) );
OR2_X1 U960 ( .A1(n1157), .A2(G902), .ZN(n1282) );
XOR2_X1 U961 ( .A(n1283), .B(n1284), .Z(n1157) );
XOR2_X1 U962 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U963 ( .A(G113), .B(G104), .Z(n1286) );
XNOR2_X1 U964 ( .A(KEYINPUT12), .B(n1275), .ZN(n1285) );
INV_X1 U965 ( .A(G122), .ZN(n1275) );
XOR2_X1 U966 ( .A(n1287), .B(n1113), .Z(n1283) );
XOR2_X1 U967 ( .A(G125), .B(n1288), .Z(n1113) );
XOR2_X1 U968 ( .A(n1289), .B(n1290), .Z(n1287) );
NOR2_X1 U969 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U970 ( .A(n1241), .B(n1293), .ZN(n1292) );
AND2_X1 U971 ( .A1(n1294), .A2(G214), .ZN(n1293) );
XNOR2_X1 U972 ( .A(KEYINPUT53), .B(KEYINPUT24), .ZN(n1291) );
NAND2_X1 U973 ( .A1(KEYINPUT45), .A2(n1295), .ZN(n1289) );
XOR2_X1 U974 ( .A(n1296), .B(G478), .Z(n1239) );
NAND2_X1 U975 ( .A1(n1153), .A2(n1195), .ZN(n1296) );
XNOR2_X1 U976 ( .A(n1297), .B(n1298), .ZN(n1153) );
XOR2_X1 U977 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U978 ( .A(n1301), .B(n1302), .ZN(n1300) );
NOR2_X1 U979 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
INV_X1 U980 ( .A(G217), .ZN(n1304) );
XOR2_X1 U981 ( .A(n1305), .B(n1306), .Z(n1297) );
XNOR2_X1 U982 ( .A(KEYINPUT51), .B(n1241), .ZN(n1306) );
INV_X1 U983 ( .A(G143), .ZN(n1241) );
XNOR2_X1 U984 ( .A(G116), .B(G134), .ZN(n1305) );
NAND2_X1 U985 ( .A1(n1307), .A2(n1308), .ZN(n1256) );
NAND2_X1 U986 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
INV_X1 U987 ( .A(KEYINPUT14), .ZN(n1310) );
NAND2_X1 U988 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
NAND2_X1 U989 ( .A1(n1102), .A2(n1101), .ZN(n1312) );
INV_X1 U990 ( .A(n1098), .ZN(n1311) );
NOR2_X1 U991 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U992 ( .A1(KEYINPUT14), .A2(n1313), .ZN(n1307) );
XNOR2_X1 U993 ( .A(n1102), .B(n1149), .ZN(n1313) );
INV_X1 U994 ( .A(n1101), .ZN(n1149) );
NAND2_X1 U995 ( .A1(G217), .A2(n1314), .ZN(n1101) );
NOR2_X1 U996 ( .A1(n1148), .A2(G902), .ZN(n1102) );
XOR2_X1 U997 ( .A(n1315), .B(n1316), .Z(n1148) );
NOR2_X1 U998 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NOR2_X1 U999 ( .A1(KEYINPUT19), .A2(n1319), .ZN(n1318) );
AND2_X1 U1000 ( .A1(KEYINPUT9), .A2(n1319), .ZN(n1317) );
XNOR2_X1 U1001 ( .A(n1320), .B(n1321), .ZN(n1319) );
XOR2_X1 U1002 ( .A(G140), .B(G125), .Z(n1321) );
XNOR2_X1 U1003 ( .A(n1295), .B(n1322), .ZN(n1320) );
NOR2_X1 U1004 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1005 ( .A(n1325), .B(KEYINPUT18), .Z(n1324) );
NAND2_X1 U1006 ( .A1(n1326), .A2(G110), .ZN(n1325) );
NOR2_X1 U1007 ( .A1(G110), .A2(n1326), .ZN(n1323) );
XNOR2_X1 U1008 ( .A(G119), .B(n1301), .ZN(n1326) );
XOR2_X1 U1009 ( .A(G146), .B(KEYINPUT60), .Z(n1295) );
XNOR2_X1 U1010 ( .A(G137), .B(n1327), .ZN(n1315) );
NOR2_X1 U1011 ( .A1(n1303), .A2(n1328), .ZN(n1327) );
INV_X1 U1012 ( .A(G221), .ZN(n1328) );
NAND2_X1 U1013 ( .A1(G234), .A2(n1329), .ZN(n1303) );
INV_X1 U1014 ( .A(n1208), .ZN(n1264) );
NAND2_X1 U1015 ( .A1(n1330), .A2(n1050), .ZN(n1208) );
NAND2_X1 U1016 ( .A1(G237), .A2(n1331), .ZN(n1050) );
NAND2_X1 U1017 ( .A1(n1267), .A2(n1332), .ZN(n1330) );
NAND3_X1 U1018 ( .A1(n1333), .A2(n1125), .A3(G902), .ZN(n1332) );
INV_X1 U1019 ( .A(G898), .ZN(n1125) );
XOR2_X1 U1020 ( .A(KEYINPUT22), .B(n1124), .Z(n1333) );
XNOR2_X1 U1021 ( .A(n1069), .B(KEYINPUT52), .ZN(n1124) );
NAND2_X1 U1022 ( .A1(G952), .A2(n1069), .ZN(n1267) );
INV_X1 U1023 ( .A(n1263), .ZN(n1066) );
NOR2_X1 U1024 ( .A1(n1092), .A2(n1334), .ZN(n1263) );
AND2_X1 U1025 ( .A1(n1096), .A2(n1095), .ZN(n1334) );
NOR2_X1 U1026 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
AND2_X1 U1027 ( .A1(n1335), .A2(n1195), .ZN(n1096) );
XNOR2_X1 U1028 ( .A(n1336), .B(n1166), .ZN(n1335) );
XNOR2_X1 U1029 ( .A(n1337), .B(n1338), .ZN(n1166) );
XNOR2_X1 U1030 ( .A(n1339), .B(n1340), .ZN(n1338) );
XNOR2_X1 U1031 ( .A(n1192), .B(n1341), .ZN(n1337) );
XOR2_X1 U1032 ( .A(G131), .B(n1342), .Z(n1341) );
NOR2_X1 U1033 ( .A1(G116), .A2(KEYINPUT36), .ZN(n1342) );
NAND2_X1 U1034 ( .A1(KEYINPUT43), .A2(n1162), .ZN(n1336) );
AND2_X1 U1035 ( .A1(n1343), .A2(n1344), .ZN(n1162) );
NAND2_X1 U1036 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
INV_X1 U1037 ( .A(G101), .ZN(n1346) );
NAND2_X1 U1038 ( .A1(G210), .A2(n1294), .ZN(n1345) );
NAND3_X1 U1039 ( .A1(G210), .A2(n1294), .A3(G101), .ZN(n1343) );
AND2_X1 U1040 ( .A1(n1329), .A2(n1347), .ZN(n1294) );
INV_X1 U1041 ( .A(G472), .ZN(n1095) );
INV_X1 U1042 ( .A(n1232), .ZN(n1209) );
NOR2_X1 U1043 ( .A1(n1075), .A2(n1222), .ZN(n1232) );
NAND2_X1 U1044 ( .A1(n1059), .A2(n1060), .ZN(n1222) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1348), .ZN(n1060) );
XNOR2_X1 U1046 ( .A(n1349), .B(n1194), .ZN(n1059) );
AND2_X1 U1047 ( .A1(G210), .A2(n1348), .ZN(n1194) );
NAND2_X1 U1048 ( .A1(n1347), .A2(n1195), .ZN(n1348) );
INV_X1 U1049 ( .A(G237), .ZN(n1347) );
NAND2_X1 U1050 ( .A1(n1350), .A2(n1195), .ZN(n1349) );
XOR2_X1 U1051 ( .A(n1186), .B(n1351), .Z(n1350) );
XNOR2_X1 U1052 ( .A(KEYINPUT13), .B(n1190), .ZN(n1351) );
INV_X1 U1053 ( .A(n1192), .ZN(n1190) );
XNOR2_X1 U1054 ( .A(n1352), .B(n1353), .ZN(n1192) );
XNOR2_X1 U1055 ( .A(n1229), .B(n1301), .ZN(n1353) );
XOR2_X1 U1056 ( .A(n1354), .B(n1355), .Z(n1186) );
XOR2_X1 U1057 ( .A(n1356), .B(n1357), .Z(n1355) );
XNOR2_X1 U1058 ( .A(G125), .B(G110), .ZN(n1357) );
NAND2_X1 U1059 ( .A1(G224), .A2(n1329), .ZN(n1356) );
XNOR2_X1 U1060 ( .A(n1358), .B(n1136), .ZN(n1354) );
INV_X1 U1061 ( .A(n1132), .ZN(n1136) );
XOR2_X1 U1062 ( .A(G116), .B(n1340), .Z(n1132) );
XOR2_X1 U1063 ( .A(G113), .B(G119), .Z(n1340) );
XOR2_X1 U1064 ( .A(n1299), .B(n1141), .Z(n1358) );
XNOR2_X1 U1065 ( .A(n1359), .B(KEYINPUT2), .ZN(n1141) );
XNOR2_X1 U1066 ( .A(G107), .B(G122), .ZN(n1299) );
INV_X1 U1067 ( .A(n1248), .ZN(n1075) );
NOR2_X1 U1068 ( .A1(n1360), .A2(n1078), .ZN(n1248) );
NOR2_X1 U1069 ( .A1(n1361), .A2(n1091), .ZN(n1078) );
NOR2_X1 U1070 ( .A1(n1362), .A2(G469), .ZN(n1091) );
XNOR2_X1 U1071 ( .A(KEYINPUT17), .B(n1090), .ZN(n1361) );
AND2_X1 U1072 ( .A1(G469), .A2(n1362), .ZN(n1090) );
NAND2_X1 U1073 ( .A1(n1363), .A2(n1195), .ZN(n1362) );
XOR2_X1 U1074 ( .A(n1181), .B(n1364), .Z(n1363) );
XOR2_X1 U1075 ( .A(n1365), .B(n1112), .Z(n1364) );
XOR2_X1 U1076 ( .A(n1352), .B(n1366), .Z(n1112) );
XNOR2_X1 U1077 ( .A(n1367), .B(n1368), .ZN(n1366) );
NOR2_X1 U1078 ( .A1(KEYINPUT31), .A2(n1369), .ZN(n1368) );
INV_X1 U1079 ( .A(n1301), .ZN(n1369) );
XOR2_X1 U1080 ( .A(G128), .B(KEYINPUT29), .Z(n1301) );
NAND2_X1 U1081 ( .A1(KEYINPUT30), .A2(n1229), .ZN(n1367) );
INV_X1 U1082 ( .A(G146), .ZN(n1229) );
XNOR2_X1 U1083 ( .A(G143), .B(KEYINPUT0), .ZN(n1352) );
NAND2_X1 U1084 ( .A1(KEYINPUT32), .A2(n1179), .ZN(n1365) );
XNOR2_X1 U1085 ( .A(n1370), .B(n1371), .ZN(n1181) );
XOR2_X1 U1086 ( .A(n1372), .B(n1373), .Z(n1371) );
XOR2_X1 U1087 ( .A(n1374), .B(KEYINPUT63), .Z(n1373) );
NAND2_X1 U1088 ( .A1(G227), .A2(n1375), .ZN(n1374) );
XOR2_X1 U1089 ( .A(KEYINPUT39), .B(n1329), .Z(n1375) );
XNOR2_X1 U1090 ( .A(n1069), .B(KEYINPUT62), .ZN(n1329) );
INV_X1 U1091 ( .A(G953), .ZN(n1069) );
NAND2_X1 U1092 ( .A1(KEYINPUT34), .A2(n1034), .ZN(n1372) );
INV_X1 U1093 ( .A(G107), .ZN(n1034) );
XNOR2_X1 U1094 ( .A(n1288), .B(n1376), .ZN(n1370) );
XOR2_X1 U1095 ( .A(n1339), .B(n1359), .Z(n1376) );
XNOR2_X1 U1096 ( .A(G104), .B(G101), .ZN(n1359) );
XNOR2_X1 U1097 ( .A(G137), .B(n1377), .ZN(n1339) );
NOR2_X1 U1098 ( .A1(G134), .A2(KEYINPUT26), .ZN(n1377) );
XOR2_X1 U1099 ( .A(G131), .B(G140), .Z(n1288) );
INV_X1 U1100 ( .A(n1278), .ZN(n1360) );
XNOR2_X1 U1101 ( .A(n1079), .B(KEYINPUT37), .ZN(n1278) );
AND2_X1 U1102 ( .A1(G221), .A2(n1314), .ZN(n1079) );
NAND2_X1 U1103 ( .A1(n1331), .A2(n1195), .ZN(n1314) );
INV_X1 U1104 ( .A(G902), .ZN(n1195) );
XNOR2_X1 U1105 ( .A(G234), .B(KEYINPUT42), .ZN(n1331) );
NAND2_X1 U1106 ( .A1(KEYINPUT54), .A2(n1179), .ZN(n1281) );
INV_X1 U1107 ( .A(G110), .ZN(n1179) );
endmodule


