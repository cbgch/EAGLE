//Key = 1101100111101101110101011101010010100001000110001010000101110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390;

XNOR2_X1 U767 ( .A(G107), .B(n1058), .ZN(G9) );
NOR2_X1 U768 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR3_X1 U769 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR2_X1 U770 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
XOR2_X1 U771 ( .A(n1066), .B(KEYINPUT11), .Z(n1064) );
NAND3_X1 U772 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1061) );
NAND3_X1 U773 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U774 ( .A1(n1073), .A2(n1066), .ZN(n1071) );
NAND4_X1 U775 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1066) );
NAND2_X1 U776 ( .A1(n1078), .A2(n1079), .ZN(n1070) );
NAND2_X1 U777 ( .A1(n1080), .A2(n1077), .ZN(n1078) );
NAND2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U779 ( .A1(n1076), .A2(n1083), .ZN(n1082) );
NAND2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U781 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U782 ( .A(n1075), .B(KEYINPUT0), .ZN(n1086) );
NAND2_X1 U783 ( .A1(n1075), .A2(n1088), .ZN(n1084) );
NAND2_X1 U784 ( .A1(n1074), .A2(n1089), .ZN(n1081) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U786 ( .A1(n1076), .A2(n1092), .ZN(n1091) );
OR2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U788 ( .A1(n1075), .A2(n1095), .ZN(n1090) );
NAND3_X1 U789 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
OR3_X1 U790 ( .A1(n1099), .A2(n1100), .A3(KEYINPUT2), .ZN(n1097) );
NAND2_X1 U791 ( .A1(KEYINPUT2), .A2(n1100), .ZN(n1096) );
NOR3_X1 U792 ( .A1(n1101), .A2(G953), .A3(G952), .ZN(n1059) );
INV_X1 U793 ( .A(n1067), .ZN(n1101) );
NAND4_X1 U794 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1067) );
NOR3_X1 U795 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
XOR2_X1 U796 ( .A(n1109), .B(KEYINPUT5), .Z(n1108) );
NAND4_X1 U797 ( .A1(n1110), .A2(n1111), .A3(n1099), .A4(n1079), .ZN(n1109) );
XOR2_X1 U798 ( .A(n1112), .B(n1113), .Z(n1111) );
NAND2_X1 U799 ( .A1(KEYINPUT29), .A2(n1114), .ZN(n1113) );
XOR2_X1 U800 ( .A(n1115), .B(n1116), .Z(n1110) );
XOR2_X1 U801 ( .A(KEYINPUT6), .B(G469), .Z(n1116) );
NOR2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(n1107) );
XOR2_X1 U803 ( .A(n1119), .B(KEYINPUT17), .Z(n1106) );
XOR2_X1 U804 ( .A(n1120), .B(KEYINPUT28), .Z(n1104) );
NAND2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1120) );
INV_X1 U806 ( .A(G478), .ZN(n1118) );
XOR2_X1 U807 ( .A(n1121), .B(KEYINPUT54), .Z(n1102) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(G72) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1068), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U812 ( .A1(n1129), .A2(n1130), .ZN(n1124) );
NAND2_X1 U813 ( .A1(G953), .A2(n1128), .ZN(n1130) );
XOR2_X1 U814 ( .A(n1131), .B(n1132), .Z(n1129) );
XOR2_X1 U815 ( .A(G134), .B(n1133), .Z(n1132) );
XNOR2_X1 U816 ( .A(n1134), .B(n1135), .ZN(n1131) );
NAND2_X1 U817 ( .A1(n1068), .A2(n1136), .ZN(n1122) );
NAND2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(G69) );
XOR2_X1 U820 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U821 ( .A1(n1068), .A2(n1143), .ZN(n1142) );
NAND2_X1 U822 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XNOR2_X1 U823 ( .A(n1146), .B(KEYINPUT25), .ZN(n1144) );
NAND3_X1 U824 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1141) );
NAND2_X1 U825 ( .A1(n1150), .A2(G953), .ZN(n1149) );
XOR2_X1 U826 ( .A(n1151), .B(KEYINPUT60), .Z(n1150) );
OR2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
NAND2_X1 U828 ( .A1(n1152), .A2(n1154), .ZN(n1147) );
NAND2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U830 ( .A1(KEYINPUT10), .A2(n1153), .ZN(n1156) );
OR2_X1 U831 ( .A1(KEYINPUT18), .A2(n1157), .ZN(n1153) );
OR2_X1 U832 ( .A1(n1157), .A2(KEYINPUT10), .ZN(n1155) );
XNOR2_X1 U833 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR2_X1 U834 ( .A1(n1160), .A2(n1068), .ZN(n1139) );
NOR2_X1 U835 ( .A1(n1161), .A2(n1151), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1162), .A2(n1163), .ZN(G66) );
XOR2_X1 U837 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U838 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
NOR2_X1 U839 ( .A1(n1162), .A2(n1168), .ZN(G63) );
XOR2_X1 U840 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U841 ( .A(n1171), .B(KEYINPUT33), .ZN(n1170) );
NAND3_X1 U842 ( .A1(n1172), .A2(G478), .A3(KEYINPUT58), .ZN(n1171) );
NOR2_X1 U843 ( .A1(n1162), .A2(n1173), .ZN(G60) );
XOR2_X1 U844 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND3_X1 U845 ( .A1(G475), .A2(n1176), .A3(n1177), .ZN(n1174) );
XOR2_X1 U846 ( .A(n1063), .B(KEYINPUT49), .Z(n1177) );
XNOR2_X1 U847 ( .A(G104), .B(n1178), .ZN(G6) );
NOR2_X1 U848 ( .A1(n1162), .A2(n1179), .ZN(G57) );
XOR2_X1 U849 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U850 ( .A(G101), .B(n1182), .ZN(n1181) );
NAND2_X1 U851 ( .A1(n1183), .A2(n1184), .ZN(n1180) );
NAND4_X1 U852 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
AND2_X1 U853 ( .A1(n1189), .A2(G472), .ZN(n1188) );
NAND2_X1 U854 ( .A1(n1190), .A2(n1191), .ZN(n1183) );
NAND3_X1 U855 ( .A1(n1185), .A2(n1186), .A3(G472), .ZN(n1191) );
NAND2_X1 U856 ( .A1(n1167), .A2(n1192), .ZN(n1186) );
INV_X1 U857 ( .A(KEYINPUT36), .ZN(n1192) );
NAND2_X1 U858 ( .A1(KEYINPUT36), .A2(n1193), .ZN(n1185) );
NAND2_X1 U859 ( .A1(n1194), .A2(n1063), .ZN(n1193) );
NAND2_X1 U860 ( .A1(n1187), .A2(n1189), .ZN(n1190) );
INV_X1 U861 ( .A(n1195), .ZN(n1187) );
NOR2_X1 U862 ( .A1(n1162), .A2(n1196), .ZN(G54) );
XOR2_X1 U863 ( .A(n1197), .B(n1198), .Z(n1196) );
XNOR2_X1 U864 ( .A(n1199), .B(n1200), .ZN(n1198) );
XNOR2_X1 U865 ( .A(n1201), .B(n1202), .ZN(n1197) );
NAND3_X1 U866 ( .A1(n1172), .A2(G469), .A3(KEYINPUT15), .ZN(n1202) );
INV_X1 U867 ( .A(n1167), .ZN(n1172) );
NAND2_X1 U868 ( .A1(KEYINPUT59), .A2(n1203), .ZN(n1201) );
NOR2_X1 U869 ( .A1(n1162), .A2(n1204), .ZN(G51) );
XOR2_X1 U870 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U871 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U872 ( .A1(n1112), .A2(n1167), .ZN(n1208) );
NAND2_X1 U873 ( .A1(n1176), .A2(n1063), .ZN(n1167) );
NAND4_X1 U874 ( .A1(n1209), .A2(n1146), .A3(n1137), .A4(n1145), .ZN(n1063) );
AND4_X1 U875 ( .A1(n1178), .A2(n1058), .A3(n1210), .A4(n1211), .ZN(n1145) );
NAND3_X1 U876 ( .A1(n1087), .A2(n1075), .A3(n1212), .ZN(n1058) );
NAND3_X1 U877 ( .A1(n1075), .A2(n1088), .A3(n1212), .ZN(n1178) );
AND4_X1 U878 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1137) );
NOR4_X1 U879 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
INV_X1 U880 ( .A(n1221), .ZN(n1220) );
NAND2_X1 U881 ( .A1(n1222), .A2(n1223), .ZN(n1215) );
XNOR2_X1 U882 ( .A(n1087), .B(KEYINPUT12), .ZN(n1222) );
AND4_X1 U883 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1146) );
NAND3_X1 U884 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1225) );
INV_X1 U885 ( .A(n1231), .ZN(n1230) );
OR2_X1 U886 ( .A1(n1232), .A2(KEYINPUT52), .ZN(n1229) );
NAND2_X1 U887 ( .A1(KEYINPUT52), .A2(n1233), .ZN(n1228) );
NAND3_X1 U888 ( .A1(n1076), .A2(n1065), .A3(n1234), .ZN(n1233) );
NAND3_X1 U889 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1224) );
OR2_X1 U890 ( .A1(n1232), .A2(KEYINPUT20), .ZN(n1236) );
NAND2_X1 U891 ( .A1(KEYINPUT20), .A2(n1238), .ZN(n1235) );
NAND2_X1 U892 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XOR2_X1 U893 ( .A(n1138), .B(KEYINPUT22), .Z(n1209) );
INV_X1 U894 ( .A(n1194), .ZN(n1176) );
XOR2_X1 U895 ( .A(n1241), .B(KEYINPUT46), .Z(n1194) );
NAND3_X1 U896 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1207) );
INV_X1 U897 ( .A(n1245), .ZN(n1244) );
NAND2_X1 U898 ( .A1(n1246), .A2(n1247), .ZN(n1243) );
INV_X1 U899 ( .A(KEYINPUT16), .ZN(n1247) );
XNOR2_X1 U900 ( .A(n1248), .B(n1249), .ZN(n1246) );
NOR2_X1 U901 ( .A1(G125), .A2(n1250), .ZN(n1249) );
NAND2_X1 U902 ( .A1(KEYINPUT16), .A2(n1251), .ZN(n1242) );
NOR2_X1 U903 ( .A1(n1068), .A2(G952), .ZN(n1162) );
XOR2_X1 U904 ( .A(n1213), .B(n1252), .Z(G48) );
NAND2_X1 U905 ( .A1(KEYINPUT24), .A2(G146), .ZN(n1252) );
NAND2_X1 U906 ( .A1(n1223), .A2(n1088), .ZN(n1213) );
XOR2_X1 U907 ( .A(n1253), .B(n1254), .Z(G45) );
XOR2_X1 U908 ( .A(KEYINPUT38), .B(G143), .Z(n1254) );
NAND2_X1 U909 ( .A1(KEYINPUT50), .A2(n1214), .ZN(n1253) );
NAND4_X1 U910 ( .A1(n1093), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1214) );
AND3_X1 U911 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1257) );
XNOR2_X1 U912 ( .A(G140), .B(n1261), .ZN(G42) );
NAND2_X1 U913 ( .A1(KEYINPUT61), .A2(n1219), .ZN(n1261) );
AND3_X1 U914 ( .A1(n1262), .A2(n1088), .A3(n1094), .ZN(n1219) );
XNOR2_X1 U915 ( .A(n1263), .B(n1138), .ZN(G39) );
NAND2_X1 U916 ( .A1(n1262), .A2(n1237), .ZN(n1138) );
INV_X1 U917 ( .A(n1264), .ZN(n1237) );
XOR2_X1 U918 ( .A(n1265), .B(KEYINPUT55), .Z(n1263) );
XOR2_X1 U919 ( .A(G134), .B(n1218), .Z(G36) );
AND3_X1 U920 ( .A1(n1093), .A2(n1087), .A3(n1262), .ZN(n1218) );
XOR2_X1 U921 ( .A(G131), .B(n1217), .Z(G33) );
AND3_X1 U922 ( .A1(n1093), .A2(n1088), .A3(n1262), .ZN(n1217) );
AND4_X1 U923 ( .A1(n1256), .A2(n1258), .A3(n1072), .A4(n1079), .ZN(n1262) );
XOR2_X1 U924 ( .A(G128), .B(n1266), .Z(G30) );
AND2_X1 U925 ( .A1(n1087), .A2(n1223), .ZN(n1266) );
AND3_X1 U926 ( .A1(n1256), .A2(n1255), .A3(n1267), .ZN(n1223) );
NOR3_X1 U927 ( .A1(n1098), .A2(n1119), .A3(n1121), .ZN(n1267) );
XNOR2_X1 U928 ( .A(G101), .B(n1210), .ZN(G3) );
NAND3_X1 U929 ( .A1(n1074), .A2(n1212), .A3(n1093), .ZN(n1210) );
XOR2_X1 U930 ( .A(n1268), .B(n1221), .Z(G27) );
NAND4_X1 U931 ( .A1(n1094), .A2(n1256), .A3(n1239), .A4(n1088), .ZN(n1221) );
AND2_X1 U932 ( .A1(n1269), .A2(n1077), .ZN(n1256) );
NAND2_X1 U933 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND3_X1 U934 ( .A1(G902), .A2(n1128), .A3(G953), .ZN(n1271) );
INV_X1 U935 ( .A(G900), .ZN(n1128) );
XOR2_X1 U936 ( .A(G122), .B(n1272), .Z(G24) );
NOR3_X1 U937 ( .A1(n1231), .A2(KEYINPUT37), .A3(n1273), .ZN(n1272) );
NAND3_X1 U938 ( .A1(n1260), .A2(n1259), .A3(n1075), .ZN(n1231) );
NOR2_X1 U939 ( .A1(n1274), .A2(n1275), .ZN(n1075) );
XOR2_X1 U940 ( .A(KEYINPUT47), .B(n1276), .Z(n1260) );
XOR2_X1 U941 ( .A(G119), .B(n1277), .Z(G21) );
NOR2_X1 U942 ( .A1(n1273), .A2(n1264), .ZN(n1277) );
NAND3_X1 U943 ( .A1(n1275), .A2(n1274), .A3(n1074), .ZN(n1264) );
XOR2_X1 U944 ( .A(n1278), .B(n1226), .Z(G18) );
NAND3_X1 U945 ( .A1(n1093), .A2(n1087), .A3(n1232), .ZN(n1226) );
AND2_X1 U946 ( .A1(n1103), .A2(n1259), .ZN(n1087) );
XOR2_X1 U947 ( .A(n1279), .B(n1227), .Z(G15) );
NAND3_X1 U948 ( .A1(n1093), .A2(n1088), .A3(n1232), .ZN(n1227) );
INV_X1 U949 ( .A(n1273), .ZN(n1232) );
NAND2_X1 U950 ( .A1(n1239), .A2(n1234), .ZN(n1273) );
INV_X1 U951 ( .A(n1240), .ZN(n1234) );
AND2_X1 U952 ( .A1(n1255), .A2(n1076), .ZN(n1239) );
NAND2_X1 U953 ( .A1(n1280), .A2(n1281), .ZN(n1076) );
OR3_X1 U954 ( .A1(n1100), .A2(n1282), .A3(KEYINPUT2), .ZN(n1281) );
INV_X1 U955 ( .A(n1099), .ZN(n1282) );
NAND2_X1 U956 ( .A1(KEYINPUT2), .A2(n1258), .ZN(n1280) );
INV_X1 U957 ( .A(n1098), .ZN(n1258) );
NAND2_X1 U958 ( .A1(n1283), .A2(n1284), .ZN(n1088) );
OR3_X1 U959 ( .A1(n1103), .A2(n1259), .A3(KEYINPUT47), .ZN(n1284) );
NAND2_X1 U960 ( .A1(KEYINPUT47), .A2(n1074), .ZN(n1283) );
NOR2_X1 U961 ( .A1(n1274), .A2(n1121), .ZN(n1093) );
INV_X1 U962 ( .A(n1119), .ZN(n1274) );
XNOR2_X1 U963 ( .A(n1285), .B(n1211), .ZN(G12) );
NAND3_X1 U964 ( .A1(n1074), .A2(n1212), .A3(n1094), .ZN(n1211) );
NOR2_X1 U965 ( .A1(n1275), .A2(n1119), .ZN(n1094) );
XNOR2_X1 U966 ( .A(n1286), .B(n1166), .ZN(n1119) );
NAND2_X1 U967 ( .A1(G217), .A2(n1287), .ZN(n1166) );
OR2_X1 U968 ( .A1(n1165), .A2(G902), .ZN(n1286) );
XNOR2_X1 U969 ( .A(n1288), .B(n1289), .ZN(n1165) );
XOR2_X1 U970 ( .A(n1265), .B(n1290), .Z(n1289) );
XNOR2_X1 U971 ( .A(KEYINPUT39), .B(KEYINPUT13), .ZN(n1290) );
XOR2_X1 U972 ( .A(n1291), .B(n1292), .Z(n1288) );
XOR2_X1 U973 ( .A(n1293), .B(n1294), .Z(n1291) );
AND3_X1 U974 ( .A1(n1295), .A2(n1068), .A3(G221), .ZN(n1294) );
NAND4_X1 U975 ( .A1(n1296), .A2(n1297), .A3(n1298), .A4(n1299), .ZN(n1293) );
NAND3_X1 U976 ( .A1(KEYINPUT35), .A2(n1300), .A3(n1301), .ZN(n1299) );
OR2_X1 U977 ( .A1(n1302), .A2(KEYINPUT3), .ZN(n1300) );
OR3_X1 U978 ( .A1(n1303), .A2(KEYINPUT35), .A3(n1301), .ZN(n1298) );
AND2_X1 U979 ( .A1(KEYINPUT3), .A2(n1203), .ZN(n1303) );
NAND2_X1 U980 ( .A1(KEYINPUT51), .A2(n1302), .ZN(n1297) );
NAND3_X1 U981 ( .A1(n1304), .A2(n1305), .A3(n1203), .ZN(n1296) );
INV_X1 U982 ( .A(KEYINPUT51), .ZN(n1305) );
XNOR2_X1 U983 ( .A(KEYINPUT3), .B(n1301), .ZN(n1304) );
NAND2_X1 U984 ( .A1(n1306), .A2(n1307), .ZN(n1301) );
NAND2_X1 U985 ( .A1(G128), .A2(n1308), .ZN(n1307) );
XOR2_X1 U986 ( .A(n1309), .B(KEYINPUT41), .Z(n1306) );
NAND2_X1 U987 ( .A1(G119), .A2(n1310), .ZN(n1309) );
INV_X1 U988 ( .A(n1121), .ZN(n1275) );
XOR2_X1 U989 ( .A(n1311), .B(G472), .Z(n1121) );
NAND2_X1 U990 ( .A1(n1312), .A2(n1241), .ZN(n1311) );
XNOR2_X1 U991 ( .A(n1313), .B(n1182), .ZN(n1312) );
NAND3_X1 U992 ( .A1(n1314), .A2(n1068), .A3(G210), .ZN(n1182) );
XOR2_X1 U993 ( .A(KEYINPUT8), .B(G237), .Z(n1314) );
XOR2_X1 U994 ( .A(n1315), .B(n1316), .Z(n1313) );
NOR2_X1 U995 ( .A1(KEYINPUT53), .A2(G101), .ZN(n1316) );
NAND3_X1 U996 ( .A1(n1317), .A2(n1318), .A3(n1189), .ZN(n1315) );
OR3_X1 U997 ( .A1(n1250), .A2(n1319), .A3(n1320), .ZN(n1189) );
NAND2_X1 U998 ( .A1(n1321), .A2(n1322), .ZN(n1318) );
INV_X1 U999 ( .A(KEYINPUT19), .ZN(n1322) );
XOR2_X1 U1000 ( .A(n1323), .B(n1319), .Z(n1321) );
NAND2_X1 U1001 ( .A1(n1320), .A2(n1250), .ZN(n1323) );
NAND2_X1 U1002 ( .A1(KEYINPUT19), .A2(n1195), .ZN(n1317) );
NAND2_X1 U1003 ( .A1(n1324), .A2(n1325), .ZN(n1195) );
NAND2_X1 U1004 ( .A1(n1326), .A2(n1250), .ZN(n1325) );
INV_X1 U1005 ( .A(n1327), .ZN(n1250) );
XOR2_X1 U1006 ( .A(n1320), .B(n1319), .Z(n1326) );
NAND3_X1 U1007 ( .A1(n1320), .A2(n1319), .A3(n1327), .ZN(n1324) );
XOR2_X1 U1008 ( .A(n1328), .B(G113), .Z(n1319) );
NAND3_X1 U1009 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1328) );
OR2_X1 U1010 ( .A1(n1278), .A2(KEYINPUT1), .ZN(n1331) );
NAND3_X1 U1011 ( .A1(KEYINPUT1), .A2(n1278), .A3(G119), .ZN(n1330) );
INV_X1 U1012 ( .A(G116), .ZN(n1278) );
NAND2_X1 U1013 ( .A1(n1332), .A2(n1308), .ZN(n1329) );
INV_X1 U1014 ( .A(G119), .ZN(n1308) );
NAND2_X1 U1015 ( .A1(KEYINPUT1), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1016 ( .A(KEYINPUT4), .B(G116), .Z(n1333) );
NOR3_X1 U1017 ( .A1(n1098), .A2(n1240), .A3(n1065), .ZN(n1212) );
INV_X1 U1018 ( .A(n1255), .ZN(n1065) );
NOR2_X1 U1019 ( .A1(n1072), .A2(n1073), .ZN(n1255) );
INV_X1 U1020 ( .A(n1079), .ZN(n1073) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1334), .ZN(n1079) );
XOR2_X1 U1022 ( .A(n1335), .B(n1112), .Z(n1072) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1334), .ZN(n1112) );
NAND2_X1 U1024 ( .A1(n1336), .A2(n1241), .ZN(n1334) );
XOR2_X1 U1025 ( .A(n1114), .B(KEYINPUT21), .Z(n1335) );
NAND2_X1 U1026 ( .A1(n1337), .A2(n1241), .ZN(n1114) );
XOR2_X1 U1027 ( .A(n1205), .B(n1338), .Z(n1337) );
XOR2_X1 U1028 ( .A(KEYINPUT31), .B(n1339), .Z(n1338) );
NOR2_X1 U1029 ( .A1(n1245), .A2(n1251), .ZN(n1339) );
NAND2_X1 U1030 ( .A1(n1340), .A2(n1341), .ZN(n1251) );
NAND2_X1 U1031 ( .A1(n1342), .A2(n1268), .ZN(n1341) );
XOR2_X1 U1032 ( .A(n1248), .B(n1327), .Z(n1342) );
NAND3_X1 U1033 ( .A1(n1248), .A2(n1327), .A3(G125), .ZN(n1340) );
NOR3_X1 U1034 ( .A1(n1327), .A2(n1248), .A3(n1268), .ZN(n1245) );
INV_X1 U1035 ( .A(G125), .ZN(n1268) );
NOR2_X1 U1036 ( .A1(n1161), .A2(G953), .ZN(n1248) );
INV_X1 U1037 ( .A(G224), .ZN(n1161) );
XNOR2_X1 U1038 ( .A(n1343), .B(n1344), .ZN(n1327) );
XOR2_X1 U1039 ( .A(n1310), .B(KEYINPUT43), .Z(n1343) );
INV_X1 U1040 ( .A(G128), .ZN(n1310) );
XOR2_X1 U1041 ( .A(n1345), .B(n1152), .Z(n1205) );
XNOR2_X1 U1042 ( .A(n1346), .B(n1203), .ZN(n1152) );
INV_X1 U1043 ( .A(G122), .ZN(n1346) );
XOR2_X1 U1044 ( .A(n1158), .B(n1347), .Z(n1345) );
NOR2_X1 U1045 ( .A1(KEYINPUT14), .A2(n1159), .ZN(n1347) );
XNOR2_X1 U1046 ( .A(n1348), .B(n1349), .ZN(n1159) );
XNOR2_X1 U1047 ( .A(G104), .B(KEYINPUT23), .ZN(n1348) );
XOR2_X1 U1048 ( .A(n1350), .B(n1351), .Z(n1158) );
XOR2_X1 U1049 ( .A(KEYINPUT32), .B(G119), .Z(n1351) );
XOR2_X1 U1050 ( .A(n1279), .B(G116), .Z(n1350) );
NAND2_X1 U1051 ( .A1(n1077), .A2(n1352), .ZN(n1240) );
NAND2_X1 U1052 ( .A1(n1353), .A2(n1270), .ZN(n1352) );
NAND2_X1 U1053 ( .A1(n1354), .A2(n1068), .ZN(n1270) );
XOR2_X1 U1054 ( .A(KEYINPUT42), .B(G952), .Z(n1354) );
NAND3_X1 U1055 ( .A1(G902), .A2(n1151), .A3(G953), .ZN(n1353) );
INV_X1 U1056 ( .A(G898), .ZN(n1151) );
NAND2_X1 U1057 ( .A1(G237), .A2(G234), .ZN(n1077) );
NAND2_X1 U1058 ( .A1(n1100), .A2(n1099), .ZN(n1098) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1287), .ZN(n1099) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1241), .ZN(n1287) );
XNOR2_X1 U1061 ( .A(n1115), .B(n1355), .ZN(n1100) );
NOR2_X1 U1062 ( .A1(KEYINPUT40), .A2(n1356), .ZN(n1355) );
INV_X1 U1063 ( .A(G469), .ZN(n1356) );
NAND2_X1 U1064 ( .A1(n1357), .A2(n1241), .ZN(n1115) );
XOR2_X1 U1065 ( .A(n1358), .B(n1359), .Z(n1357) );
XOR2_X1 U1066 ( .A(n1203), .B(n1200), .Z(n1359) );
XOR2_X1 U1067 ( .A(G140), .B(n1360), .Z(n1200) );
NOR2_X1 U1068 ( .A1(G953), .A2(n1127), .ZN(n1360) );
INV_X1 U1069 ( .A(G227), .ZN(n1127) );
INV_X1 U1070 ( .A(n1302), .ZN(n1203) );
XOR2_X1 U1071 ( .A(n1361), .B(KEYINPUT57), .Z(n1302) );
NOR2_X1 U1072 ( .A1(n1362), .A2(n1363), .ZN(n1358) );
AND2_X1 U1073 ( .A1(KEYINPUT62), .A2(n1199), .ZN(n1363) );
NOR2_X1 U1074 ( .A1(KEYINPUT44), .A2(n1199), .ZN(n1362) );
XOR2_X1 U1075 ( .A(n1364), .B(n1365), .Z(n1199) );
XOR2_X1 U1076 ( .A(n1135), .B(n1349), .Z(n1365) );
XOR2_X1 U1077 ( .A(G107), .B(G101), .Z(n1349) );
XOR2_X1 U1078 ( .A(G128), .B(n1366), .Z(n1135) );
NOR2_X1 U1079 ( .A1(KEYINPUT56), .A2(n1344), .ZN(n1366) );
XNOR2_X1 U1080 ( .A(G146), .B(G143), .ZN(n1344) );
XOR2_X1 U1081 ( .A(n1367), .B(n1320), .Z(n1364) );
XOR2_X1 U1082 ( .A(n1133), .B(n1368), .Z(n1320) );
NOR2_X1 U1083 ( .A1(G134), .A2(KEYINPUT45), .ZN(n1368) );
XOR2_X1 U1084 ( .A(n1369), .B(n1265), .Z(n1133) );
INV_X1 U1085 ( .A(G137), .ZN(n1265) );
INV_X1 U1086 ( .A(G131), .ZN(n1369) );
NAND2_X1 U1087 ( .A1(KEYINPUT63), .A2(G104), .ZN(n1367) );
NOR2_X1 U1088 ( .A1(n1259), .A2(n1276), .ZN(n1074) );
INV_X1 U1089 ( .A(n1103), .ZN(n1276) );
XOR2_X1 U1090 ( .A(n1370), .B(G475), .Z(n1103) );
NAND2_X1 U1091 ( .A1(n1175), .A2(n1241), .ZN(n1370) );
XOR2_X1 U1092 ( .A(n1371), .B(n1372), .Z(n1175) );
XOR2_X1 U1093 ( .A(n1373), .B(n1374), .Z(n1372) );
XOR2_X1 U1094 ( .A(G131), .B(n1375), .Z(n1374) );
NOR2_X1 U1095 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
XOR2_X1 U1096 ( .A(n1378), .B(KEYINPUT7), .Z(n1377) );
NAND2_X1 U1097 ( .A1(n1379), .A2(n1380), .ZN(n1378) );
XNOR2_X1 U1098 ( .A(G104), .B(KEYINPUT9), .ZN(n1379) );
NOR2_X1 U1099 ( .A1(G104), .A2(n1380), .ZN(n1376) );
XOR2_X1 U1100 ( .A(n1381), .B(G122), .Z(n1380) );
NAND2_X1 U1101 ( .A1(KEYINPUT34), .A2(n1279), .ZN(n1381) );
INV_X1 U1102 ( .A(G113), .ZN(n1279) );
AND3_X1 U1103 ( .A1(G214), .A2(n1068), .A3(n1336), .ZN(n1373) );
INV_X1 U1104 ( .A(G237), .ZN(n1336) );
XNOR2_X1 U1105 ( .A(n1292), .B(n1382), .ZN(n1371) );
NOR2_X1 U1106 ( .A1(G143), .A2(KEYINPUT30), .ZN(n1382) );
XOR2_X1 U1107 ( .A(G146), .B(n1134), .Z(n1292) );
XOR2_X1 U1108 ( .A(G140), .B(G125), .Z(n1134) );
XOR2_X1 U1109 ( .A(n1117), .B(G478), .Z(n1259) );
AND2_X1 U1110 ( .A1(n1383), .A2(n1241), .ZN(n1117) );
INV_X1 U1111 ( .A(G902), .ZN(n1241) );
XOR2_X1 U1112 ( .A(KEYINPUT26), .B(n1384), .Z(n1383) );
INV_X1 U1113 ( .A(n1169), .ZN(n1384) );
XOR2_X1 U1114 ( .A(n1385), .B(n1386), .Z(n1169) );
XOR2_X1 U1115 ( .A(n1387), .B(n1388), .Z(n1386) );
XOR2_X1 U1116 ( .A(G128), .B(G122), .Z(n1388) );
XOR2_X1 U1117 ( .A(G143), .B(G134), .Z(n1387) );
XOR2_X1 U1118 ( .A(n1389), .B(n1390), .Z(n1385) );
XOR2_X1 U1119 ( .A(G116), .B(G107), .Z(n1390) );
NAND3_X1 U1120 ( .A1(n1295), .A2(n1068), .A3(G217), .ZN(n1389) );
INV_X1 U1121 ( .A(G953), .ZN(n1068) );
XNOR2_X1 U1122 ( .A(G234), .B(KEYINPUT27), .ZN(n1295) );
NAND2_X1 U1123 ( .A1(KEYINPUT48), .A2(n1361), .ZN(n1285) );
INV_X1 U1124 ( .A(G110), .ZN(n1361) );
endmodule


