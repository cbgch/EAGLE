//Key = 1010011100001000001000100010010111001110000011110011011010001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409;

XOR2_X1 U776 ( .A(G107), .B(n1070), .Z(G9) );
NOR2_X1 U777 ( .A1(n1071), .A2(n1072), .ZN(G75) );
NOR3_X1 U778 ( .A1(n1073), .A2(G953), .A3(G952), .ZN(n1072) );
NOR4_X1 U779 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1073), .ZN(n1071) );
AND4_X1 U780 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1073) );
NOR4_X1 U781 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1080) );
XNOR2_X1 U782 ( .A(G472), .B(n1085), .ZN(n1084) );
XOR2_X1 U783 ( .A(n1086), .B(n1087), .Z(n1083) );
NAND2_X1 U784 ( .A1(n1088), .A2(KEYINPUT18), .ZN(n1087) );
XNOR2_X1 U785 ( .A(n1089), .B(KEYINPUT22), .ZN(n1088) );
NOR2_X1 U786 ( .A1(n1090), .A2(n1091), .ZN(n1079) );
XNOR2_X1 U787 ( .A(n1092), .B(n1093), .ZN(n1078) );
NOR2_X1 U788 ( .A1(n1094), .A2(KEYINPUT20), .ZN(n1093) );
XOR2_X1 U789 ( .A(n1095), .B(n1096), .Z(n1077) );
XNOR2_X1 U790 ( .A(G475), .B(KEYINPUT44), .ZN(n1096) );
NOR3_X1 U791 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1076) );
NOR2_X1 U792 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NOR2_X1 U793 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR3_X1 U796 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1106) );
AND2_X1 U797 ( .A1(n1111), .A2(KEYINPUT23), .ZN(n1110) );
NOR3_X1 U798 ( .A1(KEYINPUT23), .A2(n1112), .A3(n1111), .ZN(n1109) );
NOR2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1104) );
NOR2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR3_X1 U801 ( .A1(n1107), .A2(n1114), .A3(n1117), .ZN(n1100) );
NAND3_X1 U802 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1075) );
NAND2_X1 U803 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND3_X1 U805 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
INV_X1 U806 ( .A(KEYINPUT13), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(n1123) );
NAND2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U809 ( .A1(KEYINPUT62), .A2(n1132), .ZN(n1131) );
NAND2_X1 U810 ( .A1(n1090), .A2(n1133), .ZN(n1130) );
INV_X1 U811 ( .A(n1134), .ZN(n1090) );
NAND3_X1 U812 ( .A1(n1135), .A2(n1136), .A3(KEYINPUT13), .ZN(n1118) );
NAND4_X1 U813 ( .A1(n1127), .A2(n1137), .A3(n1125), .A4(n1138), .ZN(n1136) );
INV_X1 U814 ( .A(n1097), .ZN(n1137) );
XNOR2_X1 U815 ( .A(n1139), .B(KEYINPUT54), .ZN(n1127) );
NAND4_X1 U816 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1074) );
NAND2_X1 U817 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND3_X1 U818 ( .A1(n1128), .A2(n1132), .A3(n1121), .ZN(n1145) );
NOR3_X1 U819 ( .A1(n1107), .A2(n1114), .A3(n1097), .ZN(n1121) );
INV_X1 U820 ( .A(n1135), .ZN(n1114) );
INV_X1 U821 ( .A(KEYINPUT62), .ZN(n1144) );
NAND2_X1 U822 ( .A1(n1146), .A2(n1147), .ZN(G72) );
NAND2_X1 U823 ( .A1(G953), .A2(n1148), .ZN(n1147) );
NAND2_X1 U824 ( .A1(G900), .A2(n1149), .ZN(n1148) );
OR2_X1 U825 ( .A1(n1150), .A2(G227), .ZN(n1149) );
XOR2_X1 U826 ( .A(n1151), .B(KEYINPUT58), .Z(n1146) );
NAND2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U828 ( .A1(G953), .A2(n1154), .ZN(n1153) );
XNOR2_X1 U829 ( .A(n1140), .B(n1150), .ZN(n1152) );
XNOR2_X1 U830 ( .A(n1155), .B(n1156), .ZN(n1150) );
XNOR2_X1 U831 ( .A(G140), .B(n1157), .ZN(n1156) );
NAND2_X1 U832 ( .A1(KEYINPUT29), .A2(n1158), .ZN(n1157) );
XOR2_X1 U833 ( .A(n1159), .B(n1160), .Z(n1155) );
NAND2_X1 U834 ( .A1(n1161), .A2(n1162), .ZN(G69) );
NAND3_X1 U835 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
OR2_X1 U836 ( .A1(n1119), .A2(G224), .ZN(n1165) );
NAND2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
NAND4_X1 U838 ( .A1(n1166), .A2(G953), .A3(n1168), .A4(n1167), .ZN(n1161) );
INV_X1 U839 ( .A(KEYINPUT19), .ZN(n1167) );
NAND2_X1 U840 ( .A1(G898), .A2(G224), .ZN(n1168) );
XOR2_X1 U841 ( .A(n1169), .B(n1170), .Z(n1166) );
AND2_X1 U842 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND2_X1 U843 ( .A1(n1141), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U844 ( .A(n1142), .B(KEYINPUT47), .ZN(n1173) );
XNOR2_X1 U845 ( .A(KEYINPUT6), .B(n1119), .ZN(n1171) );
NAND3_X1 U846 ( .A1(n1174), .A2(n1175), .A3(n1164), .ZN(n1169) );
INV_X1 U847 ( .A(n1176), .ZN(n1164) );
NAND2_X1 U848 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
INV_X1 U849 ( .A(n1179), .ZN(n1178) );
NAND2_X1 U850 ( .A1(n1180), .A2(n1179), .ZN(n1174) );
XNOR2_X1 U851 ( .A(n1177), .B(KEYINPUT24), .ZN(n1180) );
XOR2_X1 U852 ( .A(n1181), .B(n1182), .Z(n1177) );
NOR2_X1 U853 ( .A1(KEYINPUT40), .A2(n1183), .ZN(n1182) );
NOR2_X1 U854 ( .A1(n1184), .A2(n1185), .ZN(G66) );
XNOR2_X1 U855 ( .A(n1186), .B(n1187), .ZN(n1185) );
NOR3_X1 U856 ( .A1(n1188), .A2(KEYINPUT1), .A3(n1189), .ZN(n1187) );
NOR2_X1 U857 ( .A1(n1184), .A2(n1190), .ZN(G63) );
XNOR2_X1 U858 ( .A(n1191), .B(n1192), .ZN(n1190) );
AND2_X1 U859 ( .A1(G478), .A2(n1193), .ZN(n1192) );
NOR2_X1 U860 ( .A1(n1184), .A2(n1194), .ZN(G60) );
XNOR2_X1 U861 ( .A(n1195), .B(n1196), .ZN(n1194) );
NOR3_X1 U862 ( .A1(n1188), .A2(KEYINPUT42), .A3(n1197), .ZN(n1195) );
XOR2_X1 U863 ( .A(G104), .B(n1198), .Z(G6) );
NOR3_X1 U864 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(G57) );
AND2_X1 U865 ( .A1(KEYINPUT50), .A2(n1184), .ZN(n1201) );
NOR3_X1 U866 ( .A1(KEYINPUT50), .A2(G953), .A3(G952), .ZN(n1200) );
NOR2_X1 U867 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
XOR2_X1 U868 ( .A(KEYINPUT30), .B(n1204), .Z(n1203) );
NOR2_X1 U869 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U870 ( .A(n1207), .B(n1208), .Z(n1206) );
INV_X1 U871 ( .A(n1209), .ZN(n1205) );
NOR2_X1 U872 ( .A1(n1210), .A2(n1209), .ZN(n1202) );
XNOR2_X1 U873 ( .A(n1207), .B(n1208), .ZN(n1210) );
XNOR2_X1 U874 ( .A(n1211), .B(KEYINPUT48), .ZN(n1208) );
NAND2_X1 U875 ( .A1(n1193), .A2(G472), .ZN(n1211) );
NOR2_X1 U876 ( .A1(n1184), .A2(n1212), .ZN(G54) );
XOR2_X1 U877 ( .A(n1213), .B(n1214), .Z(n1212) );
XNOR2_X1 U878 ( .A(n1215), .B(n1216), .ZN(n1214) );
NAND2_X1 U879 ( .A1(KEYINPUT0), .A2(n1217), .ZN(n1215) );
XOR2_X1 U880 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U881 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U882 ( .A(n1222), .B(n1223), .Z(n1213) );
NOR2_X1 U883 ( .A1(KEYINPUT28), .A2(n1224), .ZN(n1223) );
AND2_X1 U884 ( .A1(G469), .A2(n1193), .ZN(n1222) );
INV_X1 U885 ( .A(n1188), .ZN(n1193) );
NOR2_X1 U886 ( .A1(n1184), .A2(n1225), .ZN(G51) );
XOR2_X1 U887 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U888 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
XOR2_X1 U889 ( .A(n1230), .B(KEYINPUT12), .Z(n1229) );
NAND2_X1 U890 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NOR2_X1 U891 ( .A1(n1231), .A2(n1232), .ZN(n1228) );
XOR2_X1 U892 ( .A(n1233), .B(n1234), .Z(n1231) );
XOR2_X1 U893 ( .A(n1235), .B(n1236), .Z(n1234) );
XNOR2_X1 U894 ( .A(G125), .B(KEYINPUT45), .ZN(n1233) );
NOR2_X1 U895 ( .A1(n1092), .A2(n1188), .ZN(n1226) );
NAND2_X1 U896 ( .A1(G902), .A2(n1237), .ZN(n1188) );
NAND3_X1 U897 ( .A1(n1142), .A2(n1141), .A3(n1140), .ZN(n1237) );
AND4_X1 U898 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1140) );
NOR4_X1 U899 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1241) );
NOR2_X1 U900 ( .A1(n1246), .A2(n1247), .ZN(n1240) );
INV_X1 U901 ( .A(n1248), .ZN(n1246) );
NAND3_X1 U902 ( .A1(n1249), .A2(n1115), .A3(n1250), .ZN(n1238) );
AND2_X1 U903 ( .A1(n1251), .A2(n1252), .ZN(n1141) );
NOR4_X1 U904 ( .A1(n1070), .A2(n1253), .A3(n1254), .A4(n1198), .ZN(n1252) );
AND3_X1 U905 ( .A1(n1255), .A2(n1128), .A3(n1116), .ZN(n1198) );
INV_X1 U906 ( .A(n1256), .ZN(n1254) );
INV_X1 U907 ( .A(n1257), .ZN(n1253) );
AND3_X1 U908 ( .A1(n1128), .A2(n1115), .A3(n1255), .ZN(n1070) );
NOR4_X1 U909 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1251) );
NOR2_X1 U910 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
INV_X1 U911 ( .A(KEYINPUT38), .ZN(n1263) );
AND2_X1 U912 ( .A1(n1264), .A2(KEYINPUT60), .ZN(n1260) );
NOR3_X1 U913 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1259) );
NOR2_X1 U914 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
INV_X1 U915 ( .A(KEYINPUT55), .ZN(n1269) );
NOR3_X1 U916 ( .A1(n1099), .A2(n1270), .A3(n1108), .ZN(n1268) );
NOR2_X1 U917 ( .A1(KEYINPUT55), .A2(n1271), .ZN(n1266) );
NOR4_X1 U918 ( .A1(n1272), .A2(n1273), .A3(n1107), .A4(n1274), .ZN(n1258) );
INV_X1 U919 ( .A(n1138), .ZN(n1107) );
NOR2_X1 U920 ( .A1(n1275), .A2(n1276), .ZN(n1272) );
NOR2_X1 U921 ( .A1(KEYINPUT38), .A2(n1277), .ZN(n1276) );
NOR2_X1 U922 ( .A1(KEYINPUT60), .A2(n1117), .ZN(n1275) );
INV_X1 U923 ( .A(n1249), .ZN(n1117) );
AND2_X1 U924 ( .A1(n1278), .A2(n1279), .ZN(n1142) );
NAND4_X1 U925 ( .A1(n1128), .A2(n1280), .A3(n1271), .A4(n1281), .ZN(n1279) );
INV_X1 U926 ( .A(KEYINPUT32), .ZN(n1281) );
NAND2_X1 U927 ( .A1(n1282), .A2(n1081), .ZN(n1280) );
NAND2_X1 U928 ( .A1(n1283), .A2(KEYINPUT32), .ZN(n1278) );
NOR2_X1 U929 ( .A1(n1119), .A2(G952), .ZN(n1184) );
XOR2_X1 U930 ( .A(G146), .B(n1245), .Z(G48) );
AND2_X1 U931 ( .A1(n1284), .A2(n1116), .ZN(n1245) );
XNOR2_X1 U932 ( .A(G143), .B(n1239), .ZN(G45) );
NAND4_X1 U933 ( .A1(n1282), .A2(n1285), .A3(n1108), .A4(n1081), .ZN(n1239) );
XOR2_X1 U934 ( .A(G140), .B(n1244), .Z(G42) );
AND3_X1 U935 ( .A1(n1250), .A2(n1116), .A3(n1125), .ZN(n1244) );
XOR2_X1 U936 ( .A(G137), .B(n1243), .Z(G39) );
NOR2_X1 U937 ( .A1(n1265), .A2(n1286), .ZN(n1243) );
XNOR2_X1 U938 ( .A(G134), .B(n1287), .ZN(G36) );
NAND3_X1 U939 ( .A1(n1285), .A2(n1115), .A3(n1288), .ZN(n1287) );
XNOR2_X1 U940 ( .A(n1135), .B(KEYINPUT56), .ZN(n1288) );
AND3_X1 U941 ( .A1(n1132), .A2(n1289), .A3(n1249), .ZN(n1285) );
XOR2_X1 U942 ( .A(n1242), .B(n1290), .Z(G33) );
NOR2_X1 U943 ( .A1(KEYINPUT41), .A2(n1291), .ZN(n1290) );
AND3_X1 U944 ( .A1(n1116), .A2(n1249), .A3(n1250), .ZN(n1242) );
INV_X1 U945 ( .A(n1286), .ZN(n1250) );
NAND3_X1 U946 ( .A1(n1132), .A2(n1289), .A3(n1135), .ZN(n1286) );
NOR2_X1 U947 ( .A1(n1112), .A2(n1091), .ZN(n1135) );
XNOR2_X1 U948 ( .A(n1292), .B(n1247), .ZN(G30) );
AND2_X1 U949 ( .A1(n1284), .A2(n1115), .ZN(n1247) );
AND4_X1 U950 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1289), .ZN(n1284) );
INV_X1 U951 ( .A(n1273), .ZN(n1293) );
XNOR2_X1 U952 ( .A(n1296), .B(n1264), .ZN(G3) );
AND3_X1 U953 ( .A1(n1249), .A2(n1255), .A3(n1138), .ZN(n1264) );
XNOR2_X1 U954 ( .A(G125), .B(n1248), .ZN(G27) );
NAND4_X1 U955 ( .A1(n1139), .A2(n1125), .A3(n1297), .A4(n1116), .ZN(n1248) );
AND2_X1 U956 ( .A1(n1289), .A2(n1108), .ZN(n1297) );
NAND2_X1 U957 ( .A1(n1298), .A2(n1097), .ZN(n1289) );
NAND4_X1 U958 ( .A1(G953), .A2(G902), .A3(n1299), .A4(n1300), .ZN(n1298) );
INV_X1 U959 ( .A(G900), .ZN(n1300) );
XNOR2_X1 U960 ( .A(n1283), .B(n1301), .ZN(G24) );
NAND2_X1 U961 ( .A1(KEYINPUT31), .A2(G122), .ZN(n1301) );
NOR4_X1 U962 ( .A1(n1302), .A2(n1303), .A3(n1103), .A4(n1304), .ZN(n1283) );
INV_X1 U963 ( .A(n1128), .ZN(n1103) );
NOR2_X1 U964 ( .A1(n1295), .A2(n1294), .ZN(n1128) );
XOR2_X1 U965 ( .A(G119), .B(n1305), .Z(G21) );
NOR2_X1 U966 ( .A1(n1265), .A2(n1303), .ZN(n1305) );
NAND3_X1 U967 ( .A1(n1294), .A2(n1295), .A3(n1138), .ZN(n1265) );
XNOR2_X1 U968 ( .A(G116), .B(n1256), .ZN(G18) );
NAND3_X1 U969 ( .A1(n1249), .A2(n1115), .A3(n1271), .ZN(n1256) );
NOR2_X1 U970 ( .A1(n1304), .A2(n1282), .ZN(n1115) );
INV_X1 U971 ( .A(n1081), .ZN(n1304) );
XNOR2_X1 U972 ( .A(G113), .B(n1257), .ZN(G15) );
NAND3_X1 U973 ( .A1(n1116), .A2(n1249), .A3(n1271), .ZN(n1257) );
INV_X1 U974 ( .A(n1303), .ZN(n1271) );
NAND3_X1 U975 ( .A1(n1108), .A2(n1274), .A3(n1139), .ZN(n1303) );
INV_X1 U976 ( .A(n1099), .ZN(n1139) );
NAND2_X1 U977 ( .A1(n1306), .A2(n1134), .ZN(n1099) );
XNOR2_X1 U978 ( .A(n1082), .B(KEYINPUT15), .ZN(n1306) );
NOR2_X1 U979 ( .A1(n1294), .A2(n1307), .ZN(n1249) );
NOR2_X1 U980 ( .A1(n1302), .A2(n1081), .ZN(n1116) );
XNOR2_X1 U981 ( .A(G110), .B(n1262), .ZN(G12) );
NAND3_X1 U982 ( .A1(n1138), .A2(n1255), .A3(n1125), .ZN(n1262) );
INV_X1 U983 ( .A(n1277), .ZN(n1125) );
NAND2_X1 U984 ( .A1(n1307), .A2(n1294), .ZN(n1277) );
NAND3_X1 U985 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1294) );
NAND2_X1 U986 ( .A1(n1089), .A2(n1086), .ZN(n1310) );
NAND2_X1 U987 ( .A1(KEYINPUT10), .A2(n1311), .ZN(n1309) );
NAND2_X1 U988 ( .A1(n1312), .A2(n1189), .ZN(n1311) );
XNOR2_X1 U989 ( .A(n1086), .B(n1313), .ZN(n1312) );
NAND2_X1 U990 ( .A1(n1314), .A2(n1315), .ZN(n1308) );
INV_X1 U991 ( .A(KEYINPUT10), .ZN(n1315) );
NAND2_X1 U992 ( .A1(n1316), .A2(n1317), .ZN(n1314) );
NAND2_X1 U993 ( .A1(n1086), .A2(n1313), .ZN(n1317) );
OR3_X1 U994 ( .A1(n1086), .A2(n1089), .A3(n1313), .ZN(n1316) );
INV_X1 U995 ( .A(KEYINPUT33), .ZN(n1313) );
INV_X1 U996 ( .A(n1189), .ZN(n1089) );
NAND2_X1 U997 ( .A1(G217), .A2(n1318), .ZN(n1189) );
NAND2_X1 U998 ( .A1(n1319), .A2(n1186), .ZN(n1086) );
XNOR2_X1 U999 ( .A(n1320), .B(n1321), .ZN(n1186) );
XNOR2_X1 U1000 ( .A(n1322), .B(n1323), .ZN(n1321) );
NOR2_X1 U1001 ( .A1(KEYINPUT8), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1002 ( .A(n1325), .B(n1326), .Z(n1324) );
XNOR2_X1 U1003 ( .A(G140), .B(n1158), .ZN(n1326) );
NOR2_X1 U1004 ( .A1(KEYINPUT61), .A2(n1327), .ZN(n1325) );
NAND2_X1 U1005 ( .A1(KEYINPUT37), .A2(n1328), .ZN(n1322) );
XOR2_X1 U1006 ( .A(G137), .B(n1329), .Z(n1328) );
AND4_X1 U1007 ( .A1(n1330), .A2(G234), .A3(G221), .A4(n1331), .ZN(n1329) );
INV_X1 U1008 ( .A(KEYINPUT39), .ZN(n1330) );
XNOR2_X1 U1009 ( .A(G110), .B(n1332), .ZN(n1320) );
XNOR2_X1 U1010 ( .A(n1292), .B(G119), .ZN(n1332) );
INV_X1 U1011 ( .A(n1295), .ZN(n1307) );
NAND2_X1 U1012 ( .A1(n1333), .A2(n1334), .ZN(n1295) );
NAND2_X1 U1013 ( .A1(G472), .A2(n1085), .ZN(n1334) );
XOR2_X1 U1014 ( .A(KEYINPUT5), .B(n1335), .Z(n1333) );
NOR2_X1 U1015 ( .A1(G472), .A2(n1085), .ZN(n1335) );
NAND2_X1 U1016 ( .A1(n1319), .A2(n1336), .ZN(n1085) );
XNOR2_X1 U1017 ( .A(n1337), .B(n1209), .ZN(n1336) );
NAND2_X1 U1018 ( .A1(n1338), .A2(n1339), .ZN(n1209) );
NAND2_X1 U1019 ( .A1(n1340), .A2(n1296), .ZN(n1339) );
NAND2_X1 U1020 ( .A1(n1341), .A2(G210), .ZN(n1340) );
NAND3_X1 U1021 ( .A1(n1341), .A2(G210), .A3(G101), .ZN(n1338) );
XNOR2_X1 U1022 ( .A(n1207), .B(KEYINPUT59), .ZN(n1337) );
XNOR2_X1 U1023 ( .A(n1342), .B(n1343), .ZN(n1207) );
XOR2_X1 U1024 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1025 ( .A(G119), .B(n1346), .ZN(n1345) );
NOR2_X1 U1026 ( .A1(KEYINPUT57), .A2(n1347), .ZN(n1346) );
INV_X1 U1027 ( .A(G113), .ZN(n1347) );
NAND2_X1 U1028 ( .A1(KEYINPUT7), .A2(n1348), .ZN(n1344) );
XOR2_X1 U1029 ( .A(n1236), .B(n1160), .Z(n1342) );
NOR2_X1 U1030 ( .A1(n1273), .A2(n1270), .ZN(n1255) );
INV_X1 U1031 ( .A(n1274), .ZN(n1270) );
NAND2_X1 U1032 ( .A1(n1097), .A2(n1349), .ZN(n1274) );
NAND3_X1 U1033 ( .A1(G902), .A2(n1299), .A3(n1176), .ZN(n1349) );
NOR2_X1 U1034 ( .A1(n1119), .A2(G898), .ZN(n1176) );
NAND3_X1 U1035 ( .A1(n1299), .A2(n1119), .A3(G952), .ZN(n1097) );
INV_X1 U1036 ( .A(G953), .ZN(n1119) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1299) );
NAND2_X1 U1038 ( .A1(n1132), .A2(n1108), .ZN(n1273) );
NOR2_X1 U1039 ( .A1(n1350), .A2(n1091), .ZN(n1108) );
INV_X1 U1040 ( .A(n1111), .ZN(n1091) );
NAND2_X1 U1041 ( .A1(G214), .A2(n1351), .ZN(n1111) );
INV_X1 U1042 ( .A(n1112), .ZN(n1350) );
XNOR2_X1 U1043 ( .A(n1094), .B(n1092), .ZN(n1112) );
NAND2_X1 U1044 ( .A1(G210), .A2(n1351), .ZN(n1092) );
NAND2_X1 U1045 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
INV_X1 U1046 ( .A(G237), .ZN(n1352) );
AND2_X1 U1047 ( .A1(n1319), .A2(n1354), .ZN(n1094) );
XOR2_X1 U1048 ( .A(n1355), .B(n1356), .Z(n1354) );
XNOR2_X1 U1049 ( .A(n1236), .B(n1232), .ZN(n1356) );
XNOR2_X1 U1050 ( .A(n1179), .B(n1357), .ZN(n1232) );
NOR2_X1 U1051 ( .A1(KEYINPUT25), .A2(n1358), .ZN(n1357) );
XNOR2_X1 U1052 ( .A(n1183), .B(n1359), .ZN(n1358) );
INV_X1 U1053 ( .A(n1181), .ZN(n1359) );
XNOR2_X1 U1054 ( .A(n1360), .B(n1361), .ZN(n1181) );
XNOR2_X1 U1055 ( .A(n1348), .B(n1362), .ZN(n1361) );
NOR2_X1 U1056 ( .A1(G113), .A2(KEYINPUT4), .ZN(n1362) );
XNOR2_X1 U1057 ( .A(G119), .B(KEYINPUT52), .ZN(n1360) );
NAND2_X1 U1058 ( .A1(n1363), .A2(n1364), .ZN(n1183) );
NAND2_X1 U1059 ( .A1(n1365), .A2(n1296), .ZN(n1364) );
XOR2_X1 U1060 ( .A(KEYINPUT46), .B(n1366), .Z(n1363) );
NOR2_X1 U1061 ( .A1(n1365), .A2(n1296), .ZN(n1366) );
INV_X1 U1062 ( .A(G101), .ZN(n1296) );
XNOR2_X1 U1063 ( .A(G104), .B(n1367), .ZN(n1365) );
XOR2_X1 U1064 ( .A(KEYINPUT43), .B(G107), .Z(n1367) );
NAND4_X1 U1065 ( .A1(n1368), .A2(n1369), .A3(n1370), .A4(n1371), .ZN(n1179) );
OR3_X1 U1066 ( .A1(n1372), .A2(G110), .A3(KEYINPUT51), .ZN(n1371) );
AND2_X1 U1067 ( .A1(KEYINPUT11), .A2(n1373), .ZN(n1372) );
NAND3_X1 U1068 ( .A1(G110), .A2(n1374), .A3(KEYINPUT51), .ZN(n1370) );
OR2_X1 U1069 ( .A1(G122), .A2(KEYINPUT11), .ZN(n1374) );
NAND3_X1 U1070 ( .A1(n1375), .A2(n1373), .A3(n1376), .ZN(n1369) );
INV_X1 U1071 ( .A(KEYINPUT34), .ZN(n1376) );
XNOR2_X1 U1072 ( .A(KEYINPUT11), .B(G110), .ZN(n1375) );
NAND2_X1 U1073 ( .A1(KEYINPUT34), .A2(G122), .ZN(n1368) );
XNOR2_X1 U1074 ( .A(n1220), .B(n1377), .ZN(n1236) );
NOR2_X1 U1075 ( .A1(KEYINPUT14), .A2(n1292), .ZN(n1377) );
XNOR2_X1 U1076 ( .A(n1235), .B(n1378), .ZN(n1355) );
NOR2_X1 U1077 ( .A1(G125), .A2(KEYINPUT16), .ZN(n1378) );
NAND2_X1 U1078 ( .A1(G224), .A2(n1331), .ZN(n1235) );
AND2_X1 U1079 ( .A1(n1379), .A2(n1134), .ZN(n1132) );
NAND2_X1 U1080 ( .A1(G221), .A2(n1318), .ZN(n1134) );
NAND2_X1 U1081 ( .A1(G234), .A2(n1353), .ZN(n1318) );
INV_X1 U1082 ( .A(G902), .ZN(n1353) );
XNOR2_X1 U1083 ( .A(KEYINPUT35), .B(n1133), .ZN(n1379) );
INV_X1 U1084 ( .A(n1082), .ZN(n1133) );
XNOR2_X1 U1085 ( .A(n1380), .B(G469), .ZN(n1082) );
NAND2_X1 U1086 ( .A1(n1319), .A2(n1381), .ZN(n1380) );
XOR2_X1 U1087 ( .A(n1382), .B(n1383), .Z(n1381) );
XOR2_X1 U1088 ( .A(n1218), .B(n1224), .Z(n1383) );
XNOR2_X1 U1089 ( .A(n1384), .B(n1385), .ZN(n1224) );
NOR2_X1 U1090 ( .A1(n1386), .A2(n1154), .ZN(n1385) );
INV_X1 U1091 ( .A(G227), .ZN(n1154) );
XNOR2_X1 U1092 ( .A(G140), .B(G110), .ZN(n1384) );
XOR2_X1 U1093 ( .A(G101), .B(n1387), .Z(n1218) );
NOR2_X1 U1094 ( .A1(G104), .A2(n1388), .ZN(n1387) );
XNOR2_X1 U1095 ( .A(KEYINPUT3), .B(KEYINPUT26), .ZN(n1388) );
XNOR2_X1 U1096 ( .A(n1389), .B(n1390), .ZN(n1382) );
XOR2_X1 U1097 ( .A(G107), .B(n1391), .Z(n1390) );
NOR2_X1 U1098 ( .A1(KEYINPUT21), .A2(n1159), .ZN(n1391) );
XNOR2_X1 U1099 ( .A(G128), .B(n1220), .ZN(n1159) );
INV_X1 U1100 ( .A(n1216), .ZN(n1389) );
XOR2_X1 U1101 ( .A(n1160), .B(KEYINPUT63), .Z(n1216) );
XOR2_X1 U1102 ( .A(G131), .B(n1392), .Z(n1160) );
XOR2_X1 U1103 ( .A(G137), .B(G134), .Z(n1392) );
NOR2_X1 U1104 ( .A1(n1081), .A2(n1282), .ZN(n1138) );
INV_X1 U1105 ( .A(n1302), .ZN(n1282) );
XOR2_X1 U1106 ( .A(n1393), .B(n1095), .Z(n1302) );
NAND2_X1 U1107 ( .A1(n1196), .A2(n1319), .ZN(n1095) );
XOR2_X1 U1108 ( .A(n1394), .B(n1395), .Z(n1196) );
XOR2_X1 U1109 ( .A(n1396), .B(n1397), .Z(n1395) );
XNOR2_X1 U1110 ( .A(n1373), .B(G113), .ZN(n1397) );
INV_X1 U1111 ( .A(G122), .ZN(n1373) );
XNOR2_X1 U1112 ( .A(G140), .B(n1291), .ZN(n1396) );
INV_X1 U1113 ( .A(G131), .ZN(n1291) );
XOR2_X1 U1114 ( .A(n1398), .B(n1399), .Z(n1394) );
XNOR2_X1 U1115 ( .A(G104), .B(n1400), .ZN(n1399) );
NAND2_X1 U1116 ( .A1(n1341), .A2(G214), .ZN(n1400) );
NOR2_X1 U1117 ( .A1(n1386), .A2(G237), .ZN(n1341) );
XOR2_X1 U1118 ( .A(n1401), .B(n1220), .Z(n1398) );
XOR2_X1 U1119 ( .A(G143), .B(n1327), .Z(n1220) );
XOR2_X1 U1120 ( .A(G146), .B(KEYINPUT49), .Z(n1327) );
NAND2_X1 U1121 ( .A1(KEYINPUT2), .A2(n1158), .ZN(n1401) );
INV_X1 U1122 ( .A(G125), .ZN(n1158) );
NAND2_X1 U1123 ( .A1(KEYINPUT53), .A2(n1197), .ZN(n1393) );
INV_X1 U1124 ( .A(G475), .ZN(n1197) );
XNOR2_X1 U1125 ( .A(n1402), .B(G478), .ZN(n1081) );
NAND2_X1 U1126 ( .A1(n1319), .A2(n1191), .ZN(n1402) );
XNOR2_X1 U1127 ( .A(n1403), .B(n1404), .ZN(n1191) );
XNOR2_X1 U1128 ( .A(n1221), .B(n1405), .ZN(n1404) );
XOR2_X1 U1129 ( .A(n1406), .B(n1407), .Z(n1405) );
AND3_X1 U1130 ( .A1(G217), .A2(G234), .A3(n1331), .ZN(n1407) );
INV_X1 U1131 ( .A(n1386), .ZN(n1331) );
XOR2_X1 U1132 ( .A(G953), .B(KEYINPUT17), .Z(n1386) );
NAND2_X1 U1133 ( .A1(KEYINPUT36), .A2(n1348), .ZN(n1406) );
INV_X1 U1134 ( .A(G116), .ZN(n1348) );
XNOR2_X1 U1135 ( .A(G107), .B(n1292), .ZN(n1221) );
INV_X1 U1136 ( .A(G128), .ZN(n1292) );
XOR2_X1 U1137 ( .A(n1408), .B(n1409), .Z(n1403) );
NOR2_X1 U1138 ( .A1(KEYINPUT9), .A2(G143), .ZN(n1409) );
XNOR2_X1 U1139 ( .A(G134), .B(G122), .ZN(n1408) );
XNOR2_X1 U1140 ( .A(G902), .B(KEYINPUT27), .ZN(n1319) );
endmodule


