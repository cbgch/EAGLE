//Key = 0111111100111101010100100010100001110010111110101111111000000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
n1428, n1429, n1430, n1431;

XNOR2_X1 U787 ( .A(G107), .B(n1088), .ZN(G9) );
NOR2_X1 U788 ( .A1(n1089), .A2(n1090), .ZN(G75) );
NOR4_X1 U789 ( .A1(G953), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1090) );
INV_X1 U790 ( .A(n1094), .ZN(n1093) );
NOR2_X1 U791 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NOR2_X1 U792 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR3_X1 U793 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NOR2_X1 U794 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U796 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U797 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NOR2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1106) );
NOR2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NOR3_X1 U803 ( .A1(n1115), .A2(n1120), .A3(n1109), .ZN(n1102) );
NOR2_X1 U804 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U805 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NOR4_X1 U806 ( .A1(n1125), .A2(n1109), .A3(n1105), .A4(n1115), .ZN(n1097) );
INV_X1 U807 ( .A(n1126), .ZN(n1105) );
NOR2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
INV_X1 U809 ( .A(n1129), .ZN(n1095) );
NOR3_X1 U810 ( .A1(n1091), .A2(G953), .A3(G952), .ZN(n1089) );
AND4_X1 U811 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1091) );
NOR4_X1 U812 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(n1136) );
NAND2_X1 U815 ( .A1(n1124), .A2(n1113), .ZN(n1135) );
NOR3_X1 U816 ( .A1(n1142), .A2(n1143), .A3(n1099), .ZN(n1132) );
XOR2_X1 U817 ( .A(n1144), .B(KEYINPUT63), .Z(n1143) );
NAND2_X1 U818 ( .A1(n1138), .A2(n1139), .ZN(n1144) );
XNOR2_X1 U819 ( .A(n1145), .B(G469), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1130) );
XNOR2_X1 U821 ( .A(KEYINPUT11), .B(n1148), .ZN(n1147) );
NAND2_X1 U822 ( .A1(KEYINPUT10), .A2(n1149), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1150), .B(n1151), .Z(G72) );
XOR2_X1 U824 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U825 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U826 ( .A(n1156), .B(n1157), .Z(n1155) );
XNOR2_X1 U827 ( .A(n1158), .B(n1159), .ZN(n1157) );
XNOR2_X1 U828 ( .A(n1160), .B(n1161), .ZN(n1156) );
NAND2_X1 U829 ( .A1(KEYINPUT40), .A2(n1162), .ZN(n1160) );
NOR2_X1 U830 ( .A1(G900), .A2(n1163), .ZN(n1154) );
NOR3_X1 U831 ( .A1(n1164), .A2(KEYINPUT29), .A3(G953), .ZN(n1152) );
XOR2_X1 U832 ( .A(KEYINPUT0), .B(n1165), .Z(n1164) );
NOR2_X1 U833 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR2_X1 U834 ( .A1(n1168), .A2(n1163), .ZN(n1150) );
AND2_X1 U835 ( .A1(G227), .A2(G900), .ZN(n1168) );
XOR2_X1 U836 ( .A(n1169), .B(n1170), .Z(G69) );
XOR2_X1 U837 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U838 ( .A1(n1173), .A2(n1163), .ZN(n1172) );
AND2_X1 U839 ( .A1(G224), .A2(G898), .ZN(n1173) );
NOR2_X1 U840 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
XNOR2_X1 U841 ( .A(G953), .B(KEYINPUT6), .ZN(n1175) );
NOR2_X1 U842 ( .A1(n1176), .A2(n1177), .ZN(n1174) );
XOR2_X1 U843 ( .A(KEYINPUT31), .B(n1178), .Z(n1177) );
NOR3_X1 U844 ( .A1(n1179), .A2(KEYINPUT8), .A3(n1180), .ZN(n1169) );
XOR2_X1 U845 ( .A(KEYINPUT20), .B(n1181), .Z(n1179) );
NOR2_X1 U846 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XNOR2_X1 U848 ( .A(n1186), .B(KEYINPUT33), .ZN(n1185) );
AND2_X1 U849 ( .A1(n1184), .A2(n1186), .ZN(n1182) );
XOR2_X1 U850 ( .A(n1187), .B(n1188), .Z(n1184) );
XOR2_X1 U851 ( .A(n1189), .B(KEYINPUT49), .Z(n1187) );
NOR2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(G66) );
NOR3_X1 U853 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1191) );
NOR3_X1 U854 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
NOR2_X1 U855 ( .A1(n1198), .A2(n1199), .ZN(n1193) );
NOR2_X1 U856 ( .A1(n1094), .A2(n1196), .ZN(n1198) );
NOR2_X1 U857 ( .A1(n1190), .A2(n1200), .ZN(G63) );
NOR3_X1 U858 ( .A1(n1138), .A2(n1201), .A3(n1202), .ZN(n1200) );
AND3_X1 U859 ( .A1(n1203), .A2(G478), .A3(n1204), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1205), .A2(n1203), .ZN(n1201) );
NOR2_X1 U861 ( .A1(n1094), .A2(n1139), .ZN(n1205) );
NOR2_X1 U862 ( .A1(n1190), .A2(n1206), .ZN(G60) );
NOR2_X1 U863 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U864 ( .A(KEYINPUT36), .B(n1209), .Z(n1208) );
NOR2_X1 U865 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
AND2_X1 U866 ( .A1(n1211), .A2(n1210), .ZN(n1207) );
NAND2_X1 U867 ( .A1(n1204), .A2(G475), .ZN(n1211) );
XOR2_X1 U868 ( .A(G104), .B(n1212), .Z(G6) );
NOR2_X1 U869 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NOR2_X1 U870 ( .A1(n1190), .A2(n1215), .ZN(G57) );
XNOR2_X1 U871 ( .A(n1216), .B(n1217), .ZN(n1215) );
NOR2_X1 U872 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U873 ( .A(KEYINPUT59), .B(n1220), .Z(n1219) );
NOR2_X1 U874 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
AND2_X1 U875 ( .A1(n1222), .A2(n1221), .ZN(n1218) );
NOR2_X1 U876 ( .A1(n1197), .A2(n1149), .ZN(n1221) );
XOR2_X1 U877 ( .A(n1223), .B(n1224), .Z(n1222) );
NAND2_X1 U878 ( .A1(KEYINPUT26), .A2(n1225), .ZN(n1223) );
NOR2_X1 U879 ( .A1(n1190), .A2(n1226), .ZN(G54) );
XOR2_X1 U880 ( .A(n1227), .B(n1228), .Z(n1226) );
XOR2_X1 U881 ( .A(n1229), .B(n1230), .Z(n1228) );
AND2_X1 U882 ( .A1(G469), .A2(n1204), .ZN(n1230) );
NAND2_X1 U883 ( .A1(KEYINPUT48), .A2(n1231), .ZN(n1229) );
XOR2_X1 U884 ( .A(n1232), .B(n1233), .Z(n1227) );
XOR2_X1 U885 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND3_X1 U886 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1235) );
OR2_X1 U887 ( .A1(n1239), .A2(KEYINPUT12), .ZN(n1238) );
NAND3_X1 U888 ( .A1(KEYINPUT12), .A2(n1239), .A3(G140), .ZN(n1237) );
NAND2_X1 U889 ( .A1(n1240), .A2(n1241), .ZN(n1236) );
NAND2_X1 U890 ( .A1(KEYINPUT12), .A2(n1242), .ZN(n1240) );
XNOR2_X1 U891 ( .A(KEYINPUT3), .B(n1239), .ZN(n1242) );
NAND2_X1 U892 ( .A1(n1243), .A2(n1244), .ZN(n1232) );
OR2_X1 U893 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U894 ( .A(n1247), .B(KEYINPUT47), .Z(n1243) );
NAND2_X1 U895 ( .A1(n1245), .A2(n1246), .ZN(n1247) );
NOR2_X1 U896 ( .A1(n1190), .A2(n1248), .ZN(G51) );
XOR2_X1 U897 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U898 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U899 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U900 ( .A1(KEYINPUT21), .A2(n1246), .ZN(n1254) );
NOR2_X1 U901 ( .A1(n1255), .A2(n1197), .ZN(n1253) );
INV_X1 U902 ( .A(n1204), .ZN(n1197) );
NOR2_X1 U903 ( .A1(n1256), .A2(n1094), .ZN(n1204) );
NOR4_X1 U904 ( .A1(n1176), .A2(n1167), .A3(n1257), .A4(n1178), .ZN(n1094) );
XNOR2_X1 U905 ( .A(KEYINPUT7), .B(n1166), .ZN(n1257) );
INV_X1 U906 ( .A(n1258), .ZN(n1166) );
NAND4_X1 U907 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1167) );
NOR4_X1 U908 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1262) );
INV_X1 U909 ( .A(n1267), .ZN(n1264) );
NOR3_X1 U910 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1263) );
XNOR2_X1 U911 ( .A(KEYINPUT53), .B(n1213), .ZN(n1268) );
NAND4_X1 U912 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1176) );
AND3_X1 U913 ( .A1(n1275), .A2(n1088), .A3(n1276), .ZN(n1274) );
NAND2_X1 U914 ( .A1(n1277), .A2(n1278), .ZN(n1088) );
NAND2_X1 U915 ( .A1(n1111), .A2(n1279), .ZN(n1273) );
NAND2_X1 U916 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U917 ( .A1(n1282), .A2(n1127), .ZN(n1281) );
XOR2_X1 U918 ( .A(n1214), .B(KEYINPUT58), .Z(n1280) );
NAND2_X1 U919 ( .A1(n1128), .A2(n1278), .ZN(n1214) );
NOR3_X1 U920 ( .A1(n1109), .A2(n1283), .A3(n1284), .ZN(n1278) );
NAND2_X1 U921 ( .A1(n1285), .A2(n1286), .ZN(n1271) );
XNOR2_X1 U922 ( .A(n1287), .B(KEYINPUT28), .ZN(n1285) );
XOR2_X1 U923 ( .A(n1288), .B(n1289), .Z(n1249) );
XNOR2_X1 U924 ( .A(KEYINPUT52), .B(n1290), .ZN(n1289) );
NOR2_X1 U925 ( .A1(n1163), .A2(G952), .ZN(n1190) );
XNOR2_X1 U926 ( .A(G146), .B(n1261), .ZN(G48) );
NAND3_X1 U927 ( .A1(n1128), .A2(n1111), .A3(n1291), .ZN(n1261) );
XOR2_X1 U928 ( .A(n1259), .B(n1292), .Z(G45) );
XOR2_X1 U929 ( .A(KEYINPUT4), .B(G143), .Z(n1292) );
NAND4_X1 U930 ( .A1(n1293), .A2(n1294), .A3(n1111), .A4(n1295), .ZN(n1259) );
XOR2_X1 U931 ( .A(n1260), .B(n1296), .Z(G42) );
NAND2_X1 U932 ( .A1(G140), .A2(n1297), .ZN(n1296) );
XOR2_X1 U933 ( .A(KEYINPUT42), .B(KEYINPUT32), .Z(n1297) );
NAND4_X1 U934 ( .A1(n1298), .A2(n1128), .A3(n1299), .A4(n1300), .ZN(n1260) );
XOR2_X1 U935 ( .A(G137), .B(n1266), .Z(G39) );
NOR4_X1 U936 ( .A1(n1115), .A2(n1270), .A3(n1099), .A4(n1101), .ZN(n1266) );
INV_X1 U937 ( .A(n1298), .ZN(n1115) );
NAND3_X1 U938 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(G36) );
NAND2_X1 U939 ( .A1(G134), .A2(n1304), .ZN(n1303) );
NAND2_X1 U940 ( .A1(KEYINPUT37), .A2(n1305), .ZN(n1302) );
NAND2_X1 U941 ( .A1(n1306), .A2(n1265), .ZN(n1305) );
INV_X1 U942 ( .A(n1304), .ZN(n1265) );
XNOR2_X1 U943 ( .A(KEYINPUT16), .B(G134), .ZN(n1306) );
NAND2_X1 U944 ( .A1(n1307), .A2(n1308), .ZN(n1301) );
INV_X1 U945 ( .A(KEYINPUT37), .ZN(n1308) );
NAND2_X1 U946 ( .A1(n1309), .A2(n1310), .ZN(n1307) );
OR3_X1 U947 ( .A1(n1304), .A2(G134), .A3(KEYINPUT16), .ZN(n1310) );
NAND3_X1 U948 ( .A1(n1294), .A2(n1127), .A3(n1298), .ZN(n1304) );
NAND2_X1 U949 ( .A1(KEYINPUT16), .A2(G134), .ZN(n1309) );
XNOR2_X1 U950 ( .A(G131), .B(n1267), .ZN(G33) );
NAND3_X1 U951 ( .A1(n1294), .A2(n1128), .A3(n1298), .ZN(n1267) );
NOR2_X1 U952 ( .A1(n1112), .A2(n1311), .ZN(n1298) );
INV_X1 U953 ( .A(n1113), .ZN(n1311) );
AND3_X1 U954 ( .A1(n1122), .A2(n1300), .A3(n1117), .ZN(n1294) );
XNOR2_X1 U955 ( .A(G128), .B(n1312), .ZN(G30) );
NAND2_X1 U956 ( .A1(n1291), .A2(n1277), .ZN(n1312) );
NOR2_X1 U957 ( .A1(n1269), .A2(n1213), .ZN(n1277) );
INV_X1 U958 ( .A(n1127), .ZN(n1269) );
INV_X1 U959 ( .A(n1270), .ZN(n1291) );
NAND3_X1 U960 ( .A1(n1122), .A2(n1300), .A3(n1287), .ZN(n1270) );
XNOR2_X1 U961 ( .A(G101), .B(n1272), .ZN(G3) );
NAND3_X1 U962 ( .A1(n1313), .A2(n1122), .A3(n1117), .ZN(n1272) );
INV_X1 U963 ( .A(n1284), .ZN(n1122) );
XNOR2_X1 U964 ( .A(G125), .B(n1258), .ZN(G27) );
NAND4_X1 U965 ( .A1(n1314), .A2(n1126), .A3(n1128), .A4(n1315), .ZN(n1258) );
AND3_X1 U966 ( .A1(n1111), .A2(n1316), .A3(n1300), .ZN(n1315) );
NAND2_X1 U967 ( .A1(n1317), .A2(n1318), .ZN(n1300) );
NAND4_X1 U968 ( .A1(n1319), .A2(G953), .A3(n1129), .A4(n1320), .ZN(n1318) );
INV_X1 U969 ( .A(G900), .ZN(n1320) );
XOR2_X1 U970 ( .A(n1321), .B(G122), .Z(G24) );
NAND2_X1 U971 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NAND2_X1 U972 ( .A1(n1178), .A2(n1324), .ZN(n1323) );
INV_X1 U973 ( .A(KEYINPUT45), .ZN(n1324) );
NOR2_X1 U974 ( .A1(n1325), .A2(n1213), .ZN(n1178) );
NAND3_X1 U975 ( .A1(n1111), .A2(n1325), .A3(KEYINPUT45), .ZN(n1322) );
NAND3_X1 U976 ( .A1(n1293), .A2(n1126), .A3(n1326), .ZN(n1325) );
NOR3_X1 U977 ( .A1(n1109), .A2(n1283), .A3(n1327), .ZN(n1326) );
NAND2_X1 U978 ( .A1(n1118), .A2(n1314), .ZN(n1109) );
INV_X1 U979 ( .A(n1328), .ZN(n1293) );
XNOR2_X1 U980 ( .A(G119), .B(n1329), .ZN(G21) );
NAND2_X1 U981 ( .A1(n1286), .A2(n1287), .ZN(n1329) );
NOR2_X1 U982 ( .A1(n1314), .A2(n1118), .ZN(n1287) );
AND2_X1 U983 ( .A1(n1313), .A2(n1126), .ZN(n1286) );
XNOR2_X1 U984 ( .A(G116), .B(n1330), .ZN(G18) );
NAND3_X1 U985 ( .A1(n1282), .A2(n1127), .A3(n1331), .ZN(n1330) );
XNOR2_X1 U986 ( .A(n1111), .B(KEYINPUT13), .ZN(n1331) );
NOR2_X1 U987 ( .A1(n1099), .A2(n1327), .ZN(n1127) );
INV_X1 U988 ( .A(n1295), .ZN(n1327) );
XNOR2_X1 U989 ( .A(n1101), .B(KEYINPUT50), .ZN(n1295) );
NAND2_X1 U990 ( .A1(n1332), .A2(n1333), .ZN(G15) );
NAND2_X1 U991 ( .A1(G113), .A2(n1275), .ZN(n1333) );
XOR2_X1 U992 ( .A(KEYINPUT62), .B(n1334), .Z(n1332) );
NOR2_X1 U993 ( .A1(G113), .A2(n1275), .ZN(n1334) );
NAND3_X1 U994 ( .A1(n1282), .A2(n1111), .A3(n1128), .ZN(n1275) );
NOR2_X1 U995 ( .A1(n1328), .A2(n1101), .ZN(n1128) );
XOR2_X1 U996 ( .A(n1099), .B(KEYINPUT35), .Z(n1328) );
INV_X1 U997 ( .A(n1213), .ZN(n1111) );
AND3_X1 U998 ( .A1(n1126), .A2(n1335), .A3(n1117), .ZN(n1282) );
NOR2_X1 U999 ( .A1(n1316), .A2(n1314), .ZN(n1117) );
INV_X1 U1000 ( .A(n1119), .ZN(n1314) );
NOR2_X1 U1001 ( .A1(n1123), .A2(n1336), .ZN(n1126) );
INV_X1 U1002 ( .A(n1124), .ZN(n1336) );
XNOR2_X1 U1003 ( .A(G110), .B(n1276), .ZN(G12) );
NAND2_X1 U1004 ( .A1(n1313), .A2(n1299), .ZN(n1276) );
NOR3_X1 U1005 ( .A1(n1119), .A2(n1118), .A3(n1284), .ZN(n1299) );
NAND2_X1 U1006 ( .A1(n1123), .A2(n1124), .ZN(n1284) );
NAND2_X1 U1007 ( .A1(G221), .A2(n1337), .ZN(n1124) );
XNOR2_X1 U1008 ( .A(G469), .B(n1338), .ZN(n1123) );
NOR2_X1 U1009 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NOR2_X1 U1010 ( .A1(KEYINPUT51), .A2(n1145), .ZN(n1340) );
AND2_X1 U1011 ( .A1(KEYINPUT43), .A2(n1145), .ZN(n1339) );
AND2_X1 U1012 ( .A1(n1341), .A2(n1342), .ZN(n1145) );
XOR2_X1 U1013 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1014 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1015 ( .A(n1234), .B(n1347), .Z(n1346) );
NOR2_X1 U1016 ( .A1(KEYINPUT27), .A2(n1348), .ZN(n1347) );
NAND2_X1 U1017 ( .A1(G227), .A2(n1163), .ZN(n1234) );
XNOR2_X1 U1018 ( .A(G140), .B(KEYINPUT1), .ZN(n1345) );
XNOR2_X1 U1019 ( .A(n1245), .B(n1349), .ZN(n1343) );
XNOR2_X1 U1020 ( .A(n1246), .B(n1239), .ZN(n1349) );
XNOR2_X1 U1021 ( .A(n1350), .B(n1351), .ZN(n1245) );
XNOR2_X1 U1022 ( .A(KEYINPUT60), .B(n1352), .ZN(n1351) );
XNOR2_X1 U1023 ( .A(G104), .B(n1353), .ZN(n1350) );
XNOR2_X1 U1024 ( .A(G902), .B(KEYINPUT56), .ZN(n1341) );
INV_X1 U1025 ( .A(n1316), .ZN(n1118) );
NAND3_X1 U1026 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1316) );
INV_X1 U1027 ( .A(n1134), .ZN(n1356) );
NOR2_X1 U1028 ( .A1(n1196), .A2(n1192), .ZN(n1134) );
NAND2_X1 U1029 ( .A1(KEYINPUT23), .A2(n1141), .ZN(n1355) );
OR3_X1 U1030 ( .A1(n1140), .A2(KEYINPUT23), .A3(n1141), .ZN(n1354) );
INV_X1 U1031 ( .A(n1192), .ZN(n1141) );
NOR2_X1 U1032 ( .A1(n1199), .A2(G902), .ZN(n1192) );
INV_X1 U1033 ( .A(n1195), .ZN(n1199) );
XNOR2_X1 U1034 ( .A(n1357), .B(n1358), .ZN(n1195) );
XOR2_X1 U1035 ( .A(n1359), .B(n1360), .Z(n1358) );
XNOR2_X1 U1036 ( .A(G128), .B(G137), .ZN(n1360) );
NAND3_X1 U1037 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1359) );
OR2_X1 U1038 ( .A1(n1162), .A2(KEYINPUT5), .ZN(n1363) );
NAND3_X1 U1039 ( .A1(KEYINPUT5), .A2(n1364), .A3(G146), .ZN(n1362) );
OR2_X1 U1040 ( .A1(n1364), .A2(G146), .ZN(n1361) );
AND2_X1 U1041 ( .A1(KEYINPUT46), .A2(n1162), .ZN(n1364) );
XNOR2_X1 U1042 ( .A(n1290), .B(n1241), .ZN(n1162) );
XNOR2_X1 U1043 ( .A(n1365), .B(n1366), .ZN(n1357) );
XOR2_X1 U1044 ( .A(n1367), .B(n1368), .Z(n1366) );
NOR2_X1 U1045 ( .A1(G119), .A2(KEYINPUT57), .ZN(n1368) );
AND3_X1 U1046 ( .A1(G221), .A2(n1163), .A3(G234), .ZN(n1367) );
INV_X1 U1047 ( .A(n1196), .ZN(n1140) );
NAND2_X1 U1048 ( .A1(G217), .A2(n1337), .ZN(n1196) );
NAND2_X1 U1049 ( .A1(n1369), .A2(n1256), .ZN(n1337) );
XOR2_X1 U1050 ( .A(n1148), .B(n1149), .Z(n1119) );
INV_X1 U1051 ( .A(G472), .ZN(n1149) );
NAND2_X1 U1052 ( .A1(n1370), .A2(n1256), .ZN(n1148) );
XOR2_X1 U1053 ( .A(n1224), .B(n1371), .Z(n1370) );
XNOR2_X1 U1054 ( .A(n1225), .B(n1216), .ZN(n1371) );
XNOR2_X1 U1055 ( .A(n1372), .B(n1353), .ZN(n1216) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1373), .ZN(n1372) );
XNOR2_X1 U1057 ( .A(n1348), .B(n1159), .ZN(n1225) );
INV_X1 U1058 ( .A(n1231), .ZN(n1348) );
XOR2_X1 U1059 ( .A(G131), .B(n1374), .Z(n1231) );
NOR2_X1 U1060 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
NOR3_X1 U1061 ( .A1(n1377), .A2(G137), .A3(n1378), .ZN(n1376) );
INV_X1 U1062 ( .A(KEYINPUT14), .ZN(n1377) );
NOR2_X1 U1063 ( .A1(KEYINPUT14), .A2(n1158), .ZN(n1375) );
XNOR2_X1 U1064 ( .A(G137), .B(n1378), .ZN(n1158) );
XOR2_X1 U1065 ( .A(G113), .B(n1379), .Z(n1224) );
NOR2_X1 U1066 ( .A1(KEYINPUT9), .A2(n1380), .ZN(n1379) );
NOR4_X1 U1067 ( .A1(n1099), .A2(n1213), .A3(n1101), .A4(n1283), .ZN(n1313) );
INV_X1 U1068 ( .A(n1335), .ZN(n1283) );
NAND2_X1 U1069 ( .A1(n1317), .A2(n1381), .ZN(n1335) );
NAND3_X1 U1070 ( .A1(n1319), .A2(n1129), .A3(n1180), .ZN(n1381) );
NOR2_X1 U1071 ( .A1(n1163), .A2(G898), .ZN(n1180) );
XNOR2_X1 U1072 ( .A(G902), .B(KEYINPUT38), .ZN(n1319) );
NAND3_X1 U1073 ( .A1(n1129), .A2(n1163), .A3(G952), .ZN(n1317) );
NAND2_X1 U1074 ( .A1(G237), .A2(n1369), .ZN(n1129) );
XNOR2_X1 U1075 ( .A(G234), .B(KEYINPUT22), .ZN(n1369) );
NAND3_X1 U1076 ( .A1(n1382), .A2(n1383), .A3(n1384), .ZN(n1101) );
OR2_X1 U1077 ( .A1(n1139), .A2(n1138), .ZN(n1384) );
NAND2_X1 U1078 ( .A1(KEYINPUT39), .A2(n1385), .ZN(n1383) );
NAND2_X1 U1079 ( .A1(n1386), .A2(n1139), .ZN(n1385) );
XNOR2_X1 U1080 ( .A(n1138), .B(KEYINPUT34), .ZN(n1386) );
NAND2_X1 U1081 ( .A1(n1387), .A2(n1388), .ZN(n1382) );
INV_X1 U1082 ( .A(KEYINPUT39), .ZN(n1388) );
NAND2_X1 U1083 ( .A1(n1389), .A2(n1390), .ZN(n1387) );
OR2_X1 U1084 ( .A1(n1138), .A2(KEYINPUT34), .ZN(n1390) );
NAND3_X1 U1085 ( .A1(n1138), .A2(n1139), .A3(KEYINPUT34), .ZN(n1389) );
INV_X1 U1086 ( .A(G478), .ZN(n1139) );
NOR2_X1 U1087 ( .A1(n1203), .A2(G902), .ZN(n1138) );
XOR2_X1 U1088 ( .A(n1391), .B(n1392), .Z(n1203) );
XNOR2_X1 U1089 ( .A(n1393), .B(n1394), .ZN(n1392) );
XOR2_X1 U1090 ( .A(n1395), .B(n1396), .Z(n1394) );
AND3_X1 U1091 ( .A1(G234), .A2(n1163), .A3(G217), .ZN(n1396) );
NAND2_X1 U1092 ( .A1(KEYINPUT17), .A2(G116), .ZN(n1395) );
XOR2_X1 U1093 ( .A(n1397), .B(n1398), .Z(n1391) );
NOR2_X1 U1094 ( .A1(KEYINPUT18), .A2(n1378), .ZN(n1398) );
INV_X1 U1095 ( .A(G134), .ZN(n1378) );
XNOR2_X1 U1096 ( .A(G107), .B(G122), .ZN(n1397) );
NAND2_X1 U1097 ( .A1(n1112), .A2(n1113), .ZN(n1213) );
NAND2_X1 U1098 ( .A1(G214), .A2(n1399), .ZN(n1113) );
XNOR2_X1 U1099 ( .A(n1142), .B(KEYINPUT19), .ZN(n1112) );
XOR2_X1 U1100 ( .A(n1400), .B(n1255), .Z(n1142) );
NAND2_X1 U1101 ( .A1(G210), .A2(n1399), .ZN(n1255) );
NAND2_X1 U1102 ( .A1(n1401), .A2(n1256), .ZN(n1399) );
INV_X1 U1103 ( .A(G237), .ZN(n1401) );
NAND2_X1 U1104 ( .A1(n1402), .A2(n1256), .ZN(n1400) );
XNOR2_X1 U1105 ( .A(n1251), .B(n1403), .ZN(n1402) );
XNOR2_X1 U1106 ( .A(n1288), .B(n1404), .ZN(n1403) );
NAND2_X1 U1107 ( .A1(KEYINPUT54), .A2(n1405), .ZN(n1404) );
NAND2_X1 U1108 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
NAND2_X1 U1109 ( .A1(n1159), .A2(G125), .ZN(n1407) );
INV_X1 U1110 ( .A(n1246), .ZN(n1159) );
XOR2_X1 U1111 ( .A(n1408), .B(KEYINPUT25), .Z(n1406) );
NAND2_X1 U1112 ( .A1(n1246), .A2(n1290), .ZN(n1408) );
INV_X1 U1113 ( .A(G125), .ZN(n1290) );
XOR2_X1 U1114 ( .A(G146), .B(n1393), .Z(n1246) );
XOR2_X1 U1115 ( .A(G128), .B(G143), .Z(n1393) );
AND2_X1 U1116 ( .A1(G224), .A2(n1163), .ZN(n1288) );
INV_X1 U1117 ( .A(G953), .ZN(n1163) );
XNOR2_X1 U1118 ( .A(n1409), .B(n1186), .ZN(n1251) );
XNOR2_X1 U1119 ( .A(G122), .B(n1239), .ZN(n1186) );
INV_X1 U1120 ( .A(n1365), .ZN(n1239) );
XOR2_X1 U1121 ( .A(G110), .B(KEYINPUT24), .Z(n1365) );
NAND3_X1 U1122 ( .A1(n1410), .A2(n1411), .A3(n1412), .ZN(n1409) );
OR2_X1 U1123 ( .A1(n1189), .A2(KEYINPUT41), .ZN(n1412) );
NAND3_X1 U1124 ( .A1(KEYINPUT41), .A2(n1413), .A3(n1188), .ZN(n1411) );
OR2_X1 U1125 ( .A1(n1188), .A2(n1413), .ZN(n1410) );
AND2_X1 U1126 ( .A1(KEYINPUT2), .A2(n1189), .ZN(n1413) );
XOR2_X1 U1127 ( .A(n1414), .B(n1353), .Z(n1189) );
XOR2_X1 U1128 ( .A(G101), .B(KEYINPUT30), .Z(n1353) );
XOR2_X1 U1129 ( .A(n1415), .B(KEYINPUT15), .Z(n1414) );
NAND2_X1 U1130 ( .A1(n1416), .A2(n1417), .ZN(n1415) );
NAND2_X1 U1131 ( .A1(G104), .A2(n1352), .ZN(n1417) );
XOR2_X1 U1132 ( .A(KEYINPUT44), .B(n1418), .Z(n1416) );
NOR2_X1 U1133 ( .A1(G104), .A2(n1352), .ZN(n1418) );
INV_X1 U1134 ( .A(G107), .ZN(n1352) );
XNOR2_X1 U1135 ( .A(G113), .B(n1380), .ZN(n1188) );
XNOR2_X1 U1136 ( .A(G116), .B(G119), .ZN(n1380) );
XNOR2_X1 U1137 ( .A(n1419), .B(G475), .ZN(n1099) );
NAND2_X1 U1138 ( .A1(n1210), .A2(n1256), .ZN(n1419) );
INV_X1 U1139 ( .A(G902), .ZN(n1256) );
XOR2_X1 U1140 ( .A(n1420), .B(n1421), .Z(n1210) );
XOR2_X1 U1141 ( .A(n1422), .B(n1423), .Z(n1421) );
XOR2_X1 U1142 ( .A(n1424), .B(n1425), .Z(n1423) );
AND3_X1 U1143 ( .A1(G214), .A2(n1426), .A3(n1373), .ZN(n1425) );
NOR2_X1 U1144 ( .A1(G953), .A2(G237), .ZN(n1373) );
INV_X1 U1145 ( .A(KEYINPUT55), .ZN(n1426) );
NAND2_X1 U1146 ( .A1(n1427), .A2(n1428), .ZN(n1424) );
NAND2_X1 U1147 ( .A1(G125), .A2(n1241), .ZN(n1428) );
XOR2_X1 U1148 ( .A(KEYINPUT61), .B(n1429), .Z(n1427) );
NOR2_X1 U1149 ( .A1(G125), .A2(n1241), .ZN(n1429) );
INV_X1 U1150 ( .A(G140), .ZN(n1241) );
XNOR2_X1 U1151 ( .A(G104), .B(G113), .ZN(n1422) );
XOR2_X1 U1152 ( .A(n1430), .B(n1431), .Z(n1420) );
XNOR2_X1 U1153 ( .A(n1161), .B(G122), .ZN(n1431) );
INV_X1 U1154 ( .A(G131), .ZN(n1161) );
XNOR2_X1 U1155 ( .A(G143), .B(G146), .ZN(n1430) );
endmodule


