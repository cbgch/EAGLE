//Key = 1001111111010100100001001110000101111110101000001100111010000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372;

XNOR2_X1 U747 ( .A(G107), .B(n1038), .ZN(G9) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR3_X1 U749 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR3_X1 U752 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NOR3_X1 U753 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NOR2_X1 U754 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U755 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
XNOR2_X1 U756 ( .A(KEYINPUT33), .B(n1058), .ZN(n1057) );
NOR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1049) );
NOR3_X1 U758 ( .A1(n1055), .A2(n1061), .A3(n1058), .ZN(n1060) );
AND2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR3_X1 U760 ( .A1(n1055), .A2(n1064), .A3(n1051), .ZN(n1046) );
NOR3_X1 U761 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XNOR2_X1 U763 ( .A(KEYINPUT63), .B(n1058), .ZN(n1069) );
NOR2_X1 U764 ( .A1(n1070), .A2(n1071), .ZN(n1066) );
XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n1048), .ZN(n1071) );
INV_X1 U766 ( .A(n1072), .ZN(n1070) );
AND2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1065) );
NAND3_X1 U768 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1041) );
NAND3_X1 U769 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
XOR2_X1 U770 ( .A(KEYINPUT45), .B(n1081), .Z(n1080) );
NOR4_X1 U771 ( .A1(n1058), .A2(n1048), .A3(n1051), .A4(n1045), .ZN(n1081) );
INV_X1 U772 ( .A(n1082), .ZN(n1048) );
INV_X1 U773 ( .A(n1073), .ZN(n1058) );
NAND2_X1 U774 ( .A1(KEYINPUT18), .A2(n1055), .ZN(n1079) );
INV_X1 U775 ( .A(n1083), .ZN(n1055) );
NAND2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1078) );
INV_X1 U777 ( .A(KEYINPUT18), .ZN(n1085) );
NAND2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR3_X1 U779 ( .A1(n1088), .A2(G953), .A3(G952), .ZN(n1039) );
INV_X1 U780 ( .A(n1075), .ZN(n1088) );
NAND4_X1 U781 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1075) );
NOR4_X1 U782 ( .A1(n1063), .A2(n1086), .A3(n1093), .A4(n1094), .ZN(n1092) );
XNOR2_X1 U783 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U784 ( .A1(n1097), .A2(KEYINPUT22), .ZN(n1096) );
XNOR2_X1 U785 ( .A(n1098), .B(n1099), .ZN(n1093) );
NAND2_X1 U786 ( .A1(KEYINPUT25), .A2(n1100), .ZN(n1098) );
NOR2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(n1091) );
XNOR2_X1 U788 ( .A(n1103), .B(n1104), .ZN(n1102) );
XOR2_X1 U789 ( .A(n1105), .B(KEYINPUT56), .Z(n1103) );
XNOR2_X1 U790 ( .A(n1106), .B(n1107), .ZN(n1101) );
XNOR2_X1 U791 ( .A(KEYINPUT37), .B(n1108), .ZN(n1107) );
XOR2_X1 U792 ( .A(n1109), .B(n1110), .Z(G72) );
NOR2_X1 U793 ( .A1(n1111), .A2(n1076), .ZN(n1110) );
AND2_X1 U794 ( .A1(G227), .A2(G900), .ZN(n1111) );
NAND2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
NAND2_X1 U796 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1116), .A2(n1076), .ZN(n1115) );
XOR2_X1 U798 ( .A(KEYINPUT47), .B(n1117), .Z(n1114) );
AND2_X1 U799 ( .A1(n1118), .A2(n1076), .ZN(n1117) );
NAND3_X1 U800 ( .A1(n1119), .A2(n1120), .A3(n1116), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(n1116) );
XNOR2_X1 U802 ( .A(n1123), .B(n1124), .ZN(n1122) );
XNOR2_X1 U803 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR2_X1 U804 ( .A1(KEYINPUT60), .A2(n1127), .ZN(n1126) );
NOR2_X1 U805 ( .A1(G131), .A2(KEYINPUT43), .ZN(n1125) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(n1121) );
XOR2_X1 U807 ( .A(KEYINPUT49), .B(KEYINPUT27), .Z(n1129) );
XOR2_X1 U808 ( .A(n1130), .B(G134), .Z(n1128) );
NAND2_X1 U809 ( .A1(G953), .A2(n1131), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1118), .A2(n1076), .ZN(n1119) );
NAND2_X1 U811 ( .A1(n1132), .A2(n1133), .ZN(n1118) );
XOR2_X1 U812 ( .A(n1134), .B(KEYINPUT50), .Z(n1132) );
XOR2_X1 U813 ( .A(n1135), .B(n1136), .Z(G69) );
NOR2_X1 U814 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1076), .ZN(n1138) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XNOR2_X1 U817 ( .A(KEYINPUT53), .B(n1142), .ZN(n1141) );
NOR2_X1 U818 ( .A1(G953), .A2(n1143), .ZN(n1137) );
NAND2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1135) );
OR2_X1 U820 ( .A1(KEYINPUT42), .A2(n1146), .ZN(n1145) );
NAND2_X1 U821 ( .A1(KEYINPUT48), .A2(n1146), .ZN(n1144) );
NAND2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U823 ( .A1(G953), .A2(n1142), .ZN(n1148) );
XOR2_X1 U824 ( .A(n1149), .B(n1150), .Z(n1147) );
NAND2_X1 U825 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
XNOR2_X1 U826 ( .A(KEYINPUT46), .B(KEYINPUT30), .ZN(n1151) );
NOR2_X1 U827 ( .A1(n1153), .A2(n1154), .ZN(G66) );
NOR3_X1 U828 ( .A1(n1095), .A2(n1155), .A3(n1156), .ZN(n1154) );
NOR3_X1 U829 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
NOR2_X1 U830 ( .A1(n1160), .A2(n1161), .ZN(n1155) );
NOR2_X1 U831 ( .A1(n1162), .A2(n1158), .ZN(n1160) );
INV_X1 U832 ( .A(G217), .ZN(n1158) );
NOR2_X1 U833 ( .A1(n1153), .A2(n1163), .ZN(G63) );
XNOR2_X1 U834 ( .A(n1164), .B(n1165), .ZN(n1163) );
NOR2_X1 U835 ( .A1(n1166), .A2(n1159), .ZN(n1165) );
NOR2_X1 U836 ( .A1(n1153), .A2(n1167), .ZN(G60) );
NOR3_X1 U837 ( .A1(n1106), .A2(n1168), .A3(n1169), .ZN(n1167) );
NOR3_X1 U838 ( .A1(n1170), .A2(n1108), .A3(n1159), .ZN(n1169) );
INV_X1 U839 ( .A(n1171), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1171), .ZN(n1168) );
NOR2_X1 U841 ( .A1(n1162), .A2(n1108), .ZN(n1172) );
INV_X1 U842 ( .A(n1043), .ZN(n1162) );
XNOR2_X1 U843 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U844 ( .A1(n1153), .A2(n1174), .ZN(G57) );
XOR2_X1 U845 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U846 ( .A(n1177), .B(n1178), .ZN(n1176) );
XOR2_X1 U847 ( .A(n1179), .B(n1180), .Z(n1175) );
NOR2_X1 U848 ( .A1(n1181), .A2(n1159), .ZN(n1180) );
NAND2_X1 U849 ( .A1(n1182), .A2(KEYINPUT26), .ZN(n1179) );
XOR2_X1 U850 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U851 ( .A1(KEYINPUT17), .A2(n1185), .ZN(n1184) );
NOR2_X1 U852 ( .A1(n1153), .A2(n1186), .ZN(G54) );
XOR2_X1 U853 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U854 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U855 ( .A(n1130), .B(n1191), .Z(n1190) );
NOR2_X1 U856 ( .A1(KEYINPUT29), .A2(n1192), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NOR2_X1 U859 ( .A1(G110), .A2(n1197), .ZN(n1195) );
NOR2_X1 U860 ( .A1(n1198), .A2(n1199), .ZN(n1193) );
XNOR2_X1 U861 ( .A(G110), .B(KEYINPUT31), .ZN(n1199) );
NOR2_X1 U862 ( .A1(n1200), .A2(G110), .ZN(n1198) );
NOR2_X1 U863 ( .A1(G140), .A2(n1197), .ZN(n1200) );
INV_X1 U864 ( .A(KEYINPUT24), .ZN(n1197) );
XOR2_X1 U865 ( .A(n1201), .B(n1202), .Z(n1187) );
XOR2_X1 U866 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U867 ( .A1(KEYINPUT39), .A2(n1205), .ZN(n1204) );
NOR2_X1 U868 ( .A1(n1100), .A2(n1159), .ZN(n1203) );
INV_X1 U869 ( .A(G469), .ZN(n1100) );
NOR2_X1 U870 ( .A1(n1153), .A2(n1206), .ZN(G51) );
NOR2_X1 U871 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U872 ( .A(n1209), .B(n1210), .Z(n1208) );
AND2_X1 U873 ( .A1(n1211), .A2(KEYINPUT34), .ZN(n1210) );
NOR2_X1 U874 ( .A1(n1104), .A2(n1159), .ZN(n1209) );
NAND2_X1 U875 ( .A1(G902), .A2(n1043), .ZN(n1159) );
NAND3_X1 U876 ( .A1(n1133), .A2(n1134), .A3(n1143), .ZN(n1043) );
AND4_X1 U877 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1143) );
AND4_X1 U878 ( .A1(n1038), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1215) );
NAND3_X1 U879 ( .A1(n1074), .A2(n1073), .A3(n1219), .ZN(n1038) );
AND2_X1 U880 ( .A1(n1220), .A2(n1173), .ZN(n1214) );
NAND3_X1 U881 ( .A1(n1219), .A2(n1073), .A3(n1221), .ZN(n1173) );
AND4_X1 U882 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1133) );
AND4_X1 U883 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
OR2_X1 U884 ( .A1(n1230), .A2(n1056), .ZN(n1224) );
NOR2_X1 U885 ( .A1(KEYINPUT34), .A2(n1211), .ZN(n1207) );
XNOR2_X1 U886 ( .A(n1231), .B(n1232), .ZN(n1211) );
XNOR2_X1 U887 ( .A(n1233), .B(n1234), .ZN(n1232) );
XNOR2_X1 U888 ( .A(n1235), .B(n1236), .ZN(n1231) );
NOR2_X1 U889 ( .A1(n1076), .A2(G952), .ZN(n1153) );
XNOR2_X1 U890 ( .A(n1222), .B(n1237), .ZN(G48) );
NOR2_X1 U891 ( .A1(KEYINPUT12), .A2(n1238), .ZN(n1237) );
NAND3_X1 U892 ( .A1(n1221), .A2(n1239), .A3(n1240), .ZN(n1222) );
XOR2_X1 U893 ( .A(n1241), .B(G143), .Z(G45) );
NAND2_X1 U894 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
OR2_X1 U895 ( .A1(n1134), .A2(KEYINPUT15), .ZN(n1243) );
NAND2_X1 U896 ( .A1(n1244), .A2(n1245), .ZN(n1134) );
NAND3_X1 U897 ( .A1(n1245), .A2(n1054), .A3(KEYINPUT15), .ZN(n1242) );
INV_X1 U898 ( .A(n1244), .ZN(n1054) );
AND4_X1 U899 ( .A1(n1246), .A2(n1239), .A3(n1247), .A4(n1248), .ZN(n1245) );
XNOR2_X1 U900 ( .A(G140), .B(n1223), .ZN(G42) );
NAND2_X1 U901 ( .A1(n1249), .A2(n1072), .ZN(n1223) );
XNOR2_X1 U902 ( .A(G137), .B(n1229), .ZN(G39) );
NAND3_X1 U903 ( .A1(n1083), .A2(n1082), .A3(n1240), .ZN(n1229) );
XNOR2_X1 U904 ( .A(G134), .B(n1228), .ZN(G36) );
NAND4_X1 U905 ( .A1(n1083), .A2(n1244), .A3(n1246), .A4(n1074), .ZN(n1228) );
XNOR2_X1 U906 ( .A(G131), .B(n1227), .ZN(G33) );
NAND2_X1 U907 ( .A1(n1249), .A2(n1244), .ZN(n1227) );
AND3_X1 U908 ( .A1(n1221), .A2(n1246), .A3(n1083), .ZN(n1249) );
NOR2_X1 U909 ( .A1(n1250), .A2(n1086), .ZN(n1083) );
XOR2_X1 U910 ( .A(n1251), .B(n1252), .Z(G30) );
NOR2_X1 U911 ( .A1(n1253), .A2(n1056), .ZN(n1252) );
INV_X1 U912 ( .A(n1239), .ZN(n1056) );
XOR2_X1 U913 ( .A(n1230), .B(KEYINPUT51), .Z(n1253) );
NAND2_X1 U914 ( .A1(n1240), .A2(n1074), .ZN(n1230) );
AND3_X1 U915 ( .A1(n1254), .A2(n1255), .A3(n1246), .ZN(n1240) );
AND3_X1 U916 ( .A1(n1256), .A2(n1257), .A3(n1062), .ZN(n1246) );
NAND2_X1 U917 ( .A1(KEYINPUT13), .A2(n1258), .ZN(n1251) );
XNOR2_X1 U918 ( .A(G101), .B(n1220), .ZN(G3) );
NAND3_X1 U919 ( .A1(n1244), .A2(n1219), .A3(n1082), .ZN(n1220) );
XNOR2_X1 U920 ( .A(G125), .B(n1226), .ZN(G27) );
NAND4_X1 U921 ( .A1(n1239), .A2(n1256), .A3(n1072), .A4(n1259), .ZN(n1226) );
NOR2_X1 U922 ( .A1(n1051), .A2(n1068), .ZN(n1259) );
INV_X1 U923 ( .A(n1059), .ZN(n1051) );
NAND2_X1 U924 ( .A1(n1045), .A2(n1260), .ZN(n1256) );
NAND4_X1 U925 ( .A1(G953), .A2(G902), .A3(n1261), .A4(n1131), .ZN(n1260) );
INV_X1 U926 ( .A(G900), .ZN(n1131) );
XNOR2_X1 U927 ( .A(G122), .B(n1212), .ZN(G24) );
NAND4_X1 U928 ( .A1(n1262), .A2(n1073), .A3(n1247), .A4(n1248), .ZN(n1212) );
XOR2_X1 U929 ( .A(n1263), .B(KEYINPUT1), .Z(n1247) );
NOR2_X1 U930 ( .A1(n1255), .A2(n1254), .ZN(n1073) );
XOR2_X1 U931 ( .A(n1213), .B(n1264), .Z(G21) );
XOR2_X1 U932 ( .A(KEYINPUT3), .B(G119), .Z(n1264) );
NAND4_X1 U933 ( .A1(n1262), .A2(n1082), .A3(n1254), .A4(n1255), .ZN(n1213) );
XNOR2_X1 U934 ( .A(G116), .B(n1218), .ZN(G18) );
NAND3_X1 U935 ( .A1(n1244), .A2(n1074), .A3(n1262), .ZN(n1218) );
NOR2_X1 U936 ( .A1(n1263), .A2(n1089), .ZN(n1074) );
XOR2_X1 U937 ( .A(n1217), .B(n1265), .Z(G15) );
NAND2_X1 U938 ( .A1(G113), .A2(n1266), .ZN(n1265) );
XOR2_X1 U939 ( .A(KEYINPUT6), .B(KEYINPUT57), .Z(n1266) );
NAND3_X1 U940 ( .A1(n1262), .A2(n1244), .A3(n1221), .ZN(n1217) );
INV_X1 U941 ( .A(n1068), .ZN(n1221) );
NAND2_X1 U942 ( .A1(n1089), .A2(n1263), .ZN(n1068) );
INV_X1 U943 ( .A(n1248), .ZN(n1089) );
NOR2_X1 U944 ( .A1(n1254), .A2(n1090), .ZN(n1244) );
INV_X1 U945 ( .A(n1255), .ZN(n1090) );
AND2_X1 U946 ( .A1(n1059), .A2(n1267), .ZN(n1262) );
NOR2_X1 U947 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
INV_X1 U948 ( .A(n1257), .ZN(n1063) );
XNOR2_X1 U949 ( .A(G110), .B(n1216), .ZN(G12) );
NAND3_X1 U950 ( .A1(n1072), .A2(n1219), .A3(n1082), .ZN(n1216) );
NOR2_X1 U951 ( .A1(n1248), .A2(n1263), .ZN(n1082) );
XOR2_X1 U952 ( .A(n1268), .B(n1108), .Z(n1263) );
INV_X1 U953 ( .A(G475), .ZN(n1108) );
NAND2_X1 U954 ( .A1(KEYINPUT38), .A2(n1106), .ZN(n1268) );
NOR2_X1 U955 ( .A1(n1171), .A2(G902), .ZN(n1106) );
XNOR2_X1 U956 ( .A(n1269), .B(n1270), .ZN(n1171) );
XOR2_X1 U957 ( .A(n1271), .B(n1272), .Z(n1269) );
XOR2_X1 U958 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U959 ( .A(G122), .B(n1275), .ZN(n1274) );
XOR2_X1 U960 ( .A(KEYINPUT55), .B(KEYINPUT14), .Z(n1273) );
XOR2_X1 U961 ( .A(n1276), .B(n1277), .Z(n1271) );
XNOR2_X1 U962 ( .A(G104), .B(n1278), .ZN(n1277) );
NAND2_X1 U963 ( .A1(n1279), .A2(G214), .ZN(n1278) );
XOR2_X1 U964 ( .A(n1280), .B(n1123), .Z(n1276) );
NAND2_X1 U965 ( .A1(KEYINPUT35), .A2(n1281), .ZN(n1280) );
INV_X1 U966 ( .A(G131), .ZN(n1281) );
XOR2_X1 U967 ( .A(n1282), .B(n1166), .Z(n1248) );
INV_X1 U968 ( .A(G478), .ZN(n1166) );
NAND2_X1 U969 ( .A1(n1164), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U970 ( .A(n1284), .B(n1285), .ZN(n1164) );
XOR2_X1 U971 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U972 ( .A(G107), .B(n1288), .ZN(n1287) );
AND3_X1 U973 ( .A1(G217), .A2(n1076), .A3(G234), .ZN(n1288) );
NAND2_X1 U974 ( .A1(KEYINPUT8), .A2(n1289), .ZN(n1286) );
XOR2_X1 U975 ( .A(G122), .B(G116), .Z(n1289) );
XNOR2_X1 U976 ( .A(G128), .B(n1290), .ZN(n1284) );
XOR2_X1 U977 ( .A(G143), .B(G134), .Z(n1290) );
AND3_X1 U978 ( .A1(n1062), .A2(n1257), .A3(n1267), .ZN(n1219) );
AND2_X1 U979 ( .A1(n1239), .A2(n1291), .ZN(n1267) );
NAND2_X1 U980 ( .A1(n1045), .A2(n1292), .ZN(n1291) );
NAND4_X1 U981 ( .A1(G953), .A2(G902), .A3(n1261), .A4(n1142), .ZN(n1292) );
INV_X1 U982 ( .A(G898), .ZN(n1142) );
NAND3_X1 U983 ( .A1(n1261), .A2(n1076), .A3(G952), .ZN(n1045) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1261) );
NOR2_X1 U985 ( .A1(n1087), .A2(n1086), .ZN(n1239) );
AND2_X1 U986 ( .A1(G214), .A2(n1293), .ZN(n1086) );
INV_X1 U987 ( .A(n1250), .ZN(n1087) );
NAND2_X1 U988 ( .A1(n1294), .A2(n1295), .ZN(n1250) );
NAND2_X1 U989 ( .A1(n1296), .A2(n1105), .ZN(n1295) );
XOR2_X1 U990 ( .A(n1297), .B(KEYINPUT62), .Z(n1294) );
OR2_X1 U991 ( .A1(n1105), .A2(n1296), .ZN(n1297) );
INV_X1 U992 ( .A(n1104), .ZN(n1296) );
NAND2_X1 U993 ( .A1(G210), .A2(n1293), .ZN(n1104) );
NAND2_X1 U994 ( .A1(n1298), .A2(n1283), .ZN(n1293) );
INV_X1 U995 ( .A(G237), .ZN(n1298) );
NAND3_X1 U996 ( .A1(n1299), .A2(n1300), .A3(n1283), .ZN(n1105) );
OR2_X1 U997 ( .A1(n1235), .A2(n1301), .ZN(n1300) );
NAND2_X1 U998 ( .A1(n1235), .A2(n1302), .ZN(n1299) );
NAND2_X1 U999 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U1000 ( .A1(KEYINPUT16), .A2(n1301), .ZN(n1304) );
NAND2_X1 U1001 ( .A1(KEYINPUT7), .A2(n1305), .ZN(n1301) );
NAND2_X1 U1002 ( .A1(n1305), .A2(n1306), .ZN(n1303) );
INV_X1 U1003 ( .A(KEYINPUT16), .ZN(n1306) );
AND2_X1 U1004 ( .A1(n1307), .A2(n1308), .ZN(n1305) );
NAND2_X1 U1005 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND2_X1 U1006 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND2_X1 U1007 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XNOR2_X1 U1008 ( .A(KEYINPUT44), .B(n1234), .ZN(n1314) );
XNOR2_X1 U1009 ( .A(KEYINPUT61), .B(G125), .ZN(n1313) );
NAND2_X1 U1010 ( .A1(n1234), .A2(n1315), .ZN(n1311) );
XNOR2_X1 U1011 ( .A(KEYINPUT61), .B(n1233), .ZN(n1315) );
INV_X1 U1012 ( .A(G125), .ZN(n1233) );
INV_X1 U1013 ( .A(n1236), .ZN(n1309) );
NAND2_X1 U1014 ( .A1(n1316), .A2(n1236), .ZN(n1307) );
XOR2_X1 U1015 ( .A(n1234), .B(n1317), .Z(n1316) );
NOR2_X1 U1016 ( .A1(G125), .A2(KEYINPUT44), .ZN(n1317) );
NOR2_X1 U1017 ( .A1(n1140), .A2(G953), .ZN(n1234) );
INV_X1 U1018 ( .A(G224), .ZN(n1140) );
XOR2_X1 U1019 ( .A(n1150), .B(n1152), .Z(n1235) );
XNOR2_X1 U1020 ( .A(G122), .B(G110), .ZN(n1152) );
XOR2_X1 U1021 ( .A(n1318), .B(n1319), .Z(n1150) );
XOR2_X1 U1022 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1023 ( .A(KEYINPUT52), .B(KEYINPUT4), .Z(n1321) );
NOR2_X1 U1024 ( .A1(KEYINPUT19), .A2(n1275), .ZN(n1320) );
INV_X1 U1025 ( .A(G113), .ZN(n1275) );
XOR2_X1 U1026 ( .A(n1201), .B(n1322), .Z(n1318) );
NAND2_X1 U1027 ( .A1(n1323), .A2(n1324), .ZN(n1257) );
XNOR2_X1 U1028 ( .A(G221), .B(KEYINPUT9), .ZN(n1323) );
XNOR2_X1 U1029 ( .A(n1099), .B(G469), .ZN(n1062) );
NAND2_X1 U1030 ( .A1(n1325), .A2(n1326), .ZN(n1099) );
XOR2_X1 U1031 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1032 ( .A(n1196), .B(G110), .ZN(n1328) );
INV_X1 U1033 ( .A(G140), .ZN(n1196) );
XNOR2_X1 U1034 ( .A(n1329), .B(n1189), .ZN(n1327) );
NAND2_X1 U1035 ( .A1(G227), .A2(n1076), .ZN(n1189) );
NAND2_X1 U1036 ( .A1(n1330), .A2(KEYINPUT0), .ZN(n1329) );
XOR2_X1 U1037 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1038 ( .A(n1333), .B(n1205), .ZN(n1332) );
NAND2_X1 U1039 ( .A1(KEYINPUT54), .A2(n1201), .ZN(n1333) );
XNOR2_X1 U1040 ( .A(G101), .B(n1334), .ZN(n1201) );
XNOR2_X1 U1041 ( .A(n1335), .B(G104), .ZN(n1334) );
INV_X1 U1042 ( .A(G107), .ZN(n1335) );
XOR2_X1 U1043 ( .A(n1130), .B(KEYINPUT5), .Z(n1331) );
NAND3_X1 U1044 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n1130) );
NAND2_X1 U1045 ( .A1(KEYINPUT41), .A2(G128), .ZN(n1338) );
OR3_X1 U1046 ( .A1(G128), .A2(KEYINPUT41), .A3(n1270), .ZN(n1337) );
NAND2_X1 U1047 ( .A1(n1270), .A2(n1339), .ZN(n1336) );
NAND2_X1 U1048 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
INV_X1 U1049 ( .A(KEYINPUT41), .ZN(n1341) );
XNOR2_X1 U1050 ( .A(G128), .B(KEYINPUT10), .ZN(n1340) );
XNOR2_X1 U1051 ( .A(G143), .B(n1238), .ZN(n1270) );
XNOR2_X1 U1052 ( .A(G902), .B(KEYINPUT20), .ZN(n1325) );
NOR2_X1 U1053 ( .A1(n1255), .A2(n1342), .ZN(n1072) );
INV_X1 U1054 ( .A(n1254), .ZN(n1342) );
XOR2_X1 U1055 ( .A(n1095), .B(n1097), .Z(n1254) );
AND2_X1 U1056 ( .A1(n1343), .A2(G217), .ZN(n1097) );
XOR2_X1 U1057 ( .A(n1324), .B(KEYINPUT23), .Z(n1343) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1283), .ZN(n1324) );
NOR2_X1 U1059 ( .A1(n1161), .A2(G902), .ZN(n1095) );
INV_X1 U1060 ( .A(n1157), .ZN(n1161) );
XNOR2_X1 U1061 ( .A(n1344), .B(n1345), .ZN(n1157) );
XOR2_X1 U1062 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1063 ( .A(G119), .B(G110), .Z(n1347) );
XNOR2_X1 U1064 ( .A(KEYINPUT59), .B(n1258), .ZN(n1346) );
INV_X1 U1065 ( .A(G128), .ZN(n1258) );
XNOR2_X1 U1066 ( .A(n1123), .B(n1348), .ZN(n1344) );
XNOR2_X1 U1067 ( .A(n1349), .B(n1350), .ZN(n1348) );
NOR2_X1 U1068 ( .A1(KEYINPUT28), .A2(n1238), .ZN(n1350) );
NAND2_X1 U1069 ( .A1(KEYINPUT36), .A2(n1351), .ZN(n1349) );
XNOR2_X1 U1070 ( .A(n1127), .B(n1352), .ZN(n1351) );
AND3_X1 U1071 ( .A1(G221), .A2(n1076), .A3(G234), .ZN(n1352) );
INV_X1 U1072 ( .A(G953), .ZN(n1076) );
XOR2_X1 U1073 ( .A(G140), .B(G125), .Z(n1123) );
XOR2_X1 U1074 ( .A(n1353), .B(n1181), .Z(n1255) );
INV_X1 U1075 ( .A(G472), .ZN(n1181) );
NAND2_X1 U1076 ( .A1(n1354), .A2(n1283), .ZN(n1353) );
INV_X1 U1077 ( .A(G902), .ZN(n1283) );
XOR2_X1 U1078 ( .A(n1183), .B(n1355), .Z(n1354) );
XNOR2_X1 U1079 ( .A(n1356), .B(n1185), .ZN(n1355) );
INV_X1 U1080 ( .A(G101), .ZN(n1185) );
NAND3_X1 U1081 ( .A1(n1357), .A2(n1358), .A3(n1359), .ZN(n1356) );
NAND2_X1 U1082 ( .A1(KEYINPUT58), .A2(n1360), .ZN(n1359) );
NAND3_X1 U1083 ( .A1(n1177), .A2(n1361), .A3(n1178), .ZN(n1358) );
INV_X1 U1084 ( .A(n1362), .ZN(n1178) );
NAND2_X1 U1085 ( .A1(n1362), .A2(n1363), .ZN(n1357) );
NAND2_X1 U1086 ( .A1(n1364), .A2(n1361), .ZN(n1363) );
INV_X1 U1087 ( .A(KEYINPUT58), .ZN(n1361) );
XNOR2_X1 U1088 ( .A(KEYINPUT32), .B(n1360), .ZN(n1364) );
INV_X1 U1089 ( .A(n1177), .ZN(n1360) );
XNOR2_X1 U1090 ( .A(n1365), .B(n1322), .ZN(n1177) );
XOR2_X1 U1091 ( .A(G116), .B(G119), .Z(n1322) );
XNOR2_X1 U1092 ( .A(G113), .B(KEYINPUT11), .ZN(n1365) );
XNOR2_X1 U1093 ( .A(n1236), .B(n1366), .ZN(n1362) );
INV_X1 U1094 ( .A(n1205), .ZN(n1366) );
XOR2_X1 U1095 ( .A(G131), .B(n1367), .Z(n1205) );
XNOR2_X1 U1096 ( .A(n1127), .B(G134), .ZN(n1367) );
INV_X1 U1097 ( .A(G137), .ZN(n1127) );
XNOR2_X1 U1098 ( .A(n1368), .B(n1369), .ZN(n1236) );
NOR2_X1 U1099 ( .A1(G128), .A2(KEYINPUT2), .ZN(n1369) );
NAND2_X1 U1100 ( .A1(n1370), .A2(n1371), .ZN(n1368) );
NAND2_X1 U1101 ( .A1(G143), .A2(n1238), .ZN(n1371) );
XOR2_X1 U1102 ( .A(KEYINPUT40), .B(n1372), .Z(n1370) );
NOR2_X1 U1103 ( .A1(G143), .A2(n1238), .ZN(n1372) );
INV_X1 U1104 ( .A(G146), .ZN(n1238) );
NAND2_X1 U1105 ( .A1(n1279), .A2(G210), .ZN(n1183) );
NOR2_X1 U1106 ( .A1(G953), .A2(G237), .ZN(n1279) );
endmodule


