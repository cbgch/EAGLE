//Key = 1110000001000001010100101011111000011000101100000111111100110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303;

XNOR2_X1 U727 ( .A(n996), .B(n997), .ZN(G9) );
NOR2_X1 U728 ( .A1(KEYINPUT39), .A2(n998), .ZN(n997) );
NOR2_X1 U729 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U730 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
NOR2_X1 U731 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U732 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR3_X1 U733 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
NOR3_X1 U734 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
NOR4_X1 U735 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1014) );
OR2_X1 U736 ( .A1(n1019), .A2(KEYINPUT48), .ZN(n1016) );
INV_X1 U737 ( .A(n1020), .ZN(n1015) );
NOR2_X1 U738 ( .A1(n1021), .A2(n1022), .ZN(n1012) );
NOR3_X1 U739 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1021) );
NOR2_X1 U740 ( .A1(n1019), .A2(n1026), .ZN(n1025) );
NOR2_X1 U741 ( .A1(KEYINPUT48), .A2(n1017), .ZN(n1026) );
AND3_X1 U742 ( .A1(n1019), .A2(n1027), .A3(KEYINPUT29), .ZN(n1024) );
NOR2_X1 U743 ( .A1(KEYINPUT29), .A2(n1027), .ZN(n1023) );
NOR4_X1 U744 ( .A1(n1019), .A2(n1028), .A3(n1017), .A4(n1022), .ZN(n1007) );
NOR3_X1 U745 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR3_X1 U746 ( .A1(n1032), .A2(KEYINPUT36), .A3(n1033), .ZN(n1031) );
NOR2_X1 U747 ( .A1(n1034), .A2(n1011), .ZN(n1030) );
INV_X1 U748 ( .A(n1032), .ZN(n1011) );
NOR2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
AND2_X1 U750 ( .A1(n1037), .A2(KEYINPUT36), .ZN(n1035) );
NOR2_X1 U751 ( .A1(n1038), .A2(n1009), .ZN(n1029) );
INV_X1 U752 ( .A(n1039), .ZN(n1009) );
NOR2_X1 U753 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR3_X1 U754 ( .A1(n1002), .A2(G952), .A3(n1003), .ZN(n999) );
AND4_X1 U755 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1003) );
NOR4_X1 U756 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
XOR2_X1 U757 ( .A(n1050), .B(KEYINPUT18), .Z(n1046) );
NAND2_X1 U758 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U759 ( .A(n1053), .B(KEYINPUT45), .Z(n1051) );
XNOR2_X1 U760 ( .A(n1054), .B(KEYINPUT3), .ZN(n1044) );
XNOR2_X1 U761 ( .A(n1055), .B(n1056), .ZN(n1042) );
INV_X1 U762 ( .A(n1057), .ZN(n1002) );
XOR2_X1 U763 ( .A(n1058), .B(n1059), .Z(G72) );
XOR2_X1 U764 ( .A(n1060), .B(n1061), .Z(n1059) );
NAND3_X1 U765 ( .A1(n1062), .A2(n1063), .A3(KEYINPUT0), .ZN(n1061) );
NAND2_X1 U766 ( .A1(G953), .A2(n1064), .ZN(n1063) );
XOR2_X1 U767 ( .A(n1065), .B(n1066), .Z(n1062) );
NOR2_X1 U768 ( .A1(KEYINPUT33), .A2(n1067), .ZN(n1065) );
XOR2_X1 U769 ( .A(n1068), .B(n1069), .Z(n1067) );
XOR2_X1 U770 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U771 ( .A1(G131), .A2(KEYINPUT11), .ZN(n1070) );
NAND2_X1 U772 ( .A1(n1072), .A2(n1073), .ZN(n1060) );
XNOR2_X1 U773 ( .A(KEYINPUT62), .B(n1074), .ZN(n1072) );
NOR2_X1 U774 ( .A1(n1075), .A2(n1074), .ZN(n1058) );
AND2_X1 U775 ( .A1(G227), .A2(G900), .ZN(n1075) );
XOR2_X1 U776 ( .A(n1076), .B(n1077), .Z(G69) );
XOR2_X1 U777 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR3_X1 U778 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
INV_X1 U780 ( .A(KEYINPUT40), .ZN(n1084) );
NOR2_X1 U781 ( .A1(KEYINPUT40), .A2(n1085), .ZN(n1081) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U783 ( .A1(KEYINPUT25), .A2(n1088), .ZN(n1078) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U785 ( .A1(KEYINPUT57), .A2(n1091), .ZN(n1090) );
INV_X1 U786 ( .A(n1080), .ZN(n1091) );
NOR2_X1 U787 ( .A1(n1092), .A2(n1074), .ZN(n1089) );
NOR2_X1 U788 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
AND2_X1 U789 ( .A1(G898), .A2(KEYINPUT57), .ZN(n1093) );
NOR2_X1 U790 ( .A1(n1095), .A2(G953), .ZN(n1076) );
NOR2_X1 U791 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XNOR2_X1 U792 ( .A(n1098), .B(KEYINPUT53), .ZN(n1097) );
XNOR2_X1 U793 ( .A(n1099), .B(n1100), .ZN(n1096) );
NOR2_X1 U794 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U795 ( .A1(n1098), .A2(n1103), .ZN(G63) );
XNOR2_X1 U796 ( .A(n1104), .B(n1105), .ZN(n1103) );
NOR2_X1 U797 ( .A1(n1106), .A2(n1102), .ZN(n1105) );
NOR2_X1 U798 ( .A1(n1098), .A2(n1107), .ZN(G60) );
XOR2_X1 U799 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U800 ( .A(KEYINPUT51), .B(KEYINPUT37), .Z(n1109) );
XOR2_X1 U801 ( .A(n1110), .B(n1111), .Z(n1108) );
NOR2_X1 U802 ( .A1(n1112), .A2(n1102), .ZN(n1111) );
XOR2_X1 U803 ( .A(G104), .B(n1113), .Z(G6) );
NOR2_X1 U804 ( .A1(n1098), .A2(n1114), .ZN(G57) );
XOR2_X1 U805 ( .A(n1115), .B(n1116), .Z(n1114) );
XNOR2_X1 U806 ( .A(n1117), .B(n1118), .ZN(n1116) );
XOR2_X1 U807 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U808 ( .A(n1121), .B(n1122), .Z(n1115) );
NOR2_X1 U809 ( .A1(n1056), .A2(n1102), .ZN(n1122) );
INV_X1 U810 ( .A(G472), .ZN(n1056) );
XOR2_X1 U811 ( .A(n1123), .B(KEYINPUT2), .Z(n1121) );
NOR2_X1 U812 ( .A1(n1098), .A2(n1124), .ZN(G54) );
XOR2_X1 U813 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U814 ( .A(n1127), .B(n1128), .ZN(n1126) );
XOR2_X1 U815 ( .A(n1120), .B(n1068), .Z(n1128) );
XOR2_X1 U816 ( .A(n1129), .B(n1130), .Z(n1125) );
NOR2_X1 U817 ( .A1(n1131), .A2(n1102), .ZN(n1130) );
XOR2_X1 U818 ( .A(n1132), .B(n1133), .Z(n1129) );
NAND3_X1 U819 ( .A1(n1134), .A2(n1135), .A3(KEYINPUT19), .ZN(n1132) );
NOR2_X1 U820 ( .A1(n1098), .A2(n1136), .ZN(G51) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U822 ( .A(n1083), .B(n1139), .Z(n1138) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(n1137) );
NOR3_X1 U824 ( .A1(n1102), .A2(KEYINPUT23), .A3(n1142), .ZN(n1141) );
NAND2_X1 U825 ( .A1(G902), .A2(n1001), .ZN(n1102) );
NAND2_X1 U826 ( .A1(n1095), .A2(n1143), .ZN(n1001) );
INV_X1 U827 ( .A(n1073), .ZN(n1143) );
NAND4_X1 U828 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1073) );
NOR4_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1147) );
INV_X1 U830 ( .A(n1152), .ZN(n1150) );
INV_X1 U831 ( .A(n1153), .ZN(n1149) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(n1146) );
NOR2_X1 U833 ( .A1(n1022), .A2(n1156), .ZN(n1155) );
AND3_X1 U834 ( .A1(n1157), .A2(n1041), .A3(n1036), .ZN(n1154) );
NAND3_X1 U835 ( .A1(n1158), .A2(n1040), .A3(n1159), .ZN(n1144) );
XNOR2_X1 U836 ( .A(n1160), .B(KEYINPUT59), .ZN(n1159) );
AND4_X1 U837 ( .A1(n1161), .A2(n996), .A3(n1162), .A4(n1163), .ZN(n1095) );
NOR4_X1 U838 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1113), .ZN(n1163) );
AND4_X1 U839 ( .A1(n1041), .A2(n1039), .A3(n1167), .A4(n1168), .ZN(n1113) );
NOR3_X1 U840 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1162) );
AND3_X1 U841 ( .A1(KEYINPUT7), .A2(n1172), .A3(n1173), .ZN(n1171) );
NOR2_X1 U842 ( .A1(KEYINPUT7), .A2(n1174), .ZN(n1170) );
INV_X1 U843 ( .A(n1175), .ZN(n1169) );
NAND4_X1 U844 ( .A1(n1039), .A2(n1167), .A3(n1040), .A4(n1168), .ZN(n996) );
NAND2_X1 U845 ( .A1(G224), .A2(n1074), .ZN(n1140) );
NOR2_X1 U846 ( .A1(n1074), .A2(G952), .ZN(n1098) );
XNOR2_X1 U847 ( .A(G146), .B(n1153), .ZN(G48) );
NAND3_X1 U848 ( .A1(n1160), .A2(n1041), .A3(n1158), .ZN(n1153) );
XNOR2_X1 U849 ( .A(G143), .B(n1145), .ZN(G45) );
NAND4_X1 U850 ( .A1(n1158), .A2(n1037), .A3(n1054), .A4(n1176), .ZN(n1145) );
XNOR2_X1 U851 ( .A(G140), .B(n1177), .ZN(G42) );
NAND4_X1 U852 ( .A1(KEYINPUT1), .A2(n1157), .A3(n1036), .A4(n1041), .ZN(n1177) );
XOR2_X1 U853 ( .A(G137), .B(n1178), .Z(G39) );
NOR2_X1 U854 ( .A1(n1179), .A2(n1022), .ZN(n1178) );
XOR2_X1 U855 ( .A(n1156), .B(KEYINPUT16), .Z(n1179) );
NAND3_X1 U856 ( .A1(n1160), .A2(n1032), .A3(n1180), .ZN(n1156) );
NOR3_X1 U857 ( .A1(n1181), .A2(n1027), .A3(n1019), .ZN(n1180) );
XOR2_X1 U858 ( .A(n1148), .B(n1182), .Z(G36) );
XOR2_X1 U859 ( .A(KEYINPUT8), .B(G134), .Z(n1182) );
AND3_X1 U860 ( .A1(n1037), .A2(n1040), .A3(n1157), .ZN(n1148) );
XOR2_X1 U861 ( .A(G131), .B(n1151), .Z(G33) );
AND3_X1 U862 ( .A1(n1041), .A2(n1037), .A3(n1157), .ZN(n1151) );
NOR4_X1 U863 ( .A1(n1022), .A2(n1181), .A3(n1019), .A4(n1027), .ZN(n1157) );
INV_X1 U864 ( .A(n1183), .ZN(n1019) );
INV_X1 U865 ( .A(n1184), .ZN(n1181) );
NAND2_X1 U866 ( .A1(n1020), .A2(n1018), .ZN(n1022) );
XNOR2_X1 U867 ( .A(G128), .B(n1185), .ZN(G30) );
NAND3_X1 U868 ( .A1(n1160), .A2(n1040), .A3(n1158), .ZN(n1185) );
AND2_X1 U869 ( .A1(n1167), .A2(n1184), .ZN(n1158) );
XNOR2_X1 U870 ( .A(n1186), .B(n1166), .ZN(G3) );
NOR2_X1 U871 ( .A1(n1187), .A2(n1033), .ZN(n1166) );
INV_X1 U872 ( .A(n1037), .ZN(n1033) );
XNOR2_X1 U873 ( .A(G125), .B(n1152), .ZN(G27) );
NAND4_X1 U874 ( .A1(n1036), .A2(n1041), .A3(n1013), .A4(n1184), .ZN(n1152) );
NAND2_X1 U875 ( .A1(n1006), .A2(n1188), .ZN(n1184) );
NAND4_X1 U876 ( .A1(G902), .A2(G953), .A3(n1189), .A4(n1064), .ZN(n1188) );
INV_X1 U877 ( .A(G900), .ZN(n1064) );
XOR2_X1 U878 ( .A(n1165), .B(n1190), .Z(G24) );
NOR2_X1 U879 ( .A1(KEYINPUT44), .A2(n1191), .ZN(n1190) );
AND4_X1 U880 ( .A1(n1192), .A2(n1039), .A3(n1054), .A4(n1176), .ZN(n1165) );
NOR2_X1 U881 ( .A1(n1047), .A2(n1193), .ZN(n1039) );
XOR2_X1 U882 ( .A(G119), .B(n1194), .Z(G21) );
NOR2_X1 U883 ( .A1(KEYINPUT46), .A2(n1175), .ZN(n1194) );
NAND3_X1 U884 ( .A1(n1192), .A2(n1032), .A3(n1160), .ZN(n1175) );
AND2_X1 U885 ( .A1(n1193), .A2(n1047), .ZN(n1160) );
INV_X1 U886 ( .A(n1195), .ZN(n1193) );
XOR2_X1 U887 ( .A(G116), .B(n1164), .Z(G18) );
AND3_X1 U888 ( .A1(n1192), .A2(n1040), .A3(n1037), .ZN(n1164) );
AND2_X1 U889 ( .A1(n1196), .A2(n1176), .ZN(n1040) );
XNOR2_X1 U890 ( .A(KEYINPUT55), .B(n1197), .ZN(n1196) );
XNOR2_X1 U891 ( .A(G113), .B(n1161), .ZN(G15) );
NAND3_X1 U892 ( .A1(n1037), .A2(n1192), .A3(n1041), .ZN(n1161) );
AND2_X1 U893 ( .A1(n1013), .A2(n1168), .ZN(n1192) );
NOR3_X1 U894 ( .A1(n1020), .A2(n1048), .A3(n1017), .ZN(n1013) );
NOR2_X1 U895 ( .A1(n1195), .A2(n1047), .ZN(n1037) );
XOR2_X1 U896 ( .A(n1174), .B(n1198), .Z(G12) );
XOR2_X1 U897 ( .A(KEYINPUT17), .B(G110), .Z(n1198) );
NAND2_X1 U898 ( .A1(n1036), .A2(n1173), .ZN(n1174) );
INV_X1 U899 ( .A(n1187), .ZN(n1173) );
NAND3_X1 U900 ( .A1(n1032), .A2(n1168), .A3(n1167), .ZN(n1187) );
NOR3_X1 U901 ( .A1(n1020), .A2(n1027), .A3(n1048), .ZN(n1167) );
NAND2_X1 U902 ( .A1(n1018), .A2(n1183), .ZN(n1048) );
NAND2_X1 U903 ( .A1(G221), .A2(n1199), .ZN(n1183) );
NAND2_X1 U904 ( .A1(G214), .A2(n1200), .ZN(n1018) );
INV_X1 U905 ( .A(n1017), .ZN(n1027) );
NAND2_X1 U906 ( .A1(n1053), .A2(n1052), .ZN(n1017) );
NAND3_X1 U907 ( .A1(n1131), .A2(n1201), .A3(n1202), .ZN(n1052) );
INV_X1 U908 ( .A(G469), .ZN(n1131) );
NAND2_X1 U909 ( .A1(G469), .A2(n1203), .ZN(n1053) );
NAND2_X1 U910 ( .A1(n1202), .A2(n1201), .ZN(n1203) );
XNOR2_X1 U911 ( .A(n1204), .B(n1120), .ZN(n1202) );
XOR2_X1 U912 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U913 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U914 ( .A(n1209), .B(KEYINPUT43), .Z(n1208) );
NAND3_X1 U915 ( .A1(n1210), .A2(n1135), .A3(n1133), .ZN(n1209) );
NOR2_X1 U916 ( .A1(n1211), .A2(n1133), .ZN(n1207) );
AND2_X1 U917 ( .A1(n1212), .A2(G227), .ZN(n1133) );
XNOR2_X1 U918 ( .A(G953), .B(KEYINPUT20), .ZN(n1212) );
AND2_X1 U919 ( .A1(n1135), .A2(n1210), .ZN(n1211) );
XNOR2_X1 U920 ( .A(n1134), .B(KEYINPUT54), .ZN(n1210) );
NAND2_X1 U921 ( .A1(G110), .A2(n1213), .ZN(n1134) );
OR2_X1 U922 ( .A1(n1213), .A2(G110), .ZN(n1135) );
INV_X1 U923 ( .A(G140), .ZN(n1213) );
NAND2_X1 U924 ( .A1(n1214), .A2(KEYINPUT22), .ZN(n1205) );
XOR2_X1 U925 ( .A(n1215), .B(n1068), .Z(n1214) );
XNOR2_X1 U926 ( .A(n1216), .B(n1217), .ZN(n1068) );
XNOR2_X1 U927 ( .A(G146), .B(KEYINPUT27), .ZN(n1216) );
NAND2_X1 U928 ( .A1(KEYINPUT35), .A2(n1127), .ZN(n1215) );
XOR2_X1 U929 ( .A(n1186), .B(n1218), .Z(n1127) );
XOR2_X1 U930 ( .A(n1049), .B(KEYINPUT49), .Z(n1020) );
XNOR2_X1 U931 ( .A(n1219), .B(n1220), .ZN(n1049) );
NOR2_X1 U932 ( .A1(n1142), .A2(n1221), .ZN(n1220) );
XNOR2_X1 U933 ( .A(KEYINPUT21), .B(n1200), .ZN(n1221) );
OR2_X1 U934 ( .A1(G902), .A2(G237), .ZN(n1200) );
NAND2_X1 U935 ( .A1(n1222), .A2(n1201), .ZN(n1219) );
XOR2_X1 U936 ( .A(n1083), .B(n1223), .Z(n1222) );
NOR2_X1 U937 ( .A1(KEYINPUT10), .A2(n1224), .ZN(n1223) );
XOR2_X1 U938 ( .A(n1225), .B(n1226), .Z(n1224) );
NOR2_X1 U939 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NOR3_X1 U940 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1228) );
AND2_X1 U941 ( .A1(n1229), .A2(n1139), .ZN(n1227) );
XNOR2_X1 U942 ( .A(G125), .B(n1230), .ZN(n1139) );
INV_X1 U943 ( .A(KEYINPUT60), .ZN(n1229) );
NOR3_X1 U944 ( .A1(n1094), .A2(KEYINPUT5), .A3(G953), .ZN(n1225) );
INV_X1 U945 ( .A(G224), .ZN(n1094) );
XOR2_X1 U946 ( .A(n1086), .B(n1087), .Z(n1083) );
XOR2_X1 U947 ( .A(n1191), .B(G110), .Z(n1087) );
XNOR2_X1 U948 ( .A(n1119), .B(n1232), .ZN(n1086) );
NOR2_X1 U949 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
AND3_X1 U950 ( .A1(KEYINPUT12), .A2(n998), .A3(G104), .ZN(n1234) );
NOR2_X1 U951 ( .A1(KEYINPUT12), .A2(n1218), .ZN(n1233) );
XNOR2_X1 U952 ( .A(G104), .B(n998), .ZN(n1218) );
XNOR2_X1 U953 ( .A(n1235), .B(G101), .ZN(n1119) );
NAND2_X1 U954 ( .A1(n1006), .A2(n1236), .ZN(n1168) );
NAND3_X1 U955 ( .A1(n1080), .A2(n1189), .A3(G902), .ZN(n1236) );
NOR2_X1 U956 ( .A1(n1074), .A2(G898), .ZN(n1080) );
NAND3_X1 U957 ( .A1(n1057), .A2(n1189), .A3(G952), .ZN(n1006) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1189) );
XOR2_X1 U959 ( .A(G953), .B(KEYINPUT28), .Z(n1057) );
NAND2_X1 U960 ( .A1(n1237), .A2(n1238), .ZN(n1032) );
NAND2_X1 U961 ( .A1(n1041), .A2(n1239), .ZN(n1238) );
INV_X1 U962 ( .A(KEYINPUT55), .ZN(n1239) );
NOR2_X1 U963 ( .A1(n1176), .A2(n1197), .ZN(n1041) );
NAND3_X1 U964 ( .A1(n1197), .A2(n1043), .A3(KEYINPUT55), .ZN(n1237) );
INV_X1 U965 ( .A(n1176), .ZN(n1043) );
XOR2_X1 U966 ( .A(n1240), .B(n1106), .Z(n1176) );
INV_X1 U967 ( .A(G478), .ZN(n1106) );
NAND2_X1 U968 ( .A1(n1104), .A2(n1201), .ZN(n1240) );
XNOR2_X1 U969 ( .A(n1241), .B(n1242), .ZN(n1104) );
XOR2_X1 U970 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U971 ( .A(n998), .B(n1245), .ZN(n1244) );
AND3_X1 U972 ( .A1(G217), .A2(n1074), .A3(G234), .ZN(n1245) );
INV_X1 U973 ( .A(G107), .ZN(n998) );
XNOR2_X1 U974 ( .A(n1246), .B(G116), .ZN(n1243) );
XOR2_X1 U975 ( .A(n1247), .B(n1248), .Z(n1241) );
NOR2_X1 U976 ( .A1(KEYINPUT47), .A2(n1249), .ZN(n1248) );
XOR2_X1 U977 ( .A(n1250), .B(n1251), .Z(n1247) );
NOR2_X1 U978 ( .A1(G134), .A2(KEYINPUT32), .ZN(n1251) );
NAND2_X1 U979 ( .A1(KEYINPUT9), .A2(n1191), .ZN(n1250) );
INV_X1 U980 ( .A(n1054), .ZN(n1197) );
XOR2_X1 U981 ( .A(n1252), .B(n1112), .Z(n1054) );
INV_X1 U982 ( .A(G475), .ZN(n1112) );
NAND2_X1 U983 ( .A1(n1110), .A2(n1201), .ZN(n1252) );
XOR2_X1 U984 ( .A(n1253), .B(n1254), .Z(n1110) );
XOR2_X1 U985 ( .A(n1255), .B(n1256), .Z(n1253) );
NOR2_X1 U986 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U987 ( .A(n1259), .B(KEYINPUT15), .Z(n1258) );
NAND2_X1 U988 ( .A1(n1260), .A2(G131), .ZN(n1259) );
NOR2_X1 U989 ( .A1(G131), .A2(n1260), .ZN(n1257) );
XNOR2_X1 U990 ( .A(n1261), .B(n1249), .ZN(n1260) );
INV_X1 U991 ( .A(G143), .ZN(n1249) );
NAND3_X1 U992 ( .A1(G214), .A2(n1074), .A3(n1262), .ZN(n1261) );
XNOR2_X1 U993 ( .A(G237), .B(KEYINPUT41), .ZN(n1262) );
NAND2_X1 U994 ( .A1(n1263), .A2(KEYINPUT30), .ZN(n1255) );
XOR2_X1 U995 ( .A(n1264), .B(G104), .Z(n1263) );
NAND2_X1 U996 ( .A1(KEYINPUT24), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U997 ( .A(n1266), .B(n1267), .ZN(n1265) );
XNOR2_X1 U998 ( .A(KEYINPUT61), .B(n1191), .ZN(n1267) );
INV_X1 U999 ( .A(G122), .ZN(n1191) );
INV_X1 U1000 ( .A(G113), .ZN(n1266) );
INV_X1 U1001 ( .A(n1172), .ZN(n1036) );
NAND2_X1 U1002 ( .A1(n1047), .A2(n1195), .ZN(n1172) );
XNOR2_X1 U1003 ( .A(n1055), .B(n1268), .ZN(n1195) );
NOR2_X1 U1004 ( .A1(G472), .A2(KEYINPUT14), .ZN(n1268) );
NAND3_X1 U1005 ( .A1(n1269), .A2(n1270), .A3(n1201), .ZN(n1055) );
NAND2_X1 U1006 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U1007 ( .A(n1273), .B(n1274), .Z(n1271) );
OR3_X1 U1008 ( .A1(n1273), .A2(n1274), .A3(n1272), .ZN(n1269) );
INV_X1 U1009 ( .A(KEYINPUT34), .ZN(n1272) );
XNOR2_X1 U1010 ( .A(n1275), .B(n1276), .ZN(n1274) );
XOR2_X1 U1011 ( .A(KEYINPUT6), .B(KEYINPUT13), .Z(n1276) );
XNOR2_X1 U1012 ( .A(n1123), .B(n1186), .ZN(n1275) );
INV_X1 U1013 ( .A(G101), .ZN(n1186) );
OR3_X1 U1014 ( .A1(G237), .A2(G953), .A3(n1142), .ZN(n1123) );
INV_X1 U1015 ( .A(G210), .ZN(n1142) );
XOR2_X1 U1016 ( .A(n1277), .B(n1278), .Z(n1273) );
XNOR2_X1 U1017 ( .A(n1279), .B(KEYINPUT52), .ZN(n1278) );
NAND2_X1 U1018 ( .A1(KEYINPUT58), .A2(n1120), .ZN(n1279) );
XOR2_X1 U1019 ( .A(G131), .B(n1071), .Z(n1120) );
XOR2_X1 U1020 ( .A(G134), .B(G137), .Z(n1071) );
XNOR2_X1 U1021 ( .A(n1280), .B(n1230), .ZN(n1277) );
INV_X1 U1022 ( .A(n1117), .ZN(n1230) );
XNOR2_X1 U1023 ( .A(n1281), .B(n1217), .ZN(n1117) );
XNOR2_X1 U1024 ( .A(n1246), .B(G143), .ZN(n1217) );
XOR2_X1 U1025 ( .A(n1282), .B(KEYINPUT38), .Z(n1281) );
NAND2_X1 U1026 ( .A1(KEYINPUT26), .A2(n1283), .ZN(n1282) );
INV_X1 U1027 ( .A(G146), .ZN(n1283) );
NAND2_X1 U1028 ( .A1(KEYINPUT50), .A2(n1235), .ZN(n1280) );
XOR2_X1 U1029 ( .A(G113), .B(n1284), .Z(n1235) );
XOR2_X1 U1030 ( .A(G119), .B(G116), .Z(n1284) );
XOR2_X1 U1031 ( .A(n1285), .B(n1101), .Z(n1047) );
NAND2_X1 U1032 ( .A1(G217), .A2(n1199), .ZN(n1101) );
NAND2_X1 U1033 ( .A1(G234), .A2(n1201), .ZN(n1199) );
NAND2_X1 U1034 ( .A1(n1099), .A2(n1201), .ZN(n1285) );
INV_X1 U1035 ( .A(G902), .ZN(n1201) );
XNOR2_X1 U1036 ( .A(n1286), .B(n1287), .ZN(n1099) );
AND3_X1 U1037 ( .A1(G221), .A2(n1074), .A3(G234), .ZN(n1287) );
INV_X1 U1038 ( .A(G953), .ZN(n1074) );
XOR2_X1 U1039 ( .A(n1288), .B(G137), .Z(n1286) );
NAND2_X1 U1040 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U1041 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND2_X1 U1042 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
OR2_X1 U1043 ( .A1(n1295), .A2(KEYINPUT31), .ZN(n1294) );
INV_X1 U1044 ( .A(KEYINPUT56), .ZN(n1293) );
NAND2_X1 U1045 ( .A1(n1295), .A2(n1296), .ZN(n1289) );
NAND2_X1 U1046 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
OR2_X1 U1047 ( .A1(n1291), .A2(KEYINPUT56), .ZN(n1298) );
XNOR2_X1 U1048 ( .A(n1254), .B(KEYINPUT63), .ZN(n1291) );
XOR2_X1 U1049 ( .A(G146), .B(n1066), .Z(n1254) );
XNOR2_X1 U1050 ( .A(n1231), .B(G140), .ZN(n1066) );
INV_X1 U1051 ( .A(G125), .ZN(n1231) );
INV_X1 U1052 ( .A(KEYINPUT31), .ZN(n1297) );
NAND2_X1 U1053 ( .A1(n1299), .A2(n1300), .ZN(n1295) );
NAND2_X1 U1054 ( .A1(n1301), .A2(n1246), .ZN(n1300) );
INV_X1 U1055 ( .A(G128), .ZN(n1246) );
XOR2_X1 U1056 ( .A(KEYINPUT4), .B(n1302), .Z(n1301) );
NAND2_X1 U1057 ( .A1(n1303), .A2(G128), .ZN(n1299) );
XOR2_X1 U1058 ( .A(KEYINPUT42), .B(n1302), .Z(n1303) );
XOR2_X1 U1059 ( .A(G119), .B(G110), .Z(n1302) );
endmodule


