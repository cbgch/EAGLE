//Key = 1110100100110011011111001110001000100001100100
module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, 
        G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, 
        G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, G3, G6, G9, G12, G30, 
        G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, 
        G60, G63, G66, G69, G72, G57 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921;

  XOR2_X1 U530 ( .A(n702), .B(n703), .Z(G9) );
  NOR2_X1 U531 ( .A1(n704), .A2(n705), .ZN(G75) );
  NOR4_X1 U532 ( .A1(n706), .A2(n707), .A3(n708), .A4(n709), .ZN(n705) );
  NOR3_X1 U533 ( .A1(n710), .A2(n711), .A3(n712), .ZN(n707) );
  NOR2_X1 U534 ( .A1(n713), .A2(n714), .ZN(n711) );
  NAND3_X1 U535 ( .A1(n715), .A2(n716), .A3(n717), .ZN(n710) );
  NAND2_X1 U536 ( .A1(n718), .A2(n719), .ZN(n717) );
  INV_X1 U537 ( .A(n720), .ZN(n719) );
  NAND2_X1 U538 ( .A1(n721), .A2(n722), .ZN(n718) );
  OR2_X1 U539 ( .A1(n723), .A2(n724), .ZN(n722) );
  NAND2_X1 U540 ( .A1(n725), .A2(n726), .ZN(n716) );
  INV_X1 U541 ( .A(n727), .ZN(n726) );
  NAND2_X1 U542 ( .A1(n728), .A2(n729), .ZN(n725) );
  NAND2_X1 U543 ( .A1(n730), .A2(n731), .ZN(n729) );
  NAND2_X1 U544 ( .A1(n732), .A2(n733), .ZN(n715) );
  INV_X1 U545 ( .A(n734), .ZN(n733) );
  NAND2_X1 U546 ( .A1(n735), .A2(n736), .ZN(n732) );
  OR2_X1 U547 ( .A1(n737), .A2(n738), .ZN(n736) );
  NOR3_X1 U548 ( .A1(n708), .A2(G952), .A3(n706), .ZN(n704) );
  AND2_X1 U549 ( .A1(n727), .A2(n728), .ZN(n706) );
  AND2_X1 U550 ( .A1(n735), .A2(n734), .ZN(n728) );
  XOR2_X1 U551 ( .A(n739), .B(n740), .Z(G72) );
  XOR2_X1 U552 ( .A(n741), .B(n742), .Z(n740) );
  NOR2_X1 U553 ( .A1(n743), .A2(n744), .ZN(n742) );
  NOR2_X1 U554 ( .A1(n745), .A2(n746), .ZN(n743) );
  NAND2_X1 U555 ( .A1(n747), .A2(n748), .ZN(n741) );
  NAND2_X1 U556 ( .A1(n708), .A2(n746), .ZN(n748) );
  XOR2_X1 U557 ( .A(n749), .B(n750), .Z(n747) );
  XOR2_X1 U558 ( .A(n751), .B(n752), .Z(n750) );
  NAND2_X1 U559 ( .A1(n744), .A2(n753), .ZN(n739) );
  XOR2_X1 U560 ( .A(n754), .B(n755), .Z(G69) );
  XOR2_X1 U561 ( .A(n756), .B(n757), .Z(n755) );
  NAND2_X1 U562 ( .A1(n708), .A2(n758), .ZN(n757) );
  NAND2_X1 U563 ( .A1(G898), .A2(G224), .ZN(n758) );
  NAND2_X1 U564 ( .A1(n759), .A2(n760), .ZN(n756) );
  NAND2_X1 U565 ( .A1(n708), .A2(n761), .ZN(n760) );
  XOR2_X1 U566 ( .A(n762), .B(n763), .Z(n759) );
  NOR2_X1 U567 ( .A1(n764), .A2(n708), .ZN(n754) );
  NOR2_X1 U568 ( .A1(n765), .A2(n766), .ZN(G66) );
  XOR2_X1 U569 ( .A(n767), .B(n768), .Z(n766) );
  NAND2_X1 U570 ( .A1(n769), .A2(n770), .ZN(n767) );
  NOR2_X1 U571 ( .A1(n765), .A2(n771), .ZN(G63) );
  XOR2_X1 U572 ( .A(n772), .B(n773), .Z(n771) );
  NAND2_X1 U573 ( .A1(n769), .A2(G478), .ZN(n772) );
  NOR2_X1 U574 ( .A1(n765), .A2(n774), .ZN(G60) );
  XOR2_X1 U575 ( .A(n775), .B(n776), .Z(n774) );
  NAND2_X1 U576 ( .A1(n769), .A2(G475), .ZN(n775) );
  XOR2_X1 U577 ( .A(n777), .B(n778), .Z(G6) );
  NOR2_X1 U578 ( .A1(n765), .A2(n779), .ZN(G57) );
  XOR2_X1 U579 ( .A(n780), .B(n781), .Z(n779) );
  NAND2_X1 U580 ( .A1(n769), .A2(G472), .ZN(n780) );
  NOR2_X1 U581 ( .A1(n765), .A2(n782), .ZN(G54) );
  XOR2_X1 U582 ( .A(n783), .B(n784), .Z(n782) );
  NAND2_X1 U583 ( .A1(n769), .A2(G469), .ZN(n783) );
  NOR2_X1 U584 ( .A1(n765), .A2(n785), .ZN(G51) );
  XOR2_X1 U585 ( .A(n786), .B(n787), .Z(n785) );
  NAND2_X1 U586 ( .A1(n769), .A2(n788), .ZN(n786) );
  AND2_X1 U587 ( .A1(G902), .A2(n709), .ZN(n769) );
  NAND2_X1 U588 ( .A1(n789), .A2(n764), .ZN(n709) );
  AND4_X1 U589 ( .A1(n790), .A2(n791), .A3(n792), .A4(n793), .ZN(n764) );
  AND4_X1 U590 ( .A1(n702), .A2(n794), .A3(n795), .A4(n796), .ZN(n793) );
  NAND3_X1 U591 ( .A1(n734), .A2(n797), .A3(n723), .ZN(n702) );
  AND2_X1 U592 ( .A1(n798), .A2(n777), .ZN(n792) );
  NAND3_X1 U593 ( .A1(n734), .A2(n797), .A3(n724), .ZN(n777) );
  XOR2_X1 U594 ( .A(keyinput43), .B(n799), .Z(n791) );
  XOR2_X1 U595 ( .A(n800), .B(keyinput44), .Z(n790) );
  INV_X1 U596 ( .A(n753), .ZN(n789) );
  NAND4_X1 U597 ( .A1(n801), .A2(n802), .A3(n803), .A4(n804), .ZN(n753) );
  NOR4_X1 U598 ( .A1(n805), .A2(n806), .A3(n807), .A4(n808), .ZN(n804) );
  NOR2_X1 U599 ( .A1(n809), .A2(n810), .ZN(n803) );
  XOR2_X1 U600 ( .A(keyinput42), .B(n811), .Z(n810) );
  XOR2_X1 U601 ( .A(n812), .B(keyinput45), .Z(n802) );
  XOR2_X1 U602 ( .A(n813), .B(keyinput41), .Z(n801) );
  NOR2_X1 U603 ( .A1(n744), .A2(G952), .ZN(n765) );
  XOR2_X1 U604 ( .A(n811), .B(n814), .Z(G48) );
  AND3_X1 U605 ( .A1(n724), .A2(n815), .A3(n816), .ZN(n811) );
  XNOR2_X1 U606 ( .A(n809), .B(n817), .ZN(G45) );
  AND4_X1 U607 ( .A1(n818), .A2(n815), .A3(n819), .A4(n820), .ZN(n809) );
  XOR2_X1 U608 ( .A(n821), .B(n808), .Z(G42) );
  AND3_X1 U609 ( .A1(n727), .A2(n713), .A3(n822), .ZN(n808) );
  XOR2_X1 U610 ( .A(n807), .B(n823), .Z(G39) );
  AND3_X1 U611 ( .A1(n727), .A2(n720), .A3(n816), .ZN(n807) );
  XNOR2_X1 U612 ( .A(n806), .B(n824), .ZN(G36) );
  AND3_X1 U613 ( .A1(n727), .A2(n723), .A3(n818), .ZN(n806) );
  XOR2_X1 U614 ( .A(n812), .B(n825), .Z(G33) );
  NAND3_X1 U615 ( .A1(n724), .A2(n727), .A3(n818), .ZN(n812) );
  AND3_X1 U616 ( .A1(n713), .A2(n826), .A3(n738), .ZN(n818) );
  NOR2_X1 U617 ( .A1(n730), .A2(n827), .ZN(n727) );
  AND2_X1 U618 ( .A1(G214), .A2(n828), .ZN(n827) );
  XNOR2_X1 U619 ( .A(n829), .B(n813), .ZN(G30) );
  NAND3_X1 U620 ( .A1(n723), .A2(n815), .A3(n816), .ZN(n813) );
  AND4_X1 U621 ( .A1(n713), .A2(n830), .A3(n831), .A4(n826), .ZN(n816) );
  XOR2_X1 U622 ( .A(n798), .B(n832), .Z(G3) );
  NAND3_X1 U623 ( .A1(n720), .A2(n797), .A3(n738), .ZN(n798) );
  XOR2_X1 U624 ( .A(n805), .B(n833), .Z(G27) );
  AND3_X1 U625 ( .A1(n721), .A2(n815), .A3(n822), .ZN(n805) );
  AND4_X1 U626 ( .A1(n737), .A2(n724), .A3(n831), .A4(n826), .ZN(n822) );
  NAND2_X1 U627 ( .A1(n712), .A2(n834), .ZN(n826) );
  NAND4_X1 U628 ( .A1(n708), .A2(G902), .A3(n835), .A4(n746), .ZN(n834) );
  INV_X1 U629 ( .A(G900), .ZN(n746) );
  XOR2_X1 U630 ( .A(n796), .B(n836), .Z(G24) );
  NAND4_X1 U631 ( .A1(n721), .A2(n734), .A3(n837), .A4(n838), .ZN(n796) );
  NOR2_X1 U632 ( .A1(n839), .A2(n840), .ZN(n837) );
  NOR2_X1 U633 ( .A1(n831), .A2(n830), .ZN(n734) );
  XOR2_X1 U634 ( .A(n795), .B(n841), .Z(G21) );
  NAND4_X1 U635 ( .A1(n735), .A2(n838), .A3(n830), .A4(n831), .ZN(n795) );
  AND2_X1 U636 ( .A1(n720), .A2(n721), .ZN(n735) );
  XOR2_X1 U637 ( .A(n800), .B(n842), .Z(G18) );
  NAND2_X1 U638 ( .A1(n843), .A2(n723), .ZN(n800) );
  NOR2_X1 U639 ( .A1(n819), .A2(n839), .ZN(n723) );
  INV_X1 U640 ( .A(n820), .ZN(n839) );
  XOR2_X1 U641 ( .A(n844), .B(n799), .Z(G15) );
  AND2_X1 U642 ( .A1(n843), .A2(n724), .ZN(n799) );
  NOR2_X1 U643 ( .A1(n820), .A2(n840), .ZN(n724) );
  INV_X1 U644 ( .A(n819), .ZN(n840) );
  AND3_X1 U645 ( .A1(n721), .A2(n838), .A3(n738), .ZN(n843) );
  NOR2_X1 U646 ( .A1(n831), .A2(n737), .ZN(n738) );
  AND2_X1 U647 ( .A1(n714), .A2(n845), .ZN(n721) );
  NAND2_X1 U648 ( .A1(G221), .A2(n846), .ZN(n845) );
  XOR2_X1 U649 ( .A(n794), .B(n847), .Z(G12) );
  NAND4_X1 U650 ( .A1(n720), .A2(n797), .A3(n737), .A4(n831), .ZN(n794) );
  XNOR2_X1 U651 ( .A(n848), .B(n770), .ZN(n831) );
  AND2_X1 U652 ( .A1(G217), .A2(n846), .ZN(n770) );
  NAND2_X1 U653 ( .A1(n768), .A2(n849), .ZN(n848) );
  XNOR2_X1 U654 ( .A(n850), .B(n851), .ZN(n768) );
  XOR2_X1 U655 ( .A(n749), .B(n852), .Z(n851) );
  XOR2_X1 U656 ( .A(n853), .B(n854), .Z(n852) );
  XOR2_X1 U657 ( .A(n855), .B(n856), .Z(n850) );
  XNOR2_X1 U658 ( .A(n857), .B(n858), .ZN(n856) );
  NAND2_X1 U659 ( .A1(G221), .A2(n859), .ZN(n857) );
  XNOR2_X1 U660 ( .A(n860), .B(n861), .ZN(n855) );
  INV_X1 U661 ( .A(n830), .ZN(n737) );
  XNOR2_X1 U662 ( .A(n862), .B(G472), .ZN(n830) );
  NAND2_X1 U663 ( .A1(n781), .A2(n849), .ZN(n862) );
  XNOR2_X1 U664 ( .A(n863), .B(n864), .ZN(n781) );
  INV_X1 U665 ( .A(n865), .ZN(n864) );
  XOR2_X1 U666 ( .A(n866), .B(n867), .Z(n863) );
  AND2_X1 U667 ( .A1(n868), .A2(G210), .ZN(n867) );
  AND2_X1 U668 ( .A1(n838), .A2(n713), .ZN(n797) );
  NOR2_X1 U669 ( .A1(n714), .A2(n869), .ZN(n713) );
  AND2_X1 U670 ( .A1(G221), .A2(n846), .ZN(n869) );
  NAND2_X1 U671 ( .A1(G234), .A2(n849), .ZN(n846) );
  XOR2_X1 U672 ( .A(n870), .B(G469), .Z(n714) );
  NAND2_X1 U673 ( .A1(n784), .A2(n849), .ZN(n870) );
  XOR2_X1 U674 ( .A(n871), .B(n872), .Z(n784) );
  XOR2_X1 U675 ( .A(n873), .B(n874), .Z(n872) );
  NOR2_X1 U676 ( .A1(n708), .A2(n745), .ZN(n873) );
  INV_X1 U677 ( .A(G227), .ZN(n745) );
  XOR2_X1 U678 ( .A(n866), .B(n875), .Z(n871) );
  XOR2_X1 U679 ( .A(n876), .B(n752), .Z(n866) );
  XNOR2_X1 U680 ( .A(n877), .B(n878), .ZN(n752) );
  XNOR2_X1 U681 ( .A(n879), .B(n860), .ZN(n878) );
  XNOR2_X1 U682 ( .A(n823), .B(keyinput29), .ZN(n860) );
  XOR2_X1 U683 ( .A(keyinput13), .B(G137), .Z(n823) );
  XOR2_X1 U684 ( .A(n880), .B(n881), .Z(n877) );
  XOR2_X1 U685 ( .A(keyinput40), .B(keyinput39), .Z(n881) );
  AND2_X1 U686 ( .A1(n815), .A2(n882), .ZN(n838) );
  NAND2_X1 U687 ( .A1(n712), .A2(n883), .ZN(n882) );
  NAND4_X1 U688 ( .A1(n708), .A2(G902), .A3(n835), .A4(n761), .ZN(n883) );
  INV_X1 U689 ( .A(G898), .ZN(n761) );
  NAND3_X1 U690 ( .A1(n744), .A2(n835), .A3(G952), .ZN(n712) );
  NAND2_X1 U691 ( .A1(G237), .A2(G234), .ZN(n835) );
  INV_X1 U692 ( .A(n731), .ZN(n815) );
  NAND2_X1 U693 ( .A1(n730), .A2(n884), .ZN(n731) );
  NAND2_X1 U694 ( .A1(G214), .A2(n828), .ZN(n884) );
  XNOR2_X1 U695 ( .A(n885), .B(n788), .ZN(n730) );
  AND2_X1 U696 ( .A1(G210), .A2(n828), .ZN(n788) );
  OR2_X1 U697 ( .A1(G902), .A2(G237), .ZN(n828) );
  NAND2_X1 U698 ( .A1(n787), .A2(n849), .ZN(n885) );
  XOR2_X1 U699 ( .A(n886), .B(n887), .Z(n787) );
  XOR2_X1 U700 ( .A(n888), .B(n763), .Z(n887) );
  XNOR2_X1 U701 ( .A(n889), .B(n890), .ZN(n763) );
  XNOR2_X1 U702 ( .A(n865), .B(n875), .ZN(n889) );
  XNOR2_X1 U703 ( .A(n891), .B(n892), .ZN(n875) );
  XOR2_X1 U704 ( .A(n853), .B(n893), .Z(n892) );
  XOR2_X1 U705 ( .A(n847), .B(keyinput20), .Z(n853) );
  XNOR2_X1 U706 ( .A(keyinput3), .B(G110), .ZN(n847) );
  XOR2_X1 U707 ( .A(n894), .B(n895), .Z(n891) );
  XOR2_X1 U708 ( .A(keyinput34), .B(keyinput33), .Z(n895) );
  XNOR2_X1 U709 ( .A(n896), .B(n897), .ZN(n865) );
  XNOR2_X1 U710 ( .A(n898), .B(n854), .ZN(n897) );
  XOR2_X1 U711 ( .A(n841), .B(keyinput23), .Z(n854) );
  XNOR2_X1 U712 ( .A(keyinput6), .B(G119), .ZN(n841) );
  XOR2_X1 U713 ( .A(n899), .B(n900), .Z(n896) );
  XOR2_X1 U714 ( .A(keyinput36), .B(keyinput35), .Z(n900) );
  XOR2_X1 U715 ( .A(n876), .B(n901), .Z(n886) );
  AND2_X1 U716 ( .A1(n744), .A2(G224), .ZN(n901) );
  XOR2_X1 U717 ( .A(n762), .B(n751), .Z(n876) );
  XNOR2_X1 U718 ( .A(n902), .B(n903), .ZN(n751) );
  XNOR2_X1 U719 ( .A(n904), .B(n905), .ZN(n903) );
  INV_X1 U720 ( .A(n858), .ZN(n904) );
  XNOR2_X1 U721 ( .A(keyinput38), .B(keyinput37), .ZN(n902) );
  XNOR2_X1 U722 ( .A(n832), .B(keyinput9), .ZN(n762) );
  XOR2_X1 U723 ( .A(keyinput0), .B(G101), .Z(n832) );
  NOR2_X1 U724 ( .A1(n820), .A2(n819), .ZN(n720) );
  XNOR2_X1 U725 ( .A(n906), .B(G475), .ZN(n819) );
  NAND2_X1 U726 ( .A1(n776), .A2(n849), .ZN(n906) );
  XOR2_X1 U727 ( .A(n907), .B(n908), .Z(n776) );
  XOR2_X1 U728 ( .A(n909), .B(n910), .Z(n908) );
  XOR2_X1 U729 ( .A(n893), .B(n879), .Z(n910) );
  XOR2_X1 U730 ( .A(n825), .B(keyinput27), .Z(n879) );
  XOR2_X1 U731 ( .A(keyinput11), .B(G131), .Z(n825) );
  XNOR2_X1 U732 ( .A(n778), .B(keyinput18), .ZN(n893) );
  XOR2_X1 U733 ( .A(keyinput1), .B(G104), .Z(n778) );
  XOR2_X1 U734 ( .A(n911), .B(n905), .Z(n909) );
  XNOR2_X1 U735 ( .A(n861), .B(n912), .ZN(n905) );
  XNOR2_X1 U736 ( .A(n814), .B(keyinput32), .ZN(n861) );
  XOR2_X1 U737 ( .A(keyinput16), .B(G146), .Z(n814) );
  NAND2_X1 U738 ( .A1(G214), .A2(n868), .ZN(n911) );
  NOR2_X1 U739 ( .A1(n708), .A2(G237), .ZN(n868) );
  INV_X1 U740 ( .A(n744), .ZN(n708) );
  XOR2_X1 U741 ( .A(n913), .B(n749), .Z(n907) );
  XNOR2_X1 U742 ( .A(n888), .B(n874), .ZN(n749) );
  XNOR2_X1 U743 ( .A(n821), .B(keyinput30), .ZN(n874) );
  XNOR2_X1 U744 ( .A(keyinput14), .B(G140), .ZN(n821) );
  XNOR2_X1 U745 ( .A(n833), .B(keyinput25), .ZN(n888) );
  XOR2_X1 U746 ( .A(keyinput8), .B(G125), .Z(n833) );
  XNOR2_X1 U747 ( .A(n914), .B(n898), .ZN(n913) );
  XNOR2_X1 U748 ( .A(n844), .B(keyinput21), .ZN(n898) );
  XNOR2_X1 U749 ( .A(keyinput4), .B(G113), .ZN(n844) );
  XNOR2_X1 U750 ( .A(n915), .B(G478), .ZN(n820) );
  NAND2_X1 U751 ( .A1(n773), .A2(n849), .ZN(n915) );
  INV_X1 U752 ( .A(G902), .ZN(n849) );
  XOR2_X1 U753 ( .A(n916), .B(n917), .Z(n773) );
  XNOR2_X1 U754 ( .A(n890), .B(n918), .ZN(n917) );
  XOR2_X1 U755 ( .A(n894), .B(n899), .Z(n918) );
  XOR2_X1 U756 ( .A(n842), .B(keyinput22), .Z(n899) );
  XNOR2_X1 U757 ( .A(keyinput5), .B(G116), .ZN(n842) );
  XNOR2_X1 U758 ( .A(n703), .B(keyinput19), .ZN(n894) );
  XOR2_X1 U759 ( .A(keyinput2), .B(G107), .Z(n703) );
  INV_X1 U760 ( .A(n914), .ZN(n890) );
  XOR2_X1 U761 ( .A(n836), .B(keyinput24), .Z(n914) );
  XOR2_X1 U762 ( .A(keyinput7), .B(G122), .Z(n836) );
  XOR2_X1 U763 ( .A(n919), .B(n920), .Z(n916) );
  XNOR2_X1 U764 ( .A(n921), .B(n858), .ZN(n920) );
  XNOR2_X1 U765 ( .A(n829), .B(keyinput26), .ZN(n858) );
  XNOR2_X1 U766 ( .A(keyinput10), .B(G128), .ZN(n829) );
  NAND2_X1 U767 ( .A1(G217), .A2(n859), .ZN(n921) );
  AND2_X1 U768 ( .A1(G234), .A2(n744), .ZN(n859) );
  XOR2_X1 U769 ( .A(keyinput17), .B(G953), .Z(n744) );
  XOR2_X1 U770 ( .A(n880), .B(n912), .Z(n919) );
  XOR2_X1 U771 ( .A(n817), .B(keyinput31), .Z(n912) );
  XOR2_X1 U772 ( .A(keyinput15), .B(G143), .Z(n817) );
  XOR2_X1 U773 ( .A(n824), .B(keyinput28), .Z(n880) );
  XNOR2_X1 U774 ( .A(keyinput12), .B(G134), .ZN(n824) );
endmodule

