//Key = 1000110011000001100001101101100011101010111010111111011100000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396;

XOR2_X1 U757 ( .A(G107), .B(n1061), .Z(G9) );
NOR2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR3_X1 U759 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NOR2_X1 U760 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U761 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1067) );
NOR3_X1 U762 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NOR2_X1 U763 ( .A1(KEYINPUT5), .A2(n1075), .ZN(n1074) );
AND3_X1 U764 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NOR2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1073) );
INV_X1 U766 ( .A(KEYINPUT5), .ZN(n1080) );
NOR3_X1 U767 ( .A1(n1077), .A2(n1081), .A3(n1082), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR2_X1 U769 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U770 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
XOR2_X1 U771 ( .A(n1089), .B(KEYINPUT24), .Z(n1088) );
NOR2_X1 U772 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NOR2_X1 U773 ( .A1(n1092), .A2(n1093), .ZN(n1083) );
NOR2_X1 U774 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR3_X1 U775 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1094) );
AND2_X1 U776 ( .A1(n1099), .A2(n1079), .ZN(n1069) );
NAND3_X1 U777 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1064) );
NAND3_X1 U778 ( .A1(n1103), .A2(n1104), .A3(n1079), .ZN(n1102) );
NOR3_X1 U779 ( .A1(n1093), .A2(n1086), .A3(n1077), .ZN(n1079) );
OR2_X1 U780 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
AND3_X1 U781 ( .A1(n1100), .A2(n1101), .A3(n1107), .ZN(n1062) );
NAND4_X1 U782 ( .A1(n1108), .A2(n1109), .A3(n1078), .A4(n1091), .ZN(n1100) );
XOR2_X1 U783 ( .A(n1110), .B(KEYINPUT4), .Z(n1109) );
NAND4_X1 U784 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1110) );
NOR3_X1 U785 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NOR2_X1 U786 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U787 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U788 ( .A(KEYINPUT29), .B(n1122), .Z(n1121) );
NOR3_X1 U789 ( .A1(n1123), .A2(n1122), .A3(n1120), .ZN(n1116) );
XOR2_X1 U790 ( .A(n1124), .B(n1125), .Z(n1112) );
XOR2_X1 U791 ( .A(n1126), .B(KEYINPUT50), .Z(n1125) );
NAND2_X1 U792 ( .A1(n1122), .A2(n1120), .ZN(n1111) );
INV_X1 U793 ( .A(KEYINPUT54), .ZN(n1120) );
NOR2_X1 U794 ( .A1(n1127), .A2(n1128), .ZN(n1108) );
NOR2_X1 U795 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U796 ( .A(KEYINPUT58), .B(n1131), .Z(n1130) );
NOR2_X1 U797 ( .A1(n1132), .A2(n1133), .ZN(n1127) );
XOR2_X1 U798 ( .A(KEYINPUT27), .B(n1131), .Z(n1133) );
INV_X1 U799 ( .A(n1129), .ZN(n1132) );
XOR2_X1 U800 ( .A(n1134), .B(n1135), .Z(G72) );
XOR2_X1 U801 ( .A(n1136), .B(n1137), .Z(n1135) );
NOR2_X1 U802 ( .A1(n1138), .A2(n1101), .ZN(n1137) );
AND2_X1 U803 ( .A1(G227), .A2(G900), .ZN(n1138) );
NAND2_X1 U804 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NAND2_X1 U805 ( .A1(G953), .A2(n1141), .ZN(n1140) );
XOR2_X1 U806 ( .A(n1142), .B(n1143), .Z(n1139) );
XOR2_X1 U807 ( .A(KEYINPUT39), .B(n1144), .Z(n1143) );
NOR2_X1 U808 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR2_X1 U809 ( .A1(n1147), .A2(G125), .ZN(n1146) );
NOR2_X1 U810 ( .A1(KEYINPUT26), .A2(n1148), .ZN(n1147) );
NOR2_X1 U811 ( .A1(G140), .A2(KEYINPUT20), .ZN(n1148) );
NOR2_X1 U812 ( .A1(n1149), .A2(n1150), .ZN(n1145) );
NOR2_X1 U813 ( .A1(n1151), .A2(KEYINPUT20), .ZN(n1149) );
NOR2_X1 U814 ( .A1(KEYINPUT26), .A2(n1152), .ZN(n1151) );
NAND2_X1 U815 ( .A1(n1101), .A2(n1153), .ZN(n1134) );
XOR2_X1 U816 ( .A(n1154), .B(n1155), .Z(G69) );
XOR2_X1 U817 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U818 ( .A1(G953), .A2(n1158), .ZN(n1157) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1158) );
NAND2_X1 U820 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
NAND2_X1 U821 ( .A1(G953), .A2(n1161), .ZN(n1160) );
AND2_X1 U822 ( .A1(n1162), .A2(n1101), .ZN(n1154) );
NOR2_X1 U823 ( .A1(n1163), .A2(n1164), .ZN(G66) );
NOR3_X1 U824 ( .A1(n1122), .A2(n1165), .A3(n1166), .ZN(n1164) );
NOR3_X1 U825 ( .A1(n1167), .A2(n1123), .A3(n1168), .ZN(n1166) );
INV_X1 U826 ( .A(n1169), .ZN(n1167) );
NOR2_X1 U827 ( .A1(n1170), .A2(n1169), .ZN(n1165) );
NOR2_X1 U828 ( .A1(n1171), .A2(n1123), .ZN(n1170) );
NOR2_X1 U829 ( .A1(n1163), .A2(n1172), .ZN(G63) );
XNOR2_X1 U830 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR2_X1 U831 ( .A1(n1175), .A2(n1168), .ZN(n1174) );
INV_X1 U832 ( .A(G478), .ZN(n1175) );
NOR2_X1 U833 ( .A1(n1163), .A2(n1176), .ZN(G60) );
NOR3_X1 U834 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
NOR3_X1 U835 ( .A1(n1180), .A2(n1126), .A3(n1168), .ZN(n1179) );
NOR2_X1 U836 ( .A1(n1181), .A2(n1182), .ZN(n1178) );
INV_X1 U837 ( .A(n1180), .ZN(n1182) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1126), .ZN(n1181) );
XOR2_X1 U839 ( .A(G104), .B(n1183), .Z(G6) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1184), .ZN(G57) );
XOR2_X1 U841 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U842 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U843 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
OR2_X1 U844 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U845 ( .A(n1193), .B(KEYINPUT3), .Z(n1189) );
NAND2_X1 U846 ( .A1(n1192), .A2(n1191), .ZN(n1193) );
XNOR2_X1 U847 ( .A(n1194), .B(n1195), .ZN(n1185) );
NOR2_X1 U848 ( .A1(KEYINPUT2), .A2(n1196), .ZN(n1195) );
NOR3_X1 U849 ( .A1(n1168), .A2(KEYINPUT63), .A3(n1197), .ZN(n1194) );
INV_X1 U850 ( .A(G472), .ZN(n1197) );
NOR3_X1 U851 ( .A1(n1198), .A2(n1163), .A3(n1199), .ZN(G54) );
NOR4_X1 U852 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1168), .ZN(n1199) );
NOR2_X1 U853 ( .A1(KEYINPUT14), .A2(n1203), .ZN(n1201) );
INV_X1 U854 ( .A(n1204), .ZN(n1203) );
NOR2_X1 U855 ( .A1(n1205), .A2(n1204), .ZN(n1200) );
NOR2_X1 U856 ( .A1(KEYINPUT14), .A2(n1206), .ZN(n1205) );
NOR2_X1 U857 ( .A1(n1207), .A2(n1208), .ZN(n1198) );
NOR2_X1 U858 ( .A1(n1202), .A2(n1168), .ZN(n1208) );
INV_X1 U859 ( .A(G469), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1204), .A2(n1206), .ZN(n1207) );
INV_X1 U861 ( .A(KEYINPUT21), .ZN(n1206) );
XOR2_X1 U862 ( .A(n1209), .B(n1210), .Z(n1204) );
XOR2_X1 U863 ( .A(n1211), .B(n1212), .Z(n1209) );
NAND3_X1 U864 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1211) );
NAND2_X1 U865 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U866 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
OR2_X1 U867 ( .A1(n1218), .A2(KEYINPUT44), .ZN(n1214) );
NAND3_X1 U868 ( .A1(n1220), .A2(n1218), .A3(KEYINPUT44), .ZN(n1213) );
XOR2_X1 U869 ( .A(n1221), .B(n1222), .Z(n1218) );
INV_X1 U870 ( .A(n1219), .ZN(n1220) );
XOR2_X1 U871 ( .A(n1223), .B(n1224), .Z(n1219) );
XOR2_X1 U872 ( .A(KEYINPUT61), .B(KEYINPUT15), .Z(n1224) );
NOR2_X1 U873 ( .A1(n1163), .A2(n1225), .ZN(G51) );
XOR2_X1 U874 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U875 ( .A1(n1129), .A2(n1168), .ZN(n1227) );
NAND2_X1 U876 ( .A1(G902), .A2(n1066), .ZN(n1168) );
INV_X1 U877 ( .A(n1171), .ZN(n1066) );
NOR2_X1 U878 ( .A1(n1162), .A2(n1153), .ZN(n1171) );
NAND4_X1 U879 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1153) );
NOR4_X1 U880 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1231) );
INV_X1 U881 ( .A(n1236), .ZN(n1235) );
NAND3_X1 U882 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1230) );
NAND3_X1 U883 ( .A1(n1095), .A2(n1240), .A3(n1076), .ZN(n1228) );
NAND2_X1 U884 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND3_X1 U885 ( .A1(n1105), .A2(n1237), .A3(n1243), .ZN(n1242) );
XOR2_X1 U886 ( .A(n1244), .B(KEYINPUT60), .Z(n1243) );
NAND3_X1 U887 ( .A1(n1099), .A2(n1244), .A3(n1106), .ZN(n1241) );
NAND4_X1 U888 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1162) );
NOR4_X1 U889 ( .A1(n1249), .A2(n1250), .A3(n1183), .A4(n1061), .ZN(n1248) );
NOR3_X1 U890 ( .A1(n1251), .A2(n1068), .A3(n1252), .ZN(n1061) );
NOR3_X1 U891 ( .A1(n1251), .A2(n1068), .A3(n1072), .ZN(n1183) );
INV_X1 U892 ( .A(n1253), .ZN(n1251) );
NOR2_X1 U893 ( .A1(n1254), .A2(n1255), .ZN(n1247) );
AND3_X1 U894 ( .A1(n1105), .A2(n1253), .A3(n1103), .ZN(n1255) );
NOR3_X1 U895 ( .A1(n1256), .A2(n1257), .A3(n1072), .ZN(n1254) );
NAND2_X1 U896 ( .A1(n1258), .A2(KEYINPUT51), .ZN(n1226) );
XOR2_X1 U897 ( .A(n1259), .B(n1260), .Z(n1258) );
AND2_X1 U898 ( .A1(n1261), .A2(n1107), .ZN(n1163) );
INV_X1 U899 ( .A(G952), .ZN(n1107) );
XOR2_X1 U900 ( .A(n1101), .B(KEYINPUT22), .Z(n1261) );
XOR2_X1 U901 ( .A(n1262), .B(n1263), .Z(G48) );
NAND3_X1 U902 ( .A1(n1239), .A2(n1237), .A3(n1264), .ZN(n1263) );
XOR2_X1 U903 ( .A(n1089), .B(KEYINPUT25), .Z(n1264) );
XNOR2_X1 U904 ( .A(G143), .B(n1265), .ZN(G45) );
NOR2_X1 U905 ( .A1(n1234), .A2(KEYINPUT1), .ZN(n1265) );
AND4_X1 U906 ( .A1(n1266), .A2(n1095), .A3(n1106), .A4(n1267), .ZN(n1234) );
NOR3_X1 U907 ( .A1(n1089), .A2(n1268), .A3(n1269), .ZN(n1267) );
XOR2_X1 U908 ( .A(n1150), .B(n1270), .Z(G42) );
NAND4_X1 U909 ( .A1(KEYINPUT36), .A2(n1271), .A3(n1105), .A4(n1237), .ZN(n1270) );
INV_X1 U910 ( .A(G140), .ZN(n1150) );
XOR2_X1 U911 ( .A(G137), .B(n1233), .Z(G39) );
AND3_X1 U912 ( .A1(n1076), .A2(n1103), .A3(n1239), .ZN(n1233) );
XOR2_X1 U913 ( .A(n1272), .B(n1273), .Z(G36) );
XOR2_X1 U914 ( .A(KEYINPUT9), .B(G134), .Z(n1273) );
NAND4_X1 U915 ( .A1(KEYINPUT32), .A2(n1271), .A3(n1106), .A4(n1099), .ZN(n1272) );
XNOR2_X1 U916 ( .A(G131), .B(n1229), .ZN(G33) );
NAND3_X1 U917 ( .A1(n1237), .A2(n1106), .A3(n1271), .ZN(n1229) );
NOR3_X1 U918 ( .A1(n1274), .A2(n1268), .A3(n1093), .ZN(n1271) );
INV_X1 U919 ( .A(n1076), .ZN(n1093) );
NOR2_X1 U920 ( .A1(n1090), .A2(n1275), .ZN(n1076) );
INV_X1 U921 ( .A(n1091), .ZN(n1275) );
XOR2_X1 U922 ( .A(n1276), .B(G128), .Z(G30) );
NAND2_X1 U923 ( .A1(KEYINPUT8), .A2(n1236), .ZN(n1276) );
NAND3_X1 U924 ( .A1(n1099), .A2(n1238), .A3(n1239), .ZN(n1236) );
NOR4_X1 U925 ( .A1(n1274), .A2(n1277), .A3(n1113), .A4(n1268), .ZN(n1239) );
NAND2_X1 U926 ( .A1(n1278), .A2(n1279), .ZN(G3) );
NAND2_X1 U927 ( .A1(n1250), .A2(n1192), .ZN(n1279) );
XOR2_X1 U928 ( .A(KEYINPUT40), .B(n1280), .Z(n1278) );
NOR2_X1 U929 ( .A1(n1250), .A2(n1192), .ZN(n1280) );
INV_X1 U930 ( .A(G101), .ZN(n1192) );
AND3_X1 U931 ( .A1(n1106), .A2(n1253), .A3(n1103), .ZN(n1250) );
NOR3_X1 U932 ( .A1(n1274), .A2(n1281), .A3(n1257), .ZN(n1253) );
NAND2_X1 U933 ( .A1(n1282), .A2(n1283), .ZN(G27) );
NAND2_X1 U934 ( .A1(n1232), .A2(n1284), .ZN(n1283) );
NAND2_X1 U935 ( .A1(G125), .A2(n1285), .ZN(n1284) );
OR2_X1 U936 ( .A1(KEYINPUT52), .A2(KEYINPUT53), .ZN(n1285) );
INV_X1 U937 ( .A(n1286), .ZN(n1232) );
NAND3_X1 U938 ( .A1(n1287), .A2(n1288), .A3(KEYINPUT53), .ZN(n1282) );
NAND2_X1 U939 ( .A1(n1152), .A2(n1289), .ZN(n1288) );
NAND2_X1 U940 ( .A1(G125), .A2(n1290), .ZN(n1287) );
NAND2_X1 U941 ( .A1(n1286), .A2(n1289), .ZN(n1290) );
INV_X1 U942 ( .A(KEYINPUT52), .ZN(n1289) );
NAND4_X1 U943 ( .A1(n1105), .A2(n1237), .A3(n1291), .A4(n1078), .ZN(n1286) );
NOR2_X1 U944 ( .A1(n1268), .A2(n1089), .ZN(n1291) );
INV_X1 U945 ( .A(n1244), .ZN(n1268) );
NAND2_X1 U946 ( .A1(n1077), .A2(n1292), .ZN(n1244) );
NAND4_X1 U947 ( .A1(G953), .A2(G902), .A3(n1293), .A4(n1141), .ZN(n1292) );
INV_X1 U948 ( .A(G900), .ZN(n1141) );
XOR2_X1 U949 ( .A(G122), .B(n1249), .Z(G24) );
NOR4_X1 U950 ( .A1(n1086), .A2(n1068), .A3(n1294), .A4(n1295), .ZN(n1249) );
NAND3_X1 U951 ( .A1(n1238), .A2(n1296), .A3(n1115), .ZN(n1295) );
NAND2_X1 U952 ( .A1(n1113), .A2(n1277), .ZN(n1068) );
XOR2_X1 U953 ( .A(n1245), .B(n1297), .Z(G21) );
XOR2_X1 U954 ( .A(KEYINPUT28), .B(G119), .Z(n1297) );
NAND4_X1 U955 ( .A1(n1298), .A2(n1296), .A3(n1299), .A4(n1300), .ZN(n1245) );
NOR3_X1 U956 ( .A1(n1082), .A2(n1089), .A3(n1086), .ZN(n1300) );
INV_X1 U957 ( .A(n1078), .ZN(n1086) );
XNOR2_X1 U958 ( .A(G116), .B(n1246), .ZN(G18) );
NAND3_X1 U959 ( .A1(n1099), .A2(n1238), .A3(n1301), .ZN(n1246) );
INV_X1 U960 ( .A(n1089), .ZN(n1238) );
XOR2_X1 U961 ( .A(n1257), .B(KEYINPUT57), .Z(n1089) );
INV_X1 U962 ( .A(n1252), .ZN(n1099) );
NAND2_X1 U963 ( .A1(n1115), .A2(n1294), .ZN(n1252) );
INV_X1 U964 ( .A(n1269), .ZN(n1115) );
XNOR2_X1 U965 ( .A(G113), .B(n1302), .ZN(G15) );
NAND3_X1 U966 ( .A1(n1301), .A2(n1237), .A3(n1303), .ZN(n1302) );
XOR2_X1 U967 ( .A(n1257), .B(KEYINPUT41), .Z(n1303) );
INV_X1 U968 ( .A(n1072), .ZN(n1237) );
NAND2_X1 U969 ( .A1(n1266), .A2(n1269), .ZN(n1072) );
INV_X1 U970 ( .A(n1256), .ZN(n1301) );
NAND3_X1 U971 ( .A1(n1078), .A2(n1296), .A3(n1106), .ZN(n1256) );
NOR2_X1 U972 ( .A1(n1299), .A2(n1113), .ZN(n1106) );
NOR2_X1 U973 ( .A1(n1096), .A2(n1304), .ZN(n1078) );
NOR2_X1 U974 ( .A1(n1098), .A2(n1097), .ZN(n1304) );
INV_X1 U975 ( .A(n1305), .ZN(n1097) );
XNOR2_X1 U976 ( .A(G110), .B(n1306), .ZN(G12) );
NAND4_X1 U977 ( .A1(n1105), .A2(n1103), .A3(n1307), .A4(n1095), .ZN(n1306) );
INV_X1 U978 ( .A(n1274), .ZN(n1095) );
NAND2_X1 U979 ( .A1(n1096), .A2(n1308), .ZN(n1274) );
NAND2_X1 U980 ( .A1(G221), .A2(n1305), .ZN(n1308) );
XNOR2_X1 U981 ( .A(n1309), .B(G469), .ZN(n1096) );
NAND2_X1 U982 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U983 ( .A(n1312), .B(n1313), .Z(n1310) );
XOR2_X1 U984 ( .A(n1210), .B(n1216), .Z(n1313) );
INV_X1 U985 ( .A(n1223), .ZN(n1216) );
NAND2_X1 U986 ( .A1(n1314), .A2(n1315), .ZN(n1223) );
NAND2_X1 U987 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
INV_X1 U988 ( .A(G107), .ZN(n1317) );
XOR2_X1 U989 ( .A(KEYINPUT16), .B(n1318), .Z(n1316) );
NAND2_X1 U990 ( .A1(n1318), .A2(G107), .ZN(n1314) );
XOR2_X1 U991 ( .A(G104), .B(n1319), .Z(n1318) );
XNOR2_X1 U992 ( .A(n1320), .B(n1321), .ZN(n1210) );
XOR2_X1 U993 ( .A(G140), .B(G110), .Z(n1321) );
NAND2_X1 U994 ( .A1(G227), .A2(n1101), .ZN(n1320) );
XOR2_X1 U995 ( .A(KEYINPUT18), .B(n1322), .Z(n1312) );
INV_X1 U996 ( .A(n1142), .ZN(n1322) );
XNOR2_X1 U997 ( .A(n1222), .B(n1323), .ZN(n1142) );
XNOR2_X1 U998 ( .A(n1324), .B(KEYINPUT0), .ZN(n1222) );
NOR2_X1 U999 ( .A1(n1281), .A2(n1325), .ZN(n1307) );
XOR2_X1 U1000 ( .A(n1257), .B(KEYINPUT23), .Z(n1325) );
NAND2_X1 U1001 ( .A1(n1090), .A2(n1091), .ZN(n1257) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1326), .ZN(n1091) );
XOR2_X1 U1003 ( .A(n1129), .B(n1327), .Z(n1090) );
NOR2_X1 U1004 ( .A1(n1131), .A2(KEYINPUT35), .ZN(n1327) );
AND2_X1 U1005 ( .A1(n1328), .A2(n1311), .ZN(n1131) );
XOR2_X1 U1006 ( .A(n1329), .B(n1330), .Z(n1328) );
INV_X1 U1007 ( .A(n1259), .ZN(n1330) );
XNOR2_X1 U1008 ( .A(n1159), .B(n1331), .ZN(n1259) );
XOR2_X1 U1009 ( .A(G125), .B(n1332), .Z(n1331) );
AND2_X1 U1010 ( .A1(n1101), .A2(G224), .ZN(n1332) );
XOR2_X1 U1011 ( .A(n1333), .B(n1334), .Z(n1159) );
XOR2_X1 U1012 ( .A(n1335), .B(n1336), .Z(n1333) );
XOR2_X1 U1013 ( .A(n1337), .B(n1338), .Z(n1336) );
XOR2_X1 U1014 ( .A(G116), .B(G107), .Z(n1338) );
XOR2_X1 U1015 ( .A(KEYINPUT47), .B(G122), .Z(n1337) );
XOR2_X1 U1016 ( .A(n1339), .B(n1340), .Z(n1335) );
XOR2_X1 U1017 ( .A(n1341), .B(n1319), .Z(n1340) );
XOR2_X1 U1018 ( .A(G101), .B(KEYINPUT31), .Z(n1319) );
NOR2_X1 U1019 ( .A1(G110), .A2(KEYINPUT30), .ZN(n1341) );
XOR2_X1 U1020 ( .A(n1342), .B(G104), .Z(n1339) );
NAND2_X1 U1021 ( .A1(KEYINPUT48), .A2(n1343), .ZN(n1342) );
NOR2_X1 U1022 ( .A1(KEYINPUT45), .A2(n1260), .ZN(n1329) );
XNOR2_X1 U1023 ( .A(n1221), .B(n1344), .ZN(n1260) );
NAND2_X1 U1024 ( .A1(G210), .A2(n1326), .ZN(n1129) );
NAND2_X1 U1025 ( .A1(n1345), .A2(n1311), .ZN(n1326) );
INV_X1 U1026 ( .A(n1296), .ZN(n1281) );
NAND2_X1 U1027 ( .A1(n1346), .A2(n1077), .ZN(n1296) );
NAND3_X1 U1028 ( .A1(n1293), .A2(n1101), .A3(n1347), .ZN(n1077) );
XOR2_X1 U1029 ( .A(KEYINPUT43), .B(G952), .Z(n1347) );
NAND4_X1 U1030 ( .A1(G953), .A2(G902), .A3(n1293), .A4(n1161), .ZN(n1346) );
INV_X1 U1031 ( .A(G898), .ZN(n1161) );
NAND2_X1 U1032 ( .A1(G234), .A2(G237), .ZN(n1293) );
INV_X1 U1033 ( .A(n1082), .ZN(n1103) );
NAND2_X1 U1034 ( .A1(n1269), .A2(n1294), .ZN(n1082) );
INV_X1 U1035 ( .A(n1266), .ZN(n1294) );
XOR2_X1 U1036 ( .A(n1348), .B(n1177), .Z(n1266) );
INV_X1 U1037 ( .A(n1124), .ZN(n1177) );
NAND2_X1 U1038 ( .A1(n1180), .A2(n1311), .ZN(n1124) );
XOR2_X1 U1039 ( .A(n1349), .B(n1350), .Z(n1180) );
XOR2_X1 U1040 ( .A(n1351), .B(n1352), .Z(n1350) );
NAND2_X1 U1041 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1042 ( .A(n1355), .B(n1356), .Z(n1354) );
XOR2_X1 U1043 ( .A(n1357), .B(n1358), .Z(n1356) );
NOR2_X1 U1044 ( .A1(G143), .A2(KEYINPUT62), .ZN(n1358) );
XNOR2_X1 U1045 ( .A(G131), .B(n1359), .ZN(n1355) );
AND2_X1 U1046 ( .A1(n1360), .A2(G214), .ZN(n1359) );
XNOR2_X1 U1047 ( .A(KEYINPUT46), .B(KEYINPUT33), .ZN(n1353) );
INV_X1 U1048 ( .A(G104), .ZN(n1351) );
XNOR2_X1 U1049 ( .A(G113), .B(n1361), .ZN(n1349) );
XOR2_X1 U1050 ( .A(KEYINPUT10), .B(G122), .Z(n1361) );
NAND2_X1 U1051 ( .A1(KEYINPUT38), .A2(n1126), .ZN(n1348) );
INV_X1 U1052 ( .A(G475), .ZN(n1126) );
XOR2_X1 U1053 ( .A(n1362), .B(G478), .Z(n1269) );
NAND2_X1 U1054 ( .A1(n1173), .A2(n1311), .ZN(n1362) );
XNOR2_X1 U1055 ( .A(n1363), .B(n1364), .ZN(n1173) );
XOR2_X1 U1056 ( .A(G128), .B(n1365), .Z(n1364) );
XOR2_X1 U1057 ( .A(G143), .B(G134), .Z(n1365) );
XOR2_X1 U1058 ( .A(n1366), .B(n1367), .Z(n1363) );
NOR2_X1 U1059 ( .A1(KEYINPUT37), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1060 ( .A(n1369), .B(n1370), .Z(n1368) );
XOR2_X1 U1061 ( .A(G122), .B(G107), .Z(n1370) );
NAND2_X1 U1062 ( .A1(KEYINPUT55), .A2(G116), .ZN(n1369) );
NAND3_X1 U1063 ( .A1(G217), .A2(n1101), .A3(G234), .ZN(n1366) );
NOR2_X1 U1064 ( .A1(n1298), .A2(n1277), .ZN(n1105) );
INV_X1 U1065 ( .A(n1299), .ZN(n1277) );
XOR2_X1 U1066 ( .A(n1122), .B(n1118), .Z(n1299) );
INV_X1 U1067 ( .A(n1123), .ZN(n1118) );
NAND2_X1 U1068 ( .A1(G217), .A2(n1305), .ZN(n1123) );
NAND2_X1 U1069 ( .A1(n1371), .A2(G234), .ZN(n1305) );
XOR2_X1 U1070 ( .A(n1311), .B(KEYINPUT6), .Z(n1371) );
NOR2_X1 U1071 ( .A1(n1169), .A2(G902), .ZN(n1122) );
XOR2_X1 U1072 ( .A(n1372), .B(n1373), .Z(n1169) );
XOR2_X1 U1073 ( .A(n1374), .B(n1375), .Z(n1373) );
INV_X1 U1074 ( .A(n1357), .ZN(n1375) );
XOR2_X1 U1075 ( .A(n1152), .B(n1376), .Z(n1357) );
XOR2_X1 U1076 ( .A(G146), .B(G140), .Z(n1376) );
INV_X1 U1077 ( .A(G125), .ZN(n1152) );
NOR3_X1 U1078 ( .A1(n1377), .A2(G953), .A3(n1098), .ZN(n1374) );
INV_X1 U1079 ( .A(G221), .ZN(n1098) );
XOR2_X1 U1080 ( .A(KEYINPUT42), .B(G234), .Z(n1377) );
XOR2_X1 U1081 ( .A(n1378), .B(n1379), .Z(n1372) );
NOR2_X1 U1082 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
XOR2_X1 U1083 ( .A(KEYINPUT7), .B(n1382), .Z(n1381) );
NOR2_X1 U1084 ( .A1(G110), .A2(n1383), .ZN(n1382) );
AND2_X1 U1085 ( .A1(n1383), .A2(G110), .ZN(n1380) );
XNOR2_X1 U1086 ( .A(n1343), .B(G128), .ZN(n1383) );
INV_X1 U1087 ( .A(G119), .ZN(n1343) );
XOR2_X1 U1088 ( .A(n1384), .B(KEYINPUT17), .Z(n1378) );
INV_X1 U1089 ( .A(G137), .ZN(n1384) );
INV_X1 U1090 ( .A(n1113), .ZN(n1298) );
XOR2_X1 U1091 ( .A(n1385), .B(G472), .Z(n1113) );
NAND2_X1 U1092 ( .A1(n1386), .A2(n1311), .ZN(n1385) );
INV_X1 U1093 ( .A(G902), .ZN(n1311) );
XOR2_X1 U1094 ( .A(n1387), .B(n1388), .Z(n1386) );
XOR2_X1 U1095 ( .A(G101), .B(n1389), .Z(n1388) );
NOR2_X1 U1096 ( .A1(KEYINPUT56), .A2(n1390), .ZN(n1389) );
INV_X1 U1097 ( .A(n1196), .ZN(n1390) );
XOR2_X1 U1098 ( .A(n1391), .B(n1392), .Z(n1196) );
XOR2_X1 U1099 ( .A(KEYINPUT34), .B(G119), .Z(n1392) );
XNOR2_X1 U1100 ( .A(G116), .B(n1393), .ZN(n1391) );
NOR2_X1 U1101 ( .A1(KEYINPUT11), .A2(n1334), .ZN(n1393) );
XNOR2_X1 U1102 ( .A(G113), .B(KEYINPUT19), .ZN(n1334) );
XNOR2_X1 U1103 ( .A(n1188), .B(n1191), .ZN(n1387) );
NAND2_X1 U1104 ( .A1(G210), .A2(n1360), .ZN(n1191) );
AND2_X1 U1105 ( .A1(n1394), .A2(n1101), .ZN(n1360) );
INV_X1 U1106 ( .A(G953), .ZN(n1101) );
XOR2_X1 U1107 ( .A(n1345), .B(KEYINPUT12), .Z(n1394) );
INV_X1 U1108 ( .A(G237), .ZN(n1345) );
XNOR2_X1 U1109 ( .A(n1344), .B(n1323), .ZN(n1188) );
XNOR2_X1 U1110 ( .A(n1221), .B(n1212), .ZN(n1323) );
XNOR2_X1 U1111 ( .A(n1395), .B(n1396), .ZN(n1212) );
XOR2_X1 U1112 ( .A(KEYINPUT49), .B(G137), .Z(n1396) );
XNOR2_X1 U1113 ( .A(G131), .B(G134), .ZN(n1395) );
XOR2_X1 U1114 ( .A(n1262), .B(G143), .Z(n1221) );
INV_X1 U1115 ( .A(G146), .ZN(n1262) );
NOR2_X1 U1116 ( .A1(KEYINPUT59), .A2(n1324), .ZN(n1344) );
XNOR2_X1 U1117 ( .A(G128), .B(KEYINPUT13), .ZN(n1324) );
endmodule


