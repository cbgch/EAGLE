//Key = 1111100101011010011001001111010111100110010100101100100110010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328;

XNOR2_X1 U731 ( .A(G107), .B(n1015), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U733 ( .A1(G953), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1017) );
XOR2_X1 U734 ( .A(KEYINPUT0), .B(n1021), .Z(n1020) );
NOR2_X1 U735 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR3_X1 U736 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NOR4_X1 U737 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
NOR2_X1 U738 ( .A1(n1031), .A2(KEYINPUT59), .ZN(n1030) );
NOR3_X1 U739 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NOR2_X1 U740 ( .A1(n1035), .A2(n1036), .ZN(n1029) );
NOR2_X1 U741 ( .A1(n1037), .A2(n1036), .ZN(n1028) );
NOR3_X1 U742 ( .A1(n1032), .A2(n1038), .A3(n1033), .ZN(n1027) );
NOR2_X1 U743 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
AND2_X1 U745 ( .A1(n1043), .A2(KEYINPUT59), .ZN(n1039) );
NOR3_X1 U746 ( .A1(n1033), .A2(n1044), .A3(n1045), .ZN(n1022) );
NOR3_X1 U747 ( .A1(n1025), .A2(n1046), .A3(n1047), .ZN(n1045) );
NOR2_X1 U748 ( .A1(n1048), .A2(n1036), .ZN(n1047) );
NOR2_X1 U749 ( .A1(KEYINPUT45), .A2(n1024), .ZN(n1048) );
NOR3_X1 U750 ( .A1(n1032), .A2(n1049), .A3(n1024), .ZN(n1046) );
NOR2_X1 U751 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
AND2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR3_X1 U753 ( .A1(n1042), .A2(n1054), .A3(n1055), .ZN(n1050) );
INV_X1 U754 ( .A(n1056), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1057), .A2(n1058), .ZN(n1044) );
NOR3_X1 U756 ( .A1(n1036), .A2(KEYINPUT45), .A3(n1024), .ZN(n1057) );
NAND3_X1 U757 ( .A1(n1053), .A2(n1056), .A3(n1059), .ZN(n1036) );
INV_X1 U758 ( .A(n1032), .ZN(n1059) );
NOR3_X1 U759 ( .A1(n1018), .A2(G953), .A3(G952), .ZN(n1016) );
AND4_X1 U760 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1018) );
NOR4_X1 U761 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
XNOR2_X1 U762 ( .A(G472), .B(n1068), .ZN(n1067) );
NAND2_X1 U763 ( .A1(KEYINPUT33), .A2(n1069), .ZN(n1068) );
XOR2_X1 U764 ( .A(n1070), .B(n1071), .Z(n1066) );
XNOR2_X1 U765 ( .A(KEYINPUT16), .B(n1072), .ZN(n1071) );
NOR2_X1 U766 ( .A1(KEYINPUT63), .A2(n1073), .ZN(n1070) );
XOR2_X1 U767 ( .A(KEYINPUT30), .B(n1074), .Z(n1065) );
NOR2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XNOR2_X1 U769 ( .A(n1077), .B(KEYINPUT40), .ZN(n1076) );
XNOR2_X1 U770 ( .A(n1078), .B(n1079), .ZN(n1064) );
XOR2_X1 U771 ( .A(KEYINPUT61), .B(KEYINPUT35), .Z(n1079) );
NOR3_X1 U772 ( .A1(n1080), .A2(n1081), .A3(n1025), .ZN(n1062) );
INV_X1 U773 ( .A(n1058), .ZN(n1025) );
INV_X1 U774 ( .A(n1055), .ZN(n1081) );
AND2_X1 U775 ( .A1(n1082), .A2(n1075), .ZN(n1080) );
XNOR2_X1 U776 ( .A(n1083), .B(n1084), .ZN(n1060) );
XNOR2_X1 U777 ( .A(KEYINPUT10), .B(n1085), .ZN(n1084) );
XOR2_X1 U778 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1088) );
NOR2_X1 U781 ( .A1(KEYINPUT28), .A2(n1090), .ZN(n1086) );
NOR2_X1 U782 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U784 ( .A1(n1089), .A2(n1095), .ZN(n1094) );
NAND2_X1 U785 ( .A1(KEYINPUT1), .A2(n1096), .ZN(n1093) );
NOR2_X1 U786 ( .A1(KEYINPUT1), .A2(n1096), .ZN(n1091) );
AND2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U789 ( .A(n1101), .B(n1102), .ZN(n1097) );
XNOR2_X1 U790 ( .A(n1103), .B(n1104), .ZN(n1102) );
NOR2_X1 U791 ( .A1(KEYINPUT6), .A2(n1105), .ZN(n1104) );
XOR2_X1 U792 ( .A(n1106), .B(n1107), .Z(n1105) );
XNOR2_X1 U793 ( .A(n1108), .B(n1109), .ZN(n1107) );
XNOR2_X1 U794 ( .A(G134), .B(KEYINPUT13), .ZN(n1106) );
NAND2_X1 U795 ( .A1(KEYINPUT9), .A2(n1110), .ZN(n1103) );
INV_X1 U796 ( .A(G140), .ZN(n1110) );
NAND3_X1 U797 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(G69) );
NAND2_X1 U798 ( .A1(n1114), .A2(n1089), .ZN(n1113) );
XNOR2_X1 U799 ( .A(n1115), .B(n1116), .ZN(n1114) );
NAND4_X1 U800 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1115) );
XOR2_X1 U801 ( .A(KEYINPUT22), .B(n1121), .Z(n1118) );
XOR2_X1 U802 ( .A(n1015), .B(KEYINPUT50), .Z(n1117) );
NAND3_X1 U803 ( .A1(G953), .A2(n1122), .A3(n1116), .ZN(n1112) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1122) );
NAND4_X1 U805 ( .A1(G224), .A2(G953), .A3(G898), .A4(n1123), .ZN(n1111) );
INV_X1 U806 ( .A(n1116), .ZN(n1123) );
NAND3_X1 U807 ( .A1(KEYINPUT2), .A2(n1124), .A3(n1125), .ZN(n1116) );
XNOR2_X1 U808 ( .A(n1126), .B(KEYINPUT60), .ZN(n1125) );
NOR3_X1 U809 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1130), .A2(n1131), .A3(n1089), .ZN(n1129) );
INV_X1 U811 ( .A(KEYINPUT51), .ZN(n1130) );
NOR2_X1 U812 ( .A1(KEYINPUT51), .A2(n1132), .ZN(n1128) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1127) );
NOR2_X1 U814 ( .A1(n1082), .A2(n1135), .ZN(n1133) );
NOR2_X1 U815 ( .A1(n1136), .A2(n1137), .ZN(G63) );
XOR2_X1 U816 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1135), .ZN(n1138) );
NOR2_X1 U818 ( .A1(n1136), .A2(n1141), .ZN(G60) );
NOR3_X1 U819 ( .A1(n1083), .A2(n1142), .A3(n1143), .ZN(n1141) );
NOR3_X1 U820 ( .A1(n1144), .A2(n1085), .A3(n1135), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
AND2_X1 U822 ( .A1(n1019), .A2(G475), .ZN(n1145) );
XNOR2_X1 U823 ( .A(G104), .B(n1120), .ZN(G6) );
NOR2_X1 U824 ( .A1(n1136), .A2(n1147), .ZN(G57) );
NOR2_X1 U825 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U826 ( .A(n1150), .B(KEYINPUT32), .Z(n1149) );
NAND2_X1 U827 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U828 ( .A1(n1151), .A2(n1152), .ZN(n1148) );
NAND2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U830 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
INV_X1 U831 ( .A(n1157), .ZN(n1156) );
XNOR2_X1 U832 ( .A(n1158), .B(KEYINPUT15), .ZN(n1155) );
NAND2_X1 U833 ( .A1(n1159), .A2(n1157), .ZN(n1153) );
XNOR2_X1 U834 ( .A(KEYINPUT57), .B(n1160), .ZN(n1159) );
INV_X1 U835 ( .A(n1158), .ZN(n1160) );
XOR2_X1 U836 ( .A(n1161), .B(n1162), .Z(n1158) );
XOR2_X1 U837 ( .A(n1163), .B(n1164), .Z(n1161) );
NOR2_X1 U838 ( .A1(n1165), .A2(n1135), .ZN(n1164) );
NOR2_X1 U839 ( .A1(n1136), .A2(n1166), .ZN(G54) );
XOR2_X1 U840 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U841 ( .A1(n1072), .A2(n1135), .ZN(n1168) );
NAND2_X1 U842 ( .A1(KEYINPUT37), .A2(n1169), .ZN(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U844 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U845 ( .A(n1174), .B(n1175), .Z(n1170) );
XNOR2_X1 U846 ( .A(n1176), .B(n1177), .ZN(n1175) );
NOR2_X1 U847 ( .A1(G140), .A2(KEYINPUT44), .ZN(n1177) );
NAND2_X1 U848 ( .A1(KEYINPUT21), .A2(n1178), .ZN(n1174) );
INV_X1 U849 ( .A(n1179), .ZN(n1178) );
NOR2_X1 U850 ( .A1(n1136), .A2(n1180), .ZN(G51) );
XOR2_X1 U851 ( .A(n1181), .B(n1182), .Z(n1180) );
XNOR2_X1 U852 ( .A(n1183), .B(n1184), .ZN(n1182) );
NAND2_X1 U853 ( .A1(KEYINPUT49), .A2(n1185), .ZN(n1183) );
INV_X1 U854 ( .A(n1124), .ZN(n1185) );
XOR2_X1 U855 ( .A(n1186), .B(n1187), .Z(n1181) );
NOR2_X1 U856 ( .A1(KEYINPUT53), .A2(n1101), .ZN(n1187) );
NOR2_X1 U857 ( .A1(n1188), .A2(n1135), .ZN(n1186) );
NAND2_X1 U858 ( .A1(G902), .A2(n1019), .ZN(n1135) );
NAND3_X1 U859 ( .A1(n1189), .A2(n1121), .A3(n1190), .ZN(n1019) );
AND3_X1 U860 ( .A1(n1119), .A2(n1120), .A3(n1015), .ZN(n1190) );
NAND3_X1 U861 ( .A1(n1052), .A2(n1191), .A3(n1192), .ZN(n1015) );
NAND3_X1 U862 ( .A1(n1192), .A2(n1191), .A3(n1193), .ZN(n1120) );
NAND3_X1 U863 ( .A1(n1194), .A2(n1195), .A3(n1056), .ZN(n1119) );
NAND2_X1 U864 ( .A1(n1192), .A2(n1196), .ZN(n1195) );
NAND2_X1 U865 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND2_X1 U866 ( .A1(n1035), .A2(n1199), .ZN(n1198) );
NAND2_X1 U867 ( .A1(KEYINPUT7), .A2(n1200), .ZN(n1199) );
INV_X1 U868 ( .A(n1201), .ZN(n1035) );
NAND2_X1 U869 ( .A1(n1202), .A2(n1041), .ZN(n1194) );
NAND2_X1 U870 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
INV_X1 U871 ( .A(KEYINPUT7), .ZN(n1204) );
AND4_X1 U872 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1121) );
NAND4_X1 U873 ( .A1(n1209), .A2(n1053), .A3(n1191), .A4(n1210), .ZN(n1205) );
INV_X1 U874 ( .A(n1095), .ZN(n1189) );
NAND4_X1 U875 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1095) );
NOR4_X1 U876 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NAND2_X1 U877 ( .A1(n1052), .A2(n1219), .ZN(n1213) );
NAND2_X1 U878 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND2_X1 U879 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XNOR2_X1 U880 ( .A(n1200), .B(KEYINPUT46), .ZN(n1222) );
NAND2_X1 U881 ( .A1(n1224), .A2(n1225), .ZN(n1220) );
INV_X1 U882 ( .A(n1132), .ZN(n1136) );
NAND2_X1 U883 ( .A1(n1131), .A2(G953), .ZN(n1132) );
XNOR2_X1 U884 ( .A(G952), .B(KEYINPUT20), .ZN(n1131) );
XNOR2_X1 U885 ( .A(G146), .B(n1211), .ZN(G48) );
NAND3_X1 U886 ( .A1(n1225), .A2(n1193), .A3(n1224), .ZN(n1211) );
XNOR2_X1 U887 ( .A(G143), .B(n1212), .ZN(G45) );
NAND4_X1 U888 ( .A1(n1224), .A2(n1200), .A3(n1209), .A4(n1210), .ZN(n1212) );
XOR2_X1 U889 ( .A(n1226), .B(n1218), .Z(G42) );
AND3_X1 U890 ( .A1(n1201), .A2(n1193), .A3(n1223), .ZN(n1218) );
XNOR2_X1 U891 ( .A(G140), .B(KEYINPUT17), .ZN(n1226) );
XOR2_X1 U892 ( .A(G137), .B(n1217), .Z(G39) );
AND3_X1 U893 ( .A1(n1223), .A2(n1056), .A3(n1225), .ZN(n1217) );
NAND2_X1 U894 ( .A1(n1227), .A2(n1228), .ZN(G36) );
NAND2_X1 U895 ( .A1(G134), .A2(n1229), .ZN(n1228) );
XOR2_X1 U896 ( .A(KEYINPUT27), .B(n1230), .Z(n1227) );
NOR2_X1 U897 ( .A1(G134), .A2(n1229), .ZN(n1230) );
NAND3_X1 U898 ( .A1(n1200), .A2(n1052), .A3(n1223), .ZN(n1229) );
XOR2_X1 U899 ( .A(G131), .B(n1216), .Z(G33) );
AND3_X1 U900 ( .A1(n1200), .A2(n1193), .A3(n1223), .ZN(n1216) );
AND4_X1 U901 ( .A1(n1061), .A2(n1192), .A3(n1231), .A4(n1058), .ZN(n1223) );
INV_X1 U902 ( .A(n1024), .ZN(n1061) );
INV_X1 U903 ( .A(n1037), .ZN(n1200) );
XNOR2_X1 U904 ( .A(G128), .B(n1232), .ZN(G30) );
NAND4_X1 U905 ( .A1(n1225), .A2(n1052), .A3(n1233), .A4(n1234), .ZN(n1232) );
OR2_X1 U906 ( .A1(n1224), .A2(KEYINPUT39), .ZN(n1234) );
AND2_X1 U907 ( .A1(n1235), .A2(n1192), .ZN(n1224) );
NAND2_X1 U908 ( .A1(KEYINPUT39), .A2(n1236), .ZN(n1233) );
NAND2_X1 U909 ( .A1(n1235), .A2(n1041), .ZN(n1236) );
INV_X1 U910 ( .A(n1192), .ZN(n1041) );
XNOR2_X1 U911 ( .A(G101), .B(n1237), .ZN(G3) );
NAND3_X1 U912 ( .A1(n1203), .A2(n1192), .A3(n1056), .ZN(n1237) );
XNOR2_X1 U913 ( .A(G125), .B(n1238), .ZN(G27) );
NAND2_X1 U914 ( .A1(KEYINPUT38), .A2(n1215), .ZN(n1238) );
AND3_X1 U915 ( .A1(n1235), .A2(n1043), .A3(n1201), .ZN(n1215) );
AND3_X1 U916 ( .A1(n1231), .A2(n1058), .A3(n1024), .ZN(n1235) );
NAND2_X1 U917 ( .A1(n1032), .A2(n1239), .ZN(n1231) );
NAND4_X1 U918 ( .A1(n1099), .A2(G902), .A3(n1240), .A4(n1100), .ZN(n1239) );
INV_X1 U919 ( .A(G900), .ZN(n1100) );
INV_X1 U920 ( .A(n1241), .ZN(n1099) );
XNOR2_X1 U921 ( .A(G122), .B(n1242), .ZN(G24) );
NAND4_X1 U922 ( .A1(n1209), .A2(n1191), .A3(n1243), .A4(n1210), .ZN(n1242) );
XOR2_X1 U923 ( .A(KEYINPUT36), .B(n1053), .Z(n1243) );
NOR2_X1 U924 ( .A1(n1244), .A2(n1033), .ZN(n1191) );
NAND2_X1 U925 ( .A1(n1245), .A2(n1246), .ZN(n1033) );
XNOR2_X1 U926 ( .A(G119), .B(n1206), .ZN(G21) );
NAND4_X1 U927 ( .A1(n1225), .A2(n1053), .A3(n1056), .A4(n1197), .ZN(n1206) );
NOR2_X1 U928 ( .A1(n1246), .A2(n1245), .ZN(n1225) );
INV_X1 U929 ( .A(n1247), .ZN(n1245) );
XNOR2_X1 U930 ( .A(G116), .B(n1207), .ZN(G18) );
NAND3_X1 U931 ( .A1(n1203), .A2(n1052), .A3(n1053), .ZN(n1207) );
NOR2_X1 U932 ( .A1(n1078), .A2(n1209), .ZN(n1052) );
XNOR2_X1 U933 ( .A(G113), .B(n1208), .ZN(G15) );
NAND2_X1 U934 ( .A1(n1043), .A2(n1203), .ZN(n1208) );
NOR2_X1 U935 ( .A1(n1037), .A2(n1244), .ZN(n1203) );
NAND2_X1 U936 ( .A1(n1246), .A2(n1247), .ZN(n1037) );
INV_X1 U937 ( .A(n1034), .ZN(n1043) );
NAND2_X1 U938 ( .A1(n1053), .A2(n1193), .ZN(n1034) );
AND2_X1 U939 ( .A1(n1209), .A2(n1078), .ZN(n1193) );
INV_X1 U940 ( .A(n1210), .ZN(n1078) );
NOR2_X1 U941 ( .A1(n1248), .A2(n1054), .ZN(n1053) );
XNOR2_X1 U942 ( .A(G110), .B(n1249), .ZN(G12) );
NAND4_X1 U943 ( .A1(n1250), .A2(n1201), .A3(n1056), .A4(n1197), .ZN(n1249) );
INV_X1 U944 ( .A(n1244), .ZN(n1197) );
NAND3_X1 U945 ( .A1(n1251), .A2(n1058), .A3(n1024), .ZN(n1244) );
XOR2_X1 U946 ( .A(n1252), .B(n1188), .Z(n1024) );
NAND2_X1 U947 ( .A1(G210), .A2(n1253), .ZN(n1188) );
NAND2_X1 U948 ( .A1(n1254), .A2(n1255), .ZN(n1252) );
XNOR2_X1 U949 ( .A(n1256), .B(n1257), .ZN(n1254) );
INV_X1 U950 ( .A(n1184), .ZN(n1257) );
XNOR2_X1 U951 ( .A(n1163), .B(n1258), .ZN(n1184) );
AND2_X1 U952 ( .A1(n1089), .A2(G224), .ZN(n1258) );
XNOR2_X1 U953 ( .A(n1124), .B(n1101), .ZN(n1256) );
XNOR2_X1 U954 ( .A(n1259), .B(n1260), .ZN(n1124) );
XNOR2_X1 U955 ( .A(G122), .B(n1261), .ZN(n1260) );
XNOR2_X1 U956 ( .A(KEYINPUT34), .B(KEYINPUT31), .ZN(n1261) );
XOR2_X1 U957 ( .A(n1262), .B(n1263), .Z(n1259) );
XOR2_X1 U958 ( .A(n1264), .B(n1265), .Z(n1262) );
NOR2_X1 U959 ( .A1(G104), .A2(KEYINPUT42), .ZN(n1265) );
NAND2_X1 U960 ( .A1(G214), .A2(n1253), .ZN(n1058) );
NAND2_X1 U961 ( .A1(n1266), .A2(n1255), .ZN(n1253) );
NAND2_X1 U962 ( .A1(n1032), .A2(n1267), .ZN(n1251) );
NAND3_X1 U963 ( .A1(n1126), .A2(n1240), .A3(G902), .ZN(n1267) );
NOR2_X1 U964 ( .A1(n1241), .A2(G898), .ZN(n1126) );
XOR2_X1 U965 ( .A(G953), .B(KEYINPUT18), .Z(n1241) );
NAND3_X1 U966 ( .A1(n1240), .A2(n1089), .A3(G952), .ZN(n1032) );
NAND2_X1 U967 ( .A1(G237), .A2(G234), .ZN(n1240) );
NOR2_X1 U968 ( .A1(n1210), .A2(n1209), .ZN(n1056) );
XNOR2_X1 U969 ( .A(n1268), .B(n1269), .ZN(n1209) );
INV_X1 U970 ( .A(n1083), .ZN(n1269) );
NOR2_X1 U971 ( .A1(n1146), .A2(G902), .ZN(n1083) );
INV_X1 U972 ( .A(n1144), .ZN(n1146) );
XNOR2_X1 U973 ( .A(n1270), .B(n1271), .ZN(n1144) );
XOR2_X1 U974 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U975 ( .A(G113), .B(G104), .Z(n1273) );
XNOR2_X1 U976 ( .A(G131), .B(n1274), .ZN(n1272) );
XOR2_X1 U977 ( .A(n1275), .B(n1276), .Z(n1270) );
XOR2_X1 U978 ( .A(n1277), .B(n1278), .Z(n1275) );
AND3_X1 U979 ( .A1(G214), .A2(n1089), .A3(n1266), .ZN(n1278) );
NAND2_X1 U980 ( .A1(KEYINPUT4), .A2(n1279), .ZN(n1277) );
NAND2_X1 U981 ( .A1(KEYINPUT55), .A2(n1085), .ZN(n1268) );
INV_X1 U982 ( .A(G475), .ZN(n1085) );
XOR2_X1 U983 ( .A(n1280), .B(n1140), .Z(n1210) );
INV_X1 U984 ( .A(G478), .ZN(n1140) );
NAND2_X1 U985 ( .A1(n1281), .A2(n1255), .ZN(n1280) );
XNOR2_X1 U986 ( .A(n1139), .B(KEYINPUT54), .ZN(n1281) );
XNOR2_X1 U987 ( .A(n1282), .B(KEYINPUT8), .ZN(n1139) );
XOR2_X1 U988 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U989 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U990 ( .A(n1287), .B(G116), .ZN(n1286) );
XOR2_X1 U991 ( .A(KEYINPUT29), .B(G143), .Z(n1285) );
XOR2_X1 U992 ( .A(n1288), .B(n1289), .Z(n1283) );
XNOR2_X1 U993 ( .A(n1290), .B(n1291), .ZN(n1289) );
NOR2_X1 U994 ( .A1(G128), .A2(KEYINPUT23), .ZN(n1291) );
NAND2_X1 U995 ( .A1(KEYINPUT3), .A2(n1274), .ZN(n1290) );
INV_X1 U996 ( .A(G122), .ZN(n1274) );
XOR2_X1 U997 ( .A(n1292), .B(G107), .Z(n1288) );
NAND2_X1 U998 ( .A1(G217), .A2(n1293), .ZN(n1292) );
NOR2_X1 U999 ( .A1(n1247), .A2(n1246), .ZN(n1201) );
XOR2_X1 U1000 ( .A(n1294), .B(n1075), .Z(n1246) );
NOR2_X1 U1001 ( .A1(n1134), .A2(G902), .ZN(n1075) );
XNOR2_X1 U1002 ( .A(n1295), .B(n1296), .ZN(n1134) );
XOR2_X1 U1003 ( .A(n1297), .B(n1298), .Z(n1296) );
XNOR2_X1 U1004 ( .A(n1299), .B(G119), .ZN(n1298) );
XOR2_X1 U1005 ( .A(KEYINPUT56), .B(G146), .Z(n1297) );
XOR2_X1 U1006 ( .A(n1300), .B(n1301), .Z(n1295) );
XNOR2_X1 U1007 ( .A(G110), .B(n1302), .ZN(n1301) );
NAND3_X1 U1008 ( .A1(n1293), .A2(G221), .A3(KEYINPUT24), .ZN(n1302) );
AND2_X1 U1009 ( .A1(G234), .A2(n1089), .ZN(n1293) );
XNOR2_X1 U1010 ( .A(n1279), .B(n1303), .ZN(n1300) );
XNOR2_X1 U1011 ( .A(G140), .B(n1304), .ZN(n1279) );
INV_X1 U1012 ( .A(n1101), .ZN(n1304) );
XOR2_X1 U1013 ( .A(G125), .B(KEYINPUT5), .Z(n1101) );
NAND2_X1 U1014 ( .A1(KEYINPUT26), .A2(n1077), .ZN(n1294) );
INV_X1 U1015 ( .A(n1082), .ZN(n1077) );
NAND2_X1 U1016 ( .A1(G217), .A2(n1305), .ZN(n1082) );
XOR2_X1 U1017 ( .A(n1069), .B(n1306), .Z(n1247) );
NOR2_X1 U1018 ( .A1(KEYINPUT47), .A2(n1165), .ZN(n1306) );
INV_X1 U1019 ( .A(G472), .ZN(n1165) );
AND2_X1 U1020 ( .A1(n1307), .A2(n1255), .ZN(n1069) );
XNOR2_X1 U1021 ( .A(n1151), .B(n1308), .ZN(n1307) );
XNOR2_X1 U1022 ( .A(n1157), .B(n1309), .ZN(n1308) );
NOR2_X1 U1023 ( .A1(KEYINPUT58), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1024 ( .A(n1311), .B(n1163), .Z(n1310) );
XNOR2_X1 U1025 ( .A(G128), .B(n1276), .ZN(n1163) );
XOR2_X1 U1026 ( .A(G143), .B(G146), .Z(n1276) );
NAND2_X1 U1027 ( .A1(KEYINPUT25), .A2(n1162), .ZN(n1311) );
XNOR2_X1 U1028 ( .A(n1264), .B(KEYINPUT14), .ZN(n1157) );
XNOR2_X1 U1029 ( .A(G113), .B(n1312), .ZN(n1264) );
XOR2_X1 U1030 ( .A(G119), .B(G116), .Z(n1312) );
AND2_X1 U1031 ( .A1(n1313), .A2(n1314), .ZN(n1151) );
NAND2_X1 U1032 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND3_X1 U1033 ( .A1(n1266), .A2(n1089), .A3(G210), .ZN(n1315) );
NAND4_X1 U1034 ( .A1(n1266), .A2(n1089), .A3(G210), .A4(G101), .ZN(n1313) );
INV_X1 U1035 ( .A(G237), .ZN(n1266) );
XNOR2_X1 U1036 ( .A(n1192), .B(KEYINPUT11), .ZN(n1250) );
NOR2_X1 U1037 ( .A1(n1317), .A2(n1248), .ZN(n1192) );
XOR2_X1 U1038 ( .A(n1055), .B(KEYINPUT48), .Z(n1248) );
NAND2_X1 U1039 ( .A1(G221), .A2(n1305), .ZN(n1055) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1255), .ZN(n1305) );
INV_X1 U1041 ( .A(n1054), .ZN(n1317) );
XNOR2_X1 U1042 ( .A(n1318), .B(n1072), .ZN(n1054) );
INV_X1 U1043 ( .A(G469), .ZN(n1072) );
NAND2_X1 U1044 ( .A1(KEYINPUT41), .A2(n1073), .ZN(n1318) );
NAND2_X1 U1045 ( .A1(n1319), .A2(n1255), .ZN(n1073) );
INV_X1 U1046 ( .A(G902), .ZN(n1255) );
XOR2_X1 U1047 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1048 ( .A(G140), .B(n1179), .ZN(n1321) );
NAND2_X1 U1049 ( .A1(G227), .A2(n1322), .ZN(n1179) );
XNOR2_X1 U1050 ( .A(KEYINPUT43), .B(n1089), .ZN(n1322) );
INV_X1 U1051 ( .A(G953), .ZN(n1089) );
XOR2_X1 U1052 ( .A(n1172), .B(n1263), .Z(n1320) );
XNOR2_X1 U1053 ( .A(n1176), .B(n1173), .ZN(n1263) );
XNOR2_X1 U1054 ( .A(G107), .B(n1316), .ZN(n1173) );
INV_X1 U1055 ( .A(G101), .ZN(n1316) );
INV_X1 U1056 ( .A(G110), .ZN(n1176) );
XNOR2_X1 U1057 ( .A(n1323), .B(n1324), .ZN(n1172) );
INV_X1 U1058 ( .A(n1108), .ZN(n1324) );
XNOR2_X1 U1059 ( .A(n1325), .B(n1326), .ZN(n1108) );
NOR2_X1 U1060 ( .A1(G146), .A2(KEYINPUT19), .ZN(n1326) );
XOR2_X1 U1061 ( .A(n1327), .B(G143), .Z(n1325) );
NAND2_X1 U1062 ( .A1(KEYINPUT12), .A2(n1299), .ZN(n1327) );
INV_X1 U1063 ( .A(G128), .ZN(n1299) );
XOR2_X1 U1064 ( .A(n1162), .B(G104), .Z(n1323) );
XOR2_X1 U1065 ( .A(n1328), .B(n1109), .Z(n1162) );
XOR2_X1 U1066 ( .A(G131), .B(n1303), .Z(n1109) );
XOR2_X1 U1067 ( .A(G137), .B(KEYINPUT62), .Z(n1303) );
NAND2_X1 U1068 ( .A1(KEYINPUT52), .A2(n1287), .ZN(n1328) );
INV_X1 U1069 ( .A(G134), .ZN(n1287) );
endmodule


