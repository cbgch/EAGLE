//Key = 0010100101101101000011100100010100000010101110101001001000011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378;

XOR2_X1 U764 ( .A(G107), .B(n1051), .Z(G9) );
NOR2_X1 U765 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U766 ( .A1(n1054), .A2(n1055), .ZN(G75) );
NOR4_X1 U767 ( .A1(n1056), .A2(n1057), .A3(G953), .A4(n1058), .ZN(n1055) );
NOR3_X1 U768 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1057) );
NOR2_X1 U769 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U770 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U771 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
AND2_X1 U772 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR3_X1 U773 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1066) );
NOR2_X1 U774 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U775 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1071) );
NOR3_X1 U777 ( .A1(n1079), .A2(n1080), .A3(n1070), .ZN(n1062) );
NAND2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1056) );
XOR2_X1 U779 ( .A(KEYINPUT24), .B(n1083), .Z(n1082) );
NOR2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR4_X1 U781 ( .A1(n1086), .A2(n1087), .A3(n1061), .A4(n1070), .ZN(n1085) );
OR2_X1 U782 ( .A1(n1059), .A2(n1079), .ZN(n1086) );
NOR4_X1 U783 ( .A1(n1088), .A2(n1089), .A3(n1065), .A4(n1059), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1091), .ZN(n1088) );
NAND2_X1 U786 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND3_X1 U787 ( .A1(n1095), .A2(n1096), .A3(n1069), .ZN(n1094) );
INV_X1 U788 ( .A(n1079), .ZN(n1069) );
NAND2_X1 U789 ( .A1(n1077), .A2(n1078), .ZN(n1079) );
NAND3_X1 U790 ( .A1(n1097), .A2(n1092), .A3(n1077), .ZN(n1093) );
NOR3_X1 U791 ( .A1(n1058), .A2(G953), .A3(G952), .ZN(n1054) );
AND4_X1 U792 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1058) );
NOR4_X1 U793 ( .A1(n1102), .A2(n1073), .A3(n1103), .A4(n1104), .ZN(n1101) );
XOR2_X1 U794 ( .A(n1105), .B(n1106), .Z(n1103) );
NOR2_X1 U795 ( .A1(n1107), .A2(KEYINPUT39), .ZN(n1106) );
XOR2_X1 U796 ( .A(n1108), .B(KEYINPUT47), .Z(n1105) );
NOR3_X1 U797 ( .A1(n1065), .A2(n1109), .A3(n1110), .ZN(n1100) );
AND2_X1 U798 ( .A1(n1111), .A2(KEYINPUT15), .ZN(n1110) );
NOR2_X1 U799 ( .A1(KEYINPUT15), .A2(n1112), .ZN(n1109) );
NOR2_X1 U800 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
INV_X1 U801 ( .A(G472), .ZN(n1114) );
OR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(n1099) );
NAND2_X1 U803 ( .A1(n1117), .A2(n1115), .ZN(n1098) );
XOR2_X1 U804 ( .A(KEYINPUT18), .B(n1116), .Z(n1117) );
INV_X1 U805 ( .A(n1118), .ZN(n1116) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(G72) );
XOR2_X1 U807 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U809 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
XOR2_X1 U810 ( .A(KEYINPUT2), .B(G227), .Z(n1126) );
NAND2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(n1121) );
XOR2_X1 U812 ( .A(KEYINPUT25), .B(G953), .Z(n1127) );
NAND2_X1 U813 ( .A1(n1129), .A2(n1130), .ZN(n1119) );
XOR2_X1 U814 ( .A(n1131), .B(n1132), .Z(n1129) );
XOR2_X1 U815 ( .A(KEYINPUT51), .B(n1133), .Z(n1132) );
XOR2_X1 U816 ( .A(n1134), .B(n1135), .Z(n1131) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(G69) );
NAND2_X1 U818 ( .A1(G953), .A2(n1138), .ZN(n1137) );
NAND2_X1 U819 ( .A1(G898), .A2(G224), .ZN(n1138) );
NAND2_X1 U820 ( .A1(n1139), .A2(KEYINPUT7), .ZN(n1136) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U822 ( .A1(KEYINPUT63), .A2(n1142), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1143), .A2(G953), .ZN(n1142) );
NOR2_X1 U824 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND3_X1 U825 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1140) );
XOR2_X1 U826 ( .A(KEYINPUT21), .B(n1149), .Z(n1148) );
NOR2_X1 U827 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U828 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
XNOR2_X1 U829 ( .A(n1152), .B(KEYINPUT29), .ZN(n1150) );
NAND2_X1 U830 ( .A1(G953), .A2(n1153), .ZN(n1146) );
NOR2_X1 U831 ( .A1(n1154), .A2(n1155), .ZN(G66) );
NOR3_X1 U832 ( .A1(n1107), .A2(n1156), .A3(n1157), .ZN(n1155) );
NOR3_X1 U833 ( .A1(n1158), .A2(n1108), .A3(n1159), .ZN(n1157) );
NOR2_X1 U834 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
NOR2_X1 U835 ( .A1(n1081), .A2(n1108), .ZN(n1160) );
NOR2_X1 U836 ( .A1(n1154), .A2(n1162), .ZN(G63) );
XOR2_X1 U837 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U838 ( .A1(KEYINPUT27), .A2(n1165), .ZN(n1164) );
AND2_X1 U839 ( .A1(G478), .A2(n1166), .ZN(n1163) );
NOR2_X1 U840 ( .A1(n1167), .A2(n1168), .ZN(G60) );
XOR2_X1 U841 ( .A(n1169), .B(n1170), .Z(n1168) );
NAND2_X1 U842 ( .A1(n1166), .A2(G475), .ZN(n1169) );
NOR2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1167) );
XOR2_X1 U844 ( .A(KEYINPUT59), .B(G953), .Z(n1172) );
XOR2_X1 U845 ( .A(KEYINPUT16), .B(G952), .Z(n1171) );
XNOR2_X1 U846 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U847 ( .A1(n1154), .A2(n1174), .ZN(G57) );
XOR2_X1 U848 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U849 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U850 ( .A1(n1166), .A2(G472), .ZN(n1178) );
NAND2_X1 U851 ( .A1(n1179), .A2(KEYINPUT4), .ZN(n1177) );
XOR2_X1 U852 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U853 ( .A(n1182), .B(n1183), .Z(n1175) );
XOR2_X1 U854 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U855 ( .A1(n1154), .A2(n1186), .ZN(G54) );
XOR2_X1 U856 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U857 ( .A(n1180), .B(n1189), .Z(n1188) );
XOR2_X1 U858 ( .A(n1190), .B(n1191), .Z(n1187) );
XOR2_X1 U859 ( .A(n1192), .B(KEYINPUT35), .Z(n1191) );
NAND2_X1 U860 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U861 ( .A(n1195), .ZN(n1193) );
NAND2_X1 U862 ( .A1(n1166), .A2(G469), .ZN(n1190) );
NOR2_X1 U863 ( .A1(n1196), .A2(n1197), .ZN(G51) );
XOR2_X1 U864 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U865 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR3_X1 U866 ( .A1(n1159), .A2(KEYINPUT52), .A3(n1202), .ZN(n1200) );
INV_X1 U867 ( .A(n1166), .ZN(n1159) );
NOR2_X1 U868 ( .A1(n1203), .A2(n1081), .ZN(n1166) );
NOR3_X1 U869 ( .A1(n1128), .A2(n1204), .A3(n1145), .ZN(n1081) );
NAND4_X1 U870 ( .A1(n1205), .A2(n1173), .A3(n1206), .A4(n1207), .ZN(n1145) );
NAND3_X1 U871 ( .A1(n1208), .A2(n1092), .A3(n1209), .ZN(n1173) );
NAND2_X1 U872 ( .A1(n1210), .A2(n1211), .ZN(n1205) );
XNOR2_X1 U873 ( .A(KEYINPUT32), .B(n1052), .ZN(n1211) );
NAND4_X1 U874 ( .A1(n1097), .A2(n1092), .A3(n1212), .A4(n1213), .ZN(n1052) );
XOR2_X1 U875 ( .A(KEYINPUT17), .B(n1144), .Z(n1204) );
NAND4_X1 U876 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1144) );
NAND3_X1 U877 ( .A1(n1090), .A2(n1218), .A3(n1219), .ZN(n1214) );
XNOR2_X1 U878 ( .A(KEYINPUT38), .B(n1213), .ZN(n1218) );
NAND3_X1 U879 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1128) );
AND3_X1 U880 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1222) );
NAND4_X1 U881 ( .A1(n1226), .A2(n1227), .A3(n1210), .A4(n1228), .ZN(n1221) );
NAND2_X1 U882 ( .A1(n1087), .A2(n1080), .ZN(n1228) );
NAND2_X1 U883 ( .A1(n1077), .A2(n1229), .ZN(n1220) );
NAND3_X1 U884 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1229) );
XNOR2_X1 U885 ( .A(n1233), .B(KEYINPUT34), .ZN(n1232) );
XOR2_X1 U886 ( .A(n1234), .B(KEYINPUT37), .Z(n1230) );
XOR2_X1 U887 ( .A(n1235), .B(n1236), .Z(n1198) );
NOR2_X1 U888 ( .A1(KEYINPUT57), .A2(n1237), .ZN(n1236) );
XNOR2_X1 U889 ( .A(n1154), .B(KEYINPUT60), .ZN(n1196) );
AND2_X1 U890 ( .A1(n1238), .A2(G953), .ZN(n1154) );
XNOR2_X1 U891 ( .A(KEYINPUT16), .B(G952), .ZN(n1238) );
NAND2_X1 U892 ( .A1(n1239), .A2(n1240), .ZN(G48) );
NAND2_X1 U893 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U894 ( .A(KEYINPUT20), .B(n1243), .Z(n1239) );
NOR2_X1 U895 ( .A1(n1241), .A2(n1242), .ZN(n1243) );
INV_X1 U896 ( .A(G146), .ZN(n1242) );
AND4_X1 U897 ( .A1(n1226), .A2(n1227), .A3(n1210), .A4(n1244), .ZN(n1241) );
XOR2_X1 U898 ( .A(KEYINPUT3), .B(n1209), .Z(n1244) );
XNOR2_X1 U899 ( .A(n1223), .B(n1245), .ZN(G45) );
NOR2_X1 U900 ( .A1(KEYINPUT6), .A2(n1246), .ZN(n1245) );
NAND3_X1 U901 ( .A1(n1227), .A2(n1210), .A3(n1247), .ZN(n1223) );
NOR3_X1 U902 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
XNOR2_X1 U903 ( .A(G140), .B(n1251), .ZN(G42) );
NAND2_X1 U904 ( .A1(n1233), .A2(n1077), .ZN(n1251) );
AND3_X1 U905 ( .A1(n1209), .A2(n1068), .A3(n1227), .ZN(n1233) );
NAND2_X1 U906 ( .A1(n1252), .A2(n1253), .ZN(G39) );
OR2_X1 U907 ( .A1(G137), .A2(KEYINPUT43), .ZN(n1253) );
XOR2_X1 U908 ( .A(n1254), .B(n1255), .Z(n1252) );
NOR2_X1 U909 ( .A1(n1256), .A2(n1234), .ZN(n1255) );
NAND3_X1 U910 ( .A1(n1227), .A2(n1257), .A3(n1226), .ZN(n1234) );
INV_X1 U911 ( .A(n1077), .ZN(n1256) );
NAND2_X1 U912 ( .A1(KEYINPUT43), .A2(G137), .ZN(n1254) );
XNOR2_X1 U913 ( .A(G134), .B(n1258), .ZN(G36) );
NAND2_X1 U914 ( .A1(n1077), .A2(n1259), .ZN(n1258) );
XNOR2_X1 U915 ( .A(KEYINPUT55), .B(n1231), .ZN(n1259) );
NAND2_X1 U916 ( .A1(n1219), .A2(n1227), .ZN(n1231) );
NAND2_X1 U917 ( .A1(n1260), .A2(n1261), .ZN(G33) );
NAND2_X1 U918 ( .A1(n1262), .A2(G131), .ZN(n1261) );
XOR2_X1 U919 ( .A(n1225), .B(KEYINPUT50), .Z(n1262) );
XOR2_X1 U920 ( .A(KEYINPUT12), .B(n1263), .Z(n1260) );
NOR2_X1 U921 ( .A1(G131), .A2(n1264), .ZN(n1263) );
XOR2_X1 U922 ( .A(n1225), .B(KEYINPUT28), .Z(n1264) );
NAND4_X1 U923 ( .A1(n1227), .A2(n1077), .A3(n1209), .A4(n1095), .ZN(n1225) );
NOR2_X1 U924 ( .A1(n1075), .A2(n1102), .ZN(n1077) );
INV_X1 U925 ( .A(n1076), .ZN(n1102) );
AND2_X1 U926 ( .A1(n1097), .A2(n1265), .ZN(n1227) );
XOR2_X1 U927 ( .A(n1266), .B(n1267), .Z(G30) );
NAND4_X1 U928 ( .A1(n1268), .A2(n1265), .A3(n1212), .A4(n1269), .ZN(n1267) );
AND2_X1 U929 ( .A1(n1210), .A2(n1226), .ZN(n1269) );
INV_X1 U930 ( .A(n1080), .ZN(n1212) );
XOR2_X1 U931 ( .A(KEYINPUT58), .B(n1097), .Z(n1268) );
XOR2_X1 U932 ( .A(n1185), .B(n1206), .Z(G3) );
NAND3_X1 U933 ( .A1(n1257), .A2(n1095), .A3(n1208), .ZN(n1206) );
XNOR2_X1 U934 ( .A(G125), .B(n1224), .ZN(G27) );
NAND4_X1 U935 ( .A1(n1090), .A2(n1209), .A3(n1068), .A4(n1265), .ZN(n1224) );
NAND2_X1 U936 ( .A1(n1059), .A2(n1270), .ZN(n1265) );
NAND3_X1 U937 ( .A1(G902), .A2(n1271), .A3(n1272), .ZN(n1270) );
INV_X1 U938 ( .A(n1130), .ZN(n1272) );
NAND2_X1 U939 ( .A1(G953), .A2(n1125), .ZN(n1130) );
INV_X1 U940 ( .A(G900), .ZN(n1125) );
NAND2_X1 U941 ( .A1(n1273), .A2(n1274), .ZN(G24) );
OR2_X1 U942 ( .A1(n1215), .A2(G122), .ZN(n1274) );
XOR2_X1 U943 ( .A(n1275), .B(KEYINPUT23), .Z(n1273) );
NAND2_X1 U944 ( .A1(G122), .A2(n1215), .ZN(n1275) );
NAND4_X1 U945 ( .A1(n1276), .A2(n1092), .A3(n1277), .A4(n1278), .ZN(n1215) );
XNOR2_X1 U946 ( .A(G119), .B(n1216), .ZN(G21) );
NAND3_X1 U947 ( .A1(n1226), .A2(n1257), .A3(n1276), .ZN(n1216) );
NOR2_X1 U948 ( .A1(n1279), .A2(n1280), .ZN(n1226) );
XOR2_X1 U949 ( .A(n1281), .B(n1282), .Z(G18) );
NAND2_X1 U950 ( .A1(n1276), .A2(n1219), .ZN(n1282) );
NOR2_X1 U951 ( .A1(n1080), .A2(n1248), .ZN(n1219) );
INV_X1 U952 ( .A(n1095), .ZN(n1248) );
NAND2_X1 U953 ( .A1(n1249), .A2(n1277), .ZN(n1080) );
INV_X1 U954 ( .A(n1250), .ZN(n1277) );
XOR2_X1 U955 ( .A(n1283), .B(n1217), .Z(G15) );
NAND3_X1 U956 ( .A1(n1209), .A2(n1095), .A3(n1276), .ZN(n1217) );
AND2_X1 U957 ( .A1(n1090), .A2(n1213), .ZN(n1276) );
NOR3_X1 U958 ( .A1(n1061), .A2(n1073), .A3(n1053), .ZN(n1090) );
NAND2_X1 U959 ( .A1(n1284), .A2(n1285), .ZN(n1095) );
OR3_X1 U960 ( .A1(n1280), .A2(n1286), .A3(KEYINPUT8), .ZN(n1285) );
NAND2_X1 U961 ( .A1(KEYINPUT8), .A2(n1092), .ZN(n1284) );
INV_X1 U962 ( .A(n1070), .ZN(n1092) );
NAND2_X1 U963 ( .A1(n1280), .A2(n1279), .ZN(n1070) );
INV_X1 U964 ( .A(n1111), .ZN(n1280) );
INV_X1 U965 ( .A(n1087), .ZN(n1209) );
NAND2_X1 U966 ( .A1(n1250), .A2(n1278), .ZN(n1087) );
INV_X1 U967 ( .A(n1249), .ZN(n1278) );
XNOR2_X1 U968 ( .A(G110), .B(n1207), .ZN(G12) );
NAND3_X1 U969 ( .A1(n1068), .A2(n1257), .A3(n1208), .ZN(n1207) );
AND3_X1 U970 ( .A1(n1097), .A2(n1213), .A3(n1210), .ZN(n1208) );
INV_X1 U971 ( .A(n1053), .ZN(n1210) );
NAND2_X1 U972 ( .A1(n1075), .A2(n1076), .ZN(n1053) );
NAND2_X1 U973 ( .A1(G214), .A2(n1287), .ZN(n1076) );
XOR2_X1 U974 ( .A(n1118), .B(n1115), .Z(n1075) );
NAND2_X1 U975 ( .A1(G210), .A2(n1287), .ZN(n1115) );
NAND2_X1 U976 ( .A1(n1288), .A2(n1203), .ZN(n1287) );
NAND2_X1 U977 ( .A1(n1289), .A2(n1203), .ZN(n1118) );
XOR2_X1 U978 ( .A(n1201), .B(n1290), .Z(n1289) );
XOR2_X1 U979 ( .A(n1235), .B(n1237), .Z(n1290) );
XNOR2_X1 U980 ( .A(n1181), .B(G125), .ZN(n1237) );
NAND2_X1 U981 ( .A1(G224), .A2(n1124), .ZN(n1235) );
XNOR2_X1 U982 ( .A(n1291), .B(n1152), .ZN(n1201) );
XNOR2_X1 U983 ( .A(n1292), .B(n1293), .ZN(n1152) );
XNOR2_X1 U984 ( .A(n1294), .B(n1295), .ZN(n1293) );
XOR2_X1 U985 ( .A(n1296), .B(n1297), .Z(n1292) );
XNOR2_X1 U986 ( .A(KEYINPUT40), .B(KEYINPUT36), .ZN(n1296) );
NAND2_X1 U987 ( .A1(KEYINPUT54), .A2(n1298), .ZN(n1291) );
INV_X1 U988 ( .A(n1151), .ZN(n1298) );
XOR2_X1 U989 ( .A(G110), .B(G122), .Z(n1151) );
NAND2_X1 U990 ( .A1(n1059), .A2(n1299), .ZN(n1213) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1271), .A4(n1153), .ZN(n1299) );
INV_X1 U992 ( .A(G898), .ZN(n1153) );
NAND3_X1 U993 ( .A1(n1271), .A2(n1124), .A3(G952), .ZN(n1059) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1271) );
NOR2_X1 U995 ( .A1(n1096), .A2(n1073), .ZN(n1097) );
INV_X1 U996 ( .A(n1078), .ZN(n1073) );
NAND2_X1 U997 ( .A1(G221), .A2(n1300), .ZN(n1078) );
INV_X1 U998 ( .A(n1061), .ZN(n1096) );
XNOR2_X1 U999 ( .A(n1104), .B(KEYINPUT9), .ZN(n1061) );
XNOR2_X1 U1000 ( .A(n1301), .B(G469), .ZN(n1104) );
NAND2_X1 U1001 ( .A1(n1302), .A2(n1203), .ZN(n1301) );
XOR2_X1 U1002 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1003 ( .A(n1305), .B(n1189), .Z(n1304) );
XOR2_X1 U1004 ( .A(n1306), .B(n1307), .Z(n1189) );
XOR2_X1 U1005 ( .A(KEYINPUT0), .B(n1308), .Z(n1307) );
NOR2_X1 U1006 ( .A1(G104), .A2(KEYINPUT11), .ZN(n1308) );
XOR2_X1 U1007 ( .A(n1134), .B(n1295), .Z(n1306) );
XOR2_X1 U1008 ( .A(G107), .B(G101), .Z(n1295) );
XOR2_X1 U1009 ( .A(n1309), .B(n1310), .Z(n1134) );
NAND2_X1 U1010 ( .A1(KEYINPUT44), .A2(G146), .ZN(n1309) );
NAND2_X1 U1011 ( .A1(KEYINPUT62), .A2(n1311), .ZN(n1305) );
INV_X1 U1012 ( .A(n1180), .ZN(n1311) );
XOR2_X1 U1013 ( .A(KEYINPUT48), .B(n1312), .Z(n1303) );
NOR2_X1 U1014 ( .A1(n1195), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1015 ( .A(n1194), .B(KEYINPUT10), .Z(n1313) );
NAND2_X1 U1016 ( .A1(n1314), .A2(n1315), .ZN(n1194) );
NAND2_X1 U1017 ( .A1(G227), .A2(n1124), .ZN(n1315) );
NOR3_X1 U1018 ( .A1(n1314), .A2(G953), .A3(n1316), .ZN(n1195) );
INV_X1 U1019 ( .A(G227), .ZN(n1316) );
XOR2_X1 U1020 ( .A(G140), .B(G110), .Z(n1314) );
INV_X1 U1021 ( .A(n1065), .ZN(n1257) );
NAND2_X1 U1022 ( .A1(n1250), .A2(n1249), .ZN(n1065) );
XOR2_X1 U1023 ( .A(n1317), .B(G475), .Z(n1249) );
NAND2_X1 U1024 ( .A1(n1170), .A2(n1203), .ZN(n1317) );
XNOR2_X1 U1025 ( .A(n1318), .B(n1319), .ZN(n1170) );
XNOR2_X1 U1026 ( .A(n1320), .B(n1297), .ZN(n1319) );
XOR2_X1 U1027 ( .A(G104), .B(G113), .Z(n1297) );
NAND2_X1 U1028 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U1029 ( .A(n1323), .B(KEYINPUT53), .Z(n1321) );
XNOR2_X1 U1030 ( .A(G122), .B(n1324), .ZN(n1318) );
NOR2_X1 U1031 ( .A1(KEYINPUT1), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1032 ( .A(G131), .B(n1326), .ZN(n1325) );
NOR3_X1 U1033 ( .A1(KEYINPUT49), .A2(n1327), .A3(n1328), .ZN(n1326) );
NOR3_X1 U1034 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1328) );
NOR2_X1 U1035 ( .A1(n1332), .A2(n1333), .ZN(n1327) );
NOR2_X1 U1036 ( .A1(n1330), .A2(n1331), .ZN(n1332) );
INV_X1 U1037 ( .A(G214), .ZN(n1330) );
XOR2_X1 U1038 ( .A(n1334), .B(G478), .Z(n1250) );
NAND2_X1 U1039 ( .A1(n1165), .A2(n1203), .ZN(n1334) );
XNOR2_X1 U1040 ( .A(n1335), .B(n1336), .ZN(n1165) );
XOR2_X1 U1041 ( .A(G116), .B(n1337), .Z(n1336) );
XOR2_X1 U1042 ( .A(G134), .B(G122), .Z(n1337) );
XNOR2_X1 U1043 ( .A(n1310), .B(n1338), .ZN(n1335) );
XOR2_X1 U1044 ( .A(n1339), .B(n1340), .Z(n1338) );
NAND2_X1 U1045 ( .A1(KEYINPUT31), .A2(n1341), .ZN(n1340) );
INV_X1 U1046 ( .A(G107), .ZN(n1341) );
NAND2_X1 U1047 ( .A1(G217), .A2(n1342), .ZN(n1339) );
XNOR2_X1 U1048 ( .A(n1266), .B(n1329), .ZN(n1310) );
INV_X1 U1049 ( .A(n1333), .ZN(n1329) );
NOR2_X1 U1050 ( .A1(n1111), .A2(n1279), .ZN(n1068) );
INV_X1 U1051 ( .A(n1286), .ZN(n1279) );
NAND2_X1 U1052 ( .A1(n1343), .A2(n1344), .ZN(n1286) );
NAND2_X1 U1053 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1054 ( .A(n1108), .B(KEYINPUT46), .Z(n1345) );
NAND2_X1 U1055 ( .A1(n1347), .A2(n1107), .ZN(n1343) );
INV_X1 U1056 ( .A(n1346), .ZN(n1107) );
NAND2_X1 U1057 ( .A1(n1158), .A2(n1203), .ZN(n1346) );
INV_X1 U1058 ( .A(n1161), .ZN(n1158) );
XOR2_X1 U1059 ( .A(n1348), .B(n1349), .Z(n1161) );
XNOR2_X1 U1060 ( .A(n1350), .B(n1351), .ZN(n1349) );
NOR2_X1 U1061 ( .A1(KEYINPUT45), .A2(n1352), .ZN(n1351) );
INV_X1 U1062 ( .A(G137), .ZN(n1352) );
NAND2_X1 U1063 ( .A1(KEYINPUT13), .A2(n1353), .ZN(n1350) );
XOR2_X1 U1064 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1065 ( .A(G110), .B(n1356), .ZN(n1355) );
NAND2_X1 U1066 ( .A1(n1357), .A2(n1322), .ZN(n1356) );
NAND2_X1 U1067 ( .A1(G146), .A2(n1133), .ZN(n1322) );
XOR2_X1 U1068 ( .A(n1323), .B(KEYINPUT41), .Z(n1357) );
OR2_X1 U1069 ( .A1(n1133), .A2(G146), .ZN(n1323) );
XOR2_X1 U1070 ( .A(G125), .B(G140), .Z(n1133) );
XOR2_X1 U1071 ( .A(G128), .B(G119), .Z(n1354) );
NAND2_X1 U1072 ( .A1(n1342), .A2(G221), .ZN(n1348) );
AND2_X1 U1073 ( .A1(G234), .A2(n1124), .ZN(n1342) );
XNOR2_X1 U1074 ( .A(KEYINPUT42), .B(n1108), .ZN(n1347) );
NAND2_X1 U1075 ( .A1(G217), .A2(n1300), .ZN(n1108) );
NAND2_X1 U1076 ( .A1(G234), .A2(n1203), .ZN(n1300) );
XOR2_X1 U1077 ( .A(n1113), .B(G472), .Z(n1111) );
AND2_X1 U1078 ( .A1(n1358), .A2(n1203), .ZN(n1113) );
INV_X1 U1079 ( .A(G902), .ZN(n1203) );
XOR2_X1 U1080 ( .A(n1359), .B(n1360), .Z(n1358) );
XOR2_X1 U1081 ( .A(n1361), .B(n1181), .Z(n1360) );
XOR2_X1 U1082 ( .A(n1362), .B(n1333), .Z(n1181) );
XOR2_X1 U1083 ( .A(n1246), .B(KEYINPUT22), .Z(n1333) );
INV_X1 U1084 ( .A(G143), .ZN(n1246) );
XNOR2_X1 U1085 ( .A(n1363), .B(n1364), .ZN(n1362) );
NOR2_X1 U1086 ( .A1(KEYINPUT19), .A2(n1266), .ZN(n1364) );
INV_X1 U1087 ( .A(G128), .ZN(n1266) );
NOR2_X1 U1088 ( .A1(G146), .A2(KEYINPUT14), .ZN(n1363) );
NOR2_X1 U1089 ( .A1(KEYINPUT56), .A2(n1180), .ZN(n1361) );
XNOR2_X1 U1090 ( .A(n1135), .B(KEYINPUT26), .ZN(n1180) );
XOR2_X1 U1091 ( .A(G131), .B(n1365), .Z(n1135) );
XOR2_X1 U1092 ( .A(G137), .B(G134), .Z(n1365) );
XOR2_X1 U1093 ( .A(n1366), .B(n1182), .Z(n1359) );
NAND2_X1 U1094 ( .A1(n1367), .A2(n1368), .ZN(n1182) );
NAND2_X1 U1095 ( .A1(n1369), .A2(n1283), .ZN(n1368) );
XOR2_X1 U1096 ( .A(n1370), .B(KEYINPUT30), .Z(n1367) );
OR2_X1 U1097 ( .A1(n1369), .A2(n1283), .ZN(n1370) );
INV_X1 U1098 ( .A(G113), .ZN(n1283) );
NAND2_X1 U1099 ( .A1(n1371), .A2(n1372), .ZN(n1369) );
NAND2_X1 U1100 ( .A1(KEYINPUT61), .A2(n1294), .ZN(n1372) );
XNOR2_X1 U1101 ( .A(G116), .B(G119), .ZN(n1294) );
OR3_X1 U1102 ( .A1(n1281), .A2(G119), .A3(KEYINPUT61), .ZN(n1371) );
INV_X1 U1103 ( .A(G116), .ZN(n1281) );
NAND3_X1 U1104 ( .A1(n1373), .A2(n1374), .A3(n1375), .ZN(n1366) );
OR2_X1 U1105 ( .A1(n1376), .A2(n1184), .ZN(n1375) );
NAND3_X1 U1106 ( .A1(n1184), .A2(n1376), .A3(G101), .ZN(n1374) );
NAND2_X1 U1107 ( .A1(n1377), .A2(n1185), .ZN(n1373) );
INV_X1 U1108 ( .A(G101), .ZN(n1185) );
NAND2_X1 U1109 ( .A1(n1378), .A2(n1376), .ZN(n1377) );
INV_X1 U1110 ( .A(KEYINPUT5), .ZN(n1376) );
XOR2_X1 U1111 ( .A(KEYINPUT33), .B(n1184), .Z(n1378) );
NOR2_X1 U1112 ( .A1(n1331), .A2(n1202), .ZN(n1184) );
INV_X1 U1113 ( .A(G210), .ZN(n1202) );
NAND2_X1 U1114 ( .A1(n1288), .A2(n1124), .ZN(n1331) );
INV_X1 U1115 ( .A(G953), .ZN(n1124) );
INV_X1 U1116 ( .A(G237), .ZN(n1288) );
endmodule


