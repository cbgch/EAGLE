//Key = 1010101001101000011010000011111100010010010001001000101110110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350;

XOR2_X1 U745 ( .A(G107), .B(n1016), .Z(G9) );
NOR2_X1 U746 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR2_X1 U747 ( .A1(G952), .A2(n1019), .ZN(n1018) );
NOR4_X1 U748 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1017) );
NAND3_X1 U749 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1020) );
INV_X1 U750 ( .A(n1019), .ZN(n1026) );
NAND2_X1 U751 ( .A1(n1027), .A2(n1028), .ZN(n1019) );
NAND4_X1 U752 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
NOR3_X1 U753 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
XNOR2_X1 U754 ( .A(n1036), .B(n1037), .ZN(n1035) );
NOR2_X1 U755 ( .A1(KEYINPUT50), .A2(n1038), .ZN(n1037) );
XOR2_X1 U756 ( .A(n1039), .B(KEYINPUT54), .Z(n1038) );
XOR2_X1 U757 ( .A(n1040), .B(n1041), .Z(n1034) );
NAND2_X1 U758 ( .A1(KEYINPUT0), .A2(n1042), .ZN(n1040) );
NAND3_X1 U759 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1033) );
NOR3_X1 U760 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1031) );
NOR3_X1 U761 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
INV_X1 U762 ( .A(KEYINPUT31), .ZN(n1049) );
NOR2_X1 U763 ( .A1(KEYINPUT31), .A2(G475), .ZN(n1047) );
XNOR2_X1 U764 ( .A(G469), .B(n1052), .ZN(n1046) );
XNOR2_X1 U765 ( .A(n1053), .B(n1054), .ZN(n1029) );
XNOR2_X1 U766 ( .A(KEYINPUT7), .B(KEYINPUT32), .ZN(n1053) );
NAND3_X1 U767 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1025) );
NAND2_X1 U768 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND3_X1 U769 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NAND2_X1 U770 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND2_X1 U771 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
INV_X1 U772 ( .A(n1067), .ZN(n1063) );
NAND2_X1 U773 ( .A1(n1068), .A2(n1069), .ZN(n1058) );
NAND3_X1 U774 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U775 ( .A1(n1073), .A2(n1062), .ZN(n1072) );
NAND3_X1 U776 ( .A1(n1074), .A2(n1075), .A3(n1030), .ZN(n1071) );
XOR2_X1 U777 ( .A(KEYINPUT57), .B(n1062), .Z(n1074) );
NAND2_X1 U778 ( .A1(n1060), .A2(n1076), .ZN(n1070) );
NAND2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U780 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND4_X1 U781 ( .A1(n1060), .A2(n1081), .A3(n1062), .A4(n1082), .ZN(n1024) );
AND2_X1 U782 ( .A1(n1068), .A2(n1057), .ZN(n1082) );
INV_X1 U783 ( .A(n1083), .ZN(n1057) );
OR2_X1 U784 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
XOR2_X1 U785 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U786 ( .A1(n1088), .A2(n1027), .ZN(n1087) );
AND2_X1 U787 ( .A1(G227), .A2(G900), .ZN(n1088) );
NAND2_X1 U788 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND3_X1 U789 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NAND2_X1 U790 ( .A1(G953), .A2(n1094), .ZN(n1092) );
OR2_X1 U791 ( .A1(n1091), .A2(n1093), .ZN(n1089) );
NAND2_X1 U792 ( .A1(n1027), .A2(n1095), .ZN(n1093) );
NAND2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U794 ( .A(KEYINPUT3), .B(n1023), .ZN(n1097) );
INV_X1 U795 ( .A(n1021), .ZN(n1096) );
XOR2_X1 U796 ( .A(n1098), .B(n1099), .Z(n1091) );
XOR2_X1 U797 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U798 ( .A(G134), .B(G131), .Z(n1101) );
NOR2_X1 U799 ( .A1(G137), .A2(KEYINPUT8), .ZN(n1100) );
XNOR2_X1 U800 ( .A(n1102), .B(n1103), .ZN(n1098) );
NOR2_X1 U801 ( .A1(KEYINPUT49), .A2(n1104), .ZN(n1103) );
XNOR2_X1 U802 ( .A(n1105), .B(n1106), .ZN(n1104) );
NOR2_X1 U803 ( .A1(KEYINPUT60), .A2(G125), .ZN(n1106) );
XOR2_X1 U804 ( .A(n1107), .B(n1108), .Z(G69) );
NOR3_X1 U805 ( .A1(n1022), .A2(n1109), .A3(n1110), .ZN(n1108) );
NOR2_X1 U806 ( .A1(G224), .A2(n1027), .ZN(n1110) );
NAND2_X1 U807 ( .A1(n1111), .A2(n1112), .ZN(n1107) );
INV_X1 U808 ( .A(n1109), .ZN(n1112) );
XOR2_X1 U809 ( .A(n1113), .B(n1114), .Z(n1111) );
XOR2_X1 U810 ( .A(KEYINPUT21), .B(n1115), .Z(n1114) );
XNOR2_X1 U811 ( .A(n1116), .B(n1117), .ZN(n1113) );
NOR2_X1 U812 ( .A1(n1118), .A2(n1119), .ZN(G66) );
XOR2_X1 U813 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U814 ( .A1(n1122), .A2(n1036), .ZN(n1120) );
INV_X1 U815 ( .A(n1123), .ZN(n1036) );
NOR2_X1 U816 ( .A1(n1118), .A2(n1124), .ZN(G63) );
XOR2_X1 U817 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U818 ( .A1(n1122), .A2(G478), .ZN(n1125) );
NOR2_X1 U819 ( .A1(n1118), .A2(n1127), .ZN(G60) );
XOR2_X1 U820 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U821 ( .A(n1130), .B(KEYINPUT30), .Z(n1128) );
NAND2_X1 U822 ( .A1(n1122), .A2(G475), .ZN(n1130) );
XNOR2_X1 U823 ( .A(G104), .B(n1131), .ZN(G6) );
NOR2_X1 U824 ( .A1(n1118), .A2(n1132), .ZN(G57) );
XOR2_X1 U825 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U826 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U827 ( .A1(G101), .A2(KEYINPUT42), .ZN(n1136) );
NAND3_X1 U828 ( .A1(n1137), .A2(n1138), .A3(KEYINPUT12), .ZN(n1135) );
XNOR2_X1 U829 ( .A(n1139), .B(n1140), .ZN(n1133) );
NAND2_X1 U830 ( .A1(n1122), .A2(G472), .ZN(n1139) );
NOR2_X1 U831 ( .A1(n1118), .A2(n1141), .ZN(G54) );
XOR2_X1 U832 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U833 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U834 ( .A(n1102), .B(n1146), .ZN(n1145) );
XOR2_X1 U835 ( .A(n1147), .B(n1148), .Z(n1142) );
XOR2_X1 U836 ( .A(n1149), .B(KEYINPUT47), .Z(n1148) );
NAND2_X1 U837 ( .A1(n1122), .A2(G469), .ZN(n1147) );
NOR2_X1 U838 ( .A1(n1118), .A2(n1150), .ZN(G51) );
XOR2_X1 U839 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U840 ( .A(n1153), .B(n1154), .ZN(n1152) );
XOR2_X1 U841 ( .A(n1155), .B(n1156), .Z(n1151) );
NAND2_X1 U842 ( .A1(n1122), .A2(n1041), .ZN(n1155) );
AND2_X1 U843 ( .A1(G902), .A2(n1157), .ZN(n1122) );
OR3_X1 U844 ( .A1(n1023), .A2(n1022), .A3(n1021), .ZN(n1157) );
NAND4_X1 U845 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1021) );
NAND4_X1 U846 ( .A1(n1131), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1022) );
NOR4_X1 U847 ( .A1(n1165), .A2(n1016), .A3(n1166), .A4(n1167), .ZN(n1164) );
AND3_X1 U848 ( .A1(n1060), .A2(n1085), .A3(n1168), .ZN(n1016) );
NAND2_X1 U849 ( .A1(n1169), .A2(n1170), .ZN(n1163) );
NAND2_X1 U850 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
XOR2_X1 U851 ( .A(n1085), .B(KEYINPUT29), .Z(n1172) );
NAND3_X1 U852 ( .A1(n1060), .A2(n1084), .A3(n1168), .ZN(n1131) );
NAND4_X1 U853 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1023) );
NAND2_X1 U854 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
INV_X1 U855 ( .A(KEYINPUT15), .ZN(n1178) );
NAND3_X1 U856 ( .A1(n1179), .A2(n1180), .A3(KEYINPUT15), .ZN(n1175) );
NAND2_X1 U857 ( .A1(n1181), .A2(n1085), .ZN(n1174) );
NAND3_X1 U858 ( .A1(n1073), .A2(n1182), .A3(n1183), .ZN(n1173) );
NAND2_X1 U859 ( .A1(n1171), .A2(n1184), .ZN(n1182) );
XOR2_X1 U860 ( .A(n1085), .B(KEYINPUT17), .Z(n1184) );
NOR2_X1 U861 ( .A1(n1027), .A2(G952), .ZN(n1118) );
XNOR2_X1 U862 ( .A(n1161), .B(n1185), .ZN(G48) );
NOR2_X1 U863 ( .A1(KEYINPUT14), .A2(n1186), .ZN(n1185) );
NAND2_X1 U864 ( .A1(n1181), .A2(n1084), .ZN(n1161) );
NAND2_X1 U865 ( .A1(n1187), .A2(n1188), .ZN(G45) );
NAND2_X1 U866 ( .A1(n1189), .A2(n1158), .ZN(n1188) );
NAND2_X1 U867 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U868 ( .A1(KEYINPUT33), .A2(n1192), .ZN(n1191) );
NAND3_X1 U869 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1187) );
INV_X1 U870 ( .A(KEYINPUT33), .ZN(n1195) );
NAND2_X1 U871 ( .A1(G143), .A2(n1192), .ZN(n1194) );
INV_X1 U872 ( .A(KEYINPUT13), .ZN(n1192) );
NAND2_X1 U873 ( .A1(n1196), .A2(n1190), .ZN(n1193) );
OR2_X1 U874 ( .A1(n1158), .A2(KEYINPUT13), .ZN(n1196) );
NAND4_X1 U875 ( .A1(n1197), .A2(n1073), .A3(n1198), .A4(n1199), .ZN(n1158) );
XNOR2_X1 U876 ( .A(G140), .B(n1159), .ZN(G42) );
NAND2_X1 U877 ( .A1(n1200), .A2(n1183), .ZN(n1159) );
XNOR2_X1 U878 ( .A(G137), .B(n1160), .ZN(G39) );
NAND3_X1 U879 ( .A1(n1201), .A2(n1202), .A3(n1183), .ZN(n1160) );
INV_X1 U880 ( .A(n1203), .ZN(n1183) );
NAND2_X1 U881 ( .A1(n1204), .A2(n1205), .ZN(G36) );
NAND2_X1 U882 ( .A1(KEYINPUT24), .A2(G134), .ZN(n1205) );
XOR2_X1 U883 ( .A(n1206), .B(n1207), .Z(n1204) );
NOR2_X1 U884 ( .A1(n1203), .A2(n1208), .ZN(n1207) );
NOR2_X1 U885 ( .A1(G134), .A2(KEYINPUT24), .ZN(n1206) );
XOR2_X1 U886 ( .A(G131), .B(n1209), .Z(G33) );
NOR4_X1 U887 ( .A1(KEYINPUT46), .A2(n1171), .A3(n1210), .A4(n1203), .ZN(n1209) );
NAND3_X1 U888 ( .A1(n1067), .A2(n1211), .A3(n1062), .ZN(n1203) );
NOR2_X1 U889 ( .A1(n1212), .A2(n1079), .ZN(n1062) );
INV_X1 U890 ( .A(n1073), .ZN(n1210) );
INV_X1 U891 ( .A(n1084), .ZN(n1171) );
XNOR2_X1 U892 ( .A(G128), .B(n1213), .ZN(G30) );
NAND3_X1 U893 ( .A1(n1181), .A2(n1085), .A3(KEYINPUT27), .ZN(n1213) );
AND3_X1 U894 ( .A1(n1075), .A2(n1202), .A3(n1197), .ZN(n1181) );
AND3_X1 U895 ( .A1(n1067), .A2(n1211), .A3(n1179), .ZN(n1197) );
XNOR2_X1 U896 ( .A(n1214), .B(n1165), .ZN(G3) );
AND3_X1 U897 ( .A1(n1168), .A2(n1055), .A3(n1073), .ZN(n1165) );
XOR2_X1 U898 ( .A(n1177), .B(n1215), .Z(G27) );
NOR2_X1 U899 ( .A1(KEYINPUT34), .A2(n1216), .ZN(n1215) );
NOR2_X1 U900 ( .A1(n1180), .A2(n1077), .ZN(n1177) );
INV_X1 U901 ( .A(n1179), .ZN(n1077) );
NAND3_X1 U902 ( .A1(n1068), .A2(n1211), .A3(n1200), .ZN(n1180) );
AND3_X1 U903 ( .A1(n1084), .A2(n1075), .A3(n1030), .ZN(n1200) );
NAND2_X1 U904 ( .A1(n1083), .A2(n1217), .ZN(n1211) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1218), .A4(n1094), .ZN(n1217) );
INV_X1 U906 ( .A(G900), .ZN(n1094) );
XNOR2_X1 U907 ( .A(G122), .B(n1162), .ZN(G24) );
NAND4_X1 U908 ( .A1(n1219), .A2(n1060), .A3(n1198), .A4(n1199), .ZN(n1162) );
NOR2_X1 U909 ( .A1(n1202), .A2(n1075), .ZN(n1060) );
XNOR2_X1 U910 ( .A(n1167), .B(n1220), .ZN(G21) );
XOR2_X1 U911 ( .A(KEYINPUT38), .B(G119), .Z(n1220) );
AND3_X1 U912 ( .A1(n1201), .A2(n1202), .A3(n1219), .ZN(n1167) );
XOR2_X1 U913 ( .A(n1221), .B(n1222), .Z(G18) );
NOR2_X1 U914 ( .A1(KEYINPUT36), .A2(n1223), .ZN(n1222) );
NAND2_X1 U915 ( .A1(n1224), .A2(n1225), .ZN(n1221) );
NAND3_X1 U916 ( .A1(n1179), .A2(n1226), .A3(n1227), .ZN(n1225) );
INV_X1 U917 ( .A(KEYINPUT2), .ZN(n1227) );
NAND2_X1 U918 ( .A1(n1228), .A2(n1229), .ZN(n1226) );
INV_X1 U919 ( .A(n1208), .ZN(n1228) );
NAND2_X1 U920 ( .A1(n1073), .A2(n1085), .ZN(n1208) );
NAND3_X1 U921 ( .A1(n1169), .A2(n1085), .A3(KEYINPUT2), .ZN(n1224) );
NAND2_X1 U922 ( .A1(n1230), .A2(n1231), .ZN(n1085) );
OR3_X1 U923 ( .A1(n1199), .A2(n1054), .A3(KEYINPUT1), .ZN(n1231) );
NAND2_X1 U924 ( .A1(KEYINPUT1), .A2(n1055), .ZN(n1230) );
XOR2_X1 U925 ( .A(n1232), .B(n1233), .Z(G15) );
NOR2_X1 U926 ( .A1(KEYINPUT53), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U927 ( .A(G113), .B(KEYINPUT10), .ZN(n1234) );
NAND2_X1 U928 ( .A1(n1169), .A2(n1084), .ZN(n1232) );
NAND2_X1 U929 ( .A1(n1235), .A2(n1236), .ZN(n1084) );
NAND2_X1 U930 ( .A1(n1055), .A2(n1237), .ZN(n1236) );
INV_X1 U931 ( .A(KEYINPUT52), .ZN(n1237) );
NAND3_X1 U932 ( .A1(n1054), .A2(n1199), .A3(KEYINPUT52), .ZN(n1235) );
INV_X1 U933 ( .A(n1198), .ZN(n1054) );
AND2_X1 U934 ( .A1(n1219), .A2(n1073), .ZN(n1169) );
NOR2_X1 U935 ( .A1(n1075), .A2(n1030), .ZN(n1073) );
AND2_X1 U936 ( .A1(n1229), .A2(n1179), .ZN(n1219) );
AND2_X1 U937 ( .A1(n1068), .A2(n1238), .ZN(n1229) );
NOR2_X1 U938 ( .A1(n1239), .A2(n1065), .ZN(n1068) );
XOR2_X1 U939 ( .A(G110), .B(n1166), .Z(G12) );
AND3_X1 U940 ( .A1(n1030), .A2(n1168), .A3(n1201), .ZN(n1166) );
AND2_X1 U941 ( .A1(n1055), .A2(n1075), .ZN(n1201) );
XOR2_X1 U942 ( .A(n1039), .B(n1123), .Z(n1075) );
NAND2_X1 U943 ( .A1(G217), .A2(n1240), .ZN(n1123) );
NAND2_X1 U944 ( .A1(n1241), .A2(n1121), .ZN(n1039) );
XNOR2_X1 U945 ( .A(n1242), .B(n1243), .ZN(n1121) );
XOR2_X1 U946 ( .A(G119), .B(n1244), .Z(n1243) );
XNOR2_X1 U947 ( .A(G137), .B(n1216), .ZN(n1244) );
INV_X1 U948 ( .A(G125), .ZN(n1216) );
XOR2_X1 U949 ( .A(n1245), .B(n1246), .Z(n1242) );
XNOR2_X1 U950 ( .A(n1247), .B(n1248), .ZN(n1245) );
AND2_X1 U951 ( .A1(G221), .A2(n1249), .ZN(n1248) );
NOR2_X1 U952 ( .A1(n1199), .A2(n1198), .ZN(n1055) );
XNOR2_X1 U953 ( .A(n1250), .B(n1251), .ZN(n1198) );
XOR2_X1 U954 ( .A(KEYINPUT40), .B(G478), .Z(n1251) );
NAND2_X1 U955 ( .A1(n1241), .A2(n1126), .ZN(n1250) );
XNOR2_X1 U956 ( .A(n1252), .B(n1253), .ZN(n1126) );
XOR2_X1 U957 ( .A(n1254), .B(n1255), .Z(n1253) );
NOR2_X1 U958 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U959 ( .A(n1258), .B(KEYINPUT48), .Z(n1257) );
NAND2_X1 U960 ( .A1(G107), .A2(n1259), .ZN(n1258) );
NOR2_X1 U961 ( .A1(G107), .A2(n1259), .ZN(n1256) );
XNOR2_X1 U962 ( .A(n1223), .B(n1260), .ZN(n1259) );
XOR2_X1 U963 ( .A(KEYINPUT37), .B(G122), .Z(n1260) );
NOR2_X1 U964 ( .A1(KEYINPUT16), .A2(n1261), .ZN(n1254) );
XOR2_X1 U965 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U966 ( .A(G128), .B(G134), .ZN(n1263) );
NAND2_X1 U967 ( .A1(KEYINPUT26), .A2(n1190), .ZN(n1262) );
NAND2_X1 U968 ( .A1(G217), .A2(n1249), .ZN(n1252) );
AND2_X1 U969 ( .A1(G234), .A2(n1027), .ZN(n1249) );
NAND2_X1 U970 ( .A1(n1044), .A2(n1264), .ZN(n1199) );
OR2_X1 U971 ( .A1(n1051), .A2(n1050), .ZN(n1264) );
NAND2_X1 U972 ( .A1(n1050), .A2(n1051), .ZN(n1044) );
INV_X1 U973 ( .A(G475), .ZN(n1051) );
NOR2_X1 U974 ( .A1(n1129), .A2(n1265), .ZN(n1050) );
XNOR2_X1 U975 ( .A(n1266), .B(n1267), .ZN(n1129) );
XOR2_X1 U976 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U977 ( .A(n1270), .B(KEYINPUT45), .ZN(n1269) );
NAND2_X1 U978 ( .A1(n1271), .A2(KEYINPUT20), .ZN(n1270) );
XOR2_X1 U979 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U980 ( .A(n1190), .B(G131), .ZN(n1273) );
INV_X1 U981 ( .A(G143), .ZN(n1190) );
NAND3_X1 U982 ( .A1(n1274), .A2(n1027), .A3(G214), .ZN(n1272) );
XNOR2_X1 U983 ( .A(KEYINPUT58), .B(n1275), .ZN(n1274) );
NOR2_X1 U984 ( .A1(G104), .A2(KEYINPUT39), .ZN(n1268) );
XOR2_X1 U985 ( .A(n1276), .B(n1115), .Z(n1266) );
XOR2_X1 U986 ( .A(G113), .B(G122), .Z(n1115) );
NAND2_X1 U987 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U988 ( .A1(n1279), .A2(G146), .ZN(n1278) );
XOR2_X1 U989 ( .A(KEYINPUT55), .B(n1280), .Z(n1277) );
NOR2_X1 U990 ( .A1(G146), .A2(n1279), .ZN(n1280) );
XNOR2_X1 U991 ( .A(G125), .B(n1281), .ZN(n1279) );
NOR2_X1 U992 ( .A1(KEYINPUT25), .A2(n1105), .ZN(n1281) );
AND3_X1 U993 ( .A1(n1067), .A2(n1238), .A3(n1179), .ZN(n1168) );
NOR2_X1 U994 ( .A1(n1080), .A2(n1079), .ZN(n1179) );
INV_X1 U995 ( .A(n1043), .ZN(n1079) );
NAND2_X1 U996 ( .A1(G214), .A2(n1282), .ZN(n1043) );
INV_X1 U997 ( .A(n1212), .ZN(n1080) );
XNOR2_X1 U998 ( .A(n1042), .B(n1041), .ZN(n1212) );
AND2_X1 U999 ( .A1(G210), .A2(n1282), .ZN(n1041) );
NAND2_X1 U1000 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U1001 ( .A1(n1285), .A2(n1241), .ZN(n1042) );
XNOR2_X1 U1002 ( .A(n1286), .B(n1287), .ZN(n1285) );
INV_X1 U1003 ( .A(n1153), .ZN(n1287) );
XNOR2_X1 U1004 ( .A(n1288), .B(n1289), .ZN(n1153) );
XNOR2_X1 U1005 ( .A(G122), .B(n1290), .ZN(n1289) );
XNOR2_X1 U1006 ( .A(KEYINPUT61), .B(KEYINPUT43), .ZN(n1290) );
XNOR2_X1 U1007 ( .A(n1291), .B(n1292), .ZN(n1288) );
INV_X1 U1008 ( .A(n1116), .ZN(n1292) );
XNOR2_X1 U1009 ( .A(n1146), .B(G110), .ZN(n1116) );
NAND2_X1 U1010 ( .A1(n1293), .A2(KEYINPUT56), .ZN(n1291) );
XNOR2_X1 U1011 ( .A(G113), .B(n1117), .ZN(n1293) );
NAND3_X1 U1012 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(n1286) );
NAND2_X1 U1013 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
NAND3_X1 U1014 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1298) );
NAND2_X1 U1015 ( .A1(KEYINPUT18), .A2(n1302), .ZN(n1301) );
NAND2_X1 U1016 ( .A1(KEYINPUT22), .A2(n1156), .ZN(n1300) );
NAND2_X1 U1017 ( .A1(n1303), .A2(n1304), .ZN(n1299) );
INV_X1 U1018 ( .A(KEYINPUT22), .ZN(n1304) );
NAND2_X1 U1019 ( .A1(n1156), .A2(n1305), .ZN(n1303) );
NAND2_X1 U1020 ( .A1(KEYINPUT28), .A2(n1306), .ZN(n1305) );
NAND4_X1 U1021 ( .A1(n1154), .A2(n1156), .A3(KEYINPUT18), .A4(KEYINPUT28), .ZN(n1295) );
NAND2_X1 U1022 ( .A1(n1307), .A2(n1302), .ZN(n1294) );
INV_X1 U1023 ( .A(KEYINPUT28), .ZN(n1302) );
NAND2_X1 U1024 ( .A1(n1156), .A2(n1308), .ZN(n1307) );
NAND2_X1 U1025 ( .A1(n1154), .A2(n1306), .ZN(n1308) );
INV_X1 U1026 ( .A(KEYINPUT18), .ZN(n1306) );
INV_X1 U1027 ( .A(n1297), .ZN(n1154) );
XNOR2_X1 U1028 ( .A(G125), .B(n1309), .ZN(n1297) );
AND2_X1 U1029 ( .A1(G224), .A2(n1027), .ZN(n1156) );
NAND2_X1 U1030 ( .A1(n1083), .A2(n1310), .ZN(n1238) );
NAND3_X1 U1031 ( .A1(G902), .A2(n1218), .A3(n1109), .ZN(n1310) );
NOR2_X1 U1032 ( .A1(G898), .A2(n1027), .ZN(n1109) );
NAND3_X1 U1033 ( .A1(n1218), .A2(n1027), .A3(G952), .ZN(n1083) );
NAND2_X1 U1034 ( .A1(G237), .A2(G234), .ZN(n1218) );
NOR2_X1 U1035 ( .A1(n1066), .A2(n1065), .ZN(n1067) );
INV_X1 U1036 ( .A(n1045), .ZN(n1065) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1240), .ZN(n1045) );
NAND2_X1 U1038 ( .A1(G234), .A2(n1284), .ZN(n1240) );
INV_X1 U1039 ( .A(G902), .ZN(n1284) );
INV_X1 U1040 ( .A(n1239), .ZN(n1066) );
XOR2_X1 U1041 ( .A(G469), .B(n1311), .Z(n1239) );
NOR2_X1 U1042 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
AND2_X1 U1043 ( .A1(KEYINPUT41), .A2(n1052), .ZN(n1313) );
NOR2_X1 U1044 ( .A1(KEYINPUT6), .A2(n1052), .ZN(n1312) );
NAND2_X1 U1045 ( .A1(n1314), .A2(n1241), .ZN(n1052) );
XOR2_X1 U1046 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1047 ( .A(n1317), .B(n1144), .Z(n1316) );
XNOR2_X1 U1048 ( .A(n1318), .B(n1247), .ZN(n1144) );
XNOR2_X1 U1049 ( .A(G110), .B(n1319), .ZN(n1247) );
INV_X1 U1050 ( .A(n1105), .ZN(n1319) );
XOR2_X1 U1051 ( .A(G140), .B(KEYINPUT11), .Z(n1105) );
NOR2_X1 U1052 ( .A1(KEYINPUT63), .A2(n1149), .ZN(n1317) );
NAND2_X1 U1053 ( .A1(G227), .A2(n1027), .ZN(n1149) );
XNOR2_X1 U1054 ( .A(KEYINPUT35), .B(n1320), .ZN(n1315) );
NOR2_X1 U1055 ( .A1(KEYINPUT44), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1056 ( .A(n1322), .B(n1146), .Z(n1321) );
XNOR2_X1 U1057 ( .A(G101), .B(n1323), .ZN(n1146) );
XOR2_X1 U1058 ( .A(G107), .B(G104), .Z(n1323) );
NAND2_X1 U1059 ( .A1(KEYINPUT9), .A2(n1102), .ZN(n1322) );
INV_X1 U1060 ( .A(n1202), .ZN(n1030) );
XNOR2_X1 U1061 ( .A(n1324), .B(G472), .ZN(n1202) );
NAND2_X1 U1062 ( .A1(n1241), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1063 ( .A(n1326), .B(n1327), .Z(n1325) );
NAND2_X1 U1064 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U1065 ( .A1(n1140), .A2(n1214), .ZN(n1329) );
XOR2_X1 U1066 ( .A(KEYINPUT4), .B(n1330), .Z(n1328) );
NOR2_X1 U1067 ( .A1(n1214), .A2(n1140), .ZN(n1330) );
NAND3_X1 U1068 ( .A1(G210), .A2(n1027), .A3(n1275), .ZN(n1140) );
XOR2_X1 U1069 ( .A(n1283), .B(KEYINPUT5), .Z(n1275) );
INV_X1 U1070 ( .A(G237), .ZN(n1283) );
INV_X1 U1071 ( .A(G953), .ZN(n1027) );
INV_X1 U1072 ( .A(G101), .ZN(n1214) );
NAND3_X1 U1073 ( .A1(n1331), .A2(n1332), .A3(n1138), .ZN(n1326) );
NAND2_X1 U1074 ( .A1(n1333), .A2(n1318), .ZN(n1138) );
NAND2_X1 U1075 ( .A1(KEYINPUT19), .A2(n1334), .ZN(n1332) );
NAND3_X1 U1076 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
INV_X1 U1077 ( .A(n1333), .ZN(n1337) );
NOR2_X1 U1078 ( .A1(n1338), .A2(n1309), .ZN(n1333) );
NAND2_X1 U1079 ( .A1(n1339), .A2(n1318), .ZN(n1336) );
NAND3_X1 U1080 ( .A1(n1338), .A2(n1309), .A3(n1340), .ZN(n1335) );
OR2_X1 U1081 ( .A1(n1137), .A2(KEYINPUT19), .ZN(n1331) );
AND2_X1 U1082 ( .A1(n1341), .A2(n1342), .ZN(n1137) );
NAND2_X1 U1083 ( .A1(n1343), .A2(n1309), .ZN(n1342) );
INV_X1 U1084 ( .A(n1102), .ZN(n1309) );
XNOR2_X1 U1085 ( .A(n1340), .B(n1339), .ZN(n1343) );
INV_X1 U1086 ( .A(n1338), .ZN(n1339) );
NAND3_X1 U1087 ( .A1(n1340), .A2(n1338), .A3(n1102), .ZN(n1341) );
XOR2_X1 U1088 ( .A(G143), .B(n1246), .Z(n1102) );
XNOR2_X1 U1089 ( .A(G128), .B(n1186), .ZN(n1246) );
INV_X1 U1090 ( .A(G146), .ZN(n1186) );
XNOR2_X1 U1091 ( .A(n1344), .B(n1117), .ZN(n1338) );
XNOR2_X1 U1092 ( .A(n1223), .B(G119), .ZN(n1117) );
INV_X1 U1093 ( .A(G116), .ZN(n1223) );
NAND2_X1 U1094 ( .A1(KEYINPUT62), .A2(G113), .ZN(n1344) );
INV_X1 U1095 ( .A(n1318), .ZN(n1340) );
NAND3_X1 U1096 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1318) );
NAND2_X1 U1097 ( .A1(KEYINPUT51), .A2(n1348), .ZN(n1347) );
INV_X1 U1098 ( .A(n1349), .ZN(n1348) );
OR3_X1 U1099 ( .A1(n1350), .A2(KEYINPUT51), .A3(G131), .ZN(n1346) );
NAND2_X1 U1100 ( .A1(G131), .A2(n1350), .ZN(n1345) );
NAND2_X1 U1101 ( .A1(KEYINPUT59), .A2(n1349), .ZN(n1350) );
XOR2_X1 U1102 ( .A(G134), .B(G137), .Z(n1349) );
INV_X1 U1103 ( .A(n1265), .ZN(n1241) );
XOR2_X1 U1104 ( .A(G902), .B(KEYINPUT23), .Z(n1265) );
endmodule


