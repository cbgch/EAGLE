//Key = 1100011000000110101000111101100001001111010000111110010001101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359;

XNOR2_X1 U734 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U735 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U736 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NOR2_X1 U737 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U738 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U739 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
INV_X1 U740 ( .A(KEYINPUT12), .ZN(n1040) );
NOR4_X1 U741 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1039) );
NOR2_X1 U742 ( .A1(n1045), .A2(n1044), .ZN(n1037) );
NOR2_X1 U743 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U744 ( .A1(n1048), .A2(n1042), .ZN(n1047) );
NOR2_X1 U745 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U747 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U748 ( .A1(n1055), .A2(n1041), .ZN(n1049) );
NOR2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U750 ( .A1(KEYINPUT12), .A2(n1043), .ZN(n1056) );
NOR3_X1 U751 ( .A1(n1052), .A2(n1058), .A3(n1041), .ZN(n1046) );
NAND3_X1 U752 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1031) );
NAND4_X1 U753 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
NAND2_X1 U754 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U755 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
INV_X1 U756 ( .A(n1036), .ZN(n1069) );
NAND2_X1 U757 ( .A1(n1071), .A2(n1072), .ZN(n1066) );
NAND2_X1 U758 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U759 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
INV_X1 U760 ( .A(n1044), .ZN(n1062) );
NOR3_X1 U761 ( .A1(n1077), .A2(G953), .A3(n1078), .ZN(n1029) );
INV_X1 U762 ( .A(n1059), .ZN(n1078) );
NAND3_X1 U763 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1059) );
NOR3_X1 U764 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
XOR2_X1 U765 ( .A(n1085), .B(KEYINPUT63), .Z(n1083) );
NAND3_X1 U766 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
OR2_X1 U767 ( .A1(G478), .A2(KEYINPUT36), .ZN(n1087) );
NAND3_X1 U768 ( .A1(G478), .A2(n1089), .A3(KEYINPUT36), .ZN(n1086) );
XOR2_X1 U769 ( .A(n1090), .B(KEYINPUT46), .Z(n1080) );
NAND3_X1 U770 ( .A1(n1091), .A2(n1092), .A3(n1071), .ZN(n1090) );
XOR2_X1 U771 ( .A(n1093), .B(G472), .Z(n1079) );
XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n1034), .ZN(n1077) );
XOR2_X1 U773 ( .A(n1094), .B(n1095), .Z(G72) );
XOR2_X1 U774 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U775 ( .A1(G953), .A2(n1098), .ZN(n1097) );
NAND2_X1 U776 ( .A1(G900), .A2(G227), .ZN(n1098) );
NAND2_X1 U777 ( .A1(n1099), .A2(n1100), .ZN(n1096) );
INV_X1 U778 ( .A(n1101), .ZN(n1100) );
XOR2_X1 U779 ( .A(n1102), .B(n1103), .Z(n1099) );
XOR2_X1 U780 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U781 ( .A(KEYINPUT2), .B(G131), .Z(n1105) );
NOR2_X1 U782 ( .A1(KEYINPUT20), .A2(n1106), .ZN(n1104) );
XOR2_X1 U783 ( .A(n1107), .B(KEYINPUT3), .Z(n1106) );
XNOR2_X1 U784 ( .A(n1108), .B(n1109), .ZN(n1102) );
NOR2_X1 U785 ( .A1(n1110), .A2(G953), .ZN(n1094) );
XOR2_X1 U786 ( .A(n1111), .B(n1112), .Z(G69) );
NOR2_X1 U787 ( .A1(KEYINPUT45), .A2(n1113), .ZN(n1112) );
XOR2_X1 U788 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U789 ( .A1(n1116), .A2(G953), .ZN(n1115) );
NOR2_X1 U790 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
XOR2_X1 U791 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U792 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
XOR2_X1 U793 ( .A(n1123), .B(KEYINPUT55), .Z(n1121) );
NOR2_X1 U794 ( .A1(G898), .A2(n1060), .ZN(n1117) );
NAND2_X1 U795 ( .A1(G953), .A2(n1124), .ZN(n1111) );
NAND2_X1 U796 ( .A1(G898), .A2(G224), .ZN(n1124) );
NOR2_X1 U797 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XOR2_X1 U798 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U799 ( .A1(KEYINPUT30), .A2(n1129), .ZN(n1128) );
NAND2_X1 U800 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
NOR2_X1 U801 ( .A1(n1125), .A2(n1132), .ZN(G63) );
XOR2_X1 U802 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U803 ( .A(KEYINPUT54), .B(n1135), .Z(n1134) );
NOR2_X1 U804 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR3_X1 U805 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(G60) );
NOR3_X1 U806 ( .A1(n1141), .A2(G952), .A3(n1142), .ZN(n1140) );
INV_X1 U807 ( .A(KEYINPUT7), .ZN(n1141) );
NOR2_X1 U808 ( .A1(KEYINPUT7), .A2(n1143), .ZN(n1139) );
XNOR2_X1 U809 ( .A(n1144), .B(n1145), .ZN(n1138) );
AND2_X1 U810 ( .A1(G475), .A2(n1130), .ZN(n1144) );
XNOR2_X1 U811 ( .A(G104), .B(n1146), .ZN(G6) );
NOR2_X1 U812 ( .A1(n1125), .A2(n1147), .ZN(G57) );
XOR2_X1 U813 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U814 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U815 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U816 ( .A(n1154), .B(KEYINPUT13), .Z(n1153) );
NOR2_X1 U817 ( .A1(n1155), .A2(n1154), .ZN(n1150) );
XOR2_X1 U818 ( .A(n1156), .B(n1157), .Z(n1148) );
NAND3_X1 U819 ( .A1(n1130), .A2(G472), .A3(KEYINPUT62), .ZN(n1156) );
NOR2_X1 U820 ( .A1(n1125), .A2(n1158), .ZN(G54) );
XOR2_X1 U821 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U822 ( .A1(G469), .A2(n1130), .ZN(n1160) );
INV_X1 U823 ( .A(n1137), .ZN(n1130) );
NAND2_X1 U824 ( .A1(KEYINPUT23), .A2(n1161), .ZN(n1159) );
XOR2_X1 U825 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U826 ( .A(n1164), .B(n1165), .ZN(n1163) );
XOR2_X1 U827 ( .A(n1166), .B(n1167), .Z(n1162) );
NOR2_X1 U828 ( .A1(KEYINPUT32), .A2(n1168), .ZN(n1167) );
XOR2_X1 U829 ( .A(G110), .B(n1169), .Z(n1168) );
XNOR2_X1 U830 ( .A(KEYINPUT57), .B(n1170), .ZN(n1169) );
INV_X1 U831 ( .A(G140), .ZN(n1170) );
NOR2_X1 U832 ( .A1(n1125), .A2(n1171), .ZN(G51) );
XOR2_X1 U833 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U834 ( .A1(n1174), .A2(n1137), .ZN(n1173) );
NAND2_X1 U835 ( .A1(n1175), .A2(n1032), .ZN(n1137) );
NAND2_X1 U836 ( .A1(n1110), .A2(n1116), .ZN(n1032) );
AND4_X1 U837 ( .A1(n1028), .A2(n1146), .A3(n1176), .A4(n1177), .ZN(n1116) );
NOR4_X1 U838 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR3_X1 U839 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1181) );
NOR3_X1 U840 ( .A1(n1052), .A2(n1053), .A3(n1185), .ZN(n1184) );
NOR2_X1 U841 ( .A1(KEYINPUT21), .A2(n1186), .ZN(n1185) );
INV_X1 U842 ( .A(n1054), .ZN(n1186) );
NOR2_X1 U843 ( .A1(n1063), .A2(n1187), .ZN(n1183) );
AND2_X1 U844 ( .A1(n1054), .A2(KEYINPUT21), .ZN(n1187) );
NOR2_X1 U845 ( .A1(n1188), .A2(n1189), .ZN(n1180) );
XNOR2_X1 U846 ( .A(KEYINPUT28), .B(n1190), .ZN(n1189) );
NOR2_X1 U847 ( .A1(n1191), .A2(n1192), .ZN(n1179) );
AND4_X1 U848 ( .A1(n1191), .A2(n1193), .A3(n1190), .A4(n1057), .ZN(n1178) );
INV_X1 U849 ( .A(KEYINPUT61), .ZN(n1191) );
NOR2_X1 U850 ( .A1(n1194), .A2(n1195), .ZN(n1176) );
NAND3_X1 U851 ( .A1(n1196), .A2(n1064), .A3(n1197), .ZN(n1146) );
NAND3_X1 U852 ( .A1(n1196), .A2(n1064), .A3(n1057), .ZN(n1028) );
AND4_X1 U853 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1110) );
NOR4_X1 U854 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
INV_X1 U855 ( .A(n1206), .ZN(n1205) );
INV_X1 U856 ( .A(n1207), .ZN(n1202) );
AND2_X1 U857 ( .A1(n1208), .A2(n1209), .ZN(n1200) );
XNOR2_X1 U858 ( .A(KEYINPUT10), .B(n1210), .ZN(n1175) );
NOR3_X1 U859 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1172) );
NOR2_X1 U860 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U861 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
XOR2_X1 U862 ( .A(n1218), .B(KEYINPUT26), .Z(n1216) );
NOR3_X1 U863 ( .A1(n1219), .A2(n1218), .A3(n1217), .ZN(n1212) );
AND2_X1 U864 ( .A1(n1217), .A2(n1218), .ZN(n1211) );
NAND2_X1 U865 ( .A1(n1220), .A2(n1221), .ZN(n1218) );
OR2_X1 U866 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U867 ( .A(n1224), .B(KEYINPUT40), .Z(n1220) );
NAND2_X1 U868 ( .A1(n1222), .A2(n1223), .ZN(n1224) );
INV_X1 U869 ( .A(KEYINPUT14), .ZN(n1217) );
INV_X1 U870 ( .A(n1143), .ZN(n1125) );
NAND2_X1 U871 ( .A1(n1142), .A2(n1034), .ZN(n1143) );
INV_X1 U872 ( .A(G952), .ZN(n1034) );
XNOR2_X1 U873 ( .A(G953), .B(KEYINPUT53), .ZN(n1142) );
XOR2_X1 U874 ( .A(n1209), .B(n1225), .Z(G48) );
XNOR2_X1 U875 ( .A(KEYINPUT41), .B(n1226), .ZN(n1225) );
NAND3_X1 U876 ( .A1(n1197), .A2(n1227), .A3(n1228), .ZN(n1209) );
XNOR2_X1 U877 ( .A(n1229), .B(n1230), .ZN(G45) );
NAND2_X1 U878 ( .A1(KEYINPUT49), .A2(n1208), .ZN(n1229) );
NAND4_X1 U879 ( .A1(n1231), .A2(n1227), .A3(n1053), .A4(n1232), .ZN(n1208) );
NOR3_X1 U880 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1232) );
XNOR2_X1 U881 ( .A(G140), .B(n1198), .ZN(G42) );
NAND3_X1 U882 ( .A1(n1197), .A2(n1054), .A3(n1236), .ZN(n1198) );
XNOR2_X1 U883 ( .A(G137), .B(n1199), .ZN(G39) );
NAND4_X1 U884 ( .A1(n1063), .A2(n1236), .A3(n1237), .A4(n1082), .ZN(n1199) );
XNOR2_X1 U885 ( .A(G134), .B(n1238), .ZN(G36) );
NOR2_X1 U886 ( .A1(n1204), .A2(KEYINPUT43), .ZN(n1238) );
AND3_X1 U887 ( .A1(n1236), .A2(n1057), .A3(n1053), .ZN(n1204) );
XNOR2_X1 U888 ( .A(G131), .B(n1239), .ZN(G33) );
NAND2_X1 U889 ( .A1(KEYINPUT38), .A2(n1203), .ZN(n1239) );
AND3_X1 U890 ( .A1(n1236), .A2(n1197), .A3(n1053), .ZN(n1203) );
NOR3_X1 U891 ( .A1(n1058), .A2(n1234), .A3(n1036), .ZN(n1236) );
NAND2_X1 U892 ( .A1(n1240), .A2(n1092), .ZN(n1036) );
XOR2_X1 U893 ( .A(KEYINPUT11), .B(n1076), .Z(n1240) );
INV_X1 U894 ( .A(n1227), .ZN(n1058) );
XNOR2_X1 U895 ( .A(G128), .B(n1206), .ZN(G30) );
NAND3_X1 U896 ( .A1(n1228), .A2(n1057), .A3(n1241), .ZN(n1206) );
NOR4_X1 U897 ( .A1(n1242), .A2(n1073), .A3(n1243), .A4(n1234), .ZN(n1228) );
XNOR2_X1 U898 ( .A(n1244), .B(n1245), .ZN(G3) );
NAND2_X1 U899 ( .A1(KEYINPUT5), .A2(n1246), .ZN(n1244) );
NAND4_X1 U900 ( .A1(n1063), .A2(n1053), .A3(n1247), .A4(n1248), .ZN(n1246) );
OR2_X1 U901 ( .A1(n1196), .A2(KEYINPUT8), .ZN(n1248) );
INV_X1 U902 ( .A(n1182), .ZN(n1196) );
NAND2_X1 U903 ( .A1(KEYINPUT8), .A2(n1249), .ZN(n1247) );
XNOR2_X1 U904 ( .A(G125), .B(n1207), .ZN(G27) );
NAND4_X1 U905 ( .A1(n1197), .A2(n1054), .A3(n1250), .A4(n1071), .ZN(n1207) );
NOR2_X1 U906 ( .A1(n1234), .A2(n1073), .ZN(n1250) );
INV_X1 U907 ( .A(n1231), .ZN(n1073) );
AND2_X1 U908 ( .A1(n1251), .A2(n1044), .ZN(n1234) );
NAND3_X1 U909 ( .A1(G902), .A2(n1252), .A3(n1101), .ZN(n1251) );
NOR2_X1 U910 ( .A1(n1060), .A2(G900), .ZN(n1101) );
XOR2_X1 U911 ( .A(G122), .B(n1195), .Z(G24) );
NOR4_X1 U912 ( .A1(n1253), .A2(n1041), .A3(n1233), .A4(n1235), .ZN(n1195) );
INV_X1 U913 ( .A(n1064), .ZN(n1041) );
NOR2_X1 U914 ( .A1(n1082), .A2(n1237), .ZN(n1064) );
XOR2_X1 U915 ( .A(G119), .B(n1194), .Z(G21) );
NOR4_X1 U916 ( .A1(n1253), .A2(n1052), .A3(n1242), .A4(n1243), .ZN(n1194) );
XNOR2_X1 U917 ( .A(n1254), .B(n1192), .ZN(G18) );
NAND3_X1 U918 ( .A1(n1053), .A2(n1057), .A3(n1193), .ZN(n1192) );
INV_X1 U919 ( .A(n1253), .ZN(n1193) );
NAND3_X1 U920 ( .A1(n1231), .A2(n1255), .A3(n1071), .ZN(n1253) );
NOR2_X1 U921 ( .A1(n1084), .A2(n1235), .ZN(n1057) );
NAND2_X1 U922 ( .A1(KEYINPUT60), .A2(n1256), .ZN(n1254) );
INV_X1 U923 ( .A(G116), .ZN(n1256) );
XNOR2_X1 U924 ( .A(n1257), .B(n1258), .ZN(G15) );
NOR3_X1 U925 ( .A1(n1188), .A2(KEYINPUT9), .A3(n1190), .ZN(n1258) );
INV_X1 U926 ( .A(n1053), .ZN(n1190) );
NOR2_X1 U927 ( .A1(n1242), .A2(n1082), .ZN(n1053) );
NAND4_X1 U928 ( .A1(n1197), .A2(n1071), .A3(n1259), .A4(n1255), .ZN(n1188) );
INV_X1 U929 ( .A(n1042), .ZN(n1071) );
NAND2_X1 U930 ( .A1(n1068), .A2(n1260), .ZN(n1042) );
INV_X1 U931 ( .A(n1043), .ZN(n1197) );
NAND2_X1 U932 ( .A1(n1235), .A2(n1084), .ZN(n1043) );
XNOR2_X1 U933 ( .A(G110), .B(n1261), .ZN(G12) );
NAND4_X1 U934 ( .A1(n1063), .A2(n1054), .A3(n1262), .A4(n1263), .ZN(n1261) );
NAND2_X1 U935 ( .A1(KEYINPUT48), .A2(n1182), .ZN(n1263) );
NAND2_X1 U936 ( .A1(n1264), .A2(n1259), .ZN(n1182) );
INV_X1 U937 ( .A(n1265), .ZN(n1259) );
NAND2_X1 U938 ( .A1(n1249), .A2(n1266), .ZN(n1262) );
INV_X1 U939 ( .A(KEYINPUT48), .ZN(n1266) );
NAND2_X1 U940 ( .A1(n1264), .A2(n1265), .ZN(n1249) );
XOR2_X1 U941 ( .A(n1231), .B(KEYINPUT37), .Z(n1265) );
NOR2_X1 U942 ( .A1(n1076), .A2(n1075), .ZN(n1231) );
INV_X1 U943 ( .A(n1092), .ZN(n1075) );
NAND2_X1 U944 ( .A1(G214), .A2(n1267), .ZN(n1092) );
XNOR2_X1 U945 ( .A(n1091), .B(KEYINPUT0), .ZN(n1076) );
XNOR2_X1 U946 ( .A(n1268), .B(n1174), .ZN(n1091) );
NAND2_X1 U947 ( .A1(G210), .A2(n1267), .ZN(n1174) );
NAND2_X1 U948 ( .A1(n1269), .A2(n1210), .ZN(n1267) );
INV_X1 U949 ( .A(G237), .ZN(n1269) );
NAND2_X1 U950 ( .A1(n1270), .A2(n1271), .ZN(n1268) );
XNOR2_X1 U951 ( .A(n1272), .B(n1215), .ZN(n1270) );
INV_X1 U952 ( .A(n1219), .ZN(n1215) );
XNOR2_X1 U953 ( .A(n1273), .B(n1120), .ZN(n1219) );
XOR2_X1 U954 ( .A(G122), .B(n1274), .Z(n1120) );
NOR2_X1 U955 ( .A1(G110), .A2(KEYINPUT29), .ZN(n1274) );
NAND2_X1 U956 ( .A1(n1122), .A2(n1123), .ZN(n1273) );
NAND2_X1 U957 ( .A1(n1275), .A2(n1276), .ZN(n1123) );
XNOR2_X1 U958 ( .A(G101), .B(n1277), .ZN(n1275) );
NAND2_X1 U959 ( .A1(n1278), .A2(n1279), .ZN(n1122) );
XNOR2_X1 U960 ( .A(n1245), .B(n1277), .ZN(n1279) );
NOR2_X1 U961 ( .A1(KEYINPUT17), .A2(n1280), .ZN(n1277) );
INV_X1 U962 ( .A(G101), .ZN(n1245) );
INV_X1 U963 ( .A(n1276), .ZN(n1278) );
NAND2_X1 U964 ( .A1(n1281), .A2(n1282), .ZN(n1276) );
NAND2_X1 U965 ( .A1(n1283), .A2(G113), .ZN(n1282) );
XOR2_X1 U966 ( .A(KEYINPUT18), .B(n1284), .Z(n1281) );
NOR2_X1 U967 ( .A1(G113), .A2(n1283), .ZN(n1284) );
XNOR2_X1 U968 ( .A(G119), .B(n1285), .ZN(n1283) );
NOR2_X1 U969 ( .A1(G116), .A2(KEYINPUT19), .ZN(n1285) );
XNOR2_X1 U970 ( .A(n1286), .B(n1223), .ZN(n1272) );
NAND2_X1 U971 ( .A1(G224), .A2(n1060), .ZN(n1223) );
NAND2_X1 U972 ( .A1(KEYINPUT22), .A2(n1222), .ZN(n1286) );
XNOR2_X1 U973 ( .A(n1287), .B(G125), .ZN(n1222) );
AND2_X1 U974 ( .A1(n1241), .A2(n1255), .ZN(n1264) );
NAND2_X1 U975 ( .A1(n1044), .A2(n1288), .ZN(n1255) );
NAND4_X1 U976 ( .A1(G953), .A2(G902), .A3(n1252), .A4(n1289), .ZN(n1288) );
INV_X1 U977 ( .A(G898), .ZN(n1289) );
NAND3_X1 U978 ( .A1(n1252), .A2(n1060), .A3(G952), .ZN(n1044) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1252) );
XNOR2_X1 U980 ( .A(n1227), .B(KEYINPUT24), .ZN(n1241) );
NOR2_X1 U981 ( .A1(n1068), .A2(n1070), .ZN(n1227) );
INV_X1 U982 ( .A(n1260), .ZN(n1070) );
NAND2_X1 U983 ( .A1(G221), .A2(n1290), .ZN(n1260) );
XOR2_X1 U984 ( .A(n1291), .B(G469), .Z(n1068) );
NAND2_X1 U985 ( .A1(n1271), .A2(n1292), .ZN(n1291) );
XOR2_X1 U986 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U987 ( .A(n1295), .B(n1296), .ZN(n1294) );
NAND2_X1 U988 ( .A1(KEYINPUT6), .A2(G110), .ZN(n1296) );
NAND2_X1 U989 ( .A1(n1297), .A2(KEYINPUT58), .ZN(n1295) );
XOR2_X1 U990 ( .A(n1164), .B(n1298), .Z(n1297) );
NOR2_X1 U991 ( .A1(KEYINPUT4), .A2(n1165), .ZN(n1298) );
XOR2_X1 U992 ( .A(G101), .B(n1299), .Z(n1165) );
NOR2_X1 U993 ( .A1(KEYINPUT52), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U994 ( .A(KEYINPUT47), .B(n1280), .ZN(n1300) );
XNOR2_X1 U995 ( .A(G104), .B(G107), .ZN(n1280) );
XNOR2_X1 U996 ( .A(n1107), .B(n1152), .ZN(n1164) );
NAND4_X1 U997 ( .A1(n1301), .A2(n1302), .A3(n1303), .A4(n1304), .ZN(n1107) );
NAND3_X1 U998 ( .A1(KEYINPUT31), .A2(G128), .A3(n1230), .ZN(n1304) );
NAND3_X1 U999 ( .A1(n1305), .A2(n1306), .A3(G143), .ZN(n1303) );
OR2_X1 U1000 ( .A1(KEYINPUT31), .A2(G146), .ZN(n1305) );
OR2_X1 U1001 ( .A1(n1307), .A2(KEYINPUT31), .ZN(n1301) );
XNOR2_X1 U1002 ( .A(G140), .B(n1166), .ZN(n1293) );
AND2_X1 U1003 ( .A1(G227), .A2(n1060), .ZN(n1166) );
NOR2_X1 U1004 ( .A1(n1243), .A2(n1237), .ZN(n1054) );
INV_X1 U1005 ( .A(n1242), .ZN(n1237) );
XNOR2_X1 U1006 ( .A(n1093), .B(n1308), .ZN(n1242) );
NOR2_X1 U1007 ( .A1(G472), .A2(KEYINPUT35), .ZN(n1308) );
NAND2_X1 U1008 ( .A1(n1309), .A2(n1271), .ZN(n1093) );
XOR2_X1 U1009 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1010 ( .A(KEYINPUT15), .B(n1152), .ZN(n1311) );
INV_X1 U1011 ( .A(n1155), .ZN(n1152) );
XNOR2_X1 U1012 ( .A(n1312), .B(G131), .ZN(n1155) );
NAND2_X1 U1013 ( .A1(KEYINPUT39), .A2(n1108), .ZN(n1312) );
XNOR2_X1 U1014 ( .A(G137), .B(n1313), .ZN(n1108) );
XOR2_X1 U1015 ( .A(n1154), .B(n1157), .Z(n1310) );
XNOR2_X1 U1016 ( .A(n1314), .B(G101), .ZN(n1157) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1315), .ZN(n1314) );
XNOR2_X1 U1018 ( .A(n1316), .B(n1287), .ZN(n1154) );
NAND3_X1 U1019 ( .A1(n1307), .A2(n1302), .A3(n1317), .ZN(n1287) );
NAND3_X1 U1020 ( .A1(G143), .A2(n1306), .A3(G146), .ZN(n1317) );
INV_X1 U1021 ( .A(G128), .ZN(n1306) );
NAND3_X1 U1022 ( .A1(G146), .A2(n1230), .A3(G128), .ZN(n1302) );
NAND2_X1 U1023 ( .A1(n1318), .A2(n1226), .ZN(n1307) );
INV_X1 U1024 ( .A(G146), .ZN(n1226) );
XNOR2_X1 U1025 ( .A(G128), .B(G143), .ZN(n1318) );
NAND3_X1 U1026 ( .A1(n1319), .A2(n1320), .A3(n1321), .ZN(n1316) );
NAND2_X1 U1027 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
INV_X1 U1028 ( .A(KEYINPUT50), .ZN(n1323) );
NAND3_X1 U1029 ( .A1(KEYINPUT50), .A2(n1324), .A3(n1257), .ZN(n1320) );
OR2_X1 U1030 ( .A1(n1257), .A2(n1324), .ZN(n1319) );
NOR2_X1 U1031 ( .A1(KEYINPUT44), .A2(n1322), .ZN(n1324) );
XNOR2_X1 U1032 ( .A(G116), .B(G119), .ZN(n1322) );
INV_X1 U1033 ( .A(n1082), .ZN(n1243) );
XNOR2_X1 U1034 ( .A(n1325), .B(n1131), .ZN(n1082) );
AND2_X1 U1035 ( .A1(G217), .A2(n1290), .ZN(n1131) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1210), .ZN(n1290) );
INV_X1 U1037 ( .A(G902), .ZN(n1210) );
OR2_X1 U1038 ( .A1(n1326), .A2(n1129), .ZN(n1325) );
XOR2_X1 U1039 ( .A(n1327), .B(n1328), .Z(n1129) );
XOR2_X1 U1040 ( .A(G119), .B(n1329), .Z(n1328) );
XNOR2_X1 U1041 ( .A(n1330), .B(G128), .ZN(n1329) );
INV_X1 U1042 ( .A(G137), .ZN(n1330) );
XOR2_X1 U1043 ( .A(n1331), .B(n1332), .Z(n1327) );
XOR2_X1 U1044 ( .A(n1333), .B(n1334), .Z(n1332) );
NAND2_X1 U1045 ( .A1(KEYINPUT1), .A2(G110), .ZN(n1334) );
NAND2_X1 U1046 ( .A1(G221), .A2(n1335), .ZN(n1333) );
INV_X1 U1047 ( .A(n1052), .ZN(n1063) );
NAND2_X1 U1048 ( .A1(n1235), .A2(n1233), .ZN(n1052) );
INV_X1 U1049 ( .A(n1084), .ZN(n1233) );
XNOR2_X1 U1050 ( .A(n1336), .B(G475), .ZN(n1084) );
NAND2_X1 U1051 ( .A1(n1271), .A2(n1145), .ZN(n1336) );
XOR2_X1 U1052 ( .A(n1337), .B(n1338), .Z(n1145) );
XOR2_X1 U1053 ( .A(n1339), .B(n1340), .Z(n1338) );
XNOR2_X1 U1054 ( .A(G122), .B(n1257), .ZN(n1340) );
INV_X1 U1055 ( .A(G113), .ZN(n1257) );
XOR2_X1 U1056 ( .A(KEYINPUT27), .B(G131), .Z(n1339) );
XOR2_X1 U1057 ( .A(n1341), .B(n1342), .Z(n1337) );
NOR2_X1 U1058 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NOR2_X1 U1059 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XNOR2_X1 U1060 ( .A(n1347), .B(n1230), .ZN(n1346) );
XNOR2_X1 U1061 ( .A(KEYINPUT33), .B(KEYINPUT25), .ZN(n1347) );
AND2_X1 U1062 ( .A1(n1230), .A2(n1345), .ZN(n1343) );
NAND2_X1 U1063 ( .A1(G214), .A2(n1315), .ZN(n1345) );
NOR2_X1 U1064 ( .A1(G953), .A2(G237), .ZN(n1315) );
XOR2_X1 U1065 ( .A(n1331), .B(G104), .Z(n1341) );
XNOR2_X1 U1066 ( .A(G146), .B(n1109), .ZN(n1331) );
XNOR2_X1 U1067 ( .A(n1348), .B(G140), .ZN(n1109) );
INV_X1 U1068 ( .A(G125), .ZN(n1348) );
INV_X1 U1069 ( .A(n1326), .ZN(n1271) );
AND3_X1 U1070 ( .A1(n1349), .A2(n1350), .A3(n1088), .ZN(n1235) );
NAND2_X1 U1071 ( .A1(n1351), .A2(n1136), .ZN(n1088) );
INV_X1 U1072 ( .A(G478), .ZN(n1136) );
OR2_X1 U1073 ( .A1(G478), .A2(KEYINPUT16), .ZN(n1350) );
NAND3_X1 U1074 ( .A1(G478), .A2(n1089), .A3(KEYINPUT16), .ZN(n1349) );
INV_X1 U1075 ( .A(n1351), .ZN(n1089) );
NOR2_X1 U1076 ( .A1(n1326), .A2(n1133), .ZN(n1351) );
XNOR2_X1 U1077 ( .A(n1352), .B(n1353), .ZN(n1133) );
NOR2_X1 U1078 ( .A1(KEYINPUT51), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1079 ( .A(n1355), .B(n1356), .Z(n1354) );
XOR2_X1 U1080 ( .A(n1313), .B(n1357), .Z(n1356) );
XNOR2_X1 U1081 ( .A(G107), .B(n1358), .ZN(n1357) );
NOR2_X1 U1082 ( .A1(G128), .A2(KEYINPUT42), .ZN(n1358) );
XNOR2_X1 U1083 ( .A(G134), .B(KEYINPUT59), .ZN(n1313) );
XNOR2_X1 U1084 ( .A(G116), .B(n1359), .ZN(n1355) );
XNOR2_X1 U1085 ( .A(n1230), .B(G122), .ZN(n1359) );
INV_X1 U1086 ( .A(G143), .ZN(n1230) );
NAND2_X1 U1087 ( .A1(G217), .A2(n1335), .ZN(n1352) );
AND2_X1 U1088 ( .A1(G234), .A2(n1060), .ZN(n1335) );
INV_X1 U1089 ( .A(G953), .ZN(n1060) );
XOR2_X1 U1090 ( .A(G902), .B(KEYINPUT56), .Z(n1326) );
endmodule


