//Key = 1101001001001101010100100010010010000111011100011010101010000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390;

XNOR2_X1 U754 ( .A(G107), .B(n1050), .ZN(G9) );
NAND4_X1 U755 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
XNOR2_X1 U756 ( .A(KEYINPUT32), .B(n1055), .ZN(n1054) );
NOR2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(G75) );
NOR3_X1 U758 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
XOR2_X1 U759 ( .A(n1061), .B(KEYINPUT44), .Z(n1059) );
NAND3_X1 U760 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1058) );
NAND2_X1 U761 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U762 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND4_X1 U763 ( .A1(n1069), .A2(n1070), .A3(n1053), .A4(n1071), .ZN(n1068) );
NAND2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U766 ( .A1(n1076), .A2(n1077), .A3(n1075), .ZN(n1067) );
NAND2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1080), .ZN(n1079) );
NAND2_X1 U769 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U770 ( .A1(n1083), .A2(n1053), .ZN(n1082) );
XNOR2_X1 U771 ( .A(n1084), .B(n1085), .ZN(n1083) );
NAND2_X1 U772 ( .A1(n1069), .A2(n1086), .ZN(n1081) );
NAND2_X1 U773 ( .A1(n1069), .A2(n1087), .ZN(n1078) );
INV_X1 U774 ( .A(n1088), .ZN(n1065) );
NOR3_X1 U775 ( .A1(n1089), .A2(G953), .A3(G952), .ZN(n1056) );
INV_X1 U776 ( .A(n1062), .ZN(n1089) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1062) );
NOR4_X1 U778 ( .A1(n1074), .A2(n1084), .A3(n1092), .A4(n1093), .ZN(n1091) );
XOR2_X1 U779 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U780 ( .A1(KEYINPUT0), .A2(n1096), .ZN(n1094) );
NOR2_X1 U781 ( .A1(G478), .A2(n1097), .ZN(n1092) );
NOR4_X1 U782 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1090) );
XNOR2_X1 U783 ( .A(KEYINPUT11), .B(n1102), .ZN(n1101) );
XNOR2_X1 U784 ( .A(n1103), .B(n1104), .ZN(n1100) );
XOR2_X1 U785 ( .A(n1105), .B(n1106), .Z(n1098) );
XOR2_X1 U786 ( .A(KEYINPUT60), .B(KEYINPUT46), .Z(n1106) );
XOR2_X1 U787 ( .A(n1107), .B(n1108), .Z(n1105) );
NOR2_X1 U788 ( .A1(G469), .A2(KEYINPUT4), .ZN(n1108) );
XOR2_X1 U789 ( .A(n1109), .B(n1110), .Z(G72) );
XOR2_X1 U790 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U791 ( .A1(n1113), .A2(n1063), .ZN(n1112) );
AND2_X1 U792 ( .A1(G227), .A2(G900), .ZN(n1113) );
NAND2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U794 ( .A1(G953), .A2(n1116), .ZN(n1115) );
XOR2_X1 U795 ( .A(n1117), .B(n1118), .Z(n1114) );
XNOR2_X1 U796 ( .A(G131), .B(n1119), .ZN(n1118) );
NAND2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U798 ( .A(KEYINPUT47), .B(n1122), .Z(n1120) );
NOR2_X1 U799 ( .A1(G134), .A2(n1123), .ZN(n1122) );
XOR2_X1 U800 ( .A(n1124), .B(n1125), .Z(n1117) );
NAND2_X1 U801 ( .A1(n1063), .A2(n1061), .ZN(n1109) );
NAND2_X1 U802 ( .A1(n1126), .A2(n1127), .ZN(G69) );
NAND2_X1 U803 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U804 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U805 ( .A1(G953), .A2(n1132), .ZN(n1131) );
INV_X1 U806 ( .A(n1133), .ZN(n1130) );
NAND2_X1 U807 ( .A1(n1134), .A2(n1135), .ZN(n1126) );
INV_X1 U808 ( .A(n1128), .ZN(n1135) );
NOR2_X1 U809 ( .A1(KEYINPUT16), .A2(n1136), .ZN(n1128) );
NOR3_X1 U810 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
NOR3_X1 U811 ( .A1(n1140), .A2(KEYINPUT33), .A3(n1141), .ZN(n1139) );
NOR2_X1 U812 ( .A1(n1142), .A2(n1143), .ZN(n1138) );
NOR2_X1 U813 ( .A1(n1144), .A2(KEYINPUT33), .ZN(n1143) );
NOR2_X1 U814 ( .A1(KEYINPUT24), .A2(n1145), .ZN(n1144) );
INV_X1 U815 ( .A(n1140), .ZN(n1142) );
NAND2_X1 U816 ( .A1(n1063), .A2(n1060), .ZN(n1140) );
AND2_X1 U817 ( .A1(n1145), .A2(KEYINPUT24), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1133), .ZN(n1145) );
XNOR2_X1 U819 ( .A(n1146), .B(n1147), .ZN(n1141) );
NAND2_X1 U820 ( .A1(G953), .A2(n1148), .ZN(n1134) );
NAND2_X1 U821 ( .A1(G898), .A2(G224), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1149), .A2(n1150), .ZN(G66) );
XOR2_X1 U823 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR3_X1 U824 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
XNOR2_X1 U825 ( .A(G902), .B(KEYINPUT20), .ZN(n1155) );
NAND2_X1 U826 ( .A1(KEYINPUT15), .A2(n1156), .ZN(n1151) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1157), .ZN(G63) );
XOR2_X1 U828 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U829 ( .A1(n1160), .A2(G478), .ZN(n1158) );
NOR2_X1 U830 ( .A1(n1149), .A2(n1161), .ZN(G60) );
XOR2_X1 U831 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND3_X1 U832 ( .A1(KEYINPUT13), .A2(n1160), .A3(n1164), .ZN(n1163) );
XNOR2_X1 U833 ( .A(G475), .B(KEYINPUT22), .ZN(n1164) );
XOR2_X1 U834 ( .A(G104), .B(n1165), .Z(G6) );
NOR4_X1 U835 ( .A1(KEYINPUT55), .A2(n1099), .A3(n1166), .A4(n1167), .ZN(n1165) );
INV_X1 U836 ( .A(n1053), .ZN(n1099) );
NOR2_X1 U837 ( .A1(n1149), .A2(n1168), .ZN(G57) );
XOR2_X1 U838 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U839 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U840 ( .A(n1173), .B(n1174), .ZN(n1172) );
NAND2_X1 U841 ( .A1(KEYINPUT29), .A2(n1175), .ZN(n1174) );
NAND2_X1 U842 ( .A1(KEYINPUT52), .A2(n1176), .ZN(n1173) );
XOR2_X1 U843 ( .A(n1177), .B(n1178), .Z(n1169) );
XNOR2_X1 U844 ( .A(n1179), .B(KEYINPUT57), .ZN(n1178) );
NAND2_X1 U845 ( .A1(n1160), .A2(G472), .ZN(n1177) );
NOR2_X1 U846 ( .A1(n1149), .A2(n1180), .ZN(G54) );
XOR2_X1 U847 ( .A(n1181), .B(n1182), .Z(n1180) );
XNOR2_X1 U848 ( .A(n1175), .B(n1183), .ZN(n1182) );
XOR2_X1 U849 ( .A(n1184), .B(n1185), .Z(n1181) );
XOR2_X1 U850 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U851 ( .A1(KEYINPUT8), .A2(n1188), .ZN(n1187) );
NOR2_X1 U852 ( .A1(KEYINPUT40), .A2(n1189), .ZN(n1186) );
NAND2_X1 U853 ( .A1(n1160), .A2(G469), .ZN(n1184) );
NOR2_X1 U854 ( .A1(n1149), .A2(n1190), .ZN(G51) );
XOR2_X1 U855 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U856 ( .A(n1193), .B(n1194), .Z(n1192) );
XNOR2_X1 U857 ( .A(n1195), .B(n1196), .ZN(n1193) );
NAND2_X1 U858 ( .A1(n1160), .A2(n1095), .ZN(n1195) );
NOR2_X1 U859 ( .A1(n1197), .A2(n1154), .ZN(n1160) );
NOR2_X1 U860 ( .A1(n1060), .A2(n1061), .ZN(n1154) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1061) );
NOR4_X1 U862 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
INV_X1 U863 ( .A(n1204), .ZN(n1203) );
NOR4_X1 U864 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1198) );
NOR2_X1 U865 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND4_X1 U866 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1060) );
AND3_X1 U867 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
NAND2_X1 U868 ( .A1(n1218), .A2(n1087), .ZN(n1213) );
NAND2_X1 U869 ( .A1(n1219), .A2(n1220), .ZN(n1087) );
NAND2_X1 U870 ( .A1(n1053), .A2(n1221), .ZN(n1220) );
NAND2_X1 U871 ( .A1(n1167), .A2(n1209), .ZN(n1221) );
INV_X1 U872 ( .A(n1052), .ZN(n1209) );
NAND2_X1 U873 ( .A1(n1222), .A2(n1070), .ZN(n1219) );
NAND2_X1 U874 ( .A1(n1223), .A2(n1224), .ZN(n1211) );
XOR2_X1 U875 ( .A(n1225), .B(KEYINPUT3), .Z(n1223) );
XOR2_X1 U876 ( .A(n1226), .B(n1227), .Z(n1191) );
XNOR2_X1 U877 ( .A(n1228), .B(n1229), .ZN(n1227) );
XNOR2_X1 U878 ( .A(KEYINPUT48), .B(KEYINPUT34), .ZN(n1226) );
NOR2_X1 U879 ( .A1(n1063), .A2(G952), .ZN(n1149) );
XOR2_X1 U880 ( .A(G146), .B(n1206), .Z(G48) );
AND2_X1 U881 ( .A1(n1230), .A2(n1231), .ZN(n1206) );
NAND2_X1 U882 ( .A1(n1232), .A2(n1233), .ZN(G45) );
NAND2_X1 U883 ( .A1(G143), .A2(n1234), .ZN(n1233) );
XOR2_X1 U884 ( .A(n1235), .B(KEYINPUT18), .Z(n1232) );
NAND2_X1 U885 ( .A1(n1207), .A2(n1236), .ZN(n1235) );
INV_X1 U886 ( .A(n1234), .ZN(n1207) );
NAND3_X1 U887 ( .A1(n1222), .A2(n1051), .A3(n1237), .ZN(n1234) );
NOR3_X1 U888 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1237) );
XOR2_X1 U889 ( .A(G140), .B(n1205), .Z(G42) );
AND3_X1 U890 ( .A1(n1231), .A2(n1086), .A3(n1241), .ZN(n1205) );
XNOR2_X1 U891 ( .A(G137), .B(n1204), .ZN(G39) );
NAND2_X1 U892 ( .A1(n1241), .A2(n1242), .ZN(n1204) );
XOR2_X1 U893 ( .A(G134), .B(n1243), .Z(G36) );
NOR2_X1 U894 ( .A1(n1244), .A2(n1210), .ZN(n1243) );
XNOR2_X1 U895 ( .A(n1052), .B(KEYINPUT10), .ZN(n1244) );
NAND2_X1 U896 ( .A1(n1245), .A2(n1246), .ZN(G33) );
NAND2_X1 U897 ( .A1(n1202), .A2(n1247), .ZN(n1246) );
XOR2_X1 U898 ( .A(KEYINPUT6), .B(n1248), .Z(n1245) );
NOR2_X1 U899 ( .A1(n1202), .A2(n1247), .ZN(n1248) );
INV_X1 U900 ( .A(G131), .ZN(n1247) );
NOR2_X1 U901 ( .A1(n1210), .A2(n1167), .ZN(n1202) );
NAND2_X1 U902 ( .A1(n1241), .A2(n1222), .ZN(n1210) );
AND4_X1 U903 ( .A1(n1249), .A2(n1077), .A3(n1250), .A4(n1251), .ZN(n1241) );
NOR2_X1 U904 ( .A1(n1252), .A2(n1085), .ZN(n1251) );
XNOR2_X1 U905 ( .A(n1253), .B(n1201), .ZN(G30) );
AND2_X1 U906 ( .A1(n1230), .A2(n1052), .ZN(n1201) );
AND4_X1 U907 ( .A1(n1051), .A2(n1254), .A3(n1255), .A4(n1250), .ZN(n1230) );
XNOR2_X1 U908 ( .A(G101), .B(n1256), .ZN(G3) );
NAND3_X1 U909 ( .A1(n1218), .A2(n1070), .A3(n1257), .ZN(n1256) );
XNOR2_X1 U910 ( .A(n1222), .B(KEYINPUT38), .ZN(n1257) );
NAND2_X1 U911 ( .A1(n1258), .A2(n1259), .ZN(G27) );
NAND2_X1 U912 ( .A1(n1260), .A2(n1228), .ZN(n1259) );
NAND2_X1 U913 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NAND2_X1 U914 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
OR2_X1 U915 ( .A1(n1264), .A2(n1265), .ZN(n1261) );
INV_X1 U916 ( .A(KEYINPUT54), .ZN(n1264) );
NAND2_X1 U917 ( .A1(G125), .A2(n1265), .ZN(n1258) );
NOR2_X1 U918 ( .A1(n1200), .A2(KEYINPUT23), .ZN(n1265) );
INV_X1 U919 ( .A(n1263), .ZN(n1200) );
NAND3_X1 U920 ( .A1(n1231), .A2(n1069), .A3(n1266), .ZN(n1263) );
NOR3_X1 U921 ( .A1(n1267), .A2(n1240), .A3(n1072), .ZN(n1266) );
INV_X1 U922 ( .A(n1250), .ZN(n1240) );
NAND2_X1 U923 ( .A1(n1088), .A2(n1268), .ZN(n1250) );
NAND4_X1 U924 ( .A1(G902), .A2(G953), .A3(n1269), .A4(n1116), .ZN(n1268) );
INV_X1 U925 ( .A(G900), .ZN(n1116) );
NAND2_X1 U926 ( .A1(n1270), .A2(n1271), .ZN(G24) );
NAND2_X1 U927 ( .A1(G122), .A2(n1212), .ZN(n1271) );
XOR2_X1 U928 ( .A(n1272), .B(KEYINPUT7), .Z(n1270) );
OR2_X1 U929 ( .A1(n1212), .A2(G122), .ZN(n1272) );
NAND4_X1 U930 ( .A1(n1273), .A2(n1053), .A3(n1274), .A4(n1275), .ZN(n1212) );
NOR2_X1 U931 ( .A1(n1255), .A2(n1254), .ZN(n1053) );
NAND2_X1 U932 ( .A1(n1276), .A2(n1277), .ZN(G21) );
NAND2_X1 U933 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U934 ( .A(KEYINPUT37), .B(n1280), .Z(n1276) );
NOR2_X1 U935 ( .A1(n1278), .A2(n1279), .ZN(n1280) );
XNOR2_X1 U936 ( .A(KEYINPUT12), .B(n1281), .ZN(n1279) );
INV_X1 U937 ( .A(n1215), .ZN(n1278) );
NAND2_X1 U938 ( .A1(n1242), .A2(n1273), .ZN(n1215) );
AND3_X1 U939 ( .A1(n1254), .A2(n1255), .A3(n1070), .ZN(n1242) );
XOR2_X1 U940 ( .A(G116), .B(n1282), .Z(G18) );
NOR2_X1 U941 ( .A1(n1072), .A2(n1225), .ZN(n1282) );
NAND4_X1 U942 ( .A1(n1222), .A2(n1069), .A3(n1052), .A4(n1055), .ZN(n1225) );
NOR2_X1 U943 ( .A1(n1274), .A2(n1239), .ZN(n1052) );
XNOR2_X1 U944 ( .A(G113), .B(n1217), .ZN(G15) );
NAND3_X1 U945 ( .A1(n1222), .A2(n1231), .A3(n1273), .ZN(n1217) );
AND3_X1 U946 ( .A1(n1224), .A2(n1055), .A3(n1069), .ZN(n1273) );
AND2_X1 U947 ( .A1(n1085), .A2(n1249), .ZN(n1069) );
INV_X1 U948 ( .A(n1167), .ZN(n1231) );
NAND2_X1 U949 ( .A1(n1239), .A2(n1283), .ZN(n1167) );
XNOR2_X1 U950 ( .A(KEYINPUT14), .B(n1238), .ZN(n1283) );
INV_X1 U951 ( .A(n1274), .ZN(n1238) );
INV_X1 U952 ( .A(n1275), .ZN(n1239) );
NOR2_X1 U953 ( .A1(n1254), .A2(n1284), .ZN(n1222) );
XNOR2_X1 U954 ( .A(G110), .B(n1216), .ZN(G12) );
NAND3_X1 U955 ( .A1(n1218), .A2(n1070), .A3(n1086), .ZN(n1216) );
INV_X1 U956 ( .A(n1267), .ZN(n1086) );
NAND2_X1 U957 ( .A1(n1284), .A2(n1254), .ZN(n1267) );
XOR2_X1 U958 ( .A(n1285), .B(n1153), .Z(n1254) );
NAND2_X1 U959 ( .A1(G217), .A2(n1286), .ZN(n1153) );
NAND2_X1 U960 ( .A1(n1156), .A2(n1197), .ZN(n1285) );
XOR2_X1 U961 ( .A(n1287), .B(n1288), .Z(n1156) );
XNOR2_X1 U962 ( .A(G137), .B(n1289), .ZN(n1288) );
NAND2_X1 U963 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U964 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U965 ( .A(n1294), .B(KEYINPUT25), .Z(n1290) );
OR2_X1 U966 ( .A1(n1293), .A2(n1292), .ZN(n1294) );
XOR2_X1 U967 ( .A(n1295), .B(n1296), .Z(n1292) );
NOR2_X1 U968 ( .A1(KEYINPUT49), .A2(n1281), .ZN(n1296) );
XNOR2_X1 U969 ( .A(G110), .B(G128), .ZN(n1295) );
XNOR2_X1 U970 ( .A(G146), .B(n1124), .ZN(n1293) );
NAND2_X1 U971 ( .A1(n1297), .A2(G221), .ZN(n1287) );
INV_X1 U972 ( .A(n1255), .ZN(n1284) );
XNOR2_X1 U973 ( .A(n1298), .B(G472), .ZN(n1255) );
NAND2_X1 U974 ( .A1(n1299), .A2(n1197), .ZN(n1298) );
XOR2_X1 U975 ( .A(n1171), .B(n1300), .Z(n1299) );
XNOR2_X1 U976 ( .A(KEYINPUT45), .B(n1301), .ZN(n1300) );
NOR2_X1 U977 ( .A1(KEYINPUT31), .A2(n1302), .ZN(n1301) );
XNOR2_X1 U978 ( .A(n1175), .B(n1303), .ZN(n1302) );
XNOR2_X1 U979 ( .A(n1179), .B(n1176), .ZN(n1303) );
NAND3_X1 U980 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1176) );
OR2_X1 U981 ( .A1(n1307), .A2(G113), .ZN(n1306) );
NAND2_X1 U982 ( .A1(n1308), .A2(n1309), .ZN(n1305) );
INV_X1 U983 ( .A(KEYINPUT39), .ZN(n1309) );
NAND2_X1 U984 ( .A1(n1310), .A2(n1307), .ZN(n1308) );
XNOR2_X1 U985 ( .A(KEYINPUT9), .B(G113), .ZN(n1310) );
NAND2_X1 U986 ( .A1(KEYINPUT39), .A2(n1311), .ZN(n1304) );
NAND2_X1 U987 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
OR2_X1 U988 ( .A1(G113), .A2(KEYINPUT9), .ZN(n1313) );
NAND3_X1 U989 ( .A1(G113), .A2(n1307), .A3(KEYINPUT9), .ZN(n1312) );
XOR2_X1 U990 ( .A(n1314), .B(KEYINPUT2), .Z(n1307) );
INV_X1 U991 ( .A(n1196), .ZN(n1179) );
XNOR2_X1 U992 ( .A(n1315), .B(n1316), .ZN(n1171) );
INV_X1 U993 ( .A(G101), .ZN(n1316) );
NAND2_X1 U994 ( .A1(n1317), .A2(G210), .ZN(n1315) );
NOR2_X1 U995 ( .A1(n1275), .A2(n1274), .ZN(n1070) );
XOR2_X1 U996 ( .A(n1318), .B(n1103), .Z(n1274) );
NAND2_X1 U997 ( .A1(n1319), .A2(n1197), .ZN(n1103) );
XOR2_X1 U998 ( .A(n1162), .B(KEYINPUT63), .Z(n1319) );
NAND2_X1 U999 ( .A1(n1320), .A2(n1321), .ZN(n1162) );
NAND2_X1 U1000 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1001 ( .A(KEYINPUT43), .B(n1324), .Z(n1320) );
NOR2_X1 U1002 ( .A1(n1322), .A2(n1323), .ZN(n1324) );
XOR2_X1 U1003 ( .A(G104), .B(n1325), .Z(n1323) );
XOR2_X1 U1004 ( .A(G122), .B(G113), .Z(n1325) );
XOR2_X1 U1005 ( .A(n1326), .B(n1327), .Z(n1322) );
NOR2_X1 U1006 ( .A1(KEYINPUT28), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1007 ( .A(n1329), .B(n1330), .Z(n1328) );
XNOR2_X1 U1008 ( .A(n1236), .B(G131), .ZN(n1330) );
NAND2_X1 U1009 ( .A1(n1317), .A2(G214), .ZN(n1329) );
NOR2_X1 U1010 ( .A1(G953), .A2(G237), .ZN(n1317) );
NAND2_X1 U1011 ( .A1(n1331), .A2(n1332), .ZN(n1326) );
NAND2_X1 U1012 ( .A1(n1124), .A2(n1333), .ZN(n1332) );
NAND2_X1 U1013 ( .A1(G146), .A2(n1334), .ZN(n1333) );
OR2_X1 U1014 ( .A1(KEYINPUT21), .A2(KEYINPUT41), .ZN(n1334) );
NAND3_X1 U1015 ( .A1(n1335), .A2(n1336), .A3(KEYINPUT41), .ZN(n1331) );
OR2_X1 U1016 ( .A1(G146), .A2(KEYINPUT21), .ZN(n1336) );
NAND2_X1 U1017 ( .A1(G146), .A2(n1337), .ZN(n1335) );
OR2_X1 U1018 ( .A1(n1124), .A2(KEYINPUT21), .ZN(n1337) );
XOR2_X1 U1019 ( .A(G140), .B(n1228), .Z(n1124) );
NAND2_X1 U1020 ( .A1(KEYINPUT19), .A2(n1104), .ZN(n1318) );
XOR2_X1 U1021 ( .A(G475), .B(KEYINPUT35), .Z(n1104) );
NAND2_X1 U1022 ( .A1(n1338), .A2(n1102), .ZN(n1275) );
NAND2_X1 U1023 ( .A1(G478), .A2(n1097), .ZN(n1102) );
OR2_X1 U1024 ( .A1(n1097), .A2(G478), .ZN(n1338) );
NAND2_X1 U1025 ( .A1(n1159), .A2(n1197), .ZN(n1097) );
XOR2_X1 U1026 ( .A(n1339), .B(n1340), .Z(n1159) );
XOR2_X1 U1027 ( .A(G116), .B(n1341), .Z(n1340) );
XOR2_X1 U1028 ( .A(G134), .B(G122), .Z(n1341) );
XOR2_X1 U1029 ( .A(n1342), .B(n1343), .Z(n1339) );
XOR2_X1 U1030 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1031 ( .A1(G217), .A2(n1297), .ZN(n1345) );
AND2_X1 U1032 ( .A1(G234), .A2(n1063), .ZN(n1297) );
NAND2_X1 U1033 ( .A1(KEYINPUT50), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1034 ( .A(KEYINPUT62), .B(G107), .Z(n1346) );
NAND2_X1 U1035 ( .A1(n1347), .A2(n1348), .ZN(n1342) );
XOR2_X1 U1036 ( .A(n1349), .B(KEYINPUT61), .Z(n1347) );
NAND2_X1 U1037 ( .A1(G128), .A2(n1236), .ZN(n1349) );
INV_X1 U1038 ( .A(n1166), .ZN(n1218) );
NAND2_X1 U1039 ( .A1(n1051), .A2(n1055), .ZN(n1166) );
NAND2_X1 U1040 ( .A1(n1088), .A2(n1350), .ZN(n1055) );
NAND3_X1 U1041 ( .A1(n1133), .A2(n1269), .A3(G902), .ZN(n1350) );
NOR2_X1 U1042 ( .A1(n1063), .A2(G898), .ZN(n1133) );
NAND3_X1 U1043 ( .A1(n1269), .A2(n1063), .A3(G952), .ZN(n1088) );
NAND2_X1 U1044 ( .A1(G237), .A2(G234), .ZN(n1269) );
NOR3_X1 U1045 ( .A1(n1085), .A2(n1084), .A3(n1072), .ZN(n1051) );
INV_X1 U1046 ( .A(n1224), .ZN(n1072) );
NOR2_X1 U1047 ( .A1(n1075), .A2(n1074), .ZN(n1224) );
INV_X1 U1048 ( .A(n1077), .ZN(n1074) );
NAND2_X1 U1049 ( .A1(G214), .A2(n1351), .ZN(n1077) );
INV_X1 U1050 ( .A(n1252), .ZN(n1075) );
XNOR2_X1 U1051 ( .A(n1096), .B(n1095), .ZN(n1252) );
AND2_X1 U1052 ( .A1(G210), .A2(n1351), .ZN(n1095) );
NAND2_X1 U1053 ( .A1(n1352), .A2(n1197), .ZN(n1351) );
INV_X1 U1054 ( .A(G237), .ZN(n1352) );
NAND2_X1 U1055 ( .A1(n1353), .A2(n1197), .ZN(n1096) );
XNOR2_X1 U1056 ( .A(n1194), .B(n1354), .ZN(n1353) );
NOR3_X1 U1057 ( .A1(KEYINPUT36), .A2(n1355), .A3(n1356), .ZN(n1354) );
NOR2_X1 U1058 ( .A1(G125), .A2(n1357), .ZN(n1356) );
XOR2_X1 U1059 ( .A(KEYINPUT17), .B(n1358), .Z(n1357) );
NOR2_X1 U1060 ( .A1(n1358), .A2(n1228), .ZN(n1355) );
INV_X1 U1061 ( .A(G125), .ZN(n1228) );
XNOR2_X1 U1062 ( .A(n1196), .B(n1229), .ZN(n1358) );
NOR2_X1 U1063 ( .A1(n1132), .A2(G953), .ZN(n1229) );
INV_X1 U1064 ( .A(G224), .ZN(n1132) );
NAND3_X1 U1065 ( .A1(n1359), .A2(n1360), .A3(n1361), .ZN(n1196) );
OR2_X1 U1066 ( .A1(n1348), .A2(n1362), .ZN(n1361) );
NAND2_X1 U1067 ( .A1(G143), .A2(n1253), .ZN(n1348) );
NAND3_X1 U1068 ( .A1(G128), .A2(n1362), .A3(G143), .ZN(n1360) );
NAND2_X1 U1069 ( .A1(n1363), .A2(n1236), .ZN(n1359) );
XNOR2_X1 U1070 ( .A(n1253), .B(n1362), .ZN(n1363) );
XOR2_X1 U1071 ( .A(G146), .B(KEYINPUT26), .Z(n1362) );
XOR2_X1 U1072 ( .A(n1147), .B(n1364), .Z(n1194) );
XNOR2_X1 U1073 ( .A(n1365), .B(KEYINPUT56), .ZN(n1364) );
NAND2_X1 U1074 ( .A1(KEYINPUT1), .A2(n1146), .ZN(n1365) );
XOR2_X1 U1075 ( .A(n1366), .B(n1314), .Z(n1146) );
XNOR2_X1 U1076 ( .A(G116), .B(n1281), .ZN(n1314) );
INV_X1 U1077 ( .A(G119), .ZN(n1281) );
XOR2_X1 U1078 ( .A(n1367), .B(G113), .Z(n1366) );
NAND2_X1 U1079 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
OR2_X1 U1080 ( .A1(n1370), .A2(G101), .ZN(n1369) );
XOR2_X1 U1081 ( .A(n1371), .B(KEYINPUT5), .Z(n1368) );
NAND2_X1 U1082 ( .A1(G101), .A2(n1370), .ZN(n1371) );
XOR2_X1 U1083 ( .A(G110), .B(G122), .Z(n1147) );
INV_X1 U1084 ( .A(n1249), .ZN(n1084) );
NAND2_X1 U1085 ( .A1(G221), .A2(n1286), .ZN(n1249) );
NAND2_X1 U1086 ( .A1(G234), .A2(n1197), .ZN(n1286) );
NAND2_X1 U1087 ( .A1(n1372), .A2(n1373), .ZN(n1085) );
NAND2_X1 U1088 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
INV_X1 U1089 ( .A(G469), .ZN(n1375) );
XOR2_X1 U1090 ( .A(n1107), .B(KEYINPUT27), .Z(n1374) );
NAND2_X1 U1091 ( .A1(n1376), .A2(G469), .ZN(n1372) );
XNOR2_X1 U1092 ( .A(KEYINPUT53), .B(n1107), .ZN(n1376) );
NAND2_X1 U1093 ( .A1(n1377), .A2(n1197), .ZN(n1107) );
INV_X1 U1094 ( .A(G902), .ZN(n1197) );
XOR2_X1 U1095 ( .A(n1378), .B(n1379), .Z(n1377) );
XOR2_X1 U1096 ( .A(n1188), .B(n1183), .Z(n1379) );
XOR2_X1 U1097 ( .A(G140), .B(G110), .Z(n1183) );
XOR2_X1 U1098 ( .A(n1380), .B(n1381), .Z(n1188) );
XOR2_X1 U1099 ( .A(n1125), .B(n1370), .Z(n1381) );
XOR2_X1 U1100 ( .A(G104), .B(G107), .Z(n1370) );
XNOR2_X1 U1101 ( .A(n1253), .B(n1382), .ZN(n1125) );
NOR2_X1 U1102 ( .A1(KEYINPUT51), .A2(n1383), .ZN(n1382) );
NOR3_X1 U1103 ( .A1(n1384), .A2(n1385), .A3(n1386), .ZN(n1383) );
AND2_X1 U1104 ( .A1(n1387), .A2(G146), .ZN(n1386) );
NOR3_X1 U1105 ( .A1(G146), .A2(KEYINPUT30), .A3(n1387), .ZN(n1385) );
NAND2_X1 U1106 ( .A1(KEYINPUT42), .A2(n1236), .ZN(n1387) );
INV_X1 U1107 ( .A(G143), .ZN(n1236) );
AND2_X1 U1108 ( .A1(G143), .A2(KEYINPUT30), .ZN(n1384) );
INV_X1 U1109 ( .A(G128), .ZN(n1253) );
XNOR2_X1 U1110 ( .A(G101), .B(KEYINPUT58), .ZN(n1380) );
XNOR2_X1 U1111 ( .A(n1189), .B(n1175), .ZN(n1378) );
XOR2_X1 U1112 ( .A(n1388), .B(G131), .Z(n1175) );
NAND2_X1 U1113 ( .A1(n1389), .A2(n1390), .ZN(n1388) );
OR2_X1 U1114 ( .A1(n1123), .A2(G134), .ZN(n1390) );
XOR2_X1 U1115 ( .A(n1121), .B(KEYINPUT59), .Z(n1389) );
NAND2_X1 U1116 ( .A1(G134), .A2(n1123), .ZN(n1121) );
INV_X1 U1117 ( .A(G137), .ZN(n1123) );
NAND2_X1 U1118 ( .A1(G227), .A2(n1063), .ZN(n1189) );
INV_X1 U1119 ( .A(G953), .ZN(n1063) );
endmodule


