//Key = 0110011011100000110100010100001000101001100011000100101110011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326;

NAND2_X1 U729 ( .A1(n1004), .A2(n1005), .ZN(G9) );
NAND2_X1 U730 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND2_X1 U731 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
OR2_X1 U732 ( .A1(KEYINPUT21), .A2(KEYINPUT60), .ZN(n1009) );
NAND3_X1 U733 ( .A1(n1010), .A2(n1011), .A3(KEYINPUT60), .ZN(n1004) );
OR2_X1 U734 ( .A1(n1008), .A2(KEYINPUT21), .ZN(n1011) );
NAND2_X1 U735 ( .A1(n1012), .A2(n1008), .ZN(n1010) );
OR2_X1 U736 ( .A1(n1007), .A2(KEYINPUT21), .ZN(n1012) );
NOR2_X1 U737 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR3_X1 U738 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
INV_X1 U739 ( .A(G952), .ZN(n1016) );
NAND3_X1 U740 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1015) );
NAND2_X1 U741 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U742 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND4_X1 U743 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
NAND2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1027) );
INV_X1 U746 ( .A(n1030), .ZN(n1032) );
NAND2_X1 U747 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
INV_X1 U748 ( .A(n1035), .ZN(n1034) );
NAND3_X1 U749 ( .A1(n1030), .A2(n1036), .A3(n1033), .ZN(n1023) );
NAND2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U751 ( .A1(n1026), .A2(n1039), .ZN(n1038) );
NAND2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U753 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
INV_X1 U754 ( .A(n1044), .ZN(n1040) );
NAND2_X1 U755 ( .A1(n1025), .A2(n1045), .ZN(n1037) );
NAND2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
INV_X1 U758 ( .A(n1050), .ZN(n1046) );
INV_X1 U759 ( .A(n1051), .ZN(n1021) );
NOR3_X1 U760 ( .A1(n1052), .A2(G953), .A3(n1053), .ZN(n1013) );
INV_X1 U761 ( .A(n1018), .ZN(n1053) );
NAND4_X1 U762 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1018) );
NOR4_X1 U763 ( .A1(n1042), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1057) );
AND2_X1 U764 ( .A1(n1061), .A2(G475), .ZN(n1059) );
AND2_X1 U765 ( .A1(n1026), .A2(n1062), .ZN(n1056) );
XNOR2_X1 U766 ( .A(G469), .B(n1063), .ZN(n1055) );
NOR2_X1 U767 ( .A1(KEYINPUT42), .A2(n1064), .ZN(n1063) );
XNOR2_X1 U768 ( .A(n1065), .B(n1066), .ZN(n1054) );
XNOR2_X1 U769 ( .A(G952), .B(KEYINPUT5), .ZN(n1052) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(G72) );
NAND2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
OR2_X1 U772 ( .A1(n1019), .A2(G227), .ZN(n1070) );
NAND3_X1 U773 ( .A1(G953), .A2(n1071), .A3(n1072), .ZN(n1067) );
INV_X1 U774 ( .A(n1069), .ZN(n1072) );
XNOR2_X1 U775 ( .A(n1073), .B(n1074), .ZN(n1069) );
NOR2_X1 U776 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XOR2_X1 U777 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U778 ( .A(n1079), .B(n1080), .Z(n1078) );
XNOR2_X1 U779 ( .A(G137), .B(n1081), .ZN(n1080) );
NOR2_X1 U780 ( .A1(G131), .A2(KEYINPUT33), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1082), .B(n1083), .Z(n1077) );
NAND3_X1 U782 ( .A1(n1084), .A2(n1019), .A3(KEYINPUT6), .ZN(n1073) );
NAND3_X1 U783 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
XOR2_X1 U784 ( .A(n1088), .B(KEYINPUT57), .Z(n1087) );
NAND2_X1 U785 ( .A1(G900), .A2(G227), .ZN(n1071) );
XOR2_X1 U786 ( .A(n1089), .B(n1090), .Z(G69) );
NAND2_X1 U787 ( .A1(G953), .A2(n1091), .ZN(n1090) );
NAND2_X1 U788 ( .A1(G898), .A2(G224), .ZN(n1091) );
NAND3_X1 U789 ( .A1(KEYINPUT1), .A2(n1092), .A3(n1093), .ZN(n1089) );
XNOR2_X1 U790 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U791 ( .A1(KEYINPUT53), .A2(n1096), .ZN(n1095) );
NAND2_X1 U792 ( .A1(G953), .A2(n1097), .ZN(n1092) );
NOR2_X1 U793 ( .A1(n1098), .A2(n1099), .ZN(G66) );
XOR2_X1 U794 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U795 ( .A1(n1066), .A2(n1102), .ZN(n1100) );
NOR2_X1 U796 ( .A1(n1098), .A2(n1103), .ZN(G63) );
XOR2_X1 U797 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR3_X1 U798 ( .A1(n1102), .A2(KEYINPUT11), .A3(n1106), .ZN(n1104) );
NOR2_X1 U799 ( .A1(n1098), .A2(n1107), .ZN(G60) );
XOR2_X1 U800 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND3_X1 U801 ( .A1(n1110), .A2(n1111), .A3(G475), .ZN(n1109) );
NAND2_X1 U802 ( .A1(KEYINPUT23), .A2(n1102), .ZN(n1111) );
NAND2_X1 U803 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
INV_X1 U804 ( .A(KEYINPUT23), .ZN(n1113) );
OR2_X1 U805 ( .A1(n1114), .A2(n1017), .ZN(n1112) );
XNOR2_X1 U806 ( .A(G104), .B(n1115), .ZN(G6) );
NOR2_X1 U807 ( .A1(n1098), .A2(n1116), .ZN(G57) );
XOR2_X1 U808 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U809 ( .A(KEYINPUT47), .B(n1119), .Z(n1118) );
NOR2_X1 U810 ( .A1(n1120), .A2(n1102), .ZN(n1119) );
NOR2_X1 U811 ( .A1(n1098), .A2(n1121), .ZN(G54) );
NOR3_X1 U812 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
NOR2_X1 U813 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U814 ( .A1(KEYINPUT46), .A2(n1127), .ZN(n1125) );
XOR2_X1 U815 ( .A(KEYINPUT27), .B(n1128), .Z(n1127) );
NOR3_X1 U816 ( .A1(n1129), .A2(KEYINPUT46), .A3(n1128), .ZN(n1123) );
INV_X1 U817 ( .A(n1126), .ZN(n1129) );
NOR2_X1 U818 ( .A1(n1102), .A2(n1130), .ZN(n1126) );
AND2_X1 U819 ( .A1(n1128), .A2(KEYINPUT46), .ZN(n1122) );
XNOR2_X1 U820 ( .A(n1131), .B(n1132), .ZN(n1128) );
XOR2_X1 U821 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U822 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NAND2_X1 U823 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U824 ( .A(n1139), .B(n1140), .ZN(n1137) );
XOR2_X1 U825 ( .A(n1141), .B(KEYINPUT28), .Z(n1135) );
NAND2_X1 U826 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XNOR2_X1 U827 ( .A(G110), .B(n1139), .ZN(n1143) );
NAND2_X1 U828 ( .A1(KEYINPUT16), .A2(n1144), .ZN(n1139) );
INV_X1 U829 ( .A(G140), .ZN(n1144) );
XNOR2_X1 U830 ( .A(KEYINPUT51), .B(n1145), .ZN(n1131) );
NOR3_X1 U831 ( .A1(KEYINPUT15), .A2(n1146), .A3(n1147), .ZN(n1145) );
NOR3_X1 U832 ( .A1(KEYINPUT59), .A2(n1148), .A3(n1149), .ZN(n1147) );
XOR2_X1 U833 ( .A(n1082), .B(G146), .Z(n1149) );
NOR2_X1 U834 ( .A1(n1150), .A2(n1151), .ZN(n1146) );
INV_X1 U835 ( .A(KEYINPUT59), .ZN(n1151) );
XNOR2_X1 U836 ( .A(G146), .B(n1152), .ZN(n1150) );
NOR2_X1 U837 ( .A1(n1098), .A2(n1153), .ZN(G51) );
XNOR2_X1 U838 ( .A(n1154), .B(n1096), .ZN(n1153) );
XOR2_X1 U839 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U840 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
INV_X1 U841 ( .A(n1159), .ZN(n1157) );
NAND3_X1 U842 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1155) );
NAND2_X1 U843 ( .A1(KEYINPUT49), .A2(n1102), .ZN(n1161) );
NAND2_X1 U844 ( .A1(n1163), .A2(n1017), .ZN(n1102) );
INV_X1 U845 ( .A(n1114), .ZN(n1163) );
NAND2_X1 U846 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
INV_X1 U847 ( .A(KEYINPUT49), .ZN(n1165) );
NAND2_X1 U848 ( .A1(n1114), .A2(n1017), .ZN(n1164) );
NAND4_X1 U849 ( .A1(n1166), .A2(n1094), .A3(n1085), .A4(n1088), .ZN(n1017) );
AND4_X1 U850 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1085) );
NOR3_X1 U851 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
INV_X1 U852 ( .A(n1174), .ZN(n1171) );
AND4_X1 U853 ( .A1(n1115), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1094) );
AND4_X1 U854 ( .A1(n1007), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1177) );
NAND3_X1 U855 ( .A1(n1181), .A2(n1030), .A3(n1182), .ZN(n1007) );
OR2_X1 U856 ( .A1(n1183), .A2(n1029), .ZN(n1176) );
NOR2_X1 U857 ( .A1(n1184), .A2(n1181), .ZN(n1029) );
NAND3_X1 U858 ( .A1(n1182), .A2(n1030), .A3(n1184), .ZN(n1115) );
XOR2_X1 U859 ( .A(n1086), .B(KEYINPUT41), .Z(n1166) );
XOR2_X1 U860 ( .A(G902), .B(KEYINPUT44), .Z(n1114) );
NOR2_X1 U861 ( .A1(n1019), .A2(G952), .ZN(n1098) );
XOR2_X1 U862 ( .A(n1168), .B(n1185), .Z(G48) );
NOR2_X1 U863 ( .A1(KEYINPUT3), .A2(n1186), .ZN(n1185) );
XOR2_X1 U864 ( .A(KEYINPUT22), .B(G146), .Z(n1186) );
NAND3_X1 U865 ( .A1(n1187), .A2(n1050), .A3(n1184), .ZN(n1168) );
XNOR2_X1 U866 ( .A(G143), .B(n1086), .ZN(G45) );
NAND4_X1 U867 ( .A1(n1188), .A2(n1189), .A3(n1050), .A4(n1190), .ZN(n1086) );
XNOR2_X1 U868 ( .A(G140), .B(n1174), .ZN(G42) );
NAND3_X1 U869 ( .A1(n1026), .A2(n1044), .A3(n1191), .ZN(n1174) );
XNOR2_X1 U870 ( .A(G137), .B(n1088), .ZN(G39) );
NAND3_X1 U871 ( .A1(n1187), .A2(n1026), .A3(n1033), .ZN(n1088) );
XOR2_X1 U872 ( .A(G134), .B(n1173), .Z(G36) );
AND3_X1 U873 ( .A1(n1026), .A2(n1181), .A3(n1189), .ZN(n1173) );
XOR2_X1 U874 ( .A(G131), .B(n1172), .Z(G33) );
AND3_X1 U875 ( .A1(n1184), .A2(n1026), .A3(n1189), .ZN(n1172) );
AND4_X1 U876 ( .A1(n1192), .A2(n1044), .A3(n1193), .A4(n1194), .ZN(n1189) );
NOR2_X1 U877 ( .A1(n1195), .A2(n1048), .ZN(n1026) );
XNOR2_X1 U878 ( .A(G128), .B(n1169), .ZN(G30) );
NAND3_X1 U879 ( .A1(n1181), .A2(n1050), .A3(n1187), .ZN(n1169) );
AND3_X1 U880 ( .A1(n1044), .A2(n1194), .A3(n1035), .ZN(n1187) );
XNOR2_X1 U881 ( .A(G101), .B(n1175), .ZN(G3) );
NAND4_X1 U882 ( .A1(n1033), .A2(n1182), .A3(n1192), .A4(n1193), .ZN(n1175) );
XNOR2_X1 U883 ( .A(G125), .B(n1167), .ZN(G27) );
NAND3_X1 U884 ( .A1(n1025), .A2(n1050), .A3(n1191), .ZN(n1167) );
AND4_X1 U885 ( .A1(n1062), .A2(n1184), .A3(n1196), .A4(n1194), .ZN(n1191) );
NAND2_X1 U886 ( .A1(n1197), .A2(n1051), .ZN(n1194) );
NAND3_X1 U887 ( .A1(G902), .A2(n1198), .A3(n1075), .ZN(n1197) );
NOR2_X1 U888 ( .A1(n1019), .A2(G900), .ZN(n1075) );
INV_X1 U889 ( .A(n1199), .ZN(n1184) );
XNOR2_X1 U890 ( .A(G122), .B(n1180), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1200), .A2(n1190), .A3(n1188), .A4(n1201), .ZN(n1180) );
AND2_X1 U892 ( .A1(n1030), .A2(n1025), .ZN(n1201) );
NOR2_X1 U893 ( .A1(n1196), .A2(n1193), .ZN(n1030) );
XNOR2_X1 U894 ( .A(G119), .B(n1179), .ZN(G21) );
NAND4_X1 U895 ( .A1(n1025), .A2(n1033), .A3(n1035), .A4(n1200), .ZN(n1179) );
NOR2_X1 U896 ( .A1(n1062), .A2(n1192), .ZN(n1035) );
XNOR2_X1 U897 ( .A(G116), .B(n1202), .ZN(G18) );
NAND3_X1 U898 ( .A1(n1203), .A2(n1204), .A3(KEYINPUT56), .ZN(n1202) );
XOR2_X1 U899 ( .A(KEYINPUT31), .B(n1181), .Z(n1204) );
NOR2_X1 U900 ( .A1(n1190), .A2(n1205), .ZN(n1181) );
INV_X1 U901 ( .A(n1183), .ZN(n1203) );
XNOR2_X1 U902 ( .A(n1206), .B(n1207), .ZN(G15) );
NOR2_X1 U903 ( .A1(n1199), .A2(n1183), .ZN(n1207) );
NAND4_X1 U904 ( .A1(n1192), .A2(n1025), .A3(n1200), .A4(n1193), .ZN(n1183) );
NOR2_X1 U905 ( .A1(n1208), .A2(n1042), .ZN(n1025) );
INV_X1 U906 ( .A(n1196), .ZN(n1192) );
NAND2_X1 U907 ( .A1(n1205), .A2(n1190), .ZN(n1199) );
XNOR2_X1 U908 ( .A(G110), .B(n1178), .ZN(G12) );
NAND4_X1 U909 ( .A1(n1033), .A2(n1182), .A3(n1062), .A4(n1196), .ZN(n1178) );
XNOR2_X1 U910 ( .A(n1065), .B(n1209), .ZN(n1196) );
NOR2_X1 U911 ( .A1(KEYINPUT26), .A2(n1066), .ZN(n1209) );
NAND2_X1 U912 ( .A1(G217), .A2(n1210), .ZN(n1066) );
OR2_X1 U913 ( .A1(n1101), .A2(G902), .ZN(n1065) );
XNOR2_X1 U914 ( .A(n1211), .B(n1212), .ZN(n1101) );
XOR2_X1 U915 ( .A(G137), .B(n1213), .Z(n1212) );
AND3_X1 U916 ( .A1(G221), .A2(n1019), .A3(G234), .ZN(n1213) );
NAND3_X1 U917 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1211) );
OR2_X1 U918 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U919 ( .A1(KEYINPUT7), .A2(n1219), .ZN(n1215) );
NAND2_X1 U920 ( .A1(n1220), .A2(n1217), .ZN(n1219) );
XNOR2_X1 U921 ( .A(KEYINPUT52), .B(n1218), .ZN(n1220) );
NAND2_X1 U922 ( .A1(n1221), .A2(n1222), .ZN(n1214) );
INV_X1 U923 ( .A(KEYINPUT7), .ZN(n1222) );
NAND2_X1 U924 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
OR2_X1 U925 ( .A1(n1218), .A2(KEYINPUT52), .ZN(n1224) );
NAND3_X1 U926 ( .A1(n1217), .A2(n1218), .A3(KEYINPUT52), .ZN(n1223) );
XNOR2_X1 U927 ( .A(G146), .B(n1225), .ZN(n1218) );
NOR2_X1 U928 ( .A1(KEYINPUT24), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U929 ( .A(G140), .B(n1227), .ZN(n1226) );
NAND2_X1 U930 ( .A1(KEYINPUT34), .A2(n1228), .ZN(n1227) );
XOR2_X1 U931 ( .A(n1229), .B(n1140), .Z(n1217) );
NAND4_X1 U932 ( .A1(KEYINPUT10), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1229) );
NAND3_X1 U933 ( .A1(KEYINPUT36), .A2(n1233), .A3(G128), .ZN(n1232) );
OR2_X1 U934 ( .A1(n1233), .A2(G128), .ZN(n1231) );
NOR2_X1 U935 ( .A1(KEYINPUT58), .A2(n1234), .ZN(n1233) );
OR2_X1 U936 ( .A1(G119), .A2(KEYINPUT36), .ZN(n1230) );
INV_X1 U937 ( .A(n1193), .ZN(n1062) );
XOR2_X1 U938 ( .A(n1235), .B(n1120), .Z(n1193) );
INV_X1 U939 ( .A(G472), .ZN(n1120) );
OR2_X1 U940 ( .A1(n1117), .A2(G902), .ZN(n1235) );
XNOR2_X1 U941 ( .A(n1236), .B(n1237), .ZN(n1117) );
XOR2_X1 U942 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U943 ( .A(n1134), .B(n1240), .Z(n1239) );
XOR2_X1 U944 ( .A(n1241), .B(n1242), .Z(n1236) );
AND3_X1 U945 ( .A1(G210), .A2(n1019), .A3(n1243), .ZN(n1242) );
XNOR2_X1 U946 ( .A(KEYINPUT4), .B(KEYINPUT38), .ZN(n1241) );
AND2_X1 U947 ( .A1(n1200), .A2(n1044), .ZN(n1182) );
NOR2_X1 U948 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
AND2_X1 U949 ( .A1(G221), .A2(n1210), .ZN(n1042) );
NAND2_X1 U950 ( .A1(G234), .A2(n1244), .ZN(n1210) );
XNOR2_X1 U951 ( .A(KEYINPUT45), .B(n1245), .ZN(n1244) );
INV_X1 U952 ( .A(n1208), .ZN(n1043) );
XOR2_X1 U953 ( .A(n1064), .B(n1130), .Z(n1208) );
INV_X1 U954 ( .A(G469), .ZN(n1130) );
NAND2_X1 U955 ( .A1(n1246), .A2(n1245), .ZN(n1064) );
XOR2_X1 U956 ( .A(n1247), .B(n1248), .Z(n1246) );
XNOR2_X1 U957 ( .A(n1249), .B(n1152), .ZN(n1248) );
XOR2_X1 U958 ( .A(n1082), .B(n1148), .Z(n1152) );
NAND3_X1 U959 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1148) );
NAND2_X1 U960 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND2_X1 U961 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XNOR2_X1 U962 ( .A(n1257), .B(G101), .ZN(n1253) );
NAND4_X1 U963 ( .A1(n1258), .A2(n1256), .A3(n1255), .A4(n1259), .ZN(n1251) );
INV_X1 U964 ( .A(KEYINPUT32), .ZN(n1256) );
XNOR2_X1 U965 ( .A(KEYINPUT14), .B(G101), .ZN(n1258) );
OR2_X1 U966 ( .A1(n1259), .A2(n1255), .ZN(n1250) );
XNOR2_X1 U967 ( .A(G104), .B(n1008), .ZN(n1255) );
INV_X1 U968 ( .A(KEYINPUT61), .ZN(n1259) );
NAND2_X1 U969 ( .A1(n1260), .A2(n1261), .ZN(n1082) );
NAND2_X1 U970 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XOR2_X1 U971 ( .A(KEYINPUT62), .B(n1264), .Z(n1262) );
NAND2_X1 U972 ( .A1(n1265), .A2(G143), .ZN(n1260) );
XOR2_X1 U973 ( .A(KEYINPUT12), .B(n1264), .Z(n1265) );
XNOR2_X1 U974 ( .A(n1266), .B(KEYINPUT25), .ZN(n1264) );
XOR2_X1 U975 ( .A(n1134), .B(n1267), .Z(n1247) );
XNOR2_X1 U976 ( .A(n1140), .B(n1142), .ZN(n1267) );
INV_X1 U977 ( .A(n1138), .ZN(n1142) );
NAND2_X1 U978 ( .A1(G227), .A2(n1019), .ZN(n1138) );
XOR2_X1 U979 ( .A(n1268), .B(n1269), .Z(n1134) );
XOR2_X1 U980 ( .A(KEYINPUT0), .B(G137), .Z(n1269) );
XOR2_X1 U981 ( .A(n1270), .B(G131), .Z(n1268) );
NAND2_X1 U982 ( .A1(KEYINPUT39), .A2(n1079), .ZN(n1270) );
XNOR2_X1 U983 ( .A(G134), .B(KEYINPUT55), .ZN(n1079) );
AND2_X1 U984 ( .A1(n1050), .A2(n1271), .ZN(n1200) );
NAND2_X1 U985 ( .A1(n1051), .A2(n1272), .ZN(n1271) );
NAND4_X1 U986 ( .A1(G953), .A2(G902), .A3(n1198), .A4(n1097), .ZN(n1272) );
INV_X1 U987 ( .A(G898), .ZN(n1097) );
NAND3_X1 U988 ( .A1(n1198), .A2(n1019), .A3(G952), .ZN(n1051) );
NAND2_X1 U989 ( .A1(G237), .A2(G234), .ZN(n1198) );
NOR2_X1 U990 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
AND2_X1 U991 ( .A1(G214), .A2(n1273), .ZN(n1048) );
INV_X1 U992 ( .A(n1195), .ZN(n1049) );
XNOR2_X1 U993 ( .A(n1274), .B(n1162), .ZN(n1195) );
AND2_X1 U994 ( .A1(G210), .A2(n1273), .ZN(n1162) );
NAND2_X1 U995 ( .A1(n1245), .A2(n1243), .ZN(n1273) );
NAND3_X1 U996 ( .A1(n1275), .A2(n1245), .A3(n1276), .ZN(n1274) );
NAND2_X1 U997 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U998 ( .A1(n1279), .A2(n1159), .ZN(n1278) );
XNOR2_X1 U999 ( .A(KEYINPUT30), .B(n1096), .ZN(n1277) );
NAND3_X1 U1000 ( .A1(n1280), .A2(n1159), .A3(n1279), .ZN(n1275) );
XNOR2_X1 U1001 ( .A(KEYINPUT18), .B(n1158), .ZN(n1279) );
AND2_X1 U1002 ( .A1(n1281), .A2(n1282), .ZN(n1158) );
NAND2_X1 U1003 ( .A1(G224), .A2(n1019), .ZN(n1282) );
XNOR2_X1 U1004 ( .A(G125), .B(n1240), .ZN(n1281) );
NAND3_X1 U1005 ( .A1(n1283), .A2(n1019), .A3(G224), .ZN(n1159) );
XNOR2_X1 U1006 ( .A(n1228), .B(n1240), .ZN(n1283) );
XNOR2_X1 U1007 ( .A(n1266), .B(n1284), .ZN(n1240) );
NOR3_X1 U1008 ( .A1(n1285), .A2(KEYINPUT43), .A3(n1286), .ZN(n1284) );
NOR2_X1 U1009 ( .A1(G143), .A2(n1287), .ZN(n1286) );
XOR2_X1 U1010 ( .A(KEYINPUT35), .B(n1288), .Z(n1287) );
XOR2_X1 U1011 ( .A(KEYINPUT13), .B(n1289), .Z(n1285) );
AND2_X1 U1012 ( .A1(n1288), .A2(G143), .ZN(n1289) );
XOR2_X1 U1013 ( .A(G146), .B(KEYINPUT19), .Z(n1288) );
INV_X1 U1014 ( .A(G128), .ZN(n1266) );
XNOR2_X1 U1015 ( .A(KEYINPUT50), .B(n1096), .ZN(n1280) );
XOR2_X1 U1016 ( .A(n1290), .B(n1291), .Z(n1096) );
XNOR2_X1 U1017 ( .A(n1140), .B(n1292), .ZN(n1291) );
XNOR2_X1 U1018 ( .A(n1257), .B(G122), .ZN(n1292) );
INV_X1 U1019 ( .A(KEYINPUT14), .ZN(n1257) );
INV_X1 U1020 ( .A(G110), .ZN(n1140) );
XOR2_X1 U1021 ( .A(n1238), .B(n1293), .Z(n1290) );
NOR2_X1 U1022 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XOR2_X1 U1023 ( .A(n1296), .B(KEYINPUT63), .Z(n1295) );
NAND2_X1 U1024 ( .A1(n1297), .A2(n1008), .ZN(n1296) );
NOR2_X1 U1025 ( .A1(n1298), .A2(n1297), .ZN(n1294) );
XOR2_X1 U1026 ( .A(G104), .B(KEYINPUT37), .Z(n1297) );
XNOR2_X1 U1027 ( .A(G107), .B(KEYINPUT29), .ZN(n1298) );
XOR2_X1 U1028 ( .A(n1299), .B(n1300), .Z(n1238) );
XNOR2_X1 U1029 ( .A(n1234), .B(G116), .ZN(n1300) );
INV_X1 U1030 ( .A(G119), .ZN(n1234) );
XNOR2_X1 U1031 ( .A(G113), .B(G101), .ZN(n1299) );
NOR2_X1 U1032 ( .A1(n1190), .A2(n1188), .ZN(n1033) );
INV_X1 U1033 ( .A(n1205), .ZN(n1188) );
XOR2_X1 U1034 ( .A(n1060), .B(KEYINPUT54), .Z(n1205) );
XOR2_X1 U1035 ( .A(n1301), .B(n1106), .Z(n1060) );
INV_X1 U1036 ( .A(G478), .ZN(n1106) );
OR2_X1 U1037 ( .A1(n1105), .A2(G902), .ZN(n1301) );
XNOR2_X1 U1038 ( .A(n1302), .B(n1303), .ZN(n1105) );
XOR2_X1 U1039 ( .A(n1304), .B(n1305), .Z(n1303) );
NAND3_X1 U1040 ( .A1(G234), .A2(n1019), .A3(G217), .ZN(n1305) );
NAND2_X1 U1041 ( .A1(KEYINPUT9), .A2(n1306), .ZN(n1304) );
XOR2_X1 U1042 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1043 ( .A(G116), .B(n1008), .ZN(n1308) );
INV_X1 U1044 ( .A(G107), .ZN(n1008) );
XOR2_X1 U1045 ( .A(KEYINPUT8), .B(G122), .Z(n1307) );
XNOR2_X1 U1046 ( .A(G128), .B(n1309), .ZN(n1302) );
XNOR2_X1 U1047 ( .A(n1263), .B(G134), .ZN(n1309) );
NAND3_X1 U1048 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1190) );
INV_X1 U1049 ( .A(n1058), .ZN(n1312) );
NOR2_X1 U1050 ( .A1(n1061), .A2(G475), .ZN(n1058) );
OR2_X1 U1051 ( .A1(G475), .A2(KEYINPUT2), .ZN(n1311) );
NAND3_X1 U1052 ( .A1(G475), .A2(n1061), .A3(KEYINPUT2), .ZN(n1310) );
NAND2_X1 U1053 ( .A1(n1245), .A2(n1108), .ZN(n1061) );
NAND3_X1 U1054 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1108) );
NAND2_X1 U1055 ( .A1(KEYINPUT20), .A2(n1316), .ZN(n1315) );
OR3_X1 U1056 ( .A1(n1316), .A2(KEYINPUT20), .A3(n1317), .ZN(n1314) );
NAND2_X1 U1057 ( .A1(n1317), .A2(n1318), .ZN(n1313) );
NAND2_X1 U1058 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
INV_X1 U1059 ( .A(KEYINPUT20), .ZN(n1320) );
XOR2_X1 U1060 ( .A(n1316), .B(KEYINPUT40), .Z(n1319) );
XOR2_X1 U1061 ( .A(n1321), .B(n1322), .Z(n1316) );
XNOR2_X1 U1062 ( .A(n1263), .B(G131), .ZN(n1322) );
INV_X1 U1063 ( .A(G143), .ZN(n1263) );
XNOR2_X1 U1064 ( .A(n1083), .B(n1323), .ZN(n1321) );
AND3_X1 U1065 ( .A1(G214), .A2(n1019), .A3(n1243), .ZN(n1323) );
INV_X1 U1066 ( .A(G237), .ZN(n1243) );
INV_X1 U1067 ( .A(G953), .ZN(n1019) );
XNOR2_X1 U1068 ( .A(n1228), .B(n1249), .ZN(n1083) );
XOR2_X1 U1069 ( .A(G140), .B(G146), .Z(n1249) );
INV_X1 U1070 ( .A(G125), .ZN(n1228) );
XNOR2_X1 U1071 ( .A(n1324), .B(n1325), .ZN(n1317) );
XOR2_X1 U1072 ( .A(G122), .B(n1326), .Z(n1325) );
NOR2_X1 U1073 ( .A1(G104), .A2(KEYINPUT48), .ZN(n1326) );
NAND2_X1 U1074 ( .A1(KEYINPUT17), .A2(n1206), .ZN(n1324) );
INV_X1 U1075 ( .A(G113), .ZN(n1206) );
INV_X1 U1076 ( .A(G902), .ZN(n1245) );
endmodule


