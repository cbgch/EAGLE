//Key = 1011011011010111001100100010100111000111001010101000001001000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;

XOR2_X1 U722 ( .A(n1025), .B(n1026), .Z(G9) );
NAND2_X1 U723 ( .A1(KEYINPUT39), .A2(G107), .ZN(n1026) );
NOR2_X1 U724 ( .A1(n1027), .A2(n1028), .ZN(G75) );
NOR3_X1 U725 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND3_X1 U726 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1029) );
NAND2_X1 U727 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U728 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND4_X1 U729 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1038) );
OR2_X1 U730 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U731 ( .A1(n1045), .A2(n1046), .ZN(n1037) );
NAND2_X1 U732 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U733 ( .A1(n1041), .A2(n1049), .A3(n1039), .ZN(n1048) );
NAND2_X1 U734 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U735 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U736 ( .A1(n1040), .A2(n1054), .ZN(n1047) );
NAND2_X1 U737 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U738 ( .A1(n1039), .A2(n1057), .ZN(n1056) );
NAND2_X1 U739 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U740 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U741 ( .A1(n1041), .A2(n1062), .ZN(n1055) );
NAND2_X1 U742 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U743 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
INV_X1 U744 ( .A(n1067), .ZN(n1035) );
NOR3_X1 U745 ( .A1(n1068), .A2(G953), .A3(G952), .ZN(n1027) );
INV_X1 U746 ( .A(n1032), .ZN(n1068) );
NAND4_X1 U747 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1032) );
NOR4_X1 U748 ( .A1(n1065), .A2(n1052), .A3(n1073), .A4(n1074), .ZN(n1072) );
XNOR2_X1 U749 ( .A(G478), .B(n1075), .ZN(n1074) );
NOR2_X1 U750 ( .A1(n1076), .A2(KEYINPUT41), .ZN(n1075) );
XOR2_X1 U751 ( .A(n1053), .B(KEYINPUT57), .Z(n1073) );
INV_X1 U752 ( .A(n1077), .ZN(n1052) );
NOR2_X1 U753 ( .A1(n1078), .A2(n1079), .ZN(n1071) );
XOR2_X1 U754 ( .A(KEYINPUT27), .B(n1061), .Z(n1079) );
XOR2_X1 U755 ( .A(KEYINPUT60), .B(n1080), .Z(n1070) );
NOR2_X1 U756 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U757 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
INV_X1 U758 ( .A(n1085), .ZN(n1081) );
XOR2_X1 U759 ( .A(n1086), .B(n1087), .Z(n1069) );
NAND2_X1 U760 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
XNOR2_X1 U761 ( .A(KEYINPUT51), .B(KEYINPUT24), .ZN(n1088) );
XOR2_X1 U762 ( .A(n1090), .B(n1091), .Z(G72) );
NOR2_X1 U763 ( .A1(n1092), .A2(n1033), .ZN(n1091) );
AND2_X1 U764 ( .A1(G227), .A2(G900), .ZN(n1092) );
NAND2_X1 U765 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U766 ( .A1(n1095), .A2(n1033), .ZN(n1094) );
XOR2_X1 U767 ( .A(n1031), .B(n1096), .Z(n1095) );
NAND3_X1 U768 ( .A1(n1096), .A2(G900), .A3(G953), .ZN(n1093) );
AND2_X1 U769 ( .A1(n1097), .A2(KEYINPUT33), .ZN(n1096) );
XOR2_X1 U770 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U771 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND3_X1 U772 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NAND2_X1 U773 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
INV_X1 U774 ( .A(KEYINPUT62), .ZN(n1106) );
NAND2_X1 U775 ( .A1(KEYINPUT62), .A2(G125), .ZN(n1102) );
NAND3_X1 U776 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1100) );
NAND2_X1 U777 ( .A1(KEYINPUT21), .A2(n1110), .ZN(n1109) );
OR3_X1 U778 ( .A1(n1110), .A2(KEYINPUT21), .A3(n1111), .ZN(n1108) );
NAND2_X1 U779 ( .A1(n1111), .A2(n1112), .ZN(n1107) );
NAND2_X1 U780 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
INV_X1 U781 ( .A(KEYINPUT21), .ZN(n1114) );
XOR2_X1 U782 ( .A(KEYINPUT6), .B(n1110), .Z(n1113) );
XNOR2_X1 U783 ( .A(n1115), .B(KEYINPUT3), .ZN(n1111) );
XOR2_X1 U784 ( .A(n1116), .B(n1117), .Z(G69) );
NOR3_X1 U785 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1117) );
XOR2_X1 U786 ( .A(n1121), .B(n1122), .Z(n1116) );
NOR3_X1 U787 ( .A1(n1123), .A2(KEYINPUT20), .A3(n1124), .ZN(n1122) );
INV_X1 U788 ( .A(n1030), .ZN(n1124) );
XOR2_X1 U789 ( .A(KEYINPUT43), .B(G953), .Z(n1123) );
NAND2_X1 U790 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
OR2_X1 U791 ( .A1(n1033), .A2(G224), .ZN(n1126) );
INV_X1 U792 ( .A(n1120), .ZN(n1125) );
NOR2_X1 U793 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XOR2_X1 U794 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U795 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NOR2_X1 U796 ( .A1(n1127), .A2(n1133), .ZN(G63) );
XOR2_X1 U797 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U798 ( .A1(KEYINPUT25), .A2(n1136), .ZN(n1135) );
NAND2_X1 U799 ( .A1(n1131), .A2(G478), .ZN(n1134) );
NOR2_X1 U800 ( .A1(n1127), .A2(n1137), .ZN(G60) );
XOR2_X1 U801 ( .A(n1138), .B(n1139), .Z(n1137) );
XNOR2_X1 U802 ( .A(KEYINPUT15), .B(n1140), .ZN(n1139) );
NAND2_X1 U803 ( .A1(n1131), .A2(G475), .ZN(n1138) );
XOR2_X1 U804 ( .A(n1141), .B(n1142), .Z(G6) );
NOR2_X1 U805 ( .A1(G104), .A2(KEYINPUT58), .ZN(n1142) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1143), .ZN(G57) );
XOR2_X1 U807 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U808 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U809 ( .A1(KEYINPUT59), .A2(n1148), .ZN(n1147) );
XOR2_X1 U810 ( .A(n1149), .B(n1150), .Z(n1148) );
AND2_X1 U811 ( .A1(G472), .A2(n1131), .ZN(n1150) );
NAND2_X1 U812 ( .A1(KEYINPUT11), .A2(n1151), .ZN(n1149) );
NOR2_X1 U813 ( .A1(KEYINPUT40), .A2(n1152), .ZN(n1146) );
XOR2_X1 U814 ( .A(n1153), .B(KEYINPUT23), .Z(n1144) );
NOR2_X1 U815 ( .A1(n1127), .A2(n1154), .ZN(G54) );
XOR2_X1 U816 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U817 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U818 ( .A1(n1131), .A2(G469), .ZN(n1157) );
INV_X1 U819 ( .A(n1159), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1160), .B(n1161), .Z(n1155) );
NOR2_X1 U821 ( .A1(KEYINPUT55), .A2(n1098), .ZN(n1161) );
NOR3_X1 U822 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1160) );
NOR3_X1 U823 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1164) );
AND2_X1 U824 ( .A1(n1165), .A2(n1167), .ZN(n1163) );
XNOR2_X1 U825 ( .A(n1168), .B(KEYINPUT10), .ZN(n1167) );
NAND2_X1 U826 ( .A1(G110), .A2(n1169), .ZN(n1168) );
INV_X1 U827 ( .A(n1170), .ZN(n1162) );
NOR2_X1 U828 ( .A1(n1127), .A2(n1171), .ZN(G51) );
XOR2_X1 U829 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR4_X1 U830 ( .A1(n1174), .A2(n1175), .A3(KEYINPUT63), .A4(n1176), .ZN(n1172) );
INV_X1 U831 ( .A(G210), .ZN(n1176) );
NOR2_X1 U832 ( .A1(KEYINPUT18), .A2(n1177), .ZN(n1175) );
NOR3_X1 U833 ( .A1(n1031), .A2(n1178), .A3(n1030), .ZN(n1177) );
AND2_X1 U834 ( .A1(n1159), .A2(KEYINPUT18), .ZN(n1174) );
NAND2_X1 U835 ( .A1(G902), .A2(n1179), .ZN(n1159) );
OR2_X1 U836 ( .A1(n1031), .A2(n1030), .ZN(n1179) );
NAND4_X1 U837 ( .A1(n1180), .A2(n1141), .A3(n1181), .A4(n1182), .ZN(n1030) );
AND4_X1 U838 ( .A1(n1025), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1182) );
NAND3_X1 U839 ( .A1(n1044), .A2(n1186), .A3(n1041), .ZN(n1025) );
NAND2_X1 U840 ( .A1(n1187), .A2(n1188), .ZN(n1181) );
NAND2_X1 U841 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U842 ( .A1(n1045), .A2(n1191), .ZN(n1190) );
NAND2_X1 U843 ( .A1(n1192), .A2(n1041), .ZN(n1189) );
NAND3_X1 U844 ( .A1(n1186), .A2(n1043), .A3(n1041), .ZN(n1141) );
NAND2_X1 U845 ( .A1(n1193), .A2(n1194), .ZN(n1180) );
XOR2_X1 U846 ( .A(n1195), .B(KEYINPUT48), .Z(n1193) );
NAND4_X1 U847 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1031) );
NOR4_X1 U848 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NAND2_X1 U849 ( .A1(n1194), .A2(n1204), .ZN(n1198) );
NAND2_X1 U850 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U851 ( .A1(n1207), .A2(n1192), .ZN(n1206) );
XOR2_X1 U852 ( .A(KEYINPUT14), .B(n1208), .Z(n1205) );
AND2_X1 U853 ( .A1(n1044), .A2(n1209), .ZN(n1208) );
NOR2_X1 U854 ( .A1(n1033), .A2(G952), .ZN(n1127) );
XOR2_X1 U855 ( .A(n1210), .B(n1196), .Z(G48) );
NAND3_X1 U856 ( .A1(n1194), .A2(n1043), .A3(n1209), .ZN(n1196) );
XOR2_X1 U857 ( .A(G143), .B(n1211), .Z(G45) );
NOR3_X1 U858 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
XOR2_X1 U859 ( .A(n1063), .B(KEYINPUT16), .Z(n1213) );
XOR2_X1 U860 ( .A(KEYINPUT26), .B(n1192), .Z(n1212) );
XOR2_X1 U861 ( .A(n1169), .B(n1197), .Z(G42) );
NAND4_X1 U862 ( .A1(n1215), .A2(n1039), .A3(n1043), .A4(n1216), .ZN(n1197) );
XOR2_X1 U863 ( .A(G137), .B(n1203), .Z(G39) );
AND3_X1 U864 ( .A1(n1209), .A2(n1039), .A3(n1045), .ZN(n1203) );
AND3_X1 U865 ( .A1(n1217), .A2(n1216), .A3(n1191), .ZN(n1209) );
XOR2_X1 U866 ( .A(G134), .B(n1202), .Z(G36) );
AND3_X1 U867 ( .A1(n1039), .A2(n1044), .A3(n1207), .ZN(n1202) );
XOR2_X1 U868 ( .A(G131), .B(n1201), .Z(G33) );
AND3_X1 U869 ( .A1(n1039), .A2(n1043), .A3(n1207), .ZN(n1201) );
INV_X1 U870 ( .A(n1214), .ZN(n1207) );
NAND3_X1 U871 ( .A1(n1217), .A2(n1216), .A3(n1218), .ZN(n1214) );
INV_X1 U872 ( .A(n1050), .ZN(n1217) );
NOR2_X1 U873 ( .A1(n1219), .A2(n1065), .ZN(n1039) );
INV_X1 U874 ( .A(n1066), .ZN(n1219) );
XNOR2_X1 U875 ( .A(G128), .B(n1220), .ZN(G30) );
NAND4_X1 U876 ( .A1(n1221), .A2(n1191), .A3(n1222), .A4(n1044), .ZN(n1220) );
NOR2_X1 U877 ( .A1(n1223), .A2(n1063), .ZN(n1222) );
XOR2_X1 U878 ( .A(n1050), .B(KEYINPUT8), .Z(n1221) );
XOR2_X1 U879 ( .A(n1153), .B(n1185), .Z(G3) );
NAND3_X1 U880 ( .A1(n1218), .A2(n1186), .A3(n1045), .ZN(n1185) );
NOR3_X1 U881 ( .A1(n1050), .A2(n1224), .A3(n1063), .ZN(n1186) );
XOR2_X1 U882 ( .A(n1225), .B(n1226), .Z(G27) );
NOR2_X1 U883 ( .A1(n1200), .A2(KEYINPUT50), .ZN(n1226) );
AND4_X1 U884 ( .A1(n1194), .A2(n1043), .A3(n1040), .A4(n1227), .ZN(n1200) );
NOR3_X1 U885 ( .A1(n1228), .A2(n1223), .A3(n1229), .ZN(n1227) );
INV_X1 U886 ( .A(n1216), .ZN(n1223) );
NAND2_X1 U887 ( .A1(n1067), .A2(n1230), .ZN(n1216) );
NAND4_X1 U888 ( .A1(G902), .A2(G953), .A3(n1231), .A4(n1232), .ZN(n1230) );
INV_X1 U889 ( .A(G900), .ZN(n1232) );
XOR2_X1 U890 ( .A(n1233), .B(n1234), .Z(G24) );
NAND3_X1 U891 ( .A1(n1187), .A2(n1041), .A3(n1235), .ZN(n1234) );
XNOR2_X1 U892 ( .A(n1192), .B(KEYINPUT37), .ZN(n1235) );
NOR2_X1 U893 ( .A1(n1061), .A2(n1228), .ZN(n1041) );
INV_X1 U894 ( .A(n1229), .ZN(n1061) );
XNOR2_X1 U895 ( .A(G119), .B(n1236), .ZN(G21) );
NAND4_X1 U896 ( .A1(n1045), .A2(n1191), .A3(n1237), .A4(n1238), .ZN(n1236) );
NAND2_X1 U897 ( .A1(KEYINPUT0), .A2(n1239), .ZN(n1238) );
NAND2_X1 U898 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
INV_X1 U899 ( .A(KEYINPUT0), .ZN(n1241) );
NAND3_X1 U900 ( .A1(n1040), .A2(n1194), .A3(n1224), .ZN(n1240) );
INV_X1 U901 ( .A(n1242), .ZN(n1224) );
NOR2_X1 U902 ( .A1(n1060), .A2(n1229), .ZN(n1191) );
INV_X1 U903 ( .A(n1228), .ZN(n1060) );
XNOR2_X1 U904 ( .A(G116), .B(n1243), .ZN(G18) );
NAND2_X1 U905 ( .A1(KEYINPUT38), .A2(n1244), .ZN(n1243) );
INV_X1 U906 ( .A(n1184), .ZN(n1244) );
NAND3_X1 U907 ( .A1(n1218), .A2(n1044), .A3(n1187), .ZN(n1184) );
NOR2_X1 U908 ( .A1(n1245), .A2(n1246), .ZN(n1044) );
XNOR2_X1 U909 ( .A(G113), .B(n1183), .ZN(G15) );
NAND3_X1 U910 ( .A1(n1218), .A2(n1043), .A3(n1187), .ZN(n1183) );
INV_X1 U911 ( .A(n1239), .ZN(n1187) );
NAND3_X1 U912 ( .A1(n1194), .A2(n1242), .A3(n1040), .ZN(n1239) );
AND2_X1 U913 ( .A1(n1247), .A2(n1077), .ZN(n1040) );
XOR2_X1 U914 ( .A(KEYINPUT9), .B(n1248), .Z(n1247) );
NAND2_X1 U915 ( .A1(n1249), .A2(n1250), .ZN(n1043) );
NAND3_X1 U916 ( .A1(n1246), .A2(n1245), .A3(n1251), .ZN(n1250) );
NAND2_X1 U917 ( .A1(KEYINPUT61), .A2(n1192), .ZN(n1249) );
NOR2_X1 U918 ( .A1(n1246), .A2(n1252), .ZN(n1192) );
INV_X1 U919 ( .A(n1245), .ZN(n1252) );
INV_X1 U920 ( .A(n1058), .ZN(n1218) );
NAND2_X1 U921 ( .A1(n1228), .A2(n1229), .ZN(n1058) );
XOR2_X1 U922 ( .A(G110), .B(n1253), .Z(G12) );
NOR2_X1 U923 ( .A1(n1063), .A2(n1195), .ZN(n1253) );
NAND3_X1 U924 ( .A1(n1045), .A2(n1242), .A3(n1215), .ZN(n1195) );
NOR3_X1 U925 ( .A1(n1228), .A2(n1229), .A3(n1050), .ZN(n1215) );
NAND2_X1 U926 ( .A1(n1254), .A2(n1077), .ZN(n1050) );
NAND2_X1 U927 ( .A1(G221), .A2(n1255), .ZN(n1077) );
XOR2_X1 U928 ( .A(KEYINPUT4), .B(n1248), .Z(n1254) );
INV_X1 U929 ( .A(n1053), .ZN(n1248) );
XOR2_X1 U930 ( .A(n1256), .B(G469), .Z(n1053) );
NAND2_X1 U931 ( .A1(n1257), .A2(n1178), .ZN(n1256) );
XOR2_X1 U932 ( .A(n1258), .B(n1259), .Z(n1257) );
NOR2_X1 U933 ( .A1(KEYINPUT34), .A2(n1260), .ZN(n1259) );
XOR2_X1 U934 ( .A(n1158), .B(n1261), .Z(n1260) );
INV_X1 U935 ( .A(n1098), .ZN(n1261) );
XNOR2_X1 U936 ( .A(n1262), .B(n1263), .ZN(n1098) );
XOR2_X1 U937 ( .A(n1264), .B(n1265), .Z(n1158) );
XOR2_X1 U938 ( .A(n1266), .B(n1267), .Z(n1264) );
NAND2_X1 U939 ( .A1(KEYINPUT31), .A2(n1153), .ZN(n1266) );
NAND3_X1 U940 ( .A1(n1268), .A2(n1269), .A3(n1170), .ZN(n1258) );
NAND2_X1 U941 ( .A1(n1166), .A2(n1165), .ZN(n1170) );
NOR2_X1 U942 ( .A1(n1169), .A2(G110), .ZN(n1166) );
NAND2_X1 U943 ( .A1(n1270), .A2(n1169), .ZN(n1269) );
INV_X1 U944 ( .A(G140), .ZN(n1169) );
XOR2_X1 U945 ( .A(G110), .B(n1271), .Z(n1270) );
NAND3_X1 U946 ( .A1(n1271), .A2(G110), .A3(G140), .ZN(n1268) );
INV_X1 U947 ( .A(n1165), .ZN(n1271) );
NAND2_X1 U948 ( .A1(G227), .A2(n1033), .ZN(n1165) );
XOR2_X1 U949 ( .A(n1272), .B(n1132), .Z(n1229) );
AND2_X1 U950 ( .A1(G217), .A2(n1255), .ZN(n1132) );
NAND2_X1 U951 ( .A1(G234), .A2(n1178), .ZN(n1255) );
NAND2_X1 U952 ( .A1(n1130), .A2(n1178), .ZN(n1272) );
XOR2_X1 U953 ( .A(n1273), .B(n1274), .Z(n1130) );
XOR2_X1 U954 ( .A(KEYINPUT19), .B(G137), .Z(n1274) );
XOR2_X1 U955 ( .A(n1275), .B(n1276), .Z(n1273) );
AND2_X1 U956 ( .A1(n1277), .A2(G221), .ZN(n1276) );
NAND2_X1 U957 ( .A1(KEYINPUT42), .A2(n1278), .ZN(n1275) );
XOR2_X1 U958 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U959 ( .A(n1263), .B(n1281), .Z(n1280) );
XOR2_X1 U960 ( .A(n1282), .B(n1283), .Z(n1281) );
NAND3_X1 U961 ( .A1(n1284), .A2(n1285), .A3(n1104), .ZN(n1283) );
NAND2_X1 U962 ( .A1(n1105), .A2(n1286), .ZN(n1285) );
INV_X1 U963 ( .A(KEYINPUT36), .ZN(n1286) );
NAND2_X1 U964 ( .A1(KEYINPUT36), .A2(G125), .ZN(n1284) );
XOR2_X1 U965 ( .A(G119), .B(n1287), .Z(n1279) );
XOR2_X1 U966 ( .A(KEYINPUT7), .B(G146), .Z(n1287) );
XNOR2_X1 U967 ( .A(n1078), .B(KEYINPUT44), .ZN(n1228) );
XNOR2_X1 U968 ( .A(n1288), .B(G472), .ZN(n1078) );
NAND2_X1 U969 ( .A1(n1289), .A2(n1178), .ZN(n1288) );
XOR2_X1 U970 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U971 ( .A(n1153), .B(n1292), .Z(n1291) );
XNOR2_X1 U972 ( .A(KEYINPUT53), .B(KEYINPUT1), .ZN(n1292) );
XOR2_X1 U973 ( .A(n1151), .B(n1152), .Z(n1290) );
NAND2_X1 U974 ( .A1(G210), .A2(n1293), .ZN(n1152) );
XOR2_X1 U975 ( .A(n1294), .B(n1295), .Z(n1151) );
XOR2_X1 U976 ( .A(n1296), .B(n1265), .Z(n1294) );
XNOR2_X1 U977 ( .A(n1115), .B(n1110), .ZN(n1265) );
XNOR2_X1 U978 ( .A(n1297), .B(G137), .ZN(n1110) );
INV_X1 U979 ( .A(G134), .ZN(n1297) );
NAND2_X1 U980 ( .A1(n1298), .A2(n1067), .ZN(n1242) );
NAND3_X1 U981 ( .A1(n1231), .A2(n1033), .A3(G952), .ZN(n1067) );
NAND3_X1 U982 ( .A1(n1120), .A2(n1231), .A3(G902), .ZN(n1298) );
NAND2_X1 U983 ( .A1(G237), .A2(G234), .ZN(n1231) );
NOR2_X1 U984 ( .A1(G898), .A2(n1033), .ZN(n1120) );
NOR2_X1 U985 ( .A1(n1245), .A2(n1299), .ZN(n1045) );
XOR2_X1 U986 ( .A(n1251), .B(n1246), .Z(n1299) );
XOR2_X1 U987 ( .A(n1076), .B(n1300), .Z(n1246) );
XOR2_X1 U988 ( .A(KEYINPUT2), .B(G478), .Z(n1300) );
NOR2_X1 U989 ( .A1(n1136), .A2(G902), .ZN(n1076) );
XOR2_X1 U990 ( .A(n1301), .B(n1302), .Z(n1136) );
XOR2_X1 U991 ( .A(G107), .B(n1303), .Z(n1302) );
XOR2_X1 U992 ( .A(G122), .B(G116), .Z(n1303) );
XOR2_X1 U993 ( .A(n1304), .B(n1305), .Z(n1301) );
NOR2_X1 U994 ( .A1(KEYINPUT45), .A2(n1306), .ZN(n1305) );
XOR2_X1 U995 ( .A(n1307), .B(G134), .Z(n1306) );
NAND2_X1 U996 ( .A1(KEYINPUT5), .A2(n1308), .ZN(n1307) );
XOR2_X1 U997 ( .A(G143), .B(n1263), .Z(n1308) );
NAND2_X1 U998 ( .A1(n1277), .A2(G217), .ZN(n1304) );
AND2_X1 U999 ( .A1(G234), .A2(n1033), .ZN(n1277) );
INV_X1 U1000 ( .A(KEYINPUT61), .ZN(n1251) );
NAND3_X1 U1001 ( .A1(n1309), .A2(n1310), .A3(n1085), .ZN(n1245) );
NAND2_X1 U1002 ( .A1(n1083), .A2(n1084), .ZN(n1085) );
NAND2_X1 U1003 ( .A1(n1084), .A2(n1311), .ZN(n1310) );
OR3_X1 U1004 ( .A1(n1084), .A2(n1083), .A3(n1311), .ZN(n1309) );
INV_X1 U1005 ( .A(KEYINPUT22), .ZN(n1311) );
AND2_X1 U1006 ( .A1(n1178), .A2(n1140), .ZN(n1083) );
NAND3_X1 U1007 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1140) );
NAND2_X1 U1008 ( .A1(KEYINPUT52), .A2(n1315), .ZN(n1314) );
OR3_X1 U1009 ( .A1(n1315), .A2(KEYINPUT52), .A3(n1316), .ZN(n1313) );
NAND2_X1 U1010 ( .A1(n1316), .A2(n1317), .ZN(n1312) );
NAND2_X1 U1011 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
INV_X1 U1012 ( .A(KEYINPUT52), .ZN(n1319) );
XNOR2_X1 U1013 ( .A(KEYINPUT56), .B(n1315), .ZN(n1318) );
XOR2_X1 U1014 ( .A(n1320), .B(n1321), .Z(n1315) );
NOR2_X1 U1015 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NOR2_X1 U1016 ( .A1(G146), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1017 ( .A(n1225), .B(G140), .Z(n1324) );
INV_X1 U1018 ( .A(G125), .ZN(n1225) );
NOR2_X1 U1019 ( .A1(n1325), .A2(n1210), .ZN(n1322) );
NOR2_X1 U1020 ( .A1(n1105), .A2(n1326), .ZN(n1325) );
INV_X1 U1021 ( .A(n1104), .ZN(n1326) );
NAND2_X1 U1022 ( .A1(G140), .A2(G125), .ZN(n1104) );
NOR2_X1 U1023 ( .A1(G125), .A2(G140), .ZN(n1105) );
NAND3_X1 U1024 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1320) );
NAND2_X1 U1025 ( .A1(KEYINPUT47), .A2(n1330), .ZN(n1329) );
NAND3_X1 U1026 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1328) );
INV_X1 U1027 ( .A(KEYINPUT47), .ZN(n1332) );
OR2_X1 U1028 ( .A1(n1333), .A2(n1331), .ZN(n1327) );
NOR2_X1 U1029 ( .A1(KEYINPUT49), .A2(n1330), .ZN(n1331) );
XOR2_X1 U1030 ( .A(n1115), .B(KEYINPUT29), .Z(n1330) );
XNOR2_X1 U1031 ( .A(G131), .B(KEYINPUT28), .ZN(n1115) );
XNOR2_X1 U1032 ( .A(n1334), .B(n1335), .ZN(n1333) );
NAND2_X1 U1033 ( .A1(G214), .A2(n1293), .ZN(n1334) );
NOR2_X1 U1034 ( .A1(G953), .A2(G237), .ZN(n1293) );
XNOR2_X1 U1035 ( .A(n1336), .B(n1337), .ZN(n1316) );
NOR2_X1 U1036 ( .A1(KEYINPUT30), .A2(G113), .ZN(n1337) );
XOR2_X1 U1037 ( .A(G104), .B(n1233), .Z(n1336) );
INV_X1 U1038 ( .A(G475), .ZN(n1084) );
INV_X1 U1039 ( .A(n1194), .ZN(n1063) );
NOR2_X1 U1040 ( .A1(n1066), .A2(n1065), .ZN(n1194) );
AND2_X1 U1041 ( .A1(G214), .A2(n1338), .ZN(n1065) );
XNOR2_X1 U1042 ( .A(n1087), .B(n1089), .ZN(n1066) );
NAND2_X1 U1043 ( .A1(G210), .A2(n1338), .ZN(n1089) );
NAND2_X1 U1044 ( .A1(n1339), .A2(n1178), .ZN(n1338) );
INV_X1 U1045 ( .A(G237), .ZN(n1339) );
NAND2_X1 U1046 ( .A1(n1340), .A2(n1178), .ZN(n1087) );
INV_X1 U1047 ( .A(G902), .ZN(n1178) );
XOR2_X1 U1048 ( .A(KEYINPUT13), .B(n1173), .Z(n1340) );
XNOR2_X1 U1049 ( .A(n1341), .B(n1342), .ZN(n1173) );
XOR2_X1 U1050 ( .A(n1343), .B(n1344), .Z(n1342) );
NAND3_X1 U1051 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1344) );
INV_X1 U1052 ( .A(n1119), .ZN(n1347) );
NOR3_X1 U1053 ( .A1(n1348), .A2(n1295), .A3(n1349), .ZN(n1119) );
NAND2_X1 U1054 ( .A1(n1118), .A2(n1350), .ZN(n1346) );
INV_X1 U1055 ( .A(KEYINPUT17), .ZN(n1350) );
NAND2_X1 U1056 ( .A1(n1351), .A2(n1352), .ZN(n1118) );
NAND2_X1 U1057 ( .A1(n1353), .A2(n1348), .ZN(n1352) );
XOR2_X1 U1058 ( .A(n1295), .B(n1349), .Z(n1353) );
NAND3_X1 U1059 ( .A1(n1349), .A2(n1295), .A3(n1354), .ZN(n1351) );
INV_X1 U1060 ( .A(n1348), .ZN(n1354) );
NAND2_X1 U1061 ( .A1(n1355), .A2(KEYINPUT17), .ZN(n1345) );
XOR2_X1 U1062 ( .A(n1356), .B(n1349), .Z(n1355) );
XOR2_X1 U1063 ( .A(n1357), .B(n1358), .Z(n1349) );
NOR2_X1 U1064 ( .A1(KEYINPUT12), .A2(n1359), .ZN(n1358) );
XOR2_X1 U1065 ( .A(n1282), .B(KEYINPUT46), .Z(n1359) );
INV_X1 U1066 ( .A(G110), .ZN(n1282) );
XOR2_X1 U1067 ( .A(n1233), .B(KEYINPUT54), .Z(n1357) );
INV_X1 U1068 ( .A(G122), .ZN(n1233) );
NAND2_X1 U1069 ( .A1(n1348), .A2(n1295), .ZN(n1356) );
XNOR2_X1 U1070 ( .A(G113), .B(n1360), .ZN(n1295) );
XOR2_X1 U1071 ( .A(G119), .B(G116), .Z(n1360) );
XOR2_X1 U1072 ( .A(n1153), .B(n1267), .Z(n1348) );
XOR2_X1 U1073 ( .A(G104), .B(G107), .Z(n1267) );
INV_X1 U1074 ( .A(G101), .ZN(n1153) );
NAND2_X1 U1075 ( .A1(G224), .A2(n1033), .ZN(n1343) );
INV_X1 U1076 ( .A(G953), .ZN(n1033) );
XOR2_X1 U1077 ( .A(n1296), .B(G125), .Z(n1341) );
NAND2_X1 U1078 ( .A1(n1361), .A2(n1362), .ZN(n1296) );
NAND2_X1 U1079 ( .A1(n1262), .A2(n1263), .ZN(n1362) );
XOR2_X1 U1080 ( .A(KEYINPUT32), .B(n1363), .Z(n1361) );
NOR2_X1 U1081 ( .A1(n1263), .A2(n1262), .ZN(n1363) );
XOR2_X1 U1082 ( .A(n1335), .B(n1210), .Z(n1262) );
INV_X1 U1083 ( .A(G146), .ZN(n1210) );
INV_X1 U1084 ( .A(G143), .ZN(n1335) );
XOR2_X1 U1085 ( .A(G128), .B(KEYINPUT35), .Z(n1263) );
endmodule


