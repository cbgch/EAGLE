//Key = 0100001010100110011101000010000100010110100011010111000111110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394;

XNOR2_X1 U764 ( .A(G107), .B(n1054), .ZN(G9) );
NOR2_X1 U765 ( .A1(n1055), .A2(n1056), .ZN(G75) );
NOR4_X1 U766 ( .A1(G953), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1056) );
NOR2_X1 U767 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U768 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U769 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U772 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U776 ( .A1(n1078), .A2(n1079), .ZN(n1070) );
NOR2_X1 U777 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR3_X1 U778 ( .A1(n1079), .A2(n1082), .A3(n1073), .ZN(n1066) );
NOR2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR4_X1 U781 ( .A1(n1087), .A2(n1073), .A3(n1069), .A4(n1079), .ZN(n1062) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR3_X1 U783 ( .A1(n1057), .A2(G953), .A3(G952), .ZN(n1055) );
AND4_X1 U784 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1057) );
NOR4_X1 U785 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
XOR2_X1 U786 ( .A(n1098), .B(KEYINPUT54), .Z(n1097) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U788 ( .A(n1101), .B(n1102), .Z(n1096) );
NOR2_X1 U789 ( .A1(G472), .A2(KEYINPUT16), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1104), .ZN(n1092) );
XOR2_X1 U791 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U792 ( .A(G475), .B(n1107), .ZN(n1103) );
NOR2_X1 U793 ( .A1(n1108), .A2(KEYINPUT32), .ZN(n1107) );
XOR2_X1 U794 ( .A(n1109), .B(G478), .Z(n1091) );
XOR2_X1 U795 ( .A(n1110), .B(n1111), .Z(n1090) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(G72) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
INV_X1 U799 ( .A(n1118), .ZN(n1117) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1116) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U802 ( .A(n1123), .B(KEYINPUT52), .Z(n1122) );
NAND2_X1 U803 ( .A1(KEYINPUT55), .A2(n1124), .ZN(n1121) );
XOR2_X1 U804 ( .A(n1125), .B(n1126), .Z(n1119) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1114) );
XOR2_X1 U806 ( .A(KEYINPUT47), .B(n1129), .Z(n1127) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U808 ( .A(n1132), .B(KEYINPUT49), .Z(n1130) );
NOR2_X1 U809 ( .A1(n1133), .A2(n1128), .ZN(n1112) );
AND2_X1 U810 ( .A1(G227), .A2(G900), .ZN(n1133) );
NAND2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(G69) );
NAND2_X1 U812 ( .A1(n1136), .A2(n1128), .ZN(n1135) );
XOR2_X1 U813 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U814 ( .A1(n1139), .A2(G953), .ZN(n1134) );
NAND2_X1 U815 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U816 ( .A1(n1137), .A2(n1142), .ZN(n1141) );
INV_X1 U817 ( .A(G224), .ZN(n1142) );
NAND2_X1 U818 ( .A1(G224), .A2(n1143), .ZN(n1140) );
NAND2_X1 U819 ( .A1(G898), .A2(n1137), .ZN(n1143) );
NAND3_X1 U820 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1137) );
NAND2_X1 U821 ( .A1(G953), .A2(n1147), .ZN(n1146) );
NAND4_X1 U822 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1145) );
NAND2_X1 U823 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U824 ( .A1(KEYINPUT51), .A2(n1154), .ZN(n1150) );
NAND2_X1 U825 ( .A1(n1155), .A2(n1156), .ZN(n1148) );
NAND3_X1 U826 ( .A1(n1157), .A2(n1156), .A3(n1155), .ZN(n1144) );
INV_X1 U827 ( .A(KEYINPUT9), .ZN(n1156) );
NAND3_X1 U828 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1157) );
NAND2_X1 U829 ( .A1(KEYINPUT51), .A2(n1161), .ZN(n1159) );
NAND2_X1 U830 ( .A1(n1162), .A2(n1153), .ZN(n1158) );
INV_X1 U831 ( .A(KEYINPUT51), .ZN(n1153) );
NOR2_X1 U832 ( .A1(n1163), .A2(n1164), .ZN(G66) );
XOR2_X1 U833 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND3_X1 U834 ( .A1(n1167), .A2(n1111), .A3(KEYINPUT45), .ZN(n1165) );
NOR2_X1 U835 ( .A1(n1168), .A2(n1169), .ZN(G63) );
XNOR2_X1 U836 ( .A(n1170), .B(n1171), .ZN(n1169) );
NOR2_X1 U837 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U838 ( .A1(n1174), .A2(n1128), .ZN(n1168) );
XNOR2_X1 U839 ( .A(G952), .B(KEYINPUT6), .ZN(n1174) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1175), .ZN(G60) );
XOR2_X1 U841 ( .A(n1176), .B(n1177), .Z(n1175) );
AND2_X1 U842 ( .A1(G475), .A2(n1167), .ZN(n1176) );
XNOR2_X1 U843 ( .A(G104), .B(n1178), .ZN(G6) );
NOR2_X1 U844 ( .A1(n1163), .A2(n1179), .ZN(G57) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND3_X1 U847 ( .A1(n1184), .A2(n1185), .A3(G472), .ZN(n1183) );
OR2_X1 U848 ( .A1(n1167), .A2(KEYINPUT61), .ZN(n1185) );
NAND2_X1 U849 ( .A1(KEYINPUT61), .A2(n1186), .ZN(n1184) );
NAND2_X1 U850 ( .A1(n1187), .A2(n1059), .ZN(n1186) );
NAND2_X1 U851 ( .A1(n1188), .A2(n1189), .ZN(n1182) );
OR2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XOR2_X1 U853 ( .A(n1192), .B(KEYINPUT0), .Z(n1188) );
NAND2_X1 U854 ( .A1(n1190), .A2(n1191), .ZN(n1192) );
XNOR2_X1 U855 ( .A(n1193), .B(KEYINPUT35), .ZN(n1190) );
XNOR2_X1 U856 ( .A(n1194), .B(n1195), .ZN(n1180) );
NOR2_X1 U857 ( .A1(n1163), .A2(n1196), .ZN(G54) );
XOR2_X1 U858 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U859 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U860 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XOR2_X1 U861 ( .A(KEYINPUT60), .B(n1203), .Z(n1202) );
NOR2_X1 U862 ( .A1(G140), .A2(n1204), .ZN(n1203) );
AND2_X1 U863 ( .A1(G140), .A2(n1204), .ZN(n1201) );
NAND2_X1 U864 ( .A1(KEYINPUT62), .A2(n1205), .ZN(n1199) );
NAND2_X1 U865 ( .A1(n1167), .A2(G469), .ZN(n1205) );
XOR2_X1 U866 ( .A(n1206), .B(n1207), .Z(n1197) );
NOR2_X1 U867 ( .A1(KEYINPUT4), .A2(n1208), .ZN(n1207) );
XOR2_X1 U868 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U869 ( .A(n1194), .B(n1211), .Z(n1210) );
XOR2_X1 U870 ( .A(KEYINPUT41), .B(KEYINPUT3), .Z(n1209) );
NOR2_X1 U871 ( .A1(n1163), .A2(n1212), .ZN(G51) );
XOR2_X1 U872 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U873 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND2_X1 U874 ( .A1(KEYINPUT57), .A2(n1217), .ZN(n1215) );
XOR2_X1 U875 ( .A(n1218), .B(n1219), .Z(n1213) );
XNOR2_X1 U876 ( .A(G125), .B(n1220), .ZN(n1219) );
NOR2_X1 U877 ( .A1(n1106), .A2(n1173), .ZN(n1218) );
INV_X1 U878 ( .A(n1167), .ZN(n1173) );
NOR2_X1 U879 ( .A1(n1187), .A2(n1221), .ZN(n1167) );
INV_X1 U880 ( .A(n1059), .ZN(n1221) );
NAND3_X1 U881 ( .A1(n1138), .A2(n1132), .A3(n1222), .ZN(n1059) );
INV_X1 U882 ( .A(n1131), .ZN(n1222) );
NAND4_X1 U883 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1131) );
NOR4_X1 U884 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1226) );
NOR2_X1 U885 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NOR2_X1 U886 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
NOR2_X1 U887 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NOR2_X1 U888 ( .A1(n1237), .A2(n1065), .ZN(n1233) );
XOR2_X1 U889 ( .A(n1079), .B(KEYINPUT42), .Z(n1237) );
NOR2_X1 U890 ( .A1(n1238), .A2(n1239), .ZN(n1228) );
INV_X1 U891 ( .A(KEYINPUT50), .ZN(n1238) );
NOR4_X1 U892 ( .A1(KEYINPUT50), .A2(n1240), .A3(n1079), .A4(n1241), .ZN(n1227) );
NAND3_X1 U893 ( .A1(n1088), .A2(n1084), .A3(n1081), .ZN(n1240) );
AND4_X1 U894 ( .A1(n1242), .A2(n1178), .A3(n1243), .A4(n1244), .ZN(n1138) );
AND4_X1 U895 ( .A1(n1245), .A2(n1246), .A3(n1054), .A4(n1247), .ZN(n1244) );
NAND4_X1 U896 ( .A1(n1088), .A2(n1084), .A3(n1248), .A4(n1249), .ZN(n1054) );
NOR4_X1 U897 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1243) );
NOR4_X1 U898 ( .A1(n1254), .A2(n1255), .A3(n1075), .A4(n1256), .ZN(n1253) );
INV_X1 U899 ( .A(n1257), .ZN(n1256) );
AND2_X1 U900 ( .A1(n1254), .A2(n1258), .ZN(n1252) );
INV_X1 U901 ( .A(KEYINPUT39), .ZN(n1254) );
NOR3_X1 U902 ( .A1(n1259), .A2(n1260), .A3(n1235), .ZN(n1251) );
INV_X1 U903 ( .A(KEYINPUT5), .ZN(n1259) );
NOR2_X1 U904 ( .A1(KEYINPUT5), .A2(n1261), .ZN(n1250) );
NAND4_X1 U905 ( .A1(n1089), .A2(n1084), .A3(n1248), .A4(n1249), .ZN(n1178) );
NAND2_X1 U906 ( .A1(n1262), .A2(n1089), .ZN(n1242) );
XOR2_X1 U907 ( .A(n1263), .B(KEYINPUT29), .Z(n1187) );
NOR2_X1 U908 ( .A1(n1128), .A2(G952), .ZN(n1163) );
XNOR2_X1 U909 ( .A(G146), .B(n1264), .ZN(G48) );
NAND4_X1 U910 ( .A1(KEYINPUT10), .A2(n1265), .A3(n1089), .A4(n1075), .ZN(n1264) );
XNOR2_X1 U911 ( .A(G143), .B(n1132), .ZN(G45) );
NAND4_X1 U912 ( .A1(n1081), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1132) );
NOR2_X1 U913 ( .A1(n1269), .A2(n1235), .ZN(n1267) );
XOR2_X1 U914 ( .A(G140), .B(n1229), .Z(G42) );
AND3_X1 U915 ( .A1(n1089), .A2(n1080), .A3(n1270), .ZN(n1229) );
XOR2_X1 U916 ( .A(G137), .B(n1271), .Z(G39) );
NOR3_X1 U917 ( .A1(n1065), .A2(n1232), .A3(n1079), .ZN(n1271) );
INV_X1 U918 ( .A(n1272), .ZN(n1079) );
XNOR2_X1 U919 ( .A(G134), .B(n1239), .ZN(G36) );
NAND3_X1 U920 ( .A1(n1081), .A2(n1088), .A3(n1270), .ZN(n1239) );
XOR2_X1 U921 ( .A(n1123), .B(n1225), .Z(G33) );
NAND3_X1 U922 ( .A1(n1089), .A2(n1081), .A3(n1270), .ZN(n1225) );
AND2_X1 U923 ( .A1(n1272), .A2(n1266), .ZN(n1270) );
NOR2_X1 U924 ( .A1(n1076), .A2(n1095), .ZN(n1272) );
INV_X1 U925 ( .A(n1077), .ZN(n1095) );
INV_X1 U926 ( .A(n1236), .ZN(n1089) );
XNOR2_X1 U927 ( .A(G128), .B(n1223), .ZN(G30) );
NAND3_X1 U928 ( .A1(n1088), .A2(n1075), .A3(n1265), .ZN(n1223) );
INV_X1 U929 ( .A(n1232), .ZN(n1265) );
NAND3_X1 U930 ( .A1(n1266), .A2(n1273), .A3(n1274), .ZN(n1232) );
AND2_X1 U931 ( .A1(n1084), .A2(n1241), .ZN(n1266) );
NAND2_X1 U932 ( .A1(n1275), .A2(n1276), .ZN(G3) );
NAND3_X1 U933 ( .A1(KEYINPUT58), .A2(G101), .A3(n1261), .ZN(n1276) );
NAND2_X1 U934 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
INV_X1 U935 ( .A(n1261), .ZN(n1278) );
NAND2_X1 U936 ( .A1(n1260), .A2(n1075), .ZN(n1261) );
AND4_X1 U937 ( .A1(n1279), .A2(n1081), .A3(n1084), .A4(n1257), .ZN(n1260) );
NAND2_X1 U938 ( .A1(n1280), .A2(n1281), .ZN(n1277) );
OR2_X1 U939 ( .A1(n1193), .A2(KEYINPUT38), .ZN(n1281) );
NAND2_X1 U940 ( .A1(KEYINPUT38), .A2(n1282), .ZN(n1280) );
NAND2_X1 U941 ( .A1(KEYINPUT58), .A2(G101), .ZN(n1282) );
XNOR2_X1 U942 ( .A(G125), .B(n1224), .ZN(G27) );
NAND4_X1 U943 ( .A1(n1075), .A2(n1241), .A3(n1080), .A4(n1283), .ZN(n1224) );
NOR2_X1 U944 ( .A1(n1069), .A2(n1236), .ZN(n1283) );
INV_X1 U945 ( .A(n1284), .ZN(n1069) );
NAND2_X1 U946 ( .A1(n1061), .A2(n1285), .ZN(n1241) );
NAND3_X1 U947 ( .A1(G902), .A2(n1286), .A3(n1118), .ZN(n1285) );
NOR2_X1 U948 ( .A1(n1128), .A2(G900), .ZN(n1118) );
XNOR2_X1 U949 ( .A(G122), .B(n1247), .ZN(G24) );
NAND4_X1 U950 ( .A1(n1268), .A2(n1284), .A3(n1287), .A4(n1248), .ZN(n1247) );
NOR2_X1 U951 ( .A1(n1269), .A2(n1073), .ZN(n1287) );
INV_X1 U952 ( .A(n1249), .ZN(n1073) );
NOR2_X1 U953 ( .A1(n1273), .A2(n1274), .ZN(n1249) );
XOR2_X1 U954 ( .A(n1288), .B(n1258), .Z(G21) );
NOR2_X1 U955 ( .A1(n1255), .A2(n1289), .ZN(n1258) );
NAND4_X1 U956 ( .A1(n1279), .A2(n1284), .A3(n1274), .A4(n1273), .ZN(n1255) );
INV_X1 U957 ( .A(n1290), .ZN(n1274) );
NAND2_X1 U958 ( .A1(KEYINPUT26), .A2(n1291), .ZN(n1288) );
INV_X1 U959 ( .A(G119), .ZN(n1291) );
XNOR2_X1 U960 ( .A(G116), .B(n1246), .ZN(G18) );
NAND2_X1 U961 ( .A1(n1262), .A2(n1088), .ZN(n1246) );
NOR2_X1 U962 ( .A1(n1269), .A2(n1268), .ZN(n1088) );
INV_X1 U963 ( .A(n1292), .ZN(n1262) );
XOR2_X1 U964 ( .A(G113), .B(n1293), .Z(G15) );
NOR3_X1 U965 ( .A1(n1292), .A2(KEYINPUT15), .A3(n1236), .ZN(n1293) );
NAND2_X1 U966 ( .A1(n1269), .A2(n1268), .ZN(n1236) );
NAND3_X1 U967 ( .A1(n1081), .A2(n1248), .A3(n1284), .ZN(n1292) );
NOR2_X1 U968 ( .A1(n1085), .A2(n1094), .ZN(n1284) );
INV_X1 U969 ( .A(n1086), .ZN(n1094) );
AND2_X1 U970 ( .A1(n1273), .A2(n1290), .ZN(n1081) );
XNOR2_X1 U971 ( .A(G110), .B(n1245), .ZN(G12) );
NAND4_X1 U972 ( .A1(n1279), .A2(n1080), .A3(n1084), .A4(n1248), .ZN(n1245) );
INV_X1 U973 ( .A(n1289), .ZN(n1248) );
NAND2_X1 U974 ( .A1(n1075), .A2(n1257), .ZN(n1289) );
NAND2_X1 U975 ( .A1(n1061), .A2(n1294), .ZN(n1257) );
NAND4_X1 U976 ( .A1(G902), .A2(G953), .A3(n1286), .A4(n1147), .ZN(n1294) );
INV_X1 U977 ( .A(G898), .ZN(n1147) );
NAND3_X1 U978 ( .A1(n1286), .A2(n1128), .A3(G952), .ZN(n1061) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1286) );
INV_X1 U980 ( .A(n1235), .ZN(n1075) );
NAND2_X1 U981 ( .A1(n1076), .A2(n1077), .ZN(n1235) );
NAND2_X1 U982 ( .A1(G214), .A2(n1295), .ZN(n1077) );
XNOR2_X1 U983 ( .A(n1296), .B(n1105), .ZN(n1076) );
NAND2_X1 U984 ( .A1(n1297), .A2(n1263), .ZN(n1105) );
XOR2_X1 U985 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U986 ( .A(n1216), .B(n1300), .Z(n1299) );
NOR2_X1 U987 ( .A1(G125), .A2(KEYINPUT33), .ZN(n1300) );
XOR2_X1 U988 ( .A(n1220), .B(n1217), .Z(n1298) );
AND2_X1 U989 ( .A1(n1301), .A2(n1302), .ZN(n1217) );
XOR2_X1 U990 ( .A(KEYINPUT36), .B(G224), .Z(n1301) );
NAND3_X1 U991 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1220) );
XOR2_X1 U992 ( .A(n1306), .B(KEYINPUT31), .Z(n1305) );
NAND2_X1 U993 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U994 ( .A1(n1161), .A2(n1155), .ZN(n1308) );
INV_X1 U995 ( .A(n1149), .ZN(n1161) );
NAND2_X1 U996 ( .A1(n1309), .A2(n1152), .ZN(n1149) );
NAND3_X1 U997 ( .A1(n1152), .A2(n1310), .A3(n1211), .ZN(n1307) );
NAND2_X1 U998 ( .A1(n1154), .A2(n1155), .ZN(n1304) );
INV_X1 U999 ( .A(n1160), .ZN(n1154) );
NAND2_X1 U1000 ( .A1(n1162), .A2(n1310), .ZN(n1160) );
NAND3_X1 U1001 ( .A1(n1309), .A2(n1162), .A3(n1211), .ZN(n1303) );
INV_X1 U1002 ( .A(n1152), .ZN(n1162) );
XNOR2_X1 U1003 ( .A(G122), .B(n1204), .ZN(n1152) );
INV_X1 U1004 ( .A(n1310), .ZN(n1309) );
NAND3_X1 U1005 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1310) );
NAND2_X1 U1006 ( .A1(KEYINPUT12), .A2(n1314), .ZN(n1313) );
NAND3_X1 U1007 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1312) );
INV_X1 U1008 ( .A(KEYINPUT12), .ZN(n1316) );
OR2_X1 U1009 ( .A1(n1317), .A2(n1315), .ZN(n1311) );
NOR2_X1 U1010 ( .A1(KEYINPUT23), .A2(n1314), .ZN(n1315) );
NAND2_X1 U1011 ( .A1(KEYINPUT40), .A2(n1106), .ZN(n1296) );
NAND2_X1 U1012 ( .A1(G210), .A2(n1295), .ZN(n1106) );
NAND2_X1 U1013 ( .A1(n1318), .A2(n1263), .ZN(n1295) );
AND2_X1 U1014 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1319), .ZN(n1086) );
NAND2_X1 U1016 ( .A1(n1320), .A2(n1100), .ZN(n1085) );
NAND3_X1 U1017 ( .A1(n1321), .A2(n1263), .A3(n1322), .ZN(n1100) );
INV_X1 U1018 ( .A(G469), .ZN(n1321) );
XNOR2_X1 U1019 ( .A(KEYINPUT8), .B(n1099), .ZN(n1320) );
NAND2_X1 U1020 ( .A1(G469), .A2(n1323), .ZN(n1099) );
NAND2_X1 U1021 ( .A1(n1322), .A2(n1263), .ZN(n1323) );
XNOR2_X1 U1022 ( .A(n1324), .B(n1325), .ZN(n1322) );
XOR2_X1 U1023 ( .A(n1206), .B(n1326), .Z(n1325) );
NAND2_X1 U1024 ( .A1(KEYINPUT59), .A2(n1327), .ZN(n1326) );
XNOR2_X1 U1025 ( .A(n1204), .B(n1328), .ZN(n1327) );
XOR2_X1 U1026 ( .A(KEYINPUT7), .B(G140), .Z(n1328) );
NAND2_X1 U1027 ( .A1(G227), .A2(n1302), .ZN(n1206) );
NAND2_X1 U1028 ( .A1(n1329), .A2(n1330), .ZN(n1324) );
NAND2_X1 U1029 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1030 ( .A(KEYINPUT37), .B(n1333), .Z(n1329) );
NOR2_X1 U1031 ( .A1(n1332), .A2(n1331), .ZN(n1333) );
XOR2_X1 U1032 ( .A(n1125), .B(n1211), .Z(n1331) );
INV_X1 U1033 ( .A(n1155), .ZN(n1211) );
XOR2_X1 U1034 ( .A(n1334), .B(n1335), .Z(n1155) );
XOR2_X1 U1035 ( .A(G101), .B(n1336), .Z(n1335) );
XOR2_X1 U1036 ( .A(KEYINPUT41), .B(n1216), .Z(n1125) );
INV_X1 U1037 ( .A(n1337), .ZN(n1216) );
XOR2_X1 U1038 ( .A(n1338), .B(KEYINPUT3), .Z(n1332) );
NOR2_X1 U1039 ( .A1(n1290), .A2(n1273), .ZN(n1080) );
XNOR2_X1 U1040 ( .A(n1101), .B(G472), .ZN(n1273) );
NAND2_X1 U1041 ( .A1(n1339), .A2(n1263), .ZN(n1101) );
XOR2_X1 U1042 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1043 ( .A(n1342), .B(n1194), .ZN(n1341) );
XNOR2_X1 U1044 ( .A(n1338), .B(n1337), .ZN(n1194) );
XOR2_X1 U1045 ( .A(G143), .B(n1343), .Z(n1337) );
XOR2_X1 U1046 ( .A(n1123), .B(n1124), .Z(n1338) );
XOR2_X1 U1047 ( .A(G134), .B(G137), .Z(n1124) );
NAND2_X1 U1048 ( .A1(KEYINPUT14), .A2(n1193), .ZN(n1342) );
INV_X1 U1049 ( .A(G101), .ZN(n1193) );
XOR2_X1 U1050 ( .A(n1191), .B(n1344), .Z(n1340) );
NOR2_X1 U1051 ( .A1(KEYINPUT20), .A2(n1345), .ZN(n1344) );
XNOR2_X1 U1052 ( .A(n1195), .B(KEYINPUT43), .ZN(n1345) );
XOR2_X1 U1053 ( .A(n1317), .B(n1314), .Z(n1195) );
XOR2_X1 U1054 ( .A(G116), .B(G119), .Z(n1317) );
NAND3_X1 U1055 ( .A1(n1302), .A2(n1318), .A3(G210), .ZN(n1191) );
NAND2_X1 U1056 ( .A1(n1346), .A2(n1347), .ZN(n1290) );
NAND2_X1 U1057 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
NAND2_X1 U1058 ( .A1(KEYINPUT21), .A2(n1350), .ZN(n1349) );
NAND2_X1 U1059 ( .A1(n1111), .A2(n1351), .ZN(n1350) );
INV_X1 U1060 ( .A(n1352), .ZN(n1111) );
INV_X1 U1061 ( .A(n1110), .ZN(n1348) );
NAND2_X1 U1062 ( .A1(n1353), .A2(n1352), .ZN(n1346) );
NAND2_X1 U1063 ( .A1(G217), .A2(n1319), .ZN(n1352) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1263), .ZN(n1319) );
NAND2_X1 U1065 ( .A1(n1351), .A2(n1354), .ZN(n1353) );
NAND2_X1 U1066 ( .A1(KEYINPUT21), .A2(n1110), .ZN(n1354) );
NAND2_X1 U1067 ( .A1(n1166), .A2(n1263), .ZN(n1110) );
XOR2_X1 U1068 ( .A(n1355), .B(n1356), .Z(n1166) );
XNOR2_X1 U1069 ( .A(n1204), .B(n1357), .ZN(n1356) );
XOR2_X1 U1070 ( .A(G119), .B(n1358), .Z(n1357) );
NOR2_X1 U1071 ( .A1(KEYINPUT2), .A2(n1359), .ZN(n1358) );
NOR2_X1 U1072 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
XOR2_X1 U1073 ( .A(n1362), .B(KEYINPUT56), .Z(n1361) );
NAND2_X1 U1074 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND3_X1 U1075 ( .A1(G234), .A2(n1302), .A3(n1365), .ZN(n1364) );
INV_X1 U1076 ( .A(G137), .ZN(n1363) );
AND4_X1 U1077 ( .A1(n1302), .A2(G234), .A3(G137), .A4(n1365), .ZN(n1360) );
XNOR2_X1 U1078 ( .A(G221), .B(KEYINPUT17), .ZN(n1365) );
XNOR2_X1 U1079 ( .A(G110), .B(KEYINPUT27), .ZN(n1204) );
XNOR2_X1 U1080 ( .A(n1343), .B(n1126), .ZN(n1355) );
XOR2_X1 U1081 ( .A(G128), .B(G146), .Z(n1343) );
INV_X1 U1082 ( .A(KEYINPUT34), .ZN(n1351) );
INV_X1 U1083 ( .A(n1065), .ZN(n1279) );
NAND2_X1 U1084 ( .A1(n1269), .A2(n1366), .ZN(n1065) );
INV_X1 U1085 ( .A(n1268), .ZN(n1366) );
XNOR2_X1 U1086 ( .A(n1108), .B(n1367), .ZN(n1268) );
NOR2_X1 U1087 ( .A1(G475), .A2(KEYINPUT25), .ZN(n1367) );
NOR2_X1 U1088 ( .A1(n1177), .A2(G902), .ZN(n1108) );
XNOR2_X1 U1089 ( .A(n1368), .B(n1369), .ZN(n1177) );
NOR2_X1 U1090 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1091 ( .A(n1372), .B(KEYINPUT18), .Z(n1371) );
NAND3_X1 U1092 ( .A1(n1373), .A2(n1374), .A3(n1375), .ZN(n1372) );
NOR2_X1 U1093 ( .A1(n1376), .A2(n1373), .ZN(n1370) );
XNOR2_X1 U1094 ( .A(n1377), .B(n1378), .ZN(n1373) );
NOR2_X1 U1095 ( .A1(KEYINPUT63), .A2(n1123), .ZN(n1378) );
INV_X1 U1096 ( .A(G131), .ZN(n1123) );
XNOR2_X1 U1097 ( .A(G143), .B(n1379), .ZN(n1377) );
AND4_X1 U1098 ( .A1(n1380), .A2(n1318), .A3(n1302), .A4(G214), .ZN(n1379) );
INV_X1 U1099 ( .A(G237), .ZN(n1318) );
INV_X1 U1100 ( .A(KEYINPUT46), .ZN(n1380) );
AND2_X1 U1101 ( .A1(n1374), .A2(n1375), .ZN(n1376) );
XOR2_X1 U1102 ( .A(n1381), .B(KEYINPUT22), .Z(n1375) );
OR2_X1 U1103 ( .A1(n1126), .A2(G146), .ZN(n1381) );
NAND2_X1 U1104 ( .A1(n1382), .A2(n1126), .ZN(n1374) );
XOR2_X1 U1105 ( .A(G125), .B(G140), .Z(n1126) );
XOR2_X1 U1106 ( .A(n1383), .B(G146), .Z(n1382) );
XNOR2_X1 U1107 ( .A(KEYINPUT48), .B(KEYINPUT19), .ZN(n1383) );
NAND2_X1 U1108 ( .A1(n1384), .A2(KEYINPUT13), .ZN(n1368) );
XOR2_X1 U1109 ( .A(n1385), .B(n1386), .Z(n1384) );
XOR2_X1 U1110 ( .A(n1314), .B(n1387), .Z(n1386) );
INV_X1 U1111 ( .A(n1334), .ZN(n1387) );
XNOR2_X1 U1112 ( .A(G104), .B(KEYINPUT53), .ZN(n1334) );
XOR2_X1 U1113 ( .A(G113), .B(KEYINPUT11), .Z(n1314) );
XNOR2_X1 U1114 ( .A(G122), .B(KEYINPUT24), .ZN(n1385) );
XOR2_X1 U1115 ( .A(n1109), .B(n1388), .Z(n1269) );
NOR2_X1 U1116 ( .A1(KEYINPUT28), .A2(n1172), .ZN(n1388) );
INV_X1 U1117 ( .A(G478), .ZN(n1172) );
NAND2_X1 U1118 ( .A1(n1170), .A2(n1263), .ZN(n1109) );
INV_X1 U1119 ( .A(G902), .ZN(n1263) );
XNOR2_X1 U1120 ( .A(n1389), .B(n1390), .ZN(n1170) );
XOR2_X1 U1121 ( .A(n1391), .B(n1392), .Z(n1390) );
XOR2_X1 U1122 ( .A(G128), .B(G122), .Z(n1392) );
XOR2_X1 U1123 ( .A(G143), .B(G134), .Z(n1391) );
XOR2_X1 U1124 ( .A(n1393), .B(n1336), .Z(n1389) );
XOR2_X1 U1125 ( .A(G107), .B(KEYINPUT30), .Z(n1336) );
XOR2_X1 U1126 ( .A(n1394), .B(G116), .Z(n1393) );
NAND4_X1 U1127 ( .A1(KEYINPUT44), .A2(G234), .A3(G217), .A4(n1302), .ZN(n1394) );
XNOR2_X1 U1128 ( .A(n1128), .B(KEYINPUT1), .ZN(n1302) );
INV_X1 U1129 ( .A(G953), .ZN(n1128) );
endmodule


