//Key = 0000000111000010010110110011101011100011111000010011000111010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;

XOR2_X1 U736 ( .A(G107), .B(n1015), .Z(G9) );
NOR2_X1 U737 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NOR2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
NOR2_X1 U740 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U743 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U744 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U745 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U747 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
XNOR2_X1 U748 ( .A(n1040), .B(KEYINPUT50), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1028) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1035), .ZN(n1044) );
NOR2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
AND2_X1 U753 ( .A1(n1048), .A2(KEYINPUT33), .ZN(n1046) );
NOR3_X1 U754 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1043) );
XNOR2_X1 U755 ( .A(KEYINPUT14), .B(n1031), .ZN(n1049) );
NOR3_X1 U756 ( .A1(n1042), .A2(n1052), .A3(n1035), .ZN(n1024) );
NOR3_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
AND2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR3_X1 U759 ( .A1(n1058), .A2(KEYINPUT33), .A3(n1059), .ZN(n1054) );
NOR2_X1 U760 ( .A1(n1031), .A2(n1060), .ZN(n1053) );
NOR3_X1 U761 ( .A1(n1020), .A2(G952), .A3(n1018), .ZN(n1016) );
AND4_X1 U762 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1018) );
NOR4_X1 U763 ( .A1(n1065), .A2(n1066), .A3(n1035), .A4(n1042), .ZN(n1064) );
NOR2_X1 U764 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XNOR2_X1 U765 ( .A(n1069), .B(KEYINPUT23), .ZN(n1068) );
AND2_X1 U766 ( .A1(n1067), .A2(n1069), .ZN(n1065) );
XNOR2_X1 U767 ( .A(G472), .B(n1070), .ZN(n1061) );
NAND2_X1 U768 ( .A1(KEYINPUT55), .A2(n1071), .ZN(n1070) );
INV_X1 U769 ( .A(n1072), .ZN(n1020) );
NAND3_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(G72) );
XOR2_X1 U771 ( .A(n1076), .B(KEYINPUT58), .Z(n1075) );
NAND3_X1 U772 ( .A1(n1077), .A2(n1078), .A3(G953), .ZN(n1076) );
NAND2_X1 U773 ( .A1(G900), .A2(G227), .ZN(n1077) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
XOR2_X1 U775 ( .A(n1078), .B(n1081), .Z(n1079) );
OR3_X1 U776 ( .A1(n1078), .A2(n1082), .A3(n1080), .ZN(n1073) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1084), .ZN(n1078) );
NAND2_X1 U778 ( .A1(G953), .A2(n1085), .ZN(n1084) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(n1083) );
XNOR2_X1 U780 ( .A(n1088), .B(n1089), .ZN(n1087) );
NOR2_X1 U781 ( .A1(KEYINPUT43), .A2(n1090), .ZN(n1089) );
XNOR2_X1 U782 ( .A(n1091), .B(G125), .ZN(n1090) );
XOR2_X1 U783 ( .A(n1092), .B(n1093), .Z(n1086) );
NAND3_X1 U784 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1092) );
NAND2_X1 U785 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U786 ( .A1(KEYINPUT6), .A2(n1099), .ZN(n1095) );
NAND2_X1 U787 ( .A1(G134), .A2(n1100), .ZN(n1099) );
XNOR2_X1 U788 ( .A(KEYINPUT21), .B(n1097), .ZN(n1100) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1094) );
INV_X1 U790 ( .A(KEYINPUT6), .ZN(n1102) );
NAND2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
OR3_X1 U792 ( .A1(n1098), .A2(n1097), .A3(KEYINPUT21), .ZN(n1104) );
NAND2_X1 U793 ( .A1(KEYINPUT21), .A2(n1097), .ZN(n1103) );
XNOR2_X1 U794 ( .A(G137), .B(KEYINPUT9), .ZN(n1097) );
XOR2_X1 U795 ( .A(n1105), .B(n1106), .Z(G69) );
XOR2_X1 U796 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U797 ( .A1(G953), .A2(n1109), .ZN(n1108) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
XOR2_X1 U799 ( .A(KEYINPUT56), .B(n1112), .Z(n1111) );
NOR2_X1 U800 ( .A1(G898), .A2(n1080), .ZN(n1112) );
NAND2_X1 U801 ( .A1(G953), .A2(n1113), .ZN(n1105) );
NAND2_X1 U802 ( .A1(G898), .A2(G224), .ZN(n1113) );
NOR2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(G66) );
NOR3_X1 U804 ( .A1(n1069), .A2(n1116), .A3(n1117), .ZN(n1115) );
NOR4_X1 U805 ( .A1(n1118), .A2(n1119), .A3(KEYINPUT0), .A4(n1067), .ZN(n1117) );
INV_X1 U806 ( .A(n1120), .ZN(n1118) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1120), .ZN(n1116) );
NOR3_X1 U808 ( .A1(n1067), .A2(KEYINPUT0), .A3(n1122), .ZN(n1121) );
NOR2_X1 U809 ( .A1(n1114), .A2(n1123), .ZN(G63) );
XOR2_X1 U810 ( .A(n1124), .B(n1125), .Z(n1123) );
AND2_X1 U811 ( .A1(G478), .A2(n1126), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1114), .A2(n1127), .ZN(G60) );
XOR2_X1 U813 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR3_X1 U814 ( .A1(n1119), .A2(n1130), .A3(n1131), .ZN(n1128) );
XNOR2_X1 U815 ( .A(KEYINPUT63), .B(KEYINPUT52), .ZN(n1130) );
INV_X1 U816 ( .A(n1126), .ZN(n1119) );
XOR2_X1 U817 ( .A(n1132), .B(n1133), .Z(G6) );
NOR2_X1 U818 ( .A1(KEYINPUT44), .A2(n1134), .ZN(n1133) );
NOR2_X1 U819 ( .A1(n1114), .A2(n1135), .ZN(G57) );
XNOR2_X1 U820 ( .A(n1136), .B(n1137), .ZN(n1135) );
NAND3_X1 U821 ( .A1(n1138), .A2(n1139), .A3(KEYINPUT19), .ZN(n1136) );
NAND4_X1 U822 ( .A1(n1140), .A2(G472), .A3(n1126), .A4(n1141), .ZN(n1139) );
INV_X1 U823 ( .A(KEYINPUT40), .ZN(n1141) );
NAND2_X1 U824 ( .A1(n1142), .A2(KEYINPUT40), .ZN(n1138) );
XOR2_X1 U825 ( .A(n1140), .B(n1143), .Z(n1142) );
AND2_X1 U826 ( .A1(G472), .A2(n1126), .ZN(n1143) );
XOR2_X1 U827 ( .A(n1144), .B(n1145), .Z(n1140) );
XOR2_X1 U828 ( .A(n1146), .B(KEYINPUT16), .Z(n1144) );
NOR2_X1 U829 ( .A1(n1114), .A2(n1147), .ZN(G54) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U831 ( .A(n1150), .B(n1151), .Z(n1149) );
AND2_X1 U832 ( .A1(G469), .A2(n1126), .ZN(n1150) );
XOR2_X1 U833 ( .A(n1152), .B(n1153), .Z(n1148) );
NOR2_X1 U834 ( .A1(KEYINPUT60), .A2(n1154), .ZN(n1153) );
NAND2_X1 U835 ( .A1(KEYINPUT42), .A2(n1155), .ZN(n1152) );
XOR2_X1 U836 ( .A(KEYINPUT47), .B(n1156), .Z(n1155) );
NOR2_X1 U837 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XNOR2_X1 U838 ( .A(KEYINPUT18), .B(n1159), .ZN(n1158) );
NOR2_X1 U839 ( .A1(n1114), .A2(n1160), .ZN(G51) );
XOR2_X1 U840 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U841 ( .A(n1163), .B(n1110), .ZN(n1162) );
AND2_X1 U842 ( .A1(G210), .A2(n1126), .ZN(n1163) );
NOR2_X1 U843 ( .A1(n1164), .A2(n1122), .ZN(n1126) );
INV_X1 U844 ( .A(n1021), .ZN(n1122) );
NAND2_X1 U845 ( .A1(n1081), .A2(n1109), .ZN(n1021) );
AND4_X1 U846 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1109) );
NOR4_X1 U847 ( .A1(n1169), .A2(n1170), .A3(n1132), .A4(n1171), .ZN(n1168) );
NOR3_X1 U848 ( .A1(n1060), .A2(n1172), .A3(n1031), .ZN(n1171) );
NOR3_X1 U849 ( .A1(n1172), .A2(n1027), .A3(n1058), .ZN(n1132) );
NOR2_X1 U850 ( .A1(n1015), .A2(n1173), .ZN(n1167) );
NOR3_X1 U851 ( .A1(n1174), .A2(n1027), .A3(n1172), .ZN(n1015) );
INV_X1 U852 ( .A(n1175), .ZN(n1172) );
AND4_X1 U853 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1081) );
NOR4_X1 U854 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
NOR4_X1 U855 ( .A1(n1184), .A2(n1185), .A3(n1174), .A4(n1060), .ZN(n1183) );
NOR2_X1 U856 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
INV_X1 U857 ( .A(KEYINPUT29), .ZN(n1187) );
NOR2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
NOR2_X1 U859 ( .A1(KEYINPUT29), .A2(n1190), .ZN(n1184) );
NOR3_X1 U860 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1178) );
NOR3_X1 U861 ( .A1(n1194), .A2(n1195), .A3(n1035), .ZN(n1193) );
NOR3_X1 U862 ( .A1(n1058), .A2(n1196), .A3(n1189), .ZN(n1195) );
INV_X1 U863 ( .A(KEYINPUT48), .ZN(n1194) );
NOR4_X1 U864 ( .A1(KEYINPUT48), .A2(n1058), .A3(n1196), .A4(n1197), .ZN(n1192) );
XNOR2_X1 U865 ( .A(n1198), .B(KEYINPUT3), .ZN(n1196) );
XOR2_X1 U866 ( .A(n1199), .B(n1200), .Z(n1161) );
XNOR2_X1 U867 ( .A(KEYINPUT24), .B(n1201), .ZN(n1199) );
NOR2_X1 U868 ( .A1(KEYINPUT37), .A2(n1202), .ZN(n1201) );
XOR2_X1 U869 ( .A(n1203), .B(G125), .Z(n1202) );
NAND2_X1 U870 ( .A1(KEYINPUT51), .A2(n1204), .ZN(n1203) );
NOR2_X1 U871 ( .A1(n1080), .A2(G952), .ZN(n1114) );
XOR2_X1 U872 ( .A(n1205), .B(n1191), .Z(G48) );
AND2_X1 U873 ( .A1(n1206), .A2(n1048), .ZN(n1191) );
NAND2_X1 U874 ( .A1(KEYINPUT22), .A2(n1207), .ZN(n1205) );
XNOR2_X1 U875 ( .A(G143), .B(n1208), .ZN(G45) );
NAND2_X1 U876 ( .A1(KEYINPUT41), .A2(n1182), .ZN(n1208) );
NOR4_X1 U877 ( .A1(n1209), .A2(n1060), .A3(n1210), .A4(n1211), .ZN(n1182) );
OR2_X1 U878 ( .A1(n1212), .A2(n1063), .ZN(n1210) );
XNOR2_X1 U879 ( .A(n1091), .B(n1181), .ZN(G42) );
NOR4_X1 U880 ( .A1(n1058), .A2(n1197), .A3(n1213), .A4(n1214), .ZN(n1181) );
INV_X1 U881 ( .A(n1048), .ZN(n1058) );
XOR2_X1 U882 ( .A(G137), .B(n1180), .Z(G39) );
AND3_X1 U883 ( .A1(n1057), .A2(n1213), .A3(n1190), .ZN(n1180) );
XNOR2_X1 U884 ( .A(G134), .B(n1215), .ZN(G36) );
NAND2_X1 U885 ( .A1(n1216), .A2(n1047), .ZN(n1215) );
XNOR2_X1 U886 ( .A(G131), .B(n1217), .ZN(G33) );
NAND2_X1 U887 ( .A1(n1216), .A2(n1048), .ZN(n1217) );
NOR2_X1 U888 ( .A1(n1060), .A2(n1197), .ZN(n1216) );
INV_X1 U889 ( .A(n1190), .ZN(n1197) );
NOR2_X1 U890 ( .A1(n1189), .A2(n1035), .ZN(n1190) );
INV_X1 U891 ( .A(n1188), .ZN(n1035) );
NOR2_X1 U892 ( .A1(n1051), .A2(n1218), .ZN(n1188) );
NAND2_X1 U893 ( .A1(n1037), .A2(n1219), .ZN(n1189) );
XNOR2_X1 U894 ( .A(G128), .B(n1176), .ZN(G30) );
NAND2_X1 U895 ( .A1(n1206), .A2(n1047), .ZN(n1176) );
NOR4_X1 U896 ( .A1(n1211), .A2(n1056), .A3(n1214), .A4(n1212), .ZN(n1206) );
XNOR2_X1 U897 ( .A(G101), .B(n1220), .ZN(G3) );
NAND4_X1 U898 ( .A1(n1221), .A2(KEYINPUT39), .A3(n1222), .A4(n1198), .ZN(n1220) );
NOR2_X1 U899 ( .A1(n1211), .A2(n1031), .ZN(n1222) );
XNOR2_X1 U900 ( .A(n1223), .B(KEYINPUT46), .ZN(n1221) );
XOR2_X1 U901 ( .A(n1177), .B(n1224), .Z(G27) );
XNOR2_X1 U902 ( .A(G125), .B(KEYINPUT2), .ZN(n1224) );
NAND3_X1 U903 ( .A1(n1033), .A2(n1048), .A3(n1225), .ZN(n1177) );
NOR3_X1 U904 ( .A1(n1213), .A2(n1212), .A3(n1214), .ZN(n1225) );
INV_X1 U905 ( .A(n1219), .ZN(n1212) );
NAND2_X1 U906 ( .A1(n1226), .A2(n1023), .ZN(n1219) );
NAND2_X1 U907 ( .A1(n1227), .A2(n1085), .ZN(n1226) );
INV_X1 U908 ( .A(G900), .ZN(n1085) );
XOR2_X1 U909 ( .A(G122), .B(n1170), .Z(G24) );
AND3_X1 U910 ( .A1(n1033), .A2(n1059), .A3(n1228), .ZN(n1170) );
NOR3_X1 U911 ( .A1(n1209), .A2(n1223), .A3(n1063), .ZN(n1228) );
INV_X1 U912 ( .A(n1027), .ZN(n1059) );
NAND2_X1 U913 ( .A1(n1214), .A2(n1056), .ZN(n1027) );
XNOR2_X1 U914 ( .A(G119), .B(n1165), .ZN(G21) );
NAND4_X1 U915 ( .A1(n1033), .A2(n1057), .A3(n1213), .A4(n1229), .ZN(n1165) );
XOR2_X1 U916 ( .A(G116), .B(n1169), .Z(G18) );
AND2_X1 U917 ( .A1(n1230), .A2(n1047), .ZN(n1169) );
INV_X1 U918 ( .A(n1174), .ZN(n1047) );
NAND2_X1 U919 ( .A1(n1231), .A2(n1063), .ZN(n1174) );
XOR2_X1 U920 ( .A(G113), .B(n1173), .Z(G15) );
AND2_X1 U921 ( .A1(n1230), .A2(n1048), .ZN(n1173) );
NOR2_X1 U922 ( .A1(n1063), .A2(n1231), .ZN(n1048) );
INV_X1 U923 ( .A(n1209), .ZN(n1231) );
AND3_X1 U924 ( .A1(n1198), .A2(n1229), .A3(n1033), .ZN(n1230) );
NOR3_X1 U925 ( .A1(n1232), .A2(n1218), .A3(n1042), .ZN(n1033) );
NAND2_X1 U926 ( .A1(n1233), .A2(n1039), .ZN(n1042) );
INV_X1 U927 ( .A(n1040), .ZN(n1233) );
INV_X1 U928 ( .A(n1050), .ZN(n1218) );
INV_X1 U929 ( .A(n1051), .ZN(n1232) );
INV_X1 U930 ( .A(n1060), .ZN(n1198) );
NAND2_X1 U931 ( .A1(n1214), .A2(n1213), .ZN(n1060) );
XNOR2_X1 U932 ( .A(G110), .B(n1166), .ZN(G12) );
NAND3_X1 U933 ( .A1(n1056), .A2(n1175), .A3(n1057), .ZN(n1166) );
NOR2_X1 U934 ( .A1(n1031), .A2(n1214), .ZN(n1057) );
XOR2_X1 U935 ( .A(n1069), .B(n1067), .Z(n1214) );
NAND2_X1 U936 ( .A1(G217), .A2(n1234), .ZN(n1067) );
NOR2_X1 U937 ( .A1(n1120), .A2(G902), .ZN(n1069) );
XNOR2_X1 U938 ( .A(n1235), .B(n1236), .ZN(n1120) );
XOR2_X1 U939 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U940 ( .A(G128), .B(G125), .Z(n1238) );
XNOR2_X1 U941 ( .A(n1207), .B(G137), .ZN(n1237) );
XOR2_X1 U942 ( .A(n1239), .B(n1240), .Z(n1235) );
XNOR2_X1 U943 ( .A(n1241), .B(n1242), .ZN(n1240) );
NOR2_X1 U944 ( .A1(KEYINPUT12), .A2(n1091), .ZN(n1242) );
NAND2_X1 U945 ( .A1(n1243), .A2(KEYINPUT38), .ZN(n1241) );
XNOR2_X1 U946 ( .A(G119), .B(KEYINPUT1), .ZN(n1243) );
XOR2_X1 U947 ( .A(n1244), .B(G110), .Z(n1239) );
NAND2_X1 U948 ( .A1(n1245), .A2(G221), .ZN(n1244) );
NAND2_X1 U949 ( .A1(n1063), .A2(n1209), .ZN(n1031) );
XOR2_X1 U950 ( .A(n1062), .B(KEYINPUT45), .Z(n1209) );
XNOR2_X1 U951 ( .A(n1246), .B(n1247), .ZN(n1062) );
XOR2_X1 U952 ( .A(KEYINPUT26), .B(G478), .Z(n1247) );
OR2_X1 U953 ( .A1(n1125), .A2(G902), .ZN(n1246) );
XNOR2_X1 U954 ( .A(n1248), .B(n1249), .ZN(n1125) );
XOR2_X1 U955 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U956 ( .A(G122), .B(G116), .Z(n1251) );
XNOR2_X1 U957 ( .A(KEYINPUT10), .B(n1098), .ZN(n1250) );
XOR2_X1 U958 ( .A(n1252), .B(n1253), .Z(n1248) );
XNOR2_X1 U959 ( .A(n1254), .B(n1255), .ZN(n1253) );
NOR2_X1 U960 ( .A1(KEYINPUT13), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U961 ( .A(n1257), .B(n1258), .ZN(n1256) );
NOR2_X1 U962 ( .A1(G128), .A2(KEYINPUT11), .ZN(n1258) );
NAND2_X1 U963 ( .A1(n1259), .A2(KEYINPUT61), .ZN(n1254) );
XNOR2_X1 U964 ( .A(G107), .B(KEYINPUT62), .ZN(n1259) );
NAND2_X1 U965 ( .A1(G217), .A2(n1245), .ZN(n1252) );
AND2_X1 U966 ( .A1(G234), .A2(n1080), .ZN(n1245) );
XNOR2_X1 U967 ( .A(n1260), .B(n1131), .ZN(n1063) );
INV_X1 U968 ( .A(G475), .ZN(n1131) );
OR2_X1 U969 ( .A1(n1129), .A2(G902), .ZN(n1260) );
XNOR2_X1 U970 ( .A(n1261), .B(n1262), .ZN(n1129) );
XOR2_X1 U971 ( .A(KEYINPUT20), .B(G113), .Z(n1262) );
XOR2_X1 U972 ( .A(n1263), .B(n1264), .Z(n1261) );
NAND3_X1 U973 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1263) );
NAND2_X1 U974 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U975 ( .A1(KEYINPUT25), .A2(n1270), .ZN(n1266) );
NAND2_X1 U976 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
INV_X1 U977 ( .A(n1269), .ZN(n1272) );
XNOR2_X1 U978 ( .A(KEYINPUT53), .B(n1268), .ZN(n1271) );
NAND2_X1 U979 ( .A1(n1273), .A2(n1274), .ZN(n1265) );
INV_X1 U980 ( .A(KEYINPUT25), .ZN(n1274) );
NAND2_X1 U981 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
OR3_X1 U982 ( .A1(n1268), .A2(n1269), .A3(KEYINPUT53), .ZN(n1276) );
XNOR2_X1 U983 ( .A(n1277), .B(n1278), .ZN(n1269) );
XNOR2_X1 U984 ( .A(G131), .B(n1279), .ZN(n1278) );
NAND2_X1 U985 ( .A1(n1280), .A2(G214), .ZN(n1279) );
NAND2_X1 U986 ( .A1(KEYINPUT17), .A2(n1257), .ZN(n1277) );
NAND2_X1 U987 ( .A1(KEYINPUT53), .A2(n1268), .ZN(n1275) );
XNOR2_X1 U988 ( .A(n1281), .B(n1282), .ZN(n1268) );
NOR2_X1 U989 ( .A1(KEYINPUT36), .A2(G125), .ZN(n1282) );
XNOR2_X1 U990 ( .A(G140), .B(G146), .ZN(n1281) );
NOR2_X1 U991 ( .A1(n1211), .A2(n1223), .ZN(n1175) );
INV_X1 U992 ( .A(n1229), .ZN(n1223) );
NAND2_X1 U993 ( .A1(n1023), .A2(n1283), .ZN(n1229) );
NAND2_X1 U994 ( .A1(n1227), .A2(n1284), .ZN(n1283) );
INV_X1 U995 ( .A(G898), .ZN(n1284) );
AND3_X1 U996 ( .A1(G953), .A2(n1285), .A3(n1286), .ZN(n1227) );
XNOR2_X1 U997 ( .A(G902), .B(KEYINPUT32), .ZN(n1286) );
NAND3_X1 U998 ( .A1(n1072), .A2(n1285), .A3(G952), .ZN(n1023) );
NAND2_X1 U999 ( .A1(G237), .A2(G234), .ZN(n1285) );
XOR2_X1 U1000 ( .A(G953), .B(KEYINPUT7), .Z(n1072) );
NAND3_X1 U1001 ( .A1(n1051), .A2(n1050), .A3(n1037), .ZN(n1211) );
AND2_X1 U1002 ( .A1(n1040), .A2(n1039), .ZN(n1037) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1234), .ZN(n1039) );
NAND2_X1 U1004 ( .A1(G234), .A2(n1164), .ZN(n1234) );
XOR2_X1 U1005 ( .A(G469), .B(n1287), .Z(n1040) );
NOR2_X1 U1006 ( .A1(n1288), .A2(G902), .ZN(n1287) );
NOR2_X1 U1007 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XOR2_X1 U1008 ( .A(n1291), .B(KEYINPUT30), .Z(n1290) );
NAND2_X1 U1009 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NOR2_X1 U1010 ( .A1(n1293), .A2(n1292), .ZN(n1289) );
XNOR2_X1 U1011 ( .A(n1154), .B(n1151), .ZN(n1292) );
XNOR2_X1 U1012 ( .A(n1294), .B(n1295), .ZN(n1154) );
XOR2_X1 U1013 ( .A(KEYINPUT31), .B(n1296), .Z(n1295) );
NOR2_X1 U1014 ( .A1(KEYINPUT5), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U1015 ( .A(G104), .B(KEYINPUT8), .ZN(n1297) );
XNOR2_X1 U1016 ( .A(n1093), .B(n1298), .ZN(n1294) );
XOR2_X1 U1017 ( .A(G146), .B(n1299), .Z(n1093) );
AND2_X1 U1018 ( .A1(n1300), .A2(n1159), .ZN(n1293) );
NAND2_X1 U1019 ( .A1(n1301), .A2(n1302), .ZN(n1159) );
NAND2_X1 U1020 ( .A1(G227), .A2(n1080), .ZN(n1302) );
XOR2_X1 U1021 ( .A(KEYINPUT34), .B(n1157), .Z(n1300) );
NOR3_X1 U1022 ( .A1(n1082), .A2(G953), .A3(n1301), .ZN(n1157) );
XNOR2_X1 U1023 ( .A(G110), .B(n1091), .ZN(n1301) );
INV_X1 U1024 ( .A(G140), .ZN(n1091) );
INV_X1 U1025 ( .A(G227), .ZN(n1082) );
NAND2_X1 U1026 ( .A1(G214), .A2(n1303), .ZN(n1050) );
INV_X1 U1027 ( .A(n1304), .ZN(n1303) );
XNOR2_X1 U1028 ( .A(n1305), .B(n1306), .ZN(n1051) );
NOR2_X1 U1029 ( .A1(n1304), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U1030 ( .A(G210), .B(KEYINPUT15), .ZN(n1307) );
NOR2_X1 U1031 ( .A1(G902), .A2(G237), .ZN(n1304) );
NAND2_X1 U1032 ( .A1(n1308), .A2(n1164), .ZN(n1305) );
XOR2_X1 U1033 ( .A(n1309), .B(n1310), .Z(n1308) );
XOR2_X1 U1034 ( .A(n1200), .B(n1311), .Z(n1310) );
XOR2_X1 U1035 ( .A(KEYINPUT27), .B(G125), .Z(n1311) );
AND2_X1 U1036 ( .A1(G224), .A2(n1080), .ZN(n1200) );
INV_X1 U1037 ( .A(G953), .ZN(n1080) );
XOR2_X1 U1038 ( .A(n1110), .B(n1204), .Z(n1309) );
XOR2_X1 U1039 ( .A(n1312), .B(n1313), .Z(n1110) );
XOR2_X1 U1040 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1041 ( .A(KEYINPUT8), .B(G110), .Z(n1315) );
NOR2_X1 U1042 ( .A1(KEYINPUT49), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U1043 ( .A(KEYINPUT59), .B(G116), .ZN(n1316) );
XNOR2_X1 U1044 ( .A(n1298), .B(n1317), .ZN(n1312) );
XOR2_X1 U1045 ( .A(n1318), .B(n1264), .Z(n1317) );
XNOR2_X1 U1046 ( .A(n1134), .B(G122), .ZN(n1264) );
INV_X1 U1047 ( .A(G104), .ZN(n1134) );
XOR2_X1 U1048 ( .A(G101), .B(G107), .Z(n1298) );
INV_X1 U1049 ( .A(n1213), .ZN(n1056) );
XOR2_X1 U1050 ( .A(G472), .B(n1319), .Z(n1213) );
NOR2_X1 U1051 ( .A1(KEYINPUT35), .A2(n1071), .ZN(n1319) );
NAND3_X1 U1052 ( .A1(n1320), .A2(n1321), .A3(n1164), .ZN(n1071) );
INV_X1 U1053 ( .A(G902), .ZN(n1164) );
NAND2_X1 U1054 ( .A1(KEYINPUT57), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U1055 ( .A(n1323), .B(n1324), .ZN(n1322) );
INV_X1 U1056 ( .A(n1137), .ZN(n1324) );
NAND3_X1 U1057 ( .A1(n1137), .A2(n1323), .A3(n1325), .ZN(n1320) );
INV_X1 U1058 ( .A(KEYINPUT57), .ZN(n1325) );
XOR2_X1 U1059 ( .A(n1146), .B(n1326), .Z(n1323) );
NOR2_X1 U1060 ( .A1(KEYINPUT54), .A2(n1145), .ZN(n1326) );
XOR2_X1 U1061 ( .A(n1204), .B(n1151), .Z(n1145) );
XNOR2_X1 U1062 ( .A(n1088), .B(n1327), .ZN(n1151) );
XNOR2_X1 U1063 ( .A(G137), .B(n1098), .ZN(n1327) );
INV_X1 U1064 ( .A(G134), .ZN(n1098) );
INV_X1 U1065 ( .A(G131), .ZN(n1088) );
AND2_X1 U1066 ( .A1(n1328), .A2(n1329), .ZN(n1204) );
NAND2_X1 U1067 ( .A1(n1299), .A2(G146), .ZN(n1329) );
NAND2_X1 U1068 ( .A1(n1330), .A2(n1207), .ZN(n1328) );
INV_X1 U1069 ( .A(G146), .ZN(n1207) );
XNOR2_X1 U1070 ( .A(n1299), .B(KEYINPUT4), .ZN(n1330) );
XNOR2_X1 U1071 ( .A(G128), .B(n1257), .ZN(n1299) );
INV_X1 U1072 ( .A(G143), .ZN(n1257) );
XOR2_X1 U1073 ( .A(n1331), .B(n1318), .Z(n1146) );
XOR2_X1 U1074 ( .A(G113), .B(G119), .Z(n1318) );
NAND2_X1 U1075 ( .A1(KEYINPUT28), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1076 ( .A(KEYINPUT59), .B(G116), .Z(n1332) );
XNOR2_X1 U1077 ( .A(n1333), .B(G101), .ZN(n1137) );
NAND2_X1 U1078 ( .A1(n1280), .A2(G210), .ZN(n1333) );
NOR2_X1 U1079 ( .A1(G953), .A2(G237), .ZN(n1280) );
endmodule


