//Key = 1111100100011111011100111101100111000000100000101000111010110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384;

XNOR2_X1 U762 ( .A(G107), .B(n1063), .ZN(G9) );
NOR2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(G75) );
NOR4_X1 U764 ( .A1(G953), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1065) );
NOR2_X1 U765 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR3_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR4_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1078) );
AND2_X1 U771 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
AND3_X1 U773 ( .A1(n1087), .A2(n1086), .A3(n1088), .ZN(n1080) );
NOR2_X1 U774 ( .A1(n1089), .A2(n1090), .ZN(n1076) );
NOR2_X1 U775 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NOR3_X1 U776 ( .A1(n1093), .A2(n1094), .A3(n1085), .ZN(n1091) );
XOR2_X1 U777 ( .A(KEYINPUT29), .B(KEYINPUT21), .Z(n1085) );
NOR3_X1 U778 ( .A1(n1079), .A2(n1095), .A3(n1090), .ZN(n1071) );
INV_X1 U779 ( .A(n1084), .ZN(n1090) );
NOR3_X1 U780 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
NOR2_X1 U781 ( .A1(n1099), .A2(n1075), .ZN(n1098) );
NOR2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U783 ( .A1(n1073), .A2(n1102), .ZN(n1096) );
NOR3_X1 U784 ( .A1(n1066), .A2(G953), .A3(G952), .ZN(n1064) );
AND2_X1 U785 ( .A1(n1103), .A2(n1104), .ZN(n1066) );
NOR4_X1 U786 ( .A1(n1105), .A2(n1106), .A3(n1088), .A4(n1107), .ZN(n1104) );
XOR2_X1 U787 ( .A(n1108), .B(G475), .Z(n1107) );
NAND2_X1 U788 ( .A1(KEYINPUT46), .A2(n1109), .ZN(n1108) );
NOR2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1106) );
XNOR2_X1 U790 ( .A(n1112), .B(n1113), .ZN(n1111) );
XNOR2_X1 U791 ( .A(KEYINPUT49), .B(KEYINPUT23), .ZN(n1113) );
NOR2_X1 U792 ( .A1(G902), .A2(n1114), .ZN(n1110) );
NOR4_X1 U793 ( .A1(n1115), .A2(n1116), .A3(n1079), .A4(n1117), .ZN(n1103) );
XOR2_X1 U794 ( .A(G472), .B(n1118), .Z(n1117) );
XNOR2_X1 U795 ( .A(n1119), .B(n1120), .ZN(n1115) );
NAND2_X1 U796 ( .A1(KEYINPUT61), .A2(n1121), .ZN(n1119) );
INV_X1 U797 ( .A(G469), .ZN(n1121) );
XOR2_X1 U798 ( .A(n1122), .B(n1123), .Z(G72) );
XOR2_X1 U799 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
AND2_X1 U801 ( .A1(G227), .A2(G900), .ZN(n1126) );
NAND2_X1 U802 ( .A1(n1128), .A2(n1129), .ZN(n1124) );
NAND2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U804 ( .A(KEYINPUT57), .B(G953), .Z(n1130) );
XOR2_X1 U805 ( .A(n1132), .B(n1133), .Z(n1128) );
NOR2_X1 U806 ( .A1(KEYINPUT45), .A2(G140), .ZN(n1133) );
XOR2_X1 U807 ( .A(n1134), .B(n1135), .Z(n1132) );
NOR2_X1 U808 ( .A1(KEYINPUT35), .A2(n1136), .ZN(n1135) );
XOR2_X1 U809 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U810 ( .A1(KEYINPUT44), .A2(n1139), .ZN(n1137) );
XOR2_X1 U811 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U812 ( .A1(KEYINPUT13), .A2(n1142), .ZN(n1140) );
NAND2_X1 U813 ( .A1(n1127), .A2(n1143), .ZN(n1122) );
XOR2_X1 U814 ( .A(n1144), .B(n1145), .Z(G69) );
NOR2_X1 U815 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U816 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U817 ( .A(KEYINPUT33), .B(n1150), .Z(n1149) );
NOR2_X1 U818 ( .A1(n1151), .A2(n1152), .ZN(n1148) );
NOR3_X1 U819 ( .A1(n1152), .A2(n1150), .A3(n1151), .ZN(n1146) );
AND2_X1 U820 ( .A1(n1153), .A2(n1127), .ZN(n1150) );
NAND2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U822 ( .A1(G953), .A2(n1156), .ZN(n1144) );
NAND2_X1 U823 ( .A1(G898), .A2(n1157), .ZN(n1156) );
XOR2_X1 U824 ( .A(KEYINPUT37), .B(G224), .Z(n1157) );
NOR3_X1 U825 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(G66) );
AND2_X1 U826 ( .A1(KEYINPUT56), .A2(n1161), .ZN(n1160) );
NOR3_X1 U827 ( .A1(KEYINPUT56), .A2(G953), .A3(G952), .ZN(n1159) );
XNOR2_X1 U828 ( .A(n1162), .B(n1114), .ZN(n1158) );
NAND2_X1 U829 ( .A1(n1163), .A2(n1112), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1161), .A2(n1164), .ZN(G63) );
XOR2_X1 U831 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U832 ( .A(KEYINPUT14), .B(n1167), .Z(n1166) );
AND2_X1 U833 ( .A1(G478), .A2(n1163), .ZN(n1167) );
NAND2_X1 U834 ( .A1(KEYINPUT11), .A2(n1168), .ZN(n1165) );
NOR2_X1 U835 ( .A1(n1161), .A2(n1169), .ZN(G60) );
XOR2_X1 U836 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U837 ( .A1(n1163), .A2(G475), .ZN(n1170) );
XNOR2_X1 U838 ( .A(G104), .B(n1172), .ZN(G6) );
NOR2_X1 U839 ( .A1(n1161), .A2(n1173), .ZN(G57) );
XOR2_X1 U840 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U841 ( .A(n1176), .B(n1177), .ZN(n1175) );
XOR2_X1 U842 ( .A(n1178), .B(n1179), .Z(n1174) );
INV_X1 U843 ( .A(n1180), .ZN(n1179) );
XOR2_X1 U844 ( .A(n1181), .B(n1182), .Z(n1178) );
NAND2_X1 U845 ( .A1(n1163), .A2(G472), .ZN(n1181) );
NOR2_X1 U846 ( .A1(n1161), .A2(n1183), .ZN(G54) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(n1183) );
XNOR2_X1 U848 ( .A(n1186), .B(n1187), .ZN(n1185) );
XOR2_X1 U849 ( .A(n1188), .B(n1189), .Z(n1184) );
XOR2_X1 U850 ( .A(n1190), .B(n1191), .Z(n1189) );
NAND2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NAND2_X1 U852 ( .A1(G140), .A2(n1194), .ZN(n1193) );
XOR2_X1 U853 ( .A(KEYINPUT22), .B(n1195), .Z(n1192) );
NOR2_X1 U854 ( .A1(G140), .A2(n1194), .ZN(n1195) );
NAND2_X1 U855 ( .A1(n1163), .A2(G469), .ZN(n1188) );
INV_X1 U856 ( .A(n1196), .ZN(n1163) );
NOR2_X1 U857 ( .A1(n1161), .A2(n1197), .ZN(G51) );
XOR2_X1 U858 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U859 ( .A(n1200), .B(n1201), .ZN(n1199) );
NOR3_X1 U860 ( .A1(n1196), .A2(KEYINPUT43), .A3(n1202), .ZN(n1201) );
NAND2_X1 U861 ( .A1(G902), .A2(n1068), .ZN(n1196) );
NAND3_X1 U862 ( .A1(n1154), .A2(n1203), .A3(n1204), .ZN(n1068) );
INV_X1 U863 ( .A(n1143), .ZN(n1204) );
NAND4_X1 U864 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1143) );
AND4_X1 U865 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
NOR3_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1207) );
NOR4_X1 U867 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
AND2_X1 U868 ( .A1(n1216), .A2(n1220), .ZN(n1214) );
INV_X1 U869 ( .A(KEYINPUT30), .ZN(n1216) );
NAND2_X1 U870 ( .A1(n1221), .A2(n1222), .ZN(n1205) );
XOR2_X1 U871 ( .A(n1223), .B(KEYINPUT58), .Z(n1221) );
XOR2_X1 U872 ( .A(KEYINPUT20), .B(n1155), .Z(n1203) );
AND3_X1 U873 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1155) );
NAND2_X1 U874 ( .A1(n1092), .A2(n1227), .ZN(n1226) );
NAND2_X1 U875 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND4_X1 U876 ( .A1(n1230), .A2(n1101), .A3(n1084), .A4(n1231), .ZN(n1229) );
XOR2_X1 U877 ( .A(n1232), .B(KEYINPUT55), .Z(n1228) );
AND4_X1 U878 ( .A1(n1172), .A2(n1233), .A3(n1234), .A4(n1063), .ZN(n1154) );
NAND3_X1 U879 ( .A1(n1100), .A2(n1235), .A3(n1236), .ZN(n1063) );
NAND2_X1 U880 ( .A1(n1237), .A2(n1238), .ZN(n1234) );
XOR2_X1 U881 ( .A(KEYINPUT10), .B(n1239), .Z(n1238) );
NAND4_X1 U882 ( .A1(n1097), .A2(n1082), .A3(n1240), .A4(n1231), .ZN(n1233) );
XOR2_X1 U883 ( .A(KEYINPUT5), .B(n1092), .Z(n1240) );
NAND3_X1 U884 ( .A1(n1236), .A2(n1235), .A3(n1101), .ZN(n1172) );
NOR2_X1 U885 ( .A1(KEYINPUT34), .A2(n1241), .ZN(n1200) );
XOR2_X1 U886 ( .A(n1180), .B(G125), .Z(n1241) );
NOR2_X1 U887 ( .A1(n1127), .A2(G952), .ZN(n1161) );
XOR2_X1 U888 ( .A(n1242), .B(G146), .Z(G48) );
NAND2_X1 U889 ( .A1(KEYINPUT59), .A2(n1206), .ZN(n1242) );
NAND3_X1 U890 ( .A1(n1101), .A2(n1092), .A3(n1243), .ZN(n1206) );
XNOR2_X1 U891 ( .A(G143), .B(n1244), .ZN(G45) );
NAND2_X1 U892 ( .A1(n1222), .A2(n1092), .ZN(n1244) );
NOR2_X1 U893 ( .A1(n1217), .A2(n1245), .ZN(n1222) );
INV_X1 U894 ( .A(n1246), .ZN(n1245) );
XNOR2_X1 U895 ( .A(G140), .B(n1211), .ZN(G42) );
NAND4_X1 U896 ( .A1(n1247), .A2(n1101), .A3(n1248), .A4(n1218), .ZN(n1211) );
XOR2_X1 U897 ( .A(n1142), .B(n1212), .Z(G39) );
NAND3_X1 U898 ( .A1(n1243), .A2(n1218), .A3(n1239), .ZN(n1212) );
INV_X1 U899 ( .A(n1079), .ZN(n1218) );
NAND2_X1 U900 ( .A1(n1249), .A2(n1250), .ZN(G36) );
NAND2_X1 U901 ( .A1(n1220), .A2(n1251), .ZN(n1250) );
XOR2_X1 U902 ( .A(KEYINPUT48), .B(n1252), .Z(n1249) );
NOR2_X1 U903 ( .A1(n1220), .A2(n1251), .ZN(n1252) );
INV_X1 U904 ( .A(G134), .ZN(n1251) );
NOR3_X1 U905 ( .A1(n1079), .A2(n1219), .A3(n1217), .ZN(n1220) );
XOR2_X1 U906 ( .A(n1253), .B(n1254), .Z(G33) );
NAND2_X1 U907 ( .A1(KEYINPUT54), .A2(n1213), .ZN(n1254) );
NOR3_X1 U908 ( .A1(n1255), .A2(n1079), .A3(n1217), .ZN(n1213) );
NAND3_X1 U909 ( .A1(n1082), .A2(n1256), .A3(n1230), .ZN(n1217) );
NAND2_X1 U910 ( .A1(n1257), .A2(n1093), .ZN(n1079) );
XNOR2_X1 U911 ( .A(G128), .B(n1210), .ZN(G30) );
NAND3_X1 U912 ( .A1(n1100), .A2(n1092), .A3(n1243), .ZN(n1210) );
AND2_X1 U913 ( .A1(n1247), .A2(n1258), .ZN(n1243) );
AND3_X1 U914 ( .A1(n1256), .A2(n1259), .A3(n1082), .ZN(n1247) );
XNOR2_X1 U915 ( .A(G101), .B(n1260), .ZN(G3) );
NAND2_X1 U916 ( .A1(n1237), .A2(n1239), .ZN(n1260) );
NOR2_X1 U917 ( .A1(n1102), .A2(n1261), .ZN(n1237) );
XOR2_X1 U918 ( .A(n1134), .B(n1209), .Z(G27) );
NAND4_X1 U919 ( .A1(n1248), .A2(n1092), .A3(n1101), .A4(n1262), .ZN(n1209) );
AND3_X1 U920 ( .A1(n1084), .A2(n1259), .A3(n1256), .ZN(n1262) );
NAND2_X1 U921 ( .A1(n1070), .A2(n1263), .ZN(n1256) );
NAND4_X1 U922 ( .A1(G953), .A2(G902), .A3(n1264), .A4(n1131), .ZN(n1263) );
INV_X1 U923 ( .A(G900), .ZN(n1131) );
XOR2_X1 U924 ( .A(G122), .B(n1265), .Z(G24) );
NOR2_X1 U925 ( .A1(n1223), .A2(n1232), .ZN(n1265) );
NAND4_X1 U926 ( .A1(n1235), .A2(n1246), .A3(n1084), .A4(n1231), .ZN(n1232) );
NAND2_X1 U927 ( .A1(n1266), .A2(n1267), .ZN(n1246) );
OR2_X1 U928 ( .A1(n1255), .A2(KEYINPUT15), .ZN(n1267) );
NAND3_X1 U929 ( .A1(n1268), .A2(n1269), .A3(KEYINPUT15), .ZN(n1266) );
INV_X1 U930 ( .A(n1075), .ZN(n1235) );
NAND2_X1 U931 ( .A1(n1270), .A2(n1248), .ZN(n1075) );
XOR2_X1 U932 ( .A(n1271), .B(n1224), .Z(G21) );
NAND4_X1 U933 ( .A1(n1272), .A2(n1239), .A3(n1258), .A4(n1259), .ZN(n1224) );
XOR2_X1 U934 ( .A(n1273), .B(n1225), .Z(G18) );
NAND3_X1 U935 ( .A1(n1230), .A2(n1100), .A3(n1272), .ZN(n1225) );
INV_X1 U936 ( .A(n1274), .ZN(n1272) );
INV_X1 U937 ( .A(n1219), .ZN(n1100) );
NAND2_X1 U938 ( .A1(n1275), .A2(n1276), .ZN(n1219) );
XNOR2_X1 U939 ( .A(KEYINPUT15), .B(n1268), .ZN(n1275) );
INV_X1 U940 ( .A(n1102), .ZN(n1230) );
XOR2_X1 U941 ( .A(G113), .B(n1277), .Z(G15) );
NOR4_X1 U942 ( .A1(KEYINPUT39), .A2(n1255), .A3(n1102), .A4(n1274), .ZN(n1277) );
NAND3_X1 U943 ( .A1(n1084), .A2(n1231), .A3(n1092), .ZN(n1274) );
NAND2_X1 U944 ( .A1(n1278), .A2(n1279), .ZN(n1084) );
NAND3_X1 U945 ( .A1(n1086), .A2(n1280), .A3(n1087), .ZN(n1279) );
INV_X1 U946 ( .A(KEYINPUT41), .ZN(n1087) );
NAND2_X1 U947 ( .A1(KEYINPUT41), .A2(n1082), .ZN(n1278) );
NAND2_X1 U948 ( .A1(n1270), .A2(n1258), .ZN(n1102) );
XOR2_X1 U949 ( .A(n1259), .B(KEYINPUT17), .Z(n1270) );
INV_X1 U950 ( .A(n1281), .ZN(n1259) );
INV_X1 U951 ( .A(n1101), .ZN(n1255) );
NOR2_X1 U952 ( .A1(n1268), .A2(n1276), .ZN(n1101) );
XOR2_X1 U953 ( .A(G110), .B(n1282), .Z(G12) );
AND2_X1 U954 ( .A1(n1236), .A2(n1097), .ZN(n1282) );
NOR3_X1 U955 ( .A1(n1258), .A2(n1281), .A3(n1073), .ZN(n1097) );
INV_X1 U956 ( .A(n1239), .ZN(n1073) );
NOR2_X1 U957 ( .A1(n1269), .A2(n1268), .ZN(n1239) );
XOR2_X1 U958 ( .A(n1116), .B(KEYINPUT9), .Z(n1268) );
XOR2_X1 U959 ( .A(G478), .B(n1283), .Z(n1116) );
NOR2_X1 U960 ( .A1(G902), .A2(n1168), .ZN(n1283) );
NAND3_X1 U961 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1168) );
NAND2_X1 U962 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
INV_X1 U963 ( .A(KEYINPUT1), .ZN(n1288) );
NAND3_X1 U964 ( .A1(KEYINPUT1), .A2(n1289), .A3(n1290), .ZN(n1285) );
OR2_X1 U965 ( .A1(n1290), .A2(n1289), .ZN(n1284) );
AND3_X1 U966 ( .A1(G234), .A2(n1127), .A3(G217), .ZN(n1289) );
NOR2_X1 U967 ( .A1(KEYINPUT6), .A2(n1287), .ZN(n1290) );
XNOR2_X1 U968 ( .A(n1291), .B(n1292), .ZN(n1287) );
XOR2_X1 U969 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U970 ( .A(G116), .B(G107), .Z(n1294) );
XNOR2_X1 U971 ( .A(G122), .B(n1295), .ZN(n1291) );
XOR2_X1 U972 ( .A(KEYINPUT12), .B(G134), .Z(n1295) );
INV_X1 U973 ( .A(n1276), .ZN(n1269) );
XOR2_X1 U974 ( .A(n1109), .B(G475), .Z(n1276) );
NAND2_X1 U975 ( .A1(n1296), .A2(n1297), .ZN(n1109) );
XOR2_X1 U976 ( .A(KEYINPUT4), .B(n1298), .Z(n1296) );
INV_X1 U977 ( .A(n1171), .ZN(n1298) );
XOR2_X1 U978 ( .A(n1299), .B(n1300), .Z(n1171) );
XOR2_X1 U979 ( .A(G122), .B(G113), .Z(n1300) );
XOR2_X1 U980 ( .A(n1301), .B(G104), .Z(n1299) );
NAND2_X1 U981 ( .A1(KEYINPUT18), .A2(n1302), .ZN(n1301) );
XOR2_X1 U982 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U983 ( .A(n1305), .B(n1306), .Z(n1304) );
NAND2_X1 U984 ( .A1(KEYINPUT7), .A2(n1253), .ZN(n1305) );
INV_X1 U985 ( .A(G131), .ZN(n1253) );
XOR2_X1 U986 ( .A(G143), .B(n1307), .Z(n1303) );
AND3_X1 U987 ( .A1(G214), .A2(n1127), .A3(n1308), .ZN(n1307) );
NOR2_X1 U988 ( .A1(n1309), .A2(n1105), .ZN(n1281) );
NOR3_X1 U989 ( .A1(n1112), .A2(G902), .A3(n1114), .ZN(n1105) );
AND2_X1 U990 ( .A1(n1112), .A2(n1310), .ZN(n1309) );
OR2_X1 U991 ( .A1(n1114), .A2(G902), .ZN(n1310) );
XOR2_X1 U992 ( .A(n1311), .B(n1312), .Z(n1114) );
XOR2_X1 U993 ( .A(G110), .B(n1313), .Z(n1312) );
XOR2_X1 U994 ( .A(KEYINPUT36), .B(G137), .Z(n1313) );
XOR2_X1 U995 ( .A(n1314), .B(n1315), .Z(n1311) );
NOR2_X1 U996 ( .A1(KEYINPUT47), .A2(n1306), .ZN(n1315) );
XOR2_X1 U997 ( .A(n1316), .B(n1317), .Z(n1306) );
XOR2_X1 U998 ( .A(KEYINPUT8), .B(G146), .Z(n1317) );
XOR2_X1 U999 ( .A(n1134), .B(G140), .Z(n1316) );
INV_X1 U1000 ( .A(G125), .ZN(n1134) );
XNOR2_X1 U1001 ( .A(n1318), .B(n1319), .ZN(n1314) );
NAND2_X1 U1002 ( .A1(KEYINPUT28), .A2(n1320), .ZN(n1319) );
NAND3_X1 U1003 ( .A1(G234), .A2(n1127), .A3(G221), .ZN(n1320) );
NAND2_X1 U1004 ( .A1(KEYINPUT3), .A2(n1321), .ZN(n1318) );
XOR2_X1 U1005 ( .A(G119), .B(n1322), .Z(n1321) );
XOR2_X1 U1006 ( .A(KEYINPUT32), .B(G128), .Z(n1322) );
AND2_X1 U1007 ( .A1(G217), .A2(n1323), .ZN(n1112) );
INV_X1 U1008 ( .A(n1248), .ZN(n1258) );
XOR2_X1 U1009 ( .A(n1324), .B(n1325), .Z(n1248) );
NOR2_X1 U1010 ( .A1(KEYINPUT38), .A2(n1118), .ZN(n1325) );
AND2_X1 U1011 ( .A1(n1326), .A2(n1297), .ZN(n1118) );
XOR2_X1 U1012 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1013 ( .A(n1329), .B(n1176), .Z(n1328) );
XNOR2_X1 U1014 ( .A(n1330), .B(G101), .ZN(n1176) );
NAND2_X1 U1015 ( .A1(KEYINPUT0), .A2(n1182), .ZN(n1329) );
AND3_X1 U1016 ( .A1(n1331), .A2(n1308), .A3(G210), .ZN(n1182) );
XOR2_X1 U1017 ( .A(KEYINPUT53), .B(G953), .Z(n1331) );
XNOR2_X1 U1018 ( .A(n1332), .B(n1333), .ZN(n1327) );
NAND2_X1 U1019 ( .A1(KEYINPUT27), .A2(n1180), .ZN(n1333) );
NAND2_X1 U1020 ( .A1(KEYINPUT24), .A2(n1177), .ZN(n1332) );
AND2_X1 U1021 ( .A1(n1334), .A2(n1335), .ZN(n1177) );
NAND2_X1 U1022 ( .A1(G113), .A2(n1336), .ZN(n1335) );
NAND2_X1 U1023 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND3_X1 U1024 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1334) );
XOR2_X1 U1025 ( .A(n1340), .B(KEYINPUT42), .Z(n1337) );
NAND2_X1 U1026 ( .A1(n1341), .A2(n1273), .ZN(n1340) );
INV_X1 U1027 ( .A(G116), .ZN(n1273) );
XOR2_X1 U1028 ( .A(KEYINPUT51), .B(G119), .Z(n1341) );
XNOR2_X1 U1029 ( .A(G472), .B(KEYINPUT40), .ZN(n1324) );
INV_X1 U1030 ( .A(n1261), .ZN(n1236) );
NAND3_X1 U1031 ( .A1(n1092), .A2(n1231), .A3(n1082), .ZN(n1261) );
NOR2_X1 U1032 ( .A1(n1086), .A2(n1088), .ZN(n1082) );
INV_X1 U1033 ( .A(n1280), .ZN(n1088) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1323), .ZN(n1280) );
NAND2_X1 U1035 ( .A1(G234), .A2(n1342), .ZN(n1323) );
XOR2_X1 U1036 ( .A(n1120), .B(G469), .Z(n1086) );
NAND2_X1 U1037 ( .A1(n1343), .A2(n1297), .ZN(n1120) );
XOR2_X1 U1038 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1039 ( .A(n1187), .B(n1346), .ZN(n1345) );
XNOR2_X1 U1040 ( .A(n1190), .B(n1347), .ZN(n1346) );
NOR2_X1 U1041 ( .A1(KEYINPUT16), .A2(n1186), .ZN(n1347) );
NAND2_X1 U1042 ( .A1(G227), .A2(n1127), .ZN(n1190) );
XNOR2_X1 U1043 ( .A(n1138), .B(n1330), .ZN(n1187) );
XNOR2_X1 U1044 ( .A(n1142), .B(n1141), .ZN(n1330) );
XOR2_X1 U1045 ( .A(G131), .B(G134), .Z(n1141) );
INV_X1 U1046 ( .A(G137), .ZN(n1142) );
XNOR2_X1 U1047 ( .A(n1348), .B(n1293), .ZN(n1138) );
XOR2_X1 U1048 ( .A(G128), .B(G143), .Z(n1293) );
NAND2_X1 U1049 ( .A1(KEYINPUT25), .A2(n1349), .ZN(n1348) );
XOR2_X1 U1050 ( .A(n1194), .B(n1350), .Z(n1344) );
XOR2_X1 U1051 ( .A(KEYINPUT19), .B(G140), .Z(n1350) );
NAND2_X1 U1052 ( .A1(n1070), .A2(n1351), .ZN(n1231) );
NAND3_X1 U1053 ( .A1(G902), .A2(n1264), .A3(n1151), .ZN(n1351) );
NOR2_X1 U1054 ( .A1(n1127), .A2(G898), .ZN(n1151) );
NAND3_X1 U1055 ( .A1(n1264), .A2(n1127), .A3(G952), .ZN(n1070) );
NAND2_X1 U1056 ( .A1(G237), .A2(G234), .ZN(n1264) );
INV_X1 U1057 ( .A(n1223), .ZN(n1092) );
NAND2_X1 U1058 ( .A1(n1094), .A2(n1093), .ZN(n1223) );
NAND2_X1 U1059 ( .A1(G214), .A2(n1352), .ZN(n1093) );
INV_X1 U1060 ( .A(n1257), .ZN(n1094) );
XNOR2_X1 U1061 ( .A(n1353), .B(n1202), .ZN(n1257) );
NAND2_X1 U1062 ( .A1(G210), .A2(n1352), .ZN(n1202) );
NAND2_X1 U1063 ( .A1(n1342), .A2(n1308), .ZN(n1352) );
INV_X1 U1064 ( .A(G237), .ZN(n1308) );
XOR2_X1 U1065 ( .A(G902), .B(KEYINPUT31), .Z(n1342) );
NAND2_X1 U1066 ( .A1(n1354), .A2(n1297), .ZN(n1353) );
INV_X1 U1067 ( .A(G902), .ZN(n1297) );
XOR2_X1 U1068 ( .A(n1198), .B(n1355), .Z(n1354) );
XOR2_X1 U1069 ( .A(G125), .B(n1356), .Z(n1355) );
NOR2_X1 U1070 ( .A1(KEYINPUT50), .A2(n1180), .ZN(n1356) );
XOR2_X1 U1071 ( .A(n1357), .B(G128), .Z(n1180) );
NAND3_X1 U1072 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1357) );
NAND2_X1 U1073 ( .A1(KEYINPUT63), .A2(G143), .ZN(n1360) );
NAND3_X1 U1074 ( .A1(n1361), .A2(n1362), .A3(n1349), .ZN(n1359) );
INV_X1 U1075 ( .A(KEYINPUT63), .ZN(n1362) );
OR2_X1 U1076 ( .A1(n1349), .A2(n1361), .ZN(n1358) );
NOR2_X1 U1077 ( .A1(G143), .A2(KEYINPUT26), .ZN(n1361) );
INV_X1 U1078 ( .A(G146), .ZN(n1349) );
NAND2_X1 U1079 ( .A1(n1363), .A2(n1364), .ZN(n1198) );
NAND2_X1 U1080 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
INV_X1 U1081 ( .A(KEYINPUT62), .ZN(n1366) );
XOR2_X1 U1082 ( .A(n1367), .B(n1368), .Z(n1365) );
NAND2_X1 U1083 ( .A1(KEYINPUT62), .A2(n1369), .ZN(n1363) );
XOR2_X1 U1084 ( .A(n1152), .B(n1368), .Z(n1369) );
AND2_X1 U1085 ( .A1(G224), .A2(n1127), .ZN(n1368) );
INV_X1 U1086 ( .A(G953), .ZN(n1127) );
NAND2_X1 U1087 ( .A1(n1367), .A2(n1370), .ZN(n1152) );
OR2_X1 U1088 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
NAND2_X1 U1089 ( .A1(n1372), .A2(n1371), .ZN(n1367) );
XNOR2_X1 U1090 ( .A(n1373), .B(G122), .ZN(n1371) );
NAND2_X1 U1091 ( .A1(KEYINPUT2), .A2(n1194), .ZN(n1373) );
INV_X1 U1092 ( .A(G110), .ZN(n1194) );
XNOR2_X1 U1093 ( .A(n1374), .B(n1375), .ZN(n1372) );
NOR2_X1 U1094 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
NOR2_X1 U1095 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
INV_X1 U1096 ( .A(KEYINPUT52), .ZN(n1379) );
XOR2_X1 U1097 ( .A(G119), .B(G116), .Z(n1378) );
NOR2_X1 U1098 ( .A1(KEYINPUT52), .A2(n1380), .ZN(n1376) );
NOR2_X1 U1099 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
INV_X1 U1100 ( .A(n1338), .ZN(n1382) );
NAND2_X1 U1101 ( .A1(G116), .A2(n1271), .ZN(n1338) );
NOR2_X1 U1102 ( .A1(G116), .A2(n1271), .ZN(n1381) );
INV_X1 U1103 ( .A(G119), .ZN(n1271) );
XOR2_X1 U1104 ( .A(n1339), .B(n1186), .Z(n1374) );
XNOR2_X1 U1105 ( .A(n1383), .B(n1384), .ZN(n1186) );
XOR2_X1 U1106 ( .A(KEYINPUT60), .B(G107), .Z(n1384) );
XNOR2_X1 U1107 ( .A(G101), .B(G104), .ZN(n1383) );
INV_X1 U1108 ( .A(G113), .ZN(n1339) );
endmodule


