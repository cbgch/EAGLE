//Key = 0111100011011100010011110000111101011100111001110010111110010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369;

XOR2_X1 U757 ( .A(G107), .B(n1039), .Z(G9) );
NOR2_X1 U758 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR3_X1 U759 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NOR3_X1 U760 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1043) );
NOR2_X1 U761 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U762 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U763 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
XOR2_X1 U764 ( .A(n1054), .B(KEYINPUT47), .Z(n1053) );
NAND2_X1 U765 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XNOR2_X1 U766 ( .A(n1057), .B(KEYINPUT36), .ZN(n1055) );
NOR3_X1 U767 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1048) );
NOR3_X1 U768 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR2_X1 U769 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U770 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1068), .A2(n1069), .ZN(n1062) );
NOR2_X1 U772 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR3_X1 U773 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1070) );
INV_X1 U774 ( .A(KEYINPUT52), .ZN(n1072) );
NOR2_X1 U775 ( .A1(n1075), .A2(n1076), .ZN(n1059) );
NOR4_X1 U776 ( .A1(KEYINPUT52), .A2(n1074), .A3(n1069), .A4(n1073), .ZN(n1076) );
NAND3_X1 U777 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1042) );
NAND3_X1 U778 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
INV_X1 U779 ( .A(n1051), .ZN(n1082) );
NAND3_X1 U780 ( .A1(n1083), .A2(n1084), .A3(n1075), .ZN(n1051) );
INV_X1 U781 ( .A(n1061), .ZN(n1075) );
OR2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
NOR3_X1 U783 ( .A1(n1087), .A2(G953), .A3(G952), .ZN(n1040) );
INV_X1 U784 ( .A(n1077), .ZN(n1087) );
NAND4_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1077) );
NOR4_X1 U786 ( .A1(n1092), .A2(n1056), .A3(n1093), .A4(n1094), .ZN(n1091) );
XOR2_X1 U787 ( .A(n1095), .B(KEYINPUT23), .Z(n1094) );
AND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NOR2_X1 U789 ( .A1(n1065), .A2(n1098), .ZN(n1090) );
XOR2_X1 U790 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U791 ( .A(KEYINPUT31), .B(n1045), .Z(n1089) );
XOR2_X1 U792 ( .A(n1101), .B(n1102), .Z(G72) );
XOR2_X1 U793 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U796 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1107) );
NOR2_X1 U798 ( .A1(G953), .A2(n1113), .ZN(n1103) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1078), .ZN(n1101) );
AND2_X1 U800 ( .A1(G227), .A2(G900), .ZN(n1114) );
NAND2_X1 U801 ( .A1(n1115), .A2(n1116), .ZN(G69) );
NAND2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U803 ( .A1(G953), .A2(n1119), .ZN(n1117) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1119) );
NAND2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NAND2_X1 U806 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
OR2_X1 U807 ( .A1(n1078), .A2(G224), .ZN(n1123) );
INV_X1 U808 ( .A(n1118), .ZN(n1120) );
NAND3_X1 U809 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1118) );
NAND2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
OR3_X1 U811 ( .A1(n1128), .A2(n1127), .A3(KEYINPUT7), .ZN(n1125) );
AND2_X1 U812 ( .A1(KEYINPUT45), .A2(n1129), .ZN(n1128) );
NAND2_X1 U813 ( .A1(KEYINPUT7), .A2(n1130), .ZN(n1124) );
OR2_X1 U814 ( .A1(n1129), .A2(n1127), .ZN(n1130) );
AND2_X1 U815 ( .A1(n1131), .A2(n1122), .ZN(n1127) );
INV_X1 U816 ( .A(n1132), .ZN(n1122) );
XOR2_X1 U817 ( .A(n1133), .B(n1134), .Z(n1131) );
NAND2_X1 U818 ( .A1(n1135), .A2(KEYINPUT54), .ZN(n1133) );
XOR2_X1 U819 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U820 ( .A1(n1078), .A2(n1138), .ZN(n1129) );
NAND2_X1 U821 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U822 ( .A(KEYINPUT4), .B(n1141), .ZN(n1140) );
NOR2_X1 U823 ( .A1(n1142), .A2(n1143), .ZN(G66) );
XNOR2_X1 U824 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U825 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U826 ( .A1(n1142), .A2(n1148), .ZN(G63) );
XNOR2_X1 U827 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U828 ( .A1(n1151), .A2(n1147), .ZN(n1150) );
INV_X1 U829 ( .A(G478), .ZN(n1151) );
NOR2_X1 U830 ( .A1(n1142), .A2(n1152), .ZN(G60) );
XOR2_X1 U831 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U832 ( .A1(n1099), .A2(n1147), .ZN(n1153) );
XNOR2_X1 U833 ( .A(G104), .B(n1155), .ZN(G6) );
NOR2_X1 U834 ( .A1(n1142), .A2(n1156), .ZN(G57) );
XOR2_X1 U835 ( .A(n1157), .B(KEYINPUT21), .Z(n1156) );
NAND2_X1 U836 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U837 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U838 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U839 ( .A(n1164), .B(n1165), .ZN(n1160) );
XOR2_X1 U840 ( .A(n1166), .B(KEYINPUT48), .Z(n1158) );
NAND2_X1 U841 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U842 ( .A(n1164), .B(n1165), .Z(n1168) );
XNOR2_X1 U843 ( .A(n1169), .B(n1170), .ZN(n1165) );
NOR2_X1 U844 ( .A1(n1171), .A2(n1147), .ZN(n1170) );
INV_X1 U845 ( .A(G472), .ZN(n1171) );
XOR2_X1 U846 ( .A(n1163), .B(G101), .Z(n1167) );
NOR2_X1 U847 ( .A1(n1142), .A2(n1172), .ZN(G54) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1147), .ZN(n1174) );
NAND2_X1 U850 ( .A1(G902), .A2(n1044), .ZN(n1147) );
INV_X1 U851 ( .A(G469), .ZN(n1175) );
NAND2_X1 U852 ( .A1(n1176), .A2(KEYINPUT17), .ZN(n1173) );
XOR2_X1 U853 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U854 ( .A(KEYINPUT12), .B(G110), .Z(n1178) );
XOR2_X1 U855 ( .A(n1179), .B(n1180), .Z(n1177) );
NAND2_X1 U856 ( .A1(KEYINPUT56), .A2(n1181), .ZN(n1179) );
NOR2_X1 U857 ( .A1(n1142), .A2(n1182), .ZN(G51) );
XOR2_X1 U858 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND3_X1 U859 ( .A1(G902), .A2(n1185), .A3(n1097), .ZN(n1184) );
XNOR2_X1 U860 ( .A(KEYINPUT50), .B(n1044), .ZN(n1185) );
NAND3_X1 U861 ( .A1(n1139), .A2(n1141), .A3(n1113), .ZN(n1044) );
AND4_X1 U862 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1113) );
NOR4_X1 U863 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
NOR2_X1 U864 ( .A1(n1058), .A2(n1194), .ZN(n1193) );
XNOR2_X1 U865 ( .A(n1195), .B(KEYINPUT19), .ZN(n1194) );
INV_X1 U866 ( .A(n1080), .ZN(n1058) );
NOR2_X1 U867 ( .A1(n1196), .A2(n1197), .ZN(n1188) );
INV_X1 U868 ( .A(n1198), .ZN(n1197) );
NAND2_X1 U869 ( .A1(n1052), .A2(n1199), .ZN(n1187) );
NAND2_X1 U870 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND3_X1 U871 ( .A1(n1086), .A2(n1084), .A3(n1202), .ZN(n1201) );
NOR3_X1 U872 ( .A1(n1203), .A2(KEYINPUT42), .A3(n1066), .ZN(n1202) );
XOR2_X1 U873 ( .A(KEYINPUT22), .B(n1204), .Z(n1200) );
NAND2_X1 U874 ( .A1(KEYINPUT42), .A2(n1205), .ZN(n1186) );
AND4_X1 U875 ( .A1(n1155), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1139) );
NOR4_X1 U876 ( .A1(n1209), .A2(n1210), .A3(n1039), .A4(n1211), .ZN(n1208) );
AND4_X1 U877 ( .A1(n1095), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1039) );
AND3_X1 U878 ( .A1(n1052), .A2(n1071), .A3(n1067), .ZN(n1214) );
OR2_X1 U879 ( .A1(n1215), .A2(n1216), .ZN(n1207) );
NAND4_X1 U880 ( .A1(n1217), .A2(n1071), .A3(n1095), .A4(n1212), .ZN(n1155) );
NAND2_X1 U881 ( .A1(KEYINPUT40), .A2(n1218), .ZN(n1183) );
XOR2_X1 U882 ( .A(n1219), .B(n1220), .Z(n1218) );
XNOR2_X1 U883 ( .A(n1221), .B(n1222), .ZN(n1220) );
XOR2_X1 U884 ( .A(n1223), .B(n1224), .Z(n1219) );
XOR2_X1 U885 ( .A(n1225), .B(KEYINPUT62), .Z(n1224) );
NAND2_X1 U886 ( .A1(KEYINPUT35), .A2(n1226), .ZN(n1223) );
NOR2_X1 U887 ( .A1(n1078), .A2(G952), .ZN(n1142) );
XOR2_X1 U888 ( .A(G146), .B(n1192), .Z(G48) );
AND3_X1 U889 ( .A1(n1066), .A2(n1052), .A3(n1227), .ZN(n1192) );
NAND2_X1 U890 ( .A1(n1228), .A2(n1229), .ZN(G45) );
OR2_X1 U891 ( .A1(n1230), .A2(G143), .ZN(n1229) );
NAND2_X1 U892 ( .A1(G143), .A2(n1231), .ZN(n1228) );
NAND2_X1 U893 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND2_X1 U894 ( .A1(n1191), .A2(n1234), .ZN(n1233) );
INV_X1 U895 ( .A(KEYINPUT55), .ZN(n1234) );
NAND2_X1 U896 ( .A1(KEYINPUT55), .A2(n1230), .ZN(n1232) );
NAND2_X1 U897 ( .A1(KEYINPUT30), .A2(n1191), .ZN(n1230) );
AND3_X1 U898 ( .A1(n1085), .A2(n1235), .A3(n1236), .ZN(n1191) );
NOR3_X1 U899 ( .A1(n1237), .A2(n1088), .A3(n1216), .ZN(n1236) );
XOR2_X1 U900 ( .A(G140), .B(n1190), .Z(G42) );
AND4_X1 U901 ( .A1(n1066), .A2(n1086), .A3(n1235), .A4(n1080), .ZN(n1190) );
XNOR2_X1 U902 ( .A(G137), .B(n1238), .ZN(G39) );
NAND2_X1 U903 ( .A1(n1195), .A2(n1080), .ZN(n1238) );
AND2_X1 U904 ( .A1(n1083), .A2(n1227), .ZN(n1195) );
NAND2_X1 U905 ( .A1(n1239), .A2(n1240), .ZN(G36) );
OR2_X1 U906 ( .A1(n1198), .A2(G134), .ZN(n1240) );
XOR2_X1 U907 ( .A(n1241), .B(KEYINPUT32), .Z(n1239) );
NAND2_X1 U908 ( .A1(G134), .A2(n1198), .ZN(n1241) );
NAND2_X1 U909 ( .A1(n1242), .A2(n1067), .ZN(n1198) );
XOR2_X1 U910 ( .A(G131), .B(n1196), .Z(G33) );
AND2_X1 U911 ( .A1(n1242), .A2(n1066), .ZN(n1196) );
AND3_X1 U912 ( .A1(n1235), .A2(n1080), .A3(n1085), .ZN(n1242) );
NAND2_X1 U913 ( .A1(n1243), .A2(n1244), .ZN(n1080) );
OR2_X1 U914 ( .A1(n1216), .A2(KEYINPUT36), .ZN(n1244) );
NAND3_X1 U915 ( .A1(n1057), .A2(n1245), .A3(KEYINPUT36), .ZN(n1243) );
XNOR2_X1 U916 ( .A(G128), .B(n1246), .ZN(G30) );
NAND2_X1 U917 ( .A1(n1204), .A2(n1052), .ZN(n1246) );
AND2_X1 U918 ( .A1(n1227), .A2(n1067), .ZN(n1204) );
AND3_X1 U919 ( .A1(n1047), .A2(n1045), .A3(n1235), .ZN(n1227) );
NOR2_X1 U920 ( .A1(n1247), .A2(n1203), .ZN(n1235) );
INV_X1 U921 ( .A(n1248), .ZN(n1203) );
XOR2_X1 U922 ( .A(G101), .B(n1249), .Z(G3) );
NOR2_X1 U923 ( .A1(KEYINPUT6), .A2(n1141), .ZN(n1249) );
NAND3_X1 U924 ( .A1(n1085), .A2(n1052), .A3(n1250), .ZN(n1141) );
XNOR2_X1 U925 ( .A(n1205), .B(n1251), .ZN(G27) );
NAND2_X1 U926 ( .A1(KEYINPUT63), .A2(G125), .ZN(n1251) );
AND4_X1 U927 ( .A1(n1217), .A2(n1084), .A3(n1047), .A4(n1248), .ZN(n1205) );
NAND2_X1 U928 ( .A1(n1061), .A2(n1252), .ZN(n1248) );
NAND3_X1 U929 ( .A1(G902), .A2(n1253), .A3(n1105), .ZN(n1252) );
NOR2_X1 U930 ( .A1(n1078), .A2(G900), .ZN(n1105) );
INV_X1 U931 ( .A(n1095), .ZN(n1047) );
AND3_X1 U932 ( .A1(n1213), .A2(n1052), .A3(n1066), .ZN(n1217) );
XNOR2_X1 U933 ( .A(G122), .B(n1206), .ZN(G24) );
NAND4_X1 U934 ( .A1(n1095), .A2(n1254), .A3(n1213), .A4(n1255), .ZN(n1206) );
NOR2_X1 U935 ( .A1(n1256), .A2(n1237), .ZN(n1255) );
NAND2_X1 U936 ( .A1(n1257), .A2(n1258), .ZN(G21) );
OR2_X1 U937 ( .A1(n1259), .A2(n1211), .ZN(n1258) );
XOR2_X1 U938 ( .A(n1260), .B(KEYINPUT57), .Z(n1257) );
NAND2_X1 U939 ( .A1(n1211), .A2(n1259), .ZN(n1260) );
INV_X1 U940 ( .A(G119), .ZN(n1259) );
NOR4_X1 U941 ( .A1(n1256), .A2(n1069), .A3(n1095), .A4(n1213), .ZN(n1211) );
XOR2_X1 U942 ( .A(n1261), .B(n1210), .Z(G18) );
AND3_X1 U943 ( .A1(n1085), .A2(n1067), .A3(n1262), .ZN(n1210) );
AND2_X1 U944 ( .A1(n1237), .A2(n1254), .ZN(n1067) );
NAND2_X1 U945 ( .A1(KEYINPUT11), .A2(n1263), .ZN(n1261) );
XOR2_X1 U946 ( .A(G113), .B(n1209), .Z(G15) );
AND3_X1 U947 ( .A1(n1085), .A2(n1066), .A3(n1262), .ZN(n1209) );
INV_X1 U948 ( .A(n1256), .ZN(n1262) );
NAND3_X1 U949 ( .A1(n1052), .A2(n1212), .A3(n1084), .ZN(n1256) );
INV_X1 U950 ( .A(n1065), .ZN(n1084) );
NAND2_X1 U951 ( .A1(n1264), .A2(n1073), .ZN(n1065) );
INV_X1 U952 ( .A(n1074), .ZN(n1264) );
NOR2_X1 U953 ( .A1(n1237), .A2(n1254), .ZN(n1066) );
INV_X1 U954 ( .A(n1088), .ZN(n1254) );
AND2_X1 U955 ( .A1(n1265), .A2(n1045), .ZN(n1085) );
XOR2_X1 U956 ( .A(n1095), .B(KEYINPUT26), .Z(n1265) );
XOR2_X1 U957 ( .A(n1266), .B(n1267), .Z(G12) );
NOR2_X1 U958 ( .A1(KEYINPUT44), .A2(n1268), .ZN(n1267) );
NOR2_X1 U959 ( .A1(n1269), .A2(n1216), .ZN(n1266) );
INV_X1 U960 ( .A(n1052), .ZN(n1216) );
NOR2_X1 U961 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
AND3_X1 U962 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1057) );
INV_X1 U963 ( .A(n1092), .ZN(n1272) );
NOR2_X1 U964 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
OR2_X1 U965 ( .A1(n1097), .A2(KEYINPUT53), .ZN(n1271) );
NAND3_X1 U966 ( .A1(n1097), .A2(n1096), .A3(KEYINPUT53), .ZN(n1270) );
NAND4_X1 U967 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1096) );
NAND2_X1 U968 ( .A1(KEYINPUT5), .A2(n1277), .ZN(n1276) );
NAND2_X1 U969 ( .A1(n1222), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U970 ( .A(KEYINPUT8), .B(n1279), .ZN(n1278) );
NAND2_X1 U971 ( .A1(n1280), .A2(n1281), .ZN(n1275) );
INV_X1 U972 ( .A(KEYINPUT5), .ZN(n1281) );
NAND2_X1 U973 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
OR2_X1 U974 ( .A1(n1279), .A2(KEYINPUT8), .ZN(n1283) );
NAND3_X1 U975 ( .A1(n1279), .A2(n1222), .A3(KEYINPUT8), .ZN(n1282) );
OR2_X1 U976 ( .A1(n1279), .A2(n1222), .ZN(n1273) );
XOR2_X1 U977 ( .A(n1284), .B(n1285), .Z(n1222) );
INV_X1 U978 ( .A(n1134), .ZN(n1285) );
XOR2_X1 U979 ( .A(n1268), .B(G122), .Z(n1134) );
INV_X1 U980 ( .A(G110), .ZN(n1268) );
XOR2_X1 U981 ( .A(n1136), .B(n1286), .Z(n1284) );
NOR2_X1 U982 ( .A1(KEYINPUT10), .A2(n1137), .ZN(n1286) );
XOR2_X1 U983 ( .A(n1287), .B(n1288), .Z(n1137) );
NOR2_X1 U984 ( .A1(G101), .A2(KEYINPUT34), .ZN(n1288) );
XOR2_X1 U985 ( .A(n1289), .B(n1290), .Z(n1136) );
NOR2_X1 U986 ( .A1(G119), .A2(KEYINPUT18), .ZN(n1290) );
XOR2_X1 U987 ( .A(G113), .B(n1263), .Z(n1289) );
XOR2_X1 U988 ( .A(n1291), .B(n1292), .Z(n1279) );
XNOR2_X1 U989 ( .A(n1225), .B(n1293), .ZN(n1292) );
NOR2_X1 U990 ( .A1(KEYINPUT27), .A2(n1221), .ZN(n1293) );
NAND2_X1 U991 ( .A1(G224), .A2(n1078), .ZN(n1225) );
XOR2_X1 U992 ( .A(n1226), .B(KEYINPUT39), .Z(n1291) );
AND2_X1 U993 ( .A1(G210), .A2(n1294), .ZN(n1097) );
INV_X1 U994 ( .A(n1245), .ZN(n1056) );
NAND2_X1 U995 ( .A1(G214), .A2(n1294), .ZN(n1245) );
NAND2_X1 U996 ( .A1(n1274), .A2(n1295), .ZN(n1294) );
XOR2_X1 U997 ( .A(n1215), .B(KEYINPUT43), .Z(n1269) );
NAND2_X1 U998 ( .A1(n1250), .A2(n1086), .ZN(n1215) );
NOR2_X1 U999 ( .A1(n1045), .A2(n1095), .ZN(n1086) );
XNOR2_X1 U1000 ( .A(n1296), .B(n1146), .ZN(n1095) );
NAND2_X1 U1001 ( .A1(G217), .A2(n1297), .ZN(n1146) );
NAND2_X1 U1002 ( .A1(n1144), .A2(n1274), .ZN(n1296) );
XNOR2_X1 U1003 ( .A(n1298), .B(n1299), .ZN(n1144) );
XOR2_X1 U1004 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U1005 ( .A(G128), .B(G119), .Z(n1301) );
XOR2_X1 U1006 ( .A(G146), .B(G137), .Z(n1300) );
XOR2_X1 U1007 ( .A(n1302), .B(n1109), .Z(n1298) );
INV_X1 U1008 ( .A(n1303), .ZN(n1109) );
XOR2_X1 U1009 ( .A(n1304), .B(G110), .Z(n1302) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1305), .ZN(n1304) );
INV_X1 U1011 ( .A(n1213), .ZN(n1045) );
XOR2_X1 U1012 ( .A(n1306), .B(G472), .Z(n1213) );
NAND3_X1 U1013 ( .A1(n1307), .A2(n1308), .A3(n1274), .ZN(n1306) );
NAND2_X1 U1014 ( .A1(n1309), .A2(n1162), .ZN(n1308) );
INV_X1 U1015 ( .A(G101), .ZN(n1162) );
XOR2_X1 U1016 ( .A(n1310), .B(KEYINPUT20), .Z(n1309) );
NAND2_X1 U1017 ( .A1(n1311), .A2(G101), .ZN(n1307) );
XOR2_X1 U1018 ( .A(KEYINPUT33), .B(n1312), .Z(n1311) );
INV_X1 U1019 ( .A(n1310), .ZN(n1312) );
XOR2_X1 U1020 ( .A(n1163), .B(n1313), .Z(n1310) );
XNOR2_X1 U1021 ( .A(n1314), .B(KEYINPUT3), .ZN(n1313) );
NAND2_X1 U1022 ( .A1(n1315), .A2(KEYINPUT9), .ZN(n1314) );
XOR2_X1 U1023 ( .A(n1316), .B(n1317), .Z(n1315) );
NAND2_X1 U1024 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
OR2_X1 U1025 ( .A1(n1164), .A2(KEYINPUT60), .ZN(n1319) );
XOR2_X1 U1026 ( .A(n1221), .B(n1320), .Z(n1164) );
INV_X1 U1027 ( .A(n1321), .ZN(n1320) );
NAND3_X1 U1028 ( .A1(n1221), .A2(n1321), .A3(KEYINPUT60), .ZN(n1318) );
XOR2_X1 U1029 ( .A(n1322), .B(n1323), .Z(n1221) );
NOR2_X1 U1030 ( .A1(KEYINPUT15), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1031 ( .A1(n1325), .A2(KEYINPUT59), .ZN(n1316) );
XOR2_X1 U1032 ( .A(n1169), .B(KEYINPUT29), .Z(n1325) );
XOR2_X1 U1033 ( .A(n1326), .B(n1327), .Z(n1169) );
XOR2_X1 U1034 ( .A(G119), .B(G113), .Z(n1327) );
NAND2_X1 U1035 ( .A1(KEYINPUT61), .A2(n1263), .ZN(n1326) );
NAND3_X1 U1036 ( .A1(n1328), .A2(n1078), .A3(G210), .ZN(n1163) );
XOR2_X1 U1037 ( .A(KEYINPUT37), .B(G237), .Z(n1328) );
AND3_X1 U1038 ( .A1(n1071), .A2(n1212), .A3(n1083), .ZN(n1250) );
INV_X1 U1039 ( .A(n1069), .ZN(n1083) );
NAND2_X1 U1040 ( .A1(n1088), .A2(n1237), .ZN(n1069) );
XOR2_X1 U1041 ( .A(n1329), .B(n1100), .Z(n1237) );
NAND2_X1 U1042 ( .A1(n1330), .A2(n1274), .ZN(n1100) );
XOR2_X1 U1043 ( .A(KEYINPUT46), .B(n1154), .Z(n1330) );
XNOR2_X1 U1044 ( .A(n1331), .B(n1332), .ZN(n1154) );
XOR2_X1 U1045 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1046 ( .A(n1335), .B(n1336), .Z(n1334) );
NAND3_X1 U1047 ( .A1(n1295), .A2(n1078), .A3(G214), .ZN(n1336) );
INV_X1 U1048 ( .A(G237), .ZN(n1295) );
NAND2_X1 U1049 ( .A1(n1337), .A2(n1338), .ZN(n1335) );
NAND2_X1 U1050 ( .A1(G104), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1051 ( .A(n1340), .B(KEYINPUT16), .Z(n1337) );
OR2_X1 U1052 ( .A1(n1339), .A2(G104), .ZN(n1340) );
XOR2_X1 U1053 ( .A(G113), .B(G122), .Z(n1339) );
NOR2_X1 U1054 ( .A1(G131), .A2(KEYINPUT25), .ZN(n1333) );
XOR2_X1 U1055 ( .A(n1303), .B(n1341), .Z(n1331) );
XOR2_X1 U1056 ( .A(n1226), .B(n1181), .Z(n1303) );
INV_X1 U1057 ( .A(G125), .ZN(n1226) );
NAND2_X1 U1058 ( .A1(KEYINPUT2), .A2(n1099), .ZN(n1329) );
INV_X1 U1059 ( .A(G475), .ZN(n1099) );
XOR2_X1 U1060 ( .A(n1342), .B(G478), .Z(n1088) );
NAND2_X1 U1061 ( .A1(n1149), .A2(n1274), .ZN(n1342) );
XNOR2_X1 U1062 ( .A(n1343), .B(n1344), .ZN(n1149) );
NOR3_X1 U1063 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1344) );
NOR2_X1 U1064 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
AND3_X1 U1065 ( .A1(n1349), .A2(n1350), .A3(n1348), .ZN(n1346) );
NOR2_X1 U1066 ( .A1(KEYINPUT49), .A2(n1351), .ZN(n1348) );
INV_X1 U1067 ( .A(KEYINPUT14), .ZN(n1350) );
XNOR2_X1 U1068 ( .A(n1352), .B(n1353), .ZN(n1349) );
NOR2_X1 U1069 ( .A1(G122), .A2(KEYINPUT38), .ZN(n1353) );
XOR2_X1 U1070 ( .A(G107), .B(n1263), .Z(n1352) );
INV_X1 U1071 ( .A(G116), .ZN(n1263) );
AND2_X1 U1072 ( .A1(n1351), .A2(KEYINPUT14), .ZN(n1345) );
XOR2_X1 U1073 ( .A(G128), .B(n1354), .Z(n1351) );
XOR2_X1 U1074 ( .A(G143), .B(G134), .Z(n1354) );
NAND3_X1 U1075 ( .A1(G217), .A2(n1305), .A3(KEYINPUT1), .ZN(n1343) );
AND2_X1 U1076 ( .A1(G234), .A2(n1078), .ZN(n1305) );
NAND2_X1 U1077 ( .A1(n1355), .A2(n1061), .ZN(n1212) );
NAND3_X1 U1078 ( .A1(n1253), .A2(n1078), .A3(n1356), .ZN(n1061) );
XNOR2_X1 U1079 ( .A(G952), .B(KEYINPUT28), .ZN(n1356) );
NAND3_X1 U1080 ( .A1(n1132), .A2(n1253), .A3(G902), .ZN(n1355) );
NAND2_X1 U1081 ( .A1(G237), .A2(G234), .ZN(n1253) );
NOR2_X1 U1082 ( .A1(n1078), .A2(G898), .ZN(n1132) );
INV_X1 U1083 ( .A(n1247), .ZN(n1071) );
NAND2_X1 U1084 ( .A1(n1074), .A2(n1073), .ZN(n1247) );
NAND2_X1 U1085 ( .A1(G221), .A2(n1297), .ZN(n1073) );
NAND2_X1 U1086 ( .A1(G234), .A2(n1274), .ZN(n1297) );
XNOR2_X1 U1087 ( .A(n1357), .B(G469), .ZN(n1074) );
NAND2_X1 U1088 ( .A1(n1358), .A2(n1274), .ZN(n1357) );
INV_X1 U1089 ( .A(G902), .ZN(n1274) );
XOR2_X1 U1090 ( .A(n1180), .B(n1359), .Z(n1358) );
XOR2_X1 U1091 ( .A(G110), .B(n1181), .Z(n1359) );
XOR2_X1 U1092 ( .A(G140), .B(KEYINPUT24), .Z(n1181) );
XNOR2_X1 U1093 ( .A(n1360), .B(n1361), .ZN(n1180) );
XOR2_X1 U1094 ( .A(n1287), .B(n1362), .Z(n1361) );
XOR2_X1 U1095 ( .A(n1112), .B(n1321), .Z(n1362) );
XOR2_X1 U1096 ( .A(n1363), .B(n1110), .Z(n1321) );
XOR2_X1 U1097 ( .A(G137), .B(G134), .Z(n1110) );
NAND2_X1 U1098 ( .A1(KEYINPUT41), .A2(n1111), .ZN(n1363) );
INV_X1 U1099 ( .A(G131), .ZN(n1111) );
NAND2_X1 U1100 ( .A1(n1364), .A2(n1365), .ZN(n1112) );
NAND2_X1 U1101 ( .A1(n1366), .A2(n1322), .ZN(n1365) );
XOR2_X1 U1102 ( .A(n1367), .B(KEYINPUT0), .Z(n1364) );
OR2_X1 U1103 ( .A1(n1366), .A2(n1322), .ZN(n1367) );
XOR2_X1 U1104 ( .A(G128), .B(KEYINPUT58), .Z(n1322) );
INV_X1 U1105 ( .A(n1324), .ZN(n1366) );
XNOR2_X1 U1106 ( .A(n1341), .B(KEYINPUT51), .ZN(n1324) );
XOR2_X1 U1107 ( .A(G146), .B(G143), .Z(n1341) );
XOR2_X1 U1108 ( .A(G107), .B(G104), .Z(n1287) );
XOR2_X1 U1109 ( .A(n1368), .B(n1369), .Z(n1360) );
XOR2_X1 U1110 ( .A(KEYINPUT13), .B(G101), .Z(n1369) );
NAND2_X1 U1111 ( .A1(G227), .A2(n1078), .ZN(n1368) );
INV_X1 U1112 ( .A(G953), .ZN(n1078) );
endmodule


