//Key = 0100100000110011011010010100101111111011111101011001011101010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398;

XOR2_X1 U762 ( .A(n1068), .B(n1069), .Z(G9) );
NOR2_X1 U763 ( .A1(n1070), .A2(n1071), .ZN(G75) );
NOR4_X1 U764 ( .A1(G953), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1071) );
NOR2_X1 U765 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
INV_X1 U766 ( .A(n1077), .ZN(n1076) );
NOR2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
NOR3_X1 U768 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR3_X1 U769 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1081) );
NOR2_X1 U770 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U771 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U772 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
XOR2_X1 U773 ( .A(n1092), .B(KEYINPUT3), .Z(n1091) );
NOR3_X1 U774 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1083) );
XOR2_X1 U775 ( .A(n1096), .B(KEYINPUT24), .Z(n1095) );
NOR3_X1 U776 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1078) );
NOR4_X1 U777 ( .A1(n1087), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1098) );
AND2_X1 U778 ( .A1(n1102), .A2(KEYINPUT53), .ZN(n1101) );
NOR2_X1 U779 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
XOR2_X1 U780 ( .A(n1080), .B(KEYINPUT56), .Z(n1103) );
NOR2_X1 U781 ( .A1(n1105), .A2(n1082), .ZN(n1099) );
NOR2_X1 U782 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
AND2_X1 U783 ( .A1(n1108), .A2(KEYINPUT35), .ZN(n1107) );
INV_X1 U784 ( .A(n1109), .ZN(n1087) );
NOR3_X1 U785 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1097) );
NOR2_X1 U786 ( .A1(KEYINPUT53), .A2(n1112), .ZN(n1111) );
NOR3_X1 U787 ( .A1(n1113), .A2(KEYINPUT35), .A3(n1082), .ZN(n1110) );
NOR3_X1 U788 ( .A1(n1072), .A2(G953), .A3(G952), .ZN(n1070) );
AND4_X1 U789 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1072) );
NOR4_X1 U790 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1117) );
XOR2_X1 U791 ( .A(KEYINPUT22), .B(n1122), .Z(n1121) );
NOR2_X1 U792 ( .A1(G478), .A2(n1123), .ZN(n1122) );
XOR2_X1 U793 ( .A(n1124), .B(n1125), .Z(n1120) );
NOR2_X1 U794 ( .A1(KEYINPUT27), .A2(n1126), .ZN(n1125) );
XOR2_X1 U795 ( .A(KEYINPUT30), .B(n1127), .Z(n1119) );
NOR2_X1 U796 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U797 ( .A(KEYINPUT0), .B(n1130), .Z(n1129) );
XOR2_X1 U798 ( .A(n1131), .B(n1132), .Z(n1118) );
XOR2_X1 U799 ( .A(n1133), .B(KEYINPUT55), .Z(n1132) );
NAND2_X1 U800 ( .A1(KEYINPUT4), .A2(n1134), .ZN(n1131) );
NOR3_X1 U801 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1116) );
NOR2_X1 U802 ( .A1(n1138), .A2(n1139), .ZN(n1136) );
XOR2_X1 U803 ( .A(n1092), .B(KEYINPUT33), .Z(n1135) );
XOR2_X1 U804 ( .A(n1140), .B(n1141), .Z(G72) );
XOR2_X1 U805 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U806 ( .A1(G953), .A2(n1144), .ZN(n1143) );
NOR2_X1 U807 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U808 ( .A(KEYINPUT19), .B(n1147), .Z(n1146) );
NAND2_X1 U809 ( .A1(n1148), .A2(n1149), .ZN(n1142) );
NAND2_X1 U810 ( .A1(G953), .A2(n1150), .ZN(n1149) );
XOR2_X1 U811 ( .A(n1151), .B(n1152), .Z(n1148) );
XOR2_X1 U812 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U813 ( .A1(n1155), .A2(KEYINPUT17), .ZN(n1153) );
XOR2_X1 U814 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U815 ( .A1(KEYINPUT18), .A2(G131), .ZN(n1156) );
XOR2_X1 U816 ( .A(n1158), .B(G140), .Z(n1151) );
NAND2_X1 U817 ( .A1(G953), .A2(n1159), .ZN(n1140) );
NAND2_X1 U818 ( .A1(G900), .A2(G227), .ZN(n1159) );
XOR2_X1 U819 ( .A(n1160), .B(n1161), .Z(G69) );
NOR2_X1 U820 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U821 ( .A(KEYINPUT46), .B(n1164), .Z(n1163) );
AND2_X1 U822 ( .A1(G224), .A2(G898), .ZN(n1164) );
NAND2_X1 U823 ( .A1(n1165), .A2(n1166), .ZN(n1160) );
NAND2_X1 U824 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U825 ( .A(KEYINPUT52), .B(n1169), .Z(n1167) );
NOR2_X1 U826 ( .A1(G953), .A2(n1170), .ZN(n1169) );
OR3_X1 U827 ( .A1(n1171), .A2(n1172), .A3(n1168), .ZN(n1165) );
NOR2_X1 U828 ( .A1(n1173), .A2(n1174), .ZN(G66) );
NOR3_X1 U829 ( .A1(n1124), .A2(n1175), .A3(n1176), .ZN(n1174) );
NOR3_X1 U830 ( .A1(n1177), .A2(n1126), .A3(n1178), .ZN(n1176) );
NOR2_X1 U831 ( .A1(n1179), .A2(n1180), .ZN(n1175) );
NOR2_X1 U832 ( .A1(n1181), .A2(n1126), .ZN(n1179) );
NOR2_X1 U833 ( .A1(n1173), .A2(n1182), .ZN(G63) );
NOR3_X1 U834 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
NOR2_X1 U835 ( .A1(KEYINPUT41), .A2(n1186), .ZN(n1185) );
NOR2_X1 U836 ( .A1(n1187), .A2(n1188), .ZN(n1184) );
NOR2_X1 U837 ( .A1(n1189), .A2(n1138), .ZN(n1187) );
NOR2_X1 U838 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U839 ( .A1(n1181), .A2(n1139), .ZN(n1190) );
NOR3_X1 U840 ( .A1(n1178), .A2(n1192), .A3(n1139), .ZN(n1183) );
INV_X1 U841 ( .A(G478), .ZN(n1139) );
NOR2_X1 U842 ( .A1(n1191), .A2(n1188), .ZN(n1192) );
INV_X1 U843 ( .A(KEYINPUT41), .ZN(n1188) );
NOR2_X1 U844 ( .A1(n1173), .A2(n1193), .ZN(G60) );
XNOR2_X1 U845 ( .A(n1194), .B(n1195), .ZN(n1193) );
AND2_X1 U846 ( .A1(G475), .A2(n1196), .ZN(n1194) );
XOR2_X1 U847 ( .A(n1197), .B(n1198), .Z(G6) );
NOR2_X1 U848 ( .A1(n1173), .A2(n1199), .ZN(G57) );
XOR2_X1 U849 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U850 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
AND3_X1 U851 ( .A1(n1204), .A2(G472), .A3(n1196), .ZN(n1203) );
NOR2_X1 U852 ( .A1(n1205), .A2(n1204), .ZN(n1202) );
NAND2_X1 U853 ( .A1(n1206), .A2(n1207), .ZN(n1204) );
NAND3_X1 U854 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
INV_X1 U855 ( .A(KEYINPUT11), .ZN(n1210) );
NAND2_X1 U856 ( .A1(n1211), .A2(KEYINPUT11), .ZN(n1206) );
XOR2_X1 U857 ( .A(KEYINPUT9), .B(n1212), .Z(n1205) );
NOR2_X1 U858 ( .A1(n1134), .A2(n1178), .ZN(n1212) );
INV_X1 U859 ( .A(G472), .ZN(n1134) );
NOR2_X1 U860 ( .A1(n1173), .A2(n1213), .ZN(G54) );
XOR2_X1 U861 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U862 ( .A(n1216), .B(n1217), .Z(n1214) );
AND2_X1 U863 ( .A1(G469), .A2(n1196), .ZN(n1217) );
NAND3_X1 U864 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1216) );
NAND2_X1 U865 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
OR3_X1 U866 ( .A1(n1222), .A2(n1221), .A3(n1223), .ZN(n1219) );
INV_X1 U867 ( .A(KEYINPUT57), .ZN(n1222) );
NAND2_X1 U868 ( .A1(n1224), .A2(n1223), .ZN(n1218) );
NAND3_X1 U869 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1223) );
NAND2_X1 U870 ( .A1(KEYINPUT29), .A2(n1228), .ZN(n1227) );
OR3_X1 U871 ( .A1(n1229), .A2(KEYINPUT29), .A3(n1230), .ZN(n1226) );
NAND2_X1 U872 ( .A1(n1230), .A2(n1229), .ZN(n1225) );
NAND2_X1 U873 ( .A1(KEYINPUT51), .A2(n1154), .ZN(n1229) );
INV_X1 U874 ( .A(n1228), .ZN(n1154) );
NAND2_X1 U875 ( .A1(KEYINPUT57), .A2(n1231), .ZN(n1224) );
XOR2_X1 U876 ( .A(KEYINPUT34), .B(n1221), .Z(n1231) );
NOR2_X1 U877 ( .A1(n1173), .A2(n1232), .ZN(G51) );
XOR2_X1 U878 ( .A(n1233), .B(n1234), .Z(n1232) );
NOR2_X1 U879 ( .A1(KEYINPUT12), .A2(n1235), .ZN(n1234) );
XOR2_X1 U880 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U881 ( .A(n1170), .B(n1238), .Z(n1237) );
XOR2_X1 U882 ( .A(n1158), .B(n1239), .Z(n1236) );
NOR2_X1 U883 ( .A1(KEYINPUT7), .A2(n1240), .ZN(n1239) );
NAND3_X1 U884 ( .A1(n1196), .A2(G210), .A3(KEYINPUT45), .ZN(n1233) );
INV_X1 U885 ( .A(n1178), .ZN(n1196) );
NAND2_X1 U886 ( .A1(G902), .A2(n1074), .ZN(n1178) );
INV_X1 U887 ( .A(n1181), .ZN(n1074) );
NOR3_X1 U888 ( .A1(n1168), .A2(n1147), .A3(n1145), .ZN(n1181) );
NAND4_X1 U889 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1145) );
NOR4_X1 U890 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1244) );
NAND3_X1 U891 ( .A1(n1249), .A2(n1108), .A3(n1250), .ZN(n1243) );
XOR2_X1 U892 ( .A(n1251), .B(KEYINPUT15), .Z(n1250) );
NAND4_X1 U893 ( .A1(n1252), .A2(n1198), .A3(n1253), .A4(n1254), .ZN(n1168) );
NOR4_X1 U894 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
INV_X1 U895 ( .A(n1069), .ZN(n1258) );
NAND3_X1 U896 ( .A1(n1259), .A2(n1260), .A3(n1106), .ZN(n1069) );
NOR3_X1 U897 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1253) );
NOR2_X1 U898 ( .A1(KEYINPUT16), .A2(n1264), .ZN(n1263) );
AND4_X1 U899 ( .A1(KEYINPUT16), .A2(n1265), .A3(n1251), .A4(n1266), .ZN(n1262) );
NOR2_X1 U900 ( .A1(n1251), .A2(n1267), .ZN(n1261) );
NAND3_X1 U901 ( .A1(n1259), .A2(n1260), .A3(n1108), .ZN(n1198) );
INV_X1 U902 ( .A(n1082), .ZN(n1260) );
NAND3_X1 U903 ( .A1(n1268), .A2(n1259), .A3(n1269), .ZN(n1252) );
NOR2_X1 U904 ( .A1(n1162), .A2(G952), .ZN(n1173) );
XOR2_X1 U905 ( .A(G146), .B(n1270), .Z(G48) );
NOR3_X1 U906 ( .A1(n1271), .A2(n1251), .A3(n1113), .ZN(n1270) );
NAND2_X1 U907 ( .A1(n1272), .A2(n1273), .ZN(G45) );
OR2_X1 U908 ( .A1(n1274), .A2(G143), .ZN(n1273) );
NAND2_X1 U909 ( .A1(n1275), .A2(G143), .ZN(n1272) );
NAND2_X1 U910 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U911 ( .A1(n1248), .A2(n1278), .ZN(n1277) );
INV_X1 U912 ( .A(KEYINPUT36), .ZN(n1278) );
NAND2_X1 U913 ( .A1(KEYINPUT36), .A2(n1274), .ZN(n1276) );
NAND2_X1 U914 ( .A1(KEYINPUT43), .A2(n1248), .ZN(n1274) );
AND4_X1 U915 ( .A1(n1279), .A2(n1280), .A3(n1281), .A4(n1282), .ZN(n1248) );
XOR2_X1 U916 ( .A(n1241), .B(n1283), .Z(G42) );
XOR2_X1 U917 ( .A(KEYINPUT40), .B(G140), .Z(n1283) );
NAND4_X1 U918 ( .A1(n1284), .A2(n1109), .A3(n1285), .A4(n1108), .ZN(n1241) );
XOR2_X1 U919 ( .A(n1286), .B(n1242), .Z(G39) );
NAND3_X1 U920 ( .A1(n1249), .A2(n1109), .A3(n1269), .ZN(n1242) );
XOR2_X1 U921 ( .A(G134), .B(n1247), .Z(G36) );
AND3_X1 U922 ( .A1(n1279), .A2(n1106), .A3(n1109), .ZN(n1247) );
XOR2_X1 U923 ( .A(G131), .B(n1147), .Z(G33) );
AND3_X1 U924 ( .A1(n1279), .A2(n1108), .A3(n1109), .ZN(n1147) );
NOR2_X1 U925 ( .A1(n1094), .A2(n1137), .ZN(n1109) );
INV_X1 U926 ( .A(n1093), .ZN(n1137) );
AND3_X1 U927 ( .A1(n1089), .A2(n1287), .A3(n1268), .ZN(n1279) );
XOR2_X1 U928 ( .A(G128), .B(n1246), .Z(G30) );
AND3_X1 U929 ( .A1(n1106), .A2(n1280), .A3(n1249), .ZN(n1246) );
INV_X1 U930 ( .A(n1271), .ZN(n1249) );
NAND2_X1 U931 ( .A1(n1284), .A2(n1288), .ZN(n1271) );
AND3_X1 U932 ( .A1(n1289), .A2(n1287), .A3(n1089), .ZN(n1284) );
XNOR2_X1 U933 ( .A(G101), .B(n1290), .ZN(G3) );
NAND3_X1 U934 ( .A1(n1259), .A2(n1291), .A3(n1268), .ZN(n1290) );
XOR2_X1 U935 ( .A(KEYINPUT60), .B(n1269), .Z(n1291) );
XOR2_X1 U936 ( .A(n1245), .B(n1292), .Z(G27) );
NOR2_X1 U937 ( .A1(KEYINPUT26), .A2(n1158), .ZN(n1292) );
AND3_X1 U938 ( .A1(n1084), .A2(n1108), .A3(n1293), .ZN(n1245) );
AND3_X1 U939 ( .A1(n1285), .A2(n1287), .A3(n1289), .ZN(n1293) );
NAND2_X1 U940 ( .A1(n1294), .A2(n1295), .ZN(n1287) );
NAND4_X1 U941 ( .A1(G902), .A2(G953), .A3(n1077), .A4(n1150), .ZN(n1295) );
INV_X1 U942 ( .A(G900), .ZN(n1150) );
XOR2_X1 U943 ( .A(n1296), .B(n1264), .Z(G24) );
NAND2_X1 U944 ( .A1(n1265), .A2(n1084), .ZN(n1264) );
NOR4_X1 U945 ( .A1(n1082), .A2(n1297), .A3(n1298), .A4(n1299), .ZN(n1265) );
NAND2_X1 U946 ( .A1(n1285), .A2(n1300), .ZN(n1082) );
XOR2_X1 U947 ( .A(G119), .B(n1257), .Z(G21) );
AND3_X1 U948 ( .A1(n1269), .A2(n1084), .A3(n1301), .ZN(n1257) );
NOR3_X1 U949 ( .A1(n1285), .A2(n1298), .A3(n1302), .ZN(n1301) );
INV_X1 U950 ( .A(n1303), .ZN(n1298) );
XOR2_X1 U951 ( .A(n1256), .B(n1304), .Z(G18) );
NOR2_X1 U952 ( .A1(KEYINPUT2), .A2(n1305), .ZN(n1304) );
INV_X1 U953 ( .A(G116), .ZN(n1305) );
AND4_X1 U954 ( .A1(n1084), .A2(n1268), .A3(n1106), .A4(n1303), .ZN(n1256) );
NOR2_X1 U955 ( .A1(n1282), .A2(n1297), .ZN(n1106) );
NOR2_X1 U956 ( .A1(n1096), .A2(n1251), .ZN(n1084) );
INV_X1 U957 ( .A(n1266), .ZN(n1096) );
XOR2_X1 U958 ( .A(G113), .B(n1306), .Z(G15) );
NOR2_X1 U959 ( .A1(n1307), .A2(n1251), .ZN(n1306) );
XOR2_X1 U960 ( .A(n1267), .B(KEYINPUT5), .Z(n1307) );
NAND4_X1 U961 ( .A1(n1266), .A2(n1108), .A3(n1268), .A4(n1303), .ZN(n1267) );
INV_X1 U962 ( .A(n1104), .ZN(n1268) );
NAND2_X1 U963 ( .A1(n1288), .A2(n1300), .ZN(n1104) );
XOR2_X1 U964 ( .A(n1289), .B(KEYINPUT61), .Z(n1300) );
INV_X1 U965 ( .A(n1285), .ZN(n1288) );
INV_X1 U966 ( .A(n1113), .ZN(n1108) );
NAND2_X1 U967 ( .A1(n1308), .A2(n1282), .ZN(n1113) );
INV_X1 U968 ( .A(n1299), .ZN(n1282) );
XOR2_X1 U969 ( .A(n1281), .B(KEYINPUT14), .Z(n1308) );
NOR2_X1 U970 ( .A1(n1309), .A2(n1090), .ZN(n1266) );
XNOR2_X1 U971 ( .A(n1092), .B(KEYINPUT21), .ZN(n1309) );
XOR2_X1 U972 ( .A(n1310), .B(n1255), .Z(G12) );
AND2_X1 U973 ( .A1(n1102), .A2(n1259), .ZN(n1255) );
AND3_X1 U974 ( .A1(n1280), .A2(n1303), .A3(n1089), .ZN(n1259) );
AND2_X1 U975 ( .A1(n1090), .A2(n1092), .ZN(n1089) );
NAND2_X1 U976 ( .A1(G221), .A2(n1311), .ZN(n1092) );
XOR2_X1 U977 ( .A(n1114), .B(KEYINPUT63), .Z(n1090) );
XOR2_X1 U978 ( .A(n1312), .B(G469), .Z(n1114) );
NAND2_X1 U979 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U980 ( .A(n1315), .B(n1316), .Z(n1313) );
XOR2_X1 U981 ( .A(n1228), .B(n1215), .Z(n1316) );
XNOR2_X1 U982 ( .A(n1317), .B(n1318), .ZN(n1215) );
XOR2_X1 U983 ( .A(G140), .B(G110), .Z(n1318) );
NAND2_X1 U984 ( .A1(G227), .A2(n1162), .ZN(n1317) );
XNOR2_X1 U985 ( .A(n1319), .B(n1320), .ZN(n1228) );
NOR2_X1 U986 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NOR3_X1 U987 ( .A1(G146), .A2(KEYINPUT44), .A3(n1323), .ZN(n1322) );
NOR2_X1 U988 ( .A1(n1324), .A2(n1325), .ZN(n1321) );
NOR2_X1 U989 ( .A1(n1326), .A2(n1327), .ZN(n1324) );
INV_X1 U990 ( .A(G143), .ZN(n1327) );
NOR2_X1 U991 ( .A1(n1323), .A2(n1328), .ZN(n1326) );
INV_X1 U992 ( .A(KEYINPUT44), .ZN(n1328) );
XOR2_X1 U993 ( .A(G143), .B(KEYINPUT59), .Z(n1323) );
XNOR2_X1 U994 ( .A(n1221), .B(n1230), .ZN(n1315) );
AND2_X1 U995 ( .A1(n1329), .A2(n1330), .ZN(n1230) );
NAND3_X1 U996 ( .A1(n1331), .A2(n1332), .A3(G101), .ZN(n1330) );
XOR2_X1 U997 ( .A(KEYINPUT28), .B(n1333), .Z(n1329) );
NOR2_X1 U998 ( .A1(G101), .A2(n1334), .ZN(n1333) );
AND2_X1 U999 ( .A1(n1331), .A2(n1332), .ZN(n1334) );
NAND2_X1 U1000 ( .A1(n1335), .A2(G107), .ZN(n1332) );
XOR2_X1 U1001 ( .A(n1197), .B(KEYINPUT38), .Z(n1335) );
NAND2_X1 U1002 ( .A1(n1068), .A2(n1197), .ZN(n1331) );
INV_X1 U1003 ( .A(G104), .ZN(n1197) );
NAND2_X1 U1004 ( .A1(n1294), .A2(n1336), .ZN(n1303) );
NAND3_X1 U1005 ( .A1(n1172), .A2(n1077), .A3(G902), .ZN(n1336) );
NOR2_X1 U1006 ( .A1(n1162), .A2(G898), .ZN(n1172) );
NAND3_X1 U1007 ( .A1(n1077), .A2(n1162), .A3(n1337), .ZN(n1294) );
XNOR2_X1 U1008 ( .A(G952), .B(KEYINPUT25), .ZN(n1337) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1077) );
INV_X1 U1010 ( .A(n1251), .ZN(n1280) );
NAND2_X1 U1011 ( .A1(n1094), .A2(n1093), .ZN(n1251) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1338), .ZN(n1093) );
XOR2_X1 U1013 ( .A(n1115), .B(KEYINPUT42), .Z(n1094) );
XOR2_X1 U1014 ( .A(n1339), .B(n1340), .Z(n1115) );
AND2_X1 U1015 ( .A1(n1338), .A2(G210), .ZN(n1340) );
OR2_X1 U1016 ( .A1(G902), .A2(G237), .ZN(n1338) );
NAND4_X1 U1017 ( .A1(n1341), .A2(n1314), .A3(n1342), .A4(n1343), .ZN(n1339) );
OR3_X1 U1018 ( .A1(n1170), .A2(KEYINPUT50), .A3(n1344), .ZN(n1343) );
NAND2_X1 U1019 ( .A1(n1344), .A2(n1345), .ZN(n1342) );
NAND2_X1 U1020 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
INV_X1 U1021 ( .A(KEYINPUT50), .ZN(n1347) );
XOR2_X1 U1022 ( .A(KEYINPUT58), .B(n1171), .Z(n1346) );
INV_X1 U1023 ( .A(n1170), .ZN(n1171) );
XOR2_X1 U1024 ( .A(n1348), .B(n1238), .Z(n1344) );
XNOR2_X1 U1025 ( .A(n1349), .B(n1240), .ZN(n1348) );
NAND2_X1 U1026 ( .A1(G224), .A2(n1162), .ZN(n1240) );
NAND2_X1 U1027 ( .A1(KEYINPUT23), .A2(n1158), .ZN(n1349) );
NAND2_X1 U1028 ( .A1(KEYINPUT50), .A2(n1170), .ZN(n1341) );
XOR2_X1 U1029 ( .A(n1350), .B(n1351), .Z(n1170) );
XOR2_X1 U1030 ( .A(G101), .B(n1352), .Z(n1351) );
XOR2_X1 U1031 ( .A(G110), .B(G104), .Z(n1352) );
XOR2_X1 U1032 ( .A(n1353), .B(n1354), .Z(n1350) );
XOR2_X1 U1033 ( .A(n1355), .B(n1356), .Z(n1353) );
INV_X1 U1034 ( .A(n1357), .ZN(n1356) );
NAND2_X1 U1035 ( .A1(KEYINPUT47), .A2(n1068), .ZN(n1355) );
INV_X1 U1036 ( .A(G107), .ZN(n1068) );
INV_X1 U1037 ( .A(n1112), .ZN(n1102) );
NAND3_X1 U1038 ( .A1(n1285), .A2(n1289), .A3(n1269), .ZN(n1112) );
INV_X1 U1039 ( .A(n1080), .ZN(n1269) );
NAND2_X1 U1040 ( .A1(n1297), .A2(n1299), .ZN(n1080) );
NOR2_X1 U1041 ( .A1(n1128), .A2(n1130), .ZN(n1299) );
AND3_X1 U1042 ( .A1(n1358), .A2(n1314), .A3(n1195), .ZN(n1130) );
NOR2_X1 U1043 ( .A1(n1358), .A2(n1359), .ZN(n1128) );
AND2_X1 U1044 ( .A1(n1195), .A2(n1314), .ZN(n1359) );
XOR2_X1 U1045 ( .A(n1360), .B(n1361), .Z(n1195) );
XOR2_X1 U1046 ( .A(n1362), .B(n1363), .Z(n1361) );
XOR2_X1 U1047 ( .A(G131), .B(G104), .Z(n1363) );
XOR2_X1 U1048 ( .A(G143), .B(G140), .Z(n1362) );
XOR2_X1 U1049 ( .A(n1364), .B(n1354), .Z(n1360) );
XNOR2_X1 U1050 ( .A(G113), .B(n1296), .ZN(n1354) );
INV_X1 U1051 ( .A(G122), .ZN(n1296) );
XOR2_X1 U1052 ( .A(n1365), .B(n1366), .Z(n1364) );
AND2_X1 U1053 ( .A1(n1367), .A2(G214), .ZN(n1366) );
XOR2_X1 U1054 ( .A(G475), .B(KEYINPUT54), .Z(n1358) );
INV_X1 U1055 ( .A(n1281), .ZN(n1297) );
NAND3_X1 U1056 ( .A1(n1368), .A2(n1369), .A3(n1370), .ZN(n1281) );
OR2_X1 U1057 ( .A1(n1371), .A2(KEYINPUT10), .ZN(n1370) );
NAND3_X1 U1058 ( .A1(KEYINPUT10), .A2(n1371), .A3(n1138), .ZN(n1369) );
INV_X1 U1059 ( .A(n1123), .ZN(n1138) );
NAND2_X1 U1060 ( .A1(n1372), .A2(n1123), .ZN(n1368) );
NAND2_X1 U1061 ( .A1(n1186), .A2(n1314), .ZN(n1123) );
INV_X1 U1062 ( .A(n1191), .ZN(n1186) );
XOR2_X1 U1063 ( .A(n1373), .B(n1374), .Z(n1191) );
XOR2_X1 U1064 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1065 ( .A(G122), .B(G107), .Z(n1376) );
XOR2_X1 U1066 ( .A(G143), .B(G134), .Z(n1375) );
XOR2_X1 U1067 ( .A(n1377), .B(n1378), .Z(n1373) );
XOR2_X1 U1068 ( .A(n1379), .B(n1380), .Z(n1377) );
AND3_X1 U1069 ( .A1(G234), .A2(n1162), .A3(G217), .ZN(n1380) );
NAND2_X1 U1070 ( .A1(KEYINPUT31), .A2(n1319), .ZN(n1379) );
NAND2_X1 U1071 ( .A1(KEYINPUT10), .A2(n1381), .ZN(n1372) );
XOR2_X1 U1072 ( .A(KEYINPUT49), .B(n1371), .Z(n1381) );
XOR2_X1 U1073 ( .A(G478), .B(KEYINPUT32), .Z(n1371) );
INV_X1 U1074 ( .A(n1302), .ZN(n1289) );
XOR2_X1 U1075 ( .A(n1124), .B(n1126), .Z(n1302) );
NAND2_X1 U1076 ( .A1(G217), .A2(n1311), .ZN(n1126) );
NAND2_X1 U1077 ( .A1(G234), .A2(n1314), .ZN(n1311) );
NOR2_X1 U1078 ( .A1(n1180), .A2(G902), .ZN(n1124) );
INV_X1 U1079 ( .A(n1177), .ZN(n1180) );
XOR2_X1 U1080 ( .A(n1382), .B(n1383), .Z(n1177) );
XOR2_X1 U1081 ( .A(n1384), .B(n1385), .Z(n1383) );
XNOR2_X1 U1082 ( .A(n1386), .B(n1387), .ZN(n1385) );
NOR2_X1 U1083 ( .A1(KEYINPUT37), .A2(n1388), .ZN(n1387) );
XNOR2_X1 U1084 ( .A(n1319), .B(n1389), .ZN(n1388) );
XOR2_X1 U1085 ( .A(G110), .B(n1390), .Z(n1389) );
NOR2_X1 U1086 ( .A1(G119), .A2(KEYINPUT6), .ZN(n1390) );
NOR2_X1 U1087 ( .A1(KEYINPUT13), .A2(n1391), .ZN(n1386) );
XOR2_X1 U1088 ( .A(KEYINPUT8), .B(G140), .Z(n1391) );
NAND3_X1 U1089 ( .A1(G234), .A2(n1162), .A3(G221), .ZN(n1384) );
INV_X1 U1090 ( .A(G953), .ZN(n1162) );
XOR2_X1 U1091 ( .A(n1392), .B(n1393), .Z(n1382) );
INV_X1 U1092 ( .A(n1365), .ZN(n1393) );
XOR2_X1 U1093 ( .A(n1158), .B(n1394), .Z(n1365) );
XOR2_X1 U1094 ( .A(KEYINPUT48), .B(G146), .Z(n1394) );
INV_X1 U1095 ( .A(G125), .ZN(n1158) );
NAND2_X1 U1096 ( .A1(KEYINPUT1), .A2(n1286), .ZN(n1392) );
XOR2_X1 U1097 ( .A(n1133), .B(G472), .Z(n1285) );
NAND2_X1 U1098 ( .A1(n1395), .A2(n1314), .ZN(n1133) );
INV_X1 U1099 ( .A(G902), .ZN(n1314) );
XOR2_X1 U1100 ( .A(n1396), .B(n1211), .Z(n1395) );
XOR2_X1 U1101 ( .A(n1209), .B(n1208), .Z(n1211) );
XOR2_X1 U1102 ( .A(n1221), .B(n1238), .Z(n1208) );
XNOR2_X1 U1103 ( .A(n1397), .B(n1319), .ZN(n1238) );
XOR2_X1 U1104 ( .A(G128), .B(KEYINPUT20), .Z(n1319) );
XOR2_X1 U1105 ( .A(n1325), .B(G143), .Z(n1397) );
INV_X1 U1106 ( .A(G146), .ZN(n1325) );
XOR2_X1 U1107 ( .A(G131), .B(n1157), .Z(n1221) );
XNOR2_X1 U1108 ( .A(G134), .B(n1286), .ZN(n1157) );
INV_X1 U1109 ( .A(G137), .ZN(n1286) );
XNOR2_X1 U1110 ( .A(n1357), .B(G113), .ZN(n1209) );
XNOR2_X1 U1111 ( .A(G119), .B(n1378), .ZN(n1357) );
XOR2_X1 U1112 ( .A(G116), .B(KEYINPUT39), .Z(n1378) );
INV_X1 U1113 ( .A(n1200), .ZN(n1396) );
XOR2_X1 U1114 ( .A(n1398), .B(G101), .Z(n1200) );
NAND2_X1 U1115 ( .A1(G210), .A2(n1367), .ZN(n1398) );
NOR2_X1 U1116 ( .A1(G953), .A2(G237), .ZN(n1367) );
XNOR2_X1 U1117 ( .A(G110), .B(KEYINPUT62), .ZN(n1310) );
endmodule


