//Key = 0001100000110110100011111100001011101010000100110101001010100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427, n1428, n1429, n1430;

XNOR2_X1 U782 ( .A(n1086), .B(n1087), .ZN(G9) );
NAND2_X1 U783 ( .A1(KEYINPUT13), .A2(n1088), .ZN(n1086) );
NAND3_X1 U784 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(G75) );
NOR4_X1 U786 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
XOR2_X1 U787 ( .A(n1098), .B(KEYINPUT53), .Z(n1097) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND3_X1 U789 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND3_X1 U793 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NAND2_X1 U794 ( .A1(n1090), .A2(n1113), .ZN(n1108) );
NAND2_X1 U795 ( .A1(n1114), .A2(n1115), .ZN(n1104) );
NAND2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(n1099) );
AND2_X1 U797 ( .A1(n1089), .A2(n1116), .ZN(n1096) );
NOR3_X1 U798 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1116) );
INV_X1 U799 ( .A(n1121), .ZN(n1095) );
NAND3_X1 U800 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1094) );
NAND3_X1 U801 ( .A1(n1101), .A2(n1125), .A3(n1103), .ZN(n1124) );
NAND2_X1 U802 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
OR4_X1 U803 ( .A1(n1128), .A2(n1129), .A3(n1118), .A4(KEYINPUT1), .ZN(n1127) );
NAND2_X1 U804 ( .A1(n1106), .A2(n1130), .ZN(n1126) );
NAND2_X1 U805 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND3_X1 U806 ( .A1(n1110), .A2(n1133), .A3(n1134), .ZN(n1132) );
NAND2_X1 U807 ( .A1(n1090), .A2(n1135), .ZN(n1131) );
NAND2_X1 U808 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U809 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XNOR2_X1 U810 ( .A(n1140), .B(KEYINPUT27), .ZN(n1138) );
NAND2_X1 U811 ( .A1(KEYINPUT1), .A2(n1110), .ZN(n1136) );
NOR3_X1 U812 ( .A1(n1141), .A2(G953), .A3(G952), .ZN(n1092) );
INV_X1 U813 ( .A(n1122), .ZN(n1141) );
NAND4_X1 U814 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1122) );
NOR3_X1 U815 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1145) );
XNOR2_X1 U816 ( .A(n1140), .B(KEYINPUT47), .ZN(n1148) );
XOR2_X1 U817 ( .A(n1149), .B(n1150), .Z(n1147) );
NAND2_X1 U818 ( .A1(KEYINPUT49), .A2(n1151), .ZN(n1149) );
NAND3_X1 U819 ( .A1(n1129), .A2(n1152), .A3(n1153), .ZN(n1146) );
XOR2_X1 U820 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U821 ( .A1(KEYINPUT10), .A2(n1156), .ZN(n1155) );
NOR3_X1 U822 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1144) );
NOR2_X1 U823 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
INV_X1 U824 ( .A(KEYINPUT41), .ZN(n1161) );
NOR2_X1 U825 ( .A1(G472), .A2(n1162), .ZN(n1160) );
NOR3_X1 U826 ( .A1(KEYINPUT41), .A2(G472), .A3(n1163), .ZN(n1158) );
XNOR2_X1 U827 ( .A(G475), .B(n1164), .ZN(n1157) );
NAND2_X1 U828 ( .A1(n1163), .A2(G472), .ZN(n1143) );
NOR2_X1 U829 ( .A1(n1165), .A2(KEYINPUT5), .ZN(n1163) );
INV_X1 U830 ( .A(n1133), .ZN(n1142) );
XOR2_X1 U831 ( .A(n1166), .B(n1167), .Z(G72) );
NOR2_X1 U832 ( .A1(n1168), .A2(n1123), .ZN(n1167) );
AND2_X1 U833 ( .A1(G227), .A2(G900), .ZN(n1168) );
NAND2_X1 U834 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
NAND2_X1 U835 ( .A1(n1171), .A2(n1123), .ZN(n1170) );
XOR2_X1 U836 ( .A(n1172), .B(n1173), .Z(n1171) );
NAND3_X1 U837 ( .A1(G900), .A2(n1173), .A3(G953), .ZN(n1169) );
XOR2_X1 U838 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U839 ( .A1(G125), .A2(KEYINPUT6), .ZN(n1175) );
XOR2_X1 U840 ( .A(n1176), .B(G140), .Z(n1174) );
NAND2_X1 U841 ( .A1(KEYINPUT36), .A2(n1177), .ZN(n1176) );
XOR2_X1 U842 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U843 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U844 ( .A1(KEYINPUT51), .A2(n1182), .ZN(n1181) );
XOR2_X1 U845 ( .A(KEYINPUT54), .B(G131), .Z(n1178) );
XOR2_X1 U846 ( .A(n1183), .B(n1184), .Z(G69) );
XOR2_X1 U847 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND2_X1 U848 ( .A1(G953), .A2(n1187), .ZN(n1186) );
NAND2_X1 U849 ( .A1(G898), .A2(G224), .ZN(n1187) );
NAND4_X1 U850 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1185) );
NAND2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
INV_X1 U852 ( .A(KEYINPUT4), .ZN(n1193) );
XNOR2_X1 U853 ( .A(n1194), .B(n1195), .ZN(n1192) );
AND2_X1 U854 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U855 ( .A1(KEYINPUT4), .A2(n1198), .ZN(n1190) );
INV_X1 U856 ( .A(n1199), .ZN(n1189) );
NAND2_X1 U857 ( .A1(G953), .A2(n1200), .ZN(n1188) );
AND2_X1 U858 ( .A1(n1201), .A2(n1123), .ZN(n1183) );
NOR2_X1 U859 ( .A1(n1202), .A2(n1203), .ZN(G66) );
NOR2_X1 U860 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XOR2_X1 U861 ( .A(KEYINPUT61), .B(n1206), .Z(n1205) );
NOR2_X1 U862 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
AND2_X1 U863 ( .A1(n1207), .A2(n1208), .ZN(n1204) );
NAND2_X1 U864 ( .A1(n1209), .A2(G217), .ZN(n1208) );
NOR2_X1 U865 ( .A1(n1202), .A2(n1210), .ZN(G63) );
NOR3_X1 U866 ( .A1(n1150), .A2(n1211), .A3(n1212), .ZN(n1210) );
AND3_X1 U867 ( .A1(n1213), .A2(G478), .A3(n1209), .ZN(n1212) );
NOR2_X1 U868 ( .A1(n1214), .A2(n1213), .ZN(n1211) );
NOR2_X1 U869 ( .A1(n1121), .A2(n1151), .ZN(n1214) );
NOR2_X1 U870 ( .A1(n1202), .A2(n1215), .ZN(G60) );
NOR3_X1 U871 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NOR3_X1 U872 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1218) );
NOR2_X1 U873 ( .A1(n1222), .A2(n1223), .ZN(n1217) );
NOR2_X1 U874 ( .A1(n1121), .A2(n1220), .ZN(n1222) );
XNOR2_X1 U875 ( .A(G104), .B(n1224), .ZN(G6) );
NAND4_X1 U876 ( .A1(n1117), .A2(n1090), .A3(n1225), .A4(n1113), .ZN(n1224) );
NOR2_X1 U877 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XNOR2_X1 U878 ( .A(n1115), .B(KEYINPUT55), .ZN(n1227) );
NOR2_X1 U879 ( .A1(n1202), .A2(n1228), .ZN(G57) );
XOR2_X1 U880 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U881 ( .A(n1231), .B(n1232), .Z(n1229) );
AND2_X1 U882 ( .A1(G472), .A2(n1209), .ZN(n1232) );
NAND2_X1 U883 ( .A1(KEYINPUT43), .A2(n1233), .ZN(n1231) );
NOR3_X1 U884 ( .A1(n1202), .A2(n1234), .A3(n1235), .ZN(G54) );
NOR2_X1 U885 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
XOR2_X1 U886 ( .A(n1238), .B(n1239), .Z(n1237) );
NOR2_X1 U887 ( .A1(KEYINPUT50), .A2(n1240), .ZN(n1239) );
NOR2_X1 U888 ( .A1(n1241), .A2(n1242), .ZN(n1234) );
XOR2_X1 U889 ( .A(n1238), .B(n1243), .Z(n1242) );
NOR2_X1 U890 ( .A1(KEYINPUT50), .A2(n1244), .ZN(n1243) );
XOR2_X1 U891 ( .A(n1245), .B(n1246), .Z(n1238) );
XOR2_X1 U892 ( .A(n1247), .B(n1248), .Z(n1246) );
AND2_X1 U893 ( .A1(G469), .A2(n1209), .ZN(n1247) );
NOR2_X1 U894 ( .A1(n1202), .A2(n1249), .ZN(G51) );
XOR2_X1 U895 ( .A(n1250), .B(n1251), .Z(n1249) );
NOR3_X1 U896 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
NOR2_X1 U897 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
INV_X1 U898 ( .A(n1257), .ZN(n1256) );
NOR2_X1 U899 ( .A1(KEYINPUT37), .A2(n1258), .ZN(n1255) );
XOR2_X1 U900 ( .A(n1259), .B(KEYINPUT45), .Z(n1258) );
NOR3_X1 U901 ( .A1(n1257), .A2(KEYINPUT37), .A3(n1259), .ZN(n1253) );
XOR2_X1 U902 ( .A(n1233), .B(n1260), .Z(n1257) );
AND2_X1 U903 ( .A1(n1259), .A2(KEYINPUT37), .ZN(n1252) );
XNOR2_X1 U904 ( .A(n1261), .B(n1262), .ZN(n1250) );
NOR2_X1 U905 ( .A1(n1156), .A2(n1221), .ZN(n1262) );
INV_X1 U906 ( .A(n1209), .ZN(n1221) );
NOR2_X1 U907 ( .A1(n1263), .A2(n1121), .ZN(n1209) );
NOR2_X1 U908 ( .A1(n1201), .A2(n1172), .ZN(n1121) );
NAND4_X1 U909 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1172) );
NOR4_X1 U910 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1267) );
NAND2_X1 U911 ( .A1(n1115), .A2(n1272), .ZN(n1266) );
NAND2_X1 U912 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U913 ( .A1(n1275), .A2(n1110), .ZN(n1274) );
NAND4_X1 U914 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1201) );
NOR4_X1 U915 ( .A1(n1280), .A2(n1281), .A3(n1282), .A4(n1283), .ZN(n1279) );
NOR2_X1 U916 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NOR2_X1 U917 ( .A1(n1286), .A2(n1287), .ZN(n1284) );
AND2_X1 U918 ( .A1(n1090), .A2(n1117), .ZN(n1287) );
NOR2_X1 U919 ( .A1(n1288), .A2(n1289), .ZN(n1286) );
XNOR2_X1 U920 ( .A(n1090), .B(KEYINPUT48), .ZN(n1288) );
NOR2_X1 U921 ( .A1(n1290), .A2(n1291), .ZN(n1282) );
NOR2_X1 U922 ( .A1(n1089), .A2(n1117), .ZN(n1290) );
NOR2_X1 U923 ( .A1(n1292), .A2(n1293), .ZN(n1281) );
INV_X1 U924 ( .A(KEYINPUT46), .ZN(n1292) );
NOR2_X1 U925 ( .A1(KEYINPUT46), .A2(n1294), .ZN(n1280) );
NAND4_X1 U926 ( .A1(n1295), .A2(n1110), .A3(n1296), .A4(n1297), .ZN(n1294) );
NOR2_X1 U927 ( .A1(n1123), .A2(G952), .ZN(n1202) );
XNOR2_X1 U928 ( .A(G146), .B(n1264), .ZN(G48) );
NAND3_X1 U929 ( .A1(n1117), .A2(n1115), .A3(n1298), .ZN(n1264) );
XNOR2_X1 U930 ( .A(G143), .B(n1265), .ZN(G45) );
NAND4_X1 U931 ( .A1(n1299), .A2(n1300), .A3(n1115), .A4(n1296), .ZN(n1265) );
XOR2_X1 U932 ( .A(G140), .B(n1270), .Z(G42) );
AND3_X1 U933 ( .A1(n1106), .A2(n1113), .A3(n1275), .ZN(n1270) );
INV_X1 U934 ( .A(n1301), .ZN(n1275) );
XNOR2_X1 U935 ( .A(n1269), .B(n1302), .ZN(G39) );
XOR2_X1 U936 ( .A(KEYINPUT33), .B(G137), .Z(n1302) );
AND3_X1 U937 ( .A1(n1106), .A2(n1103), .A3(n1298), .ZN(n1269) );
XNOR2_X1 U938 ( .A(G134), .B(n1303), .ZN(G36) );
NOR2_X1 U939 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NOR3_X1 U940 ( .A1(n1306), .A2(n1307), .A3(n1120), .ZN(n1305) );
NOR2_X1 U941 ( .A1(n1289), .A2(n1308), .ZN(n1307) );
AND2_X1 U942 ( .A1(n1306), .A2(n1271), .ZN(n1304) );
NOR3_X1 U943 ( .A1(n1308), .A2(n1289), .A3(n1120), .ZN(n1271) );
INV_X1 U944 ( .A(KEYINPUT28), .ZN(n1306) );
XNOR2_X1 U945 ( .A(G131), .B(n1309), .ZN(G33) );
NAND2_X1 U946 ( .A1(KEYINPUT56), .A2(n1268), .ZN(n1309) );
AND3_X1 U947 ( .A1(n1300), .A2(n1117), .A3(n1106), .ZN(n1268) );
INV_X1 U948 ( .A(n1120), .ZN(n1106) );
NAND2_X1 U949 ( .A1(n1310), .A2(n1129), .ZN(n1120) );
INV_X1 U950 ( .A(n1308), .ZN(n1300) );
NAND2_X1 U951 ( .A1(n1311), .A2(n1112), .ZN(n1308) );
XNOR2_X1 U952 ( .A(G128), .B(n1312), .ZN(G30) );
NAND2_X1 U953 ( .A1(n1313), .A2(n1115), .ZN(n1312) );
XOR2_X1 U954 ( .A(n1273), .B(KEYINPUT22), .Z(n1313) );
NAND2_X1 U955 ( .A1(n1298), .A2(n1089), .ZN(n1273) );
AND2_X1 U956 ( .A1(n1311), .A2(n1133), .ZN(n1298) );
AND3_X1 U957 ( .A1(n1111), .A2(n1314), .A3(n1113), .ZN(n1311) );
XNOR2_X1 U958 ( .A(G101), .B(n1315), .ZN(G3) );
NAND2_X1 U959 ( .A1(KEYINPUT25), .A2(n1316), .ZN(n1315) );
INV_X1 U960 ( .A(n1277), .ZN(n1316) );
NAND4_X1 U961 ( .A1(n1103), .A2(n1091), .A3(n1112), .A4(n1111), .ZN(n1277) );
XOR2_X1 U962 ( .A(G125), .B(n1317), .Z(G27) );
NOR3_X1 U963 ( .A1(n1318), .A2(n1319), .A3(n1301), .ZN(n1317) );
NAND4_X1 U964 ( .A1(n1134), .A2(n1117), .A3(n1133), .A4(n1314), .ZN(n1301) );
NAND2_X1 U965 ( .A1(n1119), .A2(n1320), .ZN(n1314) );
NAND4_X1 U966 ( .A1(G953), .A2(G902), .A3(n1321), .A4(n1322), .ZN(n1320) );
INV_X1 U967 ( .A(G900), .ZN(n1322) );
XNOR2_X1 U968 ( .A(KEYINPUT34), .B(n1323), .ZN(n1318) );
XNOR2_X1 U969 ( .A(G122), .B(n1293), .ZN(G24) );
NAND3_X1 U970 ( .A1(n1295), .A2(n1296), .A3(n1114), .ZN(n1293) );
INV_X1 U971 ( .A(n1118), .ZN(n1114) );
NAND2_X1 U972 ( .A1(n1090), .A2(n1110), .ZN(n1118) );
INV_X1 U973 ( .A(n1297), .ZN(n1090) );
NAND2_X1 U974 ( .A1(n1112), .A2(n1134), .ZN(n1297) );
NOR3_X1 U975 ( .A1(n1323), .A2(n1226), .A3(n1324), .ZN(n1295) );
XNOR2_X1 U976 ( .A(G119), .B(n1278), .ZN(G21) );
NAND3_X1 U977 ( .A1(n1103), .A2(n1133), .A3(n1325), .ZN(n1278) );
XOR2_X1 U978 ( .A(n1326), .B(n1327), .Z(G18) );
NOR2_X1 U979 ( .A1(KEYINPUT9), .A2(n1328), .ZN(n1327) );
NOR2_X1 U980 ( .A1(n1329), .A2(n1291), .ZN(n1326) );
XNOR2_X1 U981 ( .A(n1089), .B(KEYINPUT62), .ZN(n1329) );
INV_X1 U982 ( .A(n1289), .ZN(n1089) );
NAND2_X1 U983 ( .A1(n1296), .A2(n1324), .ZN(n1289) );
XNOR2_X1 U984 ( .A(G113), .B(n1330), .ZN(G15) );
NAND2_X1 U985 ( .A1(n1117), .A2(n1331), .ZN(n1330) );
INV_X1 U986 ( .A(n1291), .ZN(n1331) );
NAND2_X1 U987 ( .A1(n1325), .A2(n1112), .ZN(n1291) );
XNOR2_X1 U988 ( .A(n1133), .B(KEYINPUT57), .ZN(n1112) );
NOR4_X1 U989 ( .A1(n1323), .A2(n1319), .A3(n1134), .A4(n1226), .ZN(n1325) );
INV_X1 U990 ( .A(n1332), .ZN(n1226) );
INV_X1 U991 ( .A(n1110), .ZN(n1319) );
NAND2_X1 U992 ( .A1(n1333), .A2(n1334), .ZN(n1110) );
OR3_X1 U993 ( .A1(n1140), .A2(n1139), .A3(KEYINPUT27), .ZN(n1334) );
NAND2_X1 U994 ( .A1(KEYINPUT27), .A2(n1113), .ZN(n1333) );
NOR2_X1 U995 ( .A1(n1324), .A2(n1296), .ZN(n1117) );
XNOR2_X1 U996 ( .A(G110), .B(n1276), .ZN(G12) );
NAND4_X1 U997 ( .A1(n1103), .A2(n1091), .A3(n1134), .A4(n1133), .ZN(n1276) );
XNOR2_X1 U998 ( .A(n1335), .B(n1336), .ZN(n1133) );
AND2_X1 U999 ( .A1(n1337), .A2(G217), .ZN(n1336) );
NAND2_X1 U1000 ( .A1(n1338), .A2(n1263), .ZN(n1335) );
XOR2_X1 U1001 ( .A(n1207), .B(KEYINPUT42), .Z(n1338) );
NAND2_X1 U1002 ( .A1(n1339), .A2(n1340), .ZN(n1207) );
NAND2_X1 U1003 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1004 ( .A(KEYINPUT11), .B(n1343), .Z(n1339) );
NOR2_X1 U1005 ( .A1(n1341), .A2(n1342), .ZN(n1343) );
XNOR2_X1 U1006 ( .A(n1344), .B(n1345), .ZN(n1342) );
XNOR2_X1 U1007 ( .A(n1346), .B(n1347), .ZN(n1345) );
XNOR2_X1 U1008 ( .A(KEYINPUT24), .B(n1348), .ZN(n1347) );
XNOR2_X1 U1009 ( .A(n1349), .B(n1350), .ZN(n1344) );
NOR2_X1 U1010 ( .A1(KEYINPUT12), .A2(n1351), .ZN(n1350) );
NOR2_X1 U1011 ( .A1(G128), .A2(KEYINPUT7), .ZN(n1349) );
XNOR2_X1 U1012 ( .A(n1352), .B(n1353), .ZN(n1341) );
NAND3_X1 U1013 ( .A1(G234), .A2(n1123), .A3(G221), .ZN(n1352) );
INV_X1 U1014 ( .A(n1111), .ZN(n1134) );
XOR2_X1 U1015 ( .A(n1165), .B(G472), .Z(n1111) );
INV_X1 U1016 ( .A(n1162), .ZN(n1165) );
NAND2_X1 U1017 ( .A1(n1354), .A2(n1263), .ZN(n1162) );
XOR2_X1 U1018 ( .A(n1355), .B(n1356), .Z(n1354) );
XOR2_X1 U1019 ( .A(KEYINPUT30), .B(KEYINPUT18), .Z(n1356) );
XNOR2_X1 U1020 ( .A(n1230), .B(n1233), .ZN(n1355) );
XNOR2_X1 U1021 ( .A(n1357), .B(n1358), .ZN(n1230) );
XOR2_X1 U1022 ( .A(n1359), .B(n1360), .Z(n1358) );
NOR2_X1 U1023 ( .A1(KEYINPUT26), .A2(n1348), .ZN(n1360) );
INV_X1 U1024 ( .A(G119), .ZN(n1348) );
AND2_X1 U1025 ( .A1(G210), .A2(n1361), .ZN(n1359) );
XNOR2_X1 U1026 ( .A(n1248), .B(n1362), .ZN(n1357) );
XOR2_X1 U1027 ( .A(n1363), .B(n1364), .Z(n1248) );
INV_X1 U1028 ( .A(n1285), .ZN(n1091) );
NAND3_X1 U1029 ( .A1(n1115), .A2(n1332), .A3(n1113), .ZN(n1285) );
NOR2_X1 U1030 ( .A1(n1365), .A2(n1139), .ZN(n1113) );
INV_X1 U1031 ( .A(n1152), .ZN(n1139) );
NAND2_X1 U1032 ( .A1(G221), .A2(n1337), .ZN(n1152) );
NAND2_X1 U1033 ( .A1(n1366), .A2(n1263), .ZN(n1337) );
XOR2_X1 U1034 ( .A(KEYINPUT35), .B(G234), .Z(n1366) );
INV_X1 U1035 ( .A(n1140), .ZN(n1365) );
XOR2_X1 U1036 ( .A(G469), .B(n1367), .Z(n1140) );
NOR2_X1 U1037 ( .A1(G902), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1038 ( .A(n1369), .B(n1370), .Z(n1368) );
XOR2_X1 U1039 ( .A(n1364), .B(n1371), .Z(n1370) );
NOR2_X1 U1040 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
AND3_X1 U1041 ( .A1(KEYINPUT44), .A2(n1346), .A3(G140), .ZN(n1373) );
NOR2_X1 U1042 ( .A1(KEYINPUT44), .A2(n1244), .ZN(n1372) );
INV_X1 U1043 ( .A(n1240), .ZN(n1244) );
XOR2_X1 U1044 ( .A(G140), .B(n1346), .Z(n1240) );
XOR2_X1 U1045 ( .A(n1182), .B(n1374), .Z(n1364) );
XOR2_X1 U1046 ( .A(KEYINPUT20), .B(G131), .Z(n1374) );
XOR2_X1 U1047 ( .A(G134), .B(n1353), .Z(n1182) );
XOR2_X1 U1048 ( .A(G137), .B(KEYINPUT60), .Z(n1353) );
XNOR2_X1 U1049 ( .A(n1241), .B(n1375), .ZN(n1369) );
NOR2_X1 U1050 ( .A1(KEYINPUT52), .A2(n1376), .ZN(n1375) );
XOR2_X1 U1051 ( .A(n1245), .B(n1363), .Z(n1376) );
XOR2_X1 U1052 ( .A(n1180), .B(n1377), .Z(n1245) );
NAND2_X1 U1053 ( .A1(n1378), .A2(n1379), .ZN(n1180) );
NAND2_X1 U1054 ( .A1(G128), .A2(n1380), .ZN(n1379) );
XOR2_X1 U1055 ( .A(KEYINPUT21), .B(n1381), .Z(n1378) );
NOR2_X1 U1056 ( .A1(G128), .A2(n1380), .ZN(n1381) );
XNOR2_X1 U1057 ( .A(G146), .B(n1382), .ZN(n1380) );
INV_X1 U1058 ( .A(n1236), .ZN(n1241) );
NAND2_X1 U1059 ( .A1(G227), .A2(n1123), .ZN(n1236) );
NAND2_X1 U1060 ( .A1(n1383), .A2(n1384), .ZN(n1332) );
NAND4_X1 U1061 ( .A1(G953), .A2(G902), .A3(n1321), .A4(n1200), .ZN(n1384) );
INV_X1 U1062 ( .A(G898), .ZN(n1200) );
XNOR2_X1 U1063 ( .A(n1101), .B(KEYINPUT8), .ZN(n1383) );
INV_X1 U1064 ( .A(n1119), .ZN(n1101) );
NAND3_X1 U1065 ( .A1(n1321), .A2(n1123), .A3(G952), .ZN(n1119) );
NAND2_X1 U1066 ( .A1(G237), .A2(G234), .ZN(n1321) );
INV_X1 U1067 ( .A(n1323), .ZN(n1115) );
NAND2_X1 U1068 ( .A1(n1128), .A2(n1129), .ZN(n1323) );
NAND2_X1 U1069 ( .A1(G214), .A2(n1385), .ZN(n1129) );
INV_X1 U1070 ( .A(n1310), .ZN(n1128) );
XNOR2_X1 U1071 ( .A(n1154), .B(n1156), .ZN(n1310) );
NAND2_X1 U1072 ( .A1(G210), .A2(n1385), .ZN(n1156) );
NAND2_X1 U1073 ( .A1(n1386), .A2(n1263), .ZN(n1385) );
INV_X1 U1074 ( .A(G237), .ZN(n1386) );
NAND2_X1 U1075 ( .A1(n1387), .A2(n1263), .ZN(n1154) );
INV_X1 U1076 ( .A(G902), .ZN(n1263) );
XOR2_X1 U1077 ( .A(n1388), .B(n1389), .Z(n1387) );
XNOR2_X1 U1078 ( .A(n1259), .B(n1233), .ZN(n1389) );
XNOR2_X1 U1079 ( .A(n1390), .B(n1391), .ZN(n1233) );
XOR2_X1 U1080 ( .A(G146), .B(G128), .Z(n1391) );
NAND2_X1 U1081 ( .A1(KEYINPUT16), .A2(n1382), .ZN(n1390) );
NAND2_X1 U1082 ( .A1(G224), .A2(n1123), .ZN(n1259) );
XOR2_X1 U1083 ( .A(n1392), .B(n1261), .Z(n1388) );
NOR2_X1 U1084 ( .A1(n1198), .A2(n1199), .ZN(n1261) );
NOR3_X1 U1085 ( .A1(n1197), .A2(n1194), .A3(n1196), .ZN(n1199) );
NAND2_X1 U1086 ( .A1(n1393), .A2(n1394), .ZN(n1198) );
NAND2_X1 U1087 ( .A1(n1194), .A2(n1395), .ZN(n1394) );
XOR2_X1 U1088 ( .A(n1197), .B(n1196), .Z(n1395) );
INV_X1 U1089 ( .A(n1396), .ZN(n1194) );
NAND3_X1 U1090 ( .A1(n1196), .A2(n1197), .A3(n1396), .ZN(n1393) );
NAND3_X1 U1091 ( .A1(n1397), .A2(n1398), .A3(n1399), .ZN(n1396) );
NAND2_X1 U1092 ( .A1(KEYINPUT31), .A2(n1400), .ZN(n1399) );
NAND3_X1 U1093 ( .A1(G122), .A2(n1401), .A3(n1346), .ZN(n1398) );
INV_X1 U1094 ( .A(G110), .ZN(n1346) );
NAND2_X1 U1095 ( .A1(G110), .A2(n1402), .ZN(n1397) );
NAND2_X1 U1096 ( .A1(n1403), .A2(n1401), .ZN(n1402) );
INV_X1 U1097 ( .A(KEYINPUT31), .ZN(n1401) );
XNOR2_X1 U1098 ( .A(KEYINPUT39), .B(n1400), .ZN(n1403) );
INV_X1 U1099 ( .A(G122), .ZN(n1400) );
XNOR2_X1 U1100 ( .A(n1362), .B(n1404), .ZN(n1197) );
NOR2_X1 U1101 ( .A1(G119), .A2(KEYINPUT2), .ZN(n1404) );
XNOR2_X1 U1102 ( .A(G113), .B(n1328), .ZN(n1362) );
INV_X1 U1103 ( .A(G116), .ZN(n1328) );
XNOR2_X1 U1104 ( .A(n1405), .B(n1377), .ZN(n1196) );
XNOR2_X1 U1105 ( .A(n1406), .B(n1407), .ZN(n1377) );
XNOR2_X1 U1106 ( .A(G107), .B(KEYINPUT14), .ZN(n1406) );
XNOR2_X1 U1107 ( .A(KEYINPUT0), .B(n1408), .ZN(n1405) );
NOR2_X1 U1108 ( .A1(KEYINPUT17), .A2(n1363), .ZN(n1408) );
XOR2_X1 U1109 ( .A(G101), .B(KEYINPUT29), .Z(n1363) );
NAND2_X1 U1110 ( .A1(KEYINPUT38), .A2(n1260), .ZN(n1392) );
XNOR2_X1 U1111 ( .A(G125), .B(KEYINPUT15), .ZN(n1260) );
NOR2_X1 U1112 ( .A1(n1296), .A2(n1299), .ZN(n1103) );
INV_X1 U1113 ( .A(n1324), .ZN(n1299) );
XOR2_X1 U1114 ( .A(n1409), .B(n1164), .Z(n1324) );
INV_X1 U1115 ( .A(n1216), .ZN(n1164) );
NOR2_X1 U1116 ( .A1(n1223), .A2(G902), .ZN(n1216) );
INV_X1 U1117 ( .A(n1219), .ZN(n1223) );
XNOR2_X1 U1118 ( .A(n1410), .B(n1411), .ZN(n1219) );
XNOR2_X1 U1119 ( .A(n1412), .B(n1407), .ZN(n1411) );
XOR2_X1 U1120 ( .A(G104), .B(KEYINPUT40), .Z(n1407) );
NAND2_X1 U1121 ( .A1(KEYINPUT63), .A2(n1413), .ZN(n1412) );
XNOR2_X1 U1122 ( .A(n1351), .B(n1414), .ZN(n1413) );
XOR2_X1 U1123 ( .A(n1415), .B(G131), .Z(n1414) );
NAND3_X1 U1124 ( .A1(n1416), .A2(n1417), .A3(KEYINPUT32), .ZN(n1415) );
NAND3_X1 U1125 ( .A1(n1418), .A2(n1419), .A3(n1420), .ZN(n1417) );
INV_X1 U1126 ( .A(KEYINPUT3), .ZN(n1420) );
NAND2_X1 U1127 ( .A1(n1421), .A2(KEYINPUT3), .ZN(n1416) );
XOR2_X1 U1128 ( .A(n1419), .B(n1418), .Z(n1421) );
XNOR2_X1 U1129 ( .A(G143), .B(KEYINPUT19), .ZN(n1418) );
NAND2_X1 U1130 ( .A1(n1361), .A2(G214), .ZN(n1419) );
NOR2_X1 U1131 ( .A1(G953), .A2(G237), .ZN(n1361) );
XOR2_X1 U1132 ( .A(G125), .B(n1422), .Z(n1351) );
XOR2_X1 U1133 ( .A(G146), .B(G140), .Z(n1422) );
XNOR2_X1 U1134 ( .A(G122), .B(n1423), .ZN(n1410) );
NOR2_X1 U1135 ( .A1(G113), .A2(KEYINPUT59), .ZN(n1423) );
NAND2_X1 U1136 ( .A1(KEYINPUT23), .A2(n1220), .ZN(n1409) );
INV_X1 U1137 ( .A(G475), .ZN(n1220) );
XNOR2_X1 U1138 ( .A(n1150), .B(n1151), .ZN(n1296) );
INV_X1 U1139 ( .A(G478), .ZN(n1151) );
NOR2_X1 U1140 ( .A1(n1213), .A2(G902), .ZN(n1150) );
XNOR2_X1 U1141 ( .A(n1424), .B(n1425), .ZN(n1213) );
XOR2_X1 U1142 ( .A(G128), .B(n1426), .Z(n1425) );
XNOR2_X1 U1143 ( .A(n1382), .B(G134), .ZN(n1426) );
INV_X1 U1144 ( .A(G143), .ZN(n1382) );
XOR2_X1 U1145 ( .A(n1427), .B(n1428), .Z(n1424) );
XNOR2_X1 U1146 ( .A(n1087), .B(n1429), .ZN(n1428) );
AND3_X1 U1147 ( .A1(G217), .A2(n1123), .A3(G234), .ZN(n1429) );
INV_X1 U1148 ( .A(G953), .ZN(n1123) );
INV_X1 U1149 ( .A(G107), .ZN(n1087) );
NAND2_X1 U1150 ( .A1(n1430), .A2(KEYINPUT58), .ZN(n1427) );
XNOR2_X1 U1151 ( .A(G116), .B(G122), .ZN(n1430) );
endmodule


