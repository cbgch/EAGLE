//Key = 0100010100000110011011111101000010011001000011101011000100011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413;

NAND3_X1 U784 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(G9) );
NAND2_X1 U785 ( .A1(KEYINPUT30), .A2(n1078), .ZN(n1077) );
OR3_X1 U786 ( .A1(n1078), .A2(KEYINPUT30), .A3(G107), .ZN(n1076) );
NAND2_X1 U787 ( .A1(G107), .A2(n1079), .ZN(n1075) );
NAND2_X1 U788 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
INV_X1 U789 ( .A(KEYINPUT30), .ZN(n1081) );
XNOR2_X1 U790 ( .A(KEYINPUT54), .B(n1078), .ZN(n1080) );
NOR2_X1 U791 ( .A1(n1082), .A2(n1083), .ZN(G75) );
NOR4_X1 U792 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1083) );
XOR2_X1 U793 ( .A(n1088), .B(KEYINPUT55), .Z(n1086) );
NAND4_X1 U794 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1088) );
INV_X1 U795 ( .A(n1093), .ZN(n1089) );
NAND4_X1 U796 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1084) );
NAND3_X1 U797 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1095) );
NAND2_X1 U798 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NAND3_X1 U799 ( .A1(n1103), .A2(n1104), .A3(n1090), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U801 ( .A1(n1107), .A2(n1108), .ZN(n1101) );
NAND2_X1 U802 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U803 ( .A1(n1090), .A2(n1111), .ZN(n1110) );
NAND2_X1 U804 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U805 ( .A1(n1103), .A2(n1114), .ZN(n1109) );
NAND2_X1 U806 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
OR2_X1 U807 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U808 ( .A1(n1090), .A2(n1119), .ZN(n1094) );
XOR2_X1 U809 ( .A(KEYINPUT2), .B(n1120), .Z(n1119) );
NOR3_X1 U810 ( .A1(n1093), .A2(n1092), .A3(n1091), .ZN(n1120) );
NAND3_X1 U811 ( .A1(n1107), .A2(n1103), .A3(n1100), .ZN(n1093) );
INV_X1 U812 ( .A(n1121), .ZN(n1100) );
NOR3_X1 U813 ( .A1(n1122), .A2(G953), .A3(G952), .ZN(n1082) );
INV_X1 U814 ( .A(n1096), .ZN(n1122) );
NAND4_X1 U815 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1096) );
NOR4_X1 U816 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
XOR2_X1 U817 ( .A(n1131), .B(n1132), .Z(n1127) );
NOR2_X1 U818 ( .A1(G472), .A2(n1133), .ZN(n1132) );
XNOR2_X1 U819 ( .A(KEYINPUT59), .B(KEYINPUT15), .ZN(n1133) );
NOR3_X1 U820 ( .A1(n1092), .A2(n1134), .A3(n1135), .ZN(n1125) );
NAND2_X1 U821 ( .A1(n1136), .A2(n1137), .ZN(n1124) );
XNOR2_X1 U822 ( .A(G478), .B(KEYINPUT20), .ZN(n1136) );
XOR2_X1 U823 ( .A(n1138), .B(n1139), .Z(n1123) );
XNOR2_X1 U824 ( .A(KEYINPUT62), .B(n1140), .ZN(n1139) );
XOR2_X1 U825 ( .A(n1141), .B(n1142), .Z(G72) );
NOR2_X1 U826 ( .A1(n1143), .A2(n1097), .ZN(n1142) );
AND2_X1 U827 ( .A1(G227), .A2(G900), .ZN(n1143) );
NAND2_X1 U828 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
NAND2_X1 U829 ( .A1(n1146), .A2(n1097), .ZN(n1145) );
XOR2_X1 U830 ( .A(n1147), .B(n1087), .Z(n1146) );
NAND3_X1 U831 ( .A1(G900), .A2(n1147), .A3(G953), .ZN(n1144) );
XNOR2_X1 U832 ( .A(n1148), .B(n1149), .ZN(n1147) );
XOR2_X1 U833 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U834 ( .A(n1152), .B(n1153), .Z(n1148) );
NOR3_X1 U835 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
NOR2_X1 U836 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
AND3_X1 U837 ( .A1(n1158), .A2(n1157), .A3(KEYINPUT50), .ZN(n1155) );
AND2_X1 U838 ( .A1(KEYINPUT60), .A2(n1159), .ZN(n1157) );
NOR2_X1 U839 ( .A1(KEYINPUT50), .A2(n1159), .ZN(n1154) );
NAND2_X1 U840 ( .A1(n1160), .A2(KEYINPUT45), .ZN(n1152) );
XNOR2_X1 U841 ( .A(n1161), .B(KEYINPUT34), .ZN(n1160) );
XOR2_X1 U842 ( .A(n1162), .B(n1163), .Z(G69) );
NAND2_X1 U843 ( .A1(G953), .A2(n1164), .ZN(n1163) );
NAND2_X1 U844 ( .A1(G898), .A2(G224), .ZN(n1164) );
NAND2_X1 U845 ( .A1(KEYINPUT17), .A2(n1165), .ZN(n1162) );
XOR2_X1 U846 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U847 ( .A1(n1097), .A2(n1085), .ZN(n1167) );
NAND2_X1 U848 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NAND2_X1 U849 ( .A1(G953), .A2(n1170), .ZN(n1169) );
XOR2_X1 U850 ( .A(n1171), .B(n1172), .Z(n1168) );
NOR2_X1 U851 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NOR3_X1 U852 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
NOR2_X1 U853 ( .A1(n1178), .A2(n1179), .ZN(n1173) );
INV_X1 U854 ( .A(n1175), .ZN(n1179) );
NOR2_X1 U855 ( .A1(n1176), .A2(n1177), .ZN(n1178) );
INV_X1 U856 ( .A(KEYINPUT5), .ZN(n1177) );
NOR2_X1 U857 ( .A1(n1180), .A2(n1181), .ZN(G66) );
XNOR2_X1 U858 ( .A(n1182), .B(n1183), .ZN(n1181) );
NOR2_X1 U859 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U860 ( .A1(n1180), .A2(n1186), .ZN(G63) );
XOR2_X1 U861 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND3_X1 U862 ( .A1(n1189), .A2(G478), .A3(KEYINPUT51), .ZN(n1187) );
NOR2_X1 U863 ( .A1(n1180), .A2(n1190), .ZN(G60) );
NOR3_X1 U864 ( .A1(n1138), .A2(n1191), .A3(n1192), .ZN(n1190) );
NOR2_X1 U865 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U866 ( .A1(n1195), .A2(n1140), .ZN(n1193) );
INV_X1 U867 ( .A(G475), .ZN(n1140) );
NOR2_X1 U868 ( .A1(n1087), .A2(n1085), .ZN(n1195) );
AND3_X1 U869 ( .A1(n1194), .A2(G475), .A3(n1189), .ZN(n1191) );
XOR2_X1 U870 ( .A(G104), .B(n1196), .Z(G6) );
NOR2_X1 U871 ( .A1(n1180), .A2(n1197), .ZN(G57) );
XOR2_X1 U872 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U873 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U874 ( .A1(KEYINPUT43), .A2(n1202), .ZN(n1200) );
XNOR2_X1 U875 ( .A(n1203), .B(n1204), .ZN(n1198) );
NAND2_X1 U876 ( .A1(KEYINPUT25), .A2(n1205), .ZN(n1204) );
NAND3_X1 U877 ( .A1(n1189), .A2(G472), .A3(KEYINPUT35), .ZN(n1203) );
NOR2_X1 U878 ( .A1(n1180), .A2(n1206), .ZN(G54) );
XOR2_X1 U879 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U880 ( .A(n1209), .B(n1210), .Z(n1208) );
AND2_X1 U881 ( .A1(G469), .A2(n1189), .ZN(n1210) );
INV_X1 U882 ( .A(n1185), .ZN(n1189) );
NOR2_X1 U883 ( .A1(G140), .A2(KEYINPUT10), .ZN(n1209) );
XNOR2_X1 U884 ( .A(n1211), .B(n1212), .ZN(n1207) );
XOR2_X1 U885 ( .A(G110), .B(n1213), .Z(n1212) );
NOR2_X1 U886 ( .A1(KEYINPUT38), .A2(n1214), .ZN(n1213) );
XOR2_X1 U887 ( .A(n1215), .B(n1216), .Z(n1214) );
NOR2_X1 U888 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
XOR2_X1 U889 ( .A(n1219), .B(KEYINPUT22), .Z(n1218) );
NAND2_X1 U890 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NOR2_X1 U891 ( .A1(n1220), .A2(n1221), .ZN(n1217) );
NOR2_X1 U892 ( .A1(n1180), .A2(n1222), .ZN(G51) );
NOR2_X1 U893 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U894 ( .A(n1225), .B(n1226), .Z(n1224) );
NOR2_X1 U895 ( .A1(KEYINPUT0), .A2(n1227), .ZN(n1226) );
XNOR2_X1 U896 ( .A(n1228), .B(n1229), .ZN(n1227) );
NOR2_X1 U897 ( .A1(n1230), .A2(n1185), .ZN(n1225) );
NAND2_X1 U898 ( .A1(G902), .A2(n1231), .ZN(n1185) );
OR2_X1 U899 ( .A1(n1085), .A2(n1087), .ZN(n1231) );
NAND4_X1 U900 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1087) );
NOR4_X1 U901 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
INV_X1 U902 ( .A(n1240), .ZN(n1239) );
NOR2_X1 U903 ( .A1(n1241), .A2(n1242), .ZN(n1234) );
NAND2_X1 U904 ( .A1(n1243), .A2(n1090), .ZN(n1233) );
XOR2_X1 U905 ( .A(n1244), .B(KEYINPUT18), .Z(n1243) );
NAND3_X1 U906 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
NAND2_X1 U907 ( .A1(n1248), .A2(n1249), .ZN(n1232) );
XOR2_X1 U908 ( .A(KEYINPUT47), .B(n1250), .Z(n1249) );
NAND4_X1 U909 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1085) );
NOR4_X1 U910 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1196), .ZN(n1254) );
AND3_X1 U911 ( .A1(n1258), .A2(n1103), .A3(n1245), .ZN(n1196) );
AND2_X1 U912 ( .A1(n1078), .A2(n1259), .ZN(n1253) );
NAND3_X1 U913 ( .A1(n1103), .A2(n1260), .A3(n1258), .ZN(n1078) );
NAND3_X1 U914 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1251) );
XNOR2_X1 U915 ( .A(n1248), .B(KEYINPUT39), .ZN(n1263) );
XNOR2_X1 U916 ( .A(G210), .B(KEYINPUT42), .ZN(n1230) );
NOR2_X1 U917 ( .A1(n1264), .A2(n1265), .ZN(n1223) );
INV_X1 U918 ( .A(KEYINPUT0), .ZN(n1265) );
XNOR2_X1 U919 ( .A(n1228), .B(n1266), .ZN(n1264) );
NAND2_X1 U920 ( .A1(n1267), .A2(n1268), .ZN(n1228) );
NOR2_X1 U921 ( .A1(n1097), .A2(G952), .ZN(n1180) );
XNOR2_X1 U922 ( .A(G146), .B(n1269), .ZN(G48) );
NAND2_X1 U923 ( .A1(n1250), .A2(n1248), .ZN(n1269) );
AND2_X1 U924 ( .A1(n1270), .A2(n1245), .ZN(n1250) );
NAND3_X1 U925 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(G45) );
NAND2_X1 U926 ( .A1(KEYINPUT61), .A2(n1242), .ZN(n1273) );
NAND3_X1 U927 ( .A1(n1274), .A2(n1275), .A3(G143), .ZN(n1272) );
NAND2_X1 U928 ( .A1(n1276), .A2(n1277), .ZN(n1271) );
NAND2_X1 U929 ( .A1(n1278), .A2(n1275), .ZN(n1276) );
INV_X1 U930 ( .A(KEYINPUT61), .ZN(n1275) );
XNOR2_X1 U931 ( .A(n1242), .B(KEYINPUT3), .ZN(n1278) );
INV_X1 U932 ( .A(n1274), .ZN(n1242) );
NAND3_X1 U933 ( .A1(n1279), .A2(n1280), .A3(n1247), .ZN(n1274) );
XNOR2_X1 U934 ( .A(G140), .B(n1281), .ZN(G42) );
NAND4_X1 U935 ( .A1(n1090), .A2(n1247), .A3(n1245), .A4(n1282), .ZN(n1281) );
XNOR2_X1 U936 ( .A(KEYINPUT49), .B(n1112), .ZN(n1282) );
XNOR2_X1 U937 ( .A(n1158), .B(n1241), .ZN(G39) );
AND3_X1 U938 ( .A1(n1270), .A2(n1107), .A3(n1090), .ZN(n1241) );
XNOR2_X1 U939 ( .A(G134), .B(n1240), .ZN(G36) );
NAND2_X1 U940 ( .A1(n1283), .A2(n1260), .ZN(n1240) );
XOR2_X1 U941 ( .A(n1238), .B(n1284), .Z(G33) );
NOR2_X1 U942 ( .A1(KEYINPUT12), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U943 ( .A(G131), .B(KEYINPUT53), .ZN(n1285) );
AND2_X1 U944 ( .A1(n1283), .A2(n1245), .ZN(n1238) );
AND3_X1 U945 ( .A1(n1247), .A2(n1280), .A3(n1090), .ZN(n1283) );
NOR2_X1 U946 ( .A1(n1118), .A2(n1135), .ZN(n1090) );
XNOR2_X1 U947 ( .A(n1130), .B(KEYINPUT46), .ZN(n1118) );
XOR2_X1 U948 ( .A(G128), .B(n1237), .Z(G30) );
AND3_X1 U949 ( .A1(n1260), .A2(n1248), .A3(n1270), .ZN(n1237) );
AND3_X1 U950 ( .A1(n1286), .A2(n1287), .A3(n1247), .ZN(n1270) );
NOR3_X1 U951 ( .A1(n1288), .A2(n1092), .A3(n1091), .ZN(n1247) );
NAND2_X1 U952 ( .A1(KEYINPUT8), .A2(n1112), .ZN(n1287) );
INV_X1 U953 ( .A(n1246), .ZN(n1112) );
NAND2_X1 U954 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
INV_X1 U955 ( .A(KEYINPUT8), .ZN(n1290) );
NAND2_X1 U956 ( .A1(n1128), .A2(n1291), .ZN(n1289) );
XOR2_X1 U957 ( .A(G101), .B(n1257), .Z(G3) );
AND3_X1 U958 ( .A1(n1107), .A2(n1258), .A3(n1280), .ZN(n1257) );
XOR2_X1 U959 ( .A(G125), .B(n1236), .Z(G27) );
AND4_X1 U960 ( .A1(n1245), .A2(n1098), .A3(n1292), .A4(n1246), .ZN(n1236) );
NOR2_X1 U961 ( .A1(n1288), .A2(n1115), .ZN(n1292) );
AND2_X1 U962 ( .A1(n1121), .A2(n1293), .ZN(n1288) );
NAND4_X1 U963 ( .A1(G953), .A2(G902), .A3(n1294), .A4(n1295), .ZN(n1293) );
INV_X1 U964 ( .A(G900), .ZN(n1295) );
XNOR2_X1 U965 ( .A(G122), .B(n1252), .ZN(G24) );
NAND3_X1 U966 ( .A1(n1296), .A2(n1103), .A3(n1279), .ZN(n1252) );
AND3_X1 U967 ( .A1(n1248), .A2(n1297), .A3(n1298), .ZN(n1279) );
NOR2_X1 U968 ( .A1(n1291), .A2(n1128), .ZN(n1103) );
XNOR2_X1 U969 ( .A(n1299), .B(n1300), .ZN(G21) );
AND3_X1 U970 ( .A1(n1261), .A2(n1262), .A3(n1248), .ZN(n1300) );
XOR2_X1 U971 ( .A(KEYINPUT8), .B(n1291), .Z(n1262) );
AND3_X1 U972 ( .A1(n1107), .A2(n1128), .A3(n1296), .ZN(n1261) );
NAND2_X1 U973 ( .A1(n1301), .A2(n1302), .ZN(G18) );
OR2_X1 U974 ( .A1(n1259), .A2(G116), .ZN(n1302) );
XOR2_X1 U975 ( .A(n1303), .B(KEYINPUT19), .Z(n1301) );
NAND2_X1 U976 ( .A1(G116), .A2(n1259), .ZN(n1303) );
NAND4_X1 U977 ( .A1(n1280), .A2(n1296), .A3(n1260), .A4(n1248), .ZN(n1259) );
INV_X1 U978 ( .A(n1106), .ZN(n1260) );
NAND2_X1 U979 ( .A1(n1304), .A2(n1297), .ZN(n1106) );
INV_X1 U980 ( .A(n1305), .ZN(n1297) );
XOR2_X1 U981 ( .A(G113), .B(n1256), .Z(G15) );
AND4_X1 U982 ( .A1(n1280), .A2(n1245), .A3(n1296), .A4(n1248), .ZN(n1256) );
AND2_X1 U983 ( .A1(n1098), .A2(n1306), .ZN(n1296) );
AND2_X1 U984 ( .A1(n1307), .A2(n1091), .ZN(n1098) );
INV_X1 U985 ( .A(n1129), .ZN(n1091) );
XNOR2_X1 U986 ( .A(n1092), .B(KEYINPUT41), .ZN(n1307) );
INV_X1 U987 ( .A(n1308), .ZN(n1092) );
INV_X1 U988 ( .A(n1105), .ZN(n1245) );
NAND2_X1 U989 ( .A1(n1309), .A2(n1305), .ZN(n1105) );
XOR2_X1 U990 ( .A(n1298), .B(KEYINPUT33), .Z(n1309) );
INV_X1 U991 ( .A(n1113), .ZN(n1280) );
NAND2_X1 U992 ( .A1(n1310), .A2(n1291), .ZN(n1113) );
XOR2_X1 U993 ( .A(G110), .B(n1255), .Z(G12) );
AND3_X1 U994 ( .A1(n1246), .A2(n1258), .A3(n1107), .ZN(n1255) );
AND2_X1 U995 ( .A1(n1304), .A2(n1305), .ZN(n1107) );
NOR2_X1 U996 ( .A1(n1311), .A2(n1134), .ZN(n1305) );
NOR2_X1 U997 ( .A1(n1137), .A2(G478), .ZN(n1134) );
AND2_X1 U998 ( .A1(G478), .A2(n1137), .ZN(n1311) );
NAND2_X1 U999 ( .A1(n1188), .A2(n1312), .ZN(n1137) );
XOR2_X1 U1000 ( .A(n1313), .B(n1314), .Z(n1188) );
XOR2_X1 U1001 ( .A(G128), .B(n1315), .Z(n1314) );
XNOR2_X1 U1002 ( .A(n1277), .B(G134), .ZN(n1315) );
XOR2_X1 U1003 ( .A(n1316), .B(n1317), .Z(n1313) );
AND2_X1 U1004 ( .A1(G217), .A2(n1318), .ZN(n1317) );
NAND2_X1 U1005 ( .A1(KEYINPUT13), .A2(n1319), .ZN(n1316) );
XNOR2_X1 U1006 ( .A(G107), .B(n1320), .ZN(n1319) );
NAND2_X1 U1007 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
OR2_X1 U1008 ( .A1(n1323), .A2(G116), .ZN(n1322) );
XOR2_X1 U1009 ( .A(n1324), .B(KEYINPUT52), .Z(n1321) );
NAND2_X1 U1010 ( .A1(G116), .A2(n1323), .ZN(n1324) );
XOR2_X1 U1011 ( .A(n1298), .B(KEYINPUT23), .Z(n1304) );
XNOR2_X1 U1012 ( .A(n1138), .B(n1325), .ZN(n1298) );
NOR2_X1 U1013 ( .A1(G475), .A2(KEYINPUT56), .ZN(n1325) );
NOR2_X1 U1014 ( .A1(n1194), .A2(G902), .ZN(n1138) );
XNOR2_X1 U1015 ( .A(n1326), .B(n1327), .ZN(n1194) );
XOR2_X1 U1016 ( .A(n1328), .B(n1329), .Z(n1327) );
NAND2_X1 U1017 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1018 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
INV_X1 U1019 ( .A(n1334), .ZN(n1333) );
NAND2_X1 U1020 ( .A1(n1335), .A2(n1336), .ZN(n1332) );
NAND2_X1 U1021 ( .A1(G104), .A2(n1323), .ZN(n1336) );
NAND2_X1 U1022 ( .A1(n1337), .A2(G122), .ZN(n1335) );
NAND2_X1 U1023 ( .A1(n1334), .A2(n1338), .ZN(n1330) );
NAND2_X1 U1024 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
NAND2_X1 U1025 ( .A1(G104), .A2(G122), .ZN(n1340) );
NAND2_X1 U1026 ( .A1(n1337), .A2(n1323), .ZN(n1339) );
INV_X1 U1027 ( .A(G122), .ZN(n1323) );
XNOR2_X1 U1028 ( .A(G104), .B(KEYINPUT6), .ZN(n1337) );
NOR2_X1 U1029 ( .A1(G113), .A2(KEYINPUT26), .ZN(n1334) );
NAND2_X1 U1030 ( .A1(n1341), .A2(G214), .ZN(n1328) );
XOR2_X1 U1031 ( .A(n1342), .B(n1343), .Z(n1326) );
NOR2_X1 U1032 ( .A1(KEYINPUT9), .A2(n1344), .ZN(n1343) );
XNOR2_X1 U1033 ( .A(n1345), .B(n1161), .ZN(n1344) );
XOR2_X1 U1034 ( .A(G125), .B(G140), .Z(n1161) );
XNOR2_X1 U1035 ( .A(G131), .B(G143), .ZN(n1342) );
AND4_X1 U1036 ( .A1(n1248), .A2(n1129), .A3(n1306), .A4(n1308), .ZN(n1258) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1346), .ZN(n1308) );
NAND2_X1 U1038 ( .A1(n1121), .A2(n1347), .ZN(n1306) );
NAND4_X1 U1039 ( .A1(G953), .A2(G902), .A3(n1294), .A4(n1170), .ZN(n1347) );
INV_X1 U1040 ( .A(G898), .ZN(n1170) );
NAND3_X1 U1041 ( .A1(n1294), .A2(n1097), .A3(G952), .ZN(n1121) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1294) );
XNOR2_X1 U1043 ( .A(n1348), .B(G469), .ZN(n1129) );
NAND2_X1 U1044 ( .A1(n1349), .A2(n1312), .ZN(n1348) );
XOR2_X1 U1045 ( .A(n1350), .B(n1351), .Z(n1349) );
XOR2_X1 U1046 ( .A(n1352), .B(n1353), .Z(n1351) );
NAND2_X1 U1047 ( .A1(KEYINPUT27), .A2(n1221), .ZN(n1353) );
XNOR2_X1 U1048 ( .A(n1354), .B(n1355), .ZN(n1221) );
NOR2_X1 U1049 ( .A1(KEYINPUT31), .A2(G104), .ZN(n1355) );
XNOR2_X1 U1050 ( .A(G101), .B(G107), .ZN(n1354) );
NAND2_X1 U1051 ( .A1(KEYINPUT21), .A2(n1356), .ZN(n1352) );
NAND2_X1 U1052 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
NAND2_X1 U1053 ( .A1(n1359), .A2(n1211), .ZN(n1358) );
XOR2_X1 U1054 ( .A(KEYINPUT48), .B(n1360), .Z(n1357) );
NOR2_X1 U1055 ( .A1(n1359), .A2(n1211), .ZN(n1360) );
NAND2_X1 U1056 ( .A1(G227), .A2(n1097), .ZN(n1211) );
XOR2_X1 U1057 ( .A(n1220), .B(n1361), .Z(n1350) );
NOR2_X1 U1058 ( .A1(KEYINPUT28), .A2(n1216), .ZN(n1361) );
XNOR2_X1 U1059 ( .A(n1362), .B(G131), .ZN(n1216) );
XOR2_X1 U1060 ( .A(n1151), .B(G128), .Z(n1220) );
XOR2_X1 U1061 ( .A(n1363), .B(n1364), .Z(n1151) );
XNOR2_X1 U1062 ( .A(KEYINPUT36), .B(n1345), .ZN(n1364) );
NAND2_X1 U1063 ( .A1(KEYINPUT32), .A2(n1277), .ZN(n1363) );
INV_X1 U1064 ( .A(n1115), .ZN(n1248) );
NAND2_X1 U1065 ( .A1(n1130), .A2(n1117), .ZN(n1115) );
INV_X1 U1066 ( .A(n1135), .ZN(n1117) );
NOR2_X1 U1067 ( .A1(n1365), .A2(n1366), .ZN(n1135) );
INV_X1 U1068 ( .A(G214), .ZN(n1365) );
XNOR2_X1 U1069 ( .A(n1367), .B(n1368), .ZN(n1130) );
NOR2_X1 U1070 ( .A1(n1366), .A2(n1369), .ZN(n1368) );
INV_X1 U1071 ( .A(G210), .ZN(n1369) );
NOR2_X1 U1072 ( .A1(G902), .A2(G237), .ZN(n1366) );
NAND2_X1 U1073 ( .A1(n1370), .A2(n1312), .ZN(n1367) );
XNOR2_X1 U1074 ( .A(n1371), .B(n1266), .ZN(n1370) );
INV_X1 U1075 ( .A(n1229), .ZN(n1266) );
XOR2_X1 U1076 ( .A(n1172), .B(n1372), .Z(n1229) );
XNOR2_X1 U1077 ( .A(n1176), .B(n1175), .ZN(n1372) );
NAND2_X1 U1078 ( .A1(n1373), .A2(n1374), .ZN(n1176) );
NAND2_X1 U1079 ( .A1(G101), .A2(n1375), .ZN(n1374) );
XOR2_X1 U1080 ( .A(KEYINPUT24), .B(n1376), .Z(n1373) );
NOR2_X1 U1081 ( .A1(G101), .A2(n1375), .ZN(n1376) );
XNOR2_X1 U1082 ( .A(G104), .B(n1377), .ZN(n1375) );
NOR2_X1 U1083 ( .A1(G107), .A2(KEYINPUT58), .ZN(n1377) );
XOR2_X1 U1084 ( .A(G122), .B(n1378), .Z(n1172) );
NOR2_X1 U1085 ( .A1(G110), .A2(KEYINPUT16), .ZN(n1378) );
NAND2_X1 U1086 ( .A1(n1379), .A2(n1268), .ZN(n1371) );
NAND3_X1 U1087 ( .A1(n1380), .A2(n1097), .A3(G224), .ZN(n1268) );
XNOR2_X1 U1088 ( .A(KEYINPUT7), .B(n1267), .ZN(n1379) );
OR2_X1 U1089 ( .A1(n1380), .A2(n1381), .ZN(n1267) );
AND2_X1 U1090 ( .A1(G224), .A2(n1097), .ZN(n1381) );
XNOR2_X1 U1091 ( .A(n1382), .B(n1383), .ZN(n1380) );
XOR2_X1 U1092 ( .A(G128), .B(G125), .Z(n1383) );
NOR2_X1 U1093 ( .A1(n1291), .A2(n1310), .ZN(n1246) );
INV_X1 U1094 ( .A(n1128), .ZN(n1310) );
XOR2_X1 U1095 ( .A(n1384), .B(n1184), .Z(n1128) );
NAND2_X1 U1096 ( .A1(G217), .A2(n1346), .ZN(n1184) );
NAND2_X1 U1097 ( .A1(G234), .A2(n1312), .ZN(n1346) );
NAND2_X1 U1098 ( .A1(n1182), .A2(n1312), .ZN(n1384) );
XNOR2_X1 U1099 ( .A(n1385), .B(n1386), .ZN(n1182) );
XNOR2_X1 U1100 ( .A(n1359), .B(n1387), .ZN(n1386) );
XOR2_X1 U1101 ( .A(n1388), .B(n1389), .Z(n1387) );
NOR2_X1 U1102 ( .A1(G125), .A2(KEYINPUT4), .ZN(n1389) );
NAND2_X1 U1103 ( .A1(n1318), .A2(G221), .ZN(n1388) );
AND2_X1 U1104 ( .A1(G234), .A2(n1097), .ZN(n1318) );
INV_X1 U1105 ( .A(G953), .ZN(n1097) );
XOR2_X1 U1106 ( .A(G110), .B(G140), .Z(n1359) );
XOR2_X1 U1107 ( .A(n1390), .B(n1391), .Z(n1385) );
XNOR2_X1 U1108 ( .A(n1345), .B(G137), .ZN(n1391) );
NAND3_X1 U1109 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n1390) );
OR2_X1 U1110 ( .A1(n1299), .A2(G128), .ZN(n1394) );
NAND2_X1 U1111 ( .A1(KEYINPUT40), .A2(n1395), .ZN(n1393) );
NAND2_X1 U1112 ( .A1(n1396), .A2(n1299), .ZN(n1395) );
XNOR2_X1 U1113 ( .A(G128), .B(n1397), .ZN(n1396) );
NAND2_X1 U1114 ( .A1(n1398), .A2(n1399), .ZN(n1392) );
INV_X1 U1115 ( .A(KEYINPUT40), .ZN(n1399) );
NAND2_X1 U1116 ( .A1(n1400), .A2(n1401), .ZN(n1398) );
OR2_X1 U1117 ( .A1(n1397), .A2(G128), .ZN(n1401) );
NAND3_X1 U1118 ( .A1(n1397), .A2(n1299), .A3(G128), .ZN(n1400) );
XNOR2_X1 U1119 ( .A(KEYINPUT37), .B(KEYINPUT11), .ZN(n1397) );
XNOR2_X1 U1120 ( .A(n1131), .B(G472), .ZN(n1291) );
NAND2_X1 U1121 ( .A1(n1402), .A2(n1312), .ZN(n1131) );
INV_X1 U1122 ( .A(G902), .ZN(n1312) );
XNOR2_X1 U1123 ( .A(n1201), .B(n1403), .ZN(n1402) );
XOR2_X1 U1124 ( .A(n1202), .B(n1205), .Z(n1403) );
XOR2_X1 U1125 ( .A(n1382), .B(n1404), .Z(n1205) );
XOR2_X1 U1126 ( .A(n1150), .B(n1362), .Z(n1404) );
XNOR2_X1 U1127 ( .A(n1405), .B(n1158), .ZN(n1362) );
INV_X1 U1128 ( .A(G137), .ZN(n1158) );
NAND2_X1 U1129 ( .A1(KEYINPUT14), .A2(n1159), .ZN(n1405) );
INV_X1 U1130 ( .A(G134), .ZN(n1159) );
XNOR2_X1 U1131 ( .A(G131), .B(G128), .ZN(n1150) );
XOR2_X1 U1132 ( .A(n1406), .B(KEYINPUT57), .Z(n1382) );
NAND2_X1 U1133 ( .A1(n1407), .A2(n1408), .ZN(n1406) );
NAND2_X1 U1134 ( .A1(G146), .A2(n1277), .ZN(n1408) );
INV_X1 U1135 ( .A(G143), .ZN(n1277) );
XOR2_X1 U1136 ( .A(n1409), .B(KEYINPUT29), .Z(n1407) );
NAND2_X1 U1137 ( .A1(G143), .A2(n1345), .ZN(n1409) );
INV_X1 U1138 ( .A(G146), .ZN(n1345) );
NAND2_X1 U1139 ( .A1(n1341), .A2(G210), .ZN(n1202) );
NOR2_X1 U1140 ( .A1(G953), .A2(G237), .ZN(n1341) );
XNOR2_X1 U1141 ( .A(n1410), .B(n1411), .ZN(n1201) );
XOR2_X1 U1142 ( .A(KEYINPUT63), .B(KEYINPUT1), .Z(n1411) );
XNOR2_X1 U1143 ( .A(G101), .B(n1175), .ZN(n1410) );
XNOR2_X1 U1144 ( .A(n1412), .B(n1413), .ZN(n1175) );
XNOR2_X1 U1145 ( .A(KEYINPUT44), .B(n1299), .ZN(n1413) );
INV_X1 U1146 ( .A(G119), .ZN(n1299) );
XNOR2_X1 U1147 ( .A(G113), .B(G116), .ZN(n1412) );
endmodule


