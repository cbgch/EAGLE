//Key = 0100111010010011011111000111001011111001100010011100000000000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299;

XOR2_X1 U735 ( .A(G107), .B(n1007), .Z(G9) );
NOR2_X1 U736 ( .A1(n1008), .A2(n1009), .ZN(G75) );
NOR4_X1 U737 ( .A1(G953), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1009) );
NOR2_X1 U738 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR2_X1 U739 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
AND3_X1 U740 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
OR3_X1 U741 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1018) );
NOR3_X1 U742 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1020) );
XNOR2_X1 U743 ( .A(n1026), .B(n1027), .ZN(n1024) );
NOR3_X1 U744 ( .A1(n1028), .A2(n1025), .A3(n1023), .ZN(n1015) );
NAND3_X1 U745 ( .A1(n1026), .A2(n1027), .A3(n1029), .ZN(n1028) );
NAND2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U747 ( .A1(n1019), .A2(n1032), .ZN(n1031) );
OR2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U749 ( .A1(n1017), .A2(n1035), .ZN(n1030) );
NAND2_X1 U750 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR3_X1 U751 ( .A1(n1010), .A2(G953), .A3(G952), .ZN(n1008) );
AND4_X1 U752 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1010) );
NOR4_X1 U753 ( .A1(n1042), .A2(n1025), .A3(n1043), .A4(n1044), .ZN(n1041) );
XNOR2_X1 U754 ( .A(n1045), .B(n1046), .ZN(n1044) );
XOR2_X1 U755 ( .A(n1047), .B(n1048), .Z(n1043) );
XNOR2_X1 U756 ( .A(KEYINPUT4), .B(n1049), .ZN(n1048) );
NOR2_X1 U757 ( .A1(KEYINPUT23), .A2(G469), .ZN(n1049) );
AND3_X1 U758 ( .A1(n1026), .A2(n1050), .A3(n1027), .ZN(n1040) );
NAND2_X1 U759 ( .A1(n1051), .A2(n1052), .ZN(n1039) );
INV_X1 U760 ( .A(n1053), .ZN(n1052) );
XOR2_X1 U761 ( .A(n1054), .B(KEYINPUT48), .Z(n1051) );
XOR2_X1 U762 ( .A(n1055), .B(n1056), .Z(n1038) );
NAND2_X1 U763 ( .A1(KEYINPUT39), .A2(n1057), .ZN(n1056) );
XOR2_X1 U764 ( .A(n1058), .B(n1059), .Z(G72) );
XOR2_X1 U765 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR3_X1 U766 ( .A1(n1062), .A2(KEYINPUT61), .A3(n1063), .ZN(n1061) );
NOR2_X1 U767 ( .A1(G900), .A2(n1064), .ZN(n1063) );
XOR2_X1 U768 ( .A(n1065), .B(n1066), .Z(n1062) );
XOR2_X1 U769 ( .A(n1067), .B(n1068), .Z(n1066) );
XNOR2_X1 U770 ( .A(KEYINPUT27), .B(n1069), .ZN(n1068) );
NOR2_X1 U771 ( .A1(KEYINPUT38), .A2(G140), .ZN(n1067) );
XNOR2_X1 U772 ( .A(n1070), .B(n1071), .ZN(n1065) );
NAND2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(n1060) );
NAND2_X1 U774 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XNOR2_X1 U775 ( .A(KEYINPUT25), .B(n1076), .ZN(n1075) );
NAND2_X1 U776 ( .A1(G953), .A2(n1077), .ZN(n1058) );
NAND2_X1 U777 ( .A1(G900), .A2(G227), .ZN(n1077) );
XOR2_X1 U778 ( .A(n1078), .B(n1079), .Z(G69) );
XOR2_X1 U779 ( .A(n1080), .B(n1081), .Z(n1079) );
NAND2_X1 U780 ( .A1(G953), .A2(n1082), .ZN(n1081) );
NAND2_X1 U781 ( .A1(G898), .A2(G224), .ZN(n1082) );
NAND2_X1 U782 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
OR2_X1 U783 ( .A1(n1064), .A2(G898), .ZN(n1084) );
XNOR2_X1 U784 ( .A(n1085), .B(n1086), .ZN(n1083) );
NAND2_X1 U785 ( .A1(KEYINPUT1), .A2(n1087), .ZN(n1085) );
NOR2_X1 U786 ( .A1(n1088), .A2(G953), .ZN(n1078) );
NOR2_X1 U787 ( .A1(n1089), .A2(n1090), .ZN(G66) );
XNOR2_X1 U788 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR2_X1 U789 ( .A1(n1054), .A2(n1093), .ZN(n1092) );
NOR2_X1 U790 ( .A1(n1089), .A2(n1094), .ZN(G63) );
XOR2_X1 U791 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U792 ( .A1(n1057), .A2(n1093), .ZN(n1096) );
INV_X1 U793 ( .A(G478), .ZN(n1057) );
NAND2_X1 U794 ( .A1(KEYINPUT44), .A2(n1097), .ZN(n1095) );
NOR2_X1 U795 ( .A1(n1089), .A2(n1098), .ZN(G60) );
XOR2_X1 U796 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U797 ( .A1(n1101), .A2(n1093), .ZN(n1099) );
XOR2_X1 U798 ( .A(G104), .B(n1102), .Z(G6) );
NOR2_X1 U799 ( .A1(n1089), .A2(n1103), .ZN(G57) );
XOR2_X1 U800 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U801 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U802 ( .A1(G101), .A2(KEYINPUT16), .ZN(n1106) );
XOR2_X1 U803 ( .A(n1108), .B(n1109), .Z(n1104) );
XOR2_X1 U804 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U805 ( .A1(n1045), .A2(n1093), .ZN(n1108) );
NOR3_X1 U806 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(G54) );
AND3_X1 U807 ( .A1(KEYINPUT2), .A2(G953), .A3(G952), .ZN(n1114) );
NOR2_X1 U808 ( .A1(KEYINPUT2), .A2(n1115), .ZN(n1113) );
INV_X1 U809 ( .A(n1089), .ZN(n1115) );
XOR2_X1 U810 ( .A(n1116), .B(n1117), .Z(n1112) );
XOR2_X1 U811 ( .A(n1107), .B(n1118), .Z(n1117) );
XOR2_X1 U812 ( .A(n1119), .B(n1120), .Z(n1116) );
XOR2_X1 U813 ( .A(KEYINPUT41), .B(G110), .Z(n1120) );
NOR2_X1 U814 ( .A1(n1121), .A2(n1093), .ZN(n1119) );
NOR2_X1 U815 ( .A1(n1089), .A2(n1122), .ZN(G51) );
XOR2_X1 U816 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U817 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U818 ( .A1(n1127), .A2(n1093), .ZN(n1125) );
NAND2_X1 U819 ( .A1(n1128), .A2(n1012), .ZN(n1093) );
NAND3_X1 U820 ( .A1(n1074), .A2(n1076), .A3(n1088), .ZN(n1012) );
AND2_X1 U821 ( .A1(n1129), .A2(n1130), .ZN(n1088) );
NOR4_X1 U822 ( .A1(n1131), .A2(n1132), .A3(n1102), .A4(n1007), .ZN(n1130) );
AND4_X1 U823 ( .A1(n1133), .A2(n1034), .A3(n1019), .A4(n1134), .ZN(n1007) );
AND4_X1 U824 ( .A1(n1033), .A2(n1133), .A3(n1019), .A4(n1134), .ZN(n1102) );
AND4_X1 U825 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1129) );
OR2_X1 U826 ( .A1(n1139), .A2(n1036), .ZN(n1138) );
INV_X1 U827 ( .A(n1140), .ZN(n1036) );
AND4_X1 U828 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1074) );
NOR4_X1 U829 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1144) );
NAND4_X1 U830 ( .A1(n1149), .A2(n1034), .A3(n1150), .A4(n1151), .ZN(n1143) );
XOR2_X1 U831 ( .A(KEYINPUT51), .B(n1152), .Z(n1151) );
XNOR2_X1 U832 ( .A(KEYINPUT3), .B(n1153), .ZN(n1128) );
NOR2_X1 U833 ( .A1(n1072), .A2(G952), .ZN(n1089) );
XNOR2_X1 U834 ( .A(G146), .B(n1141), .ZN(G48) );
NAND3_X1 U835 ( .A1(n1033), .A2(n1133), .A3(n1149), .ZN(n1141) );
NAND3_X1 U836 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(G45) );
NAND2_X1 U837 ( .A1(G143), .A2(n1142), .ZN(n1156) );
NAND2_X1 U838 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
INV_X1 U839 ( .A(KEYINPUT36), .ZN(n1158) );
NAND2_X1 U840 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
INV_X1 U841 ( .A(n1142), .ZN(n1160) );
XNOR2_X1 U842 ( .A(KEYINPUT29), .B(G143), .ZN(n1159) );
NAND2_X1 U843 ( .A1(KEYINPUT36), .A2(n1161), .ZN(n1154) );
NAND2_X1 U844 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
OR3_X1 U845 ( .A1(n1142), .A2(G143), .A3(KEYINPUT29), .ZN(n1163) );
NAND3_X1 U846 ( .A1(n1140), .A2(n1133), .A3(n1164), .ZN(n1142) );
AND3_X1 U847 ( .A1(n1042), .A2(n1165), .A3(n1166), .ZN(n1164) );
NAND2_X1 U848 ( .A1(KEYINPUT29), .A2(G143), .ZN(n1162) );
XNOR2_X1 U849 ( .A(G140), .B(n1167), .ZN(G42) );
NAND2_X1 U850 ( .A1(KEYINPUT32), .A2(n1147), .ZN(n1167) );
AND3_X1 U851 ( .A1(n1033), .A2(n1168), .A3(n1169), .ZN(n1147) );
XOR2_X1 U852 ( .A(n1146), .B(n1170), .Z(G39) );
NOR2_X1 U853 ( .A1(KEYINPUT50), .A2(n1171), .ZN(n1170) );
AND4_X1 U854 ( .A1(n1169), .A2(n1017), .A3(n1172), .A4(n1173), .ZN(n1146) );
XNOR2_X1 U855 ( .A(G134), .B(n1076), .ZN(G36) );
NAND3_X1 U856 ( .A1(n1140), .A2(n1034), .A3(n1169), .ZN(n1076) );
NAND2_X1 U857 ( .A1(n1174), .A2(n1175), .ZN(G33) );
NAND2_X1 U858 ( .A1(n1176), .A2(n1069), .ZN(n1175) );
NAND2_X1 U859 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U860 ( .A1(KEYINPUT42), .A2(n1179), .ZN(n1178) );
OR2_X1 U861 ( .A1(n1180), .A2(KEYINPUT42), .ZN(n1177) );
NAND2_X1 U862 ( .A1(G131), .A2(n1180), .ZN(n1174) );
NOR2_X1 U863 ( .A1(n1148), .A2(KEYINPUT24), .ZN(n1180) );
INV_X1 U864 ( .A(n1179), .ZN(n1148) );
NAND3_X1 U865 ( .A1(n1140), .A2(n1033), .A3(n1169), .ZN(n1179) );
AND2_X1 U866 ( .A1(n1022), .A2(n1166), .ZN(n1169) );
AND3_X1 U867 ( .A1(n1181), .A2(n1026), .A3(n1152), .ZN(n1022) );
INV_X1 U868 ( .A(n1025), .ZN(n1181) );
XNOR2_X1 U869 ( .A(n1182), .B(n1183), .ZN(G30) );
AND3_X1 U870 ( .A1(n1149), .A2(n1034), .A3(n1133), .ZN(n1183) );
AND3_X1 U871 ( .A1(n1166), .A2(n1173), .A3(n1172), .ZN(n1149) );
XNOR2_X1 U872 ( .A(G101), .B(n1184), .ZN(G3) );
NOR2_X1 U873 ( .A1(KEYINPUT46), .A2(n1185), .ZN(n1184) );
NOR2_X1 U874 ( .A1(n1186), .A2(n1139), .ZN(n1185) );
XNOR2_X1 U875 ( .A(n1140), .B(KEYINPUT45), .ZN(n1186) );
XOR2_X1 U876 ( .A(n1145), .B(n1187), .Z(G27) );
NOR2_X1 U877 ( .A1(KEYINPUT59), .A2(n1188), .ZN(n1187) );
AND4_X1 U878 ( .A1(n1033), .A2(n1021), .A3(n1168), .A4(n1166), .ZN(n1145) );
NAND2_X1 U879 ( .A1(n1189), .A2(n1014), .ZN(n1166) );
XOR2_X1 U880 ( .A(KEYINPUT21), .B(n1190), .Z(n1189) );
NOR4_X1 U881 ( .A1(G900), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1190) );
XNOR2_X1 U882 ( .A(KEYINPUT47), .B(n1064), .ZN(n1193) );
INV_X1 U883 ( .A(n1037), .ZN(n1168) );
XNOR2_X1 U884 ( .A(G122), .B(n1137), .ZN(G24) );
NAND4_X1 U885 ( .A1(n1194), .A2(n1019), .A3(n1042), .A4(n1165), .ZN(n1137) );
NOR2_X1 U886 ( .A1(n1173), .A2(n1172), .ZN(n1019) );
XOR2_X1 U887 ( .A(G119), .B(n1195), .Z(G21) );
NOR2_X1 U888 ( .A1(KEYINPUT58), .A2(n1136), .ZN(n1195) );
NAND4_X1 U889 ( .A1(n1194), .A2(n1017), .A3(n1172), .A4(n1173), .ZN(n1136) );
XNOR2_X1 U890 ( .A(G116), .B(n1135), .ZN(G18) );
NAND3_X1 U891 ( .A1(n1194), .A2(n1034), .A3(n1140), .ZN(n1135) );
AND2_X1 U892 ( .A1(n1196), .A2(n1165), .ZN(n1034) );
XOR2_X1 U893 ( .A(n1132), .B(n1197), .Z(G15) );
NOR2_X1 U894 ( .A1(KEYINPUT9), .A2(n1198), .ZN(n1197) );
AND3_X1 U895 ( .A1(n1033), .A2(n1194), .A3(n1140), .ZN(n1132) );
NOR2_X1 U896 ( .A1(n1173), .A2(n1199), .ZN(n1140) );
AND2_X1 U897 ( .A1(n1021), .A2(n1134), .ZN(n1194) );
AND3_X1 U898 ( .A1(n1150), .A2(n1027), .A3(n1200), .ZN(n1021) );
INV_X1 U899 ( .A(n1023), .ZN(n1200) );
NOR2_X1 U900 ( .A1(n1165), .A2(n1196), .ZN(n1033) );
INV_X1 U901 ( .A(n1042), .ZN(n1196) );
XOR2_X1 U902 ( .A(G110), .B(n1131), .Z(G12) );
NOR2_X1 U903 ( .A1(n1037), .A2(n1139), .ZN(n1131) );
NAND3_X1 U904 ( .A1(n1133), .A2(n1134), .A3(n1017), .ZN(n1139) );
NOR2_X1 U905 ( .A1(n1165), .A2(n1042), .ZN(n1017) );
XOR2_X1 U906 ( .A(n1201), .B(n1101), .Z(n1042) );
INV_X1 U907 ( .A(G475), .ZN(n1101) );
OR2_X1 U908 ( .A1(n1100), .A2(G902), .ZN(n1201) );
XNOR2_X1 U909 ( .A(n1202), .B(n1203), .ZN(n1100) );
XOR2_X1 U910 ( .A(n1204), .B(n1205), .Z(n1203) );
NOR2_X1 U911 ( .A1(KEYINPUT37), .A2(n1206), .ZN(n1204) );
XOR2_X1 U912 ( .A(n1207), .B(n1208), .Z(n1202) );
XNOR2_X1 U913 ( .A(n1069), .B(n1209), .ZN(n1208) );
NOR2_X1 U914 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U915 ( .A(n1212), .B(KEYINPUT17), .Z(n1211) );
NAND2_X1 U916 ( .A1(G104), .A2(n1213), .ZN(n1212) );
NOR2_X1 U917 ( .A1(G104), .A2(n1213), .ZN(n1210) );
XNOR2_X1 U918 ( .A(n1198), .B(n1214), .ZN(n1213) );
XOR2_X1 U919 ( .A(KEYINPUT13), .B(G122), .Z(n1214) );
INV_X1 U920 ( .A(G131), .ZN(n1069) );
NAND2_X1 U921 ( .A1(n1215), .A2(G214), .ZN(n1207) );
NAND2_X1 U922 ( .A1(n1216), .A2(n1217), .ZN(n1165) );
NAND2_X1 U923 ( .A1(G478), .A2(n1218), .ZN(n1217) );
XOR2_X1 U924 ( .A(n1219), .B(KEYINPUT0), .Z(n1216) );
OR2_X1 U925 ( .A1(n1218), .A2(G478), .ZN(n1219) );
XNOR2_X1 U926 ( .A(n1055), .B(KEYINPUT19), .ZN(n1218) );
NAND2_X1 U927 ( .A1(n1097), .A2(n1153), .ZN(n1055) );
XOR2_X1 U928 ( .A(n1220), .B(n1221), .Z(n1097) );
XOR2_X1 U929 ( .A(n1222), .B(n1223), .Z(n1221) );
AND3_X1 U930 ( .A1(G217), .A2(n1072), .A3(G234), .ZN(n1223) );
NOR2_X1 U931 ( .A1(KEYINPUT53), .A2(n1224), .ZN(n1222) );
XNOR2_X1 U932 ( .A(n1225), .B(n1226), .ZN(n1224) );
XNOR2_X1 U933 ( .A(G116), .B(G122), .ZN(n1225) );
NAND2_X1 U934 ( .A1(n1227), .A2(n1228), .ZN(n1220) );
NAND2_X1 U935 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
XOR2_X1 U936 ( .A(n1231), .B(KEYINPUT54), .Z(n1227) );
OR2_X1 U937 ( .A1(n1229), .A2(n1230), .ZN(n1231) );
XNOR2_X1 U938 ( .A(n1232), .B(n1206), .ZN(n1229) );
NAND2_X1 U939 ( .A1(KEYINPUT26), .A2(n1182), .ZN(n1232) );
INV_X1 U940 ( .A(G128), .ZN(n1182) );
NAND2_X1 U941 ( .A1(n1014), .A2(n1233), .ZN(n1134) );
OR4_X1 U942 ( .A1(n1192), .A2(n1064), .A3(n1191), .A4(G898), .ZN(n1233) );
INV_X1 U943 ( .A(n1234), .ZN(n1191) );
XOR2_X1 U944 ( .A(n1072), .B(KEYINPUT62), .Z(n1064) );
XOR2_X1 U945 ( .A(G902), .B(KEYINPUT63), .Z(n1192) );
NAND3_X1 U946 ( .A1(n1234), .A2(n1072), .A3(G952), .ZN(n1014) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1234) );
AND2_X1 U948 ( .A1(n1152), .A2(n1150), .ZN(n1133) );
AND2_X1 U949 ( .A1(n1235), .A2(n1026), .ZN(n1150) );
NAND2_X1 U950 ( .A1(G214), .A2(n1236), .ZN(n1026) );
XNOR2_X1 U951 ( .A(n1025), .B(KEYINPUT18), .ZN(n1235) );
XOR2_X1 U952 ( .A(n1237), .B(n1127), .Z(n1025) );
NAND2_X1 U953 ( .A1(G210), .A2(n1236), .ZN(n1127) );
NAND2_X1 U954 ( .A1(n1238), .A2(n1153), .ZN(n1236) );
INV_X1 U955 ( .A(G237), .ZN(n1238) );
NAND2_X1 U956 ( .A1(n1239), .A2(n1153), .ZN(n1237) );
XOR2_X1 U957 ( .A(n1240), .B(n1126), .Z(n1239) );
XNOR2_X1 U958 ( .A(n1070), .B(n1241), .ZN(n1126) );
NOR2_X1 U959 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XNOR2_X1 U960 ( .A(KEYINPUT22), .B(n1072), .ZN(n1243) );
INV_X1 U961 ( .A(G224), .ZN(n1242) );
XNOR2_X1 U962 ( .A(G125), .B(n1244), .ZN(n1070) );
NAND2_X1 U963 ( .A1(KEYINPUT8), .A2(n1123), .ZN(n1240) );
XNOR2_X1 U964 ( .A(n1087), .B(n1245), .ZN(n1123) );
INV_X1 U965 ( .A(n1086), .ZN(n1245) );
XNOR2_X1 U966 ( .A(n1246), .B(n1247), .ZN(n1086) );
XOR2_X1 U967 ( .A(G122), .B(G110), .Z(n1247) );
NAND2_X1 U968 ( .A1(n1248), .A2(n1249), .ZN(n1246) );
XOR2_X1 U969 ( .A(n1250), .B(KEYINPUT43), .Z(n1248) );
XNOR2_X1 U970 ( .A(G101), .B(n1251), .ZN(n1087) );
NOR2_X1 U971 ( .A1(KEYINPUT60), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U972 ( .A(n1253), .B(n1254), .ZN(n1252) );
NOR2_X1 U973 ( .A1(G104), .A2(KEYINPUT12), .ZN(n1254) );
AND2_X1 U974 ( .A1(n1023), .A2(n1027), .ZN(n1152) );
NAND2_X1 U975 ( .A1(G221), .A2(n1255), .ZN(n1027) );
XOR2_X1 U976 ( .A(n1047), .B(n1121), .Z(n1023) );
INV_X1 U977 ( .A(G469), .ZN(n1121) );
NAND2_X1 U978 ( .A1(n1256), .A2(n1153), .ZN(n1047) );
XOR2_X1 U979 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U980 ( .A(n1118), .B(n1259), .ZN(n1258) );
XNOR2_X1 U981 ( .A(n1260), .B(n1261), .ZN(n1118) );
XOR2_X1 U982 ( .A(G104), .B(n1262), .Z(n1261) );
XOR2_X1 U983 ( .A(KEYINPUT40), .B(G140), .Z(n1262) );
XNOR2_X1 U984 ( .A(n1263), .B(n1226), .ZN(n1260) );
INV_X1 U985 ( .A(n1253), .ZN(n1226) );
XOR2_X1 U986 ( .A(G107), .B(KEYINPUT20), .Z(n1253) );
XOR2_X1 U987 ( .A(n1264), .B(n1265), .Z(n1263) );
AND2_X1 U988 ( .A1(n1072), .A2(G227), .ZN(n1265) );
NAND2_X1 U989 ( .A1(KEYINPUT6), .A2(n1266), .ZN(n1264) );
XOR2_X1 U990 ( .A(KEYINPUT15), .B(G101), .Z(n1266) );
XOR2_X1 U991 ( .A(n1267), .B(n1268), .Z(n1257) );
NOR2_X1 U992 ( .A1(G110), .A2(KEYINPUT52), .ZN(n1268) );
NAND2_X1 U993 ( .A1(KEYINPUT5), .A2(n1244), .ZN(n1267) );
NAND2_X1 U994 ( .A1(n1199), .A2(n1173), .ZN(n1037) );
NAND2_X1 U995 ( .A1(n1269), .A2(n1050), .ZN(n1173) );
NAND2_X1 U996 ( .A1(n1053), .A2(n1054), .ZN(n1050) );
OR2_X1 U997 ( .A1(n1054), .A2(n1053), .ZN(n1269) );
NOR2_X1 U998 ( .A1(n1270), .A2(G902), .ZN(n1053) );
INV_X1 U999 ( .A(n1091), .ZN(n1270) );
XNOR2_X1 U1000 ( .A(n1271), .B(n1272), .ZN(n1091) );
NOR2_X1 U1001 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U1002 ( .A(KEYINPUT56), .B(n1275), .Z(n1274) );
AND2_X1 U1003 ( .A1(n1276), .A2(n1171), .ZN(n1275) );
NOR2_X1 U1004 ( .A1(n1171), .A2(n1276), .ZN(n1273) );
NAND3_X1 U1005 ( .A1(G234), .A2(n1072), .A3(G221), .ZN(n1276) );
INV_X1 U1006 ( .A(G953), .ZN(n1072) );
INV_X1 U1007 ( .A(G137), .ZN(n1171) );
NAND2_X1 U1008 ( .A1(KEYINPUT30), .A2(n1277), .ZN(n1271) );
XOR2_X1 U1009 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U1010 ( .A(G110), .B(n1280), .ZN(n1279) );
NOR2_X1 U1011 ( .A1(KEYINPUT7), .A2(n1281), .ZN(n1280) );
XOR2_X1 U1012 ( .A(G119), .B(n1282), .Z(n1281) );
NOR2_X1 U1013 ( .A1(G128), .A2(KEYINPUT55), .ZN(n1282) );
NAND2_X1 U1014 ( .A1(KEYINPUT34), .A2(n1205), .ZN(n1278) );
XNOR2_X1 U1015 ( .A(n1188), .B(n1283), .ZN(n1205) );
XNOR2_X1 U1016 ( .A(n1284), .B(G140), .ZN(n1283) );
INV_X1 U1017 ( .A(G146), .ZN(n1284) );
INV_X1 U1018 ( .A(G125), .ZN(n1188) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1255), .ZN(n1054) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1153), .ZN(n1255) );
INV_X1 U1021 ( .A(n1172), .ZN(n1199) );
XOR2_X1 U1022 ( .A(n1285), .B(n1045), .Z(n1172) );
INV_X1 U1023 ( .A(G472), .ZN(n1045) );
NAND2_X1 U1024 ( .A1(KEYINPUT35), .A2(n1046), .ZN(n1285) );
AND2_X1 U1025 ( .A1(n1286), .A2(n1153), .ZN(n1046) );
INV_X1 U1026 ( .A(G902), .ZN(n1153) );
XOR2_X1 U1027 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U1028 ( .A(n1110), .B(n1289), .Z(n1288) );
NOR2_X1 U1029 ( .A1(KEYINPUT28), .A2(n1290), .ZN(n1289) );
XOR2_X1 U1030 ( .A(n1291), .B(n1107), .Z(n1290) );
XOR2_X1 U1031 ( .A(n1244), .B(n1259), .Z(n1107) );
XNOR2_X1 U1032 ( .A(n1292), .B(G131), .ZN(n1259) );
NAND2_X1 U1033 ( .A1(KEYINPUT14), .A2(n1071), .ZN(n1292) );
XNOR2_X1 U1034 ( .A(G137), .B(n1230), .ZN(n1071) );
XOR2_X1 U1035 ( .A(G134), .B(KEYINPUT49), .Z(n1230) );
XNOR2_X1 U1036 ( .A(n1293), .B(n1206), .ZN(n1244) );
XOR2_X1 U1037 ( .A(G143), .B(KEYINPUT31), .Z(n1206) );
XNOR2_X1 U1038 ( .A(G146), .B(G128), .ZN(n1293) );
NAND2_X1 U1039 ( .A1(KEYINPUT33), .A2(n1294), .ZN(n1291) );
XNOR2_X1 U1040 ( .A(KEYINPUT57), .B(n1111), .ZN(n1294) );
NAND2_X1 U1041 ( .A1(n1250), .A2(n1249), .ZN(n1111) );
NAND2_X1 U1042 ( .A1(n1295), .A2(n1296), .ZN(n1249) );
XNOR2_X1 U1043 ( .A(KEYINPUT10), .B(n1198), .ZN(n1296) );
INV_X1 U1044 ( .A(G113), .ZN(n1198) );
XNOR2_X1 U1045 ( .A(G119), .B(n1297), .ZN(n1295) );
INV_X1 U1046 ( .A(G116), .ZN(n1297) );
NAND2_X1 U1047 ( .A1(n1298), .A2(n1299), .ZN(n1250) );
XNOR2_X1 U1048 ( .A(KEYINPUT10), .B(G113), .ZN(n1299) );
XNOR2_X1 U1049 ( .A(G116), .B(G119), .ZN(n1298) );
NAND2_X1 U1050 ( .A1(n1215), .A2(G210), .ZN(n1110) );
NOR2_X1 U1051 ( .A1(G953), .A2(G237), .ZN(n1215) );
NAND2_X1 U1052 ( .A1(KEYINPUT11), .A2(G101), .ZN(n1287) );
endmodule


