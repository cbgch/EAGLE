//Key = 0000111001100011000011011111111110001010100101110100000011011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376;

XOR2_X1 U751 ( .A(n1043), .B(n1044), .Z(G9) );
NOR2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1049) );
XOR2_X1 U756 ( .A(n1052), .B(KEYINPUT42), .Z(n1054) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
NAND4_X1 U758 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1047) );
NAND4_X1 U759 ( .A1(n1056), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1059) );
NAND2_X1 U760 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U761 ( .A1(KEYINPUT56), .A2(n1067), .ZN(n1066) );
NAND2_X1 U762 ( .A1(KEYINPUT56), .A2(n1057), .ZN(n1063) );
AND3_X1 U763 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1056) );
NAND4_X1 U764 ( .A1(n1070), .A2(n1062), .A3(n1057), .A4(n1071), .ZN(n1058) );
NAND2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U766 ( .A1(n1069), .A2(n1074), .ZN(n1073) );
OR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U768 ( .A1(n1068), .A2(n1077), .ZN(n1072) );
OR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
INV_X1 U770 ( .A(n1080), .ZN(n1070) );
AND3_X1 U771 ( .A1(n1060), .A2(n1061), .A3(n1081), .ZN(n1045) );
NAND4_X1 U772 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1060) );
NOR4_X1 U773 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1085) );
XOR2_X1 U774 ( .A(G475), .B(n1090), .Z(n1089) );
XOR2_X1 U775 ( .A(n1091), .B(n1092), .Z(n1088) );
XOR2_X1 U776 ( .A(n1093), .B(KEYINPUT14), .Z(n1087) );
XOR2_X1 U777 ( .A(n1094), .B(n1095), .Z(n1086) );
NOR2_X1 U778 ( .A1(KEYINPUT41), .A2(n1096), .ZN(n1095) );
XNOR2_X1 U779 ( .A(KEYINPUT52), .B(n1097), .ZN(n1096) );
NOR3_X1 U780 ( .A1(n1098), .A2(n1099), .A3(n1065), .ZN(n1084) );
NOR2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
XOR2_X1 U782 ( .A(n1102), .B(n1103), .Z(n1083) );
NOR2_X1 U783 ( .A1(KEYINPUT53), .A2(n1104), .ZN(n1103) );
XOR2_X1 U784 ( .A(n1105), .B(n1106), .Z(n1082) );
NAND2_X1 U785 ( .A1(KEYINPUT26), .A2(n1107), .ZN(n1106) );
XOR2_X1 U786 ( .A(n1108), .B(n1109), .Z(G72) );
NOR2_X1 U787 ( .A1(n1110), .A2(n1061), .ZN(n1109) );
NOR2_X1 U788 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U789 ( .A(KEYINPUT27), .B(G227), .Z(n1112) );
NAND2_X1 U790 ( .A1(n1113), .A2(n1114), .ZN(n1108) );
NAND2_X1 U791 ( .A1(n1115), .A2(n1061), .ZN(n1114) );
XNOR2_X1 U792 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND3_X1 U793 ( .A1(G900), .A2(n1117), .A3(G953), .ZN(n1113) );
XNOR2_X1 U794 ( .A(n1118), .B(n1119), .ZN(n1117) );
XOR2_X1 U795 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U796 ( .A(G140), .B(n1122), .ZN(n1121) );
NOR2_X1 U797 ( .A1(G131), .A2(KEYINPUT7), .ZN(n1122) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1118) );
XOR2_X1 U799 ( .A(n1125), .B(n1126), .Z(G69) );
NOR2_X1 U800 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U801 ( .A(n1129), .B(n1130), .ZN(n1128) );
NAND2_X1 U802 ( .A1(n1131), .A2(n1132), .ZN(n1125) );
NAND3_X1 U803 ( .A1(KEYINPUT21), .A2(n1133), .A3(n1061), .ZN(n1132) );
NAND2_X1 U804 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U805 ( .A(n1136), .B(KEYINPUT8), .Z(n1134) );
NAND3_X1 U806 ( .A1(KEYINPUT29), .A2(n1137), .A3(G953), .ZN(n1131) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1137) );
NOR2_X1 U808 ( .A1(n1138), .A2(n1139), .ZN(G66) );
XOR2_X1 U809 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR3_X1 U810 ( .A1(n1142), .A2(KEYINPUT12), .A3(n1143), .ZN(n1140) );
INV_X1 U811 ( .A(G217), .ZN(n1143) );
NOR2_X1 U812 ( .A1(n1138), .A2(n1144), .ZN(G63) );
NOR3_X1 U813 ( .A1(n1102), .A2(n1145), .A3(n1146), .ZN(n1144) );
AND3_X1 U814 ( .A1(n1147), .A2(G478), .A3(n1148), .ZN(n1146) );
NOR2_X1 U815 ( .A1(n1147), .A2(n1149), .ZN(n1145) );
AND2_X1 U816 ( .A1(n1048), .A2(G478), .ZN(n1149) );
NOR2_X1 U817 ( .A1(n1138), .A2(n1150), .ZN(G60) );
NOR3_X1 U818 ( .A1(n1090), .A2(n1151), .A3(n1152), .ZN(n1150) );
AND3_X1 U819 ( .A1(n1153), .A2(G475), .A3(n1148), .ZN(n1152) );
NOR2_X1 U820 ( .A1(n1154), .A2(n1153), .ZN(n1151) );
AND2_X1 U821 ( .A1(n1048), .A2(G475), .ZN(n1154) );
XOR2_X1 U822 ( .A(n1155), .B(n1156), .Z(G6) );
NOR2_X1 U823 ( .A1(n1138), .A2(n1157), .ZN(G57) );
XOR2_X1 U824 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U825 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U826 ( .A1(KEYINPUT36), .A2(n1162), .ZN(n1160) );
XOR2_X1 U827 ( .A(n1163), .B(n1164), .Z(n1158) );
NOR2_X1 U828 ( .A1(n1105), .A2(n1142), .ZN(n1164) );
INV_X1 U829 ( .A(G472), .ZN(n1105) );
NAND2_X1 U830 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
NAND2_X1 U831 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U832 ( .A(n1169), .B(KEYINPUT22), .Z(n1165) );
OR2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1169) );
NOR2_X1 U834 ( .A1(n1138), .A2(n1170), .ZN(G54) );
XOR2_X1 U835 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U836 ( .A(n1173), .B(n1123), .ZN(n1172) );
XOR2_X1 U837 ( .A(n1174), .B(n1175), .Z(n1171) );
XOR2_X1 U838 ( .A(KEYINPUT2), .B(n1176), .Z(n1175) );
AND2_X1 U839 ( .A1(G469), .A2(n1148), .ZN(n1176) );
INV_X1 U840 ( .A(n1142), .ZN(n1148) );
NOR3_X1 U841 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(G51) );
AND2_X1 U842 ( .A1(KEYINPUT62), .A2(n1138), .ZN(n1179) );
NOR2_X1 U843 ( .A1(n1061), .A2(G952), .ZN(n1138) );
NOR3_X1 U844 ( .A1(KEYINPUT62), .A2(n1061), .A3(n1081), .ZN(n1178) );
INV_X1 U845 ( .A(G952), .ZN(n1081) );
NOR2_X1 U846 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
XOR2_X1 U847 ( .A(n1182), .B(KEYINPUT6), .Z(n1181) );
NAND2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NOR2_X1 U849 ( .A1(n1183), .A2(n1184), .ZN(n1180) );
XOR2_X1 U850 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U851 ( .A1(n1142), .A2(n1091), .ZN(n1183) );
NAND2_X1 U852 ( .A1(G902), .A2(n1048), .ZN(n1142) );
NAND3_X1 U853 ( .A1(n1135), .A2(n1136), .A3(n1116), .ZN(n1048) );
AND4_X1 U854 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1116) );
NOR4_X1 U855 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190) );
NAND2_X1 U856 ( .A1(n1195), .A2(n1196), .ZN(n1189) );
NAND2_X1 U857 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U858 ( .A(KEYINPUT43), .B(n1199), .ZN(n1197) );
AND4_X1 U859 ( .A1(n1200), .A2(n1156), .A3(n1201), .A4(n1202), .ZN(n1135) );
AND3_X1 U860 ( .A1(n1203), .A2(n1044), .A3(n1204), .ZN(n1202) );
NAND3_X1 U861 ( .A1(n1205), .A2(n1076), .A3(n1078), .ZN(n1204) );
NAND3_X1 U862 ( .A1(n1076), .A2(n1069), .A3(n1206), .ZN(n1044) );
NAND2_X1 U863 ( .A1(n1207), .A2(n1195), .ZN(n1201) );
XOR2_X1 U864 ( .A(n1208), .B(KEYINPUT40), .Z(n1207) );
NAND3_X1 U865 ( .A1(n1206), .A2(n1069), .A3(n1075), .ZN(n1156) );
NAND2_X1 U866 ( .A1(n1068), .A2(n1209), .ZN(n1200) );
NAND2_X1 U867 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U868 ( .A1(n1078), .A2(n1206), .ZN(n1210) );
XOR2_X1 U869 ( .A(G146), .B(n1212), .Z(G48) );
NOR2_X1 U870 ( .A1(n1051), .A2(n1199), .ZN(n1212) );
NAND3_X1 U871 ( .A1(n1213), .A2(n1075), .A3(n1214), .ZN(n1199) );
XOR2_X1 U872 ( .A(G143), .B(n1215), .Z(G45) );
NOR2_X1 U873 ( .A1(n1216), .A2(n1198), .ZN(n1215) );
NAND4_X1 U874 ( .A1(n1078), .A2(n1213), .A3(n1217), .A4(n1218), .ZN(n1198) );
XOR2_X1 U875 ( .A(n1051), .B(KEYINPUT17), .Z(n1216) );
NAND2_X1 U876 ( .A1(n1219), .A2(n1220), .ZN(G42) );
OR2_X1 U877 ( .A1(n1187), .A2(G140), .ZN(n1220) );
XOR2_X1 U878 ( .A(n1221), .B(KEYINPUT35), .Z(n1219) );
NAND2_X1 U879 ( .A1(G140), .A2(n1187), .ZN(n1221) );
NAND3_X1 U880 ( .A1(n1075), .A2(n1079), .A3(n1222), .ZN(n1187) );
XOR2_X1 U881 ( .A(n1188), .B(n1223), .Z(G39) );
NAND2_X1 U882 ( .A1(KEYINPUT28), .A2(G137), .ZN(n1223) );
NAND3_X1 U883 ( .A1(n1214), .A2(n1068), .A3(n1222), .ZN(n1188) );
XNOR2_X1 U884 ( .A(n1194), .B(n1224), .ZN(G36) );
XOR2_X1 U885 ( .A(KEYINPUT25), .B(G134), .Z(n1224) );
AND3_X1 U886 ( .A1(n1222), .A2(n1076), .A3(n1078), .ZN(n1194) );
NAND3_X1 U887 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(G33) );
NAND2_X1 U888 ( .A1(G131), .A2(n1228), .ZN(n1227) );
NAND2_X1 U889 ( .A1(KEYINPUT0), .A2(n1229), .ZN(n1226) );
NAND2_X1 U890 ( .A1(n1193), .A2(n1230), .ZN(n1229) );
XOR2_X1 U891 ( .A(KEYINPUT46), .B(G131), .Z(n1230) );
NAND2_X1 U892 ( .A1(n1231), .A2(n1232), .ZN(n1225) );
INV_X1 U893 ( .A(KEYINPUT0), .ZN(n1232) );
NAND2_X1 U894 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
OR2_X1 U895 ( .A1(n1235), .A2(KEYINPUT46), .ZN(n1234) );
NAND3_X1 U896 ( .A1(n1193), .A2(n1235), .A3(KEYINPUT46), .ZN(n1233) );
INV_X1 U897 ( .A(n1228), .ZN(n1193) );
NAND3_X1 U898 ( .A1(n1222), .A2(n1075), .A3(n1078), .ZN(n1228) );
AND2_X1 U899 ( .A1(n1062), .A2(n1213), .ZN(n1222) );
NOR2_X1 U900 ( .A1(n1055), .A2(n1099), .ZN(n1062) );
INV_X1 U901 ( .A(n1053), .ZN(n1099) );
XOR2_X1 U902 ( .A(G128), .B(n1192), .Z(G30) );
AND4_X1 U903 ( .A1(n1214), .A2(n1213), .A3(n1076), .A4(n1195), .ZN(n1192) );
NOR3_X1 U904 ( .A1(n1236), .A2(n1065), .A3(n1067), .ZN(n1213) );
XOR2_X1 U905 ( .A(n1168), .B(n1237), .Z(G3) );
NAND4_X1 U906 ( .A1(n1078), .A2(n1068), .A3(n1238), .A4(n1239), .ZN(n1237) );
NOR3_X1 U907 ( .A1(n1067), .A2(n1065), .A3(n1240), .ZN(n1239) );
XOR2_X1 U908 ( .A(n1051), .B(KEYINPUT4), .Z(n1238) );
INV_X1 U909 ( .A(G101), .ZN(n1168) );
NAND2_X1 U910 ( .A1(n1241), .A2(n1242), .ZN(G27) );
NAND2_X1 U911 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
NAND2_X1 U912 ( .A1(G125), .A2(n1245), .ZN(n1241) );
NAND2_X1 U913 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U914 ( .A1(n1191), .A2(n1248), .ZN(n1247) );
INV_X1 U915 ( .A(n1249), .ZN(n1191) );
OR2_X1 U916 ( .A1(n1248), .A2(n1243), .ZN(n1246) );
NOR2_X1 U917 ( .A1(KEYINPUT11), .A2(n1249), .ZN(n1243) );
NAND4_X1 U918 ( .A1(n1075), .A2(n1057), .A3(n1250), .A4(n1079), .ZN(n1249) );
NOR2_X1 U919 ( .A1(n1236), .A2(n1051), .ZN(n1250) );
AND2_X1 U920 ( .A1(n1080), .A2(n1251), .ZN(n1236) );
NAND4_X1 U921 ( .A1(G902), .A2(G953), .A3(n1252), .A4(n1111), .ZN(n1251) );
INV_X1 U922 ( .A(G900), .ZN(n1111) );
INV_X1 U923 ( .A(KEYINPUT32), .ZN(n1248) );
XOR2_X1 U924 ( .A(n1253), .B(n1203), .Z(G24) );
NAND4_X1 U925 ( .A1(n1218), .A2(n1205), .A3(n1217), .A4(n1069), .ZN(n1203) );
NOR2_X1 U926 ( .A1(n1254), .A2(n1255), .ZN(n1069) );
XOR2_X1 U927 ( .A(G119), .B(n1256), .Z(G21) );
NOR3_X1 U928 ( .A1(n1211), .A2(KEYINPUT18), .A3(n1257), .ZN(n1256) );
INV_X1 U929 ( .A(n1068), .ZN(n1257) );
NAND2_X1 U930 ( .A1(n1205), .A2(n1214), .ZN(n1211) );
AND2_X1 U931 ( .A1(n1255), .A2(n1254), .ZN(n1214) );
NAND2_X1 U932 ( .A1(n1258), .A2(n1259), .ZN(G18) );
NAND3_X1 U933 ( .A1(KEYINPUT38), .A2(n1260), .A3(n1261), .ZN(n1259) );
NAND2_X1 U934 ( .A1(n1262), .A2(G116), .ZN(n1258) );
NAND2_X1 U935 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NAND2_X1 U936 ( .A1(n1260), .A2(n1265), .ZN(n1264) );
INV_X1 U937 ( .A(KEYINPUT45), .ZN(n1265) );
NAND2_X1 U938 ( .A1(KEYINPUT45), .A2(n1266), .ZN(n1263) );
NAND2_X1 U939 ( .A1(KEYINPUT38), .A2(n1260), .ZN(n1266) );
AND3_X1 U940 ( .A1(n1205), .A2(n1076), .A3(n1267), .ZN(n1260) );
XNOR2_X1 U941 ( .A(n1078), .B(KEYINPUT31), .ZN(n1267) );
AND2_X1 U942 ( .A1(n1217), .A2(n1268), .ZN(n1076) );
AND3_X1 U943 ( .A1(n1195), .A2(n1269), .A3(n1057), .ZN(n1205) );
INV_X1 U944 ( .A(n1051), .ZN(n1195) );
XOR2_X1 U945 ( .A(G113), .B(n1270), .Z(G15) );
NOR2_X1 U946 ( .A1(n1051), .A2(n1208), .ZN(n1270) );
NAND4_X1 U947 ( .A1(n1078), .A2(n1075), .A3(n1057), .A4(n1269), .ZN(n1208) );
NOR2_X1 U948 ( .A1(n1271), .A2(n1065), .ZN(n1057) );
INV_X1 U949 ( .A(n1067), .ZN(n1271) );
NOR2_X1 U950 ( .A1(n1268), .A2(n1217), .ZN(n1075) );
INV_X1 U951 ( .A(n1218), .ZN(n1268) );
NOR2_X1 U952 ( .A1(n1272), .A2(n1254), .ZN(n1078) );
XNOR2_X1 U953 ( .A(G110), .B(n1136), .ZN(G12) );
NAND3_X1 U954 ( .A1(n1079), .A2(n1206), .A3(n1068), .ZN(n1136) );
NOR2_X1 U955 ( .A1(n1218), .A2(n1217), .ZN(n1068) );
XNOR2_X1 U956 ( .A(n1273), .B(n1104), .ZN(n1217) );
XNOR2_X1 U957 ( .A(G478), .B(KEYINPUT49), .ZN(n1104) );
XNOR2_X1 U958 ( .A(n1102), .B(KEYINPUT63), .ZN(n1273) );
NOR2_X1 U959 ( .A1(n1147), .A2(G902), .ZN(n1102) );
AND2_X1 U960 ( .A1(n1274), .A2(n1275), .ZN(n1147) );
NAND3_X1 U961 ( .A1(G217), .A2(n1276), .A3(n1277), .ZN(n1275) );
XOR2_X1 U962 ( .A(n1278), .B(KEYINPUT10), .Z(n1277) );
NAND2_X1 U963 ( .A1(n1278), .A2(n1279), .ZN(n1274) );
NAND2_X1 U964 ( .A1(G217), .A2(n1276), .ZN(n1279) );
XOR2_X1 U965 ( .A(n1280), .B(n1281), .Z(n1278) );
XOR2_X1 U966 ( .A(G143), .B(G128), .Z(n1281) );
XOR2_X1 U967 ( .A(n1282), .B(n1283), .Z(n1280) );
NOR2_X1 U968 ( .A1(G134), .A2(KEYINPUT1), .ZN(n1283) );
NAND2_X1 U969 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND2_X1 U970 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U971 ( .A(KEYINPUT23), .B(n1288), .Z(n1284) );
NOR2_X1 U972 ( .A1(n1286), .A2(n1287), .ZN(n1288) );
NAND2_X1 U973 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
NAND2_X1 U974 ( .A1(G122), .A2(n1261), .ZN(n1290) );
INV_X1 U975 ( .A(G116), .ZN(n1261) );
XOR2_X1 U976 ( .A(n1291), .B(KEYINPUT34), .Z(n1289) );
NAND2_X1 U977 ( .A1(G116), .A2(n1253), .ZN(n1291) );
INV_X1 U978 ( .A(G122), .ZN(n1253) );
XOR2_X1 U979 ( .A(KEYINPUT5), .B(n1043), .Z(n1286) );
XNOR2_X1 U980 ( .A(n1090), .B(n1292), .ZN(n1218) );
NOR2_X1 U981 ( .A1(G475), .A2(KEYINPUT58), .ZN(n1292) );
NOR2_X1 U982 ( .A1(n1153), .A2(G902), .ZN(n1090) );
XOR2_X1 U983 ( .A(n1293), .B(G113), .Z(n1153) );
XOR2_X1 U984 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U985 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U986 ( .A(G122), .B(G104), .Z(n1297) );
XOR2_X1 U987 ( .A(G146), .B(G131), .Z(n1296) );
XOR2_X1 U988 ( .A(n1298), .B(n1299), .Z(n1294) );
XOR2_X1 U989 ( .A(n1300), .B(n1124), .Z(n1299) );
NOR2_X1 U990 ( .A1(G143), .A2(KEYINPUT44), .ZN(n1300) );
XOR2_X1 U991 ( .A(n1301), .B(n1302), .Z(n1298) );
NOR2_X1 U992 ( .A1(G140), .A2(KEYINPUT61), .ZN(n1302) );
NAND3_X1 U993 ( .A1(n1303), .A2(n1061), .A3(G214), .ZN(n1301) );
NOR4_X1 U994 ( .A1(n1051), .A2(n1067), .A3(n1240), .A4(n1065), .ZN(n1206) );
AND2_X1 U995 ( .A1(G221), .A2(n1304), .ZN(n1065) );
INV_X1 U996 ( .A(n1269), .ZN(n1240) );
NAND2_X1 U997 ( .A1(n1080), .A2(n1305), .ZN(n1269) );
NAND3_X1 U998 ( .A1(n1127), .A2(n1252), .A3(G902), .ZN(n1305) );
AND2_X1 U999 ( .A1(n1306), .A2(G953), .ZN(n1127) );
XNOR2_X1 U1000 ( .A(G898), .B(KEYINPUT13), .ZN(n1306) );
NAND3_X1 U1001 ( .A1(n1252), .A2(n1061), .A3(G952), .ZN(n1080) );
NAND2_X1 U1002 ( .A1(G237), .A2(n1307), .ZN(n1252) );
XOR2_X1 U1003 ( .A(n1097), .B(n1308), .Z(n1067) );
INV_X1 U1004 ( .A(n1094), .ZN(n1308) );
XNOR2_X1 U1005 ( .A(G469), .B(KEYINPUT37), .ZN(n1094) );
NAND2_X1 U1006 ( .A1(n1309), .A2(n1310), .ZN(n1097) );
XOR2_X1 U1007 ( .A(n1311), .B(n1174), .Z(n1309) );
XNOR2_X1 U1008 ( .A(n1312), .B(n1313), .ZN(n1174) );
XOR2_X1 U1009 ( .A(G140), .B(G110), .Z(n1313) );
NAND2_X1 U1010 ( .A1(G227), .A2(n1061), .ZN(n1312) );
NOR2_X1 U1011 ( .A1(KEYINPUT19), .A2(n1314), .ZN(n1311) );
XOR2_X1 U1012 ( .A(n1315), .B(n1173), .Z(n1314) );
XNOR2_X1 U1013 ( .A(n1316), .B(n1317), .ZN(n1173) );
XOR2_X1 U1014 ( .A(G101), .B(n1318), .Z(n1317) );
NOR2_X1 U1015 ( .A1(KEYINPUT16), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1016 ( .A(n1043), .B(n1320), .Z(n1319) );
NAND2_X1 U1017 ( .A1(KEYINPUT15), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1018 ( .A(KEYINPUT47), .B(G104), .Z(n1321) );
INV_X1 U1019 ( .A(G107), .ZN(n1043) );
NAND2_X1 U1020 ( .A1(KEYINPUT20), .A2(n1123), .ZN(n1315) );
XOR2_X1 U1021 ( .A(n1322), .B(n1323), .Z(n1123) );
NAND2_X1 U1022 ( .A1(n1055), .A2(n1053), .ZN(n1051) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1324), .ZN(n1053) );
NAND2_X1 U1024 ( .A1(n1325), .A2(n1326), .ZN(n1055) );
NAND2_X1 U1025 ( .A1(n1327), .A2(n1091), .ZN(n1326) );
NAND2_X1 U1026 ( .A1(n1092), .A2(n1328), .ZN(n1327) );
NAND2_X1 U1027 ( .A1(KEYINPUT33), .A2(KEYINPUT30), .ZN(n1328) );
NAND3_X1 U1028 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1325) );
INV_X1 U1029 ( .A(KEYINPUT33), .ZN(n1331) );
NAND2_X1 U1030 ( .A1(n1092), .A2(n1332), .ZN(n1330) );
INV_X1 U1031 ( .A(KEYINPUT30), .ZN(n1332) );
NAND2_X1 U1032 ( .A1(KEYINPUT30), .A2(n1333), .ZN(n1329) );
NAND2_X1 U1033 ( .A1(n1334), .A2(n1092), .ZN(n1333) );
NAND2_X1 U1034 ( .A1(n1335), .A2(n1310), .ZN(n1092) );
XOR2_X1 U1035 ( .A(n1336), .B(n1185), .Z(n1335) );
XOR2_X1 U1036 ( .A(n1337), .B(n1338), .Z(n1185) );
XOR2_X1 U1037 ( .A(n1339), .B(n1340), .Z(n1338) );
NAND2_X1 U1038 ( .A1(KEYINPUT9), .A2(n1129), .ZN(n1340) );
XOR2_X1 U1039 ( .A(G110), .B(n1341), .Z(n1129) );
XOR2_X1 U1040 ( .A(KEYINPUT24), .B(G122), .Z(n1341) );
NAND2_X1 U1041 ( .A1(G224), .A2(n1061), .ZN(n1339) );
XOR2_X1 U1042 ( .A(n1130), .B(n1342), .Z(n1337) );
XOR2_X1 U1043 ( .A(n1343), .B(n1344), .Z(n1130) );
XOR2_X1 U1044 ( .A(G107), .B(G101), .Z(n1344) );
XOR2_X1 U1045 ( .A(n1345), .B(n1346), .Z(n1343) );
NOR2_X1 U1046 ( .A1(KEYINPUT48), .A2(n1347), .ZN(n1346) );
XOR2_X1 U1047 ( .A(KEYINPUT47), .B(n1155), .Z(n1347) );
INV_X1 U1048 ( .A(G104), .ZN(n1155) );
NAND2_X1 U1049 ( .A1(KEYINPUT59), .A2(n1186), .ZN(n1336) );
INV_X1 U1050 ( .A(n1091), .ZN(n1334) );
NAND2_X1 U1051 ( .A1(G210), .A2(n1324), .ZN(n1091) );
NAND2_X1 U1052 ( .A1(n1310), .A2(n1303), .ZN(n1324) );
AND2_X1 U1053 ( .A1(n1272), .A2(n1254), .ZN(n1079) );
NAND2_X1 U1054 ( .A1(n1348), .A2(n1093), .ZN(n1254) );
NAND2_X1 U1055 ( .A1(n1100), .A2(n1101), .ZN(n1093) );
INV_X1 U1056 ( .A(n1349), .ZN(n1101) );
INV_X1 U1057 ( .A(n1350), .ZN(n1100) );
NAND2_X1 U1058 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1059 ( .A1(G217), .A2(n1304), .ZN(n1350) );
NAND2_X1 U1060 ( .A1(n1307), .A2(n1310), .ZN(n1304) );
XOR2_X1 U1061 ( .A(G234), .B(KEYINPUT39), .Z(n1307) );
NOR2_X1 U1062 ( .A1(n1141), .A2(G902), .ZN(n1349) );
XNOR2_X1 U1063 ( .A(n1351), .B(n1352), .ZN(n1141) );
XNOR2_X1 U1064 ( .A(n1323), .B(n1353), .ZN(n1352) );
XOR2_X1 U1065 ( .A(n1354), .B(n1355), .Z(n1353) );
NOR2_X1 U1066 ( .A1(KEYINPUT50), .A2(n1124), .ZN(n1355) );
INV_X1 U1067 ( .A(n1186), .ZN(n1124) );
XOR2_X1 U1068 ( .A(n1244), .B(KEYINPUT55), .Z(n1186) );
INV_X1 U1069 ( .A(G125), .ZN(n1244) );
NAND2_X1 U1070 ( .A1(n1276), .A2(G221), .ZN(n1354) );
AND2_X1 U1071 ( .A1(G234), .A2(n1061), .ZN(n1276) );
XOR2_X1 U1072 ( .A(G128), .B(G146), .Z(n1323) );
XOR2_X1 U1073 ( .A(n1356), .B(n1357), .Z(n1351) );
XOR2_X1 U1074 ( .A(G140), .B(G137), .Z(n1357) );
XNOR2_X1 U1075 ( .A(G119), .B(G110), .ZN(n1356) );
INV_X1 U1076 ( .A(n1255), .ZN(n1272) );
XOR2_X1 U1077 ( .A(n1358), .B(G472), .Z(n1255) );
NAND2_X1 U1078 ( .A1(KEYINPUT60), .A2(n1107), .ZN(n1358) );
NAND2_X1 U1079 ( .A1(n1359), .A2(n1310), .ZN(n1107) );
INV_X1 U1080 ( .A(G902), .ZN(n1310) );
XOR2_X1 U1081 ( .A(n1167), .B(n1360), .Z(n1359) );
XOR2_X1 U1082 ( .A(n1361), .B(G101), .Z(n1360) );
NAND2_X1 U1083 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
NAND2_X1 U1084 ( .A1(n1161), .A2(n1345), .ZN(n1363) );
XOR2_X1 U1085 ( .A(n1364), .B(KEYINPUT3), .Z(n1362) );
NAND2_X1 U1086 ( .A1(n1365), .A2(n1162), .ZN(n1364) );
INV_X1 U1087 ( .A(n1345), .ZN(n1162) );
XOR2_X1 U1088 ( .A(n1366), .B(n1367), .Z(n1345) );
XOR2_X1 U1089 ( .A(G119), .B(G116), .Z(n1367) );
INV_X1 U1090 ( .A(G113), .ZN(n1366) );
INV_X1 U1091 ( .A(n1161), .ZN(n1365) );
XOR2_X1 U1092 ( .A(n1342), .B(n1316), .Z(n1161) );
XNOR2_X1 U1093 ( .A(n1368), .B(n1120), .ZN(n1316) );
XNOR2_X1 U1094 ( .A(G134), .B(G137), .ZN(n1120) );
NAND2_X1 U1095 ( .A1(KEYINPUT57), .A2(n1235), .ZN(n1368) );
INV_X1 U1096 ( .A(G131), .ZN(n1235) );
XNOR2_X1 U1097 ( .A(n1369), .B(G128), .ZN(n1342) );
NAND3_X1 U1098 ( .A1(n1370), .A2(n1371), .A3(n1372), .ZN(n1369) );
NAND2_X1 U1099 ( .A1(KEYINPUT51), .A2(G143), .ZN(n1372) );
NAND3_X1 U1100 ( .A1(n1322), .A2(n1373), .A3(G146), .ZN(n1371) );
NAND2_X1 U1101 ( .A1(n1374), .A2(n1375), .ZN(n1370) );
INV_X1 U1102 ( .A(G146), .ZN(n1375) );
NAND2_X1 U1103 ( .A1(n1376), .A2(n1373), .ZN(n1374) );
INV_X1 U1104 ( .A(KEYINPUT51), .ZN(n1373) );
XOR2_X1 U1105 ( .A(n1322), .B(KEYINPUT54), .Z(n1376) );
INV_X1 U1106 ( .A(G143), .ZN(n1322) );
NAND3_X1 U1107 ( .A1(n1303), .A2(n1061), .A3(G210), .ZN(n1167) );
INV_X1 U1108 ( .A(G953), .ZN(n1061) );
INV_X1 U1109 ( .A(G237), .ZN(n1303) );
endmodule


