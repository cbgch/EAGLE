//Key = 0100111110001000110010011111010001001010111111011011101101000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382;

XOR2_X1 U759 ( .A(G107), .B(n1047), .Z(G9) );
NOR2_X1 U760 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U761 ( .A1(n1050), .A2(n1051), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
XOR2_X1 U763 ( .A(n1056), .B(KEYINPUT34), .Z(n1054) );
NAND3_X1 U764 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1052) );
NAND2_X1 U765 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U766 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U767 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NAND2_X1 U768 ( .A1(n1067), .A2(n1068), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U770 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
XNOR2_X1 U772 ( .A(KEYINPUT39), .B(n1076), .ZN(n1074) );
XOR2_X1 U773 ( .A(KEYINPUT53), .B(n1077), .Z(n1073) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1067) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1077), .A2(n1082), .ZN(n1081) );
NAND2_X1 U777 ( .A1(n1083), .A2(n1049), .ZN(n1082) );
NAND2_X1 U778 ( .A1(n1069), .A2(n1084), .ZN(n1080) );
OR2_X1 U779 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND3_X1 U780 ( .A1(n1087), .A2(n1088), .A3(n1077), .ZN(n1062) );
NAND2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U782 ( .A1(KEYINPUT28), .A2(n1091), .ZN(n1089) );
NAND3_X1 U783 ( .A1(n1092), .A2(n1093), .A3(n1069), .ZN(n1087) );
NAND3_X1 U784 ( .A1(n1066), .A2(n1078), .A3(n1094), .ZN(n1093) );
OR2_X1 U785 ( .A1(n1095), .A2(KEYINPUT28), .ZN(n1092) );
INV_X1 U786 ( .A(n1096), .ZN(n1060) );
NOR3_X1 U787 ( .A1(n1097), .A2(G953), .A3(G952), .ZN(n1050) );
INV_X1 U788 ( .A(n1057), .ZN(n1097) );
NAND4_X1 U789 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1057) );
NOR3_X1 U790 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NAND3_X1 U791 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1102) );
XOR2_X1 U792 ( .A(KEYINPUT63), .B(n1108), .Z(n1107) );
NAND2_X1 U793 ( .A1(G475), .A2(n1109), .ZN(n1106) );
NAND2_X1 U794 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
NOR3_X1 U795 ( .A1(n1075), .A2(n1112), .A3(n1094), .ZN(n1100) );
INV_X1 U796 ( .A(n1065), .ZN(n1094) );
XOR2_X1 U797 ( .A(n1113), .B(n1114), .Z(G72) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1058), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1113) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1058), .ZN(n1119) );
XOR2_X1 U802 ( .A(n1056), .B(n1121), .Z(n1120) );
NAND3_X1 U803 ( .A1(G900), .A2(n1121), .A3(G953), .ZN(n1118) );
XNOR2_X1 U804 ( .A(n1122), .B(n1123), .ZN(n1121) );
XNOR2_X1 U805 ( .A(n1124), .B(KEYINPUT49), .ZN(n1123) );
NAND2_X1 U806 ( .A1(n1125), .A2(KEYINPUT16), .ZN(n1124) );
XNOR2_X1 U807 ( .A(n1126), .B(n1127), .ZN(n1125) );
XOR2_X1 U808 ( .A(n1128), .B(G131), .Z(n1126) );
NAND3_X1 U809 ( .A1(n1129), .A2(n1130), .A3(KEYINPUT7), .ZN(n1128) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
INV_X1 U811 ( .A(KEYINPUT10), .ZN(n1132) );
XOR2_X1 U812 ( .A(n1133), .B(G134), .Z(n1131) );
NAND3_X1 U813 ( .A1(G134), .A2(n1133), .A3(KEYINPUT10), .ZN(n1129) );
XOR2_X1 U814 ( .A(n1134), .B(n1135), .Z(G69) );
NOR3_X1 U815 ( .A1(n1058), .A2(KEYINPUT30), .A3(n1136), .ZN(n1135) );
AND2_X1 U816 ( .A1(G224), .A2(G898), .ZN(n1136) );
NAND2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NAND2_X1 U818 ( .A1(n1139), .A2(n1058), .ZN(n1138) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
INV_X1 U821 ( .A(n1053), .ZN(n1142) );
NAND3_X1 U822 ( .A1(n1141), .A2(G898), .A3(G953), .ZN(n1137) );
NOR2_X1 U823 ( .A1(KEYINPUT13), .A2(n1144), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U825 ( .A(KEYINPUT2), .B(G110), .Z(n1146) );
NOR2_X1 U826 ( .A1(n1147), .A2(n1148), .ZN(G66) );
XOR2_X1 U827 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U828 ( .A1(KEYINPUT35), .A2(n1151), .ZN(n1150) );
NOR2_X1 U829 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
NOR2_X1 U830 ( .A1(n1147), .A2(n1154), .ZN(G63) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U832 ( .A1(n1157), .A2(n1153), .ZN(n1155) );
INV_X1 U833 ( .A(G478), .ZN(n1157) );
NOR2_X1 U834 ( .A1(n1147), .A2(n1158), .ZN(G60) );
XNOR2_X1 U835 ( .A(n1159), .B(n1160), .ZN(n1158) );
NOR2_X1 U836 ( .A1(n1161), .A2(n1153), .ZN(n1160) );
INV_X1 U837 ( .A(G475), .ZN(n1161) );
XOR2_X1 U838 ( .A(n1162), .B(n1163), .Z(G6) );
NAND2_X1 U839 ( .A1(KEYINPUT5), .A2(G104), .ZN(n1163) );
NAND2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
XOR2_X1 U841 ( .A(KEYINPUT37), .B(n1166), .Z(n1165) );
NOR2_X1 U842 ( .A1(n1147), .A2(n1167), .ZN(G57) );
NOR2_X1 U843 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U844 ( .A(KEYINPUT59), .B(n1170), .Z(n1169) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
AND2_X1 U846 ( .A1(n1172), .A2(n1171), .ZN(n1168) );
XNOR2_X1 U847 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR2_X1 U848 ( .A1(n1175), .A2(n1153), .ZN(n1174) );
INV_X1 U849 ( .A(G472), .ZN(n1175) );
NAND3_X1 U850 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1173) );
NAND3_X1 U851 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1178) );
NOR2_X1 U852 ( .A1(n1182), .A2(n1183), .ZN(G54) );
XOR2_X1 U853 ( .A(n1184), .B(n1185), .Z(n1183) );
XNOR2_X1 U854 ( .A(n1186), .B(KEYINPUT12), .ZN(n1185) );
NAND2_X1 U855 ( .A1(KEYINPUT47), .A2(n1187), .ZN(n1186) );
XOR2_X1 U856 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U857 ( .A(n1190), .B(n1127), .Z(n1189) );
XOR2_X1 U858 ( .A(n1191), .B(n1192), .Z(n1188) );
XNOR2_X1 U859 ( .A(KEYINPUT43), .B(n1193), .ZN(n1192) );
NOR2_X1 U860 ( .A1(KEYINPUT15), .A2(n1194), .ZN(n1193) );
XOR2_X1 U861 ( .A(n1195), .B(n1196), .Z(n1194) );
NAND2_X1 U862 ( .A1(KEYINPUT44), .A2(G110), .ZN(n1195) );
NAND2_X1 U863 ( .A1(KEYINPUT27), .A2(n1197), .ZN(n1191) );
NOR2_X1 U864 ( .A1(n1198), .A2(n1153), .ZN(n1184) );
INV_X1 U865 ( .A(G469), .ZN(n1198) );
NOR2_X1 U866 ( .A1(G952), .A2(n1199), .ZN(n1182) );
XOR2_X1 U867 ( .A(KEYINPUT51), .B(G953), .Z(n1199) );
NOR2_X1 U868 ( .A1(n1147), .A2(n1200), .ZN(G51) );
XNOR2_X1 U869 ( .A(n1201), .B(n1202), .ZN(n1200) );
NOR2_X1 U870 ( .A1(n1203), .A2(n1153), .ZN(n1202) );
NAND2_X1 U871 ( .A1(G902), .A2(n1204), .ZN(n1153) );
OR3_X1 U872 ( .A1(n1055), .A2(n1056), .A3(n1053), .ZN(n1204) );
NAND4_X1 U873 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1053) );
NOR4_X1 U874 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
NOR2_X1 U875 ( .A1(n1213), .A2(n1048), .ZN(n1212) );
INV_X1 U876 ( .A(n1164), .ZN(n1048) );
NOR3_X1 U877 ( .A1(n1214), .A2(n1215), .A3(n1071), .ZN(n1164) );
NAND2_X1 U878 ( .A1(n1077), .A2(n1216), .ZN(n1071) );
AND2_X1 U879 ( .A1(n1083), .A2(n1049), .ZN(n1213) );
AND3_X1 U880 ( .A1(n1085), .A2(n1216), .A3(n1217), .ZN(n1211) );
NOR2_X1 U881 ( .A1(n1218), .A2(n1219), .ZN(n1210) );
AND3_X1 U882 ( .A1(n1218), .A2(n1215), .A3(n1220), .ZN(n1209) );
INV_X1 U883 ( .A(KEYINPUT36), .ZN(n1218) );
NAND2_X1 U884 ( .A1(n1221), .A2(n1222), .ZN(n1205) );
XOR2_X1 U885 ( .A(KEYINPUT42), .B(n1215), .Z(n1222) );
NAND4_X1 U886 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1056) );
NOR3_X1 U887 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1226) );
NAND2_X1 U888 ( .A1(n1166), .A2(n1230), .ZN(n1225) );
NAND2_X1 U889 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND3_X1 U890 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1232) );
NAND2_X1 U891 ( .A1(n1085), .A2(n1236), .ZN(n1231) );
NAND2_X1 U892 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND2_X1 U893 ( .A1(n1091), .A2(n1239), .ZN(n1238) );
OR2_X1 U894 ( .A1(n1240), .A2(n1241), .ZN(n1223) );
XOR2_X1 U895 ( .A(n1143), .B(KEYINPUT57), .Z(n1055) );
AND2_X1 U896 ( .A1(n1242), .A2(n1243), .ZN(n1143) );
NAND4_X1 U897 ( .A1(n1244), .A2(n1234), .A3(n1245), .A4(n1246), .ZN(n1243) );
OR2_X1 U898 ( .A1(n1247), .A2(n1246), .ZN(n1242) );
INV_X1 U899 ( .A(KEYINPUT41), .ZN(n1246) );
NOR2_X1 U900 ( .A1(n1058), .A2(G952), .ZN(n1147) );
XOR2_X1 U901 ( .A(G146), .B(n1248), .Z(G48) );
NOR4_X1 U902 ( .A1(n1241), .A2(n1249), .A3(n1083), .A4(n1250), .ZN(n1248) );
XOR2_X1 U903 ( .A(n1251), .B(KEYINPUT22), .Z(n1249) );
XNOR2_X1 U904 ( .A(G143), .B(n1252), .ZN(G45) );
NAND2_X1 U905 ( .A1(n1253), .A2(n1234), .ZN(n1252) );
XOR2_X1 U906 ( .A(n1240), .B(KEYINPUT4), .Z(n1253) );
NAND4_X1 U907 ( .A1(n1254), .A2(n1235), .A3(n1086), .A4(n1255), .ZN(n1240) );
XNOR2_X1 U908 ( .A(KEYINPUT23), .B(n1104), .ZN(n1254) );
NAND2_X1 U909 ( .A1(n1256), .A2(n1257), .ZN(G42) );
NAND2_X1 U910 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U911 ( .A(KEYINPUT3), .B(G140), .Z(n1258) );
XOR2_X1 U912 ( .A(n1260), .B(KEYINPUT46), .Z(n1256) );
NAND2_X1 U913 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
INV_X1 U914 ( .A(n1259), .ZN(n1262) );
NAND3_X1 U915 ( .A1(n1263), .A2(n1166), .A3(n1264), .ZN(n1259) );
XNOR2_X1 U916 ( .A(n1085), .B(KEYINPUT52), .ZN(n1264) );
XNOR2_X1 U917 ( .A(G140), .B(KEYINPUT18), .ZN(n1261) );
XOR2_X1 U918 ( .A(n1224), .B(n1265), .Z(G39) );
XOR2_X1 U919 ( .A(KEYINPUT38), .B(G137), .Z(n1265) );
NAND3_X1 U920 ( .A1(n1233), .A2(n1069), .A3(n1263), .ZN(n1224) );
INV_X1 U921 ( .A(n1237), .ZN(n1263) );
INV_X1 U922 ( .A(n1251), .ZN(n1233) );
XOR2_X1 U923 ( .A(G134), .B(n1227), .Z(G36) );
NOR3_X1 U924 ( .A1(n1266), .A2(n1049), .A3(n1237), .ZN(n1227) );
XOR2_X1 U925 ( .A(G131), .B(n1229), .Z(G33) );
NOR3_X1 U926 ( .A1(n1266), .A2(n1083), .A3(n1237), .ZN(n1229) );
NAND3_X1 U927 ( .A1(n1066), .A2(n1065), .A3(n1235), .ZN(n1237) );
INV_X1 U928 ( .A(n1250), .ZN(n1235) );
INV_X1 U929 ( .A(n1267), .ZN(n1066) );
XOR2_X1 U930 ( .A(G128), .B(n1228), .Z(G30) );
NOR4_X1 U931 ( .A1(n1250), .A2(n1251), .A3(n1049), .A4(n1241), .ZN(n1228) );
NAND2_X1 U932 ( .A1(n1216), .A2(n1239), .ZN(n1250) );
XNOR2_X1 U933 ( .A(G101), .B(n1207), .ZN(G3) );
NAND3_X1 U934 ( .A1(n1086), .A2(n1216), .A3(n1217), .ZN(n1207) );
INV_X1 U935 ( .A(n1266), .ZN(n1086) );
XNOR2_X1 U936 ( .A(G125), .B(n1268), .ZN(G27) );
NAND4_X1 U937 ( .A1(KEYINPUT24), .A2(n1085), .A3(n1269), .A4(n1166), .ZN(n1268) );
AND2_X1 U938 ( .A1(n1239), .A2(n1091), .ZN(n1269) );
NAND2_X1 U939 ( .A1(n1096), .A2(n1270), .ZN(n1239) );
NAND4_X1 U940 ( .A1(G953), .A2(G902), .A3(n1271), .A4(n1117), .ZN(n1270) );
INV_X1 U941 ( .A(G900), .ZN(n1117) );
XOR2_X1 U942 ( .A(n1206), .B(n1272), .Z(G24) );
NAND2_X1 U943 ( .A1(KEYINPUT17), .A2(G122), .ZN(n1272) );
NAND4_X1 U944 ( .A1(n1273), .A2(n1274), .A3(n1091), .A4(n1275), .ZN(n1206) );
NOR2_X1 U945 ( .A1(n1215), .A2(n1103), .ZN(n1275) );
INV_X1 U946 ( .A(n1077), .ZN(n1103) );
NOR2_X1 U947 ( .A1(n1276), .A2(n1277), .ZN(n1077) );
OR2_X1 U948 ( .A1(n1166), .A2(KEYINPUT23), .ZN(n1274) );
NAND2_X1 U949 ( .A1(KEYINPUT23), .A2(n1278), .ZN(n1273) );
NAND2_X1 U950 ( .A1(n1104), .A2(n1255), .ZN(n1278) );
XNOR2_X1 U951 ( .A(G119), .B(n1219), .ZN(G21) );
NAND2_X1 U952 ( .A1(n1220), .A2(n1279), .ZN(n1219) );
NOR3_X1 U953 ( .A1(n1090), .A2(n1095), .A3(n1251), .ZN(n1220) );
NAND2_X1 U954 ( .A1(n1277), .A2(n1276), .ZN(n1251) );
INV_X1 U955 ( .A(n1280), .ZN(n1277) );
XOR2_X1 U956 ( .A(n1281), .B(n1247), .Z(G18) );
NAND2_X1 U957 ( .A1(n1245), .A2(n1091), .ZN(n1247) );
INV_X1 U958 ( .A(n1095), .ZN(n1091) );
NAND2_X1 U959 ( .A1(n1078), .A2(n1234), .ZN(n1095) );
INV_X1 U960 ( .A(n1241), .ZN(n1234) );
XOR2_X1 U961 ( .A(n1214), .B(KEYINPUT60), .Z(n1241) );
NOR3_X1 U962 ( .A1(n1049), .A2(n1215), .A3(n1266), .ZN(n1245) );
NAND2_X1 U963 ( .A1(n1282), .A2(n1104), .ZN(n1049) );
XOR2_X1 U964 ( .A(G113), .B(n1283), .Z(G15) );
NOR3_X1 U965 ( .A1(n1284), .A2(KEYINPUT56), .A3(n1215), .ZN(n1283) );
INV_X1 U966 ( .A(n1221), .ZN(n1284) );
NOR4_X1 U967 ( .A1(n1266), .A2(n1083), .A3(n1214), .A4(n1244), .ZN(n1221) );
INV_X1 U968 ( .A(n1078), .ZN(n1244) );
NAND2_X1 U969 ( .A1(n1285), .A2(n1286), .ZN(n1078) );
OR3_X1 U970 ( .A1(n1076), .A2(n1075), .A3(KEYINPUT39), .ZN(n1286) );
INV_X1 U971 ( .A(n1287), .ZN(n1075) );
NAND2_X1 U972 ( .A1(KEYINPUT39), .A2(n1216), .ZN(n1285) );
INV_X1 U973 ( .A(n1166), .ZN(n1083) );
NOR2_X1 U974 ( .A1(n1104), .A2(n1282), .ZN(n1166) );
NAND2_X1 U975 ( .A1(n1280), .A2(n1276), .ZN(n1266) );
XNOR2_X1 U976 ( .A(G110), .B(n1288), .ZN(G12) );
NAND3_X1 U977 ( .A1(n1085), .A2(n1217), .A3(n1289), .ZN(n1288) );
XNOR2_X1 U978 ( .A(n1216), .B(KEYINPUT8), .ZN(n1289) );
AND2_X1 U979 ( .A1(n1287), .A2(n1076), .ZN(n1216) );
NAND2_X1 U980 ( .A1(n1290), .A2(n1098), .ZN(n1076) );
NAND2_X1 U981 ( .A1(G469), .A2(n1291), .ZN(n1098) );
XOR2_X1 U982 ( .A(n1099), .B(KEYINPUT14), .Z(n1290) );
OR2_X1 U983 ( .A1(n1291), .A2(G469), .ZN(n1099) );
NAND2_X1 U984 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U985 ( .A(n1294), .B(n1295), .Z(n1292) );
XNOR2_X1 U986 ( .A(n1127), .B(n1197), .ZN(n1295) );
XNOR2_X1 U987 ( .A(n1296), .B(n1297), .ZN(n1197) );
XOR2_X1 U988 ( .A(KEYINPUT6), .B(G107), .Z(n1297) );
XOR2_X1 U989 ( .A(G101), .B(n1298), .Z(n1296) );
XNOR2_X1 U990 ( .A(n1299), .B(n1181), .ZN(n1127) );
XNOR2_X1 U991 ( .A(KEYINPUT61), .B(KEYINPUT54), .ZN(n1299) );
XOR2_X1 U992 ( .A(n1300), .B(n1301), .Z(n1294) );
INV_X1 U993 ( .A(n1196), .ZN(n1301) );
XNOR2_X1 U994 ( .A(G140), .B(n1302), .ZN(n1196) );
NOR2_X1 U995 ( .A1(G953), .A2(n1116), .ZN(n1302) );
INV_X1 U996 ( .A(G227), .ZN(n1116) );
XOR2_X1 U997 ( .A(n1303), .B(G110), .Z(n1300) );
NAND2_X1 U998 ( .A1(KEYINPUT26), .A2(n1190), .ZN(n1303) );
NAND2_X1 U999 ( .A1(G221), .A2(n1304), .ZN(n1287) );
NOR3_X1 U1000 ( .A1(n1214), .A2(n1215), .A3(n1090), .ZN(n1217) );
INV_X1 U1001 ( .A(n1069), .ZN(n1090) );
NOR2_X1 U1002 ( .A1(n1104), .A2(n1255), .ZN(n1069) );
INV_X1 U1003 ( .A(n1282), .ZN(n1255) );
NOR2_X1 U1004 ( .A1(n1108), .A2(n1305), .ZN(n1282) );
AND2_X1 U1005 ( .A1(G475), .A2(n1109), .ZN(n1305) );
NOR2_X1 U1006 ( .A1(n1109), .A2(G475), .ZN(n1108) );
NAND2_X1 U1007 ( .A1(n1159), .A2(n1293), .ZN(n1109) );
XNOR2_X1 U1008 ( .A(n1306), .B(n1307), .ZN(n1159) );
XNOR2_X1 U1009 ( .A(n1308), .B(n1309), .ZN(n1307) );
XOR2_X1 U1010 ( .A(n1310), .B(n1311), .Z(n1309) );
AND2_X1 U1011 ( .A1(n1312), .A2(G214), .ZN(n1311) );
NAND2_X1 U1012 ( .A1(KEYINPUT50), .A2(n1313), .ZN(n1310) );
XNOR2_X1 U1013 ( .A(n1314), .B(n1122), .ZN(n1313) );
XNOR2_X1 U1014 ( .A(G125), .B(G140), .ZN(n1122) );
NOR2_X1 U1015 ( .A1(G146), .A2(KEYINPUT11), .ZN(n1314) );
XOR2_X1 U1016 ( .A(n1315), .B(n1316), .Z(n1306) );
NOR2_X1 U1017 ( .A1(KEYINPUT32), .A2(G143), .ZN(n1316) );
XOR2_X1 U1018 ( .A(G131), .B(n1298), .Z(n1315) );
XNOR2_X1 U1019 ( .A(n1317), .B(G478), .ZN(n1104) );
OR2_X1 U1020 ( .A1(n1156), .A2(G902), .ZN(n1317) );
XNOR2_X1 U1021 ( .A(n1318), .B(n1319), .ZN(n1156) );
XOR2_X1 U1022 ( .A(n1320), .B(n1321), .Z(n1319) );
NAND2_X1 U1023 ( .A1(KEYINPUT29), .A2(n1322), .ZN(n1321) );
NAND2_X1 U1024 ( .A1(n1323), .A2(n1324), .ZN(n1320) );
OR2_X1 U1025 ( .A1(n1325), .A2(G134), .ZN(n1324) );
XOR2_X1 U1026 ( .A(n1326), .B(KEYINPUT0), .Z(n1323) );
NAND2_X1 U1027 ( .A1(G134), .A2(n1325), .ZN(n1326) );
XOR2_X1 U1028 ( .A(n1327), .B(n1328), .Z(n1318) );
XOR2_X1 U1029 ( .A(G116), .B(G107), .Z(n1328) );
NAND2_X1 U1030 ( .A1(G217), .A2(n1329), .ZN(n1327) );
INV_X1 U1031 ( .A(n1279), .ZN(n1215) );
NAND2_X1 U1032 ( .A1(n1096), .A2(n1330), .ZN(n1279) );
NAND4_X1 U1033 ( .A1(n1331), .A2(G953), .A3(G902), .A4(n1271), .ZN(n1330) );
XNOR2_X1 U1034 ( .A(G898), .B(KEYINPUT9), .ZN(n1331) );
NAND3_X1 U1035 ( .A1(n1271), .A2(n1058), .A3(G952), .ZN(n1096) );
NAND2_X1 U1036 ( .A1(G237), .A2(G234), .ZN(n1271) );
NAND2_X1 U1037 ( .A1(n1267), .A2(n1065), .ZN(n1214) );
NAND2_X1 U1038 ( .A1(G214), .A2(n1332), .ZN(n1065) );
NAND3_X1 U1039 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1267) );
INV_X1 U1040 ( .A(n1112), .ZN(n1335) );
NOR2_X1 U1041 ( .A1(n1111), .A2(n1110), .ZN(n1112) );
NAND2_X1 U1042 ( .A1(KEYINPUT31), .A2(n1203), .ZN(n1334) );
NAND3_X1 U1043 ( .A1(n1111), .A2(n1336), .A3(n1110), .ZN(n1333) );
INV_X1 U1044 ( .A(n1203), .ZN(n1110) );
NAND2_X1 U1045 ( .A1(G210), .A2(n1332), .ZN(n1203) );
NAND2_X1 U1046 ( .A1(n1337), .A2(n1293), .ZN(n1332) );
INV_X1 U1047 ( .A(G237), .ZN(n1337) );
INV_X1 U1048 ( .A(KEYINPUT31), .ZN(n1336) );
NAND2_X1 U1049 ( .A1(n1201), .A2(n1293), .ZN(n1111) );
XNOR2_X1 U1050 ( .A(n1338), .B(n1339), .ZN(n1201) );
XOR2_X1 U1051 ( .A(n1340), .B(n1341), .Z(n1339) );
AND2_X1 U1052 ( .A1(n1058), .A2(G224), .ZN(n1340) );
XNOR2_X1 U1053 ( .A(n1342), .B(n1145), .ZN(n1338) );
XNOR2_X1 U1054 ( .A(n1343), .B(n1344), .ZN(n1145) );
XOR2_X1 U1055 ( .A(n1345), .B(n1346), .Z(n1344) );
XOR2_X1 U1056 ( .A(n1347), .B(KEYINPUT21), .Z(n1346) );
NAND3_X1 U1057 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1347) );
OR2_X1 U1058 ( .A1(n1298), .A2(KEYINPUT20), .ZN(n1350) );
NAND3_X1 U1059 ( .A1(KEYINPUT20), .A2(n1298), .A3(G107), .ZN(n1349) );
INV_X1 U1060 ( .A(G104), .ZN(n1298) );
NAND2_X1 U1061 ( .A1(n1351), .A2(n1352), .ZN(n1348) );
INV_X1 U1062 ( .A(G107), .ZN(n1352) );
NAND2_X1 U1063 ( .A1(KEYINPUT20), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1064 ( .A(KEYINPUT45), .B(G104), .Z(n1353) );
NAND2_X1 U1065 ( .A1(KEYINPUT55), .A2(n1354), .ZN(n1345) );
XOR2_X1 U1066 ( .A(KEYINPUT48), .B(G101), .Z(n1354) );
XOR2_X1 U1067 ( .A(n1355), .B(n1308), .Z(n1343) );
XNOR2_X1 U1068 ( .A(n1322), .B(G113), .ZN(n1308) );
INV_X1 U1069 ( .A(G122), .ZN(n1322) );
NOR2_X1 U1070 ( .A1(n1276), .A2(n1280), .ZN(n1085) );
XNOR2_X1 U1071 ( .A(n1356), .B(n1152), .ZN(n1280) );
NAND2_X1 U1072 ( .A1(G217), .A2(n1304), .ZN(n1152) );
NAND2_X1 U1073 ( .A1(G234), .A2(n1293), .ZN(n1304) );
NAND2_X1 U1074 ( .A1(n1151), .A2(n1293), .ZN(n1356) );
XOR2_X1 U1075 ( .A(n1357), .B(n1358), .Z(n1151) );
XOR2_X1 U1076 ( .A(n1342), .B(n1359), .Z(n1358) );
XNOR2_X1 U1077 ( .A(n1360), .B(n1361), .ZN(n1359) );
NOR2_X1 U1078 ( .A1(G140), .A2(KEYINPUT19), .ZN(n1361) );
NAND2_X1 U1079 ( .A1(KEYINPUT25), .A2(G146), .ZN(n1360) );
XOR2_X1 U1080 ( .A(G125), .B(G110), .Z(n1342) );
XOR2_X1 U1081 ( .A(n1362), .B(n1363), .Z(n1357) );
XOR2_X1 U1082 ( .A(G137), .B(G128), .Z(n1363) );
XOR2_X1 U1083 ( .A(n1364), .B(G119), .Z(n1362) );
NAND3_X1 U1084 ( .A1(KEYINPUT40), .A2(n1329), .A3(n1365), .ZN(n1364) );
XNOR2_X1 U1085 ( .A(G221), .B(KEYINPUT33), .ZN(n1365) );
AND2_X1 U1086 ( .A1(G234), .A2(n1058), .ZN(n1329) );
INV_X1 U1087 ( .A(G953), .ZN(n1058) );
XNOR2_X1 U1088 ( .A(n1366), .B(G472), .ZN(n1276) );
NAND2_X1 U1089 ( .A1(n1367), .A2(n1293), .ZN(n1366) );
INV_X1 U1090 ( .A(G902), .ZN(n1293) );
XOR2_X1 U1091 ( .A(n1368), .B(n1171), .Z(n1367) );
XOR2_X1 U1092 ( .A(n1369), .B(G101), .Z(n1171) );
NAND2_X1 U1093 ( .A1(G210), .A2(n1312), .ZN(n1369) );
NOR2_X1 U1094 ( .A1(G953), .A2(G237), .ZN(n1312) );
NAND4_X1 U1095 ( .A1(n1370), .A2(n1176), .A3(n1371), .A4(n1372), .ZN(n1368) );
NAND3_X1 U1096 ( .A1(n1373), .A2(n1374), .A3(n1341), .ZN(n1372) );
NAND3_X1 U1097 ( .A1(n1375), .A2(n1180), .A3(n1181), .ZN(n1371) );
NAND2_X1 U1098 ( .A1(KEYINPUT62), .A2(n1190), .ZN(n1375) );
NAND3_X1 U1099 ( .A1(n1179), .A2(n1341), .A3(n1373), .ZN(n1176) );
INV_X1 U1100 ( .A(n1180), .ZN(n1373) );
INV_X1 U1101 ( .A(n1190), .ZN(n1179) );
OR2_X1 U1102 ( .A1(n1177), .A2(n1374), .ZN(n1370) );
INV_X1 U1103 ( .A(KEYINPUT62), .ZN(n1374) );
NAND2_X1 U1104 ( .A1(n1190), .A2(n1376), .ZN(n1177) );
XOR2_X1 U1105 ( .A(n1180), .B(n1181), .Z(n1376) );
INV_X1 U1106 ( .A(n1341), .ZN(n1181) );
XOR2_X1 U1107 ( .A(G146), .B(n1325), .Z(n1341) );
XOR2_X1 U1108 ( .A(G128), .B(G143), .Z(n1325) );
NAND2_X1 U1109 ( .A1(n1377), .A2(n1378), .ZN(n1180) );
NAND2_X1 U1110 ( .A1(n1355), .A2(n1379), .ZN(n1378) );
XOR2_X1 U1111 ( .A(KEYINPUT1), .B(n1380), .Z(n1377) );
NOR2_X1 U1112 ( .A1(n1355), .A2(n1379), .ZN(n1380) );
INV_X1 U1113 ( .A(G113), .ZN(n1379) );
XOR2_X1 U1114 ( .A(n1281), .B(G119), .Z(n1355) );
INV_X1 U1115 ( .A(G116), .ZN(n1281) );
XOR2_X1 U1116 ( .A(n1381), .B(n1382), .Z(n1190) );
NOR2_X1 U1117 ( .A1(KEYINPUT58), .A2(G134), .ZN(n1382) );
XOR2_X1 U1118 ( .A(G131), .B(n1133), .Z(n1381) );
INV_X1 U1119 ( .A(G137), .ZN(n1133) );
endmodule


