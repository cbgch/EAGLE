//Key = 0101110110011011111111010010110011000110110000110111001101110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399;

XOR2_X1 U757 ( .A(n1053), .B(n1054), .Z(G9) );
XOR2_X1 U758 ( .A(KEYINPUT36), .B(G107), .Z(n1054) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(G75) );
XOR2_X1 U761 ( .A(KEYINPUT25), .B(n1059), .Z(n1058) );
NOR3_X1 U762 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U764 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U766 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR3_X1 U768 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1071) );
NOR2_X1 U769 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR3_X1 U772 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1074) );
XNOR2_X1 U773 ( .A(KEYINPUT51), .B(n1085), .ZN(n1082) );
AND2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1073) );
NOR3_X1 U775 ( .A1(n1085), .A2(n1088), .A3(n1077), .ZN(n1069) );
NOR2_X1 U776 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
AND2_X1 U777 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NOR4_X1 U778 ( .A1(n1093), .A2(n1094), .A3(n1077), .A4(n1085), .ZN(n1065) );
NOR3_X1 U779 ( .A1(n1072), .A2(n1095), .A3(n1096), .ZN(n1094) );
NOR2_X1 U780 ( .A1(KEYINPUT22), .A2(n1097), .ZN(n1096) );
NOR2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1093) );
AND2_X1 U782 ( .A1(n1100), .A2(KEYINPUT22), .ZN(n1099) );
NOR2_X1 U783 ( .A1(G952), .A2(n1062), .ZN(n1057) );
NAND2_X1 U784 ( .A1(n1101), .A2(n1102), .ZN(n1062) );
NAND4_X1 U785 ( .A1(n1091), .A2(n1103), .A3(n1086), .A4(n1104), .ZN(n1102) );
NOR4_X1 U786 ( .A1(n1105), .A2(n1106), .A3(n1092), .A4(n1107), .ZN(n1104) );
XOR2_X1 U787 ( .A(n1108), .B(n1109), .Z(n1107) );
XNOR2_X1 U788 ( .A(KEYINPUT17), .B(n1110), .ZN(n1109) );
INV_X1 U789 ( .A(n1111), .ZN(n1106) );
NAND2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(G72) );
NAND2_X1 U791 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U792 ( .A(KEYINPUT18), .B(n1116), .Z(n1112) );
NOR2_X1 U793 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U794 ( .A(n1114), .B(KEYINPUT11), .ZN(n1118) );
AND2_X1 U795 ( .A1(G953), .A2(n1119), .ZN(n1114) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1119) );
NOR2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
INV_X1 U798 ( .A(n1115), .ZN(n1121) );
NAND3_X1 U799 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1115) );
XOR2_X1 U800 ( .A(n1125), .B(KEYINPUT45), .Z(n1124) );
NAND2_X1 U801 ( .A1(n1101), .A2(n1126), .ZN(n1125) );
OR2_X1 U802 ( .A1(n1101), .A2(G900), .ZN(n1123) );
NOR3_X1 U803 ( .A1(n1127), .A2(G953), .A3(n1122), .ZN(n1120) );
AND2_X1 U804 ( .A1(n1128), .A2(n1129), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U806 ( .A(KEYINPUT3), .B(n1132), .Z(n1128) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1132) );
XOR2_X1 U808 ( .A(n1133), .B(n1134), .Z(n1131) );
NOR2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NOR2_X1 U810 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U811 ( .A(G131), .B(KEYINPUT31), .ZN(n1138) );
INV_X1 U812 ( .A(n1139), .ZN(n1137) );
INV_X1 U813 ( .A(n1140), .ZN(n1130) );
NAND3_X1 U814 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(G69) );
XOR2_X1 U815 ( .A(n1144), .B(KEYINPUT43), .Z(n1143) );
NAND2_X1 U816 ( .A1(G953), .A2(n1145), .ZN(n1144) );
NAND2_X1 U817 ( .A1(G898), .A2(n1146), .ZN(n1145) );
NAND2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U819 ( .A1(n1149), .A2(n1101), .ZN(n1142) );
XNOR2_X1 U820 ( .A(n1150), .B(n1147), .ZN(n1149) );
NAND2_X1 U821 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U822 ( .A(n1153), .B(KEYINPUT13), .Z(n1151) );
NAND4_X1 U823 ( .A1(G224), .A2(n1154), .A3(G898), .A4(G953), .ZN(n1141) );
NOR2_X1 U824 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XOR2_X1 U825 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U826 ( .A1(KEYINPUT0), .A2(n1159), .ZN(n1158) );
OR2_X1 U827 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1162), .ZN(G63) );
XOR2_X1 U829 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND3_X1 U830 ( .A1(n1165), .A2(n1166), .A3(G478), .ZN(n1163) );
NAND2_X1 U831 ( .A1(KEYINPUT47), .A2(n1160), .ZN(n1166) );
NAND2_X1 U832 ( .A1(n1167), .A2(n1168), .ZN(n1165) );
INV_X1 U833 ( .A(KEYINPUT47), .ZN(n1168) );
OR2_X1 U834 ( .A1(n1060), .A2(n1169), .ZN(n1167) );
NOR3_X1 U835 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(G60) );
AND3_X1 U836 ( .A1(KEYINPUT48), .A2(n1101), .A3(n1173), .ZN(n1172) );
NOR2_X1 U837 ( .A1(KEYINPUT48), .A2(n1174), .ZN(n1171) );
INV_X1 U838 ( .A(n1155), .ZN(n1174) );
XOR2_X1 U839 ( .A(n1175), .B(n1176), .Z(n1170) );
NOR2_X1 U840 ( .A1(n1177), .A2(n1160), .ZN(n1176) );
XNOR2_X1 U841 ( .A(G104), .B(n1178), .ZN(G6) );
NAND2_X1 U842 ( .A1(n1179), .A2(n1079), .ZN(n1178) );
XOR2_X1 U843 ( .A(n1180), .B(KEYINPUT1), .Z(n1179) );
NOR2_X1 U844 ( .A1(n1155), .A2(n1181), .ZN(G57) );
XOR2_X1 U845 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U846 ( .A(KEYINPUT56), .B(KEYINPUT19), .Z(n1183) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(n1182) );
NOR2_X1 U848 ( .A1(n1110), .A2(n1160), .ZN(n1185) );
NOR3_X1 U849 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(G54) );
AND2_X1 U850 ( .A1(n1155), .A2(KEYINPUT58), .ZN(n1188) );
NOR3_X1 U851 ( .A1(KEYINPUT58), .A2(n1101), .A3(n1173), .ZN(n1187) );
INV_X1 U852 ( .A(G952), .ZN(n1173) );
XOR2_X1 U853 ( .A(n1189), .B(n1190), .Z(n1186) );
XOR2_X1 U854 ( .A(n1191), .B(n1192), .Z(n1190) );
NOR2_X1 U855 ( .A1(n1193), .A2(n1160), .ZN(n1191) );
XOR2_X1 U856 ( .A(n1194), .B(n1195), .Z(n1189) );
XOR2_X1 U857 ( .A(n1133), .B(n1196), .Z(n1195) );
NAND2_X1 U858 ( .A1(KEYINPUT49), .A2(n1197), .ZN(n1194) );
XNOR2_X1 U859 ( .A(n1198), .B(n1199), .ZN(n1197) );
NAND2_X1 U860 ( .A1(KEYINPUT26), .A2(n1200), .ZN(n1198) );
XNOR2_X1 U861 ( .A(KEYINPUT7), .B(n1201), .ZN(n1200) );
NOR2_X1 U862 ( .A1(n1155), .A2(n1202), .ZN(G51) );
XOR2_X1 U863 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U864 ( .A1(n1205), .A2(n1160), .ZN(n1204) );
NAND2_X1 U865 ( .A1(G902), .A2(n1060), .ZN(n1160) );
NAND3_X1 U866 ( .A1(n1152), .A2(n1153), .A3(n1127), .ZN(n1060) );
INV_X1 U867 ( .A(n1126), .ZN(n1127) );
NAND4_X1 U868 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1126) );
AND4_X1 U869 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1209) );
NAND2_X1 U870 ( .A1(n1087), .A2(n1214), .ZN(n1208) );
NAND2_X1 U871 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND3_X1 U872 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1216) );
NAND2_X1 U873 ( .A1(n1220), .A2(n1100), .ZN(n1215) );
NAND3_X1 U874 ( .A1(n1221), .A2(n1079), .A3(n1222), .ZN(n1153) );
XOR2_X1 U875 ( .A(n1223), .B(KEYINPUT9), .Z(n1222) );
INV_X1 U876 ( .A(n1055), .ZN(n1221) );
NAND3_X1 U877 ( .A1(n1224), .A2(n1095), .A3(n1090), .ZN(n1055) );
AND4_X1 U878 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1152) );
NOR3_X1 U879 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1228) );
NOR2_X1 U880 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NOR2_X1 U881 ( .A1(n1095), .A2(n1100), .ZN(n1232) );
NOR2_X1 U882 ( .A1(n1234), .A2(n1180), .ZN(n1229) );
NAND4_X1 U883 ( .A1(n1100), .A2(n1090), .A3(n1224), .A4(n1223), .ZN(n1180) );
XOR2_X1 U884 ( .A(n1235), .B(n1236), .Z(n1203) );
NOR2_X1 U885 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U886 ( .A(n1239), .B(KEYINPUT5), .ZN(n1238) );
NAND2_X1 U887 ( .A1(KEYINPUT21), .A2(n1154), .ZN(n1235) );
NOR2_X1 U888 ( .A1(n1101), .A2(G952), .ZN(n1155) );
XOR2_X1 U889 ( .A(n1206), .B(n1240), .Z(G48) );
NAND2_X1 U890 ( .A1(KEYINPUT57), .A2(G146), .ZN(n1240) );
NAND4_X1 U891 ( .A1(n1100), .A2(n1219), .A3(n1084), .A4(n1241), .ZN(n1206) );
XNOR2_X1 U892 ( .A(G143), .B(n1242), .ZN(G45) );
NAND3_X1 U893 ( .A1(KEYINPUT37), .A2(n1087), .A3(n1243), .ZN(n1242) );
NOR3_X1 U894 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
XNOR2_X1 U895 ( .A(G140), .B(n1207), .ZN(G42) );
NAND2_X1 U896 ( .A1(n1220), .A2(n1247), .ZN(n1207) );
XNOR2_X1 U897 ( .A(G137), .B(n1213), .ZN(G39) );
NAND4_X1 U898 ( .A1(n1084), .A2(n1220), .A3(n1103), .A4(n1241), .ZN(n1213) );
XNOR2_X1 U899 ( .A(G134), .B(n1212), .ZN(G36) );
NAND3_X1 U900 ( .A1(n1220), .A2(n1095), .A3(n1087), .ZN(n1212) );
XNOR2_X1 U901 ( .A(G131), .B(n1248), .ZN(G33) );
NAND4_X1 U902 ( .A1(KEYINPUT32), .A2(n1087), .A3(n1220), .A4(n1100), .ZN(n1248) );
AND3_X1 U903 ( .A1(n1090), .A2(n1249), .A3(n1086), .ZN(n1220) );
INV_X1 U904 ( .A(n1085), .ZN(n1086) );
NAND2_X1 U905 ( .A1(n1250), .A2(n1081), .ZN(n1085) );
INV_X1 U906 ( .A(n1080), .ZN(n1250) );
XNOR2_X1 U907 ( .A(G128), .B(n1210), .ZN(G30) );
NAND4_X1 U908 ( .A1(n1084), .A2(n1219), .A3(n1095), .A4(n1241), .ZN(n1210) );
INV_X1 U909 ( .A(n1244), .ZN(n1219) );
NAND2_X1 U910 ( .A1(n1251), .A2(n1090), .ZN(n1244) );
XNOR2_X1 U911 ( .A(G101), .B(n1226), .ZN(G3) );
NAND4_X1 U912 ( .A1(n1087), .A2(n1103), .A3(n1252), .A4(n1090), .ZN(n1226) );
XNOR2_X1 U913 ( .A(G125), .B(n1211), .ZN(G27) );
NAND3_X1 U914 ( .A1(n1247), .A2(n1251), .A3(n1098), .ZN(n1211) );
AND2_X1 U915 ( .A1(n1079), .A2(n1249), .ZN(n1251) );
NAND2_X1 U916 ( .A1(n1064), .A2(n1253), .ZN(n1249) );
NAND4_X1 U917 ( .A1(n1254), .A2(G953), .A3(G902), .A4(n1255), .ZN(n1253) );
XNOR2_X1 U918 ( .A(G900), .B(KEYINPUT62), .ZN(n1254) );
NOR3_X1 U919 ( .A1(n1084), .A2(n1083), .A3(n1097), .ZN(n1247) );
XOR2_X1 U920 ( .A(G122), .B(n1230), .Z(G24) );
AND3_X1 U921 ( .A1(n1098), .A2(n1252), .A3(n1256), .ZN(n1230) );
NOR3_X1 U922 ( .A1(n1077), .A2(n1245), .A3(n1246), .ZN(n1256) );
INV_X1 U923 ( .A(n1224), .ZN(n1077) );
NOR2_X1 U924 ( .A1(n1241), .A2(n1084), .ZN(n1224) );
XNOR2_X1 U925 ( .A(G119), .B(n1227), .ZN(G21) );
NAND3_X1 U926 ( .A1(n1084), .A2(n1098), .A3(n1257), .ZN(n1227) );
INV_X1 U927 ( .A(n1258), .ZN(n1084) );
XOR2_X1 U928 ( .A(G116), .B(n1259), .Z(G18) );
NOR2_X1 U929 ( .A1(n1260), .A2(n1233), .ZN(n1259) );
INV_X1 U930 ( .A(n1095), .ZN(n1260) );
NOR2_X1 U931 ( .A1(n1218), .A2(n1246), .ZN(n1095) );
INV_X1 U932 ( .A(n1217), .ZN(n1246) );
XOR2_X1 U933 ( .A(G113), .B(n1261), .Z(G15) );
NOR2_X1 U934 ( .A1(n1233), .A2(n1262), .ZN(n1261) );
XNOR2_X1 U935 ( .A(KEYINPUT59), .B(n1097), .ZN(n1262) );
INV_X1 U936 ( .A(n1100), .ZN(n1097) );
NOR2_X1 U937 ( .A1(n1217), .A2(n1245), .ZN(n1100) );
NAND3_X1 U938 ( .A1(n1098), .A2(n1252), .A3(n1087), .ZN(n1233) );
NOR2_X1 U939 ( .A1(n1258), .A2(n1241), .ZN(n1087) );
INV_X1 U940 ( .A(n1056), .ZN(n1252) );
INV_X1 U941 ( .A(n1072), .ZN(n1098) );
NAND2_X1 U942 ( .A1(n1091), .A2(n1263), .ZN(n1072) );
XOR2_X1 U943 ( .A(KEYINPUT38), .B(n1092), .Z(n1263) );
NAND2_X1 U944 ( .A1(n1264), .A2(n1265), .ZN(G12) );
NAND2_X1 U945 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
INV_X1 U946 ( .A(G110), .ZN(n1267) );
XNOR2_X1 U947 ( .A(KEYINPUT52), .B(n1225), .ZN(n1266) );
NAND2_X1 U948 ( .A1(G110), .A2(n1268), .ZN(n1264) );
XOR2_X1 U949 ( .A(n1225), .B(KEYINPUT27), .Z(n1268) );
NAND3_X1 U950 ( .A1(n1090), .A2(n1258), .A3(n1257), .ZN(n1225) );
NOR3_X1 U951 ( .A1(n1056), .A2(n1083), .A3(n1068), .ZN(n1257) );
INV_X1 U952 ( .A(n1103), .ZN(n1068) );
NOR2_X1 U953 ( .A1(n1217), .A2(n1218), .ZN(n1103) );
INV_X1 U954 ( .A(n1245), .ZN(n1218) );
XOR2_X1 U955 ( .A(n1177), .B(n1269), .Z(n1245) );
NOR2_X1 U956 ( .A1(G902), .A2(n1175), .ZN(n1269) );
NAND3_X1 U957 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1175) );
OR2_X1 U958 ( .A1(n1273), .A2(KEYINPUT12), .ZN(n1272) );
NAND3_X1 U959 ( .A1(KEYINPUT12), .A2(n1274), .A3(n1275), .ZN(n1271) );
OR2_X1 U960 ( .A1(n1275), .A2(n1274), .ZN(n1270) );
AND2_X1 U961 ( .A1(KEYINPUT20), .A2(n1273), .ZN(n1274) );
XNOR2_X1 U962 ( .A(n1276), .B(n1277), .ZN(n1273) );
XOR2_X1 U963 ( .A(KEYINPUT33), .B(G122), .Z(n1277) );
XNOR2_X1 U964 ( .A(G104), .B(G113), .ZN(n1276) );
XNOR2_X1 U965 ( .A(n1278), .B(n1279), .ZN(n1275) );
XNOR2_X1 U966 ( .A(G131), .B(n1280), .ZN(n1279) );
NAND2_X1 U967 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U968 ( .A1(G146), .A2(n1140), .ZN(n1282) );
XOR2_X1 U969 ( .A(KEYINPUT28), .B(n1283), .Z(n1281) );
NOR2_X1 U970 ( .A1(G146), .A2(n1140), .ZN(n1283) );
NAND2_X1 U971 ( .A1(n1284), .A2(KEYINPUT61), .ZN(n1278) );
XNOR2_X1 U972 ( .A(G143), .B(n1285), .ZN(n1284) );
NOR3_X1 U973 ( .A1(n1286), .A2(G953), .A3(G237), .ZN(n1285) );
INV_X1 U974 ( .A(G214), .ZN(n1286) );
INV_X1 U975 ( .A(G475), .ZN(n1177) );
XNOR2_X1 U976 ( .A(n1287), .B(G478), .ZN(n1217) );
NAND2_X1 U977 ( .A1(n1288), .A2(n1164), .ZN(n1287) );
XNOR2_X1 U978 ( .A(n1289), .B(n1290), .ZN(n1164) );
XNOR2_X1 U979 ( .A(n1291), .B(n1292), .ZN(n1290) );
NOR2_X1 U980 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U981 ( .A(n1295), .B(KEYINPUT40), .Z(n1294) );
NAND2_X1 U982 ( .A1(G107), .A2(n1296), .ZN(n1295) );
NOR2_X1 U983 ( .A1(G107), .A2(n1296), .ZN(n1293) );
XOR2_X1 U984 ( .A(G122), .B(n1297), .Z(n1296) );
INV_X1 U985 ( .A(G134), .ZN(n1291) );
XOR2_X1 U986 ( .A(n1298), .B(n1299), .Z(n1289) );
NAND2_X1 U987 ( .A1(n1300), .A2(G217), .ZN(n1298) );
XNOR2_X1 U988 ( .A(KEYINPUT16), .B(n1169), .ZN(n1288) );
INV_X1 U989 ( .A(n1241), .ZN(n1083) );
NAND2_X1 U990 ( .A1(n1301), .A2(n1111), .ZN(n1241) );
NAND2_X1 U991 ( .A1(n1302), .A2(n1161), .ZN(n1111) );
XNOR2_X1 U992 ( .A(n1105), .B(KEYINPUT24), .ZN(n1301) );
NOR2_X1 U993 ( .A1(n1161), .A2(n1302), .ZN(n1105) );
NOR2_X1 U994 ( .A1(n1159), .A2(G902), .ZN(n1302) );
XOR2_X1 U995 ( .A(n1303), .B(n1304), .Z(n1159) );
XOR2_X1 U996 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U997 ( .A(n1307), .B(G137), .ZN(n1306) );
NOR2_X1 U998 ( .A1(KEYINPUT6), .A2(n1308), .ZN(n1305) );
XNOR2_X1 U999 ( .A(G119), .B(G128), .ZN(n1308) );
XNOR2_X1 U1000 ( .A(n1309), .B(n1201), .ZN(n1303) );
XNOR2_X1 U1001 ( .A(n1140), .B(n1310), .ZN(n1309) );
AND2_X1 U1002 ( .A1(G221), .A2(n1300), .ZN(n1310) );
AND2_X1 U1003 ( .A1(G234), .A2(n1101), .ZN(n1300) );
XNOR2_X1 U1004 ( .A(G125), .B(n1311), .ZN(n1140) );
INV_X1 U1005 ( .A(n1199), .ZN(n1311) );
NAND2_X1 U1006 ( .A1(G217), .A2(n1312), .ZN(n1161) );
NAND2_X1 U1007 ( .A1(n1079), .A2(n1223), .ZN(n1056) );
NAND2_X1 U1008 ( .A1(n1064), .A2(n1313), .ZN(n1223) );
NAND4_X1 U1009 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1314), .ZN(n1313) );
INV_X1 U1010 ( .A(G898), .ZN(n1314) );
NAND3_X1 U1011 ( .A1(n1255), .A2(n1101), .A3(G952), .ZN(n1064) );
NAND2_X1 U1012 ( .A1(G234), .A2(G237), .ZN(n1255) );
INV_X1 U1013 ( .A(n1234), .ZN(n1079) );
NAND2_X1 U1014 ( .A1(n1080), .A2(n1081), .ZN(n1234) );
NAND2_X1 U1015 ( .A1(G214), .A2(n1315), .ZN(n1081) );
XOR2_X1 U1016 ( .A(n1316), .B(n1205), .Z(n1080) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1315), .ZN(n1205) );
NAND2_X1 U1018 ( .A1(n1317), .A2(n1169), .ZN(n1315) );
XNOR2_X1 U1019 ( .A(G237), .B(KEYINPUT60), .ZN(n1317) );
NAND2_X1 U1020 ( .A1(n1318), .A2(n1169), .ZN(n1316) );
XNOR2_X1 U1021 ( .A(n1319), .B(n1147), .ZN(n1318) );
INV_X1 U1022 ( .A(n1154), .ZN(n1147) );
XNOR2_X1 U1023 ( .A(n1320), .B(n1321), .ZN(n1154) );
XOR2_X1 U1024 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1025 ( .A(n1324), .B(n1201), .ZN(n1323) );
NAND2_X1 U1026 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1027 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1028 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1029 ( .A1(KEYINPUT35), .A2(n1331), .ZN(n1330) );
NAND3_X1 U1030 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1325) );
INV_X1 U1031 ( .A(KEYINPUT35), .ZN(n1334) );
NAND2_X1 U1032 ( .A1(G119), .A2(n1331), .ZN(n1333) );
NAND2_X1 U1033 ( .A1(n1335), .A2(n1329), .ZN(n1332) );
NAND2_X1 U1034 ( .A1(n1336), .A2(n1331), .ZN(n1335) );
INV_X1 U1035 ( .A(KEYINPUT2), .ZN(n1331) );
XNOR2_X1 U1036 ( .A(G101), .B(n1337), .ZN(n1320) );
XOR2_X1 U1037 ( .A(G122), .B(G113), .Z(n1337) );
NOR3_X1 U1038 ( .A1(n1239), .A2(KEYINPUT53), .A3(n1237), .ZN(n1319) );
NOR3_X1 U1039 ( .A1(n1338), .A2(G953), .A3(n1148), .ZN(n1237) );
INV_X1 U1040 ( .A(G224), .ZN(n1148) );
AND2_X1 U1041 ( .A1(n1338), .A2(n1339), .ZN(n1239) );
NAND2_X1 U1042 ( .A1(G224), .A2(n1101), .ZN(n1339) );
XNOR2_X1 U1043 ( .A(n1340), .B(n1341), .ZN(n1338) );
INV_X1 U1044 ( .A(G125), .ZN(n1341) );
XOR2_X1 U1045 ( .A(n1342), .B(n1110), .Z(n1258) );
INV_X1 U1046 ( .A(G472), .ZN(n1110) );
NAND2_X1 U1047 ( .A1(KEYINPUT14), .A2(n1108), .ZN(n1342) );
NAND2_X1 U1048 ( .A1(n1343), .A2(n1169), .ZN(n1108) );
XOR2_X1 U1049 ( .A(n1184), .B(KEYINPUT44), .Z(n1343) );
XOR2_X1 U1050 ( .A(n1344), .B(n1345), .Z(n1184) );
XOR2_X1 U1051 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1052 ( .A(n1348), .B(n1349), .ZN(n1347) );
XNOR2_X1 U1053 ( .A(n1329), .B(G113), .ZN(n1346) );
INV_X1 U1054 ( .A(G119), .ZN(n1329) );
XNOR2_X1 U1055 ( .A(n1350), .B(n1351), .ZN(n1344) );
INV_X1 U1056 ( .A(n1340), .ZN(n1351) );
XOR2_X1 U1057 ( .A(G146), .B(n1299), .Z(n1340) );
XNOR2_X1 U1058 ( .A(n1352), .B(G143), .ZN(n1299) );
XNOR2_X1 U1059 ( .A(n1353), .B(n1336), .ZN(n1350) );
INV_X1 U1060 ( .A(n1327), .ZN(n1336) );
XOR2_X1 U1061 ( .A(n1297), .B(KEYINPUT4), .Z(n1327) );
XOR2_X1 U1062 ( .A(G116), .B(KEYINPUT63), .Z(n1297) );
NAND3_X1 U1063 ( .A1(n1354), .A2(n1101), .A3(G210), .ZN(n1353) );
XOR2_X1 U1064 ( .A(KEYINPUT23), .B(G237), .Z(n1354) );
NOR2_X1 U1065 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
AND2_X1 U1066 ( .A1(G221), .A2(n1312), .ZN(n1092) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1355), .ZN(n1312) );
XNOR2_X1 U1068 ( .A(KEYINPUT54), .B(n1169), .ZN(n1355) );
XNOR2_X1 U1069 ( .A(n1356), .B(n1193), .ZN(n1091) );
INV_X1 U1070 ( .A(G469), .ZN(n1193) );
NAND3_X1 U1071 ( .A1(n1357), .A2(n1358), .A3(n1169), .ZN(n1356) );
INV_X1 U1072 ( .A(G902), .ZN(n1169) );
NAND2_X1 U1073 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
INV_X1 U1074 ( .A(KEYINPUT42), .ZN(n1360) );
XOR2_X1 U1075 ( .A(n1361), .B(n1362), .Z(n1359) );
NAND2_X1 U1076 ( .A1(n1363), .A2(n1364), .ZN(n1361) );
INV_X1 U1077 ( .A(KEYINPUT39), .ZN(n1364) );
NAND3_X1 U1078 ( .A1(n1365), .A2(n1363), .A3(KEYINPUT42), .ZN(n1357) );
XNOR2_X1 U1079 ( .A(n1192), .B(n1366), .ZN(n1363) );
XNOR2_X1 U1080 ( .A(n1367), .B(KEYINPUT8), .ZN(n1366) );
NAND2_X1 U1081 ( .A1(KEYINPUT29), .A2(n1133), .ZN(n1367) );
AND3_X1 U1082 ( .A1(n1368), .A2(n1369), .A3(n1370), .ZN(n1133) );
NAND3_X1 U1083 ( .A1(n1371), .A2(n1307), .A3(n1372), .ZN(n1370) );
XNOR2_X1 U1084 ( .A(KEYINPUT46), .B(G128), .ZN(n1372) );
INV_X1 U1085 ( .A(G146), .ZN(n1307) );
XNOR2_X1 U1086 ( .A(KEYINPUT30), .B(n1373), .ZN(n1371) );
NAND4_X1 U1087 ( .A1(G146), .A2(n1373), .A3(KEYINPUT46), .A4(G128), .ZN(n1369) );
NAND2_X1 U1088 ( .A1(n1374), .A2(n1352), .ZN(n1368) );
INV_X1 U1089 ( .A(G128), .ZN(n1352) );
NAND3_X1 U1090 ( .A1(n1375), .A2(n1376), .A3(n1377), .ZN(n1374) );
NAND2_X1 U1091 ( .A1(KEYINPUT30), .A2(G143), .ZN(n1377) );
OR3_X1 U1092 ( .A1(G143), .A2(KEYINPUT30), .A3(G146), .ZN(n1376) );
NAND2_X1 U1093 ( .A1(G146), .A2(n1378), .ZN(n1375) );
NAND2_X1 U1094 ( .A1(KEYINPUT46), .A2(n1373), .ZN(n1378) );
INV_X1 U1095 ( .A(G143), .ZN(n1373) );
XNOR2_X1 U1096 ( .A(n1379), .B(n1349), .ZN(n1192) );
NOR2_X1 U1097 ( .A1(n1380), .A2(n1135), .ZN(n1349) );
NOR2_X1 U1098 ( .A1(n1139), .A2(G131), .ZN(n1135) );
AND2_X1 U1099 ( .A1(G131), .A2(n1139), .ZN(n1380) );
XOR2_X1 U1100 ( .A(G134), .B(G137), .Z(n1139) );
NAND3_X1 U1101 ( .A1(n1381), .A2(n1382), .A3(n1383), .ZN(n1379) );
NAND2_X1 U1102 ( .A1(n1384), .A2(n1348), .ZN(n1383) );
INV_X1 U1103 ( .A(G101), .ZN(n1348) );
NAND2_X1 U1104 ( .A1(n1385), .A2(n1386), .ZN(n1382) );
INV_X1 U1105 ( .A(KEYINPUT15), .ZN(n1386) );
NAND2_X1 U1106 ( .A1(n1387), .A2(n1388), .ZN(n1385) );
XNOR2_X1 U1107 ( .A(KEYINPUT41), .B(G101), .ZN(n1387) );
NAND2_X1 U1108 ( .A1(KEYINPUT15), .A2(n1389), .ZN(n1381) );
NAND2_X1 U1109 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
OR2_X1 U1110 ( .A1(G101), .A2(KEYINPUT41), .ZN(n1391) );
NAND3_X1 U1111 ( .A1(G101), .A2(n1388), .A3(KEYINPUT41), .ZN(n1390) );
INV_X1 U1112 ( .A(n1384), .ZN(n1388) );
NAND2_X1 U1113 ( .A1(n1392), .A2(n1393), .ZN(n1384) );
NAND2_X1 U1114 ( .A1(KEYINPUT55), .A2(n1322), .ZN(n1393) );
XNOR2_X1 U1115 ( .A(G104), .B(G107), .ZN(n1322) );
OR3_X1 U1116 ( .A1(n1394), .A2(G107), .A3(KEYINPUT55), .ZN(n1392) );
INV_X1 U1117 ( .A(G104), .ZN(n1394) );
XNOR2_X1 U1118 ( .A(KEYINPUT39), .B(n1362), .ZN(n1365) );
NAND2_X1 U1119 ( .A1(n1395), .A2(n1396), .ZN(n1362) );
NAND2_X1 U1120 ( .A1(n1397), .A2(n1201), .ZN(n1396) );
INV_X1 U1121 ( .A(n1398), .ZN(n1201) );
NAND2_X1 U1122 ( .A1(n1399), .A2(n1398), .ZN(n1395) );
XOR2_X1 U1123 ( .A(G110), .B(KEYINPUT10), .Z(n1398) );
XOR2_X1 U1124 ( .A(KEYINPUT50), .B(n1397), .Z(n1399) );
XNOR2_X1 U1125 ( .A(n1196), .B(n1199), .ZN(n1397) );
XOR2_X1 U1126 ( .A(G140), .B(KEYINPUT34), .Z(n1199) );
NAND2_X1 U1127 ( .A1(G227), .A2(n1101), .ZN(n1196) );
INV_X1 U1128 ( .A(G953), .ZN(n1101) );
endmodule


