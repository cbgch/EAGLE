//Key = 1110000101110001110011101111010111110110010011111010101111101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362;

XOR2_X1 U749 ( .A(n1041), .B(n1042), .Z(G9) );
NAND2_X1 U750 ( .A1(KEYINPUT31), .A2(n1043), .ZN(n1041) );
INV_X1 U751 ( .A(G107), .ZN(n1043) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NOR2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NOR3_X1 U757 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NOR2_X1 U758 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U759 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U761 ( .A1(n1065), .A2(n1066), .ZN(n1057) );
NOR2_X1 U762 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
AND2_X1 U764 ( .A1(n1071), .A2(KEYINPUT2), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1054) );
NOR3_X1 U766 ( .A1(n1066), .A2(KEYINPUT2), .A3(n1074), .ZN(n1073) );
NOR3_X1 U767 ( .A1(n1060), .A2(n1075), .A3(n1066), .ZN(n1051) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1053), .ZN(n1077) );
NOR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NOR2_X1 U771 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NOR2_X1 U772 ( .A1(n1083), .A2(n1056), .ZN(n1076) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
INV_X1 U774 ( .A(n1086), .ZN(n1049) );
NAND3_X1 U775 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1046) );
NAND3_X1 U776 ( .A1(n1090), .A2(n1064), .A3(n1072), .ZN(n1089) );
INV_X1 U777 ( .A(KEYINPUT20), .ZN(n1064) );
NAND4_X1 U778 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1086), .ZN(n1090) );
NOR3_X1 U779 ( .A1(n1094), .A2(G953), .A3(G952), .ZN(n1044) );
INV_X1 U780 ( .A(n1087), .ZN(n1094) );
NAND4_X1 U781 ( .A1(n1095), .A2(n1093), .A3(n1096), .A4(n1097), .ZN(n1087) );
NOR4_X1 U782 ( .A1(n1098), .A2(n1099), .A3(n1056), .A4(n1100), .ZN(n1097) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
AND3_X1 U784 ( .A1(KEYINPUT54), .A2(n1103), .A3(G478), .ZN(n1102) );
NOR2_X1 U785 ( .A1(KEYINPUT54), .A2(G478), .ZN(n1101) );
XNOR2_X1 U786 ( .A(n1104), .B(n1105), .ZN(n1095) );
XOR2_X1 U787 ( .A(n1106), .B(KEYINPUT13), .Z(n1104) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(G72) );
XOR2_X1 U789 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U790 ( .A1(G953), .A2(n1111), .ZN(n1110) );
XOR2_X1 U791 ( .A(n1112), .B(KEYINPUT37), .Z(n1111) );
NOR2_X1 U792 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
AND2_X1 U793 ( .A1(G227), .A2(G900), .ZN(n1113) );
NOR2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1107) );
XOR2_X1 U795 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U796 ( .A(G125), .B(G140), .ZN(n1118) );
NAND2_X1 U797 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NAND2_X1 U798 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U799 ( .A(n1123), .B(KEYINPUT23), .Z(n1119) );
OR2_X1 U800 ( .A1(n1122), .A2(n1121), .ZN(n1123) );
AND2_X1 U801 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
NAND2_X1 U802 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U803 ( .A(KEYINPUT58), .B(n1128), .Z(n1126) );
NAND2_X1 U804 ( .A1(n1129), .A2(G131), .ZN(n1124) );
XOR2_X1 U805 ( .A(KEYINPUT39), .B(n1128), .Z(n1129) );
XNOR2_X1 U806 ( .A(n1130), .B(G137), .ZN(n1128) );
NAND2_X1 U807 ( .A1(KEYINPUT45), .A2(n1131), .ZN(n1130) );
XOR2_X1 U808 ( .A(n1132), .B(n1133), .Z(G69) );
XOR2_X1 U809 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U810 ( .A1(G953), .A2(n1136), .ZN(n1135) );
XNOR2_X1 U811 ( .A(KEYINPUT49), .B(n1137), .ZN(n1136) );
NAND2_X1 U812 ( .A1(n1138), .A2(n1139), .ZN(n1134) );
NAND2_X1 U813 ( .A1(G898), .A2(G224), .ZN(n1139) );
INV_X1 U814 ( .A(n1114), .ZN(n1138) );
XOR2_X1 U815 ( .A(n1088), .B(KEYINPUT53), .Z(n1114) );
NAND2_X1 U816 ( .A1(n1140), .A2(n1141), .ZN(n1132) );
NAND2_X1 U817 ( .A1(G953), .A2(n1142), .ZN(n1141) );
XNOR2_X1 U818 ( .A(n1143), .B(n1144), .ZN(n1140) );
XNOR2_X1 U819 ( .A(n1145), .B(n1146), .ZN(n1143) );
NOR2_X1 U820 ( .A1(KEYINPUT36), .A2(n1147), .ZN(n1146) );
NOR2_X1 U821 ( .A1(n1148), .A2(KEYINPUT28), .ZN(n1145) );
NOR2_X1 U822 ( .A1(n1149), .A2(n1150), .ZN(G66) );
NOR3_X1 U823 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR4_X1 U824 ( .A1(n1154), .A2(n1155), .A3(n1105), .A4(n1156), .ZN(n1153) );
NOR2_X1 U825 ( .A1(n1157), .A2(n1158), .ZN(n1152) );
NOR3_X1 U826 ( .A1(n1155), .A2(n1159), .A3(n1105), .ZN(n1157) );
INV_X1 U827 ( .A(KEYINPUT11), .ZN(n1155) );
NOR2_X1 U828 ( .A1(n1149), .A2(n1160), .ZN(G63) );
XOR2_X1 U829 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND2_X1 U830 ( .A1(n1163), .A2(G478), .ZN(n1161) );
NOR2_X1 U831 ( .A1(n1149), .A2(n1164), .ZN(G60) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U833 ( .A1(n1163), .A2(G475), .ZN(n1165) );
XNOR2_X1 U834 ( .A(G104), .B(n1167), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1168), .A2(KEYINPUT19), .ZN(n1167) );
NOR2_X1 U836 ( .A1(n1149), .A2(n1169), .ZN(G57) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U838 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U839 ( .A(n1174), .B(KEYINPUT29), .Z(n1173) );
NAND2_X1 U840 ( .A1(n1175), .A2(G101), .ZN(n1174) );
NOR2_X1 U841 ( .A1(n1175), .A2(n1176), .ZN(n1172) );
XNOR2_X1 U842 ( .A(G101), .B(KEYINPUT33), .ZN(n1176) );
NOR2_X1 U843 ( .A1(KEYINPUT3), .A2(n1177), .ZN(n1170) );
XOR2_X1 U844 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U846 ( .A(n1182), .B(KEYINPUT32), .Z(n1178) );
NAND2_X1 U847 ( .A1(n1163), .A2(G472), .ZN(n1182) );
NOR2_X1 U848 ( .A1(n1149), .A2(n1183), .ZN(G54) );
XOR2_X1 U849 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U850 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1184) );
NOR2_X1 U852 ( .A1(KEYINPUT61), .A2(n1144), .ZN(n1189) );
XOR2_X1 U853 ( .A(n1190), .B(KEYINPUT21), .Z(n1188) );
NAND2_X1 U854 ( .A1(n1191), .A2(n1163), .ZN(n1190) );
XNOR2_X1 U855 ( .A(G469), .B(KEYINPUT52), .ZN(n1191) );
NOR2_X1 U856 ( .A1(n1149), .A2(n1192), .ZN(G51) );
XOR2_X1 U857 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U858 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U859 ( .A(n1197), .B(n1198), .Z(n1193) );
NAND2_X1 U860 ( .A1(n1163), .A2(n1199), .ZN(n1197) );
INV_X1 U861 ( .A(n1156), .ZN(n1163) );
NAND2_X1 U862 ( .A1(G902), .A2(n1048), .ZN(n1156) );
INV_X1 U863 ( .A(n1159), .ZN(n1048) );
NOR2_X1 U864 ( .A1(n1137), .A2(n1112), .ZN(n1159) );
NAND4_X1 U865 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1112) );
NOR4_X1 U866 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
NOR2_X1 U867 ( .A1(n1063), .A2(n1208), .ZN(n1206) );
INV_X1 U868 ( .A(n1091), .ZN(n1063) );
NOR3_X1 U869 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1202) );
NOR2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
INV_X1 U871 ( .A(KEYINPUT60), .ZN(n1212) );
NOR2_X1 U872 ( .A1(KEYINPUT60), .A2(n1214), .ZN(n1210) );
NAND4_X1 U873 ( .A1(n1215), .A2(n1099), .A3(n1216), .A4(n1217), .ZN(n1214) );
AND2_X1 U874 ( .A1(n1085), .A2(n1218), .ZN(n1209) );
NAND2_X1 U875 ( .A1(n1219), .A2(n1220), .ZN(n1200) );
INV_X1 U876 ( .A(n1208), .ZN(n1220) );
XOR2_X1 U877 ( .A(n1221), .B(KEYINPUT56), .Z(n1219) );
NAND4_X1 U878 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1137) );
NOR4_X1 U879 ( .A1(n1226), .A2(n1168), .A3(n1227), .A4(n1042), .ZN(n1225) );
AND3_X1 U880 ( .A1(n1084), .A2(n1228), .A3(n1229), .ZN(n1042) );
NOR4_X1 U881 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1053), .ZN(n1227) );
AND3_X1 U882 ( .A1(n1229), .A2(n1228), .A3(n1085), .ZN(n1168) );
AND2_X1 U883 ( .A1(n1233), .A2(n1234), .ZN(n1224) );
NOR2_X1 U884 ( .A1(n1088), .A2(G952), .ZN(n1149) );
XOR2_X1 U885 ( .A(G146), .B(n1235), .Z(G48) );
NOR4_X1 U886 ( .A1(n1236), .A2(n1217), .A3(n1237), .A4(n1238), .ZN(n1235) );
XOR2_X1 U887 ( .A(n1074), .B(KEYINPUT8), .Z(n1236) );
XNOR2_X1 U888 ( .A(G143), .B(n1213), .ZN(G45) );
NAND4_X1 U889 ( .A1(n1215), .A2(n1080), .A3(n1099), .A4(n1216), .ZN(n1213) );
INV_X1 U890 ( .A(n1217), .ZN(n1080) );
XNOR2_X1 U891 ( .A(G140), .B(n1239), .ZN(G42) );
NAND3_X1 U892 ( .A1(n1240), .A2(n1091), .A3(n1241), .ZN(n1239) );
XOR2_X1 U893 ( .A(n1074), .B(KEYINPUT27), .Z(n1241) );
XOR2_X1 U894 ( .A(G137), .B(n1205), .Z(G39) );
NOR4_X1 U895 ( .A1(n1238), .A2(n1053), .A3(n1056), .A4(n1074), .ZN(n1205) );
INV_X1 U896 ( .A(n1092), .ZN(n1053) );
XOR2_X1 U897 ( .A(n1242), .B(n1243), .Z(G36) );
XOR2_X1 U898 ( .A(KEYINPUT44), .B(G134), .Z(n1243) );
NAND2_X1 U899 ( .A1(KEYINPUT35), .A2(n1244), .ZN(n1242) );
INV_X1 U900 ( .A(n1201), .ZN(n1244) );
NAND3_X1 U901 ( .A1(n1072), .A2(n1084), .A3(n1215), .ZN(n1201) );
NOR3_X1 U902 ( .A1(n1074), .A2(n1245), .A3(n1221), .ZN(n1215) );
XOR2_X1 U903 ( .A(n1246), .B(n1247), .Z(G33) );
NOR2_X1 U904 ( .A1(KEYINPUT40), .A2(n1127), .ZN(n1247) );
INV_X1 U905 ( .A(G131), .ZN(n1127) );
NOR2_X1 U906 ( .A1(n1221), .A2(n1208), .ZN(n1246) );
NAND2_X1 U907 ( .A1(n1240), .A2(n1071), .ZN(n1208) );
INV_X1 U908 ( .A(n1074), .ZN(n1071) );
NOR3_X1 U909 ( .A1(n1056), .A2(n1245), .A3(n1237), .ZN(n1240) );
INV_X1 U910 ( .A(n1072), .ZN(n1056) );
NOR2_X1 U911 ( .A1(n1081), .A2(n1248), .ZN(n1072) );
INV_X1 U912 ( .A(n1082), .ZN(n1248) );
NAND2_X1 U913 ( .A1(n1249), .A2(n1250), .ZN(G30) );
NAND2_X1 U914 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U915 ( .A(G128), .ZN(n1252) );
NAND2_X1 U916 ( .A1(G128), .A2(n1253), .ZN(n1249) );
NAND2_X1 U917 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U918 ( .A1(n1207), .A2(n1256), .ZN(n1255) );
INV_X1 U919 ( .A(n1257), .ZN(n1207) );
OR2_X1 U920 ( .A1(n1256), .A2(n1251), .ZN(n1254) );
NOR2_X1 U921 ( .A1(KEYINPUT43), .A2(n1257), .ZN(n1251) );
NAND2_X1 U922 ( .A1(n1218), .A2(n1084), .ZN(n1257) );
NOR3_X1 U923 ( .A1(n1217), .A2(n1074), .A3(n1238), .ZN(n1218) );
OR3_X1 U924 ( .A1(n1230), .A2(n1245), .A3(n1231), .ZN(n1238) );
INV_X1 U925 ( .A(KEYINPUT9), .ZN(n1256) );
XNOR2_X1 U926 ( .A(G101), .B(n1233), .ZN(G3) );
NAND3_X1 U927 ( .A1(n1062), .A2(n1229), .A3(n1092), .ZN(n1233) );
XNOR2_X1 U928 ( .A(n1204), .B(n1258), .ZN(G27) );
XOR2_X1 U929 ( .A(KEYINPUT7), .B(G125), .Z(n1258) );
AND4_X1 U930 ( .A1(n1091), .A2(n1085), .A3(n1259), .A4(n1093), .ZN(n1204) );
NOR2_X1 U931 ( .A1(n1245), .A2(n1217), .ZN(n1259) );
AND2_X1 U932 ( .A1(n1260), .A2(n1261), .ZN(n1245) );
NAND3_X1 U933 ( .A1(G902), .A2(n1086), .A3(n1115), .ZN(n1261) );
NOR2_X1 U934 ( .A1(n1088), .A2(G900), .ZN(n1115) );
XOR2_X1 U935 ( .A(n1262), .B(n1222), .Z(G24) );
NAND4_X1 U936 ( .A1(n1263), .A2(n1228), .A3(n1099), .A4(n1216), .ZN(n1222) );
INV_X1 U937 ( .A(n1066), .ZN(n1228) );
NAND2_X1 U938 ( .A1(n1264), .A2(n1230), .ZN(n1066) );
XOR2_X1 U939 ( .A(n1265), .B(n1266), .Z(G21) );
NAND4_X1 U940 ( .A1(n1092), .A2(n1093), .A3(n1267), .A4(n1268), .ZN(n1266) );
NOR3_X1 U941 ( .A1(n1231), .A2(n1269), .A3(n1230), .ZN(n1268) );
XOR2_X1 U942 ( .A(n1217), .B(KEYINPUT63), .Z(n1267) );
XOR2_X1 U943 ( .A(n1270), .B(G116), .Z(G18) );
NAND2_X1 U944 ( .A1(KEYINPUT22), .A2(n1234), .ZN(n1270) );
NAND3_X1 U945 ( .A1(n1062), .A2(n1084), .A3(n1263), .ZN(n1234) );
AND2_X1 U946 ( .A1(n1271), .A2(n1216), .ZN(n1084) );
XOR2_X1 U947 ( .A(KEYINPUT1), .B(n1099), .Z(n1271) );
INV_X1 U948 ( .A(n1221), .ZN(n1062) );
XNOR2_X1 U949 ( .A(n1226), .B(n1272), .ZN(G15) );
XOR2_X1 U950 ( .A(n1273), .B(KEYINPUT14), .Z(n1272) );
NOR3_X1 U951 ( .A1(n1232), .A2(n1221), .A3(n1237), .ZN(n1226) );
INV_X1 U952 ( .A(n1085), .ZN(n1237) );
NOR2_X1 U953 ( .A1(n1216), .A2(n1274), .ZN(n1085) );
NAND2_X1 U954 ( .A1(n1264), .A2(n1100), .ZN(n1221) );
XNOR2_X1 U955 ( .A(n1231), .B(KEYINPUT46), .ZN(n1264) );
INV_X1 U956 ( .A(n1263), .ZN(n1232) );
NOR3_X1 U957 ( .A1(n1217), .A2(n1269), .A3(n1060), .ZN(n1263) );
INV_X1 U958 ( .A(n1093), .ZN(n1060) );
NOR2_X1 U959 ( .A1(n1069), .A2(n1275), .ZN(n1093) );
INV_X1 U960 ( .A(n1070), .ZN(n1275) );
XOR2_X1 U961 ( .A(n1276), .B(n1223), .Z(G12) );
NAND3_X1 U962 ( .A1(n1092), .A2(n1229), .A3(n1091), .ZN(n1223) );
NOR2_X1 U963 ( .A1(n1100), .A2(n1231), .ZN(n1091) );
XNOR2_X1 U964 ( .A(n1277), .B(n1151), .ZN(n1231) );
INV_X1 U965 ( .A(n1106), .ZN(n1151) );
NAND2_X1 U966 ( .A1(n1154), .A2(n1278), .ZN(n1106) );
INV_X1 U967 ( .A(n1158), .ZN(n1154) );
XOR2_X1 U968 ( .A(n1279), .B(n1280), .Z(n1158) );
XOR2_X1 U969 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U970 ( .A(n1283), .B(n1284), .ZN(n1282) );
NOR2_X1 U971 ( .A1(G119), .A2(KEYINPUT4), .ZN(n1284) );
NAND2_X1 U972 ( .A1(KEYINPUT50), .A2(G137), .ZN(n1283) );
XOR2_X1 U973 ( .A(n1285), .B(n1286), .Z(n1279) );
XOR2_X1 U974 ( .A(G128), .B(G125), .Z(n1286) );
XOR2_X1 U975 ( .A(n1287), .B(n1288), .Z(n1285) );
NOR2_X1 U976 ( .A1(KEYINPUT42), .A2(G146), .ZN(n1288) );
NAND2_X1 U977 ( .A1(n1289), .A2(G221), .ZN(n1287) );
NAND2_X1 U978 ( .A1(KEYINPUT10), .A2(n1105), .ZN(n1277) );
NAND2_X1 U979 ( .A1(G217), .A2(n1290), .ZN(n1105) );
INV_X1 U980 ( .A(n1230), .ZN(n1100) );
XOR2_X1 U981 ( .A(n1291), .B(G472), .Z(n1230) );
NAND2_X1 U982 ( .A1(n1292), .A2(n1278), .ZN(n1291) );
XOR2_X1 U983 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U984 ( .A(n1295), .B(n1181), .Z(n1294) );
XNOR2_X1 U985 ( .A(n1296), .B(n1297), .ZN(n1181) );
XOR2_X1 U986 ( .A(G116), .B(n1298), .Z(n1297) );
NOR2_X1 U987 ( .A1(KEYINPUT18), .A2(n1273), .ZN(n1298) );
INV_X1 U988 ( .A(G113), .ZN(n1273) );
NAND2_X1 U989 ( .A1(KEYINPUT0), .A2(G119), .ZN(n1296) );
NOR2_X1 U990 ( .A1(KEYINPUT51), .A2(n1299), .ZN(n1295) );
XNOR2_X1 U991 ( .A(n1175), .B(n1300), .ZN(n1299) );
XNOR2_X1 U992 ( .A(G101), .B(KEYINPUT34), .ZN(n1300) );
AND3_X1 U993 ( .A1(n1301), .A2(n1088), .A3(G210), .ZN(n1175) );
NAND2_X1 U994 ( .A1(n1302), .A2(n1303), .ZN(n1293) );
NAND2_X1 U995 ( .A1(KEYINPUT57), .A2(n1180), .ZN(n1303) );
XOR2_X1 U996 ( .A(n1198), .B(n1304), .Z(n1180) );
OR3_X1 U997 ( .A1(n1198), .A2(n1304), .A3(KEYINPUT57), .ZN(n1302) );
NOR3_X1 U998 ( .A1(n1074), .A2(n1269), .A3(n1217), .ZN(n1229) );
NAND2_X1 U999 ( .A1(n1081), .A2(n1082), .ZN(n1217) );
NAND2_X1 U1000 ( .A1(G214), .A2(n1305), .ZN(n1082) );
XNOR2_X1 U1001 ( .A(n1306), .B(n1199), .ZN(n1081) );
AND2_X1 U1002 ( .A1(G210), .A2(n1305), .ZN(n1199) );
NAND2_X1 U1003 ( .A1(n1301), .A2(n1278), .ZN(n1305) );
NAND2_X1 U1004 ( .A1(n1307), .A2(n1278), .ZN(n1306) );
XOR2_X1 U1005 ( .A(n1308), .B(n1195), .Z(n1307) );
XNOR2_X1 U1006 ( .A(n1309), .B(n1147), .ZN(n1195) );
XOR2_X1 U1007 ( .A(n1310), .B(n1311), .Z(n1147) );
XOR2_X1 U1008 ( .A(G116), .B(G113), .Z(n1311) );
NAND2_X1 U1009 ( .A1(KEYINPUT26), .A2(n1265), .ZN(n1310) );
INV_X1 U1010 ( .A(G119), .ZN(n1265) );
XOR2_X1 U1011 ( .A(n1148), .B(n1144), .Z(n1309) );
AND3_X1 U1012 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1148) );
NAND2_X1 U1013 ( .A1(G122), .A2(n1315), .ZN(n1314) );
NAND2_X1 U1014 ( .A1(KEYINPUT48), .A2(n1276), .ZN(n1315) );
NAND4_X1 U1015 ( .A1(KEYINPUT48), .A2(n1262), .A3(KEYINPUT55), .A4(n1276), .ZN(n1313) );
INV_X1 U1016 ( .A(G122), .ZN(n1262) );
OR2_X1 U1017 ( .A1(n1276), .A2(KEYINPUT55), .ZN(n1312) );
NAND2_X1 U1018 ( .A1(n1316), .A2(KEYINPUT16), .ZN(n1308) );
XOR2_X1 U1019 ( .A(KEYINPUT30), .B(n1317), .Z(n1316) );
NOR2_X1 U1020 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NOR2_X1 U1021 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
XOR2_X1 U1022 ( .A(KEYINPUT62), .B(n1322), .Z(n1321) );
INV_X1 U1023 ( .A(n1198), .ZN(n1320) );
NOR2_X1 U1024 ( .A1(n1198), .A2(n1322), .ZN(n1318) );
INV_X1 U1025 ( .A(n1196), .ZN(n1322) );
XNOR2_X1 U1026 ( .A(G125), .B(n1323), .ZN(n1196) );
AND2_X1 U1027 ( .A1(n1088), .A2(G224), .ZN(n1323) );
XOR2_X1 U1028 ( .A(n1324), .B(n1325), .Z(n1198) );
XOR2_X1 U1029 ( .A(G146), .B(G128), .Z(n1325) );
NAND2_X1 U1030 ( .A1(KEYINPUT38), .A2(G143), .ZN(n1324) );
AND2_X1 U1031 ( .A1(n1326), .A2(n1260), .ZN(n1269) );
NAND3_X1 U1032 ( .A1(G952), .A2(n1086), .A3(n1327), .ZN(n1260) );
XOR2_X1 U1033 ( .A(n1088), .B(KEYINPUT12), .Z(n1327) );
NAND4_X1 U1034 ( .A1(G902), .A2(G953), .A3(n1086), .A4(n1142), .ZN(n1326) );
INV_X1 U1035 ( .A(G898), .ZN(n1142) );
NAND2_X1 U1036 ( .A1(G237), .A2(G234), .ZN(n1086) );
NAND2_X1 U1037 ( .A1(n1069), .A2(n1070), .ZN(n1074) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1290), .ZN(n1070) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1278), .ZN(n1290) );
XNOR2_X1 U1040 ( .A(n1328), .B(G469), .ZN(n1069) );
NAND2_X1 U1041 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XNOR2_X1 U1042 ( .A(n1187), .B(n1331), .ZN(n1330) );
XNOR2_X1 U1043 ( .A(n1332), .B(KEYINPUT17), .ZN(n1331) );
NAND2_X1 U1044 ( .A1(KEYINPUT15), .A2(n1333), .ZN(n1332) );
XOR2_X1 U1045 ( .A(n1186), .B(n1144), .Z(n1333) );
XNOR2_X1 U1046 ( .A(G101), .B(n1334), .ZN(n1144) );
XOR2_X1 U1047 ( .A(G107), .B(G104), .Z(n1334) );
XNOR2_X1 U1048 ( .A(n1122), .B(n1304), .ZN(n1186) );
XNOR2_X1 U1049 ( .A(n1335), .B(n1336), .ZN(n1304) );
NOR2_X1 U1050 ( .A1(KEYINPUT5), .A2(G131), .ZN(n1336) );
XOR2_X1 U1051 ( .A(n1131), .B(G137), .Z(n1335) );
INV_X1 U1052 ( .A(G134), .ZN(n1131) );
XNOR2_X1 U1053 ( .A(n1337), .B(n1338), .ZN(n1122) );
XOR2_X1 U1054 ( .A(KEYINPUT59), .B(G143), .Z(n1338) );
XOR2_X1 U1055 ( .A(n1339), .B(G128), .Z(n1337) );
NAND2_X1 U1056 ( .A1(KEYINPUT41), .A2(n1340), .ZN(n1339) );
INV_X1 U1057 ( .A(G146), .ZN(n1340) );
XNOR2_X1 U1058 ( .A(n1341), .B(n1281), .ZN(n1187) );
XOR2_X1 U1059 ( .A(G110), .B(G140), .Z(n1281) );
NAND2_X1 U1060 ( .A1(G227), .A2(n1088), .ZN(n1341) );
XOR2_X1 U1061 ( .A(n1278), .B(KEYINPUT6), .Z(n1329) );
NOR2_X1 U1062 ( .A1(n1216), .A2(n1099), .ZN(n1092) );
INV_X1 U1063 ( .A(n1274), .ZN(n1099) );
XOR2_X1 U1064 ( .A(n1342), .B(G475), .Z(n1274) );
NAND2_X1 U1065 ( .A1(n1166), .A2(n1278), .ZN(n1342) );
XOR2_X1 U1066 ( .A(n1343), .B(n1344), .Z(n1166) );
XOR2_X1 U1067 ( .A(G113), .B(n1345), .Z(n1344) );
XOR2_X1 U1068 ( .A(KEYINPUT25), .B(G122), .Z(n1345) );
XOR2_X1 U1069 ( .A(n1346), .B(G104), .Z(n1343) );
NAND2_X1 U1070 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NAND2_X1 U1071 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
XOR2_X1 U1072 ( .A(KEYINPUT24), .B(n1351), .Z(n1347) );
NOR2_X1 U1073 ( .A1(n1349), .A2(n1350), .ZN(n1351) );
XOR2_X1 U1074 ( .A(n1352), .B(n1353), .Z(n1350) );
XOR2_X1 U1075 ( .A(G143), .B(G131), .Z(n1353) );
NAND3_X1 U1076 ( .A1(n1301), .A2(n1088), .A3(G214), .ZN(n1352) );
INV_X1 U1077 ( .A(G237), .ZN(n1301) );
XOR2_X1 U1078 ( .A(n1354), .B(n1355), .Z(n1349) );
XOR2_X1 U1079 ( .A(G146), .B(G140), .Z(n1355) );
NAND2_X1 U1080 ( .A1(KEYINPUT47), .A2(G125), .ZN(n1354) );
OR2_X1 U1081 ( .A1(n1098), .A2(n1356), .ZN(n1216) );
AND2_X1 U1082 ( .A1(G478), .A2(n1103), .ZN(n1356) );
NOR2_X1 U1083 ( .A1(n1103), .A2(G478), .ZN(n1098) );
NAND2_X1 U1084 ( .A1(n1162), .A2(n1278), .ZN(n1103) );
INV_X1 U1085 ( .A(G902), .ZN(n1278) );
XNOR2_X1 U1086 ( .A(n1357), .B(n1358), .ZN(n1162) );
XOR2_X1 U1087 ( .A(n1359), .B(n1360), .Z(n1358) );
XOR2_X1 U1088 ( .A(G128), .B(G122), .Z(n1360) );
XOR2_X1 U1089 ( .A(G143), .B(G134), .Z(n1359) );
XOR2_X1 U1090 ( .A(n1361), .B(n1362), .Z(n1357) );
XOR2_X1 U1091 ( .A(G116), .B(G107), .Z(n1362) );
NAND2_X1 U1092 ( .A1(G217), .A2(n1289), .ZN(n1361) );
AND2_X1 U1093 ( .A1(G234), .A2(n1088), .ZN(n1289) );
INV_X1 U1094 ( .A(G953), .ZN(n1088) );
INV_X1 U1095 ( .A(G110), .ZN(n1276) );
endmodule


