//Key = 0111100001110100010001111011100100101100100110011101100001111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;

XNOR2_X1 U742 ( .A(G107), .B(n1026), .ZN(G9) );
NOR2_X1 U743 ( .A1(n1027), .A2(KEYINPUT46), .ZN(n1026) );
NOR2_X1 U744 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U745 ( .A1(G953), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
NOR2_X1 U746 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U748 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR3_X1 U749 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR3_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1041) );
NOR2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U755 ( .A1(n1044), .A2(n1053), .ZN(n1048) );
INV_X1 U756 ( .A(KEYINPUT27), .ZN(n1053) );
NOR2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1038) );
NOR3_X1 U758 ( .A1(n1044), .A2(n1056), .A3(n1047), .ZN(n1055) );
NOR2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR4_X1 U760 ( .A1(n1059), .A2(n1047), .A3(n1044), .A4(n1040), .ZN(n1035) );
NOR2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR3_X1 U762 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n1028) );
AND4_X1 U763 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1030) );
NOR4_X1 U764 ( .A1(n1066), .A2(n1067), .A3(n1044), .A4(n1068), .ZN(n1065) );
XOR2_X1 U765 ( .A(G472), .B(n1069), .Z(n1068) );
NOR2_X1 U766 ( .A1(KEYINPUT54), .A2(n1070), .ZN(n1069) );
XNOR2_X1 U767 ( .A(n1071), .B(n1072), .ZN(n1066) );
NAND2_X1 U768 ( .A1(KEYINPUT40), .A2(n1073), .ZN(n1071) );
INV_X1 U769 ( .A(G469), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1064) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1063) );
XNOR2_X1 U772 ( .A(n1078), .B(n1079), .ZN(n1062) );
NAND2_X1 U773 ( .A1(KEYINPUT37), .A2(n1080), .ZN(n1079) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(G72) );
NOR2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U776 ( .A(n1085), .B(KEYINPUT17), .Z(n1084) );
NAND3_X1 U777 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
NOR2_X1 U778 ( .A1(n1089), .A2(n1088), .ZN(n1083) );
NAND2_X1 U779 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NAND2_X1 U780 ( .A1(G953), .A2(n1092), .ZN(n1091) );
XOR2_X1 U781 ( .A(n1093), .B(n1094), .Z(n1090) );
XNOR2_X1 U782 ( .A(n1095), .B(n1096), .ZN(n1093) );
INV_X1 U783 ( .A(n1097), .ZN(n1096) );
NAND2_X1 U784 ( .A1(KEYINPUT36), .A2(n1098), .ZN(n1095) );
XOR2_X1 U785 ( .A(KEYINPUT2), .B(n1099), .Z(n1098) );
NOR2_X1 U786 ( .A1(G953), .A2(n1100), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(n1081) );
XOR2_X1 U788 ( .A(n1103), .B(KEYINPUT30), .Z(n1101) );
NAND2_X1 U789 ( .A1(G900), .A2(G227), .ZN(n1103) );
XOR2_X1 U790 ( .A(n1104), .B(n1105), .Z(G69) );
NOR2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U792 ( .A(KEYINPUT12), .B(n1108), .Z(n1107) );
NOR2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
AND3_X1 U794 ( .A1(n1109), .A2(n1087), .A3(n1110), .ZN(n1106) );
NAND2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U796 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1111) );
XNOR2_X1 U798 ( .A(n1116), .B(n1117), .ZN(n1115) );
NOR2_X1 U799 ( .A1(KEYINPUT8), .A2(n1118), .ZN(n1117) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1109) );
NAND2_X1 U802 ( .A1(n1102), .A2(n1123), .ZN(n1104) );
NAND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1123) );
XNOR2_X1 U804 ( .A(G953), .B(KEYINPUT9), .ZN(n1102) );
NOR2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U807 ( .A1(n1128), .A2(G217), .ZN(n1126) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1129), .ZN(G63) );
XOR2_X1 U809 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U810 ( .A1(n1128), .A2(G478), .ZN(n1130) );
NOR2_X1 U811 ( .A1(n1124), .A2(n1132), .ZN(G60) );
NOR3_X1 U812 ( .A1(n1078), .A2(n1133), .A3(n1134), .ZN(n1132) );
AND3_X1 U813 ( .A1(n1135), .A2(G475), .A3(n1128), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1135), .ZN(n1133) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1080), .ZN(n1136) );
NAND2_X1 U816 ( .A1(n1138), .A2(n1139), .ZN(G6) );
NAND2_X1 U817 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U818 ( .A1(n1142), .A2(G104), .ZN(n1138) );
NAND2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U820 ( .A1(KEYINPUT45), .A2(n1145), .ZN(n1144) );
INV_X1 U821 ( .A(n1122), .ZN(n1145) );
OR2_X1 U822 ( .A1(n1140), .A2(KEYINPUT45), .ZN(n1143) );
NOR2_X1 U823 ( .A1(KEYINPUT18), .A2(n1122), .ZN(n1140) );
NOR2_X1 U824 ( .A1(n1124), .A2(n1146), .ZN(G57) );
XOR2_X1 U825 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U826 ( .A(n1097), .B(n1149), .ZN(n1148) );
XOR2_X1 U827 ( .A(n1150), .B(n1151), .Z(n1147) );
XOR2_X1 U828 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U829 ( .A1(n1128), .A2(G472), .ZN(n1153) );
NAND3_X1 U830 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1152) );
NAND2_X1 U831 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
OR3_X1 U832 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1155) );
INV_X1 U833 ( .A(KEYINPUT47), .ZN(n1159) );
NAND2_X1 U834 ( .A1(KEYINPUT49), .A2(n1160), .ZN(n1157) );
OR2_X1 U835 ( .A1(n1160), .A2(KEYINPUT47), .ZN(n1154) );
XNOR2_X1 U836 ( .A(G101), .B(KEYINPUT56), .ZN(n1160) );
NOR3_X1 U837 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(G54) );
AND3_X1 U838 ( .A1(KEYINPUT29), .A2(G953), .A3(G952), .ZN(n1163) );
NOR2_X1 U839 ( .A1(KEYINPUT29), .A2(n1164), .ZN(n1162) );
INV_X1 U840 ( .A(n1124), .ZN(n1164) );
XOR2_X1 U841 ( .A(n1165), .B(n1166), .Z(n1161) );
NOR3_X1 U842 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
NOR3_X1 U843 ( .A1(n1170), .A2(n1097), .A3(n1171), .ZN(n1169) );
AND3_X1 U844 ( .A1(n1170), .A2(n1172), .A3(n1097), .ZN(n1168) );
NOR2_X1 U845 ( .A1(n1172), .A2(n1173), .ZN(n1167) );
XNOR2_X1 U846 ( .A(n1170), .B(n1097), .ZN(n1173) );
NAND3_X1 U847 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1170) );
NAND3_X1 U848 ( .A1(n1177), .A2(n1087), .A3(G227), .ZN(n1176) );
NAND2_X1 U849 ( .A1(KEYINPUT31), .A2(n1178), .ZN(n1177) );
OR2_X1 U850 ( .A1(n1179), .A2(KEYINPUT16), .ZN(n1178) );
OR2_X1 U851 ( .A1(n1179), .A2(KEYINPUT31), .ZN(n1175) );
NAND3_X1 U852 ( .A1(n1179), .A2(n1180), .A3(KEYINPUT31), .ZN(n1174) );
NAND3_X1 U853 ( .A1(n1087), .A2(n1181), .A3(G227), .ZN(n1180) );
INV_X1 U854 ( .A(KEYINPUT16), .ZN(n1181) );
XOR2_X1 U855 ( .A(G110), .B(n1182), .Z(n1179) );
NOR2_X1 U856 ( .A1(KEYINPUT0), .A2(n1183), .ZN(n1182) );
NAND2_X1 U857 ( .A1(KEYINPUT58), .A2(n1184), .ZN(n1165) );
NAND2_X1 U858 ( .A1(G469), .A2(n1128), .ZN(n1184) );
NOR2_X1 U859 ( .A1(n1124), .A2(n1185), .ZN(G51) );
XOR2_X1 U860 ( .A(n1186), .B(n1187), .Z(n1185) );
XNOR2_X1 U861 ( .A(n1188), .B(n1189), .ZN(n1187) );
XOR2_X1 U862 ( .A(n1190), .B(n1191), .Z(n1186) );
NOR2_X1 U863 ( .A1(KEYINPUT20), .A2(n1192), .ZN(n1191) );
NAND2_X1 U864 ( .A1(n1128), .A2(n1193), .ZN(n1190) );
NOR2_X1 U865 ( .A1(n1194), .A2(n1137), .ZN(n1128) );
INV_X1 U866 ( .A(n1032), .ZN(n1137) );
NAND3_X1 U867 ( .A1(n1100), .A2(n1195), .A3(n1121), .ZN(n1032) );
AND4_X1 U868 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1121) );
NOR4_X1 U869 ( .A1(n1200), .A2(n1201), .A3(n1027), .A4(n1202), .ZN(n1199) );
INV_X1 U870 ( .A(n1203), .ZN(n1202) );
AND3_X1 U871 ( .A1(n1060), .A2(n1204), .A3(n1205), .ZN(n1027) );
XNOR2_X1 U872 ( .A(KEYINPUT62), .B(n1122), .ZN(n1195) );
NAND3_X1 U873 ( .A1(n1205), .A2(n1204), .A3(n1061), .ZN(n1122) );
INV_X1 U874 ( .A(n1086), .ZN(n1100) );
NAND4_X1 U875 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1086) );
AND3_X1 U876 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1209) );
NAND2_X1 U877 ( .A1(n1213), .A2(n1214), .ZN(n1208) );
NAND2_X1 U878 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U879 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U880 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND2_X1 U881 ( .A1(n1045), .A2(n1060), .ZN(n1220) );
NAND2_X1 U882 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
XOR2_X1 U883 ( .A(n1223), .B(KEYINPUT63), .Z(n1215) );
NAND3_X1 U884 ( .A1(n1222), .A2(n1061), .A3(n1224), .ZN(n1206) );
NOR2_X1 U885 ( .A1(n1087), .A2(G952), .ZN(n1124) );
XOR2_X1 U886 ( .A(n1225), .B(n1226), .Z(G48) );
NOR2_X1 U887 ( .A1(KEYINPUT19), .A2(n1227), .ZN(n1226) );
AND3_X1 U888 ( .A1(n1224), .A2(n1228), .A3(n1061), .ZN(n1225) );
XNOR2_X1 U889 ( .A(n1229), .B(KEYINPUT6), .ZN(n1228) );
XNOR2_X1 U890 ( .A(G143), .B(n1207), .ZN(G45) );
NAND4_X1 U891 ( .A1(n1224), .A2(n1045), .A3(n1067), .A4(n1230), .ZN(n1207) );
NAND2_X1 U892 ( .A1(n1231), .A2(n1232), .ZN(G42) );
OR2_X1 U893 ( .A1(G140), .A2(KEYINPUT1), .ZN(n1232) );
XOR2_X1 U894 ( .A(n1233), .B(n1234), .Z(n1231) );
NOR2_X1 U895 ( .A1(n1044), .A2(n1223), .ZN(n1234) );
NAND3_X1 U896 ( .A1(n1061), .A2(n1046), .A3(n1217), .ZN(n1223) );
NAND2_X1 U897 ( .A1(KEYINPUT1), .A2(G140), .ZN(n1233) );
XOR2_X1 U898 ( .A(G137), .B(n1235), .Z(G39) );
NOR3_X1 U899 ( .A1(n1236), .A2(KEYINPUT14), .A3(n1044), .ZN(n1235) );
INV_X1 U900 ( .A(n1213), .ZN(n1044) );
XOR2_X1 U901 ( .A(KEYINPUT13), .B(n1237), .Z(n1236) );
NOR3_X1 U902 ( .A1(n1238), .A2(n1239), .A3(n1037), .ZN(n1237) );
INV_X1 U903 ( .A(n1221), .ZN(n1037) );
XNOR2_X1 U904 ( .A(n1222), .B(KEYINPUT15), .ZN(n1239) );
XNOR2_X1 U905 ( .A(G134), .B(n1240), .ZN(G36) );
NAND4_X1 U906 ( .A1(n1241), .A2(n1217), .A3(n1045), .A4(n1060), .ZN(n1240) );
XNOR2_X1 U907 ( .A(n1213), .B(KEYINPUT21), .ZN(n1241) );
XNOR2_X1 U908 ( .A(G131), .B(n1210), .ZN(G33) );
NAND4_X1 U909 ( .A1(n1217), .A2(n1061), .A3(n1045), .A4(n1213), .ZN(n1210) );
NOR2_X1 U910 ( .A1(n1052), .A2(n1242), .ZN(n1213) );
XNOR2_X1 U911 ( .A(G128), .B(n1212), .ZN(G30) );
NAND3_X1 U912 ( .A1(n1222), .A2(n1060), .A3(n1224), .ZN(n1212) );
NOR3_X1 U913 ( .A1(n1243), .A2(n1242), .A3(n1238), .ZN(n1224) );
INV_X1 U914 ( .A(n1217), .ZN(n1238) );
NOR3_X1 U915 ( .A1(n1244), .A2(n1075), .A3(n1057), .ZN(n1217) );
XNOR2_X1 U916 ( .A(G101), .B(n1198), .ZN(G3) );
NAND3_X1 U917 ( .A1(n1045), .A2(n1205), .A3(n1221), .ZN(n1198) );
XNOR2_X1 U918 ( .A(G125), .B(n1211), .ZN(G27) );
NAND4_X1 U919 ( .A1(n1054), .A2(n1046), .A3(n1061), .A4(n1245), .ZN(n1211) );
NOR3_X1 U920 ( .A1(n1243), .A2(n1242), .A3(n1244), .ZN(n1245) );
AND2_X1 U921 ( .A1(n1034), .A2(n1246), .ZN(n1244) );
NAND3_X1 U922 ( .A1(n1247), .A2(n1092), .A3(n1248), .ZN(n1246) );
INV_X1 U923 ( .A(G900), .ZN(n1092) );
INV_X1 U924 ( .A(n1051), .ZN(n1242) );
INV_X1 U925 ( .A(n1052), .ZN(n1243) );
NAND2_X1 U926 ( .A1(n1249), .A2(n1250), .ZN(G24) );
OR2_X1 U927 ( .A1(n1196), .A2(G122), .ZN(n1250) );
XOR2_X1 U928 ( .A(n1251), .B(KEYINPUT25), .Z(n1249) );
NAND2_X1 U929 ( .A1(G122), .A2(n1196), .ZN(n1251) );
NAND3_X1 U930 ( .A1(n1054), .A2(n1204), .A3(n1252), .ZN(n1196) );
NOR3_X1 U931 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1252) );
INV_X1 U932 ( .A(n1047), .ZN(n1204) );
NAND2_X1 U933 ( .A1(n1256), .A2(n1257), .ZN(n1047) );
XNOR2_X1 U934 ( .A(KEYINPUT44), .B(n1258), .ZN(n1257) );
XNOR2_X1 U935 ( .A(G119), .B(n1197), .ZN(G21) );
NAND4_X1 U936 ( .A1(n1221), .A2(n1222), .A3(n1054), .A4(n1259), .ZN(n1197) );
XOR2_X1 U937 ( .A(G116), .B(n1201), .Z(G18) );
AND2_X1 U938 ( .A1(n1260), .A2(n1060), .ZN(n1201) );
NOR2_X1 U939 ( .A1(n1230), .A2(n1255), .ZN(n1060) );
INV_X1 U940 ( .A(n1067), .ZN(n1255) );
XOR2_X1 U941 ( .A(G113), .B(n1200), .Z(G15) );
AND2_X1 U942 ( .A1(n1260), .A2(n1061), .ZN(n1200) );
NOR2_X1 U943 ( .A1(n1067), .A2(n1254), .ZN(n1061) );
AND3_X1 U944 ( .A1(n1054), .A2(n1259), .A3(n1045), .ZN(n1260) );
AND2_X1 U945 ( .A1(n1261), .A2(n1256), .ZN(n1045) );
XNOR2_X1 U946 ( .A(n1262), .B(KEYINPUT28), .ZN(n1261) );
INV_X1 U947 ( .A(n1253), .ZN(n1259) );
INV_X1 U948 ( .A(n1040), .ZN(n1054) );
NAND2_X1 U949 ( .A1(n1057), .A2(n1058), .ZN(n1040) );
XNOR2_X1 U950 ( .A(G110), .B(n1203), .ZN(G12) );
NAND3_X1 U951 ( .A1(n1205), .A2(n1046), .A3(n1221), .ZN(n1203) );
NOR2_X1 U952 ( .A1(n1067), .A2(n1230), .ZN(n1221) );
INV_X1 U953 ( .A(n1254), .ZN(n1230) );
XOR2_X1 U954 ( .A(n1078), .B(n1080), .Z(n1254) );
INV_X1 U955 ( .A(G475), .ZN(n1080) );
NOR2_X1 U956 ( .A1(n1135), .A2(G902), .ZN(n1078) );
XOR2_X1 U957 ( .A(n1263), .B(n1264), .Z(n1135) );
NOR2_X1 U958 ( .A1(KEYINPUT53), .A2(n1265), .ZN(n1264) );
XOR2_X1 U959 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U960 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U961 ( .A(n1270), .B(n1271), .ZN(n1269) );
NOR2_X1 U962 ( .A1(KEYINPUT7), .A2(n1272), .ZN(n1271) );
NAND2_X1 U963 ( .A1(KEYINPUT23), .A2(n1273), .ZN(n1270) );
INV_X1 U964 ( .A(G131), .ZN(n1273) );
NOR2_X1 U965 ( .A1(KEYINPUT50), .A2(n1274), .ZN(n1268) );
XOR2_X1 U966 ( .A(n1275), .B(n1276), .Z(n1266) );
AND3_X1 U967 ( .A1(G214), .A2(n1087), .A3(n1277), .ZN(n1276) );
XNOR2_X1 U968 ( .A(G146), .B(G140), .ZN(n1275) );
NAND3_X1 U969 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1263) );
NAND2_X1 U970 ( .A1(G104), .A2(n1281), .ZN(n1280) );
NAND3_X1 U971 ( .A1(n1282), .A2(n1141), .A3(KEYINPUT48), .ZN(n1279) );
INV_X1 U972 ( .A(n1281), .ZN(n1282) );
NAND2_X1 U973 ( .A1(KEYINPUT60), .A2(n1283), .ZN(n1281) );
OR2_X1 U974 ( .A1(n1283), .A2(KEYINPUT48), .ZN(n1278) );
XNOR2_X1 U975 ( .A(G113), .B(n1116), .ZN(n1283) );
INV_X1 U976 ( .A(G122), .ZN(n1116) );
XNOR2_X1 U977 ( .A(n1284), .B(G478), .ZN(n1067) );
NAND2_X1 U978 ( .A1(n1131), .A2(n1194), .ZN(n1284) );
XNOR2_X1 U979 ( .A(n1285), .B(n1286), .ZN(n1131) );
XOR2_X1 U980 ( .A(G134), .B(n1287), .Z(n1286) );
XNOR2_X1 U981 ( .A(KEYINPUT24), .B(n1274), .ZN(n1287) );
XNOR2_X1 U982 ( .A(n1288), .B(n1289), .ZN(n1285) );
INV_X1 U983 ( .A(n1290), .ZN(n1289) );
XOR2_X1 U984 ( .A(n1291), .B(n1292), .Z(n1288) );
AND3_X1 U985 ( .A1(G217), .A2(n1087), .A3(G234), .ZN(n1292) );
NAND2_X1 U986 ( .A1(KEYINPUT43), .A2(n1293), .ZN(n1291) );
NAND2_X1 U987 ( .A1(n1294), .A2(n1295), .ZN(n1046) );
OR2_X1 U988 ( .A1(n1229), .A2(KEYINPUT44), .ZN(n1295) );
INV_X1 U989 ( .A(n1222), .ZN(n1229) );
NOR2_X1 U990 ( .A1(n1258), .A2(n1256), .ZN(n1222) );
INV_X1 U991 ( .A(n1296), .ZN(n1256) );
NAND3_X1 U992 ( .A1(n1258), .A2(n1296), .A3(KEYINPUT44), .ZN(n1294) );
NAND3_X1 U993 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1296) );
INV_X1 U994 ( .A(n1074), .ZN(n1299) );
NOR2_X1 U995 ( .A1(n1077), .A2(n1076), .ZN(n1074) );
OR2_X1 U996 ( .A1(n1076), .A2(KEYINPUT11), .ZN(n1298) );
NAND3_X1 U997 ( .A1(n1076), .A2(n1077), .A3(KEYINPUT11), .ZN(n1297) );
NAND2_X1 U998 ( .A1(n1300), .A2(n1194), .ZN(n1077) );
XOR2_X1 U999 ( .A(KEYINPUT35), .B(n1127), .Z(n1300) );
XNOR2_X1 U1000 ( .A(n1301), .B(n1302), .ZN(n1127) );
AND3_X1 U1001 ( .A1(G221), .A2(n1087), .A3(G234), .ZN(n1302) );
XOR2_X1 U1002 ( .A(n1303), .B(G137), .Z(n1301) );
NAND2_X1 U1003 ( .A1(n1304), .A2(KEYINPUT3), .ZN(n1303) );
XOR2_X1 U1004 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1005 ( .A(n1293), .B(G119), .ZN(n1306) );
INV_X1 U1006 ( .A(G128), .ZN(n1293) );
XOR2_X1 U1007 ( .A(n1307), .B(n1308), .Z(n1305) );
NOR2_X1 U1008 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U1009 ( .A(n1311), .B(KEYINPUT52), .Z(n1310) );
NAND2_X1 U1010 ( .A1(n1312), .A2(n1227), .ZN(n1311) );
NOR2_X1 U1011 ( .A1(n1227), .A2(n1312), .ZN(n1309) );
XOR2_X1 U1012 ( .A(KEYINPUT59), .B(n1099), .Z(n1312) );
XNOR2_X1 U1013 ( .A(n1272), .B(G140), .ZN(n1099) );
INV_X1 U1014 ( .A(G125), .ZN(n1272) );
INV_X1 U1015 ( .A(G146), .ZN(n1227) );
NAND2_X1 U1016 ( .A1(KEYINPUT57), .A2(n1313), .ZN(n1307) );
INV_X1 U1017 ( .A(G110), .ZN(n1313) );
AND2_X1 U1018 ( .A1(n1314), .A2(n1315), .ZN(n1076) );
XNOR2_X1 U1019 ( .A(G217), .B(KEYINPUT22), .ZN(n1314) );
INV_X1 U1020 ( .A(n1262), .ZN(n1258) );
XNOR2_X1 U1021 ( .A(n1070), .B(G472), .ZN(n1262) );
NAND2_X1 U1022 ( .A1(n1316), .A2(n1194), .ZN(n1070) );
XOR2_X1 U1023 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U1024 ( .A(G101), .B(n1158), .ZN(n1318) );
NAND3_X1 U1025 ( .A1(n1277), .A2(n1087), .A3(G210), .ZN(n1158) );
NOR2_X1 U1026 ( .A1(n1319), .A2(n1320), .ZN(n1317) );
XOR2_X1 U1027 ( .A(KEYINPUT39), .B(n1321), .Z(n1320) );
NOR2_X1 U1028 ( .A1(n1149), .A2(n1322), .ZN(n1321) );
AND2_X1 U1029 ( .A1(n1322), .A2(n1149), .ZN(n1319) );
XOR2_X1 U1030 ( .A(G116), .B(n1323), .Z(n1149) );
NAND2_X1 U1031 ( .A1(n1324), .A2(n1325), .ZN(n1322) );
NAND2_X1 U1032 ( .A1(n1097), .A2(n1150), .ZN(n1325) );
XOR2_X1 U1033 ( .A(n1326), .B(KEYINPUT41), .Z(n1324) );
OR2_X1 U1034 ( .A1(n1097), .A2(n1150), .ZN(n1326) );
NOR3_X1 U1035 ( .A1(n1057), .A2(n1075), .A3(n1253), .ZN(n1205) );
NAND3_X1 U1036 ( .A1(n1327), .A2(n1051), .A3(n1052), .ZN(n1253) );
XNOR2_X1 U1037 ( .A(n1328), .B(n1193), .ZN(n1052) );
AND2_X1 U1038 ( .A1(G210), .A2(n1329), .ZN(n1193) );
NAND2_X1 U1039 ( .A1(n1330), .A2(n1194), .ZN(n1328) );
XOR2_X1 U1040 ( .A(n1188), .B(n1331), .Z(n1330) );
XNOR2_X1 U1041 ( .A(n1332), .B(n1192), .ZN(n1331) );
NAND2_X1 U1042 ( .A1(G224), .A2(n1087), .ZN(n1192) );
NAND2_X1 U1043 ( .A1(KEYINPUT34), .A2(n1189), .ZN(n1332) );
XOR2_X1 U1044 ( .A(n1333), .B(n1150), .Z(n1189) );
XOR2_X1 U1045 ( .A(G128), .B(n1334), .Z(n1150) );
NOR2_X1 U1046 ( .A1(KEYINPUT5), .A2(n1335), .ZN(n1334) );
XNOR2_X1 U1047 ( .A(G125), .B(KEYINPUT4), .ZN(n1333) );
XOR2_X1 U1048 ( .A(n1336), .B(n1120), .Z(n1188) );
XNOR2_X1 U1049 ( .A(n1323), .B(n1337), .ZN(n1120) );
XNOR2_X1 U1050 ( .A(G113), .B(G119), .ZN(n1323) );
XNOR2_X1 U1051 ( .A(n1290), .B(n1114), .ZN(n1336) );
AND2_X1 U1052 ( .A1(KEYINPUT51), .A2(G110), .ZN(n1114) );
XOR2_X1 U1053 ( .A(G122), .B(n1119), .Z(n1290) );
XOR2_X1 U1054 ( .A(G107), .B(G116), .Z(n1119) );
NAND2_X1 U1055 ( .A1(G214), .A2(n1329), .ZN(n1051) );
NAND2_X1 U1056 ( .A1(n1194), .A2(n1277), .ZN(n1329) );
INV_X1 U1057 ( .A(G237), .ZN(n1277) );
NAND2_X1 U1058 ( .A1(n1034), .A2(n1338), .ZN(n1327) );
NAND3_X1 U1059 ( .A1(n1248), .A2(n1113), .A3(n1339), .ZN(n1338) );
XOR2_X1 U1060 ( .A(n1247), .B(KEYINPUT32), .Z(n1339) );
INV_X1 U1061 ( .A(G898), .ZN(n1113) );
NOR2_X1 U1062 ( .A1(n1087), .A2(n1194), .ZN(n1248) );
NAND3_X1 U1063 ( .A1(n1247), .A2(n1087), .A3(G952), .ZN(n1034) );
INV_X1 U1064 ( .A(G953), .ZN(n1087) );
NAND2_X1 U1065 ( .A1(G237), .A2(G234), .ZN(n1247) );
INV_X1 U1066 ( .A(n1058), .ZN(n1075) );
NAND2_X1 U1067 ( .A1(G221), .A2(n1315), .ZN(n1058) );
NAND2_X1 U1068 ( .A1(G234), .A2(n1194), .ZN(n1315) );
XNOR2_X1 U1069 ( .A(n1072), .B(n1340), .ZN(n1057) );
NOR2_X1 U1070 ( .A1(G469), .A2(KEYINPUT55), .ZN(n1340) );
NAND2_X1 U1071 ( .A1(n1341), .A2(n1194), .ZN(n1072) );
INV_X1 U1072 ( .A(G902), .ZN(n1194) );
XOR2_X1 U1073 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1074 ( .A(n1344), .B(n1345), .ZN(n1343) );
NOR3_X1 U1075 ( .A1(KEYINPUT33), .A2(n1346), .A3(n1347), .ZN(n1345) );
NOR3_X1 U1076 ( .A1(n1172), .A2(KEYINPUT42), .A3(n1348), .ZN(n1347) );
INV_X1 U1077 ( .A(n1171), .ZN(n1172) );
NOR2_X1 U1078 ( .A1(n1349), .A2(n1171), .ZN(n1346) );
XNOR2_X1 U1079 ( .A(n1350), .B(n1351), .ZN(n1171) );
XOR2_X1 U1080 ( .A(KEYINPUT38), .B(G107), .Z(n1351) );
XNOR2_X1 U1081 ( .A(n1337), .B(n1094), .ZN(n1350) );
XOR2_X1 U1082 ( .A(n1352), .B(n1335), .Z(n1094) );
XOR2_X1 U1083 ( .A(n1274), .B(G146), .Z(n1335) );
INV_X1 U1084 ( .A(G143), .ZN(n1274) );
XNOR2_X1 U1085 ( .A(G128), .B(KEYINPUT61), .ZN(n1352) );
XNOR2_X1 U1086 ( .A(G101), .B(n1141), .ZN(n1337) );
INV_X1 U1087 ( .A(G104), .ZN(n1141) );
NOR2_X1 U1088 ( .A1(n1353), .A2(n1097), .ZN(n1349) );
NOR2_X1 U1089 ( .A1(n1348), .A2(n1354), .ZN(n1353) );
INV_X1 U1090 ( .A(KEYINPUT42), .ZN(n1354) );
XNOR2_X1 U1091 ( .A(n1097), .B(KEYINPUT26), .ZN(n1348) );
XOR2_X1 U1092 ( .A(G131), .B(n1355), .Z(n1097) );
XOR2_X1 U1093 ( .A(G137), .B(G134), .Z(n1355) );
NAND2_X1 U1094 ( .A1(KEYINPUT10), .A2(G227), .ZN(n1344) );
XNOR2_X1 U1095 ( .A(n1183), .B(G110), .ZN(n1342) );
INV_X1 U1096 ( .A(G140), .ZN(n1183) );
endmodule


