//Key = 1011111110001001000101001110011100000100111000001010001110111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;

XOR2_X1 U737 ( .A(G107), .B(n1018), .Z(G9) );
NOR2_X1 U738 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U739 ( .A1(G953), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1020) );
NOR2_X1 U740 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
INV_X1 U743 ( .A(n1030), .ZN(n1029) );
NOR2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
XOR2_X1 U750 ( .A(n1043), .B(KEYINPUT0), .Z(n1041) );
NOR2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(n1035) );
NOR2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1048), .A2(n1045), .ZN(n1031) );
NOR2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
AND2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U756 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1049) );
XOR2_X1 U757 ( .A(KEYINPUT62), .B(n1052), .Z(n1053) );
NOR4_X1 U758 ( .A1(n1056), .A2(n1045), .A3(n1038), .A4(n1034), .ZN(n1026) );
INV_X1 U759 ( .A(n1057), .ZN(n1045) );
NOR2_X1 U760 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR3_X1 U761 ( .A1(n1021), .A2(G953), .A3(G952), .ZN(n1019) );
AND4_X1 U762 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1021) );
NOR4_X1 U763 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
XNOR2_X1 U764 ( .A(n1068), .B(n1069), .ZN(n1067) );
NAND2_X1 U765 ( .A1(KEYINPUT19), .A2(n1070), .ZN(n1068) );
XNOR2_X1 U766 ( .A(KEYINPUT42), .B(n1071), .ZN(n1070) );
XOR2_X1 U767 ( .A(n1072), .B(KEYINPUT55), .Z(n1066) );
INV_X1 U768 ( .A(n1042), .ZN(n1065) );
NOR2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1062) );
XOR2_X1 U770 ( .A(KEYINPUT36), .B(n1055), .Z(n1074) );
INV_X1 U771 ( .A(n1075), .ZN(n1055) );
XOR2_X1 U772 ( .A(KEYINPUT2), .B(n1076), .Z(n1061) );
NAND2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(G72) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U776 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NAND2_X1 U777 ( .A1(G900), .A2(G227), .ZN(n1083) );
NAND2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND2_X1 U779 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NAND2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1077) );
NAND2_X1 U781 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND3_X1 U782 ( .A1(n1086), .A2(n1087), .A3(n1085), .ZN(n1091) );
NAND2_X1 U783 ( .A1(G227), .A2(G953), .ZN(n1090) );
INV_X1 U784 ( .A(n1080), .ZN(n1088) );
NAND3_X1 U785 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1080) );
XOR2_X1 U786 ( .A(KEYINPUT12), .B(n1095), .Z(n1094) );
NOR2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NAND2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U790 ( .A1(G140), .A2(n1100), .ZN(n1099) );
XOR2_X1 U791 ( .A(n1101), .B(KEYINPUT18), .Z(n1098) );
NAND2_X1 U792 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U793 ( .A(KEYINPUT1), .B(G125), .Z(n1102) );
XOR2_X1 U794 ( .A(n1104), .B(n1105), .Z(n1096) );
XOR2_X1 U795 ( .A(n1106), .B(n1107), .Z(n1105) );
XNOR2_X1 U796 ( .A(G131), .B(KEYINPUT25), .ZN(n1107) );
NAND2_X1 U797 ( .A1(KEYINPUT7), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U798 ( .A(n1109), .B(n1110), .ZN(n1104) );
NAND2_X1 U799 ( .A1(G953), .A2(n1111), .ZN(n1092) );
NAND2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(G69) );
NAND2_X1 U801 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND3_X1 U802 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1114) );
XNOR2_X1 U803 ( .A(KEYINPUT48), .B(n1119), .ZN(n1118) );
NAND2_X1 U804 ( .A1(G953), .A2(n1120), .ZN(n1116) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1112) );
NAND2_X1 U806 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
OR2_X1 U807 ( .A1(n1119), .A2(KEYINPUT48), .ZN(n1124) );
NAND2_X1 U808 ( .A1(KEYINPUT48), .A2(n1125), .ZN(n1123) );
NAND2_X1 U809 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U810 ( .A1(n1119), .A2(n1085), .ZN(n1127) );
NAND2_X1 U811 ( .A1(G953), .A2(G224), .ZN(n1126) );
INV_X1 U812 ( .A(n1115), .ZN(n1121) );
NAND2_X1 U813 ( .A1(n1128), .A2(n1117), .ZN(n1115) );
INV_X1 U814 ( .A(n1129), .ZN(n1117) );
XOR2_X1 U815 ( .A(n1130), .B(n1131), .Z(n1128) );
NOR2_X1 U816 ( .A1(KEYINPUT39), .A2(n1132), .ZN(n1131) );
NOR2_X1 U817 ( .A1(n1133), .A2(n1134), .ZN(G66) );
XOR2_X1 U818 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U819 ( .A(KEYINPUT32), .B(n1137), .Z(n1136) );
NOR2_X1 U820 ( .A1(n1069), .A2(n1138), .ZN(n1137) );
NOR2_X1 U821 ( .A1(n1133), .A2(n1139), .ZN(G63) );
XNOR2_X1 U822 ( .A(n1140), .B(n1141), .ZN(n1139) );
AND2_X1 U823 ( .A1(G478), .A2(n1142), .ZN(n1141) );
NOR2_X1 U824 ( .A1(n1133), .A2(n1143), .ZN(G60) );
NOR2_X1 U825 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U826 ( .A(KEYINPUT52), .B(n1146), .Z(n1145) );
NOR2_X1 U827 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XNOR2_X1 U828 ( .A(KEYINPUT9), .B(n1149), .ZN(n1148) );
NOR2_X1 U829 ( .A1(n1149), .A2(n1150), .ZN(n1144) );
XNOR2_X1 U830 ( .A(KEYINPUT33), .B(n1147), .ZN(n1150) );
NAND2_X1 U831 ( .A1(n1142), .A2(G475), .ZN(n1149) );
NAND2_X1 U832 ( .A1(n1151), .A2(n1152), .ZN(G6) );
NAND2_X1 U833 ( .A1(G104), .A2(n1153), .ZN(n1152) );
XOR2_X1 U834 ( .A(n1154), .B(KEYINPUT35), .Z(n1151) );
OR2_X1 U835 ( .A1(n1153), .A2(G104), .ZN(n1154) );
NAND4_X1 U836 ( .A1(n1059), .A2(n1052), .A3(n1155), .A4(n1156), .ZN(n1153) );
XOR2_X1 U837 ( .A(KEYINPUT47), .B(n1051), .Z(n1156) );
NOR2_X1 U838 ( .A1(n1133), .A2(n1157), .ZN(G57) );
XOR2_X1 U839 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U840 ( .A(n1160), .B(n1161), .Z(n1158) );
AND2_X1 U841 ( .A1(G472), .A2(n1142), .ZN(n1161) );
NAND2_X1 U842 ( .A1(n1162), .A2(n1163), .ZN(n1160) );
NAND2_X1 U843 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XOR2_X1 U844 ( .A(n1166), .B(KEYINPUT20), .Z(n1162) );
NAND2_X1 U845 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U846 ( .A(KEYINPUT16), .B(n1169), .Z(n1168) );
NOR2_X1 U847 ( .A1(n1133), .A2(n1170), .ZN(G54) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U849 ( .A(n1169), .B(n1173), .Z(n1172) );
XOR2_X1 U850 ( .A(n1174), .B(n1175), .Z(n1171) );
AND2_X1 U851 ( .A1(G469), .A2(n1142), .ZN(n1175) );
INV_X1 U852 ( .A(n1138), .ZN(n1142) );
NAND3_X1 U853 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1174) );
NAND2_X1 U854 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
OR3_X1 U855 ( .A1(n1179), .A2(n1180), .A3(KEYINPUT63), .ZN(n1177) );
OR2_X1 U856 ( .A1(KEYINPUT23), .A2(n1181), .ZN(n1179) );
NAND2_X1 U857 ( .A1(KEYINPUT63), .A2(n1181), .ZN(n1176) );
XOR2_X1 U858 ( .A(n1182), .B(G140), .Z(n1181) );
NOR2_X1 U859 ( .A1(n1133), .A2(n1183), .ZN(G51) );
XOR2_X1 U860 ( .A(n1184), .B(n1185), .Z(n1183) );
XOR2_X1 U861 ( .A(n1186), .B(n1187), .Z(n1184) );
NOR2_X1 U862 ( .A1(n1188), .A2(n1138), .ZN(n1187) );
NAND2_X1 U863 ( .A1(G902), .A2(n1023), .ZN(n1138) );
NAND3_X1 U864 ( .A1(n1119), .A2(n1086), .A3(n1189), .ZN(n1023) );
XOR2_X1 U865 ( .A(n1087), .B(KEYINPUT10), .Z(n1189) );
AND4_X1 U866 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1086) );
AND4_X1 U867 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NAND3_X1 U868 ( .A1(n1058), .A2(n1040), .A3(n1198), .ZN(n1192) );
AND4_X1 U869 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1119) );
NOR4_X1 U870 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
NOR2_X1 U871 ( .A1(n1207), .A2(n1018), .ZN(n1201) );
NOR3_X1 U872 ( .A1(n1208), .A2(n1038), .A3(n1209), .ZN(n1018) );
AND3_X1 U873 ( .A1(n1059), .A2(n1052), .A3(n1210), .ZN(n1207) );
INV_X1 U874 ( .A(n1038), .ZN(n1052) );
OR2_X1 U875 ( .A1(n1211), .A2(n1212), .ZN(n1199) );
NAND2_X1 U876 ( .A1(n1213), .A2(n1214), .ZN(n1186) );
NAND2_X1 U877 ( .A1(n1165), .A2(n1215), .ZN(n1214) );
NAND2_X1 U878 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U879 ( .A1(KEYINPUT24), .A2(n1100), .ZN(n1217) );
INV_X1 U880 ( .A(n1167), .ZN(n1165) );
NAND2_X1 U881 ( .A1(G125), .A2(n1218), .ZN(n1213) );
NAND2_X1 U882 ( .A1(KEYINPUT24), .A2(n1219), .ZN(n1218) );
NAND2_X1 U883 ( .A1(n1167), .A2(n1216), .ZN(n1219) );
INV_X1 U884 ( .A(KEYINPUT28), .ZN(n1216) );
NOR2_X1 U885 ( .A1(n1085), .A2(G952), .ZN(n1133) );
XNOR2_X1 U886 ( .A(G146), .B(n1190), .ZN(G48) );
NAND3_X1 U887 ( .A1(n1059), .A2(n1040), .A3(n1198), .ZN(n1190) );
XNOR2_X1 U888 ( .A(G143), .B(n1191), .ZN(G45) );
NAND4_X1 U889 ( .A1(n1220), .A2(n1047), .A3(n1221), .A4(n1222), .ZN(n1191) );
NOR2_X1 U890 ( .A1(n1223), .A2(n1212), .ZN(n1221) );
XOR2_X1 U891 ( .A(n1103), .B(n1197), .Z(G42) );
NAND4_X1 U892 ( .A1(n1220), .A2(n1059), .A3(n1046), .A4(n1057), .ZN(n1197) );
XNOR2_X1 U893 ( .A(G137), .B(n1087), .ZN(G39) );
NAND3_X1 U894 ( .A1(n1030), .A2(n1057), .A3(n1198), .ZN(n1087) );
INV_X1 U895 ( .A(n1224), .ZN(n1198) );
XNOR2_X1 U896 ( .A(G134), .B(n1196), .ZN(G36) );
NAND4_X1 U897 ( .A1(n1220), .A2(n1047), .A3(n1058), .A4(n1057), .ZN(n1196) );
XNOR2_X1 U898 ( .A(G131), .B(n1195), .ZN(G33) );
NAND4_X1 U899 ( .A1(n1220), .A2(n1059), .A3(n1047), .A4(n1057), .ZN(n1195) );
NAND2_X1 U900 ( .A1(n1225), .A2(n1226), .ZN(n1057) );
OR2_X1 U901 ( .A1(n1212), .A2(KEYINPUT0), .ZN(n1226) );
NAND3_X1 U902 ( .A1(n1043), .A2(n1042), .A3(KEYINPUT0), .ZN(n1225) );
XOR2_X1 U903 ( .A(n1227), .B(n1228), .Z(G30) );
NAND2_X1 U904 ( .A1(n1040), .A2(n1229), .ZN(n1228) );
XOR2_X1 U905 ( .A(KEYINPUT14), .B(n1230), .Z(n1229) );
NOR2_X1 U906 ( .A1(n1208), .A2(n1224), .ZN(n1230) );
NAND3_X1 U907 ( .A1(n1073), .A2(n1231), .A3(n1220), .ZN(n1224) );
AND2_X1 U908 ( .A1(n1051), .A2(n1232), .ZN(n1220) );
XOR2_X1 U909 ( .A(G101), .B(n1206), .Z(G3) );
AND3_X1 U910 ( .A1(n1030), .A2(n1210), .A3(n1047), .ZN(n1206) );
XNOR2_X1 U911 ( .A(n1233), .B(n1194), .ZN(G27) );
NAND4_X1 U912 ( .A1(n1059), .A2(n1234), .A3(n1235), .A4(n1046), .ZN(n1194) );
AND2_X1 U913 ( .A1(n1232), .A2(n1040), .ZN(n1235) );
NAND2_X1 U914 ( .A1(n1236), .A2(n1025), .ZN(n1232) );
XOR2_X1 U915 ( .A(n1237), .B(KEYINPUT11), .Z(n1236) );
NAND4_X1 U916 ( .A1(G902), .A2(G953), .A3(n1238), .A4(n1111), .ZN(n1237) );
INV_X1 U917 ( .A(G900), .ZN(n1111) );
NAND2_X1 U918 ( .A1(KEYINPUT30), .A2(n1100), .ZN(n1233) );
XOR2_X1 U919 ( .A(G122), .B(n1205), .Z(G24) );
AND4_X1 U920 ( .A1(n1155), .A2(n1239), .A3(n1222), .A4(n1240), .ZN(n1205) );
NOR2_X1 U921 ( .A1(n1038), .A2(n1034), .ZN(n1240) );
NAND2_X1 U922 ( .A1(n1241), .A2(n1242), .ZN(n1038) );
INV_X1 U923 ( .A(n1223), .ZN(n1239) );
XOR2_X1 U924 ( .A(G119), .B(n1204), .Z(G21) );
AND4_X1 U925 ( .A1(n1234), .A2(n1030), .A3(n1243), .A4(n1155), .ZN(n1204) );
NOR2_X1 U926 ( .A1(n1241), .A2(n1242), .ZN(n1243) );
XNOR2_X1 U927 ( .A(G116), .B(n1200), .ZN(G18) );
NAND4_X1 U928 ( .A1(n1047), .A2(n1234), .A3(n1058), .A4(n1155), .ZN(n1200) );
INV_X1 U929 ( .A(n1208), .ZN(n1058) );
NAND2_X1 U930 ( .A1(n1222), .A2(n1072), .ZN(n1208) );
XOR2_X1 U931 ( .A(n1244), .B(n1245), .Z(G15) );
NAND2_X1 U932 ( .A1(n1246), .A2(n1040), .ZN(n1245) );
XOR2_X1 U933 ( .A(n1211), .B(KEYINPUT4), .Z(n1246) );
NAND4_X1 U934 ( .A1(n1059), .A2(n1047), .A3(n1234), .A4(n1247), .ZN(n1211) );
INV_X1 U935 ( .A(n1034), .ZN(n1234) );
NAND2_X1 U936 ( .A1(n1075), .A2(n1248), .ZN(n1034) );
XOR2_X1 U937 ( .A(KEYINPUT41), .B(n1064), .Z(n1248) );
NOR2_X1 U938 ( .A1(n1231), .A2(n1242), .ZN(n1047) );
NOR2_X1 U939 ( .A1(n1223), .A2(n1222), .ZN(n1059) );
XOR2_X1 U940 ( .A(n1072), .B(KEYINPUT27), .Z(n1223) );
INV_X1 U941 ( .A(n1249), .ZN(n1072) );
XOR2_X1 U942 ( .A(n1182), .B(n1250), .Z(G12) );
NAND2_X1 U943 ( .A1(KEYINPUT59), .A2(n1203), .ZN(n1250) );
AND3_X1 U944 ( .A1(n1030), .A2(n1210), .A3(n1046), .ZN(n1203) );
NOR2_X1 U945 ( .A1(n1073), .A2(n1241), .ZN(n1046) );
INV_X1 U946 ( .A(n1231), .ZN(n1241) );
XOR2_X1 U947 ( .A(n1071), .B(n1069), .Z(n1231) );
NAND2_X1 U948 ( .A1(G217), .A2(n1251), .ZN(n1069) );
NAND2_X1 U949 ( .A1(n1252), .A2(n1253), .ZN(n1071) );
XOR2_X1 U950 ( .A(KEYINPUT34), .B(n1254), .Z(n1252) );
INV_X1 U951 ( .A(n1135), .ZN(n1254) );
XOR2_X1 U952 ( .A(n1255), .B(n1256), .Z(n1135) );
XNOR2_X1 U953 ( .A(n1257), .B(n1258), .ZN(n1256) );
XOR2_X1 U954 ( .A(n1259), .B(n1109), .Z(n1258) );
XOR2_X1 U955 ( .A(G137), .B(G128), .Z(n1109) );
NAND2_X1 U956 ( .A1(n1260), .A2(G221), .ZN(n1259) );
XOR2_X1 U957 ( .A(n1261), .B(n1262), .Z(n1255) );
XOR2_X1 U958 ( .A(KEYINPUT38), .B(G119), .Z(n1262) );
XOR2_X1 U959 ( .A(n1182), .B(n1263), .Z(n1261) );
NOR2_X1 U960 ( .A1(KEYINPUT51), .A2(n1264), .ZN(n1263) );
INV_X1 U961 ( .A(n1242), .ZN(n1073) );
XOR2_X1 U962 ( .A(n1265), .B(G472), .Z(n1242) );
NAND2_X1 U963 ( .A1(n1266), .A2(n1253), .ZN(n1265) );
XOR2_X1 U964 ( .A(n1167), .B(n1267), .Z(n1266) );
XOR2_X1 U965 ( .A(n1159), .B(n1169), .Z(n1267) );
INV_X1 U966 ( .A(n1164), .ZN(n1169) );
XNOR2_X1 U967 ( .A(n1268), .B(n1269), .ZN(n1159) );
XOR2_X1 U968 ( .A(KEYINPUT29), .B(n1270), .Z(n1269) );
AND2_X1 U969 ( .A1(G210), .A2(n1271), .ZN(n1270) );
INV_X1 U970 ( .A(n1209), .ZN(n1210) );
NAND2_X1 U971 ( .A1(n1155), .A2(n1051), .ZN(n1209) );
NOR2_X1 U972 ( .A1(n1075), .A2(n1064), .ZN(n1051) );
INV_X1 U973 ( .A(n1054), .ZN(n1064) );
NAND2_X1 U974 ( .A1(G221), .A2(n1251), .ZN(n1054) );
NAND2_X1 U975 ( .A1(G234), .A2(n1253), .ZN(n1251) );
XOR2_X1 U976 ( .A(n1272), .B(G469), .Z(n1075) );
NAND2_X1 U977 ( .A1(n1273), .A2(n1253), .ZN(n1272) );
XOR2_X1 U978 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U979 ( .A(n1276), .B(n1164), .Z(n1275) );
XOR2_X1 U980 ( .A(n1277), .B(n1278), .Z(n1164) );
NOR2_X1 U981 ( .A1(KEYINPUT61), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U982 ( .A(G137), .B(n1280), .ZN(n1279) );
NAND2_X1 U983 ( .A1(KEYINPUT26), .A2(n1108), .ZN(n1280) );
XNOR2_X1 U984 ( .A(G134), .B(KEYINPUT46), .ZN(n1108) );
XNOR2_X1 U985 ( .A(G131), .B(KEYINPUT49), .ZN(n1277) );
NAND2_X1 U986 ( .A1(KEYINPUT3), .A2(n1182), .ZN(n1276) );
XOR2_X1 U987 ( .A(n1281), .B(n1282), .Z(n1274) );
XOR2_X1 U988 ( .A(n1103), .B(n1180), .Z(n1282) );
NAND2_X1 U989 ( .A1(G227), .A2(n1085), .ZN(n1180) );
NAND2_X1 U990 ( .A1(KEYINPUT37), .A2(n1173), .ZN(n1281) );
XNOR2_X1 U991 ( .A(n1283), .B(n1284), .ZN(n1173) );
XOR2_X1 U992 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U993 ( .A(G107), .B(G101), .Z(n1286) );
XOR2_X1 U994 ( .A(n1287), .B(G128), .Z(n1283) );
XNOR2_X1 U995 ( .A(KEYINPUT22), .B(KEYINPUT17), .ZN(n1287) );
AND2_X1 U996 ( .A1(n1040), .A2(n1247), .ZN(n1155) );
NAND2_X1 U997 ( .A1(n1025), .A2(n1288), .ZN(n1247) );
NAND3_X1 U998 ( .A1(n1129), .A2(n1238), .A3(G902), .ZN(n1288) );
NOR2_X1 U999 ( .A1(G898), .A2(n1085), .ZN(n1129) );
NAND3_X1 U1000 ( .A1(n1238), .A2(n1085), .A3(G952), .ZN(n1025) );
NAND2_X1 U1001 ( .A1(G237), .A2(G234), .ZN(n1238) );
INV_X1 U1002 ( .A(n1212), .ZN(n1040) );
NAND2_X1 U1003 ( .A1(n1076), .A2(n1042), .ZN(n1212) );
NAND2_X1 U1004 ( .A1(G214), .A2(n1289), .ZN(n1042) );
INV_X1 U1005 ( .A(n1043), .ZN(n1076) );
XNOR2_X1 U1006 ( .A(n1290), .B(n1188), .ZN(n1043) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1289), .ZN(n1188) );
NAND2_X1 U1008 ( .A1(n1291), .A2(n1253), .ZN(n1289) );
INV_X1 U1009 ( .A(G237), .ZN(n1291) );
NAND3_X1 U1010 ( .A1(n1292), .A2(n1293), .A3(n1253), .ZN(n1290) );
NAND2_X1 U1011 ( .A1(n1294), .A2(n1100), .ZN(n1293) );
XOR2_X1 U1012 ( .A(n1295), .B(KEYINPUT6), .Z(n1294) );
NAND2_X1 U1013 ( .A1(n1296), .A2(G125), .ZN(n1292) );
XOR2_X1 U1014 ( .A(n1295), .B(KEYINPUT45), .Z(n1296) );
XOR2_X1 U1015 ( .A(n1185), .B(n1167), .Z(n1295) );
XOR2_X1 U1016 ( .A(n1297), .B(G128), .Z(n1167) );
NAND2_X1 U1017 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U1018 ( .A1(n1264), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1019 ( .A(KEYINPUT15), .B(n1301), .Z(n1298) );
NOR2_X1 U1020 ( .A1(n1264), .A2(n1300), .ZN(n1301) );
XOR2_X1 U1021 ( .A(n1302), .B(n1132), .Z(n1185) );
XOR2_X1 U1022 ( .A(n1268), .B(n1303), .Z(n1132) );
XOR2_X1 U1023 ( .A(KEYINPUT43), .B(n1304), .Z(n1303) );
NOR2_X1 U1024 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U1025 ( .A(n1307), .B(KEYINPUT31), .Z(n1306) );
NAND2_X1 U1026 ( .A1(G107), .A2(n1308), .ZN(n1307) );
NOR2_X1 U1027 ( .A1(G107), .A2(n1308), .ZN(n1305) );
XOR2_X1 U1028 ( .A(n1309), .B(n1310), .Z(n1268) );
XOR2_X1 U1029 ( .A(G113), .B(G101), .Z(n1310) );
XNOR2_X1 U1030 ( .A(G116), .B(n1311), .ZN(n1309) );
XOR2_X1 U1031 ( .A(KEYINPUT54), .B(G119), .Z(n1311) );
XOR2_X1 U1032 ( .A(n1130), .B(n1312), .Z(n1302) );
NOR2_X1 U1033 ( .A1(G953), .A2(n1120), .ZN(n1312) );
INV_X1 U1034 ( .A(G224), .ZN(n1120) );
XOR2_X1 U1035 ( .A(n1313), .B(KEYINPUT50), .Z(n1130) );
NAND2_X1 U1036 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND2_X1 U1037 ( .A1(G110), .A2(n1316), .ZN(n1315) );
XOR2_X1 U1038 ( .A(KEYINPUT58), .B(n1317), .Z(n1314) );
NOR2_X1 U1039 ( .A1(G110), .A2(n1316), .ZN(n1317) );
XOR2_X1 U1040 ( .A(KEYINPUT56), .B(G122), .Z(n1316) );
NOR2_X1 U1041 ( .A1(n1249), .A2(n1222), .ZN(n1030) );
XOR2_X1 U1042 ( .A(n1060), .B(KEYINPUT5), .Z(n1222) );
XOR2_X1 U1043 ( .A(n1318), .B(G478), .Z(n1060) );
NAND2_X1 U1044 ( .A1(n1140), .A2(n1253), .ZN(n1318) );
INV_X1 U1045 ( .A(G902), .ZN(n1253) );
XNOR2_X1 U1046 ( .A(n1319), .B(n1320), .ZN(n1140) );
XNOR2_X1 U1047 ( .A(n1300), .B(n1321), .ZN(n1320) );
XOR2_X1 U1048 ( .A(n1322), .B(n1323), .Z(n1321) );
NOR2_X1 U1049 ( .A1(KEYINPUT57), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1050 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1051 ( .A(G116), .B(G107), .Z(n1326) );
XOR2_X1 U1052 ( .A(n1327), .B(G122), .Z(n1325) );
XNOR2_X1 U1053 ( .A(KEYINPUT8), .B(KEYINPUT44), .ZN(n1327) );
NAND2_X1 U1054 ( .A1(G217), .A2(n1260), .ZN(n1322) );
AND2_X1 U1055 ( .A1(G234), .A2(n1085), .ZN(n1260) );
INV_X1 U1056 ( .A(G953), .ZN(n1085) );
XOR2_X1 U1057 ( .A(n1227), .B(n1328), .Z(n1319) );
XOR2_X1 U1058 ( .A(KEYINPUT60), .B(G134), .Z(n1328) );
INV_X1 U1059 ( .A(G128), .ZN(n1227) );
XNOR2_X1 U1060 ( .A(n1329), .B(G475), .ZN(n1249) );
OR2_X1 U1061 ( .A1(n1147), .A2(G902), .ZN(n1329) );
XOR2_X1 U1062 ( .A(n1330), .B(n1331), .Z(n1147) );
XOR2_X1 U1063 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1064 ( .A(G131), .B(G122), .Z(n1333) );
XOR2_X1 U1065 ( .A(KEYINPUT40), .B(KEYINPUT21), .Z(n1332) );
XOR2_X1 U1066 ( .A(n1334), .B(n1335), .Z(n1330) );
XOR2_X1 U1067 ( .A(n1244), .B(n1336), .Z(n1335) );
NAND2_X1 U1068 ( .A1(n1271), .A2(G214), .ZN(n1336) );
NOR2_X1 U1069 ( .A1(G953), .A2(G237), .ZN(n1271) );
INV_X1 U1070 ( .A(G113), .ZN(n1244) );
XNOR2_X1 U1071 ( .A(n1285), .B(n1257), .ZN(n1334) );
XOR2_X1 U1072 ( .A(n1103), .B(n1100), .Z(n1257) );
INV_X1 U1073 ( .A(G125), .ZN(n1100) );
INV_X1 U1074 ( .A(G140), .ZN(n1103) );
XNOR2_X1 U1075 ( .A(n1308), .B(n1110), .ZN(n1285) );
XNOR2_X1 U1076 ( .A(n1264), .B(n1300), .ZN(n1110) );
XOR2_X1 U1077 ( .A(G143), .B(KEYINPUT13), .Z(n1300) );
XNOR2_X1 U1078 ( .A(G146), .B(KEYINPUT53), .ZN(n1264) );
INV_X1 U1079 ( .A(G104), .ZN(n1308) );
INV_X1 U1080 ( .A(G110), .ZN(n1182) );
endmodule


