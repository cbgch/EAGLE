//Key = 0011101101111111000110110001101010101110011110111111101011101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366;

XNOR2_X1 U753 ( .A(G107), .B(n1034), .ZN(G9) );
NAND2_X1 U754 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U755 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR3_X1 U756 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NAND3_X1 U757 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1039) );
NAND2_X1 U758 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U759 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U760 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND2_X1 U761 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NAND2_X1 U762 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U763 ( .A(KEYINPUT18), .B(n1056), .Z(n1055) );
NAND2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
NAND2_X1 U765 ( .A1(n1058), .A2(n1059), .ZN(n1047) );
NAND3_X1 U766 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NAND2_X1 U767 ( .A1(n1049), .A2(n1063), .ZN(n1062) );
NAND2_X1 U768 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U769 ( .A1(n1056), .A2(n1066), .ZN(n1065) );
OR2_X1 U770 ( .A1(n1067), .A2(n1035), .ZN(n1066) );
NAND2_X1 U771 ( .A1(n1051), .A2(n1068), .ZN(n1064) );
NAND2_X1 U772 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND4_X1 U774 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1061) );
XOR2_X1 U775 ( .A(KEYINPUT40), .B(n1056), .Z(n1076) );
XOR2_X1 U776 ( .A(KEYINPUT25), .B(n1051), .Z(n1075) );
NAND3_X1 U777 ( .A1(n1056), .A2(n1077), .A3(n1051), .ZN(n1060) );
INV_X1 U778 ( .A(n1078), .ZN(n1045) );
NOR3_X1 U779 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1037) );
INV_X1 U780 ( .A(n1042), .ZN(n1079) );
NAND4_X1 U781 ( .A1(n1080), .A2(n1049), .A3(n1072), .A4(n1081), .ZN(n1042) );
XOR2_X1 U782 ( .A(n1082), .B(KEYINPUT37), .Z(n1080) );
NAND4_X1 U783 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
XOR2_X1 U784 ( .A(n1087), .B(KEYINPUT1), .Z(n1083) );
XOR2_X1 U785 ( .A(n1088), .B(n1089), .Z(G72) );
NOR2_X1 U786 ( .A1(n1090), .A2(n1043), .ZN(n1089) );
AND2_X1 U787 ( .A1(G227), .A2(G900), .ZN(n1090) );
NAND2_X1 U788 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
NAND2_X1 U789 ( .A1(n1093), .A2(n1043), .ZN(n1092) );
XOR2_X1 U790 ( .A(n1041), .B(n1094), .Z(n1093) );
NAND3_X1 U791 ( .A1(G900), .A2(n1094), .A3(G953), .ZN(n1091) );
XOR2_X1 U792 ( .A(n1095), .B(n1096), .Z(n1094) );
XNOR2_X1 U793 ( .A(n1097), .B(n1098), .ZN(n1095) );
NOR2_X1 U794 ( .A1(KEYINPUT0), .A2(n1099), .ZN(n1098) );
XOR2_X1 U795 ( .A(n1100), .B(n1101), .Z(G69) );
NOR2_X1 U796 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
AND4_X1 U797 ( .A1(n1104), .A2(G898), .A3(G953), .A4(G224), .ZN(n1103) );
NOR2_X1 U798 ( .A1(n1105), .A2(n1104), .ZN(n1102) );
INV_X1 U799 ( .A(KEYINPUT7), .ZN(n1104) );
NOR2_X1 U800 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U801 ( .A1(G224), .A2(n1043), .ZN(n1106) );
NAND2_X1 U802 ( .A1(KEYINPUT43), .A2(n1108), .ZN(n1100) );
XOR2_X1 U803 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U804 ( .A1(n1111), .A2(G953), .ZN(n1110) );
NOR3_X1 U805 ( .A1(n1107), .A2(n1112), .A3(n1113), .ZN(n1109) );
NOR3_X1 U806 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
NOR2_X1 U807 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
NOR2_X1 U808 ( .A1(n1115), .A2(n1116), .ZN(n1117) );
AND2_X1 U809 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
XNOR2_X1 U810 ( .A(n1121), .B(KEYINPUT2), .ZN(n1119) );
NOR2_X1 U811 ( .A1(n1122), .A2(n1123), .ZN(G66) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U813 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NOR3_X1 U814 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(G63) );
AND3_X1 U815 ( .A1(KEYINPUT55), .A2(G953), .A3(G952), .ZN(n1130) );
NOR2_X1 U816 ( .A1(KEYINPUT55), .A2(n1131), .ZN(n1129) );
XOR2_X1 U817 ( .A(n1132), .B(n1133), .Z(n1128) );
AND2_X1 U818 ( .A1(G478), .A2(n1134), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1122), .A2(n1135), .ZN(G60) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U821 ( .A1(n1134), .A2(G475), .ZN(n1137) );
NAND2_X1 U822 ( .A1(n1138), .A2(KEYINPUT32), .ZN(n1136) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U824 ( .A(G104), .B(n1141), .Z(G6) );
NOR2_X1 U825 ( .A1(n1142), .A2(n1143), .ZN(G57) );
XOR2_X1 U826 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U828 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U829 ( .A1(KEYINPUT5), .A2(n1150), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1144) );
AND2_X1 U831 ( .A1(G472), .A2(n1134), .ZN(n1152) );
XOR2_X1 U832 ( .A(n1153), .B(G101), .Z(n1151) );
XOR2_X1 U833 ( .A(n1131), .B(KEYINPUT30), .Z(n1142) );
INV_X1 U834 ( .A(n1122), .ZN(n1131) );
NOR2_X1 U835 ( .A1(n1122), .A2(n1154), .ZN(G54) );
XOR2_X1 U836 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U837 ( .A(n1157), .B(n1096), .Z(n1156) );
XOR2_X1 U838 ( .A(n1158), .B(n1159), .Z(n1157) );
AND2_X1 U839 ( .A1(G469), .A2(n1134), .ZN(n1159) );
INV_X1 U840 ( .A(n1127), .ZN(n1134) );
XOR2_X1 U841 ( .A(n1160), .B(n1161), .Z(n1155) );
XOR2_X1 U842 ( .A(G140), .B(G110), .Z(n1161) );
NAND3_X1 U843 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1160) );
OR2_X1 U844 ( .A1(n1165), .A2(KEYINPUT48), .ZN(n1164) );
NAND3_X1 U845 ( .A1(KEYINPUT48), .A2(n1166), .A3(n1099), .ZN(n1163) );
OR2_X1 U846 ( .A1(n1099), .A2(n1166), .ZN(n1162) );
AND2_X1 U847 ( .A1(KEYINPUT57), .A2(n1165), .ZN(n1166) );
XOR2_X1 U848 ( .A(n1167), .B(n1168), .Z(n1165) );
XNOR2_X1 U849 ( .A(n1169), .B(n1170), .ZN(n1099) );
NOR2_X1 U850 ( .A1(n1122), .A2(n1171), .ZN(G51) );
XOR2_X1 U851 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U852 ( .A1(n1174), .A2(n1127), .ZN(n1173) );
NAND2_X1 U853 ( .A1(G902), .A2(n1175), .ZN(n1127) );
NAND2_X1 U854 ( .A1(n1176), .A2(n1111), .ZN(n1175) );
INV_X1 U855 ( .A(n1040), .ZN(n1111) );
NAND4_X1 U856 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1040) );
NOR4_X1 U857 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1141), .ZN(n1180) );
AND2_X1 U858 ( .A1(n1067), .A2(n1036), .ZN(n1141) );
NOR2_X1 U859 ( .A1(n1184), .A2(n1185), .ZN(n1036) );
NOR3_X1 U860 ( .A1(n1186), .A2(n1184), .A3(n1187), .ZN(n1182) );
XOR2_X1 U861 ( .A(n1058), .B(KEYINPUT47), .Z(n1186) );
INV_X1 U862 ( .A(n1188), .ZN(n1181) );
NAND2_X1 U863 ( .A1(n1057), .A2(n1189), .ZN(n1179) );
NAND2_X1 U864 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND3_X1 U865 ( .A1(n1049), .A2(n1192), .A3(n1067), .ZN(n1191) );
INV_X1 U866 ( .A(n1193), .ZN(n1190) );
NAND2_X1 U867 ( .A1(n1194), .A2(n1193), .ZN(n1178) );
XOR2_X1 U868 ( .A(n1195), .B(KEYINPUT13), .Z(n1194) );
NAND2_X1 U869 ( .A1(n1196), .A2(n1197), .ZN(n1177) );
XNOR2_X1 U870 ( .A(n1198), .B(KEYINPUT62), .ZN(n1196) );
XOR2_X1 U871 ( .A(n1041), .B(KEYINPUT20), .Z(n1176) );
NAND4_X1 U872 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1041) );
AND4_X1 U873 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
NOR2_X1 U874 ( .A1(n1207), .A2(n1208), .ZN(n1201) );
NOR2_X1 U875 ( .A1(n1209), .A2(n1069), .ZN(n1208) );
XOR2_X1 U876 ( .A(n1210), .B(KEYINPUT63), .Z(n1209) );
NOR2_X1 U877 ( .A1(n1211), .A2(n1212), .ZN(n1172) );
XOR2_X1 U878 ( .A(n1213), .B(KEYINPUT41), .Z(n1212) );
NAND2_X1 U879 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U880 ( .A1(n1214), .A2(n1216), .ZN(n1211) );
XNOR2_X1 U881 ( .A(KEYINPUT44), .B(n1215), .ZN(n1216) );
NAND3_X1 U882 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1215) );
NAND2_X1 U883 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND3_X1 U884 ( .A1(n1222), .A2(n1146), .A3(G125), .ZN(n1218) );
NAND2_X1 U885 ( .A1(n1223), .A2(n1224), .ZN(n1217) );
XOR2_X1 U886 ( .A(n1146), .B(n1222), .Z(n1223) );
INV_X1 U887 ( .A(n1221), .ZN(n1222) );
NOR2_X1 U888 ( .A1(n1043), .A2(G952), .ZN(n1122) );
NAND2_X1 U889 ( .A1(n1225), .A2(n1226), .ZN(G48) );
NAND2_X1 U890 ( .A1(n1207), .A2(n1227), .ZN(n1226) );
XOR2_X1 U891 ( .A(KEYINPUT46), .B(n1228), .Z(n1225) );
NOR2_X1 U892 ( .A1(n1207), .A2(n1227), .ZN(n1228) );
AND3_X1 U893 ( .A1(n1067), .A2(n1197), .A3(n1229), .ZN(n1207) );
XOR2_X1 U894 ( .A(G143), .B(n1230), .Z(G45) );
NOR2_X1 U895 ( .A1(n1069), .A2(n1210), .ZN(n1230) );
NAND3_X1 U896 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1210) );
XOR2_X1 U897 ( .A(n1199), .B(n1234), .Z(G42) );
NAND2_X1 U898 ( .A1(KEYINPUT19), .A2(G140), .ZN(n1234) );
NAND3_X1 U899 ( .A1(n1235), .A2(n1077), .A3(n1056), .ZN(n1199) );
XNOR2_X1 U900 ( .A(G137), .B(n1200), .ZN(G39) );
NAND3_X1 U901 ( .A1(n1056), .A2(n1229), .A3(n1051), .ZN(n1200) );
XNOR2_X1 U902 ( .A(G134), .B(n1206), .ZN(G36) );
NAND3_X1 U903 ( .A1(n1233), .A2(n1035), .A3(n1056), .ZN(n1206) );
XNOR2_X1 U904 ( .A(G131), .B(n1205), .ZN(G33) );
NAND3_X1 U905 ( .A1(n1233), .A2(n1067), .A3(n1056), .ZN(n1205) );
AND2_X1 U906 ( .A1(n1072), .A2(n1236), .ZN(n1056) );
XOR2_X1 U907 ( .A(KEYINPUT50), .B(n1071), .Z(n1236) );
AND3_X1 U908 ( .A1(n1077), .A2(n1237), .A3(n1057), .ZN(n1233) );
XOR2_X1 U909 ( .A(n1238), .B(G128), .Z(G30) );
NAND2_X1 U910 ( .A1(KEYINPUT12), .A2(n1204), .ZN(n1238) );
NAND3_X1 U911 ( .A1(n1035), .A2(n1197), .A3(n1229), .ZN(n1204) );
AND4_X1 U912 ( .A1(n1239), .A2(n1077), .A3(n1240), .A4(n1237), .ZN(n1229) );
XOR2_X1 U913 ( .A(n1167), .B(n1241), .Z(G3) );
NAND4_X1 U914 ( .A1(n1051), .A2(n1057), .A3(KEYINPUT23), .A4(n1242), .ZN(n1241) );
NOR3_X1 U915 ( .A1(n1243), .A2(n1244), .A3(n1069), .ZN(n1242) );
XOR2_X1 U916 ( .A(n1245), .B(KEYINPUT36), .Z(n1244) );
INV_X1 U917 ( .A(n1077), .ZN(n1243) );
XOR2_X1 U918 ( .A(n1224), .B(n1203), .Z(G27) );
NAND3_X1 U919 ( .A1(n1049), .A2(n1197), .A3(n1235), .ZN(n1203) );
AND3_X1 U920 ( .A1(n1054), .A2(n1237), .A3(n1067), .ZN(n1235) );
NAND2_X1 U921 ( .A1(n1078), .A2(n1246), .ZN(n1237) );
NAND4_X1 U922 ( .A1(G902), .A2(G953), .A3(n1247), .A4(n1248), .ZN(n1246) );
INV_X1 U923 ( .A(G900), .ZN(n1248) );
XOR2_X1 U924 ( .A(n1249), .B(n1188), .Z(G24) );
NAND4_X1 U925 ( .A1(n1049), .A2(n1192), .A3(n1250), .A4(n1231), .ZN(n1188) );
NOR2_X1 U926 ( .A1(n1251), .A2(n1185), .ZN(n1250) );
INV_X1 U927 ( .A(n1058), .ZN(n1185) );
NAND2_X1 U928 ( .A1(n1252), .A2(n1253), .ZN(n1058) );
OR2_X1 U929 ( .A1(n1195), .A2(KEYINPUT10), .ZN(n1253) );
NAND3_X1 U930 ( .A1(n1254), .A2(n1084), .A3(KEYINPUT10), .ZN(n1252) );
INV_X1 U931 ( .A(n1239), .ZN(n1254) );
XOR2_X1 U932 ( .A(n1255), .B(n1256), .Z(G21) );
NAND2_X1 U933 ( .A1(KEYINPUT6), .A2(G119), .ZN(n1256) );
NAND2_X1 U934 ( .A1(n1198), .A2(n1197), .ZN(n1255) );
AND4_X1 U935 ( .A1(n1240), .A2(n1245), .A3(n1239), .A4(n1257), .ZN(n1198) );
AND2_X1 U936 ( .A1(n1049), .A2(n1051), .ZN(n1257) );
XOR2_X1 U937 ( .A(G116), .B(n1183), .Z(G18) );
AND3_X1 U938 ( .A1(n1035), .A2(n1197), .A3(n1258), .ZN(n1183) );
INV_X1 U939 ( .A(n1187), .ZN(n1035) );
NAND2_X1 U940 ( .A1(n1231), .A2(n1259), .ZN(n1187) );
XOR2_X1 U941 ( .A(KEYINPUT49), .B(n1232), .Z(n1259) );
XOR2_X1 U942 ( .A(n1260), .B(n1261), .Z(G15) );
NAND2_X1 U943 ( .A1(KEYINPUT15), .A2(n1262), .ZN(n1261) );
XOR2_X1 U944 ( .A(KEYINPUT53), .B(G113), .Z(n1262) );
NAND3_X1 U945 ( .A1(n1258), .A2(n1067), .A3(n1263), .ZN(n1260) );
XOR2_X1 U946 ( .A(n1069), .B(KEYINPUT38), .Z(n1263) );
INV_X1 U947 ( .A(n1197), .ZN(n1069) );
NOR2_X1 U948 ( .A1(n1251), .A2(n1231), .ZN(n1067) );
AND3_X1 U949 ( .A1(n1049), .A2(n1245), .A3(n1057), .ZN(n1258) );
AND2_X1 U950 ( .A1(n1264), .A2(n1240), .ZN(n1057) );
INV_X1 U951 ( .A(n1084), .ZN(n1240) );
XOR2_X1 U952 ( .A(n1239), .B(KEYINPUT10), .Z(n1264) );
NOR2_X1 U953 ( .A1(n1265), .A2(n1074), .ZN(n1049) );
INV_X1 U954 ( .A(n1073), .ZN(n1265) );
XNOR2_X1 U955 ( .A(G110), .B(n1266), .ZN(G12) );
NAND2_X1 U956 ( .A1(n1193), .A2(n1054), .ZN(n1266) );
INV_X1 U957 ( .A(n1195), .ZN(n1054) );
NAND2_X1 U958 ( .A1(n1239), .A2(n1084), .ZN(n1195) );
XOR2_X1 U959 ( .A(n1267), .B(G472), .Z(n1084) );
NAND2_X1 U960 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U961 ( .A(n1270), .B(n1271), .Z(n1268) );
XOR2_X1 U962 ( .A(n1272), .B(n1273), .Z(n1271) );
NOR2_X1 U963 ( .A1(KEYINPUT45), .A2(n1153), .ZN(n1272) );
NAND3_X1 U964 ( .A1(n1274), .A2(n1275), .A3(G210), .ZN(n1153) );
XOR2_X1 U965 ( .A(KEYINPUT9), .B(G953), .Z(n1274) );
XOR2_X1 U966 ( .A(n1276), .B(n1277), .Z(n1270) );
XOR2_X1 U967 ( .A(n1278), .B(G101), .Z(n1277) );
NAND2_X1 U968 ( .A1(KEYINPUT27), .A2(n1279), .ZN(n1278) );
XOR2_X1 U969 ( .A(KEYINPUT42), .B(n1096), .Z(n1279) );
INV_X1 U970 ( .A(n1148), .ZN(n1096) );
NAND2_X1 U971 ( .A1(KEYINPUT3), .A2(n1150), .ZN(n1276) );
XOR2_X1 U972 ( .A(G113), .B(n1280), .Z(n1150) );
NOR2_X1 U973 ( .A1(KEYINPUT35), .A2(n1281), .ZN(n1280) );
XOR2_X1 U974 ( .A(n1087), .B(KEYINPUT58), .Z(n1239) );
XOR2_X1 U975 ( .A(n1282), .B(n1283), .Z(n1087) );
NOR2_X1 U976 ( .A1(n1124), .A2(G902), .ZN(n1283) );
AND2_X1 U977 ( .A1(n1284), .A2(n1285), .ZN(n1124) );
NAND2_X1 U978 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U979 ( .A(KEYINPUT56), .B(n1288), .Z(n1284) );
NOR2_X1 U980 ( .A1(n1286), .A2(n1287), .ZN(n1288) );
XOR2_X1 U981 ( .A(n1289), .B(n1290), .Z(n1287) );
XOR2_X1 U982 ( .A(n1291), .B(n1097), .Z(n1290) );
XNOR2_X1 U983 ( .A(n1292), .B(G125), .ZN(n1097) );
NAND2_X1 U984 ( .A1(KEYINPUT34), .A2(n1227), .ZN(n1291) );
XOR2_X1 U985 ( .A(n1293), .B(n1294), .Z(n1289) );
NOR2_X1 U986 ( .A1(G110), .A2(KEYINPUT33), .ZN(n1294) );
XOR2_X1 U987 ( .A(G119), .B(n1169), .Z(n1293) );
XNOR2_X1 U988 ( .A(G137), .B(n1295), .ZN(n1286) );
NOR4_X1 U989 ( .A1(KEYINPUT31), .A2(G953), .A3(n1296), .A4(n1297), .ZN(n1295) );
NAND2_X1 U990 ( .A1(G217), .A2(n1298), .ZN(n1282) );
XOR2_X1 U991 ( .A(KEYINPUT22), .B(n1299), .Z(n1298) );
NOR2_X1 U992 ( .A1(n1300), .A2(n1184), .ZN(n1193) );
NAND2_X1 U993 ( .A1(n1077), .A2(n1192), .ZN(n1184) );
AND2_X1 U994 ( .A1(n1197), .A2(n1245), .ZN(n1192) );
NAND2_X1 U995 ( .A1(n1078), .A2(n1301), .ZN(n1245) );
NAND3_X1 U996 ( .A1(n1107), .A2(n1247), .A3(G902), .ZN(n1301) );
NOR2_X1 U997 ( .A1(n1043), .A2(G898), .ZN(n1107) );
NAND3_X1 U998 ( .A1(n1247), .A2(n1043), .A3(G952), .ZN(n1078) );
NAND2_X1 U999 ( .A1(G237), .A2(G234), .ZN(n1247) );
NOR2_X1 U1000 ( .A1(n1072), .A2(n1071), .ZN(n1197) );
INV_X1 U1001 ( .A(n1081), .ZN(n1071) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1302), .ZN(n1081) );
AND2_X1 U1003 ( .A1(n1303), .A2(n1304), .ZN(n1072) );
NAND2_X1 U1004 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND2_X1 U1005 ( .A1(n1307), .A2(n1269), .ZN(n1306) );
INV_X1 U1006 ( .A(n1174), .ZN(n1305) );
NAND3_X1 U1007 ( .A1(n1307), .A2(n1269), .A3(n1174), .ZN(n1303) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1302), .ZN(n1174) );
NAND2_X1 U1009 ( .A1(n1275), .A2(n1269), .ZN(n1302) );
XOR2_X1 U1010 ( .A(n1308), .B(n1221), .Z(n1307) );
NAND2_X1 U1011 ( .A1(n1309), .A2(n1043), .ZN(n1221) );
XOR2_X1 U1012 ( .A(KEYINPUT29), .B(G224), .Z(n1309) );
XNOR2_X1 U1013 ( .A(n1214), .B(n1310), .ZN(n1308) );
NOR3_X1 U1014 ( .A1(n1220), .A2(n1311), .A3(n1312), .ZN(n1310) );
NOR2_X1 U1015 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
INV_X1 U1016 ( .A(KEYINPUT60), .ZN(n1314) );
NOR2_X1 U1017 ( .A1(n1315), .A2(n1316), .ZN(n1313) );
AND2_X1 U1018 ( .A1(G125), .A2(KEYINPUT24), .ZN(n1316) );
NOR3_X1 U1019 ( .A1(KEYINPUT24), .A2(G125), .A3(n1273), .ZN(n1315) );
NOR2_X1 U1020 ( .A1(KEYINPUT60), .A2(n1317), .ZN(n1311) );
NOR2_X1 U1021 ( .A1(n1273), .A2(n1318), .ZN(n1317) );
XOR2_X1 U1022 ( .A(KEYINPUT24), .B(G125), .Z(n1318) );
INV_X1 U1023 ( .A(n1146), .ZN(n1273) );
NOR2_X1 U1024 ( .A1(n1224), .A2(n1146), .ZN(n1220) );
XOR2_X1 U1025 ( .A(n1319), .B(G128), .Z(n1146) );
NAND2_X1 U1026 ( .A1(KEYINPUT11), .A2(n1170), .ZN(n1319) );
AND2_X1 U1027 ( .A1(n1320), .A2(n1321), .ZN(n1214) );
NAND2_X1 U1028 ( .A1(n1114), .A2(n1322), .ZN(n1321) );
NAND2_X1 U1029 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1030 ( .A(n1325), .B(KEYINPUT26), .Z(n1320) );
NAND3_X1 U1031 ( .A1(n1323), .A2(n1324), .A3(n1118), .ZN(n1325) );
INV_X1 U1032 ( .A(n1114), .ZN(n1118) );
XNOR2_X1 U1033 ( .A(G110), .B(n1326), .ZN(n1114) );
XOR2_X1 U1034 ( .A(KEYINPUT52), .B(G122), .Z(n1326) );
INV_X1 U1035 ( .A(n1115), .ZN(n1324) );
NOR2_X1 U1036 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NAND2_X1 U1037 ( .A1(n1121), .A2(n1120), .ZN(n1323) );
NAND3_X1 U1038 ( .A1(n1327), .A2(n1328), .A3(n1329), .ZN(n1120) );
NAND2_X1 U1039 ( .A1(KEYINPUT21), .A2(n1168), .ZN(n1329) );
NAND3_X1 U1040 ( .A1(n1330), .A2(n1331), .A3(n1167), .ZN(n1328) );
INV_X1 U1041 ( .A(KEYINPUT21), .ZN(n1331) );
OR2_X1 U1042 ( .A1(n1167), .A2(n1330), .ZN(n1327) );
NOR2_X1 U1043 ( .A1(KEYINPUT39), .A2(n1168), .ZN(n1330) );
XNOR2_X1 U1044 ( .A(G104), .B(G107), .ZN(n1168) );
XNOR2_X1 U1045 ( .A(G113), .B(n1281), .ZN(n1121) );
XNOR2_X1 U1046 ( .A(G116), .B(G119), .ZN(n1281) );
NOR2_X1 U1047 ( .A1(n1073), .A2(n1074), .ZN(n1077) );
NOR2_X1 U1048 ( .A1(n1297), .A2(n1299), .ZN(n1074) );
NOR2_X1 U1049 ( .A1(n1296), .A2(G902), .ZN(n1299) );
INV_X1 U1050 ( .A(G221), .ZN(n1297) );
XOR2_X1 U1051 ( .A(n1332), .B(G469), .Z(n1073) );
NAND2_X1 U1052 ( .A1(n1333), .A2(n1269), .ZN(n1332) );
XOR2_X1 U1053 ( .A(n1148), .B(n1334), .Z(n1333) );
XOR2_X1 U1054 ( .A(n1335), .B(n1336), .Z(n1334) );
NAND2_X1 U1055 ( .A1(KEYINPUT28), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1056 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1057 ( .A(n1340), .B(n1167), .Z(n1339) );
INV_X1 U1058 ( .A(G101), .ZN(n1167) );
NAND2_X1 U1059 ( .A1(n1341), .A2(n1342), .ZN(n1335) );
NAND2_X1 U1060 ( .A1(n1158), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1061 ( .A(n1344), .B(n1345), .Z(n1341) );
NOR2_X1 U1062 ( .A1(KEYINPUT8), .A2(n1292), .ZN(n1345) );
XNOR2_X1 U1063 ( .A(G110), .B(n1346), .ZN(n1344) );
NOR2_X1 U1064 ( .A1(n1158), .A2(n1343), .ZN(n1346) );
INV_X1 U1065 ( .A(KEYINPUT4), .ZN(n1343) );
NAND2_X1 U1066 ( .A1(n1347), .A2(n1043), .ZN(n1158) );
INV_X1 U1067 ( .A(G953), .ZN(n1043) );
XOR2_X1 U1068 ( .A(KEYINPUT17), .B(G227), .Z(n1347) );
XNOR2_X1 U1069 ( .A(G131), .B(n1348), .ZN(n1148) );
XOR2_X1 U1070 ( .A(G137), .B(G134), .Z(n1348) );
INV_X1 U1071 ( .A(n1051), .ZN(n1300) );
NOR2_X1 U1072 ( .A1(n1232), .A2(n1231), .ZN(n1051) );
XOR2_X1 U1073 ( .A(n1085), .B(KEYINPUT54), .Z(n1231) );
XNOR2_X1 U1074 ( .A(G478), .B(n1349), .ZN(n1085) );
NOR2_X1 U1075 ( .A1(G902), .A2(n1133), .ZN(n1349) );
XNOR2_X1 U1076 ( .A(n1350), .B(n1351), .ZN(n1133) );
XOR2_X1 U1077 ( .A(n1338), .B(n1352), .Z(n1351) );
XOR2_X1 U1078 ( .A(n1353), .B(n1354), .Z(n1352) );
NOR3_X1 U1079 ( .A1(n1296), .A2(G953), .A3(n1126), .ZN(n1354) );
INV_X1 U1080 ( .A(G217), .ZN(n1126) );
INV_X1 U1081 ( .A(G234), .ZN(n1296) );
NAND2_X1 U1082 ( .A1(KEYINPUT51), .A2(n1355), .ZN(n1353) );
INV_X1 U1083 ( .A(G116), .ZN(n1355) );
XOR2_X1 U1084 ( .A(G107), .B(n1169), .Z(n1338) );
INV_X1 U1085 ( .A(G128), .ZN(n1169) );
XOR2_X1 U1086 ( .A(n1249), .B(n1356), .Z(n1350) );
XOR2_X1 U1087 ( .A(G143), .B(G134), .Z(n1356) );
INV_X1 U1088 ( .A(G122), .ZN(n1249) );
INV_X1 U1089 ( .A(n1251), .ZN(n1232) );
XOR2_X1 U1090 ( .A(n1086), .B(KEYINPUT16), .Z(n1251) );
XOR2_X1 U1091 ( .A(n1357), .B(G475), .Z(n1086) );
NAND2_X1 U1092 ( .A1(n1358), .A2(n1269), .ZN(n1357) );
INV_X1 U1093 ( .A(G902), .ZN(n1269) );
XOR2_X1 U1094 ( .A(n1359), .B(n1140), .Z(n1358) );
XNOR2_X1 U1095 ( .A(n1360), .B(n1340), .ZN(n1140) );
XNOR2_X1 U1096 ( .A(G104), .B(n1170), .ZN(n1340) );
XOR2_X1 U1097 ( .A(G143), .B(n1227), .Z(n1170) );
INV_X1 U1098 ( .A(G146), .ZN(n1227) );
XOR2_X1 U1099 ( .A(n1361), .B(n1362), .Z(n1360) );
NOR2_X1 U1100 ( .A1(KEYINPUT61), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1101 ( .A(n1224), .B(n1364), .Z(n1363) );
NOR2_X1 U1102 ( .A1(KEYINPUT59), .A2(n1292), .ZN(n1364) );
INV_X1 U1103 ( .A(G140), .ZN(n1292) );
INV_X1 U1104 ( .A(G125), .ZN(n1224) );
NAND3_X1 U1105 ( .A1(n1365), .A2(n1275), .A3(G214), .ZN(n1361) );
INV_X1 U1106 ( .A(G237), .ZN(n1275) );
XOR2_X1 U1107 ( .A(KEYINPUT14), .B(G953), .Z(n1365) );
INV_X1 U1108 ( .A(n1139), .ZN(n1359) );
XNOR2_X1 U1109 ( .A(G113), .B(n1366), .ZN(n1139) );
XOR2_X1 U1110 ( .A(G131), .B(G122), .Z(n1366) );
endmodule


