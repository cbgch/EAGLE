//Key = 0110100001010000101101011100110010101111100111101101100011100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269;

XOR2_X1 U704 ( .A(G107), .B(n968), .Z(G9) );
NOR2_X1 U705 ( .A1(n969), .A2(n970), .ZN(G75) );
XOR2_X1 U706 ( .A(n971), .B(KEYINPUT45), .Z(n970) );
OR3_X1 U707 ( .A1(G952), .A2(G953), .A3(n972), .ZN(n971) );
NOR4_X1 U708 ( .A1(n973), .A2(n974), .A3(G953), .A4(n972), .ZN(n969) );
AND4_X1 U709 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .ZN(n972) );
NOR4_X1 U710 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(n978) );
XOR2_X1 U711 ( .A(n983), .B(n984), .Z(n981) );
XOR2_X1 U712 ( .A(KEYINPUT49), .B(G478), .Z(n984) );
XOR2_X1 U713 ( .A(n985), .B(n986), .Z(n980) );
XOR2_X1 U714 ( .A(KEYINPUT1), .B(G469), .Z(n986) );
NOR2_X1 U715 ( .A1(n987), .A2(n988), .ZN(n977) );
NOR2_X1 U716 ( .A1(n989), .A2(n990), .ZN(n988) );
XOR2_X1 U717 ( .A(KEYINPUT8), .B(n991), .Z(n990) );
INV_X1 U718 ( .A(G475), .ZN(n989) );
NOR2_X1 U719 ( .A1(G475), .A2(n992), .ZN(n987) );
XOR2_X1 U720 ( .A(KEYINPUT63), .B(n991), .Z(n992) );
XOR2_X1 U721 ( .A(n993), .B(KEYINPUT42), .Z(n975) );
NOR2_X1 U722 ( .A1(n994), .A2(n995), .ZN(n974) );
NOR2_X1 U723 ( .A1(n996), .A2(n997), .ZN(n994) );
NOR2_X1 U724 ( .A1(n998), .A2(n999), .ZN(n997) );
INV_X1 U725 ( .A(n1000), .ZN(n999) );
NOR2_X1 U726 ( .A1(n1001), .A2(n1002), .ZN(n998) );
NOR4_X1 U727 ( .A1(n1003), .A2(n1004), .A3(n979), .A4(n1005), .ZN(n1002) );
NOR3_X1 U728 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1004) );
NOR2_X1 U729 ( .A1(n1009), .A2(n1010), .ZN(n1003) );
NOR4_X1 U730 ( .A1(n1011), .A2(n1012), .A3(n1006), .A4(n1013), .ZN(n1001) );
NOR3_X1 U731 ( .A1(n979), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR2_X1 U732 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U733 ( .A1(n976), .A2(n1018), .ZN(n1011) );
NOR3_X1 U734 ( .A1(n1005), .A2(n1019), .A3(n1013), .ZN(n996) );
NOR2_X1 U735 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
AND3_X1 U736 ( .A1(n1022), .A2(n1018), .A3(n1010), .ZN(n1020) );
NAND2_X1 U737 ( .A1(n1023), .A2(G952), .ZN(n973) );
XOR2_X1 U738 ( .A(n1024), .B(n1025), .Z(G72) );
XOR2_X1 U739 ( .A(n1026), .B(n1027), .Z(n1025) );
NAND3_X1 U740 ( .A1(n1028), .A2(n1029), .A3(KEYINPUT2), .ZN(n1027) );
NAND2_X1 U741 ( .A1(n1030), .A2(n1031), .ZN(n1026) );
NAND2_X1 U742 ( .A1(G953), .A2(n1032), .ZN(n1031) );
XOR2_X1 U743 ( .A(n1033), .B(n1034), .Z(n1030) );
XNOR2_X1 U744 ( .A(KEYINPUT62), .B(n1035), .ZN(n1033) );
NOR2_X1 U745 ( .A1(KEYINPUT53), .A2(n1036), .ZN(n1035) );
XOR2_X1 U746 ( .A(n1037), .B(KEYINPUT10), .Z(n1036) );
NOR3_X1 U747 ( .A1(n1029), .A2(KEYINPUT33), .A3(n1038), .ZN(n1024) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1032), .ZN(n1038) );
XOR2_X1 U749 ( .A(n1040), .B(n1041), .Z(G69) );
NOR2_X1 U750 ( .A1(n1042), .A2(n1029), .ZN(n1041) );
AND2_X1 U751 ( .A1(G224), .A2(G898), .ZN(n1042) );
NAND2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1040) );
NAND2_X1 U753 ( .A1(n1045), .A2(n1029), .ZN(n1044) );
XOR2_X1 U754 ( .A(n1046), .B(n1047), .Z(n1045) );
NAND3_X1 U755 ( .A1(n1046), .A2(G898), .A3(G953), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
INV_X1 U757 ( .A(KEYINPUT39), .ZN(n1048) );
NOR2_X1 U758 ( .A1(n1050), .A2(n1051), .ZN(G66) );
XOR2_X1 U759 ( .A(n1052), .B(n1053), .Z(n1051) );
NOR2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U761 ( .A1(n1050), .A2(n1056), .ZN(G63) );
XOR2_X1 U762 ( .A(n1057), .B(n1058), .Z(n1056) );
XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n1059), .ZN(n1058) );
NAND2_X1 U764 ( .A1(n1060), .A2(G478), .ZN(n1057) );
NOR2_X1 U765 ( .A1(n1050), .A2(n1061), .ZN(G60) );
XOR2_X1 U766 ( .A(n1062), .B(n1063), .Z(n1061) );
NOR2_X1 U767 ( .A1(KEYINPUT22), .A2(n1064), .ZN(n1063) );
NAND2_X1 U768 ( .A1(n1060), .A2(G475), .ZN(n1062) );
XOR2_X1 U769 ( .A(n1065), .B(n1066), .Z(G6) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1014), .ZN(n1066) );
XOR2_X1 U771 ( .A(n1068), .B(KEYINPUT34), .Z(n1067) );
NOR2_X1 U772 ( .A1(n1050), .A2(n1069), .ZN(G57) );
XOR2_X1 U773 ( .A(n1070), .B(n1071), .Z(n1069) );
XOR2_X1 U774 ( .A(n1072), .B(n1073), .Z(n1071) );
XOR2_X1 U775 ( .A(n1074), .B(n1075), .Z(n1070) );
XNOR2_X1 U776 ( .A(n1076), .B(KEYINPUT44), .ZN(n1075) );
NAND2_X1 U777 ( .A1(KEYINPUT57), .A2(n1077), .ZN(n1076) );
AND2_X1 U778 ( .A1(G472), .A2(n1060), .ZN(n1074) );
NOR2_X1 U779 ( .A1(n1050), .A2(n1078), .ZN(G54) );
XOR2_X1 U780 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U781 ( .A1(KEYINPUT20), .A2(n1081), .ZN(n1080) );
NAND2_X1 U782 ( .A1(n1060), .A2(G469), .ZN(n1079) );
NOR2_X1 U783 ( .A1(n1029), .A2(G952), .ZN(n1050) );
NOR2_X1 U784 ( .A1(n1082), .A2(n1083), .ZN(G51) );
XOR2_X1 U785 ( .A(n1084), .B(n1085), .Z(n1083) );
XOR2_X1 U786 ( .A(n1086), .B(n1049), .Z(n1085) );
NOR2_X1 U787 ( .A1(n1087), .A2(n1055), .ZN(n1086) );
INV_X1 U788 ( .A(n1060), .ZN(n1055) );
NOR2_X1 U789 ( .A1(n1088), .A2(n1023), .ZN(n1060) );
NOR2_X1 U790 ( .A1(n1047), .A2(n1028), .ZN(n1023) );
NAND4_X1 U791 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1028) );
AND4_X1 U792 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1092) );
NOR2_X1 U793 ( .A1(n1097), .A2(n1098), .ZN(n1091) );
NOR2_X1 U794 ( .A1(n1005), .A2(n1099), .ZN(n1098) );
NOR2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
XOR2_X1 U796 ( .A(n1102), .B(KEYINPUT15), .Z(n1100) );
NAND2_X1 U797 ( .A1(n1103), .A2(n1104), .ZN(n1089) );
XNOR2_X1 U798 ( .A(n1007), .B(KEYINPUT19), .ZN(n1103) );
NAND4_X1 U799 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1047) );
NOR4_X1 U800 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n968), .ZN(n1108) );
AND4_X1 U801 ( .A1(n1112), .A2(n1022), .A3(n1006), .A4(n1009), .ZN(n968) );
NAND2_X1 U802 ( .A1(n1014), .A2(n1113), .ZN(n1107) );
NAND2_X1 U803 ( .A1(n1068), .A2(n1114), .ZN(n1113) );
NAND3_X1 U804 ( .A1(n1007), .A2(n1115), .A3(n1021), .ZN(n1114) );
NAND4_X1 U805 ( .A1(n1116), .A2(n1009), .A3(n1117), .A4(n1006), .ZN(n1068) );
NOR2_X1 U806 ( .A1(n1118), .A2(n979), .ZN(n1117) );
NOR2_X1 U807 ( .A1(n1119), .A2(n1120), .ZN(n1084) );
NOR2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XNOR2_X1 U809 ( .A(n1123), .B(n1124), .ZN(n1122) );
XOR2_X1 U810 ( .A(KEYINPUT46), .B(KEYINPUT24), .Z(n1124) );
NOR2_X1 U811 ( .A1(n1125), .A2(n1123), .ZN(n1119) );
XNOR2_X1 U812 ( .A(n1126), .B(n1127), .ZN(n1123) );
NOR2_X1 U813 ( .A1(KEYINPUT47), .A2(n1128), .ZN(n1127) );
NOR2_X1 U814 ( .A1(G952), .A2(n1129), .ZN(n1082) );
XOR2_X1 U815 ( .A(KEYINPUT32), .B(G953), .Z(n1129) );
XOR2_X1 U816 ( .A(n1093), .B(n1130), .Z(G48) );
XNOR2_X1 U817 ( .A(G146), .B(KEYINPUT14), .ZN(n1130) );
NAND3_X1 U818 ( .A1(n1116), .A2(n1014), .A3(n1131), .ZN(n1093) );
XOR2_X1 U819 ( .A(G143), .B(n1132), .Z(G45) );
NOR2_X1 U820 ( .A1(n1101), .A2(n1102), .ZN(n1132) );
NAND4_X1 U821 ( .A1(n1133), .A2(n1007), .A3(n1134), .A4(n1135), .ZN(n1102) );
XNOR2_X1 U822 ( .A(G140), .B(n1090), .ZN(G42) );
NAND2_X1 U823 ( .A1(n1104), .A2(n1008), .ZN(n1090) );
XOR2_X1 U824 ( .A(G137), .B(n1136), .Z(G39) );
NOR3_X1 U825 ( .A1(n1137), .A2(KEYINPUT7), .A3(n1005), .ZN(n1136) );
XNOR2_X1 U826 ( .A(KEYINPUT48), .B(n1099), .ZN(n1137) );
NAND2_X1 U827 ( .A1(n1131), .A2(n1000), .ZN(n1099) );
XOR2_X1 U828 ( .A(G134), .B(n1138), .Z(G36) );
NOR2_X1 U829 ( .A1(KEYINPUT26), .A2(n1096), .ZN(n1138) );
NAND4_X1 U830 ( .A1(n1133), .A2(n1007), .A3(n976), .A4(n1022), .ZN(n1096) );
XOR2_X1 U831 ( .A(G131), .B(n1139), .Z(G33) );
AND2_X1 U832 ( .A1(n1007), .A2(n1104), .ZN(n1139) );
AND3_X1 U833 ( .A1(n1116), .A2(n976), .A3(n1133), .ZN(n1104) );
INV_X1 U834 ( .A(n1005), .ZN(n976) );
NAND2_X1 U835 ( .A1(n1140), .A2(n1017), .ZN(n1005) );
INV_X1 U836 ( .A(n1016), .ZN(n1140) );
XOR2_X1 U837 ( .A(n1141), .B(G128), .Z(G30) );
NAND2_X1 U838 ( .A1(KEYINPUT18), .A2(n1095), .ZN(n1141) );
NAND3_X1 U839 ( .A1(n1022), .A2(n1014), .A3(n1131), .ZN(n1095) );
AND3_X1 U840 ( .A1(n1142), .A2(n982), .A3(n1133), .ZN(n1131) );
AND3_X1 U841 ( .A1(n1018), .A2(n1143), .A3(n1006), .ZN(n1133) );
NAND2_X1 U842 ( .A1(n1144), .A2(n1145), .ZN(G3) );
NAND2_X1 U843 ( .A1(n1111), .A2(n1146), .ZN(n1145) );
XOR2_X1 U844 ( .A(KEYINPUT23), .B(n1147), .Z(n1144) );
NOR2_X1 U845 ( .A1(n1111), .A2(n1146), .ZN(n1147) );
AND2_X1 U846 ( .A1(n1007), .A2(n1148), .ZN(n1111) );
XOR2_X1 U847 ( .A(n1128), .B(n1094), .Z(G27) );
NAND4_X1 U848 ( .A1(n1021), .A2(n1008), .A3(n1014), .A4(n1143), .ZN(n1094) );
NAND2_X1 U849 ( .A1(n1149), .A2(n995), .ZN(n1143) );
NAND2_X1 U850 ( .A1(n1150), .A2(n1032), .ZN(n1149) );
INV_X1 U851 ( .A(G900), .ZN(n1032) );
INV_X1 U852 ( .A(G125), .ZN(n1128) );
XNOR2_X1 U853 ( .A(G122), .B(n1105), .ZN(G24) );
NAND3_X1 U854 ( .A1(n1112), .A2(n1009), .A3(n1151), .ZN(n1105) );
NOR3_X1 U855 ( .A1(n1152), .A2(n1006), .A3(n1153), .ZN(n1151) );
INV_X1 U856 ( .A(n1013), .ZN(n1009) );
NAND2_X1 U857 ( .A1(n1154), .A2(n993), .ZN(n1013) );
XNOR2_X1 U858 ( .A(n1155), .B(n1106), .ZN(G21) );
NAND3_X1 U859 ( .A1(n1000), .A2(n1112), .A3(n1156), .ZN(n1106) );
NOR3_X1 U860 ( .A1(n1006), .A2(n1154), .A3(n993), .ZN(n1156) );
NAND2_X1 U861 ( .A1(KEYINPUT51), .A2(n1157), .ZN(n1155) );
XOR2_X1 U862 ( .A(n1110), .B(n1158), .Z(G18) );
NOR2_X1 U863 ( .A1(KEYINPUT59), .A2(n1159), .ZN(n1158) );
INV_X1 U864 ( .A(G116), .ZN(n1159) );
AND4_X1 U865 ( .A1(n1007), .A2(n1112), .A3(n1022), .A4(n1010), .ZN(n1110) );
NOR2_X1 U866 ( .A1(n1135), .A2(n1152), .ZN(n1022) );
INV_X1 U867 ( .A(n1134), .ZN(n1152) );
XOR2_X1 U868 ( .A(n1160), .B(KEYINPUT6), .Z(n1134) );
XNOR2_X1 U869 ( .A(G113), .B(n1161), .ZN(G15) );
NAND4_X1 U870 ( .A1(n1162), .A2(n1021), .A3(n1007), .A4(n1014), .ZN(n1161) );
INV_X1 U871 ( .A(n1101), .ZN(n1014) );
NOR2_X1 U872 ( .A1(n982), .A2(n993), .ZN(n1007) );
AND3_X1 U873 ( .A1(n1010), .A2(n1018), .A3(n1116), .ZN(n1021) );
NOR2_X1 U874 ( .A1(n1160), .A2(n1153), .ZN(n1116) );
INV_X1 U875 ( .A(n1006), .ZN(n1010) );
XOR2_X1 U876 ( .A(n1115), .B(KEYINPUT17), .Z(n1162) );
XOR2_X1 U877 ( .A(G110), .B(n1109), .Z(G12) );
AND2_X1 U878 ( .A1(n1148), .A2(n1008), .ZN(n1109) );
NOR2_X1 U879 ( .A1(n1142), .A2(n1154), .ZN(n1008) );
INV_X1 U880 ( .A(n982), .ZN(n1154) );
NAND3_X1 U881 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n982) );
NAND2_X1 U882 ( .A1(n1052), .A2(n1166), .ZN(n1165) );
OR3_X1 U883 ( .A1(n1166), .A2(n1052), .A3(G902), .ZN(n1164) );
AND2_X1 U884 ( .A1(n1167), .A2(n1168), .ZN(n1052) );
NAND2_X1 U885 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U886 ( .A(n1171), .B(KEYINPUT27), .Z(n1167) );
OR2_X1 U887 ( .A1(n1170), .A2(n1169), .ZN(n1171) );
XOR2_X1 U888 ( .A(n1172), .B(n1173), .Z(n1169) );
XOR2_X1 U889 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U890 ( .A1(KEYINPUT58), .A2(n1176), .ZN(n1175) );
XOR2_X1 U891 ( .A(G128), .B(G119), .Z(n1176) );
INV_X1 U892 ( .A(G110), .ZN(n1174) );
NAND2_X1 U893 ( .A1(KEYINPUT43), .A2(n1177), .ZN(n1172) );
XOR2_X1 U894 ( .A(n1178), .B(n1034), .Z(n1177) );
XNOR2_X1 U895 ( .A(n1179), .B(G137), .ZN(n1170) );
NAND3_X1 U896 ( .A1(G234), .A2(n1029), .A3(G221), .ZN(n1179) );
NOR2_X1 U897 ( .A1(n1054), .A2(G234), .ZN(n1166) );
INV_X1 U898 ( .A(G217), .ZN(n1054) );
NAND2_X1 U899 ( .A1(G217), .A2(G902), .ZN(n1163) );
INV_X1 U900 ( .A(n993), .ZN(n1142) );
XOR2_X1 U901 ( .A(n1180), .B(G472), .Z(n993) );
NAND2_X1 U902 ( .A1(n1181), .A2(n1088), .ZN(n1180) );
XNOR2_X1 U903 ( .A(n1077), .B(n1182), .ZN(n1181) );
XOR2_X1 U904 ( .A(n1183), .B(n1072), .Z(n1182) );
XNOR2_X1 U905 ( .A(n1184), .B(n1185), .ZN(n1072) );
XOR2_X1 U906 ( .A(n1146), .B(n1186), .Z(n1185) );
NAND2_X1 U907 ( .A1(n1187), .A2(G210), .ZN(n1186) );
INV_X1 U908 ( .A(G101), .ZN(n1146) );
NAND2_X1 U909 ( .A1(KEYINPUT29), .A2(n1073), .ZN(n1183) );
XNOR2_X1 U910 ( .A(n1188), .B(n1189), .ZN(n1073) );
NOR2_X1 U911 ( .A1(G113), .A2(KEYINPUT5), .ZN(n1189) );
XNOR2_X1 U912 ( .A(n1126), .B(KEYINPUT13), .ZN(n1077) );
AND3_X1 U913 ( .A1(n1006), .A2(n1112), .A3(n1000), .ZN(n1148) );
NOR2_X1 U914 ( .A1(n1135), .A2(n1160), .ZN(n1000) );
NAND3_X1 U915 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1160) );
NAND2_X1 U916 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U917 ( .A(G478), .ZN(n1194) );
NAND2_X1 U918 ( .A1(KEYINPUT61), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U919 ( .A(KEYINPUT36), .B(n983), .ZN(n1195) );
NAND3_X1 U920 ( .A1(KEYINPUT61), .A2(G478), .A3(n983), .ZN(n1191) );
OR2_X1 U921 ( .A1(n983), .A2(KEYINPUT61), .ZN(n1190) );
NAND2_X1 U922 ( .A1(n1088), .A2(n1059), .ZN(n983) );
NAND3_X1 U923 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1059) );
NAND2_X1 U924 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U925 ( .A1(n1201), .A2(KEYINPUT16), .ZN(n1200) );
XNOR2_X1 U926 ( .A(n1202), .B(KEYINPUT38), .ZN(n1201) );
NAND3_X1 U927 ( .A1(KEYINPUT16), .A2(n1203), .A3(n1202), .ZN(n1197) );
INV_X1 U928 ( .A(n1199), .ZN(n1203) );
XOR2_X1 U929 ( .A(n1204), .B(n1205), .Z(n1199) );
XOR2_X1 U930 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U931 ( .A(G128), .B(G116), .Z(n1207) );
XOR2_X1 U932 ( .A(KEYINPUT50), .B(G143), .Z(n1206) );
XNOR2_X1 U933 ( .A(n1208), .B(n1209), .ZN(n1204) );
XOR2_X1 U934 ( .A(G107), .B(n1210), .Z(n1209) );
NOR2_X1 U935 ( .A1(KEYINPUT31), .A2(n1211), .ZN(n1210) );
INV_X1 U936 ( .A(G134), .ZN(n1211) );
OR2_X1 U937 ( .A1(n1202), .A2(KEYINPUT16), .ZN(n1196) );
AND3_X1 U938 ( .A1(G234), .A2(n1029), .A3(G217), .ZN(n1202) );
INV_X1 U939 ( .A(n1153), .ZN(n1135) );
XOR2_X1 U940 ( .A(n1212), .B(G475), .Z(n1153) );
NAND2_X1 U941 ( .A1(KEYINPUT40), .A2(n991), .ZN(n1212) );
NOR2_X1 U942 ( .A1(n1064), .A2(G902), .ZN(n991) );
XNOR2_X1 U943 ( .A(n1213), .B(n1214), .ZN(n1064) );
XOR2_X1 U944 ( .A(n1215), .B(n1216), .Z(n1214) );
XOR2_X1 U945 ( .A(G104), .B(n1217), .Z(n1216) );
NOR2_X1 U946 ( .A1(KEYINPUT3), .A2(n1218), .ZN(n1217) );
XNOR2_X1 U947 ( .A(G113), .B(n1219), .ZN(n1218) );
NAND2_X1 U948 ( .A1(KEYINPUT4), .A2(n1208), .ZN(n1219) );
XOR2_X1 U949 ( .A(G143), .B(G131), .Z(n1215) );
XNOR2_X1 U950 ( .A(n1034), .B(n1220), .ZN(n1213) );
XNOR2_X1 U951 ( .A(n1221), .B(n1222), .ZN(n1220) );
AND3_X1 U952 ( .A1(n1187), .A2(n1223), .A3(G214), .ZN(n1222) );
INV_X1 U953 ( .A(KEYINPUT0), .ZN(n1223) );
NOR2_X1 U954 ( .A1(G953), .A2(G237), .ZN(n1187) );
NAND2_X1 U955 ( .A1(KEYINPUT56), .A2(n1224), .ZN(n1221) );
XOR2_X1 U956 ( .A(G140), .B(G125), .Z(n1034) );
NOR3_X1 U957 ( .A1(n979), .A2(n1118), .A3(n1101), .ZN(n1112) );
NAND2_X1 U958 ( .A1(n1016), .A2(n1017), .ZN(n1101) );
NAND2_X1 U959 ( .A1(G214), .A2(n1225), .ZN(n1017) );
NAND2_X1 U960 ( .A1(n1226), .A2(n1088), .ZN(n1225) );
NAND3_X1 U961 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1016) );
NAND2_X1 U962 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
OR3_X1 U963 ( .A1(n1231), .A2(n1230), .A3(G902), .ZN(n1228) );
NOR2_X1 U964 ( .A1(n1087), .A2(n1226), .ZN(n1230) );
INV_X1 U965 ( .A(G237), .ZN(n1226) );
INV_X1 U966 ( .A(G210), .ZN(n1087) );
XNOR2_X1 U967 ( .A(n1232), .B(n1233), .ZN(n1231) );
XOR2_X1 U968 ( .A(G125), .B(n1125), .Z(n1233) );
INV_X1 U969 ( .A(n1121), .ZN(n1125) );
NAND2_X1 U970 ( .A1(G224), .A2(n1029), .ZN(n1121) );
XNOR2_X1 U971 ( .A(n1049), .B(n1234), .ZN(n1232) );
NOR2_X1 U972 ( .A1(KEYINPUT60), .A2(n1126), .ZN(n1234) );
XOR2_X1 U973 ( .A(n1235), .B(n1236), .Z(n1126) );
NOR2_X1 U974 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NOR2_X1 U975 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
XOR2_X1 U976 ( .A(KEYINPUT30), .B(n1178), .Z(n1240) );
XNOR2_X1 U977 ( .A(n1241), .B(n1242), .ZN(n1049) );
XNOR2_X1 U978 ( .A(n1188), .B(n1208), .ZN(n1242) );
XOR2_X1 U979 ( .A(G122), .B(KEYINPUT9), .Z(n1208) );
XOR2_X1 U980 ( .A(G116), .B(n1157), .Z(n1188) );
INV_X1 U981 ( .A(G119), .ZN(n1157) );
XOR2_X1 U982 ( .A(n1243), .B(n1244), .Z(n1241) );
XNOR2_X1 U983 ( .A(KEYINPUT35), .B(n1245), .ZN(n1243) );
NOR2_X1 U984 ( .A1(G113), .A2(KEYINPUT41), .ZN(n1245) );
NAND2_X1 U985 ( .A1(G210), .A2(G902), .ZN(n1227) );
INV_X1 U986 ( .A(n1115), .ZN(n1118) );
NAND2_X1 U987 ( .A1(n1246), .A2(n995), .ZN(n1115) );
NAND3_X1 U988 ( .A1(n1247), .A2(n1029), .A3(n1248), .ZN(n995) );
XNOR2_X1 U989 ( .A(G952), .B(KEYINPUT37), .ZN(n1248) );
INV_X1 U990 ( .A(G953), .ZN(n1029) );
NAND2_X1 U991 ( .A1(n1150), .A2(n1249), .ZN(n1246) );
INV_X1 U992 ( .A(G898), .ZN(n1249) );
AND3_X1 U993 ( .A1(G902), .A2(n1247), .A3(G953), .ZN(n1150) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1247) );
INV_X1 U995 ( .A(n1018), .ZN(n979) );
NAND2_X1 U996 ( .A1(G221), .A2(n1250), .ZN(n1018) );
NAND2_X1 U997 ( .A1(G234), .A2(n1088), .ZN(n1250) );
INV_X1 U998 ( .A(G902), .ZN(n1088) );
XOR2_X1 U999 ( .A(n1251), .B(G469), .Z(n1006) );
NAND2_X1 U1000 ( .A1(KEYINPUT52), .A2(n985), .ZN(n1251) );
NAND2_X1 U1001 ( .A1(n1252), .A2(n1253), .ZN(n985) );
XOR2_X1 U1002 ( .A(KEYINPUT11), .B(G902), .Z(n1253) );
INV_X1 U1003 ( .A(n1081), .ZN(n1252) );
XOR2_X1 U1004 ( .A(n1254), .B(n1255), .Z(n1081) );
XOR2_X1 U1005 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U1006 ( .A(KEYINPUT25), .B(G140), .Z(n1257) );
NOR2_X1 U1007 ( .A1(G953), .A2(n1039), .ZN(n1256) );
INV_X1 U1008 ( .A(G227), .ZN(n1039) );
XOR2_X1 U1009 ( .A(n1037), .B(n1244), .Z(n1254) );
XNOR2_X1 U1010 ( .A(n1258), .B(n1259), .ZN(n1244) );
XOR2_X1 U1011 ( .A(G110), .B(G107), .Z(n1259) );
XOR2_X1 U1012 ( .A(n1065), .B(G101), .Z(n1258) );
INV_X1 U1013 ( .A(G104), .ZN(n1065) );
XOR2_X1 U1014 ( .A(n1260), .B(n1261), .Z(n1037) );
NOR2_X1 U1015 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NOR2_X1 U1016 ( .A1(KEYINPUT55), .A2(n1264), .ZN(n1263) );
XOR2_X1 U1017 ( .A(G143), .B(n1178), .Z(n1264) );
NOR2_X1 U1018 ( .A1(n1265), .A2(n1266), .ZN(n1262) );
INV_X1 U1019 ( .A(KEYINPUT55), .ZN(n1266) );
NOR2_X1 U1020 ( .A1(n1267), .A2(n1238), .ZN(n1265) );
NOR2_X1 U1021 ( .A1(n1224), .A2(G143), .ZN(n1238) );
NOR2_X1 U1022 ( .A1(n1178), .A2(n1239), .ZN(n1267) );
INV_X1 U1023 ( .A(G143), .ZN(n1239) );
INV_X1 U1024 ( .A(n1224), .ZN(n1178) );
XNOR2_X1 U1025 ( .A(G146), .B(KEYINPUT54), .ZN(n1224) );
XNOR2_X1 U1026 ( .A(n1268), .B(n1184), .ZN(n1260) );
XNOR2_X1 U1027 ( .A(G131), .B(n1269), .ZN(n1184) );
XOR2_X1 U1028 ( .A(G137), .B(G134), .Z(n1269) );
NAND2_X1 U1029 ( .A1(KEYINPUT28), .A2(n1235), .ZN(n1268) );
XNOR2_X1 U1030 ( .A(G128), .B(KEYINPUT12), .ZN(n1235) );
endmodule


