//Key = 1000011001100000011011101011101100100010100001101100010110110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268;

XOR2_X1 U696 ( .A(G107), .B(n961), .Z(G9) );
NOR2_X1 U697 ( .A1(n962), .A2(n963), .ZN(G75) );
NOR3_X1 U698 ( .A1(n964), .A2(n965), .A3(n966), .ZN(n963) );
NOR2_X1 U699 ( .A1(n967), .A2(n968), .ZN(n965) );
NOR2_X1 U700 ( .A1(n969), .A2(n970), .ZN(n967) );
XOR2_X1 U701 ( .A(KEYINPUT32), .B(n971), .Z(n970) );
NOR4_X1 U702 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(n971) );
NAND2_X1 U703 ( .A1(n976), .A2(n977), .ZN(n973) );
XOR2_X1 U704 ( .A(KEYINPUT23), .B(n978), .Z(n976) );
AND4_X1 U705 ( .A1(n979), .A2(n980), .A3(n981), .A4(n978), .ZN(n969) );
NAND3_X1 U706 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n964) );
NAND3_X1 U707 ( .A1(n985), .A2(n986), .A3(n978), .ZN(n984) );
INV_X1 U708 ( .A(n987), .ZN(n978) );
NAND2_X1 U709 ( .A1(n988), .A2(n989), .ZN(n986) );
NAND2_X1 U710 ( .A1(n980), .A2(n990), .ZN(n989) );
NAND3_X1 U711 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n990) );
NAND2_X1 U712 ( .A1(n994), .A2(n995), .ZN(n993) );
XOR2_X1 U713 ( .A(n974), .B(KEYINPUT53), .Z(n994) );
NAND3_X1 U714 ( .A1(n996), .A2(n981), .A3(n997), .ZN(n992) );
NAND2_X1 U715 ( .A1(n998), .A2(n999), .ZN(n991) );
NAND2_X1 U716 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND2_X1 U717 ( .A1(n981), .A2(n1002), .ZN(n988) );
NAND2_X1 U718 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U719 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
XOR2_X1 U720 ( .A(n968), .B(KEYINPUT27), .Z(n1005) );
INV_X1 U721 ( .A(n998), .ZN(n968) );
NAND2_X1 U722 ( .A1(n998), .A2(n1007), .ZN(n1003) );
NOR3_X1 U723 ( .A1(n1008), .A2(G953), .A3(G952), .ZN(n962) );
INV_X1 U724 ( .A(n982), .ZN(n1008) );
NAND4_X1 U725 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n982) );
NOR4_X1 U726 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
XOR2_X1 U727 ( .A(G469), .B(n1017), .Z(n1016) );
XOR2_X1 U728 ( .A(KEYINPUT57), .B(n1018), .Z(n1015) );
XOR2_X1 U729 ( .A(KEYINPUT11), .B(n1019), .Z(n1014) );
XOR2_X1 U730 ( .A(KEYINPUT54), .B(n1020), .Z(n1013) );
NOR3_X1 U731 ( .A1(n1021), .A2(n1022), .A3(n997), .ZN(n1011) );
XNOR2_X1 U732 ( .A(KEYINPUT56), .B(n1023), .ZN(n1010) );
XOR2_X1 U733 ( .A(n1024), .B(G475), .Z(n1009) );
NAND2_X1 U734 ( .A1(n1025), .A2(n1026), .ZN(G72) );
NAND2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XNOR2_X1 U736 ( .A(n1029), .B(n1030), .ZN(n1028) );
NAND2_X1 U737 ( .A1(KEYINPUT26), .A2(n1031), .ZN(n1029) );
NAND2_X1 U738 ( .A1(n983), .A2(n1032), .ZN(n1031) );
NAND2_X1 U739 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
XOR2_X1 U740 ( .A(n1035), .B(KEYINPUT39), .Z(n1033) );
XOR2_X1 U741 ( .A(n1036), .B(KEYINPUT2), .Z(n1027) );
XOR2_X1 U742 ( .A(KEYINPUT61), .B(n1037), .Z(n1025) );
NOR2_X1 U743 ( .A1(n1038), .A2(n1036), .ZN(n1037) );
NAND2_X1 U744 ( .A1(n1039), .A2(G953), .ZN(n1036) );
XOR2_X1 U745 ( .A(n1040), .B(KEYINPUT62), .Z(n1039) );
NAND2_X1 U746 ( .A1(G900), .A2(G227), .ZN(n1040) );
XOR2_X1 U747 ( .A(n1030), .B(KEYINPUT26), .Z(n1038) );
NAND2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1030) );
NAND2_X1 U749 ( .A1(G953), .A2(n1043), .ZN(n1042) );
XOR2_X1 U750 ( .A(n1044), .B(n1045), .Z(n1041) );
XOR2_X1 U751 ( .A(n1046), .B(n1047), .Z(n1045) );
NOR2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U753 ( .A(n1050), .B(KEYINPUT28), .Z(n1049) );
NAND2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1051), .ZN(n1048) );
XOR2_X1 U756 ( .A(G134), .B(n1053), .Z(n1051) );
XOR2_X1 U757 ( .A(KEYINPUT46), .B(G137), .Z(n1053) );
NOR2_X1 U758 ( .A1(KEYINPUT52), .A2(n1054), .ZN(n1046) );
XOR2_X1 U759 ( .A(n1055), .B(n1056), .Z(G69) );
XOR2_X1 U760 ( .A(n1057), .B(n1058), .Z(n1056) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U762 ( .A(n1061), .B(n1062), .Z(n1060) );
XOR2_X1 U763 ( .A(KEYINPUT9), .B(n1063), .Z(n1062) );
NOR2_X1 U764 ( .A1(KEYINPUT51), .A2(n1064), .ZN(n1063) );
XOR2_X1 U765 ( .A(n1065), .B(n1066), .Z(n1061) );
NOR2_X1 U766 ( .A1(G898), .A2(n983), .ZN(n1059) );
NAND2_X1 U767 ( .A1(n1067), .A2(n983), .ZN(n1057) );
XOR2_X1 U768 ( .A(KEYINPUT40), .B(n1068), .Z(n1067) );
NAND2_X1 U769 ( .A1(G953), .A2(n1069), .ZN(n1055) );
NAND2_X1 U770 ( .A1(G898), .A2(G224), .ZN(n1069) );
NOR2_X1 U771 ( .A1(n1070), .A2(n1071), .ZN(G66) );
XOR2_X1 U772 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U774 ( .A1(n1070), .A2(n1076), .ZN(G63) );
XOR2_X1 U775 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U776 ( .A(KEYINPUT35), .B(n1079), .Z(n1078) );
NOR2_X1 U777 ( .A1(n1080), .A2(n1075), .ZN(n1079) );
INV_X1 U778 ( .A(G478), .ZN(n1080) );
NOR2_X1 U779 ( .A1(n1070), .A2(n1081), .ZN(G60) );
NOR3_X1 U780 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NOR3_X1 U781 ( .A1(n1085), .A2(n1086), .A3(n1075), .ZN(n1084) );
NOR2_X1 U782 ( .A1(n1087), .A2(n1088), .ZN(n1083) );
INV_X1 U783 ( .A(n1085), .ZN(n1088) );
AND2_X1 U784 ( .A1(n966), .A2(G475), .ZN(n1087) );
XOR2_X1 U785 ( .A(n1089), .B(n1090), .Z(G6) );
NOR2_X1 U786 ( .A1(KEYINPUT15), .A2(n1091), .ZN(n1090) );
NOR4_X1 U787 ( .A1(n1092), .A2(n1093), .A3(n972), .A4(n1000), .ZN(n1089) );
NOR2_X1 U788 ( .A1(KEYINPUT49), .A2(n1094), .ZN(n1093) );
NOR2_X1 U789 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
AND2_X1 U790 ( .A1(n1097), .A2(KEYINPUT49), .ZN(n1092) );
NOR2_X1 U791 ( .A1(n1070), .A2(n1098), .ZN(G57) );
XOR2_X1 U792 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U793 ( .A(n1101), .B(G101), .Z(n1100) );
NAND2_X1 U794 ( .A1(n1102), .A2(KEYINPUT38), .ZN(n1099) );
XOR2_X1 U795 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U796 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U797 ( .A1(KEYINPUT19), .A2(n1107), .ZN(n1106) );
NOR2_X1 U798 ( .A1(n1108), .A2(n1075), .ZN(n1105) );
INV_X1 U799 ( .A(G472), .ZN(n1108) );
NOR2_X1 U800 ( .A1(n1070), .A2(n1109), .ZN(G54) );
XOR2_X1 U801 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U802 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U803 ( .A(KEYINPUT31), .B(G134), .Z(n1113) );
NOR2_X1 U804 ( .A1(n1114), .A2(n1075), .ZN(n1112) );
INV_X1 U805 ( .A(G469), .ZN(n1114) );
XNOR2_X1 U806 ( .A(n1115), .B(n1116), .ZN(n1110) );
XOR2_X1 U807 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND3_X1 U808 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1117) );
NAND2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
OR3_X1 U810 ( .A1(n1123), .A2(n1122), .A3(n1124), .ZN(n1120) );
NAND2_X1 U811 ( .A1(KEYINPUT6), .A2(n1044), .ZN(n1123) );
INV_X1 U812 ( .A(n1125), .ZN(n1044) );
NAND2_X1 U813 ( .A1(n1125), .A2(n1124), .ZN(n1119) );
INV_X1 U814 ( .A(KEYINPUT17), .ZN(n1124) );
XOR2_X1 U815 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U816 ( .A1(n1070), .A2(n1128), .ZN(G51) );
XOR2_X1 U817 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U818 ( .A(n1131), .B(n1132), .ZN(n1130) );
NOR2_X1 U819 ( .A1(KEYINPUT44), .A2(n1133), .ZN(n1131) );
XNOR2_X1 U820 ( .A(n1134), .B(KEYINPUT7), .ZN(n1133) );
NOR2_X1 U821 ( .A1(n1135), .A2(n1075), .ZN(n1129) );
NAND2_X1 U822 ( .A1(G902), .A2(n966), .ZN(n1075) );
NAND3_X1 U823 ( .A1(n1034), .A2(n1035), .A3(n1068), .ZN(n966) );
AND2_X1 U824 ( .A1(n1136), .A2(n1137), .ZN(n1068) );
NOR4_X1 U825 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1137) );
NOR4_X1 U826 ( .A1(n1142), .A2(n961), .A3(n1143), .A4(n1144), .ZN(n1136) );
NOR3_X1 U827 ( .A1(n1000), .A2(n972), .A3(n1097), .ZN(n1144) );
NOR3_X1 U828 ( .A1(n1001), .A2(n972), .A3(n1097), .ZN(n961) );
NAND3_X1 U829 ( .A1(n1145), .A2(n1007), .A3(n1146), .ZN(n1035) );
AND4_X1 U830 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1034) );
NOR4_X1 U831 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
INV_X1 U832 ( .A(n1155), .ZN(n1152) );
NAND3_X1 U833 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1149) );
XOR2_X1 U834 ( .A(KEYINPUT16), .B(n998), .Z(n1157) );
NOR2_X1 U835 ( .A1(n983), .A2(G952), .ZN(n1070) );
XNOR2_X1 U836 ( .A(G146), .B(n1159), .ZN(G48) );
NOR2_X1 U837 ( .A1(n1160), .A2(KEYINPUT43), .ZN(n1159) );
INV_X1 U838 ( .A(n1147), .ZN(n1160) );
NAND4_X1 U839 ( .A1(n1145), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1147) );
XNOR2_X1 U840 ( .A(G143), .B(n1164), .ZN(G45) );
NAND2_X1 U841 ( .A1(KEYINPUT45), .A2(n1165), .ZN(n1164) );
INV_X1 U842 ( .A(n1148), .ZN(n1165) );
NAND4_X1 U843 ( .A1(n1166), .A2(n1158), .A3(n995), .A4(n1020), .ZN(n1148) );
AND3_X1 U844 ( .A1(n979), .A2(n1163), .A3(n1006), .ZN(n1158) );
XNOR2_X1 U845 ( .A(G140), .B(n1167), .ZN(G42) );
NAND4_X1 U846 ( .A1(n998), .A2(n1145), .A3(n1168), .A4(n979), .ZN(n1167) );
NOR2_X1 U847 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U848 ( .A(n1163), .B(KEYINPUT20), .Z(n1170) );
XOR2_X1 U849 ( .A(G137), .B(n1153), .Z(G39) );
AND3_X1 U850 ( .A1(n981), .A2(n1162), .A3(n1146), .ZN(n1153) );
XNOR2_X1 U851 ( .A(G134), .B(n1171), .ZN(G36) );
NAND4_X1 U852 ( .A1(KEYINPUT21), .A2(n1146), .A3(n1006), .A4(n1156), .ZN(n1171) );
XOR2_X1 U853 ( .A(G131), .B(n1154), .Z(G33) );
AND3_X1 U854 ( .A1(n1145), .A2(n1006), .A3(n1146), .ZN(n1154) );
AND3_X1 U855 ( .A1(n979), .A2(n1163), .A3(n998), .ZN(n1146) );
NOR2_X1 U856 ( .A1(n1172), .A2(n997), .ZN(n998) );
XOR2_X1 U857 ( .A(n1126), .B(n1155), .Z(G30) );
NAND4_X1 U858 ( .A1(n1156), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1155) );
XOR2_X1 U859 ( .A(G101), .B(n1142), .Z(G3) );
NOR3_X1 U860 ( .A1(n1173), .A2(n1097), .A3(n974), .ZN(n1142) );
XOR2_X1 U861 ( .A(G125), .B(n1151), .Z(G27) );
AND4_X1 U862 ( .A1(n1007), .A2(n1163), .A3(n995), .A4(n1174), .ZN(n1151) );
NOR2_X1 U863 ( .A1(n1175), .A2(n1000), .ZN(n1174) );
NAND2_X1 U864 ( .A1(n987), .A2(n1176), .ZN(n1163) );
NAND4_X1 U865 ( .A1(G953), .A2(G902), .A3(n1177), .A4(n1043), .ZN(n1176) );
INV_X1 U866 ( .A(G900), .ZN(n1043) );
XOR2_X1 U867 ( .A(n1143), .B(n1178), .Z(G24) );
NOR2_X1 U868 ( .A1(KEYINPUT3), .A2(n1179), .ZN(n1178) );
AND4_X1 U869 ( .A1(n1166), .A2(n1180), .A3(n980), .A4(n1020), .ZN(n1143) );
INV_X1 U870 ( .A(n972), .ZN(n980) );
NAND2_X1 U871 ( .A1(n1181), .A2(n1182), .ZN(n972) );
XOR2_X1 U872 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U873 ( .A(n1141), .B(n1185), .Z(G21) );
XOR2_X1 U874 ( .A(KEYINPUT50), .B(G119), .Z(n1185) );
AND3_X1 U875 ( .A1(n981), .A2(n1162), .A3(n1180), .ZN(n1141) );
INV_X1 U876 ( .A(n974), .ZN(n981) );
XOR2_X1 U877 ( .A(G116), .B(n1140), .Z(G18) );
AND3_X1 U878 ( .A1(n1006), .A2(n1156), .A3(n1180), .ZN(n1140) );
INV_X1 U879 ( .A(n1001), .ZN(n1156) );
NAND2_X1 U880 ( .A1(n1020), .A2(n1186), .ZN(n1001) );
INV_X1 U881 ( .A(n1187), .ZN(n1020) );
XNOR2_X1 U882 ( .A(G113), .B(n1188), .ZN(G15) );
NAND2_X1 U883 ( .A1(KEYINPUT30), .A2(n1139), .ZN(n1188) );
AND3_X1 U884 ( .A1(n1145), .A2(n1006), .A3(n1180), .ZN(n1139) );
AND3_X1 U885 ( .A1(n995), .A2(n1096), .A3(n985), .ZN(n1180) );
INV_X1 U886 ( .A(n1175), .ZN(n985) );
NAND2_X1 U887 ( .A1(n977), .A2(n975), .ZN(n1175) );
INV_X1 U888 ( .A(n1000), .ZN(n1145) );
NAND2_X1 U889 ( .A1(n1166), .A2(n1187), .ZN(n1000) );
XOR2_X1 U890 ( .A(G110), .B(n1138), .Z(G12) );
NOR3_X1 U891 ( .A1(n1097), .A2(n1169), .A3(n974), .ZN(n1138) );
NAND2_X1 U892 ( .A1(n1187), .A2(n1186), .ZN(n974) );
INV_X1 U893 ( .A(n1166), .ZN(n1186) );
XOR2_X1 U894 ( .A(n1189), .B(n1082), .Z(n1166) );
INV_X1 U895 ( .A(n1024), .ZN(n1082) );
NAND2_X1 U896 ( .A1(n1085), .A2(n1190), .ZN(n1024) );
XOR2_X1 U897 ( .A(n1191), .B(n1192), .Z(n1085) );
XOR2_X1 U898 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U899 ( .A(G122), .B(G113), .Z(n1194) );
XOR2_X1 U900 ( .A(KEYINPUT34), .B(G131), .Z(n1193) );
XOR2_X1 U901 ( .A(n1195), .B(n1196), .Z(n1191) );
NOR2_X1 U902 ( .A1(KEYINPUT1), .A2(n1197), .ZN(n1196) );
XOR2_X1 U903 ( .A(n1091), .B(n1198), .Z(n1195) );
NOR2_X1 U904 ( .A1(KEYINPUT8), .A2(n1199), .ZN(n1198) );
XOR2_X1 U905 ( .A(G143), .B(n1200), .Z(n1199) );
AND3_X1 U906 ( .A1(n1201), .A2(n983), .A3(G214), .ZN(n1200) );
INV_X1 U907 ( .A(G104), .ZN(n1091) );
NAND2_X1 U908 ( .A1(KEYINPUT18), .A2(n1086), .ZN(n1189) );
INV_X1 U909 ( .A(G475), .ZN(n1086) );
XOR2_X1 U910 ( .A(n1202), .B(G478), .Z(n1187) );
OR2_X1 U911 ( .A1(n1077), .A2(G902), .ZN(n1202) );
XNOR2_X1 U912 ( .A(n1203), .B(n1204), .ZN(n1077) );
XOR2_X1 U913 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U914 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U915 ( .A1(G107), .A2(KEYINPUT14), .ZN(n1207) );
XOR2_X1 U916 ( .A(n1209), .B(n1210), .Z(n1203) );
XOR2_X1 U917 ( .A(KEYINPUT24), .B(G143), .Z(n1210) );
XOR2_X1 U918 ( .A(n1211), .B(G122), .Z(n1209) );
NAND2_X1 U919 ( .A1(G217), .A2(n1212), .ZN(n1211) );
INV_X1 U920 ( .A(n1007), .ZN(n1169) );
NAND2_X1 U921 ( .A1(n1213), .A2(n1214), .ZN(n1007) );
NAND2_X1 U922 ( .A1(n1162), .A2(n1183), .ZN(n1214) );
INV_X1 U923 ( .A(KEYINPUT0), .ZN(n1183) );
NAND2_X1 U924 ( .A1(n1215), .A2(n1216), .ZN(n1162) );
OR3_X1 U925 ( .A1(n1184), .A2(n1181), .A3(KEYINPUT13), .ZN(n1216) );
NAND2_X1 U926 ( .A1(KEYINPUT13), .A2(n1006), .ZN(n1215) );
INV_X1 U927 ( .A(n1173), .ZN(n1006) );
NAND2_X1 U928 ( .A1(n1181), .A2(n1019), .ZN(n1173) );
INV_X1 U929 ( .A(n1184), .ZN(n1019) );
NAND3_X1 U930 ( .A1(n1217), .A2(n1184), .A3(KEYINPUT0), .ZN(n1213) );
XOR2_X1 U931 ( .A(n1218), .B(G472), .Z(n1184) );
NAND2_X1 U932 ( .A1(n1219), .A2(n1190), .ZN(n1218) );
XOR2_X1 U933 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U934 ( .A(n1064), .B(n1107), .Z(n1221) );
XNOR2_X1 U935 ( .A(n1222), .B(n1223), .ZN(n1107) );
XNOR2_X1 U936 ( .A(n1101), .B(n1224), .ZN(n1220) );
NOR2_X1 U937 ( .A1(G101), .A2(KEYINPUT4), .ZN(n1224) );
NAND3_X1 U938 ( .A1(G210), .A2(n983), .A3(n1201), .ZN(n1101) );
XNOR2_X1 U939 ( .A(G237), .B(KEYINPUT12), .ZN(n1201) );
XNOR2_X1 U940 ( .A(KEYINPUT13), .B(n1181), .ZN(n1217) );
XNOR2_X1 U941 ( .A(n1018), .B(KEYINPUT33), .ZN(n1181) );
XOR2_X1 U942 ( .A(n1225), .B(n1074), .Z(n1018) );
NAND2_X1 U943 ( .A1(G217), .A2(n1226), .ZN(n1074) );
OR2_X1 U944 ( .A1(n1073), .A2(G902), .ZN(n1225) );
XNOR2_X1 U945 ( .A(n1227), .B(n1228), .ZN(n1073) );
XOR2_X1 U946 ( .A(G110), .B(n1229), .Z(n1228) );
XOR2_X1 U947 ( .A(G137), .B(G119), .Z(n1229) );
XNOR2_X1 U948 ( .A(n1197), .B(n1230), .ZN(n1227) );
XOR2_X1 U949 ( .A(n1231), .B(n1232), .Z(n1230) );
NAND2_X1 U950 ( .A1(KEYINPUT48), .A2(n1126), .ZN(n1232) );
NAND2_X1 U951 ( .A1(n1212), .A2(G221), .ZN(n1231) );
AND2_X1 U952 ( .A1(G234), .A2(n983), .ZN(n1212) );
XOR2_X1 U953 ( .A(G146), .B(n1054), .Z(n1197) );
XOR2_X1 U954 ( .A(G125), .B(G140), .Z(n1054) );
NAND2_X1 U955 ( .A1(n1161), .A2(n1096), .ZN(n1097) );
NAND2_X1 U956 ( .A1(n987), .A2(n1233), .ZN(n1096) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1177), .A4(n1234), .ZN(n1233) );
INV_X1 U958 ( .A(G898), .ZN(n1234) );
NAND3_X1 U959 ( .A1(n1177), .A2(n983), .A3(n1235), .ZN(n987) );
XNOR2_X1 U960 ( .A(G952), .B(KEYINPUT55), .ZN(n1235) );
NAND2_X1 U961 ( .A1(G237), .A2(G234), .ZN(n1177) );
INV_X1 U962 ( .A(n1095), .ZN(n1161) );
NAND2_X1 U963 ( .A1(n995), .A2(n979), .ZN(n1095) );
NOR2_X1 U964 ( .A1(n977), .A2(n1021), .ZN(n979) );
INV_X1 U965 ( .A(n975), .ZN(n1021) );
NAND2_X1 U966 ( .A1(n1236), .A2(G221), .ZN(n975) );
XOR2_X1 U967 ( .A(n1226), .B(KEYINPUT42), .Z(n1236) );
NAND2_X1 U968 ( .A1(G234), .A2(n1190), .ZN(n1226) );
XOR2_X1 U969 ( .A(n1017), .B(n1237), .Z(n977) );
NOR2_X1 U970 ( .A1(G469), .A2(KEYINPUT63), .ZN(n1237) );
AND2_X1 U971 ( .A1(n1238), .A2(n1190), .ZN(n1017) );
XOR2_X1 U972 ( .A(n1239), .B(n1240), .Z(n1238) );
XNOR2_X1 U973 ( .A(n1122), .B(n1115), .ZN(n1240) );
XNOR2_X1 U974 ( .A(n1241), .B(n1242), .ZN(n1115) );
XOR2_X1 U975 ( .A(G140), .B(G110), .Z(n1242) );
NAND2_X1 U976 ( .A1(G227), .A2(n983), .ZN(n1241) );
XNOR2_X1 U977 ( .A(n1243), .B(n1244), .ZN(n1122) );
NOR2_X1 U978 ( .A1(KEYINPUT41), .A2(n1245), .ZN(n1244) );
XOR2_X1 U979 ( .A(G107), .B(G104), .Z(n1245) );
XOR2_X1 U980 ( .A(n1222), .B(n1127), .Z(n1239) );
NOR2_X1 U981 ( .A1(KEYINPUT36), .A2(n1246), .ZN(n1127) );
XOR2_X1 U982 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U983 ( .A1(G146), .A2(KEYINPUT47), .ZN(n1247) );
XOR2_X1 U984 ( .A(n1118), .B(n1205), .Z(n1222) );
XOR2_X1 U985 ( .A(G128), .B(G134), .Z(n1205) );
XOR2_X1 U986 ( .A(n1052), .B(G137), .Z(n1118) );
INV_X1 U987 ( .A(G131), .ZN(n1052) );
NOR2_X1 U988 ( .A1(n997), .A2(n996), .ZN(n995) );
INV_X1 U989 ( .A(n1172), .ZN(n996) );
NAND2_X1 U990 ( .A1(n1249), .A2(n1023), .ZN(n1172) );
NAND2_X1 U991 ( .A1(n1250), .A2(n1251), .ZN(n1023) );
XOR2_X1 U992 ( .A(KEYINPUT5), .B(n1022), .Z(n1249) );
NOR2_X1 U993 ( .A1(n1251), .A2(n1250), .ZN(n1022) );
INV_X1 U994 ( .A(n1135), .ZN(n1250) );
NAND2_X1 U995 ( .A1(G210), .A2(n1252), .ZN(n1135) );
NAND2_X1 U996 ( .A1(n1253), .A2(n1190), .ZN(n1251) );
XOR2_X1 U997 ( .A(n1132), .B(n1134), .Z(n1253) );
XNOR2_X1 U998 ( .A(n1254), .B(n1255), .ZN(n1134) );
XOR2_X1 U999 ( .A(n1223), .B(n1256), .Z(n1255) );
AND2_X1 U1000 ( .A1(n983), .A2(G224), .ZN(n1256) );
INV_X1 U1001 ( .A(G953), .ZN(n983) );
NOR2_X1 U1002 ( .A1(KEYINPUT29), .A2(n1257), .ZN(n1223) );
XNOR2_X1 U1003 ( .A(G146), .B(n1248), .ZN(n1257) );
XOR2_X1 U1004 ( .A(G143), .B(KEYINPUT60), .Z(n1248) );
XOR2_X1 U1005 ( .A(G125), .B(n1126), .Z(n1254) );
INV_X1 U1006 ( .A(G128), .ZN(n1126) );
NAND2_X1 U1007 ( .A1(n1258), .A2(n1259), .ZN(n1132) );
NAND2_X1 U1008 ( .A1(n1260), .A2(n1066), .ZN(n1259) );
XOR2_X1 U1009 ( .A(n1261), .B(KEYINPUT37), .Z(n1258) );
OR2_X1 U1010 ( .A1(n1066), .A2(n1260), .ZN(n1261) );
XNOR2_X1 U1011 ( .A(n1065), .B(n1064), .ZN(n1260) );
INV_X1 U1012 ( .A(n1103), .ZN(n1064) );
XOR2_X1 U1013 ( .A(n1262), .B(n1208), .Z(n1103) );
XOR2_X1 U1014 ( .A(G116), .B(KEYINPUT22), .Z(n1208) );
XNOR2_X1 U1015 ( .A(G113), .B(G119), .ZN(n1262) );
XOR2_X1 U1016 ( .A(n1263), .B(n1264), .Z(n1065) );
XOR2_X1 U1017 ( .A(n1265), .B(n1266), .Z(n1264) );
INV_X1 U1018 ( .A(n1243), .ZN(n1266) );
XNOR2_X1 U1019 ( .A(G101), .B(KEYINPUT59), .ZN(n1243) );
NOR2_X1 U1020 ( .A1(G104), .A2(KEYINPUT25), .ZN(n1265) );
XNOR2_X1 U1021 ( .A(G107), .B(KEYINPUT58), .ZN(n1263) );
XNOR2_X1 U1022 ( .A(n1267), .B(G110), .ZN(n1066) );
NAND2_X1 U1023 ( .A1(KEYINPUT10), .A2(n1179), .ZN(n1267) );
INV_X1 U1024 ( .A(G122), .ZN(n1179) );
AND2_X1 U1025 ( .A1(G214), .A2(n1252), .ZN(n997) );
NAND2_X1 U1026 ( .A1(n1268), .A2(n1190), .ZN(n1252) );
INV_X1 U1027 ( .A(G902), .ZN(n1190) );
INV_X1 U1028 ( .A(G237), .ZN(n1268) );
endmodule


