//Key = 0110110100000110101010100110001000001100110001001110111011101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372;

XNOR2_X1 U758 ( .A(G107), .B(n1032), .ZN(G9) );
NAND2_X1 U759 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
XOR2_X1 U760 ( .A(n1035), .B(KEYINPUT54), .Z(n1033) );
NAND4_X1 U761 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
XNOR2_X1 U762 ( .A(n1040), .B(KEYINPUT5), .ZN(n1036) );
NOR2_X1 U763 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR3_X1 U764 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
NOR2_X1 U765 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR3_X1 U766 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1046) );
NAND3_X1 U767 ( .A1(n1051), .A2(n1038), .A3(n1037), .ZN(n1048) );
NAND3_X1 U768 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1043) );
NAND2_X1 U769 ( .A1(n1051), .A2(n1055), .ZN(n1054) );
NAND2_X1 U770 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND3_X1 U771 ( .A1(n1038), .A2(n1058), .A3(n1059), .ZN(n1057) );
NAND2_X1 U772 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U773 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U774 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U775 ( .A1(n1037), .A2(n1047), .ZN(n1065) );
INV_X1 U776 ( .A(KEYINPUT38), .ZN(n1047) );
INV_X1 U777 ( .A(n1066), .ZN(n1064) );
NAND2_X1 U778 ( .A1(n1067), .A2(n1068), .ZN(n1060) );
NAND2_X1 U779 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U780 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U781 ( .A1(n1062), .A2(n1073), .A3(n1067), .ZN(n1056) );
NAND3_X1 U782 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NAND2_X1 U783 ( .A1(n1077), .A2(n1059), .ZN(n1076) );
INV_X1 U784 ( .A(n1078), .ZN(n1075) );
NAND2_X1 U785 ( .A1(n1038), .A2(n1079), .ZN(n1074) );
NAND2_X1 U786 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U787 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U788 ( .A1(n1084), .A2(G953), .A3(G952), .ZN(n1041) );
INV_X1 U789 ( .A(n1052), .ZN(n1084) );
NAND4_X1 U790 ( .A1(n1085), .A2(n1062), .A3(n1086), .A4(n1087), .ZN(n1052) );
NOR4_X1 U791 ( .A1(n1088), .A2(n1089), .A3(n1049), .A4(n1090), .ZN(n1087) );
NOR2_X1 U792 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
XOR2_X1 U793 ( .A(n1093), .B(G475), .Z(n1086) );
XNOR2_X1 U794 ( .A(n1094), .B(n1095), .ZN(n1085) );
XOR2_X1 U795 ( .A(n1096), .B(n1097), .Z(G72) );
XOR2_X1 U796 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR3_X1 U797 ( .A1(n1100), .A2(KEYINPUT11), .A3(n1101), .ZN(n1099) );
XOR2_X1 U798 ( .A(n1102), .B(n1103), .Z(n1100) );
NAND2_X1 U799 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U801 ( .A(n1108), .B(n1109), .ZN(n1107) );
XNOR2_X1 U802 ( .A(n1110), .B(KEYINPUT18), .ZN(n1106) );
NAND2_X1 U803 ( .A1(n1111), .A2(n1112), .ZN(n1104) );
XNOR2_X1 U804 ( .A(n1108), .B(n1113), .ZN(n1112) );
INV_X1 U805 ( .A(n1109), .ZN(n1113) );
NAND2_X1 U806 ( .A1(n1114), .A2(n1115), .ZN(n1108) );
NAND2_X1 U807 ( .A1(G137), .A2(n1116), .ZN(n1115) );
XOR2_X1 U808 ( .A(KEYINPUT36), .B(n1117), .Z(n1114) );
NOR2_X1 U809 ( .A1(G137), .A2(n1116), .ZN(n1117) );
XNOR2_X1 U810 ( .A(n1110), .B(KEYINPUT28), .ZN(n1111) );
NAND2_X1 U811 ( .A1(n1118), .A2(n1119), .ZN(n1098) );
XNOR2_X1 U812 ( .A(G953), .B(KEYINPUT31), .ZN(n1118) );
NAND2_X1 U813 ( .A1(G953), .A2(n1120), .ZN(n1096) );
NAND2_X1 U814 ( .A1(G900), .A2(G227), .ZN(n1120) );
XOR2_X1 U815 ( .A(n1121), .B(n1122), .Z(G69) );
NOR2_X1 U816 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U817 ( .A(KEYINPUT12), .B(n1125), .Z(n1124) );
NOR3_X1 U818 ( .A1(n1126), .A2(G953), .A3(n1127), .ZN(n1125) );
INV_X1 U819 ( .A(n1128), .ZN(n1127) );
NOR3_X1 U820 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1123) );
NOR2_X1 U821 ( .A1(G953), .A2(n1126), .ZN(n1130) );
AND2_X1 U822 ( .A1(n1131), .A2(n1132), .ZN(n1126) );
NOR2_X1 U823 ( .A1(G898), .A2(n1053), .ZN(n1129) );
NAND2_X1 U824 ( .A1(n1133), .A2(n1134), .ZN(n1128) );
OR2_X1 U825 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U826 ( .A(n1137), .B(KEYINPUT29), .Z(n1133) );
NAND2_X1 U827 ( .A1(n1136), .A2(n1135), .ZN(n1137) );
NAND2_X1 U828 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
NAND2_X1 U829 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U830 ( .A(KEYINPUT45), .B(n1142), .Z(n1138) );
NOR2_X1 U831 ( .A1(n1140), .A2(n1141), .ZN(n1142) );
XNOR2_X1 U832 ( .A(KEYINPUT53), .B(n1143), .ZN(n1141) );
NAND3_X1 U833 ( .A1(G953), .A2(n1144), .A3(KEYINPUT25), .ZN(n1121) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1144) );
NOR2_X1 U835 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XNOR2_X1 U836 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U837 ( .A(n1149), .B(KEYINPUT7), .Z(n1148) );
NAND2_X1 U838 ( .A1(n1150), .A2(n1091), .ZN(n1149) );
INV_X1 U839 ( .A(n1151), .ZN(n1091) );
NOR2_X1 U840 ( .A1(n1145), .A2(n1152), .ZN(G63) );
XNOR2_X1 U841 ( .A(n1153), .B(n1154), .ZN(n1152) );
NAND2_X1 U842 ( .A1(n1150), .A2(G478), .ZN(n1153) );
NOR2_X1 U843 ( .A1(n1145), .A2(n1155), .ZN(G60) );
XOR2_X1 U844 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U845 ( .A1(n1158), .A2(KEYINPUT59), .ZN(n1157) );
AND2_X1 U846 ( .A1(G475), .A2(n1150), .ZN(n1158) );
XNOR2_X1 U847 ( .A(G104), .B(n1159), .ZN(G6) );
NOR2_X1 U848 ( .A1(n1145), .A2(n1160), .ZN(G57) );
XOR2_X1 U849 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U850 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U851 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
INV_X1 U852 ( .A(n1167), .ZN(n1166) );
XNOR2_X1 U853 ( .A(n1168), .B(n1169), .ZN(n1165) );
XNOR2_X1 U854 ( .A(KEYINPUT62), .B(KEYINPUT58), .ZN(n1169) );
NOR2_X1 U855 ( .A1(n1168), .A2(n1167), .ZN(n1163) );
XNOR2_X1 U856 ( .A(n1170), .B(n1171), .ZN(n1167) );
NAND2_X1 U857 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
OR2_X1 U858 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U859 ( .A(n1176), .B(KEYINPUT33), .Z(n1172) );
NAND2_X1 U860 ( .A1(n1175), .A2(n1174), .ZN(n1176) );
NOR2_X1 U861 ( .A1(n1177), .A2(n1095), .ZN(n1168) );
NAND3_X1 U862 ( .A1(n1178), .A2(n1179), .A3(KEYINPUT56), .ZN(n1161) );
OR3_X1 U863 ( .A1(n1180), .A2(G101), .A3(KEYINPUT48), .ZN(n1179) );
NAND2_X1 U864 ( .A1(n1181), .A2(KEYINPUT48), .ZN(n1178) );
XNOR2_X1 U865 ( .A(G101), .B(n1182), .ZN(n1181) );
NAND2_X1 U866 ( .A1(KEYINPUT52), .A2(n1180), .ZN(n1182) );
NOR2_X1 U867 ( .A1(n1145), .A2(n1183), .ZN(G54) );
XOR2_X1 U868 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND2_X1 U869 ( .A1(n1150), .A2(G469), .ZN(n1185) );
NAND2_X1 U870 ( .A1(n1186), .A2(n1187), .ZN(n1184) );
NAND2_X1 U871 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U872 ( .A(n1190), .B(KEYINPUT47), .Z(n1186) );
OR2_X1 U873 ( .A1(n1189), .A2(n1188), .ZN(n1190) );
XOR2_X1 U874 ( .A(n1191), .B(n1192), .Z(n1188) );
NOR2_X1 U875 ( .A1(KEYINPUT39), .A2(G110), .ZN(n1192) );
XNOR2_X1 U876 ( .A(G140), .B(n1193), .ZN(n1191) );
NAND2_X1 U877 ( .A1(n1194), .A2(n1195), .ZN(n1189) );
NOR2_X1 U878 ( .A1(n1145), .A2(n1196), .ZN(G51) );
XNOR2_X1 U879 ( .A(n1197), .B(n1198), .ZN(n1196) );
XOR2_X1 U880 ( .A(n1199), .B(KEYINPUT35), .Z(n1198) );
NAND2_X1 U881 ( .A1(n1150), .A2(G210), .ZN(n1199) );
INV_X1 U882 ( .A(n1177), .ZN(n1150) );
NAND2_X1 U883 ( .A1(G902), .A2(n1045), .ZN(n1177) );
NAND3_X1 U884 ( .A1(n1200), .A2(n1201), .A3(n1131), .ZN(n1045) );
AND4_X1 U885 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1131) );
XOR2_X1 U886 ( .A(KEYINPUT0), .B(n1132), .Z(n1201) );
AND4_X1 U887 ( .A1(n1159), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1132) );
NAND3_X1 U888 ( .A1(n1209), .A2(n1038), .A3(n1210), .ZN(n1206) );
XNOR2_X1 U889 ( .A(KEYINPUT4), .B(n1039), .ZN(n1209) );
NAND3_X1 U890 ( .A1(n1066), .A2(n1038), .A3(n1211), .ZN(n1159) );
INV_X1 U891 ( .A(n1119), .ZN(n1200) );
NAND4_X1 U892 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1119) );
AND4_X1 U893 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1215) );
NAND2_X1 U894 ( .A1(n1034), .A2(n1220), .ZN(n1214) );
NAND2_X1 U895 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND3_X1 U896 ( .A1(n1223), .A2(n1037), .A3(n1224), .ZN(n1222) );
XOR2_X1 U897 ( .A(n1225), .B(KEYINPUT51), .Z(n1221) );
NAND3_X1 U898 ( .A1(n1226), .A2(n1077), .A3(n1227), .ZN(n1212) );
XNOR2_X1 U899 ( .A(n1059), .B(KEYINPUT1), .ZN(n1227) );
NOR2_X1 U900 ( .A1(n1053), .A2(G952), .ZN(n1145) );
XOR2_X1 U901 ( .A(n1228), .B(n1229), .Z(G48) );
NOR2_X1 U902 ( .A1(KEYINPUT15), .A2(n1230), .ZN(n1229) );
INV_X1 U903 ( .A(G146), .ZN(n1230) );
NOR2_X1 U904 ( .A1(n1080), .A2(n1225), .ZN(n1228) );
NAND2_X1 U905 ( .A1(n1226), .A2(n1223), .ZN(n1225) );
XNOR2_X1 U906 ( .A(G143), .B(n1213), .ZN(G45) );
NAND3_X1 U907 ( .A1(n1224), .A2(n1034), .A3(n1231), .ZN(n1213) );
NOR3_X1 U908 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
XNOR2_X1 U909 ( .A(G140), .B(n1235), .ZN(G42) );
NAND4_X1 U910 ( .A1(KEYINPUT60), .A2(n1226), .A3(n1077), .A4(n1059), .ZN(n1235) );
XNOR2_X1 U911 ( .A(G137), .B(n1219), .ZN(G39) );
NAND4_X1 U912 ( .A1(n1224), .A2(n1067), .A3(n1223), .A4(n1059), .ZN(n1219) );
INV_X1 U913 ( .A(n1049), .ZN(n1059) );
XNOR2_X1 U914 ( .A(G134), .B(n1218), .ZN(G36) );
NAND3_X1 U915 ( .A1(n1224), .A2(n1037), .A3(n1078), .ZN(n1218) );
XNOR2_X1 U916 ( .A(G131), .B(n1236), .ZN(G33) );
NAND2_X1 U917 ( .A1(KEYINPUT57), .A2(n1237), .ZN(n1236) );
INV_X1 U918 ( .A(n1217), .ZN(n1237) );
NAND2_X1 U919 ( .A1(n1078), .A2(n1226), .ZN(n1217) );
AND2_X1 U920 ( .A1(n1224), .A2(n1066), .ZN(n1226) );
AND2_X1 U921 ( .A1(n1040), .A2(n1238), .ZN(n1224) );
NOR2_X1 U922 ( .A1(n1049), .A2(n1232), .ZN(n1078) );
NAND2_X1 U923 ( .A1(n1083), .A2(n1239), .ZN(n1049) );
INV_X1 U924 ( .A(n1082), .ZN(n1239) );
XNOR2_X1 U925 ( .A(G128), .B(n1240), .ZN(G30) );
NAND3_X1 U926 ( .A1(n1223), .A2(n1241), .A3(n1210), .ZN(n1240) );
AND3_X1 U927 ( .A1(n1037), .A2(n1040), .A3(n1034), .ZN(n1210) );
XNOR2_X1 U928 ( .A(KEYINPUT13), .B(n1238), .ZN(n1241) );
XNOR2_X1 U929 ( .A(G101), .B(n1207), .ZN(G3) );
NAND3_X1 U930 ( .A1(n1067), .A2(n1242), .A3(n1211), .ZN(n1207) );
XNOR2_X1 U931 ( .A(G125), .B(n1216), .ZN(G27) );
NAND4_X1 U932 ( .A1(n1034), .A2(n1238), .A3(n1062), .A4(n1243), .ZN(n1216) );
AND2_X1 U933 ( .A1(n1066), .A2(n1077), .ZN(n1243) );
INV_X1 U934 ( .A(n1050), .ZN(n1062) );
NAND2_X1 U935 ( .A1(n1244), .A2(n1245), .ZN(n1238) );
NAND3_X1 U936 ( .A1(G902), .A2(n1246), .A3(n1101), .ZN(n1245) );
NOR2_X1 U937 ( .A1(n1053), .A2(G900), .ZN(n1101) );
XOR2_X1 U938 ( .A(G122), .B(n1247), .Z(G24) );
NOR2_X1 U939 ( .A1(KEYINPUT21), .A2(n1202), .ZN(n1247) );
NAND4_X1 U940 ( .A1(n1248), .A2(n1249), .A3(n1038), .A4(n1250), .ZN(n1202) );
NAND2_X1 U941 ( .A1(n1251), .A2(n1252), .ZN(n1038) );
OR2_X1 U942 ( .A1(n1232), .A2(KEYINPUT22), .ZN(n1252) );
NAND3_X1 U943 ( .A1(n1253), .A2(n1254), .A3(KEYINPUT22), .ZN(n1251) );
XNOR2_X1 U944 ( .A(G119), .B(n1203), .ZN(G21) );
NAND3_X1 U945 ( .A1(n1223), .A2(n1249), .A3(n1067), .ZN(n1203) );
NOR2_X1 U946 ( .A1(n1254), .A2(n1253), .ZN(n1223) );
INV_X1 U947 ( .A(n1255), .ZN(n1254) );
XNOR2_X1 U948 ( .A(G116), .B(n1204), .ZN(G18) );
NAND3_X1 U949 ( .A1(n1037), .A2(n1242), .A3(n1249), .ZN(n1204) );
NOR2_X1 U950 ( .A1(n1250), .A2(n1234), .ZN(n1037) );
XNOR2_X1 U951 ( .A(G113), .B(n1205), .ZN(G15) );
NAND3_X1 U952 ( .A1(n1249), .A2(n1242), .A3(n1066), .ZN(n1205) );
NOR2_X1 U953 ( .A1(n1248), .A2(n1233), .ZN(n1066) );
INV_X1 U954 ( .A(n1250), .ZN(n1233) );
INV_X1 U955 ( .A(n1232), .ZN(n1242) );
NAND2_X1 U956 ( .A1(n1253), .A2(n1255), .ZN(n1232) );
NOR3_X1 U957 ( .A1(n1080), .A2(n1256), .A3(n1050), .ZN(n1249) );
NAND2_X1 U958 ( .A1(n1072), .A2(n1257), .ZN(n1050) );
XNOR2_X1 U959 ( .A(G110), .B(n1208), .ZN(G12) );
NAND3_X1 U960 ( .A1(n1077), .A2(n1067), .A3(n1211), .ZN(n1208) );
NOR3_X1 U961 ( .A1(n1069), .A2(n1256), .A3(n1080), .ZN(n1211) );
INV_X1 U962 ( .A(n1034), .ZN(n1080) );
NOR2_X1 U963 ( .A1(n1083), .A2(n1082), .ZN(n1034) );
NOR2_X1 U964 ( .A1(n1258), .A2(n1259), .ZN(n1082) );
XOR2_X1 U965 ( .A(n1260), .B(n1261), .Z(n1083) );
NOR2_X1 U966 ( .A1(n1259), .A2(n1262), .ZN(n1261) );
XOR2_X1 U967 ( .A(KEYINPUT2), .B(G210), .Z(n1262) );
NOR2_X1 U968 ( .A1(G902), .A2(G237), .ZN(n1259) );
NAND2_X1 U969 ( .A1(n1263), .A2(n1264), .ZN(n1260) );
XNOR2_X1 U970 ( .A(KEYINPUT37), .B(n1265), .ZN(n1263) );
INV_X1 U971 ( .A(n1197), .ZN(n1265) );
XNOR2_X1 U972 ( .A(n1266), .B(n1267), .ZN(n1197) );
XNOR2_X1 U973 ( .A(n1268), .B(n1110), .ZN(n1267) );
NAND2_X1 U974 ( .A1(G224), .A2(n1053), .ZN(n1268) );
XOR2_X1 U975 ( .A(n1269), .B(G125), .Z(n1266) );
NAND3_X1 U976 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1269) );
OR2_X1 U977 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U978 ( .A1(KEYINPUT44), .A2(n1275), .ZN(n1271) );
NAND2_X1 U979 ( .A1(n1276), .A2(n1274), .ZN(n1275) );
XNOR2_X1 U980 ( .A(n1273), .B(KEYINPUT26), .ZN(n1276) );
NAND2_X1 U981 ( .A1(n1277), .A2(n1278), .ZN(n1270) );
INV_X1 U982 ( .A(KEYINPUT44), .ZN(n1278) );
NAND2_X1 U983 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
OR2_X1 U984 ( .A1(n1273), .A2(KEYINPUT26), .ZN(n1280) );
NAND3_X1 U985 ( .A1(n1273), .A2(n1274), .A3(KEYINPUT26), .ZN(n1279) );
INV_X1 U986 ( .A(n1136), .ZN(n1274) );
XOR2_X1 U987 ( .A(G110), .B(n1281), .Z(n1136) );
XNOR2_X1 U988 ( .A(n1143), .B(n1282), .ZN(n1273) );
NOR2_X1 U989 ( .A1(KEYINPUT32), .A2(n1140), .ZN(n1282) );
XNOR2_X1 U990 ( .A(G101), .B(n1283), .ZN(n1140) );
NOR2_X1 U991 ( .A1(KEYINPUT34), .A2(n1284), .ZN(n1283) );
NAND2_X1 U992 ( .A1(n1285), .A2(n1286), .ZN(n1143) );
NAND2_X1 U993 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U994 ( .A(KEYINPUT20), .B(n1289), .Z(n1285) );
NOR2_X1 U995 ( .A1(n1287), .A2(n1288), .ZN(n1289) );
XOR2_X1 U996 ( .A(KEYINPUT23), .B(n1290), .Z(n1287) );
INV_X1 U997 ( .A(n1039), .ZN(n1256) );
NAND2_X1 U998 ( .A1(n1291), .A2(n1292), .ZN(n1039) );
NAND4_X1 U999 ( .A1(G953), .A2(G902), .A3(n1246), .A4(n1293), .ZN(n1292) );
INV_X1 U1000 ( .A(G898), .ZN(n1293) );
XNOR2_X1 U1001 ( .A(n1051), .B(KEYINPUT42), .ZN(n1291) );
INV_X1 U1002 ( .A(n1244), .ZN(n1051) );
NAND3_X1 U1003 ( .A1(n1246), .A2(n1053), .A3(G952), .ZN(n1244) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1246) );
INV_X1 U1005 ( .A(n1040), .ZN(n1069) );
NOR2_X1 U1006 ( .A1(n1072), .A2(n1071), .ZN(n1040) );
INV_X1 U1007 ( .A(n1257), .ZN(n1071) );
NAND2_X1 U1008 ( .A1(G221), .A2(n1294), .ZN(n1257) );
XOR2_X1 U1009 ( .A(n1295), .B(G469), .Z(n1072) );
NAND2_X1 U1010 ( .A1(n1296), .A2(n1264), .ZN(n1295) );
XOR2_X1 U1011 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U1012 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1013 ( .A(n1301), .B(KEYINPUT30), .Z(n1300) );
NAND2_X1 U1014 ( .A1(G110), .A2(n1302), .ZN(n1301) );
NOR2_X1 U1015 ( .A1(G110), .A2(n1302), .ZN(n1299) );
XOR2_X1 U1016 ( .A(n1303), .B(n1193), .Z(n1297) );
AND2_X1 U1017 ( .A1(G227), .A2(n1053), .ZN(n1193) );
NAND3_X1 U1018 ( .A1(n1304), .A2(n1305), .A3(n1195), .ZN(n1303) );
NAND2_X1 U1019 ( .A1(n1306), .A2(n1307), .ZN(n1195) );
NAND2_X1 U1020 ( .A1(KEYINPUT43), .A2(n1308), .ZN(n1305) );
NAND3_X1 U1021 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1308) );
INV_X1 U1022 ( .A(n1306), .ZN(n1311) );
NOR2_X1 U1023 ( .A1(n1312), .A2(n1110), .ZN(n1306) );
NAND2_X1 U1024 ( .A1(n1313), .A2(n1307), .ZN(n1310) );
INV_X1 U1025 ( .A(n1314), .ZN(n1307) );
NAND3_X1 U1026 ( .A1(n1314), .A2(n1110), .A3(n1312), .ZN(n1309) );
OR2_X1 U1027 ( .A1(n1194), .A2(KEYINPUT43), .ZN(n1304) );
AND2_X1 U1028 ( .A1(n1315), .A2(n1316), .ZN(n1194) );
NAND3_X1 U1029 ( .A1(n1314), .A2(n1312), .A3(n1175), .ZN(n1316) );
NAND2_X1 U1030 ( .A1(n1317), .A2(n1110), .ZN(n1315) );
INV_X1 U1031 ( .A(n1175), .ZN(n1110) );
XNOR2_X1 U1032 ( .A(n1314), .B(n1313), .ZN(n1317) );
INV_X1 U1033 ( .A(n1312), .ZN(n1313) );
XOR2_X1 U1034 ( .A(n1174), .B(KEYINPUT14), .Z(n1312) );
XOR2_X1 U1035 ( .A(n1318), .B(n1284), .Z(n1314) );
XNOR2_X1 U1036 ( .A(G104), .B(G107), .ZN(n1284) );
XNOR2_X1 U1037 ( .A(G101), .B(KEYINPUT19), .ZN(n1318) );
NOR2_X1 U1038 ( .A1(n1250), .A2(n1248), .ZN(n1067) );
INV_X1 U1039 ( .A(n1234), .ZN(n1248) );
XOR2_X1 U1040 ( .A(n1090), .B(KEYINPUT63), .Z(n1234) );
XOR2_X1 U1041 ( .A(G478), .B(n1319), .Z(n1090) );
NOR2_X1 U1042 ( .A1(G902), .A2(n1154), .ZN(n1319) );
XNOR2_X1 U1043 ( .A(n1320), .B(n1321), .ZN(n1154) );
XOR2_X1 U1044 ( .A(n1281), .B(n1322), .Z(n1321) );
XOR2_X1 U1045 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR2_X1 U1046 ( .A1(G134), .A2(KEYINPUT10), .ZN(n1324) );
AND3_X1 U1047 ( .A1(G234), .A2(n1053), .A3(G217), .ZN(n1323) );
XOR2_X1 U1048 ( .A(n1325), .B(n1326), .Z(n1320) );
XNOR2_X1 U1049 ( .A(n1327), .B(G128), .ZN(n1326) );
INV_X1 U1050 ( .A(G143), .ZN(n1327) );
XNOR2_X1 U1051 ( .A(G107), .B(G116), .ZN(n1325) );
XOR2_X1 U1052 ( .A(n1328), .B(n1093), .Z(n1250) );
NAND2_X1 U1053 ( .A1(n1156), .A2(n1264), .ZN(n1093) );
XOR2_X1 U1054 ( .A(n1329), .B(n1330), .Z(n1156) );
XNOR2_X1 U1055 ( .A(n1281), .B(n1331), .ZN(n1330) );
XNOR2_X1 U1056 ( .A(n1332), .B(n1333), .ZN(n1331) );
NOR2_X1 U1057 ( .A1(KEYINPUT6), .A2(n1103), .ZN(n1333) );
XOR2_X1 U1058 ( .A(G122), .B(KEYINPUT24), .Z(n1281) );
XOR2_X1 U1059 ( .A(n1334), .B(n1335), .Z(n1329) );
XOR2_X1 U1060 ( .A(G104), .B(n1336), .Z(n1335) );
NOR3_X1 U1061 ( .A1(n1258), .A2(G953), .A3(G237), .ZN(n1336) );
INV_X1 U1062 ( .A(G214), .ZN(n1258) );
XNOR2_X1 U1063 ( .A(G131), .B(G113), .ZN(n1334) );
NAND2_X1 U1064 ( .A1(KEYINPUT41), .A2(G475), .ZN(n1328) );
NOR2_X1 U1065 ( .A1(n1255), .A2(n1253), .ZN(n1077) );
NOR2_X1 U1066 ( .A1(n1337), .A2(n1088), .ZN(n1253) );
NOR2_X1 U1067 ( .A1(n1151), .A2(n1338), .ZN(n1088) );
AND2_X1 U1068 ( .A1(n1339), .A2(n1151), .ZN(n1337) );
NAND2_X1 U1069 ( .A1(G217), .A2(n1294), .ZN(n1151) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1264), .ZN(n1294) );
XNOR2_X1 U1071 ( .A(KEYINPUT27), .B(n1092), .ZN(n1339) );
INV_X1 U1072 ( .A(n1338), .ZN(n1092) );
NOR2_X1 U1073 ( .A1(n1340), .A2(G902), .ZN(n1338) );
INV_X1 U1074 ( .A(n1147), .ZN(n1340) );
XNOR2_X1 U1075 ( .A(n1341), .B(n1342), .ZN(n1147) );
XOR2_X1 U1076 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1077 ( .A(G119), .B(n1345), .Z(n1344) );
AND3_X1 U1078 ( .A1(G221), .A2(n1053), .A3(G234), .ZN(n1345) );
INV_X1 U1079 ( .A(G953), .ZN(n1053) );
XNOR2_X1 U1080 ( .A(n1346), .B(G128), .ZN(n1343) );
INV_X1 U1081 ( .A(G137), .ZN(n1346) );
XOR2_X1 U1082 ( .A(n1347), .B(n1103), .Z(n1341) );
XNOR2_X1 U1083 ( .A(G125), .B(n1302), .ZN(n1103) );
INV_X1 U1084 ( .A(G140), .ZN(n1302) );
XNOR2_X1 U1085 ( .A(n1348), .B(n1349), .ZN(n1347) );
NOR2_X1 U1086 ( .A1(G110), .A2(KEYINPUT9), .ZN(n1349) );
NOR2_X1 U1087 ( .A1(G146), .A2(KEYINPUT3), .ZN(n1348) );
NAND3_X1 U1088 ( .A1(n1350), .A2(n1351), .A3(n1352), .ZN(n1255) );
NAND2_X1 U1089 ( .A1(G472), .A2(n1094), .ZN(n1352) );
NAND2_X1 U1090 ( .A1(n1353), .A2(n1354), .ZN(n1351) );
INV_X1 U1091 ( .A(KEYINPUT16), .ZN(n1354) );
NAND2_X1 U1092 ( .A1(n1355), .A2(n1095), .ZN(n1353) );
INV_X1 U1093 ( .A(G472), .ZN(n1095) );
XNOR2_X1 U1094 ( .A(n1094), .B(n1356), .ZN(n1355) );
NAND2_X1 U1095 ( .A1(KEYINPUT16), .A2(n1357), .ZN(n1350) );
NAND2_X1 U1096 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
NAND2_X1 U1097 ( .A1(n1094), .A2(n1356), .ZN(n1359) );
OR3_X1 U1098 ( .A1(n1094), .A2(G472), .A3(n1356), .ZN(n1358) );
INV_X1 U1099 ( .A(KEYINPUT50), .ZN(n1356) );
NAND2_X1 U1100 ( .A1(n1360), .A2(n1264), .ZN(n1094) );
INV_X1 U1101 ( .A(G902), .ZN(n1264) );
XOR2_X1 U1102 ( .A(n1361), .B(n1362), .Z(n1360) );
XNOR2_X1 U1103 ( .A(n1363), .B(n1171), .ZN(n1362) );
XOR2_X1 U1104 ( .A(n1364), .B(n1288), .Z(n1171) );
INV_X1 U1105 ( .A(G113), .ZN(n1288) );
NAND2_X1 U1106 ( .A1(KEYINPUT61), .A2(n1290), .ZN(n1364) );
XNOR2_X1 U1107 ( .A(G116), .B(G119), .ZN(n1290) );
NAND2_X1 U1108 ( .A1(KEYINPUT40), .A2(n1365), .ZN(n1363) );
INV_X1 U1109 ( .A(G101), .ZN(n1365) );
XOR2_X1 U1110 ( .A(n1366), .B(n1180), .Z(n1361) );
NOR3_X1 U1111 ( .A1(G237), .A2(G953), .A3(n1367), .ZN(n1180) );
INV_X1 U1112 ( .A(G210), .ZN(n1367) );
NAND2_X1 U1113 ( .A1(KEYINPUT49), .A2(n1368), .ZN(n1366) );
XNOR2_X1 U1114 ( .A(n1175), .B(n1174), .ZN(n1368) );
XOR2_X1 U1115 ( .A(n1109), .B(n1369), .Z(n1174) );
NOR2_X1 U1116 ( .A1(KEYINPUT8), .A2(n1370), .ZN(n1369) );
XNOR2_X1 U1117 ( .A(G137), .B(n1371), .ZN(n1370) );
NOR2_X1 U1118 ( .A1(KEYINPUT55), .A2(n1372), .ZN(n1371) );
XNOR2_X1 U1119 ( .A(KEYINPUT46), .B(n1116), .ZN(n1372) );
INV_X1 U1120 ( .A(G134), .ZN(n1116) );
XOR2_X1 U1121 ( .A(G131), .B(KEYINPUT17), .Z(n1109) );
XNOR2_X1 U1122 ( .A(G128), .B(n1332), .ZN(n1175) );
XOR2_X1 U1123 ( .A(G143), .B(G146), .Z(n1332) );
endmodule


