//Key = 1111000010001010101000111001110001001111000001000101100011010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369;

XNOR2_X1 U760 ( .A(n1043), .B(n1044), .ZN(G9) );
NOR2_X1 U761 ( .A1(n1045), .A2(n1046), .ZN(G75) );
XOR2_X1 U762 ( .A(KEYINPUT55), .B(n1047), .Z(n1046) );
AND3_X1 U763 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NOR4_X1 U764 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1049), .ZN(n1045) );
INV_X1 U765 ( .A(G952), .ZN(n1049) );
XOR2_X1 U766 ( .A(n1054), .B(KEYINPUT25), .Z(n1053) );
NAND2_X1 U767 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND3_X1 U768 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1056) );
NAND2_X1 U769 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U770 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U771 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND3_X1 U772 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NAND2_X1 U773 ( .A1(n1069), .A2(n1070), .ZN(n1060) );
NAND2_X1 U774 ( .A1(n1071), .A2(n1072), .ZN(n1055) );
INV_X1 U775 ( .A(n1073), .ZN(n1052) );
NAND4_X1 U776 ( .A1(n1048), .A2(n1074), .A3(n1075), .A4(n1050), .ZN(n1051) );
NAND4_X1 U777 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1050) );
NOR3_X1 U778 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NAND3_X1 U779 ( .A1(n1067), .A2(n1083), .A3(n1084), .ZN(n1080) );
NOR3_X1 U780 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1078) );
AND3_X1 U781 ( .A1(KEYINPUT39), .A2(n1088), .A3(G478), .ZN(n1087) );
NOR2_X1 U782 ( .A1(KEYINPUT39), .A2(G478), .ZN(n1086) );
XOR2_X1 U783 ( .A(n1089), .B(n1090), .Z(n1085) );
XNOR2_X1 U784 ( .A(n1091), .B(n1092), .ZN(n1077) );
XNOR2_X1 U785 ( .A(n1066), .B(KEYINPUT20), .ZN(n1076) );
NAND3_X1 U786 ( .A1(n1057), .A2(n1093), .A3(n1059), .ZN(n1075) );
NAND2_X1 U787 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND4_X1 U788 ( .A1(n1096), .A2(n1069), .A3(n1097), .A4(n1098), .ZN(n1095) );
INV_X1 U789 ( .A(KEYINPUT9), .ZN(n1098) );
INV_X1 U790 ( .A(n1084), .ZN(n1096) );
NAND2_X1 U791 ( .A1(n1062), .A2(n1099), .ZN(n1094) );
NAND2_X1 U792 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND3_X1 U793 ( .A1(n1102), .A2(n1068), .A3(n1103), .ZN(n1101) );
INV_X1 U794 ( .A(n1066), .ZN(n1102) );
NAND2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1100) );
NAND2_X1 U796 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U797 ( .A1(KEYINPUT9), .A2(n1068), .ZN(n1107) );
INV_X1 U798 ( .A(n1108), .ZN(n1106) );
NAND2_X1 U799 ( .A1(n1071), .A2(n1109), .ZN(n1074) );
AND3_X1 U800 ( .A1(n1069), .A2(n1062), .A3(n1059), .ZN(n1071) );
INV_X1 U801 ( .A(n1110), .ZN(n1059) );
XOR2_X1 U802 ( .A(n1111), .B(n1112), .Z(G72) );
NOR2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR2_X1 U805 ( .A1(KEYINPUT19), .A2(n1117), .ZN(n1111) );
XOR2_X1 U806 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U809 ( .A1(G900), .A2(n1114), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1114), .A2(n1124), .ZN(n1118) );
NAND2_X1 U811 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
INV_X1 U813 ( .A(n1129), .ZN(n1128) );
NAND2_X1 U814 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
NAND3_X1 U815 ( .A1(n1132), .A2(n1114), .A3(KEYINPUT18), .ZN(n1131) );
NAND3_X1 U816 ( .A1(n1133), .A2(n1134), .A3(n1129), .ZN(n1125) );
NOR3_X1 U817 ( .A1(KEYINPUT7), .A2(n1135), .A3(n1136), .ZN(n1129) );
XOR2_X1 U818 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR3_X1 U819 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NOR2_X1 U820 ( .A1(KEYINPUT47), .A2(n1142), .ZN(n1141) );
NOR2_X1 U821 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR3_X1 U822 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
NOR2_X1 U823 ( .A1(KEYINPUT37), .A2(n1148), .ZN(n1143) );
NOR2_X1 U824 ( .A1(n1149), .A2(n1150), .ZN(n1140) );
INV_X1 U825 ( .A(KEYINPUT47), .ZN(n1150) );
NOR2_X1 U826 ( .A1(n1146), .A2(n1151), .ZN(n1149) );
XNOR2_X1 U827 ( .A(n1145), .B(n1148), .ZN(n1151) );
INV_X1 U828 ( .A(KEYINPUT37), .ZN(n1145) );
AND2_X1 U829 ( .A1(n1146), .A2(n1147), .ZN(n1139) );
INV_X1 U830 ( .A(n1148), .ZN(n1147) );
XOR2_X1 U831 ( .A(G113), .B(n1152), .Z(n1148) );
XOR2_X1 U832 ( .A(G104), .B(n1153), .Z(n1146) );
NOR2_X1 U833 ( .A1(KEYINPUT48), .A2(n1154), .ZN(n1137) );
XNOR2_X1 U834 ( .A(G122), .B(G110), .ZN(n1154) );
NAND2_X1 U835 ( .A1(n1132), .A2(n1114), .ZN(n1134) );
XNOR2_X1 U836 ( .A(n1130), .B(KEYINPUT18), .ZN(n1133) );
NOR2_X1 U837 ( .A1(n1135), .A2(n1155), .ZN(n1130) );
NOR2_X1 U838 ( .A1(n1114), .A2(G224), .ZN(n1155) );
NOR2_X1 U839 ( .A1(n1156), .A2(n1157), .ZN(G66) );
NOR3_X1 U840 ( .A1(n1089), .A2(n1158), .A3(n1159), .ZN(n1157) );
AND3_X1 U841 ( .A1(n1160), .A2(G217), .A3(n1161), .ZN(n1159) );
NOR2_X1 U842 ( .A1(n1162), .A2(n1160), .ZN(n1158) );
NOR2_X1 U843 ( .A1(n1073), .A2(n1163), .ZN(n1162) );
NOR2_X1 U844 ( .A1(n1156), .A2(n1164), .ZN(G63) );
XOR2_X1 U845 ( .A(n1165), .B(n1166), .Z(n1164) );
AND2_X1 U846 ( .A1(G478), .A2(n1161), .ZN(n1166) );
NAND2_X1 U847 ( .A1(n1167), .A2(KEYINPUT14), .ZN(n1165) );
XOR2_X1 U848 ( .A(n1168), .B(KEYINPUT10), .Z(n1167) );
NOR2_X1 U849 ( .A1(n1156), .A2(n1169), .ZN(G60) );
XOR2_X1 U850 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR4_X1 U851 ( .A1(n1073), .A2(n1172), .A3(n1173), .A4(n1092), .ZN(n1170) );
INV_X1 U852 ( .A(G475), .ZN(n1092) );
XNOR2_X1 U853 ( .A(KEYINPUT41), .B(KEYINPUT3), .ZN(n1173) );
XNOR2_X1 U854 ( .A(G902), .B(KEYINPUT46), .ZN(n1172) );
XOR2_X1 U855 ( .A(G104), .B(n1174), .Z(G6) );
NOR2_X1 U856 ( .A1(n1156), .A2(n1175), .ZN(G57) );
XOR2_X1 U857 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U858 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U859 ( .A(n1180), .B(n1181), .Z(n1176) );
XOR2_X1 U860 ( .A(n1182), .B(KEYINPUT52), .Z(n1181) );
NAND3_X1 U861 ( .A1(n1183), .A2(n1184), .A3(KEYINPUT33), .ZN(n1182) );
NAND2_X1 U862 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
INV_X1 U863 ( .A(KEYINPUT23), .ZN(n1186) );
NAND2_X1 U864 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NAND3_X1 U865 ( .A1(KEYINPUT6), .A2(n1189), .A3(n1190), .ZN(n1188) );
NAND2_X1 U866 ( .A1(n1191), .A2(n1192), .ZN(n1187) );
NAND2_X1 U867 ( .A1(n1193), .A2(KEYINPUT23), .ZN(n1183) );
XNOR2_X1 U868 ( .A(n1190), .B(n1191), .ZN(n1193) );
NOR2_X1 U869 ( .A1(n1194), .A2(KEYINPUT6), .ZN(n1191) );
NAND2_X1 U870 ( .A1(n1161), .A2(G472), .ZN(n1180) );
NOR2_X1 U871 ( .A1(n1156), .A2(n1195), .ZN(G54) );
XOR2_X1 U872 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U873 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U874 ( .A(KEYINPUT26), .B(G146), .Z(n1199) );
NOR2_X1 U875 ( .A1(KEYINPUT40), .A2(n1200), .ZN(n1198) );
XOR2_X1 U876 ( .A(n1201), .B(n1202), .Z(n1200) );
XNOR2_X1 U877 ( .A(n1203), .B(G110), .ZN(n1202) );
XOR2_X1 U878 ( .A(n1204), .B(n1122), .Z(n1196) );
XOR2_X1 U879 ( .A(n1205), .B(n1206), .Z(n1122) );
XOR2_X1 U880 ( .A(n1207), .B(n1208), .Z(n1204) );
NAND2_X1 U881 ( .A1(n1161), .A2(G469), .ZN(n1207) );
NOR2_X1 U882 ( .A1(n1156), .A2(n1209), .ZN(G51) );
XOR2_X1 U883 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U884 ( .A(n1212), .B(KEYINPUT13), .Z(n1210) );
NAND2_X1 U885 ( .A1(n1161), .A2(n1213), .ZN(n1212) );
NOR2_X1 U886 ( .A1(n1214), .A2(n1073), .ZN(n1161) );
NOR2_X1 U887 ( .A1(n1124), .A2(n1132), .ZN(n1073) );
NAND4_X1 U888 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1132) );
AND4_X1 U889 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1218) );
NOR2_X1 U890 ( .A1(n1174), .A2(n1044), .ZN(n1217) );
AND3_X1 U891 ( .A1(n1109), .A2(n1068), .A3(n1223), .ZN(n1044) );
AND3_X1 U892 ( .A1(n1223), .A2(n1068), .A3(n1072), .ZN(n1174) );
NAND2_X1 U893 ( .A1(n1070), .A2(n1224), .ZN(n1216) );
NAND2_X1 U894 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND4_X1 U895 ( .A1(n1227), .A2(n1228), .A3(n1072), .A4(n1229), .ZN(n1226) );
INV_X1 U896 ( .A(n1230), .ZN(n1227) );
XNOR2_X1 U897 ( .A(n1231), .B(KEYINPUT35), .ZN(n1225) );
OR2_X1 U898 ( .A1(n1229), .A2(n1232), .ZN(n1215) );
INV_X1 U899 ( .A(KEYINPUT59), .ZN(n1229) );
NAND4_X1 U900 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1124) );
NOR4_X1 U901 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
NOR2_X1 U902 ( .A1(KEYINPUT34), .A2(n1241), .ZN(n1240) );
NOR2_X1 U903 ( .A1(KEYINPUT44), .A2(n1242), .ZN(n1239) );
NOR2_X1 U904 ( .A1(n1243), .A2(n1244), .ZN(n1238) );
NOR2_X1 U905 ( .A1(n1245), .A2(n1246), .ZN(n1243) );
AND4_X1 U906 ( .A1(n1247), .A2(n1072), .A3(n1108), .A4(KEYINPUT34), .ZN(n1246) );
NOR3_X1 U907 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1245) );
INV_X1 U908 ( .A(KEYINPUT44), .ZN(n1249) );
NAND3_X1 U909 ( .A1(n1251), .A2(n1252), .A3(n1070), .ZN(n1248) );
AND3_X1 U910 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1235) );
NOR2_X1 U911 ( .A1(n1114), .A2(G952), .ZN(n1156) );
XNOR2_X1 U912 ( .A(G146), .B(n1255), .ZN(G48) );
NAND4_X1 U913 ( .A1(n1072), .A2(n1256), .A3(n1257), .A4(n1070), .ZN(n1255) );
XOR2_X1 U914 ( .A(n1242), .B(n1258), .Z(G45) );
XNOR2_X1 U915 ( .A(G143), .B(KEYINPUT5), .ZN(n1258) );
NAND4_X1 U916 ( .A1(n1259), .A2(n1260), .A3(n1070), .A4(n1251), .ZN(n1242) );
NAND2_X1 U917 ( .A1(n1261), .A2(n1262), .ZN(G42) );
NAND2_X1 U918 ( .A1(n1263), .A2(n1203), .ZN(n1262) );
XOR2_X1 U919 ( .A(KEYINPUT28), .B(n1264), .Z(n1261) );
NOR2_X1 U920 ( .A1(n1263), .A2(n1203), .ZN(n1264) );
INV_X1 U921 ( .A(n1241), .ZN(n1263) );
NAND4_X1 U922 ( .A1(n1108), .A2(n1072), .A3(n1062), .A4(n1257), .ZN(n1241) );
XOR2_X1 U923 ( .A(n1254), .B(n1265), .Z(G39) );
NAND2_X1 U924 ( .A1(G137), .A2(n1266), .ZN(n1265) );
XOR2_X1 U925 ( .A(KEYINPUT50), .B(KEYINPUT12), .Z(n1266) );
NAND4_X1 U926 ( .A1(n1057), .A2(n1256), .A3(n1062), .A4(n1257), .ZN(n1254) );
XOR2_X1 U927 ( .A(G134), .B(n1237), .Z(G36) );
AND3_X1 U928 ( .A1(n1062), .A2(n1109), .A3(n1260), .ZN(n1237) );
XOR2_X1 U929 ( .A(n1233), .B(n1267), .Z(G33) );
NAND2_X1 U930 ( .A1(KEYINPUT27), .A2(G131), .ZN(n1267) );
NAND3_X1 U931 ( .A1(n1072), .A2(n1062), .A3(n1260), .ZN(n1233) );
NOR2_X1 U932 ( .A1(n1252), .A2(n1244), .ZN(n1260) );
INV_X1 U933 ( .A(n1247), .ZN(n1062) );
NAND2_X1 U934 ( .A1(n1097), .A2(n1084), .ZN(n1247) );
XOR2_X1 U935 ( .A(n1082), .B(KEYINPUT49), .Z(n1097) );
XNOR2_X1 U936 ( .A(G128), .B(n1234), .ZN(G30) );
NAND4_X1 U937 ( .A1(n1256), .A2(n1257), .A3(n1109), .A4(n1070), .ZN(n1234) );
INV_X1 U938 ( .A(n1244), .ZN(n1257) );
NAND3_X1 U939 ( .A1(n1268), .A2(n1067), .A3(n1066), .ZN(n1244) );
XNOR2_X1 U940 ( .A(G101), .B(n1222), .ZN(G3) );
NAND3_X1 U941 ( .A1(n1057), .A2(n1223), .A3(n1269), .ZN(n1222) );
XNOR2_X1 U942 ( .A(G125), .B(n1253), .ZN(G27) );
NAND3_X1 U943 ( .A1(n1270), .A2(n1268), .A3(n1108), .ZN(n1253) );
NAND2_X1 U944 ( .A1(n1110), .A2(n1271), .ZN(n1268) );
NAND4_X1 U945 ( .A1(G902), .A2(G953), .A3(n1272), .A4(n1116), .ZN(n1271) );
INV_X1 U946 ( .A(G900), .ZN(n1116) );
XNOR2_X1 U947 ( .A(G122), .B(n1221), .ZN(G24) );
NAND4_X1 U948 ( .A1(n1259), .A2(n1069), .A3(n1273), .A4(n1251), .ZN(n1221) );
AND2_X1 U949 ( .A1(n1104), .A2(n1068), .ZN(n1069) );
NOR2_X1 U950 ( .A1(n1081), .A2(n1274), .ZN(n1068) );
XNOR2_X1 U951 ( .A(n1275), .B(n1276), .ZN(G21) );
NAND2_X1 U952 ( .A1(KEYINPUT0), .A2(n1277), .ZN(n1275) );
NAND2_X1 U953 ( .A1(n1231), .A2(n1070), .ZN(n1277) );
AND4_X1 U954 ( .A1(n1104), .A2(n1057), .A3(n1256), .A4(n1230), .ZN(n1231) );
AND2_X1 U955 ( .A1(n1274), .A2(n1081), .ZN(n1256) );
INV_X1 U956 ( .A(n1278), .ZN(n1274) );
XOR2_X1 U957 ( .A(n1220), .B(n1279), .Z(G18) );
NAND2_X1 U958 ( .A1(KEYINPUT51), .A2(G116), .ZN(n1279) );
NAND3_X1 U959 ( .A1(n1109), .A2(n1273), .A3(n1228), .ZN(n1220) );
INV_X1 U960 ( .A(n1064), .ZN(n1228) );
NAND2_X1 U961 ( .A1(n1269), .A2(n1104), .ZN(n1064) );
AND2_X1 U962 ( .A1(n1250), .A2(n1251), .ZN(n1109) );
XNOR2_X1 U963 ( .A(G113), .B(n1232), .ZN(G15) );
NAND3_X1 U964 ( .A1(n1270), .A2(n1230), .A3(n1269), .ZN(n1232) );
INV_X1 U965 ( .A(n1252), .ZN(n1269) );
NAND2_X1 U966 ( .A1(n1278), .A2(n1081), .ZN(n1252) );
AND3_X1 U967 ( .A1(n1072), .A2(n1070), .A3(n1104), .ZN(n1270) );
NOR2_X1 U968 ( .A1(n1066), .A2(n1103), .ZN(n1104) );
INV_X1 U969 ( .A(n1067), .ZN(n1103) );
NOR2_X1 U970 ( .A1(n1250), .A2(n1251), .ZN(n1072) );
XNOR2_X1 U971 ( .A(G110), .B(n1280), .ZN(G12) );
NAND2_X1 U972 ( .A1(KEYINPUT56), .A2(n1281), .ZN(n1280) );
INV_X1 U973 ( .A(n1219), .ZN(n1281) );
NAND3_X1 U974 ( .A1(n1057), .A2(n1223), .A3(n1108), .ZN(n1219) );
NOR2_X1 U975 ( .A1(n1278), .A2(n1081), .ZN(n1108) );
XNOR2_X1 U976 ( .A(n1282), .B(G472), .ZN(n1081) );
NAND2_X1 U977 ( .A1(n1283), .A2(n1214), .ZN(n1282) );
XOR2_X1 U978 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U979 ( .A(n1286), .B(n1189), .ZN(n1285) );
NOR2_X1 U980 ( .A1(KEYINPUT4), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U981 ( .A(n1288), .B(n1178), .ZN(n1287) );
XOR2_X1 U982 ( .A(n1289), .B(n1290), .Z(n1178) );
NAND2_X1 U983 ( .A1(KEYINPUT2), .A2(n1179), .ZN(n1288) );
XNOR2_X1 U984 ( .A(G113), .B(n1291), .ZN(n1179) );
XNOR2_X1 U985 ( .A(n1192), .B(KEYINPUT17), .ZN(n1284) );
INV_X1 U986 ( .A(n1190), .ZN(n1192) );
NAND3_X1 U987 ( .A1(n1292), .A2(n1114), .A3(G210), .ZN(n1190) );
XNOR2_X1 U988 ( .A(n1293), .B(n1090), .ZN(n1278) );
AND2_X1 U989 ( .A1(n1294), .A2(G217), .ZN(n1090) );
XOR2_X1 U990 ( .A(n1295), .B(KEYINPUT15), .Z(n1294) );
XNOR2_X1 U991 ( .A(KEYINPUT31), .B(n1296), .ZN(n1293) );
NOR2_X1 U992 ( .A1(n1089), .A2(KEYINPUT54), .ZN(n1296) );
NOR2_X1 U993 ( .A1(n1160), .A2(G902), .ZN(n1089) );
XOR2_X1 U994 ( .A(n1123), .B(n1297), .Z(n1160) );
XOR2_X1 U995 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR3_X1 U996 ( .A1(n1300), .A2(KEYINPUT53), .A3(n1301), .ZN(n1299) );
NOR2_X1 U997 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XOR2_X1 U998 ( .A(n1304), .B(KEYINPUT1), .Z(n1300) );
NAND2_X1 U999 ( .A1(n1302), .A2(n1303), .ZN(n1304) );
XNOR2_X1 U1000 ( .A(G119), .B(G128), .ZN(n1302) );
NOR2_X1 U1001 ( .A1(n1305), .A2(n1306), .ZN(n1298) );
XOR2_X1 U1002 ( .A(KEYINPUT30), .B(n1307), .Z(n1306) );
NOR3_X1 U1003 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1307) );
NOR2_X1 U1004 ( .A1(n1311), .A2(G137), .ZN(n1305) );
NOR2_X1 U1005 ( .A1(n1309), .A2(n1308), .ZN(n1311) );
INV_X1 U1006 ( .A(G221), .ZN(n1309) );
AND3_X1 U1007 ( .A1(n1066), .A2(n1067), .A3(n1273), .ZN(n1223) );
AND2_X1 U1008 ( .A1(n1070), .A2(n1230), .ZN(n1273) );
NAND2_X1 U1009 ( .A1(n1110), .A2(n1312), .ZN(n1230) );
NAND3_X1 U1010 ( .A1(n1135), .A2(n1272), .A3(G902), .ZN(n1312) );
NOR2_X1 U1011 ( .A1(G898), .A2(n1114), .ZN(n1135) );
NAND3_X1 U1012 ( .A1(n1048), .A2(n1272), .A3(G952), .ZN(n1110) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1272) );
XOR2_X1 U1014 ( .A(G953), .B(KEYINPUT22), .Z(n1048) );
AND2_X1 U1015 ( .A1(n1082), .A2(n1084), .ZN(n1070) );
NAND2_X1 U1016 ( .A1(G214), .A2(n1313), .ZN(n1084) );
XNOR2_X1 U1017 ( .A(n1314), .B(n1213), .ZN(n1082) );
AND2_X1 U1018 ( .A1(G210), .A2(n1313), .ZN(n1213) );
NAND2_X1 U1019 ( .A1(n1292), .A2(n1214), .ZN(n1313) );
NAND2_X1 U1020 ( .A1(n1211), .A2(n1214), .ZN(n1314) );
XNOR2_X1 U1021 ( .A(n1315), .B(n1316), .ZN(n1211) );
XOR2_X1 U1022 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1023 ( .A(n1319), .B(n1152), .Z(n1318) );
NOR2_X1 U1024 ( .A1(KEYINPUT42), .A2(n1291), .ZN(n1152) );
XOR2_X1 U1025 ( .A(G116), .B(n1276), .Z(n1291) );
INV_X1 U1026 ( .A(G119), .ZN(n1276) );
NAND2_X1 U1027 ( .A1(G224), .A2(n1114), .ZN(n1319) );
XNOR2_X1 U1028 ( .A(G125), .B(G110), .ZN(n1317) );
XOR2_X1 U1029 ( .A(n1289), .B(n1320), .Z(n1315) );
XOR2_X1 U1030 ( .A(n1321), .B(n1153), .Z(n1320) );
NAND2_X1 U1031 ( .A1(n1322), .A2(n1323), .ZN(n1289) );
NAND2_X1 U1032 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
XOR2_X1 U1033 ( .A(n1326), .B(KEYINPUT58), .Z(n1324) );
NAND2_X1 U1034 ( .A1(G128), .A2(n1327), .ZN(n1322) );
XOR2_X1 U1035 ( .A(n1326), .B(KEYINPUT8), .Z(n1327) );
XNOR2_X1 U1036 ( .A(G143), .B(n1328), .ZN(n1326) );
NOR2_X1 U1037 ( .A1(G146), .A2(KEYINPUT61), .ZN(n1328) );
NAND2_X1 U1038 ( .A1(G221), .A2(n1295), .ZN(n1067) );
NAND2_X1 U1039 ( .A1(G234), .A2(n1214), .ZN(n1295) );
XNOR2_X1 U1040 ( .A(n1329), .B(G469), .ZN(n1066) );
NAND2_X1 U1041 ( .A1(n1330), .A2(n1214), .ZN(n1329) );
XOR2_X1 U1042 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U1043 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1044 ( .A(n1335), .B(n1290), .ZN(n1334) );
INV_X1 U1045 ( .A(n1205), .ZN(n1290) );
XOR2_X1 U1046 ( .A(G131), .B(n1336), .Z(n1205) );
XNOR2_X1 U1047 ( .A(n1310), .B(G134), .ZN(n1336) );
INV_X1 U1048 ( .A(G137), .ZN(n1310) );
NAND2_X1 U1049 ( .A1(KEYINPUT16), .A2(n1201), .ZN(n1335) );
NOR2_X1 U1050 ( .A1(n1115), .A2(G953), .ZN(n1201) );
INV_X1 U1051 ( .A(G227), .ZN(n1115) );
NAND2_X1 U1052 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
NAND2_X1 U1053 ( .A1(KEYINPUT43), .A2(n1303), .ZN(n1338) );
INV_X1 U1054 ( .A(G110), .ZN(n1303) );
NAND2_X1 U1055 ( .A1(KEYINPUT36), .A2(G110), .ZN(n1337) );
XOR2_X1 U1056 ( .A(n1339), .B(n1340), .Z(n1331) );
XOR2_X1 U1057 ( .A(KEYINPUT29), .B(KEYINPUT26), .Z(n1340) );
XNOR2_X1 U1058 ( .A(n1341), .B(n1203), .ZN(n1339) );
NAND2_X1 U1059 ( .A1(n1342), .A2(KEYINPUT45), .ZN(n1341) );
XNOR2_X1 U1060 ( .A(n1206), .B(n1343), .ZN(n1342) );
XOR2_X1 U1061 ( .A(G146), .B(n1344), .Z(n1343) );
NOR2_X1 U1062 ( .A1(KEYINPUT60), .A2(n1208), .ZN(n1344) );
XOR2_X1 U1063 ( .A(n1153), .B(n1345), .Z(n1208) );
NOR2_X1 U1064 ( .A1(G104), .A2(KEYINPUT63), .ZN(n1345) );
XNOR2_X1 U1065 ( .A(G107), .B(n1189), .ZN(n1153) );
INV_X1 U1066 ( .A(n1194), .ZN(n1189) );
XOR2_X1 U1067 ( .A(G101), .B(KEYINPUT38), .Z(n1194) );
XOR2_X1 U1068 ( .A(G143), .B(n1346), .Z(n1206) );
NOR2_X1 U1069 ( .A1(G128), .A2(KEYINPUT32), .ZN(n1346) );
NOR2_X1 U1070 ( .A1(n1251), .A2(n1259), .ZN(n1057) );
INV_X1 U1071 ( .A(n1250), .ZN(n1259) );
XNOR2_X1 U1072 ( .A(n1091), .B(n1347), .ZN(n1250) );
NOR2_X1 U1073 ( .A1(G475), .A2(KEYINPUT62), .ZN(n1347) );
OR2_X1 U1074 ( .A1(n1171), .A2(G902), .ZN(n1091) );
XNOR2_X1 U1075 ( .A(n1348), .B(n1349), .ZN(n1171) );
XNOR2_X1 U1076 ( .A(n1350), .B(n1321), .ZN(n1349) );
XOR2_X1 U1077 ( .A(G104), .B(n1351), .Z(n1321) );
XOR2_X1 U1078 ( .A(G122), .B(G113), .Z(n1351) );
NAND2_X1 U1079 ( .A1(KEYINPUT57), .A2(n1123), .ZN(n1350) );
XNOR2_X1 U1080 ( .A(G125), .B(n1352), .ZN(n1123) );
XNOR2_X1 U1081 ( .A(G146), .B(n1203), .ZN(n1352) );
INV_X1 U1082 ( .A(G140), .ZN(n1203) );
XOR2_X1 U1083 ( .A(n1353), .B(n1354), .Z(n1348) );
XOR2_X1 U1084 ( .A(G143), .B(G131), .Z(n1354) );
NAND3_X1 U1085 ( .A1(n1292), .A2(n1114), .A3(G214), .ZN(n1353) );
INV_X1 U1086 ( .A(G237), .ZN(n1292) );
NAND2_X1 U1087 ( .A1(n1083), .A2(n1355), .ZN(n1251) );
NAND2_X1 U1088 ( .A1(G478), .A2(n1088), .ZN(n1355) );
OR2_X1 U1089 ( .A1(n1088), .A2(G478), .ZN(n1083) );
NAND2_X1 U1090 ( .A1(n1168), .A2(n1214), .ZN(n1088) );
INV_X1 U1091 ( .A(G902), .ZN(n1214) );
XOR2_X1 U1092 ( .A(n1356), .B(n1357), .Z(n1168) );
NOR2_X1 U1093 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
XOR2_X1 U1094 ( .A(KEYINPUT11), .B(n1360), .Z(n1359) );
NOR2_X1 U1095 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
AND2_X1 U1096 ( .A1(n1362), .A2(n1361), .ZN(n1358) );
XOR2_X1 U1097 ( .A(n1325), .B(n1363), .Z(n1361) );
XOR2_X1 U1098 ( .A(G143), .B(G134), .Z(n1363) );
INV_X1 U1099 ( .A(G128), .ZN(n1325) );
NAND3_X1 U1100 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1362) );
OR2_X1 U1101 ( .A1(n1043), .A2(n1367), .ZN(n1366) );
NAND3_X1 U1102 ( .A1(n1367), .A2(n1043), .A3(KEYINPUT24), .ZN(n1365) );
INV_X1 U1103 ( .A(G107), .ZN(n1043) );
NOR2_X1 U1104 ( .A1(KEYINPUT21), .A2(n1368), .ZN(n1367) );
NAND2_X1 U1105 ( .A1(n1368), .A2(n1369), .ZN(n1364) );
INV_X1 U1106 ( .A(KEYINPUT24), .ZN(n1369) );
XNOR2_X1 U1107 ( .A(G116), .B(G122), .ZN(n1368) );
OR2_X1 U1108 ( .A1(n1163), .A2(n1308), .ZN(n1356) );
NAND2_X1 U1109 ( .A1(G234), .A2(n1114), .ZN(n1308) );
INV_X1 U1110 ( .A(G953), .ZN(n1114) );
INV_X1 U1111 ( .A(G217), .ZN(n1163) );
endmodule


