//Key = 0011001001111111101101001011101001101000110100100001101000110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404;

XNOR2_X1 U761 ( .A(G107), .B(n1049), .ZN(G9) );
NOR2_X1 U762 ( .A1(n1050), .A2(n1051), .ZN(G75) );
XOR2_X1 U763 ( .A(n1052), .B(KEYINPUT58), .Z(n1051) );
NAND4_X1 U764 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NAND2_X1 U765 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND4_X1 U767 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
NAND2_X1 U768 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
OR2_X1 U769 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1059) );
NAND2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U772 ( .A1(n1061), .A2(n1073), .A3(n1074), .ZN(n1072) );
XNOR2_X1 U773 ( .A(n1062), .B(KEYINPUT54), .ZN(n1074) );
NAND2_X1 U774 ( .A1(n1063), .A2(n1075), .ZN(n1071) );
NAND2_X1 U775 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U776 ( .A1(n1061), .A2(n1078), .ZN(n1077) );
NAND2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U778 ( .A1(KEYINPUT12), .A2(n1081), .ZN(n1080) );
NAND2_X1 U779 ( .A1(n1062), .A2(n1082), .ZN(n1076) );
NAND2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U781 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U782 ( .A1(n1061), .A2(n1087), .ZN(n1055) );
NAND2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND4_X1 U784 ( .A1(n1069), .A2(n1081), .A3(n1090), .A4(n1063), .ZN(n1089) );
NOR2_X1 U785 ( .A1(KEYINPUT12), .A2(n1057), .ZN(n1090) );
INV_X1 U786 ( .A(n1091), .ZN(n1057) );
XOR2_X1 U787 ( .A(n1092), .B(KEYINPUT23), .Z(n1088) );
NAND4_X1 U788 ( .A1(n1093), .A2(n1094), .A3(n1069), .A4(n1095), .ZN(n1092) );
NOR2_X1 U789 ( .A1(n1096), .A2(n1091), .ZN(n1095) );
INV_X1 U790 ( .A(n1097), .ZN(n1054) );
NOR2_X1 U791 ( .A1(G952), .A2(n1097), .ZN(n1050) );
NAND2_X1 U792 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND4_X1 U793 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
NOR4_X1 U794 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1103) );
AND2_X1 U795 ( .A1(n1108), .A2(KEYINPUT61), .ZN(n1107) );
NOR3_X1 U796 ( .A1(KEYINPUT61), .A2(n1109), .A3(n1108), .ZN(n1106) );
XNOR2_X1 U797 ( .A(KEYINPUT4), .B(n1110), .ZN(n1105) );
NAND4_X1 U798 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1104) );
NAND3_X1 U799 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
OR2_X1 U800 ( .A1(n1117), .A2(n1115), .ZN(n1113) );
INV_X1 U801 ( .A(KEYINPUT39), .ZN(n1117) );
NAND3_X1 U802 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1112) );
INV_X1 U803 ( .A(KEYINPUT25), .ZN(n1120) );
NAND2_X1 U804 ( .A1(KEYINPUT25), .A2(n1121), .ZN(n1111) );
NOR3_X1 U805 ( .A1(n1122), .A2(n1123), .A3(n1085), .ZN(n1102) );
NOR2_X1 U806 ( .A1(G902), .A2(n1124), .ZN(n1122) );
NOR4_X1 U807 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1124) );
NOR2_X1 U808 ( .A1(G469), .A2(n1129), .ZN(n1128) );
AND2_X1 U809 ( .A1(n1121), .A2(n1130), .ZN(n1127) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1115), .ZN(n1126) );
XNOR2_X1 U811 ( .A(n1132), .B(KEYINPUT63), .ZN(n1115) );
NOR2_X1 U812 ( .A1(n1133), .A2(n1134), .ZN(n1125) );
XNOR2_X1 U813 ( .A(G475), .B(KEYINPUT27), .ZN(n1133) );
XNOR2_X1 U814 ( .A(n1135), .B(n1136), .ZN(n1100) );
XOR2_X1 U815 ( .A(n1137), .B(n1138), .Z(G72) );
XOR2_X1 U816 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U817 ( .A1(n1141), .A2(n1098), .ZN(n1140) );
AND2_X1 U818 ( .A1(G227), .A2(G900), .ZN(n1141) );
NAND2_X1 U819 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
NAND2_X1 U820 ( .A1(G953), .A2(n1144), .ZN(n1143) );
XOR2_X1 U821 ( .A(n1145), .B(n1146), .Z(n1142) );
XNOR2_X1 U822 ( .A(n1147), .B(n1148), .ZN(n1146) );
NAND2_X1 U823 ( .A1(KEYINPUT3), .A2(n1149), .ZN(n1147) );
XOR2_X1 U824 ( .A(n1150), .B(n1151), .Z(n1145) );
XNOR2_X1 U825 ( .A(G125), .B(KEYINPUT59), .ZN(n1151) );
NAND3_X1 U826 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1150) );
NAND2_X1 U827 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND3_X1 U828 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1155) );
NAND2_X1 U829 ( .A1(KEYINPUT24), .A2(KEYINPUT50), .ZN(n1159) );
NAND2_X1 U830 ( .A1(G137), .A2(n1160), .ZN(n1158) );
NAND2_X1 U831 ( .A1(n1161), .A2(n1162), .ZN(n1157) );
NAND2_X1 U832 ( .A1(n1160), .A2(n1163), .ZN(n1161) );
NAND2_X1 U833 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
INV_X1 U834 ( .A(KEYINPUT1), .ZN(n1160) );
NAND4_X1 U835 ( .A1(G134), .A2(n1162), .A3(KEYINPUT24), .A4(n1165), .ZN(n1153) );
INV_X1 U836 ( .A(KEYINPUT50), .ZN(n1165) );
NAND2_X1 U837 ( .A1(KEYINPUT50), .A2(n1166), .ZN(n1152) );
NAND2_X1 U838 ( .A1(n1162), .A2(n1167), .ZN(n1166) );
NAND2_X1 U839 ( .A1(G134), .A2(n1164), .ZN(n1167) );
INV_X1 U840 ( .A(KEYINPUT24), .ZN(n1164) );
NAND2_X1 U841 ( .A1(n1098), .A2(n1168), .ZN(n1137) );
XOR2_X1 U842 ( .A(n1169), .B(n1170), .Z(G69) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U844 ( .A1(n1173), .A2(n1098), .ZN(n1172) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NAND2_X1 U846 ( .A1(n1176), .A2(n1177), .ZN(n1171) );
NAND2_X1 U847 ( .A1(G953), .A2(n1175), .ZN(n1177) );
XOR2_X1 U848 ( .A(n1178), .B(KEYINPUT13), .Z(n1176) );
NAND2_X1 U849 ( .A1(n1098), .A2(n1179), .ZN(n1169) );
NOR2_X1 U850 ( .A1(n1180), .A2(n1181), .ZN(G66) );
XNOR2_X1 U851 ( .A(n1182), .B(n1131), .ZN(n1181) );
NAND2_X1 U852 ( .A1(n1183), .A2(G217), .ZN(n1182) );
NOR2_X1 U853 ( .A1(G952), .A2(n1184), .ZN(n1180) );
XNOR2_X1 U854 ( .A(G953), .B(KEYINPUT53), .ZN(n1184) );
NOR2_X1 U855 ( .A1(n1185), .A2(n1186), .ZN(G63) );
XOR2_X1 U856 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U857 ( .A1(n1183), .A2(G478), .ZN(n1187) );
NOR2_X1 U858 ( .A1(n1185), .A2(n1189), .ZN(G60) );
XNOR2_X1 U859 ( .A(n1190), .B(n1134), .ZN(n1189) );
NAND2_X1 U860 ( .A1(n1183), .A2(G475), .ZN(n1190) );
XNOR2_X1 U861 ( .A(G104), .B(n1191), .ZN(G6) );
NAND2_X1 U862 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U863 ( .A1(n1185), .A2(n1194), .ZN(G57) );
XOR2_X1 U864 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U865 ( .A(n1197), .B(n1198), .Z(n1196) );
NAND2_X1 U866 ( .A1(n1183), .A2(G472), .ZN(n1197) );
NOR2_X1 U867 ( .A1(n1185), .A2(n1199), .ZN(G54) );
NOR2_X1 U868 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U869 ( .A(n1202), .B(KEYINPUT11), .Z(n1201) );
NAND2_X1 U870 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
XNOR2_X1 U871 ( .A(n1205), .B(KEYINPUT18), .ZN(n1203) );
NOR2_X1 U872 ( .A1(n1204), .A2(n1205), .ZN(n1200) );
XNOR2_X1 U873 ( .A(n1206), .B(n1207), .ZN(n1205) );
NOR2_X1 U874 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NOR2_X1 U875 ( .A1(n1210), .A2(n1211), .ZN(n1208) );
XNOR2_X1 U876 ( .A(KEYINPUT17), .B(n1212), .ZN(n1211) );
NAND2_X1 U877 ( .A1(n1213), .A2(n1214), .ZN(n1206) );
NAND2_X1 U878 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U879 ( .A(KEYINPUT16), .B(n1217), .Z(n1213) );
NOR2_X1 U880 ( .A1(n1215), .A2(n1216), .ZN(n1217) );
XNOR2_X1 U881 ( .A(n1218), .B(n1219), .ZN(n1216) );
XOR2_X1 U882 ( .A(n1220), .B(n1221), .Z(n1215) );
XNOR2_X1 U883 ( .A(G131), .B(KEYINPUT55), .ZN(n1220) );
AND2_X1 U884 ( .A1(n1183), .A2(n1222), .ZN(n1204) );
XNOR2_X1 U885 ( .A(KEYINPUT38), .B(n1108), .ZN(n1222) );
NOR2_X1 U886 ( .A1(n1185), .A2(n1223), .ZN(G51) );
XNOR2_X1 U887 ( .A(n1224), .B(n1225), .ZN(n1223) );
AND3_X1 U888 ( .A1(n1183), .A2(n1226), .A3(G210), .ZN(n1225) );
INV_X1 U889 ( .A(KEYINPUT32), .ZN(n1226) );
NOR2_X1 U890 ( .A1(n1227), .A2(n1053), .ZN(n1183) );
NOR2_X1 U891 ( .A1(n1179), .A2(n1168), .ZN(n1053) );
NAND4_X1 U892 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1168) );
NOR4_X1 U893 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1231) );
NAND2_X1 U894 ( .A1(n1236), .A2(n1237), .ZN(n1230) );
NAND2_X1 U895 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U896 ( .A1(n1061), .A2(n1240), .ZN(n1238) );
NAND4_X1 U897 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1179) );
AND4_X1 U898 ( .A1(n1245), .A2(n1049), .A3(n1246), .A4(n1247), .ZN(n1244) );
NAND2_X1 U899 ( .A1(n1081), .A2(n1193), .ZN(n1049) );
NOR2_X1 U900 ( .A1(n1248), .A2(n1249), .ZN(n1193) );
NOR2_X1 U901 ( .A1(n1250), .A2(n1251), .ZN(n1243) );
NOR3_X1 U902 ( .A1(n1252), .A2(n1249), .A3(n1079), .ZN(n1251) );
XOR2_X1 U903 ( .A(KEYINPUT6), .B(n1063), .Z(n1252) );
NAND2_X1 U904 ( .A1(n1062), .A2(n1253), .ZN(n1242) );
NAND2_X1 U905 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
OR3_X1 U906 ( .A1(n1249), .A2(KEYINPUT44), .A3(n1256), .ZN(n1255) );
NAND3_X1 U907 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1254) );
NAND2_X1 U908 ( .A1(n1260), .A2(n1083), .ZN(n1258) );
INV_X1 U909 ( .A(n1261), .ZN(n1083) );
NAND4_X1 U910 ( .A1(n1069), .A2(n1262), .A3(n1094), .A4(n1263), .ZN(n1260) );
INV_X1 U911 ( .A(KEYINPUT43), .ZN(n1263) );
NAND2_X1 U912 ( .A1(n1261), .A2(n1264), .ZN(n1257) );
NAND3_X1 U913 ( .A1(n1073), .A2(n1065), .A3(KEYINPUT44), .ZN(n1264) );
NAND2_X1 U914 ( .A1(KEYINPUT43), .A2(n1265), .ZN(n1241) );
NAND2_X1 U915 ( .A1(KEYINPUT51), .A2(n1266), .ZN(n1224) );
XOR2_X1 U916 ( .A(n1267), .B(n1268), .Z(n1266) );
NOR2_X1 U917 ( .A1(KEYINPUT45), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U918 ( .A(n1270), .B(KEYINPUT47), .ZN(n1269) );
NOR2_X1 U919 ( .A1(n1098), .A2(G952), .ZN(n1185) );
XNOR2_X1 U920 ( .A(G146), .B(n1228), .ZN(G48) );
NAND3_X1 U921 ( .A1(n1192), .A2(n1261), .A3(n1271), .ZN(n1228) );
NAND2_X1 U922 ( .A1(n1272), .A2(n1273), .ZN(G45) );
NAND2_X1 U923 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
INV_X1 U924 ( .A(G143), .ZN(n1275) );
XOR2_X1 U925 ( .A(n1276), .B(KEYINPUT19), .Z(n1274) );
NAND2_X1 U926 ( .A1(G143), .A2(n1277), .ZN(n1272) );
XOR2_X1 U927 ( .A(n1276), .B(KEYINPUT5), .Z(n1277) );
NAND3_X1 U928 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1276) );
INV_X1 U929 ( .A(n1239), .ZN(n1280) );
NAND4_X1 U930 ( .A1(n1073), .A2(n1261), .A3(n1281), .A4(n1282), .ZN(n1239) );
XNOR2_X1 U931 ( .A(KEYINPUT31), .B(n1065), .ZN(n1278) );
XNOR2_X1 U932 ( .A(G140), .B(n1283), .ZN(G42) );
NAND4_X1 U933 ( .A1(n1284), .A2(n1061), .A3(n1240), .A4(n1279), .ZN(n1283) );
XNOR2_X1 U934 ( .A(n1285), .B(KEYINPUT15), .ZN(n1284) );
XOR2_X1 U935 ( .A(n1229), .B(n1286), .Z(G39) );
NAND2_X1 U936 ( .A1(KEYINPUT41), .A2(G137), .ZN(n1286) );
NAND3_X1 U937 ( .A1(n1061), .A2(n1062), .A3(n1271), .ZN(n1229) );
XNOR2_X1 U938 ( .A(n1156), .B(n1234), .ZN(G36) );
AND2_X1 U939 ( .A1(n1287), .A2(n1081), .ZN(n1234) );
XNOR2_X1 U940 ( .A(n1288), .B(n1233), .ZN(G33) );
AND2_X1 U941 ( .A1(n1287), .A2(n1192), .ZN(n1233) );
AND3_X1 U942 ( .A1(n1061), .A2(n1073), .A3(n1236), .ZN(n1287) );
AND2_X1 U943 ( .A1(n1086), .A2(n1289), .ZN(n1061) );
XNOR2_X1 U944 ( .A(n1290), .B(n1291), .ZN(G30) );
NOR2_X1 U945 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NOR2_X1 U946 ( .A1(KEYINPUT0), .A2(n1235), .ZN(n1293) );
INV_X1 U947 ( .A(n1294), .ZN(n1235) );
NOR2_X1 U948 ( .A1(KEYINPUT9), .A2(n1294), .ZN(n1292) );
NAND3_X1 U949 ( .A1(n1081), .A2(n1261), .A3(n1271), .ZN(n1294) );
AND3_X1 U950 ( .A1(n1262), .A2(n1094), .A3(n1236), .ZN(n1271) );
AND2_X1 U951 ( .A1(n1285), .A2(n1279), .ZN(n1236) );
XOR2_X1 U952 ( .A(G101), .B(n1295), .Z(G3) );
AND2_X1 U953 ( .A1(n1073), .A2(n1296), .ZN(n1295) );
XOR2_X1 U954 ( .A(G125), .B(n1232), .Z(G27) );
AND4_X1 U955 ( .A1(n1240), .A2(n1069), .A3(n1261), .A4(n1279), .ZN(n1232) );
NAND2_X1 U956 ( .A1(n1091), .A2(n1297), .ZN(n1279) );
NAND4_X1 U957 ( .A1(G902), .A2(G953), .A3(n1298), .A4(n1144), .ZN(n1297) );
INV_X1 U958 ( .A(G900), .ZN(n1144) );
NOR3_X1 U959 ( .A1(n1299), .A2(n1300), .A3(n1079), .ZN(n1240) );
XOR2_X1 U960 ( .A(G122), .B(n1250), .Z(G24) );
AND4_X1 U961 ( .A1(n1301), .A2(n1063), .A3(n1281), .A4(n1282), .ZN(n1250) );
INV_X1 U962 ( .A(n1248), .ZN(n1063) );
NAND2_X1 U963 ( .A1(n1300), .A2(n1093), .ZN(n1248) );
NAND3_X1 U964 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(G21) );
NAND2_X1 U965 ( .A1(G119), .A2(n1305), .ZN(n1304) );
NAND2_X1 U966 ( .A1(KEYINPUT22), .A2(n1306), .ZN(n1303) );
NAND2_X1 U967 ( .A1(n1307), .A2(n1265), .ZN(n1306) );
INV_X1 U968 ( .A(n1305), .ZN(n1265) );
XNOR2_X1 U969 ( .A(KEYINPUT56), .B(G119), .ZN(n1307) );
NAND2_X1 U970 ( .A1(n1308), .A2(n1309), .ZN(n1302) );
INV_X1 U971 ( .A(KEYINPUT22), .ZN(n1309) );
NAND2_X1 U972 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
OR3_X1 U973 ( .A1(n1305), .A2(G119), .A3(KEYINPUT56), .ZN(n1311) );
NAND4_X1 U974 ( .A1(n1062), .A2(n1301), .A3(n1262), .A4(n1094), .ZN(n1305) );
NAND2_X1 U975 ( .A1(KEYINPUT56), .A2(G119), .ZN(n1310) );
XNOR2_X1 U976 ( .A(G116), .B(n1245), .ZN(G18) );
NAND3_X1 U977 ( .A1(n1073), .A2(n1081), .A3(n1301), .ZN(n1245) );
NOR2_X1 U978 ( .A1(n1282), .A2(n1101), .ZN(n1081) );
NAND3_X1 U979 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(G15) );
NAND2_X1 U980 ( .A1(G113), .A2(n1315), .ZN(n1314) );
NAND2_X1 U981 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
INV_X1 U982 ( .A(KEYINPUT57), .ZN(n1317) );
XOR2_X1 U983 ( .A(n1247), .B(KEYINPUT30), .Z(n1316) );
OR3_X1 U984 ( .A1(n1247), .A2(G113), .A3(KEYINPUT57), .ZN(n1313) );
NAND2_X1 U985 ( .A1(KEYINPUT57), .A2(n1247), .ZN(n1312) );
NAND3_X1 U986 ( .A1(n1301), .A2(n1073), .A3(n1192), .ZN(n1247) );
INV_X1 U987 ( .A(n1079), .ZN(n1192) );
NAND2_X1 U988 ( .A1(n1101), .A2(n1282), .ZN(n1079) );
INV_X1 U989 ( .A(n1281), .ZN(n1101) );
INV_X1 U990 ( .A(n1256), .ZN(n1073) );
NAND2_X1 U991 ( .A1(n1300), .A2(n1262), .ZN(n1256) );
XNOR2_X1 U992 ( .A(n1299), .B(KEYINPUT33), .ZN(n1262) );
INV_X1 U993 ( .A(n1093), .ZN(n1299) );
INV_X1 U994 ( .A(n1094), .ZN(n1300) );
AND3_X1 U995 ( .A1(n1261), .A2(n1259), .A3(n1069), .ZN(n1301) );
NOR2_X1 U996 ( .A1(n1068), .A2(n1123), .ZN(n1069) );
INV_X1 U997 ( .A(n1067), .ZN(n1123) );
XNOR2_X1 U998 ( .A(G110), .B(n1246), .ZN(G12) );
NAND3_X1 U999 ( .A1(n1093), .A2(n1094), .A3(n1296), .ZN(n1246) );
NOR2_X1 U1000 ( .A1(n1096), .A2(n1249), .ZN(n1296) );
NAND3_X1 U1001 ( .A1(n1285), .A2(n1259), .A3(n1261), .ZN(n1249) );
NOR2_X1 U1002 ( .A1(n1086), .A2(n1085), .ZN(n1261) );
INV_X1 U1003 ( .A(n1289), .ZN(n1085) );
NAND2_X1 U1004 ( .A1(G214), .A2(n1318), .ZN(n1289) );
XNOR2_X1 U1005 ( .A(n1119), .B(n1319), .ZN(n1086) );
NOR2_X1 U1006 ( .A1(n1118), .A2(KEYINPUT49), .ZN(n1319) );
INV_X1 U1007 ( .A(n1121), .ZN(n1118) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1318), .ZN(n1121) );
NAND2_X1 U1009 ( .A1(n1320), .A2(n1227), .ZN(n1318) );
INV_X1 U1010 ( .A(G237), .ZN(n1320) );
NAND2_X1 U1011 ( .A1(n1130), .A2(n1227), .ZN(n1119) );
XOR2_X1 U1012 ( .A(n1268), .B(n1321), .Z(n1130) );
XNOR2_X1 U1013 ( .A(KEYINPUT52), .B(n1322), .ZN(n1321) );
INV_X1 U1014 ( .A(n1270), .ZN(n1322) );
XNOR2_X1 U1015 ( .A(G125), .B(n1219), .ZN(n1270) );
XNOR2_X1 U1016 ( .A(n1178), .B(n1323), .ZN(n1268) );
NOR2_X1 U1017 ( .A1(n1324), .A2(n1174), .ZN(n1323) );
INV_X1 U1018 ( .A(G224), .ZN(n1174) );
XOR2_X1 U1019 ( .A(n1325), .B(n1326), .Z(n1178) );
XOR2_X1 U1020 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1021 ( .A(G110), .B(G107), .ZN(n1328) );
NAND2_X1 U1022 ( .A1(KEYINPUT21), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1023 ( .A(n1198), .B(n1330), .Z(n1325) );
XNOR2_X1 U1024 ( .A(G101), .B(n1331), .ZN(n1198) );
NAND2_X1 U1025 ( .A1(n1091), .A2(n1332), .ZN(n1259) );
NAND4_X1 U1026 ( .A1(G902), .A2(G953), .A3(n1298), .A4(n1175), .ZN(n1332) );
INV_X1 U1027 ( .A(G898), .ZN(n1175) );
NAND3_X1 U1028 ( .A1(n1298), .A2(n1098), .A3(G952), .ZN(n1091) );
INV_X1 U1029 ( .A(G953), .ZN(n1098) );
NAND2_X1 U1030 ( .A1(n1333), .A2(G237), .ZN(n1298) );
XNOR2_X1 U1031 ( .A(G234), .B(KEYINPUT10), .ZN(n1333) );
INV_X1 U1032 ( .A(n1065), .ZN(n1285) );
NAND2_X1 U1033 ( .A1(n1334), .A2(n1067), .ZN(n1065) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1335), .ZN(n1067) );
XOR2_X1 U1035 ( .A(KEYINPUT48), .B(n1068), .Z(n1334) );
XNOR2_X1 U1036 ( .A(n1109), .B(n1108), .ZN(n1068) );
INV_X1 U1037 ( .A(G469), .ZN(n1108) );
NOR2_X1 U1038 ( .A1(n1129), .A2(G902), .ZN(n1109) );
XOR2_X1 U1039 ( .A(n1336), .B(n1337), .Z(n1129) );
XNOR2_X1 U1040 ( .A(n1338), .B(n1339), .ZN(n1336) );
INV_X1 U1041 ( .A(n1218), .ZN(n1339) );
XNOR2_X1 U1042 ( .A(n1340), .B(n1341), .ZN(n1218) );
XNOR2_X1 U1043 ( .A(n1329), .B(G101), .ZN(n1341) );
NAND2_X1 U1044 ( .A1(KEYINPUT46), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1045 ( .A1(n1343), .A2(n1344), .ZN(n1338) );
NAND2_X1 U1046 ( .A1(n1345), .A2(n1212), .ZN(n1344) );
INV_X1 U1047 ( .A(n1209), .ZN(n1343) );
NOR2_X1 U1048 ( .A1(n1212), .A2(n1345), .ZN(n1209) );
INV_X1 U1049 ( .A(n1210), .ZN(n1345) );
XOR2_X1 U1050 ( .A(G110), .B(n1149), .Z(n1210) );
NAND2_X1 U1051 ( .A1(G227), .A2(n1346), .ZN(n1212) );
INV_X1 U1052 ( .A(n1062), .ZN(n1096) );
NOR2_X1 U1053 ( .A1(n1281), .A2(n1282), .ZN(n1062) );
NAND2_X1 U1054 ( .A1(n1110), .A2(n1347), .ZN(n1282) );
OR3_X1 U1055 ( .A1(G475), .A2(G902), .A3(n1134), .ZN(n1347) );
NAND2_X1 U1056 ( .A1(G475), .A2(n1348), .ZN(n1110) );
NAND2_X1 U1057 ( .A1(n1349), .A2(n1227), .ZN(n1348) );
INV_X1 U1058 ( .A(n1134), .ZN(n1349) );
XNOR2_X1 U1059 ( .A(n1350), .B(n1351), .ZN(n1134) );
XOR2_X1 U1060 ( .A(n1352), .B(n1353), .Z(n1351) );
XNOR2_X1 U1061 ( .A(G113), .B(n1329), .ZN(n1353) );
INV_X1 U1062 ( .A(G104), .ZN(n1329) );
XNOR2_X1 U1063 ( .A(n1288), .B(G122), .ZN(n1352) );
INV_X1 U1064 ( .A(G131), .ZN(n1288) );
XOR2_X1 U1065 ( .A(n1354), .B(n1355), .Z(n1350) );
XNOR2_X1 U1066 ( .A(n1356), .B(n1357), .ZN(n1354) );
NAND2_X1 U1067 ( .A1(KEYINPUT26), .A2(G125), .ZN(n1357) );
NAND2_X1 U1068 ( .A1(n1358), .A2(KEYINPUT2), .ZN(n1356) );
XNOR2_X1 U1069 ( .A(G143), .B(n1359), .ZN(n1358) );
AND2_X1 U1070 ( .A1(n1360), .A2(G214), .ZN(n1359) );
XNOR2_X1 U1071 ( .A(n1361), .B(G478), .ZN(n1281) );
NAND2_X1 U1072 ( .A1(n1362), .A2(n1227), .ZN(n1361) );
XOR2_X1 U1073 ( .A(KEYINPUT60), .B(n1188), .Z(n1362) );
XNOR2_X1 U1074 ( .A(n1363), .B(n1364), .ZN(n1188) );
XOR2_X1 U1075 ( .A(n1365), .B(n1366), .Z(n1364) );
NOR2_X1 U1076 ( .A1(n1367), .A2(n1368), .ZN(n1365) );
XNOR2_X1 U1077 ( .A(n1369), .B(n1156), .ZN(n1363) );
NAND3_X1 U1078 ( .A1(n1370), .A2(n1371), .A3(n1372), .ZN(n1369) );
NAND2_X1 U1079 ( .A1(G107), .A2(n1330), .ZN(n1372) );
NAND2_X1 U1080 ( .A1(n1373), .A2(n1374), .ZN(n1371) );
INV_X1 U1081 ( .A(KEYINPUT28), .ZN(n1374) );
NAND2_X1 U1082 ( .A1(n1375), .A2(n1342), .ZN(n1373) );
INV_X1 U1083 ( .A(G107), .ZN(n1342) );
XNOR2_X1 U1084 ( .A(KEYINPUT35), .B(n1330), .ZN(n1375) );
NAND2_X1 U1085 ( .A1(KEYINPUT28), .A2(n1376), .ZN(n1370) );
NAND2_X1 U1086 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
OR3_X1 U1087 ( .A1(n1330), .A2(G107), .A3(KEYINPUT35), .ZN(n1378) );
NAND2_X1 U1088 ( .A1(KEYINPUT35), .A2(n1330), .ZN(n1377) );
XOR2_X1 U1089 ( .A(G116), .B(G122), .Z(n1330) );
NAND2_X1 U1090 ( .A1(n1379), .A2(n1380), .ZN(n1094) );
NAND2_X1 U1091 ( .A1(KEYINPUT20), .A2(n1132), .ZN(n1380) );
XOR2_X1 U1092 ( .A(n1116), .B(n1381), .Z(n1379) );
NOR2_X1 U1093 ( .A1(KEYINPUT20), .A2(n1132), .ZN(n1381) );
NAND2_X1 U1094 ( .A1(n1382), .A2(n1335), .ZN(n1132) );
NAND2_X1 U1095 ( .A1(G234), .A2(n1227), .ZN(n1335) );
XNOR2_X1 U1096 ( .A(KEYINPUT42), .B(n1368), .ZN(n1382) );
INV_X1 U1097 ( .A(G217), .ZN(n1368) );
NAND2_X1 U1098 ( .A1(n1383), .A2(n1227), .ZN(n1116) );
INV_X1 U1099 ( .A(n1131), .ZN(n1383) );
XNOR2_X1 U1100 ( .A(n1384), .B(n1385), .ZN(n1131) );
XNOR2_X1 U1101 ( .A(n1386), .B(n1387), .ZN(n1385) );
NOR3_X1 U1102 ( .A1(n1388), .A2(KEYINPUT62), .A3(n1367), .ZN(n1387) );
NAND2_X1 U1103 ( .A1(G234), .A2(n1346), .ZN(n1367) );
INV_X1 U1104 ( .A(G221), .ZN(n1388) );
NAND2_X1 U1105 ( .A1(n1389), .A2(KEYINPUT40), .ZN(n1386) );
XOR2_X1 U1106 ( .A(n1390), .B(n1355), .Z(n1389) );
XNOR2_X1 U1107 ( .A(G146), .B(n1149), .ZN(n1355) );
INV_X1 U1108 ( .A(G140), .ZN(n1149) );
XNOR2_X1 U1109 ( .A(G125), .B(KEYINPUT14), .ZN(n1390) );
XOR2_X1 U1110 ( .A(n1391), .B(n1392), .Z(n1384) );
XNOR2_X1 U1111 ( .A(n1162), .B(G110), .ZN(n1392) );
INV_X1 U1112 ( .A(G137), .ZN(n1162) );
NAND2_X1 U1113 ( .A1(n1393), .A2(n1394), .ZN(n1391) );
NAND2_X1 U1114 ( .A1(G119), .A2(n1290), .ZN(n1394) );
XOR2_X1 U1115 ( .A(n1395), .B(KEYINPUT7), .Z(n1393) );
NAND2_X1 U1116 ( .A1(G128), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1117 ( .A(n1397), .B(n1135), .Z(n1093) );
NAND2_X1 U1118 ( .A1(n1398), .A2(n1227), .ZN(n1135) );
INV_X1 U1119 ( .A(G902), .ZN(n1227) );
XOR2_X1 U1120 ( .A(n1195), .B(n1399), .Z(n1398) );
XOR2_X1 U1121 ( .A(n1400), .B(n1331), .Z(n1399) );
XNOR2_X1 U1122 ( .A(G113), .B(n1396), .ZN(n1331) );
INV_X1 U1123 ( .A(G119), .ZN(n1396) );
NOR2_X1 U1124 ( .A1(G101), .A2(KEYINPUT37), .ZN(n1400) );
XOR2_X1 U1125 ( .A(n1401), .B(n1402), .Z(n1195) );
XOR2_X1 U1126 ( .A(KEYINPUT8), .B(G116), .Z(n1402) );
XOR2_X1 U1127 ( .A(n1403), .B(n1337), .Z(n1401) );
XOR2_X1 U1128 ( .A(n1221), .B(n1148), .Z(n1337) );
XNOR2_X1 U1129 ( .A(G131), .B(n1219), .ZN(n1148) );
XNOR2_X1 U1130 ( .A(G146), .B(n1366), .ZN(n1219) );
XNOR2_X1 U1131 ( .A(n1290), .B(G143), .ZN(n1366) );
INV_X1 U1132 ( .A(G128), .ZN(n1290) );
XOR2_X1 U1133 ( .A(G137), .B(n1404), .Z(n1221) );
NOR2_X1 U1134 ( .A1(KEYINPUT29), .A2(n1156), .ZN(n1404) );
INV_X1 U1135 ( .A(G134), .ZN(n1156) );
NAND2_X1 U1136 ( .A1(G210), .A2(n1360), .ZN(n1403) );
NOR2_X1 U1137 ( .A1(n1324), .A2(G237), .ZN(n1360) );
INV_X1 U1138 ( .A(n1346), .ZN(n1324) );
XOR2_X1 U1139 ( .A(G953), .B(KEYINPUT36), .Z(n1346) );
NAND2_X1 U1140 ( .A1(KEYINPUT34), .A2(n1136), .ZN(n1397) );
INV_X1 U1141 ( .A(G472), .ZN(n1136) );
endmodule


