//Key = 1101100110110100011111100011000001110111010101001100010111100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327;

XNOR2_X1 U735 ( .A(G107), .B(n1008), .ZN(G9) );
NAND4_X1 U736 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1008) );
NOR2_X1 U737 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
XNOR2_X1 U738 ( .A(n1015), .B(KEYINPUT61), .ZN(n1014) );
NOR2_X1 U739 ( .A1(n1016), .A2(n1017), .ZN(G75) );
XOR2_X1 U740 ( .A(KEYINPUT59), .B(n1018), .Z(n1017) );
NOR3_X1 U741 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
XOR2_X1 U742 ( .A(KEYINPUT57), .B(n1022), .Z(n1021) );
NAND3_X1 U743 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1019) );
NAND2_X1 U744 ( .A1(n1026), .A2(n1027), .ZN(n1023) );
NAND2_X1 U745 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND4_X1 U746 ( .A1(n1030), .A2(n1031), .A3(n1010), .A4(n1032), .ZN(n1029) );
NAND2_X1 U747 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(n1028) );
NAND2_X1 U749 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U750 ( .A1(n1010), .A2(n1039), .ZN(n1038) );
NAND2_X1 U751 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND3_X1 U752 ( .A1(n1042), .A2(n1030), .A3(n1043), .ZN(n1041) );
NAND2_X1 U753 ( .A1(n1031), .A2(n1044), .ZN(n1037) );
NAND3_X1 U754 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NAND2_X1 U755 ( .A1(n1010), .A2(n1048), .ZN(n1047) );
NAND2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U758 ( .A1(n1030), .A2(n1053), .ZN(n1046) );
NAND2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U760 ( .A1(KEYINPUT21), .A2(n1056), .ZN(n1055) );
OR3_X1 U761 ( .A1(n1057), .A2(KEYINPUT21), .A3(n1030), .ZN(n1045) );
INV_X1 U762 ( .A(n1058), .ZN(n1030) );
INV_X1 U763 ( .A(n1059), .ZN(n1026) );
NOR3_X1 U764 ( .A1(n1060), .A2(G953), .A3(G952), .ZN(n1016) );
INV_X1 U765 ( .A(n1025), .ZN(n1060) );
NAND4_X1 U766 ( .A1(n1010), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1025) );
NOR4_X1 U767 ( .A1(n1043), .A2(n1051), .A3(n1064), .A4(n1065), .ZN(n1063) );
XNOR2_X1 U768 ( .A(G475), .B(n1066), .ZN(n1065) );
NOR2_X1 U769 ( .A1(n1067), .A2(KEYINPUT44), .ZN(n1066) );
NOR3_X1 U770 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1064) );
NOR2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
AND3_X1 U772 ( .A1(n1072), .A2(n1071), .A3(KEYINPUT13), .ZN(n1069) );
AND2_X1 U773 ( .A1(KEYINPUT39), .A2(n1073), .ZN(n1071) );
NOR2_X1 U774 ( .A1(KEYINPUT13), .A2(n1073), .ZN(n1068) );
XNOR2_X1 U775 ( .A(G469), .B(n1074), .ZN(n1061) );
NAND2_X1 U776 ( .A1(KEYINPUT48), .A2(n1075), .ZN(n1074) );
XOR2_X1 U777 ( .A(n1076), .B(n1077), .Z(G72) );
NOR2_X1 U778 ( .A1(n1078), .A2(n1024), .ZN(n1077) );
NOR2_X1 U779 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND3_X1 U780 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1076) );
NAND2_X1 U781 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
OR3_X1 U782 ( .A1(n1085), .A2(n1084), .A3(n1086), .ZN(n1082) );
INV_X1 U783 ( .A(n1087), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1088), .A2(KEYINPUT5), .ZN(n1085) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1086), .ZN(n1081) );
INV_X1 U786 ( .A(KEYINPUT37), .ZN(n1086) );
NAND2_X1 U787 ( .A1(n1088), .A2(n1087), .ZN(n1089) );
NAND2_X1 U788 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND2_X1 U789 ( .A1(G953), .A2(n1080), .ZN(n1091) );
XOR2_X1 U790 ( .A(n1092), .B(n1093), .Z(n1090) );
XNOR2_X1 U791 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U792 ( .A1(KEYINPUT16), .A2(n1096), .ZN(n1095) );
XNOR2_X1 U793 ( .A(n1097), .B(n1098), .ZN(n1092) );
NAND2_X1 U794 ( .A1(KEYINPUT49), .A2(n1099), .ZN(n1098) );
NAND2_X1 U795 ( .A1(KEYINPUT43), .A2(n1100), .ZN(n1097) );
NOR2_X1 U796 ( .A1(G953), .A2(n1101), .ZN(n1088) );
XOR2_X1 U797 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U798 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U799 ( .A1(n1022), .A2(G953), .ZN(n1105) );
NOR2_X1 U800 ( .A1(KEYINPUT25), .A2(n1106), .ZN(n1104) );
NOR3_X1 U801 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
NOR2_X1 U802 ( .A1(G898), .A2(n1024), .ZN(n1109) );
NOR2_X1 U803 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
XOR2_X1 U804 ( .A(n1112), .B(KEYINPUT56), .Z(n1107) );
NAND2_X1 U805 ( .A1(n1110), .A2(n1111), .ZN(n1112) );
XOR2_X1 U806 ( .A(n1113), .B(n1114), .Z(n1110) );
NAND2_X1 U807 ( .A1(G953), .A2(n1115), .ZN(n1102) );
NAND2_X1 U808 ( .A1(G898), .A2(G224), .ZN(n1115) );
NOR2_X1 U809 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XOR2_X1 U810 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U811 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NOR2_X1 U812 ( .A1(n1116), .A2(n1122), .ZN(G63) );
XNOR2_X1 U813 ( .A(n1123), .B(n1124), .ZN(n1122) );
NOR2_X1 U814 ( .A1(n1125), .A2(n1121), .ZN(n1124) );
XNOR2_X1 U815 ( .A(G478), .B(KEYINPUT52), .ZN(n1125) );
NOR2_X1 U816 ( .A1(n1116), .A2(n1126), .ZN(G60) );
XOR2_X1 U817 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U818 ( .A(KEYINPUT15), .B(n1129), .Z(n1128) );
NOR2_X1 U819 ( .A1(n1130), .A2(n1121), .ZN(n1129) );
XOR2_X1 U820 ( .A(G104), .B(n1131), .Z(G6) );
NOR3_X1 U821 ( .A1(n1132), .A2(n1133), .A3(n1033), .ZN(n1131) );
NOR2_X1 U822 ( .A1(n1116), .A2(n1134), .ZN(G57) );
XOR2_X1 U823 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U824 ( .A(n1137), .B(n1138), .Z(n1136) );
AND2_X1 U825 ( .A1(G472), .A2(n1139), .ZN(n1138) );
NOR2_X1 U826 ( .A1(KEYINPUT24), .A2(n1140), .ZN(n1137) );
XNOR2_X1 U827 ( .A(n1141), .B(n1142), .ZN(n1140) );
NOR2_X1 U828 ( .A1(n1116), .A2(n1143), .ZN(G54) );
XOR2_X1 U829 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U830 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U831 ( .A1(n1148), .A2(n1121), .ZN(n1147) );
XOR2_X1 U832 ( .A(n1149), .B(n1150), .Z(n1144) );
NAND2_X1 U833 ( .A1(KEYINPUT45), .A2(n1096), .ZN(n1149) );
XNOR2_X1 U834 ( .A(n1151), .B(KEYINPUT18), .ZN(n1096) );
NOR2_X1 U835 ( .A1(n1116), .A2(n1152), .ZN(G51) );
NOR2_X1 U836 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U837 ( .A(n1155), .B(KEYINPUT7), .Z(n1154) );
NAND3_X1 U838 ( .A1(n1139), .A2(n1156), .A3(n1157), .ZN(n1155) );
XOR2_X1 U839 ( .A(n1158), .B(KEYINPUT54), .Z(n1157) );
INV_X1 U840 ( .A(n1121), .ZN(n1139) );
NOR2_X1 U841 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
XOR2_X1 U842 ( .A(n1158), .B(KEYINPUT12), .Z(n1160) );
XNOR2_X1 U843 ( .A(n1161), .B(n1162), .ZN(n1158) );
NOR2_X1 U844 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U845 ( .A1(n1151), .A2(n1165), .ZN(n1164) );
XNOR2_X1 U846 ( .A(G125), .B(n1166), .ZN(n1165) );
XNOR2_X1 U847 ( .A(KEYINPUT63), .B(KEYINPUT40), .ZN(n1166) );
NOR2_X1 U848 ( .A1(n1072), .A2(n1121), .ZN(n1159) );
NAND2_X1 U849 ( .A1(G902), .A2(n1167), .ZN(n1121) );
NAND2_X1 U850 ( .A1(n1101), .A2(n1022), .ZN(n1167) );
AND4_X1 U851 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1022) );
AND4_X1 U852 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
OR4_X1 U853 ( .A1(n1176), .A2(n1177), .A3(n1133), .A4(n1033), .ZN(n1174) );
NOR2_X1 U854 ( .A1(KEYINPUT4), .A2(n1178), .ZN(n1177) );
NOR3_X1 U855 ( .A1(n1179), .A2(n1009), .A3(n1013), .ZN(n1178) );
AND2_X1 U856 ( .A1(n1132), .A2(KEYINPUT4), .ZN(n1176) );
NOR2_X1 U857 ( .A1(n1180), .A2(n1181), .ZN(n1170) );
NOR3_X1 U858 ( .A1(n1132), .A2(n1034), .A3(n1133), .ZN(n1181) );
INV_X1 U859 ( .A(n1182), .ZN(n1132) );
INV_X1 U860 ( .A(n1020), .ZN(n1101) );
NAND2_X1 U861 ( .A1(n1183), .A2(n1184), .ZN(n1020) );
NOR4_X1 U862 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
NOR4_X1 U863 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1183) );
NOR3_X1 U864 ( .A1(n1193), .A2(n1033), .A3(n1194), .ZN(n1192) );
NOR3_X1 U865 ( .A1(n1195), .A2(n1196), .A3(n1057), .ZN(n1191) );
AND2_X1 U866 ( .A1(G953), .A2(n1197), .ZN(n1116) );
XOR2_X1 U867 ( .A(KEYINPUT55), .B(G952), .Z(n1197) );
XNOR2_X1 U868 ( .A(G146), .B(n1198), .ZN(G48) );
NAND2_X1 U869 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U870 ( .A(KEYINPUT14), .B(n1201), .Z(n1200) );
NOR2_X1 U871 ( .A1(n1193), .A2(n1202), .ZN(n1201) );
XNOR2_X1 U872 ( .A(KEYINPUT19), .B(n1033), .ZN(n1202) );
XOR2_X1 U873 ( .A(G143), .B(n1188), .Z(G45) );
AND4_X1 U874 ( .A1(n1199), .A2(n1009), .A3(n1056), .A4(n1203), .ZN(n1188) );
NOR3_X1 U875 ( .A1(n1062), .A2(n1196), .A3(n1204), .ZN(n1203) );
INV_X1 U876 ( .A(n1194), .ZN(n1199) );
XNOR2_X1 U877 ( .A(n1187), .B(n1205), .ZN(G42) );
XOR2_X1 U878 ( .A(KEYINPUT26), .B(G140), .Z(n1205) );
NOR3_X1 U879 ( .A1(n1054), .A2(n1196), .A3(n1195), .ZN(n1187) );
XOR2_X1 U880 ( .A(G137), .B(n1190), .Z(G39) );
AND3_X1 U881 ( .A1(n1035), .A2(n1031), .A3(n1206), .ZN(n1190) );
XOR2_X1 U882 ( .A(G134), .B(n1189), .Z(G36) );
AND4_X1 U883 ( .A1(n1056), .A2(n1031), .A3(n1207), .A4(n1009), .ZN(n1189) );
NOR2_X1 U884 ( .A1(n1196), .A2(n1034), .ZN(n1207) );
XNOR2_X1 U885 ( .A(G131), .B(n1208), .ZN(G33) );
NAND3_X1 U886 ( .A1(n1056), .A2(n1209), .A3(n1210), .ZN(n1208) );
INV_X1 U887 ( .A(n1195), .ZN(n1210) );
NAND3_X1 U888 ( .A1(n1031), .A2(n1009), .A3(n1211), .ZN(n1195) );
NOR2_X1 U889 ( .A1(n1212), .A2(n1043), .ZN(n1031) );
INV_X1 U890 ( .A(n1042), .ZN(n1212) );
XOR2_X1 U891 ( .A(KEYINPUT27), .B(n1196), .Z(n1209) );
XOR2_X1 U892 ( .A(G128), .B(n1186), .Z(G30) );
NOR3_X1 U893 ( .A1(n1194), .A2(n1034), .A3(n1193), .ZN(n1186) );
INV_X1 U894 ( .A(n1206), .ZN(n1193) );
NOR4_X1 U895 ( .A1(n1049), .A2(n1213), .A3(n1214), .A4(n1196), .ZN(n1206) );
NAND3_X1 U896 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(G3) );
NAND2_X1 U897 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U898 ( .A1(n1220), .A2(n1221), .ZN(n1216) );
INV_X1 U899 ( .A(KEYINPUT35), .ZN(n1221) );
NAND2_X1 U900 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
XNOR2_X1 U901 ( .A(n1218), .B(KEYINPUT2), .ZN(n1222) );
NAND2_X1 U902 ( .A1(KEYINPUT35), .A2(n1224), .ZN(n1215) );
NAND2_X1 U903 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
OR3_X1 U904 ( .A1(n1219), .A2(n1218), .A3(KEYINPUT2), .ZN(n1226) );
INV_X1 U905 ( .A(n1223), .ZN(n1219) );
XOR2_X1 U906 ( .A(G101), .B(KEYINPUT31), .Z(n1223) );
NAND2_X1 U907 ( .A1(KEYINPUT2), .A2(n1218), .ZN(n1225) );
INV_X1 U908 ( .A(n1173), .ZN(n1218) );
NAND3_X1 U909 ( .A1(n1035), .A2(n1056), .A3(n1182), .ZN(n1173) );
XNOR2_X1 U910 ( .A(n1227), .B(n1185), .ZN(G27) );
NOR4_X1 U911 ( .A1(n1040), .A2(n1054), .A3(n1033), .A4(n1196), .ZN(n1185) );
AND2_X1 U912 ( .A1(n1059), .A2(n1228), .ZN(n1196) );
NAND4_X1 U913 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1080), .ZN(n1228) );
INV_X1 U914 ( .A(G900), .ZN(n1080) );
INV_X1 U915 ( .A(n1211), .ZN(n1033) );
INV_X1 U916 ( .A(n1230), .ZN(n1054) );
INV_X1 U917 ( .A(n1231), .ZN(n1040) );
XNOR2_X1 U918 ( .A(G122), .B(n1172), .ZN(G24) );
NAND4_X1 U919 ( .A1(n1231), .A2(n1010), .A3(n1232), .A4(n1233), .ZN(n1172) );
NOR2_X1 U920 ( .A1(n1013), .A2(n1204), .ZN(n1232) );
INV_X1 U921 ( .A(n1133), .ZN(n1010) );
NAND2_X1 U922 ( .A1(n1214), .A2(n1213), .ZN(n1133) );
XNOR2_X1 U923 ( .A(n1180), .B(n1234), .ZN(G21) );
NAND2_X1 U924 ( .A1(KEYINPUT8), .A2(G119), .ZN(n1234) );
AND3_X1 U925 ( .A1(n1231), .A2(n1035), .A3(n1235), .ZN(n1180) );
NOR3_X1 U926 ( .A1(n1213), .A2(n1013), .A3(n1214), .ZN(n1235) );
INV_X1 U927 ( .A(n1236), .ZN(n1214) );
XNOR2_X1 U928 ( .A(G116), .B(n1168), .ZN(G18) );
NAND4_X1 U929 ( .A1(n1231), .A2(n1056), .A3(n1012), .A4(n1237), .ZN(n1168) );
INV_X1 U930 ( .A(n1034), .ZN(n1012) );
NAND2_X1 U931 ( .A1(n1204), .A2(n1233), .ZN(n1034) );
NOR2_X1 U932 ( .A1(n1194), .A2(n1058), .ZN(n1231) );
XOR2_X1 U933 ( .A(n1015), .B(KEYINPUT41), .Z(n1194) );
XNOR2_X1 U934 ( .A(n1169), .B(n1238), .ZN(G15) );
NOR2_X1 U935 ( .A1(KEYINPUT29), .A2(n1239), .ZN(n1238) );
INV_X1 U936 ( .A(G113), .ZN(n1239) );
NAND3_X1 U937 ( .A1(n1211), .A2(n1056), .A3(n1240), .ZN(n1169) );
NOR3_X1 U938 ( .A1(n1058), .A2(n1013), .A3(n1179), .ZN(n1240) );
NAND2_X1 U939 ( .A1(n1052), .A2(n1241), .ZN(n1058) );
INV_X1 U940 ( .A(n1057), .ZN(n1056) );
NAND2_X1 U941 ( .A1(n1213), .A2(n1236), .ZN(n1057) );
NOR2_X1 U942 ( .A1(n1233), .A2(n1204), .ZN(n1211) );
XNOR2_X1 U943 ( .A(G110), .B(n1175), .ZN(G12) );
NAND3_X1 U944 ( .A1(n1230), .A2(n1035), .A3(n1182), .ZN(n1175) );
NOR3_X1 U945 ( .A1(n1179), .A2(n1013), .A3(n1049), .ZN(n1182) );
INV_X1 U946 ( .A(n1009), .ZN(n1049) );
NOR2_X1 U947 ( .A1(n1052), .A2(n1051), .ZN(n1009) );
INV_X1 U948 ( .A(n1241), .ZN(n1051) );
NAND2_X1 U949 ( .A1(G221), .A2(n1242), .ZN(n1241) );
XNOR2_X1 U950 ( .A(n1075), .B(n1148), .ZN(n1052) );
INV_X1 U951 ( .A(G469), .ZN(n1148) );
NAND2_X1 U952 ( .A1(n1243), .A2(n1244), .ZN(n1075) );
XOR2_X1 U953 ( .A(n1245), .B(n1246), .Z(n1243) );
XOR2_X1 U954 ( .A(n1247), .B(n1150), .Z(n1246) );
XNOR2_X1 U955 ( .A(n1248), .B(n1249), .ZN(n1150) );
XOR2_X1 U956 ( .A(G110), .B(n1250), .Z(n1249) );
XOR2_X1 U957 ( .A(KEYINPUT11), .B(G140), .Z(n1250) );
XOR2_X1 U958 ( .A(n1251), .B(n1252), .Z(n1248) );
XNOR2_X1 U959 ( .A(n1141), .B(n1253), .ZN(n1252) );
NOR2_X1 U960 ( .A1(G953), .A2(n1079), .ZN(n1253) );
INV_X1 U961 ( .A(G227), .ZN(n1079) );
INV_X1 U962 ( .A(G101), .ZN(n1141) );
NAND3_X1 U963 ( .A1(n1254), .A2(n1255), .A3(n1256), .ZN(n1251) );
NAND2_X1 U964 ( .A1(G107), .A2(n1257), .ZN(n1256) );
OR3_X1 U965 ( .A1(n1257), .A2(G107), .A3(n1258), .ZN(n1255) );
INV_X1 U966 ( .A(KEYINPUT20), .ZN(n1257) );
NAND2_X1 U967 ( .A1(n1258), .A2(n1259), .ZN(n1254) );
NAND2_X1 U968 ( .A1(n1260), .A2(KEYINPUT20), .ZN(n1259) );
XNOR2_X1 U969 ( .A(G107), .B(KEYINPUT23), .ZN(n1260) );
XOR2_X1 U970 ( .A(KEYINPUT42), .B(KEYINPUT18), .Z(n1245) );
INV_X1 U971 ( .A(n1237), .ZN(n1013) );
NAND2_X1 U972 ( .A1(n1059), .A2(n1261), .ZN(n1237) );
NAND4_X1 U973 ( .A1(G953), .A2(G902), .A3(n1262), .A4(n1263), .ZN(n1261) );
INV_X1 U974 ( .A(G898), .ZN(n1263) );
XNOR2_X1 U975 ( .A(KEYINPUT1), .B(n1229), .ZN(n1262) );
NAND3_X1 U976 ( .A1(n1229), .A2(n1024), .A3(G952), .ZN(n1059) );
NAND2_X1 U977 ( .A1(G237), .A2(G234), .ZN(n1229) );
INV_X1 U978 ( .A(n1015), .ZN(n1179) );
NOR2_X1 U979 ( .A1(n1042), .A2(n1043), .ZN(n1015) );
AND2_X1 U980 ( .A1(G214), .A2(n1264), .ZN(n1043) );
XOR2_X1 U981 ( .A(n1156), .B(n1073), .Z(n1042) );
NAND2_X1 U982 ( .A1(n1265), .A2(n1244), .ZN(n1073) );
XNOR2_X1 U983 ( .A(n1266), .B(n1267), .ZN(n1265) );
INV_X1 U984 ( .A(n1161), .ZN(n1267) );
XNOR2_X1 U985 ( .A(n1268), .B(n1269), .ZN(n1161) );
XOR2_X1 U986 ( .A(n1113), .B(n1111), .Z(n1269) );
XOR2_X1 U987 ( .A(G110), .B(n1270), .Z(n1111) );
XOR2_X1 U988 ( .A(KEYINPUT46), .B(G122), .Z(n1270) );
XOR2_X1 U989 ( .A(n1271), .B(n1272), .Z(n1268) );
XOR2_X1 U990 ( .A(KEYINPUT33), .B(n1273), .Z(n1272) );
AND2_X1 U991 ( .A1(n1024), .A2(G224), .ZN(n1273) );
NAND2_X1 U992 ( .A1(KEYINPUT22), .A2(n1114), .ZN(n1271) );
XOR2_X1 U993 ( .A(n1274), .B(n1258), .Z(n1114) );
XOR2_X1 U994 ( .A(G104), .B(KEYINPUT17), .Z(n1258) );
XNOR2_X1 U995 ( .A(G101), .B(G107), .ZN(n1274) );
NOR4_X1 U996 ( .A1(n1275), .A2(n1276), .A3(KEYINPUT9), .A4(n1163), .ZN(n1266) );
NOR2_X1 U997 ( .A1(n1227), .A2(n1277), .ZN(n1163) );
INV_X1 U998 ( .A(G125), .ZN(n1227) );
NOR3_X1 U999 ( .A1(n1151), .A2(KEYINPUT51), .A3(G125), .ZN(n1276) );
AND2_X1 U1000 ( .A1(n1151), .A2(KEYINPUT51), .ZN(n1275) );
INV_X1 U1001 ( .A(n1072), .ZN(n1156) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1264), .ZN(n1072) );
NAND2_X1 U1003 ( .A1(n1278), .A2(n1244), .ZN(n1264) );
AND2_X1 U1004 ( .A1(n1062), .A2(n1204), .ZN(n1035) );
XNOR2_X1 U1005 ( .A(n1067), .B(n1279), .ZN(n1204) );
XNOR2_X1 U1006 ( .A(KEYINPUT50), .B(n1130), .ZN(n1279) );
INV_X1 U1007 ( .A(G475), .ZN(n1130) );
NOR2_X1 U1008 ( .A1(n1127), .A2(G902), .ZN(n1067) );
XNOR2_X1 U1009 ( .A(n1280), .B(n1281), .ZN(n1127) );
XNOR2_X1 U1010 ( .A(n1282), .B(n1283), .ZN(n1281) );
NAND2_X1 U1011 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND2_X1 U1012 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U1013 ( .A(KEYINPUT34), .B(n1288), .Z(n1284) );
NOR2_X1 U1014 ( .A1(n1287), .A2(n1286), .ZN(n1288) );
XNOR2_X1 U1015 ( .A(G131), .B(n1289), .ZN(n1286) );
NOR2_X1 U1016 ( .A1(KEYINPUT60), .A2(n1290), .ZN(n1289) );
XOR2_X1 U1017 ( .A(n1291), .B(n1292), .Z(n1290) );
AND3_X1 U1018 ( .A1(G214), .A2(n1024), .A3(n1278), .ZN(n1292) );
NAND2_X1 U1019 ( .A1(KEYINPUT62), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U1020 ( .A(G104), .B(n1294), .ZN(n1280) );
XOR2_X1 U1021 ( .A(KEYINPUT28), .B(G122), .Z(n1294) );
INV_X1 U1022 ( .A(n1233), .ZN(n1062) );
XNOR2_X1 U1023 ( .A(n1295), .B(G478), .ZN(n1233) );
NAND2_X1 U1024 ( .A1(n1123), .A2(n1244), .ZN(n1295) );
XNOR2_X1 U1025 ( .A(n1296), .B(n1297), .ZN(n1123) );
XOR2_X1 U1026 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U1027 ( .A1(KEYINPUT36), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U1028 ( .A(n1301), .B(G134), .ZN(n1300) );
AND3_X1 U1029 ( .A1(n1302), .A2(n1024), .A3(G217), .ZN(n1298) );
XNOR2_X1 U1030 ( .A(G107), .B(n1303), .ZN(n1296) );
XOR2_X1 U1031 ( .A(G122), .B(G116), .Z(n1303) );
NOR2_X1 U1032 ( .A1(n1236), .A2(n1213), .ZN(n1230) );
XNOR2_X1 U1033 ( .A(n1304), .B(n1120), .ZN(n1213) );
NAND2_X1 U1034 ( .A1(G217), .A2(n1242), .ZN(n1120) );
NAND2_X1 U1035 ( .A1(G234), .A2(n1244), .ZN(n1242) );
OR2_X1 U1036 ( .A1(n1119), .A2(G902), .ZN(n1304) );
XNOR2_X1 U1037 ( .A(n1305), .B(n1306), .ZN(n1119) );
XOR2_X1 U1038 ( .A(n1307), .B(n1287), .Z(n1306) );
XNOR2_X1 U1039 ( .A(n1308), .B(n1099), .ZN(n1287) );
XNOR2_X1 U1040 ( .A(G140), .B(G125), .ZN(n1099) );
XNOR2_X1 U1041 ( .A(G146), .B(KEYINPUT58), .ZN(n1308) );
NAND2_X1 U1042 ( .A1(KEYINPUT38), .A2(n1309), .ZN(n1307) );
XOR2_X1 U1043 ( .A(G110), .B(n1310), .Z(n1309) );
XOR2_X1 U1044 ( .A(G128), .B(G119), .Z(n1310) );
XOR2_X1 U1045 ( .A(n1311), .B(G137), .Z(n1305) );
NAND3_X1 U1046 ( .A1(G221), .A2(n1024), .A3(n1302), .ZN(n1311) );
XNOR2_X1 U1047 ( .A(G234), .B(KEYINPUT10), .ZN(n1302) );
XNOR2_X1 U1048 ( .A(n1312), .B(G472), .ZN(n1236) );
NAND2_X1 U1049 ( .A1(n1313), .A2(n1244), .ZN(n1312) );
INV_X1 U1050 ( .A(G902), .ZN(n1244) );
XOR2_X1 U1051 ( .A(n1314), .B(n1135), .Z(n1313) );
XNOR2_X1 U1052 ( .A(n1315), .B(n1247), .ZN(n1135) );
XNOR2_X1 U1053 ( .A(n1151), .B(n1146), .ZN(n1247) );
AND2_X1 U1054 ( .A1(n1316), .A2(n1317), .ZN(n1146) );
NAND2_X1 U1055 ( .A1(n1318), .A2(n1094), .ZN(n1317) );
XOR2_X1 U1056 ( .A(KEYINPUT0), .B(n1319), .Z(n1316) );
NOR2_X1 U1057 ( .A1(n1318), .A2(n1094), .ZN(n1319) );
INV_X1 U1058 ( .A(G131), .ZN(n1094) );
INV_X1 U1059 ( .A(n1100), .ZN(n1318) );
XOR2_X1 U1060 ( .A(G134), .B(G137), .Z(n1100) );
INV_X1 U1061 ( .A(n1277), .ZN(n1151) );
XOR2_X1 U1062 ( .A(n1320), .B(n1321), .Z(n1277) );
INV_X1 U1063 ( .A(n1301), .ZN(n1321) );
XNOR2_X1 U1064 ( .A(G128), .B(n1293), .ZN(n1301) );
XNOR2_X1 U1065 ( .A(G143), .B(KEYINPUT6), .ZN(n1293) );
XNOR2_X1 U1066 ( .A(G146), .B(KEYINPUT53), .ZN(n1320) );
XNOR2_X1 U1067 ( .A(n1113), .B(KEYINPUT32), .ZN(n1315) );
XOR2_X1 U1068 ( .A(n1322), .B(n1323), .Z(n1113) );
INV_X1 U1069 ( .A(n1283), .ZN(n1323) );
XOR2_X1 U1070 ( .A(G113), .B(KEYINPUT3), .Z(n1283) );
XNOR2_X1 U1071 ( .A(G116), .B(G119), .ZN(n1322) );
NOR2_X1 U1072 ( .A1(n1324), .A2(n1325), .ZN(n1314) );
XOR2_X1 U1073 ( .A(KEYINPUT47), .B(n1326), .Z(n1325) );
NOR2_X1 U1074 ( .A1(G101), .A2(n1327), .ZN(n1326) );
AND2_X1 U1075 ( .A1(n1327), .A2(G101), .ZN(n1324) );
XOR2_X1 U1076 ( .A(n1142), .B(KEYINPUT30), .Z(n1327) );
AND3_X1 U1077 ( .A1(n1278), .A2(n1024), .A3(G210), .ZN(n1142) );
INV_X1 U1078 ( .A(G953), .ZN(n1024) );
INV_X1 U1079 ( .A(G237), .ZN(n1278) );
endmodule


