//Key = 0110011000011100011000010010110010111000101101110111100011100011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384;

XNOR2_X1 U745 ( .A(G107), .B(n1050), .ZN(G9) );
NAND2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U747 ( .A1(n1053), .A2(n1054), .ZN(G75) );
NOR3_X1 U748 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR2_X1 U749 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U750 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U751 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR3_X1 U752 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1062) );
AND2_X1 U753 ( .A1(n1067), .A2(KEYINPUT15), .ZN(n1066) );
NOR3_X1 U754 ( .A1(KEYINPUT15), .A2(n1068), .A3(n1069), .ZN(n1065) );
NOR3_X1 U755 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1060) );
NOR3_X1 U756 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
AND2_X1 U757 ( .A1(n1076), .A2(KEYINPUT26), .ZN(n1075) );
NOR3_X1 U758 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1074) );
NOR3_X1 U759 ( .A1(n1080), .A2(n1081), .A3(n1051), .ZN(n1079) );
NOR2_X1 U760 ( .A1(n1082), .A2(n1083), .ZN(n1078) );
INV_X1 U761 ( .A(n1067), .ZN(n1073) );
NOR2_X1 U762 ( .A1(n1067), .A2(n1084), .ZN(n1071) );
NOR2_X1 U763 ( .A1(KEYINPUT26), .A2(n1085), .ZN(n1084) );
NAND3_X1 U764 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1055) );
NAND3_X1 U765 ( .A1(n1067), .A2(n1089), .A3(n1090), .ZN(n1088) );
INV_X1 U766 ( .A(n1063), .ZN(n1090) );
NAND4_X1 U767 ( .A1(n1091), .A2(n1082), .A3(n1092), .A4(n1083), .ZN(n1063) );
INV_X1 U768 ( .A(n1070), .ZN(n1091) );
OR2_X1 U769 ( .A1(n1093), .A2(n1094), .ZN(n1089) );
NOR3_X1 U770 ( .A1(n1095), .A2(G953), .A3(G952), .ZN(n1053) );
INV_X1 U771 ( .A(n1086), .ZN(n1095) );
NAND4_X1 U772 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1086) );
NOR4_X1 U773 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
XNOR2_X1 U774 ( .A(n1104), .B(n1105), .ZN(n1103) );
XNOR2_X1 U775 ( .A(n1106), .B(n1107), .ZN(n1102) );
NOR2_X1 U776 ( .A1(KEYINPUT19), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U777 ( .A(KEYINPUT62), .B(n1109), .ZN(n1108) );
XNOR2_X1 U778 ( .A(n1110), .B(n1092), .ZN(n1100) );
XNOR2_X1 U779 ( .A(KEYINPUT47), .B(KEYINPUT37), .ZN(n1110) );
NOR3_X1 U780 ( .A1(n1080), .A2(n1111), .A3(n1112), .ZN(n1098) );
NAND2_X1 U781 ( .A1(n1113), .A2(n1114), .ZN(n1097) );
XNOR2_X1 U782 ( .A(G472), .B(n1115), .ZN(n1096) );
NAND2_X1 U783 ( .A1(KEYINPUT29), .A2(n1116), .ZN(n1115) );
XOR2_X1 U784 ( .A(n1117), .B(n1118), .Z(G72) );
XOR2_X1 U785 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U786 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U787 ( .A1(G953), .A2(n1123), .ZN(n1122) );
XOR2_X1 U788 ( .A(n1124), .B(n1125), .Z(n1121) );
XNOR2_X1 U789 ( .A(n1126), .B(G140), .ZN(n1124) );
NAND2_X1 U790 ( .A1(n1127), .A2(n1128), .ZN(n1119) );
NAND2_X1 U791 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XNOR2_X1 U792 ( .A(G953), .B(KEYINPUT4), .ZN(n1127) );
NOR2_X1 U793 ( .A1(n1131), .A2(n1087), .ZN(n1117) );
NOR2_X1 U794 ( .A1(n1132), .A2(n1123), .ZN(n1131) );
XOR2_X1 U795 ( .A(n1133), .B(n1134), .Z(G69) );
XOR2_X1 U796 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U797 ( .A1(n1137), .A2(n1087), .ZN(n1136) );
NOR2_X1 U798 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U799 ( .A1(n1140), .A2(n1141), .ZN(n1135) );
NAND2_X1 U800 ( .A1(G953), .A2(n1139), .ZN(n1141) );
XNOR2_X1 U801 ( .A(n1142), .B(n1143), .ZN(n1140) );
NAND2_X1 U802 ( .A1(n1087), .A2(n1144), .ZN(n1133) );
NOR2_X1 U803 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XNOR2_X1 U804 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U805 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U806 ( .A1(n1145), .A2(n1151), .ZN(G63) );
NOR3_X1 U807 ( .A1(n1105), .A2(n1152), .A3(n1153), .ZN(n1151) );
NOR4_X1 U808 ( .A1(n1154), .A2(n1150), .A3(KEYINPUT3), .A4(n1104), .ZN(n1153) );
NOR2_X1 U809 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
NOR3_X1 U810 ( .A1(n1104), .A2(KEYINPUT3), .A3(n1157), .ZN(n1155) );
INV_X1 U811 ( .A(G478), .ZN(n1104) );
NOR2_X1 U812 ( .A1(n1145), .A2(n1158), .ZN(G60) );
XOR2_X1 U813 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U814 ( .A(KEYINPUT57), .B(n1161), .Z(n1160) );
AND2_X1 U815 ( .A1(G475), .A2(n1162), .ZN(n1161) );
NAND2_X1 U816 ( .A1(n1163), .A2(n1164), .ZN(G6) );
NAND2_X1 U817 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U818 ( .A(KEYINPUT13), .B(n1167), .Z(n1163) );
NOR2_X1 U819 ( .A1(n1165), .A2(n1166), .ZN(n1167) );
INV_X1 U820 ( .A(n1168), .ZN(n1165) );
NOR2_X1 U821 ( .A1(n1145), .A2(n1169), .ZN(G57) );
XOR2_X1 U822 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U823 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U824 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U825 ( .A1(KEYINPUT42), .A2(n1176), .ZN(n1175) );
NOR2_X1 U826 ( .A1(KEYINPUT8), .A2(n1177), .ZN(n1172) );
XNOR2_X1 U827 ( .A(n1178), .B(n1179), .ZN(n1170) );
XOR2_X1 U828 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U829 ( .A1(KEYINPUT60), .A2(n1182), .ZN(n1181) );
NOR2_X1 U830 ( .A1(n1183), .A2(n1150), .ZN(n1180) );
NOR3_X1 U831 ( .A1(n1145), .A2(n1184), .A3(n1185), .ZN(G54) );
NOR2_X1 U832 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U833 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
NOR2_X1 U834 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U835 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
NOR2_X1 U836 ( .A1(n1194), .A2(n1195), .ZN(n1184) );
NOR2_X1 U837 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NOR2_X1 U838 ( .A1(n1193), .A2(n1191), .ZN(n1197) );
XOR2_X1 U839 ( .A(n1198), .B(n1192), .Z(n1191) );
XNOR2_X1 U840 ( .A(KEYINPUT63), .B(KEYINPUT51), .ZN(n1198) );
NOR2_X1 U841 ( .A1(n1192), .A2(n1190), .ZN(n1196) );
INV_X1 U842 ( .A(n1193), .ZN(n1190) );
NAND2_X1 U843 ( .A1(n1199), .A2(n1200), .ZN(n1193) );
NAND2_X1 U844 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND2_X1 U845 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NAND2_X1 U846 ( .A1(n1182), .A2(n1205), .ZN(n1204) );
INV_X1 U847 ( .A(n1126), .ZN(n1182) );
INV_X1 U848 ( .A(n1206), .ZN(n1201) );
NAND2_X1 U849 ( .A1(n1126), .A2(n1207), .ZN(n1199) );
NAND2_X1 U850 ( .A1(n1205), .A2(n1208), .ZN(n1207) );
NAND2_X1 U851 ( .A1(n1206), .A2(n1203), .ZN(n1208) );
INV_X1 U852 ( .A(KEYINPUT33), .ZN(n1203) );
INV_X1 U853 ( .A(KEYINPUT39), .ZN(n1205) );
AND2_X1 U854 ( .A1(n1162), .A2(G469), .ZN(n1192) );
INV_X1 U855 ( .A(n1187), .ZN(n1194) );
NAND2_X1 U856 ( .A1(KEYINPUT52), .A2(n1209), .ZN(n1187) );
XOR2_X1 U857 ( .A(n1210), .B(n1211), .Z(n1209) );
NAND2_X1 U858 ( .A1(KEYINPUT43), .A2(n1212), .ZN(n1210) );
NOR2_X1 U859 ( .A1(n1145), .A2(n1213), .ZN(G51) );
XOR2_X1 U860 ( .A(n1214), .B(n1215), .Z(n1213) );
XOR2_X1 U861 ( .A(n1216), .B(n1217), .Z(n1215) );
NOR2_X1 U862 ( .A1(n1109), .A2(n1150), .ZN(n1216) );
INV_X1 U863 ( .A(n1162), .ZN(n1150) );
NOR2_X1 U864 ( .A1(n1218), .A2(n1157), .ZN(n1162) );
INV_X1 U865 ( .A(n1057), .ZN(n1157) );
NAND3_X1 U866 ( .A1(n1129), .A2(n1219), .A3(n1220), .ZN(n1057) );
INV_X1 U867 ( .A(n1144), .ZN(n1220) );
NAND4_X1 U868 ( .A1(n1221), .A2(n1168), .A3(n1222), .A4(n1223), .ZN(n1144) );
AND4_X1 U869 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
NAND2_X1 U870 ( .A1(n1082), .A2(n1228), .ZN(n1222) );
NAND2_X1 U871 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND4_X1 U872 ( .A1(n1093), .A2(n1231), .A3(n1064), .A4(n1232), .ZN(n1230) );
NOR2_X1 U873 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U874 ( .A1(n1235), .A2(n1236), .ZN(n1229) );
NAND2_X1 U875 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND2_X1 U876 ( .A1(n1093), .A2(n1234), .ZN(n1238) );
INV_X1 U877 ( .A(KEYINPUT14), .ZN(n1234) );
INV_X1 U878 ( .A(n1094), .ZN(n1237) );
NAND2_X1 U879 ( .A1(n1081), .A2(n1052), .ZN(n1168) );
NOR2_X1 U880 ( .A1(n1059), .A2(n1239), .ZN(n1052) );
INV_X1 U881 ( .A(n1240), .ZN(n1059) );
NAND4_X1 U882 ( .A1(n1051), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1221) );
NAND2_X1 U883 ( .A1(KEYINPUT50), .A2(n1239), .ZN(n1242) );
NAND2_X1 U884 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
INV_X1 U885 ( .A(KEYINPUT50), .ZN(n1244) );
NAND3_X1 U886 ( .A1(n1245), .A2(n1233), .A3(n1231), .ZN(n1243) );
XOR2_X1 U887 ( .A(KEYINPUT22), .B(n1130), .Z(n1219) );
AND3_X1 U888 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1130) );
NAND2_X1 U889 ( .A1(n1051), .A2(n1249), .ZN(n1248) );
NAND2_X1 U890 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND3_X1 U891 ( .A1(n1064), .A2(n1231), .A3(n1252), .ZN(n1251) );
NAND2_X1 U892 ( .A1(n1253), .A2(n1067), .ZN(n1250) );
AND4_X1 U893 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1129) );
NOR2_X1 U894 ( .A1(n1258), .A2(n1259), .ZN(n1254) );
NOR2_X1 U895 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U896 ( .A(KEYINPUT18), .ZN(n1260) );
NOR3_X1 U897 ( .A1(KEYINPUT18), .A2(n1262), .A3(n1245), .ZN(n1258) );
NOR2_X1 U898 ( .A1(n1087), .A2(G952), .ZN(n1145) );
XOR2_X1 U899 ( .A(n1263), .B(G146), .Z(G48) );
NAND2_X1 U900 ( .A1(KEYINPUT23), .A2(n1261), .ZN(n1263) );
NAND2_X1 U901 ( .A1(n1262), .A2(n1064), .ZN(n1261) );
AND3_X1 U902 ( .A1(n1081), .A2(n1264), .A3(n1252), .ZN(n1262) );
XNOR2_X1 U903 ( .A(G143), .B(n1255), .ZN(G45) );
NAND4_X1 U904 ( .A1(n1253), .A2(n1064), .A3(n1265), .A4(n1101), .ZN(n1255) );
XNOR2_X1 U905 ( .A(n1266), .B(n1256), .ZN(G42) );
NAND3_X1 U906 ( .A1(n1067), .A2(n1264), .A3(n1267), .ZN(n1256) );
NAND2_X1 U907 ( .A1(KEYINPUT34), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U908 ( .A(G137), .B(n1257), .ZN(G39) );
NAND3_X1 U909 ( .A1(n1067), .A2(n1076), .A3(n1252), .ZN(n1257) );
INV_X1 U910 ( .A(n1085), .ZN(n1076) );
NAND2_X1 U911 ( .A1(n1082), .A2(n1264), .ZN(n1085) );
XOR2_X1 U912 ( .A(G134), .B(n1269), .Z(G36) );
NOR3_X1 U913 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1269) );
INV_X1 U914 ( .A(n1051), .ZN(n1272) );
XNOR2_X1 U915 ( .A(n1067), .B(KEYINPUT7), .ZN(n1271) );
XNOR2_X1 U916 ( .A(G131), .B(n1246), .ZN(G33) );
NAND3_X1 U917 ( .A1(n1067), .A2(n1081), .A3(n1253), .ZN(n1246) );
INV_X1 U918 ( .A(n1270), .ZN(n1253) );
NAND3_X1 U919 ( .A1(n1093), .A2(n1273), .A3(n1264), .ZN(n1270) );
NOR2_X1 U920 ( .A1(n1068), .A2(n1112), .ZN(n1067) );
INV_X1 U921 ( .A(n1069), .ZN(n1112) );
XNOR2_X1 U922 ( .A(G128), .B(n1274), .ZN(G30) );
NAND4_X1 U923 ( .A1(n1275), .A2(n1252), .A3(n1051), .A4(n1231), .ZN(n1274) );
AND3_X1 U924 ( .A1(n1273), .A2(n1276), .A3(n1277), .ZN(n1252) );
XNOR2_X1 U925 ( .A(n1064), .B(KEYINPUT56), .ZN(n1275) );
XNOR2_X1 U926 ( .A(G101), .B(n1278), .ZN(G3) );
NAND3_X1 U927 ( .A1(n1235), .A2(n1093), .A3(n1082), .ZN(n1278) );
XNOR2_X1 U928 ( .A(G125), .B(n1247), .ZN(G27) );
NAND4_X1 U929 ( .A1(n1092), .A2(n1267), .A3(n1064), .A4(n1083), .ZN(n1247) );
AND3_X1 U930 ( .A1(n1094), .A2(n1273), .A3(n1081), .ZN(n1267) );
NAND2_X1 U931 ( .A1(n1279), .A2(n1280), .ZN(n1273) );
NAND4_X1 U932 ( .A1(G953), .A2(G902), .A3(n1281), .A4(n1123), .ZN(n1280) );
INV_X1 U933 ( .A(G900), .ZN(n1123) );
XNOR2_X1 U934 ( .A(KEYINPUT12), .B(n1070), .ZN(n1279) );
NAND2_X1 U935 ( .A1(n1282), .A2(n1283), .ZN(G24) );
NAND2_X1 U936 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U937 ( .A(n1226), .B(KEYINPUT36), .Z(n1284) );
NAND2_X1 U938 ( .A1(G122), .A2(n1286), .ZN(n1282) );
XOR2_X1 U939 ( .A(n1226), .B(KEYINPUT16), .Z(n1286) );
NAND4_X1 U940 ( .A1(n1287), .A2(n1240), .A3(n1265), .A4(n1101), .ZN(n1226) );
XNOR2_X1 U941 ( .A(n1288), .B(n1289), .ZN(G21) );
NOR2_X1 U942 ( .A1(KEYINPUT48), .A2(n1227), .ZN(n1289) );
NAND4_X1 U943 ( .A1(n1082), .A2(n1287), .A3(n1277), .A4(n1276), .ZN(n1227) );
XOR2_X1 U944 ( .A(n1225), .B(n1290), .Z(G18) );
XNOR2_X1 U945 ( .A(KEYINPUT58), .B(n1291), .ZN(n1290) );
NAND3_X1 U946 ( .A1(n1051), .A2(n1093), .A3(n1287), .ZN(n1225) );
NOR2_X1 U947 ( .A1(n1101), .A2(n1292), .ZN(n1051) );
XNOR2_X1 U948 ( .A(G113), .B(n1224), .ZN(G15) );
NAND3_X1 U949 ( .A1(n1287), .A2(n1093), .A3(n1081), .ZN(n1224) );
AND2_X1 U950 ( .A1(n1292), .A2(n1101), .ZN(n1081) );
NAND2_X1 U951 ( .A1(n1293), .A2(n1294), .ZN(n1093) );
NAND2_X1 U952 ( .A1(n1240), .A2(n1295), .ZN(n1294) );
OR3_X1 U953 ( .A1(n1276), .A2(n1296), .A3(n1295), .ZN(n1293) );
INV_X1 U954 ( .A(KEYINPUT6), .ZN(n1295) );
AND4_X1 U955 ( .A1(n1092), .A2(n1064), .A3(n1233), .A4(n1083), .ZN(n1287) );
XNOR2_X1 U956 ( .A(G110), .B(n1297), .ZN(G12) );
NAND3_X1 U957 ( .A1(n1298), .A2(n1094), .A3(n1235), .ZN(n1297) );
INV_X1 U958 ( .A(n1239), .ZN(n1235) );
NAND3_X1 U959 ( .A1(n1231), .A2(n1233), .A3(n1064), .ZN(n1239) );
INV_X1 U960 ( .A(n1245), .ZN(n1064) );
NAND2_X1 U961 ( .A1(n1068), .A2(n1069), .ZN(n1245) );
NAND2_X1 U962 ( .A1(G214), .A2(n1299), .ZN(n1069) );
XOR2_X1 U963 ( .A(n1107), .B(n1109), .Z(n1068) );
NAND2_X1 U964 ( .A1(G210), .A2(n1299), .ZN(n1109) );
NAND2_X1 U965 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
INV_X1 U966 ( .A(G237), .ZN(n1301) );
NAND2_X1 U967 ( .A1(n1302), .A2(n1218), .ZN(n1107) );
XNOR2_X1 U968 ( .A(n1217), .B(n1303), .ZN(n1302) );
NOR2_X1 U969 ( .A1(KEYINPUT41), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U970 ( .A(n1214), .B(n1305), .ZN(n1304) );
XNOR2_X1 U971 ( .A(KEYINPUT17), .B(KEYINPUT0), .ZN(n1305) );
XOR2_X1 U972 ( .A(n1125), .B(n1306), .Z(n1214) );
NOR2_X1 U973 ( .A1(G953), .A2(n1138), .ZN(n1306) );
INV_X1 U974 ( .A(G224), .ZN(n1138) );
XOR2_X1 U975 ( .A(n1178), .B(G125), .Z(n1125) );
XOR2_X1 U976 ( .A(n1307), .B(n1142), .Z(n1217) );
XNOR2_X1 U977 ( .A(G110), .B(G122), .ZN(n1142) );
NAND2_X1 U978 ( .A1(n1308), .A2(n1143), .ZN(n1307) );
XNOR2_X1 U979 ( .A(n1309), .B(n1310), .ZN(n1143) );
XOR2_X1 U980 ( .A(n1311), .B(n1312), .Z(n1310) );
XNOR2_X1 U981 ( .A(G119), .B(n1313), .ZN(n1312) );
NAND2_X1 U982 ( .A1(KEYINPUT5), .A2(n1176), .ZN(n1313) );
NOR2_X1 U983 ( .A1(G113), .A2(KEYINPUT27), .ZN(n1311) );
XOR2_X1 U984 ( .A(n1314), .B(n1315), .Z(n1309) );
NAND2_X1 U985 ( .A1(KEYINPUT2), .A2(n1291), .ZN(n1314) );
INV_X1 U986 ( .A(G116), .ZN(n1291) );
XOR2_X1 U987 ( .A(KEYINPUT61), .B(KEYINPUT1), .Z(n1308) );
NAND2_X1 U988 ( .A1(n1070), .A2(n1316), .ZN(n1233) );
NAND4_X1 U989 ( .A1(G953), .A2(G902), .A3(n1281), .A4(n1139), .ZN(n1316) );
INV_X1 U990 ( .A(G898), .ZN(n1139) );
NAND3_X1 U991 ( .A1(n1281), .A2(n1087), .A3(G952), .ZN(n1070) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n1281) );
XOR2_X1 U993 ( .A(n1264), .B(KEYINPUT54), .Z(n1231) );
NOR2_X1 U994 ( .A1(n1092), .A2(n1080), .ZN(n1264) );
INV_X1 U995 ( .A(n1083), .ZN(n1080) );
NAND2_X1 U996 ( .A1(G221), .A2(n1317), .ZN(n1083) );
INV_X1 U997 ( .A(n1077), .ZN(n1092) );
XNOR2_X1 U998 ( .A(n1318), .B(G469), .ZN(n1077) );
NAND2_X1 U999 ( .A1(n1319), .A2(n1218), .ZN(n1318) );
XOR2_X1 U1000 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1001 ( .A(n1322), .B(n1211), .Z(n1321) );
XNOR2_X1 U1002 ( .A(G110), .B(n1323), .ZN(n1211) );
NOR2_X1 U1003 ( .A1(G953), .A2(n1132), .ZN(n1323) );
INV_X1 U1004 ( .A(G227), .ZN(n1132) );
NAND2_X1 U1005 ( .A1(KEYINPUT46), .A2(n1126), .ZN(n1322) );
XNOR2_X1 U1006 ( .A(n1324), .B(n1212), .ZN(n1320) );
XOR2_X1 U1007 ( .A(n1268), .B(KEYINPUT20), .Z(n1212) );
INV_X1 U1008 ( .A(G140), .ZN(n1268) );
NAND2_X1 U1009 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
OR2_X1 U1010 ( .A1(n1206), .A2(KEYINPUT31), .ZN(n1326) );
XOR2_X1 U1011 ( .A(n1327), .B(n1328), .Z(n1206) );
INV_X1 U1012 ( .A(n1178), .ZN(n1328) );
NAND3_X1 U1013 ( .A1(n1327), .A2(n1178), .A3(KEYINPUT31), .ZN(n1325) );
XNOR2_X1 U1014 ( .A(n1315), .B(n1176), .ZN(n1327) );
XOR2_X1 U1015 ( .A(G104), .B(n1329), .Z(n1315) );
NAND2_X1 U1016 ( .A1(n1330), .A2(n1331), .ZN(n1094) );
NAND3_X1 U1017 ( .A1(n1296), .A2(n1276), .A3(n1332), .ZN(n1331) );
INV_X1 U1018 ( .A(KEYINPUT55), .ZN(n1332) );
INV_X1 U1019 ( .A(n1277), .ZN(n1296) );
NAND2_X1 U1020 ( .A1(KEYINPUT55), .A2(n1240), .ZN(n1330) );
NOR2_X1 U1021 ( .A1(n1276), .A2(n1277), .ZN(n1240) );
XOR2_X1 U1022 ( .A(n1116), .B(n1183), .Z(n1277) );
INV_X1 U1023 ( .A(G472), .ZN(n1183) );
NAND2_X1 U1024 ( .A1(n1333), .A2(n1218), .ZN(n1116) );
XOR2_X1 U1025 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1026 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1027 ( .A(n1174), .B(n1176), .ZN(n1337) );
INV_X1 U1028 ( .A(G101), .ZN(n1176) );
NAND2_X1 U1029 ( .A1(G210), .A2(n1338), .ZN(n1174) );
XNOR2_X1 U1030 ( .A(KEYINPUT49), .B(KEYINPUT10), .ZN(n1336) );
XOR2_X1 U1031 ( .A(n1339), .B(n1177), .Z(n1334) );
XNOR2_X1 U1032 ( .A(n1340), .B(n1341), .ZN(n1177) );
XNOR2_X1 U1033 ( .A(n1288), .B(G113), .ZN(n1341) );
INV_X1 U1034 ( .A(G119), .ZN(n1288) );
NAND2_X1 U1035 ( .A1(KEYINPUT35), .A2(G116), .ZN(n1340) );
XNOR2_X1 U1036 ( .A(n1126), .B(n1178), .ZN(n1339) );
XOR2_X1 U1037 ( .A(G128), .B(n1342), .Z(n1178) );
XOR2_X1 U1038 ( .A(G146), .B(G143), .Z(n1342) );
XOR2_X1 U1039 ( .A(G131), .B(n1343), .Z(n1126) );
XOR2_X1 U1040 ( .A(G137), .B(G134), .Z(n1343) );
NAND3_X1 U1041 ( .A1(n1344), .A2(n1345), .A3(n1346), .ZN(n1276) );
INV_X1 U1042 ( .A(n1111), .ZN(n1346) );
NOR2_X1 U1043 ( .A1(n1114), .A2(n1113), .ZN(n1111) );
NAND2_X1 U1044 ( .A1(KEYINPUT25), .A2(n1149), .ZN(n1345) );
NAND3_X1 U1045 ( .A1(n1114), .A2(n1347), .A3(n1113), .ZN(n1344) );
INV_X1 U1046 ( .A(n1149), .ZN(n1113) );
NAND2_X1 U1047 ( .A1(G217), .A2(n1317), .ZN(n1149) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1300), .ZN(n1317) );
XNOR2_X1 U1049 ( .A(n1218), .B(KEYINPUT28), .ZN(n1300) );
INV_X1 U1050 ( .A(KEYINPUT25), .ZN(n1347) );
NAND2_X1 U1051 ( .A1(n1147), .A2(n1218), .ZN(n1114) );
XNOR2_X1 U1052 ( .A(n1348), .B(n1349), .ZN(n1147) );
XNOR2_X1 U1053 ( .A(G137), .B(n1350), .ZN(n1349) );
NAND3_X1 U1054 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1350) );
NAND2_X1 U1055 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
INV_X1 U1056 ( .A(KEYINPUT32), .ZN(n1355) );
NAND3_X1 U1057 ( .A1(KEYINPUT32), .A2(n1356), .A3(n1357), .ZN(n1352) );
OR2_X1 U1058 ( .A1(n1357), .A2(n1356), .ZN(n1351) );
NOR2_X1 U1059 ( .A1(n1358), .A2(n1354), .ZN(n1356) );
XOR2_X1 U1060 ( .A(G110), .B(n1359), .Z(n1354) );
NOR2_X1 U1061 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
XOR2_X1 U1062 ( .A(KEYINPUT24), .B(n1362), .Z(n1361) );
NOR2_X1 U1063 ( .A1(G119), .A2(n1363), .ZN(n1362) );
AND2_X1 U1064 ( .A1(n1363), .A2(G119), .ZN(n1360) );
XOR2_X1 U1065 ( .A(G128), .B(KEYINPUT11), .Z(n1363) );
INV_X1 U1066 ( .A(KEYINPUT40), .ZN(n1358) );
NAND2_X1 U1067 ( .A1(G221), .A2(n1364), .ZN(n1348) );
XOR2_X1 U1068 ( .A(KEYINPUT44), .B(n1082), .Z(n1298) );
NOR2_X1 U1069 ( .A1(n1101), .A2(n1265), .ZN(n1082) );
INV_X1 U1070 ( .A(n1292), .ZN(n1265) );
XOR2_X1 U1071 ( .A(n1105), .B(n1365), .Z(n1292) );
NOR2_X1 U1072 ( .A1(G478), .A2(KEYINPUT38), .ZN(n1365) );
NOR2_X1 U1073 ( .A1(n1156), .A2(G902), .ZN(n1105) );
INV_X1 U1074 ( .A(n1154), .ZN(n1156) );
XNOR2_X1 U1075 ( .A(n1366), .B(n1367), .ZN(n1154) );
NOR2_X1 U1076 ( .A1(KEYINPUT9), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1077 ( .A(n1369), .B(n1370), .Z(n1368) );
XNOR2_X1 U1078 ( .A(n1329), .B(n1371), .ZN(n1370) );
XNOR2_X1 U1079 ( .A(G116), .B(n1372), .ZN(n1371) );
NOR2_X1 U1080 ( .A1(G128), .A2(KEYINPUT59), .ZN(n1372) );
XOR2_X1 U1081 ( .A(G107), .B(KEYINPUT53), .Z(n1329) );
XNOR2_X1 U1082 ( .A(n1285), .B(n1373), .ZN(n1369) );
XOR2_X1 U1083 ( .A(G143), .B(G134), .Z(n1373) );
INV_X1 U1084 ( .A(G122), .ZN(n1285) );
NAND2_X1 U1085 ( .A1(G217), .A2(n1364), .ZN(n1366) );
AND2_X1 U1086 ( .A1(G234), .A2(n1087), .ZN(n1364) );
INV_X1 U1087 ( .A(G953), .ZN(n1087) );
XNOR2_X1 U1088 ( .A(n1374), .B(G475), .ZN(n1101) );
NAND2_X1 U1089 ( .A1(n1159), .A2(n1218), .ZN(n1374) );
INV_X1 U1090 ( .A(G902), .ZN(n1218) );
XOR2_X1 U1091 ( .A(n1375), .B(n1376), .Z(n1159) );
XNOR2_X1 U1092 ( .A(n1166), .B(n1377), .ZN(n1376) );
NOR2_X1 U1093 ( .A1(KEYINPUT30), .A2(n1378), .ZN(n1377) );
XOR2_X1 U1094 ( .A(n1379), .B(n1380), .Z(n1378) );
XOR2_X1 U1095 ( .A(n1357), .B(n1381), .Z(n1380) );
NOR2_X1 U1096 ( .A1(G131), .A2(KEYINPUT21), .ZN(n1381) );
XOR2_X1 U1097 ( .A(n1382), .B(n1383), .Z(n1357) );
XOR2_X1 U1098 ( .A(KEYINPUT45), .B(G146), .Z(n1383) );
XNOR2_X1 U1099 ( .A(G125), .B(G140), .ZN(n1382) );
XOR2_X1 U1100 ( .A(n1384), .B(G143), .Z(n1379) );
NAND2_X1 U1101 ( .A1(G214), .A2(n1338), .ZN(n1384) );
NOR2_X1 U1102 ( .A1(G953), .A2(G237), .ZN(n1338) );
INV_X1 U1103 ( .A(G104), .ZN(n1166) );
XNOR2_X1 U1104 ( .A(G113), .B(G122), .ZN(n1375) );
endmodule


