//Key = 0010100100011000101101101110101001101100111110001000111110011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372;

XNOR2_X1 U752 ( .A(n1041), .B(n1042), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U754 ( .A1(n1045), .A2(n1046), .ZN(G75) );
AND4_X1 U755 ( .A1(n1047), .A2(n1048), .A3(KEYINPUT42), .A4(n1049), .ZN(n1046) );
NOR4_X1 U756 ( .A1(G953), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1049) );
NOR4_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NOR3_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1054) );
NOR2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U763 ( .A1(KEYINPUT32), .A2(n1068), .ZN(n1067) );
NOR2_X1 U764 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
XOR2_X1 U765 ( .A(KEYINPUT18), .B(n1071), .Z(n1070) );
NOR2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1062) );
NOR2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1053) );
AND4_X1 U769 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(KEYINPUT32), .ZN(n1077) );
INV_X1 U770 ( .A(n1057), .ZN(n1076) );
NOR4_X1 U771 ( .A1(n1081), .A2(n1073), .A3(n1065), .A4(n1057), .ZN(n1051) );
INV_X1 U772 ( .A(n1080), .ZN(n1065) );
INV_X1 U773 ( .A(n1082), .ZN(n1073) );
NOR2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR2_X1 U775 ( .A1(n1085), .A2(n1061), .ZN(n1084) );
INV_X1 U776 ( .A(n1079), .ZN(n1061) );
NOR2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U778 ( .A(n1088), .B(KEYINPUT54), .ZN(n1087) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1056), .ZN(n1086) );
NOR4_X1 U780 ( .A1(n1090), .A2(n1056), .A3(n1055), .A4(n1091), .ZN(n1083) );
XNOR2_X1 U781 ( .A(n1092), .B(KEYINPUT26), .ZN(n1090) );
NOR3_X1 U782 ( .A1(n1050), .A2(G953), .A3(G952), .ZN(n1045) );
AND4_X1 U783 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1050) );
NOR4_X1 U784 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XNOR2_X1 U785 ( .A(n1056), .B(KEYINPUT30), .ZN(n1098) );
XOR2_X1 U786 ( .A(n1101), .B(KEYINPUT22), .Z(n1097) );
NOR2_X1 U787 ( .A1(n1102), .A2(n1071), .ZN(n1095) );
XNOR2_X1 U788 ( .A(n1103), .B(n1104), .ZN(n1094) );
NAND2_X1 U789 ( .A1(KEYINPUT52), .A2(n1105), .ZN(n1104) );
XNOR2_X1 U790 ( .A(n1106), .B(n1107), .ZN(n1093) );
NOR2_X1 U791 ( .A1(n1108), .A2(KEYINPUT8), .ZN(n1107) );
XOR2_X1 U792 ( .A(n1109), .B(n1110), .Z(G72) );
NOR2_X1 U793 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR3_X1 U795 ( .A1(KEYINPUT29), .A2(n1115), .A3(n1116), .ZN(n1109) );
NOR2_X1 U796 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
INV_X1 U797 ( .A(n1119), .ZN(n1118) );
NOR2_X1 U798 ( .A1(n1120), .A2(n1119), .ZN(n1115) );
XNOR2_X1 U799 ( .A(n1121), .B(n1122), .ZN(n1119) );
XOR2_X1 U800 ( .A(KEYINPUT46), .B(KEYINPUT36), .Z(n1122) );
XNOR2_X1 U801 ( .A(n1123), .B(n1124), .ZN(n1121) );
NOR2_X1 U802 ( .A1(n1125), .A2(n1117), .ZN(n1120) );
NOR2_X1 U803 ( .A1(G953), .A2(n1047), .ZN(n1117) );
NOR2_X1 U804 ( .A1(G900), .A2(n1112), .ZN(n1125) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(G69) );
NOR2_X1 U806 ( .A1(n1128), .A2(n1112), .ZN(n1127) );
NOR2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1126) );
NAND3_X1 U809 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
NAND2_X1 U810 ( .A1(n1136), .A2(n1137), .ZN(n1131) );
NAND2_X1 U811 ( .A1(n1135), .A2(n1134), .ZN(n1137) );
NAND2_X1 U812 ( .A1(n1138), .A2(n1130), .ZN(n1134) );
XNOR2_X1 U813 ( .A(KEYINPUT13), .B(n1112), .ZN(n1138) );
XOR2_X1 U814 ( .A(n1133), .B(KEYINPUT12), .Z(n1136) );
NAND2_X1 U815 ( .A1(n1112), .A2(n1139), .ZN(n1133) );
NOR3_X1 U816 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(G66) );
NOR2_X1 U817 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U818 ( .A(KEYINPUT11), .B(n1145), .Z(n1144) );
NOR2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1141) );
INV_X1 U820 ( .A(n1143), .ZN(n1146) );
NOR3_X1 U821 ( .A1(KEYINPUT38), .A2(n1147), .A3(n1148), .ZN(n1143) );
NOR2_X1 U822 ( .A1(n1140), .A2(n1149), .ZN(G63) );
XNOR2_X1 U823 ( .A(n1150), .B(n1151), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1148), .ZN(n1151) );
NOR2_X1 U825 ( .A1(n1140), .A2(n1153), .ZN(G60) );
NOR2_X1 U826 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U827 ( .A(n1156), .B(KEYINPUT55), .Z(n1155) );
NAND2_X1 U828 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U829 ( .A1(n1157), .A2(n1158), .ZN(n1154) );
NOR2_X1 U830 ( .A1(n1148), .A2(n1159), .ZN(n1157) );
INV_X1 U831 ( .A(G475), .ZN(n1159) );
XOR2_X1 U832 ( .A(G104), .B(n1160), .Z(G6) );
AND2_X1 U833 ( .A1(n1161), .A2(n1075), .ZN(n1160) );
NOR2_X1 U834 ( .A1(n1140), .A2(n1162), .ZN(G57) );
NOR2_X1 U835 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U836 ( .A(n1165), .B(KEYINPUT16), .Z(n1164) );
NAND2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR2_X1 U838 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
XNOR2_X1 U839 ( .A(n1168), .B(n1169), .ZN(n1167) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U841 ( .A(n1172), .B(n1173), .Z(n1168) );
NOR2_X1 U842 ( .A1(n1174), .A2(n1148), .ZN(n1173) );
NOR2_X1 U843 ( .A1(n1140), .A2(n1175), .ZN(G54) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U845 ( .A1(n1106), .A2(n1148), .ZN(n1177) );
NAND3_X1 U846 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1176) );
NAND2_X1 U847 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
INV_X1 U848 ( .A(KEYINPUT2), .ZN(n1182) );
NAND3_X1 U849 ( .A1(KEYINPUT2), .A2(n1183), .A3(n1184), .ZN(n1179) );
OR2_X1 U850 ( .A1(n1184), .A2(n1183), .ZN(n1178) );
NOR2_X1 U851 ( .A1(KEYINPUT23), .A2(n1181), .ZN(n1183) );
NAND2_X1 U852 ( .A1(n1185), .A2(n1186), .ZN(n1181) );
NAND2_X1 U853 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XNOR2_X1 U854 ( .A(KEYINPUT0), .B(n1189), .ZN(n1187) );
NAND2_X1 U855 ( .A1(n1190), .A2(G140), .ZN(n1185) );
XOR2_X1 U856 ( .A(n1189), .B(KEYINPUT3), .Z(n1190) );
XOR2_X1 U857 ( .A(n1191), .B(n1192), .Z(n1184) );
NAND2_X1 U858 ( .A1(n1193), .A2(n1194), .ZN(n1191) );
NAND2_X1 U859 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U860 ( .A(KEYINPUT25), .B(n1197), .Z(n1193) );
NOR2_X1 U861 ( .A1(n1198), .A2(n1196), .ZN(n1197) );
XOR2_X1 U862 ( .A(n1199), .B(n1200), .Z(n1196) );
XNOR2_X1 U863 ( .A(KEYINPUT61), .B(n1195), .ZN(n1198) );
NOR2_X1 U864 ( .A1(n1140), .A2(n1201), .ZN(G51) );
XOR2_X1 U865 ( .A(n1202), .B(n1203), .Z(n1201) );
XOR2_X1 U866 ( .A(n1204), .B(n1205), .Z(n1203) );
NOR2_X1 U867 ( .A1(n1206), .A2(n1148), .ZN(n1205) );
NAND2_X1 U868 ( .A1(G902), .A2(n1207), .ZN(n1148) );
NAND2_X1 U869 ( .A1(n1047), .A2(n1048), .ZN(n1207) );
INV_X1 U870 ( .A(n1139), .ZN(n1048) );
NAND4_X1 U871 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1139) );
AND3_X1 U872 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
NAND2_X1 U873 ( .A1(n1215), .A2(n1216), .ZN(n1210) );
NAND2_X1 U874 ( .A1(n1217), .A2(n1044), .ZN(n1216) );
XNOR2_X1 U875 ( .A(n1075), .B(KEYINPUT17), .ZN(n1217) );
NAND2_X1 U876 ( .A1(n1161), .A2(n1218), .ZN(n1208) );
NAND2_X1 U877 ( .A1(n1219), .A2(n1044), .ZN(n1218) );
XNOR2_X1 U878 ( .A(n1075), .B(KEYINPUT10), .ZN(n1219) );
INV_X1 U879 ( .A(n1043), .ZN(n1161) );
NAND3_X1 U880 ( .A1(n1220), .A2(n1221), .A3(n1089), .ZN(n1043) );
AND4_X1 U881 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1047) );
NOR4_X1 U882 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
NOR2_X1 U883 ( .A1(n1230), .A2(n1231), .ZN(n1224) );
NAND2_X1 U884 ( .A1(n1082), .A2(n1232), .ZN(n1222) );
XOR2_X1 U885 ( .A(KEYINPUT31), .B(n1233), .Z(n1232) );
XNOR2_X1 U886 ( .A(n1234), .B(n1235), .ZN(n1202) );
NOR2_X1 U887 ( .A1(n1236), .A2(G952), .ZN(n1140) );
XNOR2_X1 U888 ( .A(KEYINPUT50), .B(G953), .ZN(n1236) );
XNOR2_X1 U889 ( .A(G146), .B(n1223), .ZN(G48) );
NAND3_X1 U890 ( .A1(n1075), .A2(n1237), .A3(n1238), .ZN(n1223) );
XOR2_X1 U891 ( .A(n1230), .B(n1239), .Z(G45) );
NOR2_X1 U892 ( .A1(KEYINPUT62), .A2(n1240), .ZN(n1239) );
AND4_X1 U893 ( .A1(n1241), .A2(n1078), .A3(n1242), .A4(n1100), .ZN(n1230) );
XNOR2_X1 U894 ( .A(n1188), .B(n1229), .ZN(G42) );
AND3_X1 U895 ( .A1(n1243), .A2(n1237), .A3(n1082), .ZN(n1229) );
XOR2_X1 U896 ( .A(n1228), .B(n1244), .Z(G39) );
NOR2_X1 U897 ( .A1(KEYINPUT51), .A2(n1245), .ZN(n1244) );
AND4_X1 U898 ( .A1(n1058), .A2(n1056), .A3(n1246), .A4(n1055), .ZN(n1228) );
AND3_X1 U899 ( .A1(n1082), .A2(n1237), .A3(n1080), .ZN(n1058) );
XOR2_X1 U900 ( .A(G134), .B(n1227), .Z(G36) );
AND3_X1 U901 ( .A1(n1082), .A2(n1074), .A3(n1241), .ZN(n1227) );
XNOR2_X1 U902 ( .A(G131), .B(n1247), .ZN(G33) );
NAND2_X1 U903 ( .A1(n1233), .A2(n1082), .ZN(n1247) );
NOR2_X1 U904 ( .A1(n1248), .A2(n1069), .ZN(n1082) );
AND2_X1 U905 ( .A1(n1241), .A2(n1075), .ZN(n1233) );
AND3_X1 U906 ( .A1(n1237), .A2(n1246), .A3(n1088), .ZN(n1241) );
XNOR2_X1 U907 ( .A(n1249), .B(n1231), .ZN(G30) );
AND3_X1 U908 ( .A1(n1074), .A2(n1221), .A3(n1238), .ZN(n1231) );
AND4_X1 U909 ( .A1(n1078), .A2(n1056), .A3(n1246), .A4(n1055), .ZN(n1238) );
XNOR2_X1 U910 ( .A(G101), .B(n1209), .ZN(G3) );
NAND4_X1 U911 ( .A1(n1080), .A2(n1088), .A3(n1250), .A4(n1221), .ZN(n1209) );
XNOR2_X1 U912 ( .A(G125), .B(n1251), .ZN(G27) );
NAND2_X1 U913 ( .A1(KEYINPUT34), .A2(n1226), .ZN(n1251) );
AND3_X1 U914 ( .A1(n1243), .A2(n1078), .A3(n1079), .ZN(n1226) );
AND4_X1 U915 ( .A1(n1252), .A2(n1075), .A3(n1246), .A4(n1055), .ZN(n1243) );
NAND2_X1 U916 ( .A1(n1057), .A2(n1253), .ZN(n1246) );
NAND4_X1 U917 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1114), .ZN(n1253) );
INV_X1 U918 ( .A(G900), .ZN(n1114) );
XNOR2_X1 U919 ( .A(G122), .B(n1212), .ZN(G24) );
NAND4_X1 U920 ( .A1(n1079), .A2(n1089), .A3(n1255), .A4(n1220), .ZN(n1212) );
NOR2_X1 U921 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XNOR2_X1 U922 ( .A(G119), .B(n1214), .ZN(G21) );
NAND4_X1 U923 ( .A1(n1080), .A2(n1079), .A3(n1258), .A4(n1250), .ZN(n1214) );
NOR2_X1 U924 ( .A1(n1089), .A2(n1252), .ZN(n1258) );
INV_X1 U925 ( .A(n1055), .ZN(n1089) );
XOR2_X1 U926 ( .A(G116), .B(n1259), .Z(G18) );
NOR2_X1 U927 ( .A1(n1044), .A2(n1260), .ZN(n1259) );
INV_X1 U928 ( .A(n1074), .ZN(n1044) );
NOR2_X1 U929 ( .A1(n1100), .A2(n1257), .ZN(n1074) );
INV_X1 U930 ( .A(n1242), .ZN(n1257) );
XOR2_X1 U931 ( .A(n1261), .B(n1262), .Z(G15) );
NAND2_X1 U932 ( .A1(KEYINPUT40), .A2(G113), .ZN(n1262) );
NAND2_X1 U933 ( .A1(n1215), .A2(n1263), .ZN(n1261) );
XOR2_X1 U934 ( .A(KEYINPUT5), .B(n1075), .Z(n1263) );
NOR2_X1 U935 ( .A1(n1242), .A2(n1256), .ZN(n1075) );
INV_X1 U936 ( .A(n1260), .ZN(n1215) );
NAND3_X1 U937 ( .A1(n1079), .A2(n1250), .A3(n1088), .ZN(n1260) );
NOR2_X1 U938 ( .A1(n1055), .A2(n1252), .ZN(n1088) );
NOR2_X1 U939 ( .A1(n1092), .A2(n1102), .ZN(n1079) );
INV_X1 U940 ( .A(n1091), .ZN(n1102) );
XNOR2_X1 U941 ( .A(G110), .B(n1213), .ZN(G12) );
NAND4_X1 U942 ( .A1(n1080), .A2(n1220), .A3(n1221), .A4(n1055), .ZN(n1213) );
NAND2_X1 U943 ( .A1(n1264), .A2(n1265), .ZN(n1055) );
NAND2_X1 U944 ( .A1(n1103), .A2(n1105), .ZN(n1265) );
XOR2_X1 U945 ( .A(KEYINPUT19), .B(n1266), .Z(n1264) );
NOR2_X1 U946 ( .A1(n1103), .A2(n1105), .ZN(n1266) );
NAND2_X1 U947 ( .A1(n1267), .A2(n1268), .ZN(n1105) );
XNOR2_X1 U948 ( .A(n1145), .B(KEYINPUT58), .ZN(n1267) );
XNOR2_X1 U949 ( .A(n1269), .B(n1270), .ZN(n1145) );
XOR2_X1 U950 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U951 ( .A(n1273), .B(n1274), .Z(n1272) );
NAND2_X1 U952 ( .A1(G221), .A2(n1275), .ZN(n1274) );
INV_X1 U953 ( .A(n1276), .ZN(n1275) );
NAND2_X1 U954 ( .A1(KEYINPUT59), .A2(n1277), .ZN(n1273) );
NOR2_X1 U955 ( .A1(G146), .A2(KEYINPUT20), .ZN(n1271) );
XOR2_X1 U956 ( .A(n1278), .B(n1279), .Z(n1269) );
XNOR2_X1 U957 ( .A(n1188), .B(G125), .ZN(n1279) );
XNOR2_X1 U958 ( .A(n1280), .B(n1281), .ZN(n1278) );
NAND2_X1 U959 ( .A1(n1282), .A2(KEYINPUT41), .ZN(n1280) );
XNOR2_X1 U960 ( .A(G119), .B(G128), .ZN(n1282) );
AND2_X1 U961 ( .A1(G217), .A2(n1283), .ZN(n1103) );
XOR2_X1 U962 ( .A(n1237), .B(KEYINPUT57), .Z(n1221) );
AND2_X1 U963 ( .A1(n1092), .A2(n1091), .ZN(n1237) );
NAND2_X1 U964 ( .A1(G221), .A2(n1283), .ZN(n1091) );
NAND2_X1 U965 ( .A1(G234), .A2(n1268), .ZN(n1283) );
XNOR2_X1 U966 ( .A(n1108), .B(n1106), .ZN(n1092) );
INV_X1 U967 ( .A(G469), .ZN(n1106) );
AND2_X1 U968 ( .A1(n1284), .A2(n1268), .ZN(n1108) );
XOR2_X1 U969 ( .A(n1123), .B(n1285), .Z(n1284) );
XOR2_X1 U970 ( .A(n1189), .B(n1195), .Z(n1285) );
XNOR2_X1 U971 ( .A(G110), .B(n1286), .ZN(n1189) );
NOR2_X1 U972 ( .A1(G953), .A2(n1113), .ZN(n1286) );
INV_X1 U973 ( .A(G227), .ZN(n1113) );
XNOR2_X1 U974 ( .A(n1287), .B(n1199), .ZN(n1123) );
NAND2_X1 U975 ( .A1(n1288), .A2(n1289), .ZN(n1199) );
NAND2_X1 U976 ( .A1(KEYINPUT39), .A2(G143), .ZN(n1289) );
OR2_X1 U977 ( .A1(KEYINPUT45), .A2(G143), .ZN(n1288) );
XNOR2_X1 U978 ( .A(n1172), .B(n1188), .ZN(n1287) );
INV_X1 U979 ( .A(G140), .ZN(n1188) );
XNOR2_X1 U980 ( .A(n1290), .B(n1200), .ZN(n1172) );
AND2_X1 U981 ( .A1(n1250), .A2(n1252), .ZN(n1220) );
INV_X1 U982 ( .A(n1056), .ZN(n1252) );
XOR2_X1 U983 ( .A(n1291), .B(n1174), .Z(n1056) );
INV_X1 U984 ( .A(G472), .ZN(n1174) );
NAND2_X1 U985 ( .A1(n1292), .A2(n1268), .ZN(n1291) );
XOR2_X1 U986 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U987 ( .A(n1171), .B(n1166), .Z(n1294) );
AND2_X1 U988 ( .A1(n1295), .A2(n1296), .ZN(n1166) );
NAND2_X1 U989 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
INV_X1 U990 ( .A(G101), .ZN(n1298) );
NAND2_X1 U991 ( .A1(G210), .A2(n1299), .ZN(n1297) );
NAND3_X1 U992 ( .A1(G210), .A2(n1299), .A3(G101), .ZN(n1295) );
XOR2_X1 U993 ( .A(n1300), .B(KEYINPUT27), .Z(n1293) );
NAND3_X1 U994 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1300) );
NAND2_X1 U995 ( .A1(KEYINPUT47), .A2(n1290), .ZN(n1303) );
OR3_X1 U996 ( .A1(n1304), .A2(KEYINPUT47), .A3(n1305), .ZN(n1302) );
NAND2_X1 U997 ( .A1(n1305), .A2(n1304), .ZN(n1301) );
NAND2_X1 U998 ( .A1(KEYINPUT4), .A2(n1192), .ZN(n1304) );
INV_X1 U999 ( .A(n1290), .ZN(n1192) );
XOR2_X1 U1000 ( .A(n1306), .B(n1307), .Z(n1290) );
XNOR2_X1 U1001 ( .A(G131), .B(n1277), .ZN(n1306) );
XNOR2_X1 U1002 ( .A(n1245), .B(KEYINPUT7), .ZN(n1277) );
INV_X1 U1003 ( .A(G137), .ZN(n1245) );
AND2_X1 U1004 ( .A1(n1078), .A2(n1308), .ZN(n1250) );
NAND2_X1 U1005 ( .A1(n1057), .A2(n1309), .ZN(n1308) );
NAND4_X1 U1006 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1130), .ZN(n1309) );
INV_X1 U1007 ( .A(G898), .ZN(n1130) );
NAND3_X1 U1008 ( .A1(n1254), .A2(n1112), .A3(G952), .ZN(n1057) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1254) );
INV_X1 U1010 ( .A(n1068), .ZN(n1078) );
NAND2_X1 U1011 ( .A1(n1069), .A2(n1310), .ZN(n1068) );
INV_X1 U1012 ( .A(n1248), .ZN(n1310) );
XNOR2_X1 U1013 ( .A(n1071), .B(KEYINPUT28), .ZN(n1248) );
AND2_X1 U1014 ( .A1(G214), .A2(n1311), .ZN(n1071) );
XNOR2_X1 U1015 ( .A(n1099), .B(KEYINPUT53), .ZN(n1069) );
XOR2_X1 U1016 ( .A(n1312), .B(n1206), .Z(n1099) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1311), .ZN(n1206) );
NAND2_X1 U1018 ( .A1(n1313), .A2(n1268), .ZN(n1311) );
INV_X1 U1019 ( .A(G237), .ZN(n1313) );
NAND2_X1 U1020 ( .A1(n1314), .A2(n1268), .ZN(n1312) );
XNOR2_X1 U1021 ( .A(n1315), .B(n1135), .ZN(n1314) );
INV_X1 U1022 ( .A(n1234), .ZN(n1135) );
XNOR2_X1 U1023 ( .A(n1316), .B(n1317), .ZN(n1234) );
XNOR2_X1 U1024 ( .A(n1281), .B(n1318), .ZN(n1317) );
NOR2_X1 U1025 ( .A1(KEYINPUT6), .A2(n1319), .ZN(n1318) );
INV_X1 U1026 ( .A(G110), .ZN(n1281) );
XOR2_X1 U1027 ( .A(n1195), .B(n1171), .Z(n1316) );
XOR2_X1 U1028 ( .A(n1320), .B(n1321), .Z(n1171) );
XNOR2_X1 U1029 ( .A(G113), .B(G119), .ZN(n1320) );
XNOR2_X1 U1030 ( .A(G101), .B(n1322), .ZN(n1195) );
XNOR2_X1 U1031 ( .A(n1041), .B(G104), .ZN(n1322) );
NAND2_X1 U1032 ( .A1(n1323), .A2(n1324), .ZN(n1315) );
NAND2_X1 U1033 ( .A1(n1235), .A2(n1325), .ZN(n1324) );
NAND2_X1 U1034 ( .A1(KEYINPUT60), .A2(G224), .ZN(n1325) );
INV_X1 U1035 ( .A(n1326), .ZN(n1235) );
NAND3_X1 U1036 ( .A1(KEYINPUT60), .A2(n1204), .A3(n1326), .ZN(n1323) );
XOR2_X1 U1037 ( .A(n1305), .B(n1124), .Z(n1326) );
XOR2_X1 U1038 ( .A(n1200), .B(n1170), .Z(n1305) );
XNOR2_X1 U1039 ( .A(n1327), .B(G143), .ZN(n1170) );
XNOR2_X1 U1040 ( .A(KEYINPUT33), .B(KEYINPUT21), .ZN(n1327) );
XOR2_X1 U1041 ( .A(G128), .B(G146), .Z(n1200) );
NOR2_X1 U1042 ( .A1(n1129), .A2(G953), .ZN(n1204) );
INV_X1 U1043 ( .A(G224), .ZN(n1129) );
NOR2_X1 U1044 ( .A1(n1242), .A2(n1100), .ZN(n1080) );
INV_X1 U1045 ( .A(n1256), .ZN(n1100) );
XOR2_X1 U1046 ( .A(n1328), .B(G475), .Z(n1256) );
OR2_X1 U1047 ( .A1(n1158), .A2(G902), .ZN(n1328) );
XOR2_X1 U1048 ( .A(n1329), .B(n1330), .Z(n1158) );
XOR2_X1 U1049 ( .A(G113), .B(n1331), .Z(n1330) );
XNOR2_X1 U1050 ( .A(G146), .B(n1319), .ZN(n1331) );
XOR2_X1 U1051 ( .A(n1332), .B(n1333), .Z(n1329) );
XNOR2_X1 U1052 ( .A(G104), .B(n1334), .ZN(n1333) );
NAND2_X1 U1053 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND2_X1 U1054 ( .A1(G140), .A2(n1124), .ZN(n1336) );
XOR2_X1 U1055 ( .A(KEYINPUT56), .B(n1337), .Z(n1335) );
NOR2_X1 U1056 ( .A1(G140), .A2(n1124), .ZN(n1337) );
INV_X1 U1057 ( .A(G125), .ZN(n1124) );
NAND2_X1 U1058 ( .A1(n1338), .A2(n1339), .ZN(n1332) );
OR2_X1 U1059 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1060 ( .A(n1342), .B(KEYINPUT14), .Z(n1338) );
NAND2_X1 U1061 ( .A1(n1341), .A2(n1340), .ZN(n1342) );
INV_X1 U1062 ( .A(G131), .ZN(n1340) );
XOR2_X1 U1063 ( .A(n1343), .B(n1240), .Z(n1341) );
INV_X1 U1064 ( .A(G143), .ZN(n1240) );
NAND2_X1 U1065 ( .A1(G214), .A2(n1299), .ZN(n1343) );
NOR2_X1 U1066 ( .A1(G953), .A2(G237), .ZN(n1299) );
XNOR2_X1 U1067 ( .A(n1101), .B(KEYINPUT63), .ZN(n1242) );
XNOR2_X1 U1068 ( .A(n1344), .B(n1152), .ZN(n1101) );
INV_X1 U1069 ( .A(G478), .ZN(n1152) );
NAND2_X1 U1070 ( .A1(n1150), .A2(n1268), .ZN(n1344) );
INV_X1 U1071 ( .A(G902), .ZN(n1268) );
XNOR2_X1 U1072 ( .A(n1345), .B(n1346), .ZN(n1150) );
NOR2_X1 U1073 ( .A1(n1276), .A2(n1147), .ZN(n1346) );
INV_X1 U1074 ( .A(G217), .ZN(n1147) );
NAND2_X1 U1075 ( .A1(G234), .A2(n1112), .ZN(n1276) );
INV_X1 U1076 ( .A(G953), .ZN(n1112) );
NAND3_X1 U1077 ( .A1(n1347), .A2(n1348), .A3(KEYINPUT24), .ZN(n1345) );
NAND2_X1 U1078 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1079 ( .A1(KEYINPUT48), .A2(n1307), .ZN(n1350) );
XOR2_X1 U1080 ( .A(n1351), .B(n1352), .Z(n1349) );
NAND2_X1 U1081 ( .A1(KEYINPUT37), .A2(n1353), .ZN(n1352) );
NAND3_X1 U1082 ( .A1(n1307), .A2(n1354), .A3(KEYINPUT48), .ZN(n1347) );
XOR2_X1 U1083 ( .A(n1351), .B(n1355), .Z(n1354) );
NAND2_X1 U1084 ( .A1(n1356), .A2(KEYINPUT37), .ZN(n1355) );
INV_X1 U1085 ( .A(n1353), .ZN(n1356) );
NAND2_X1 U1086 ( .A1(n1357), .A2(n1358), .ZN(n1353) );
NAND2_X1 U1087 ( .A1(n1359), .A2(n1249), .ZN(n1358) );
XOR2_X1 U1088 ( .A(n1360), .B(KEYINPUT35), .Z(n1357) );
OR2_X1 U1089 ( .A1(n1249), .A2(n1359), .ZN(n1360) );
XOR2_X1 U1090 ( .A(G143), .B(KEYINPUT15), .Z(n1359) );
INV_X1 U1091 ( .A(G128), .ZN(n1249) );
NAND3_X1 U1092 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1351) );
NAND2_X1 U1093 ( .A1(n1364), .A2(n1041), .ZN(n1363) );
NAND2_X1 U1094 ( .A1(n1365), .A2(n1366), .ZN(n1362) );
INV_X1 U1095 ( .A(KEYINPUT43), .ZN(n1366) );
NAND2_X1 U1096 ( .A1(n1367), .A2(n1368), .ZN(n1365) );
XNOR2_X1 U1097 ( .A(KEYINPUT49), .B(n1041), .ZN(n1368) );
INV_X1 U1098 ( .A(n1364), .ZN(n1367) );
NAND2_X1 U1099 ( .A1(KEYINPUT43), .A2(n1369), .ZN(n1361) );
NAND2_X1 U1100 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
OR3_X1 U1101 ( .A1(n1041), .A2(n1364), .A3(KEYINPUT49), .ZN(n1371) );
XOR2_X1 U1102 ( .A(n1372), .B(n1319), .Z(n1364) );
INV_X1 U1103 ( .A(G122), .ZN(n1319) );
NAND2_X1 U1104 ( .A1(KEYINPUT44), .A2(n1321), .ZN(n1372) );
XNOR2_X1 U1105 ( .A(G116), .B(KEYINPUT9), .ZN(n1321) );
NAND2_X1 U1106 ( .A1(KEYINPUT49), .A2(n1041), .ZN(n1370) );
INV_X1 U1107 ( .A(G107), .ZN(n1041) );
XNOR2_X1 U1108 ( .A(G134), .B(KEYINPUT1), .ZN(n1307) );
endmodule


