//Key = 1101100110111011011100010010111110111000001000100010110111101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;

XOR2_X1 U719 ( .A(G107), .B(n998), .Z(G9) );
NOR2_X1 U720 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR3_X1 U721 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n1000) );
NOR2_X1 U722 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NOR2_X1 U723 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR4_X1 U724 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1007) );
NOR2_X1 U725 ( .A1(n1012), .A2(n1013), .ZN(n1009) );
NOR2_X1 U726 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR2_X1 U727 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U728 ( .A1(n1018), .A2(n1019), .ZN(n1014) );
NOR2_X1 U729 ( .A1(n1020), .A2(n1021), .ZN(n1008) );
AND2_X1 U730 ( .A1(n1018), .A2(n1022), .ZN(n1020) );
NOR4_X1 U731 ( .A1(n1023), .A2(n1012), .A3(n1024), .A4(n1017), .ZN(n1006) );
NOR3_X1 U732 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1023) );
NOR2_X1 U733 ( .A1(n1028), .A2(n1010), .ZN(n1027) );
NOR2_X1 U734 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NOR2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U736 ( .A1(n1033), .A2(n1034), .ZN(n1026) );
XNOR2_X1 U737 ( .A(n1035), .B(KEYINPUT59), .ZN(n1033) );
NOR2_X1 U738 ( .A1(n1036), .A2(n1011), .ZN(n1025) );
NAND3_X1 U739 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1001) );
NAND4_X1 U740 ( .A1(n1040), .A2(n1035), .A3(n1041), .A4(n1042), .ZN(n1039) );
NOR4_X1 U741 ( .A1(n1010), .A2(n1012), .A3(n1005), .A4(n1017), .ZN(n1042) );
XNOR2_X1 U742 ( .A(n1043), .B(n1044), .ZN(n1041) );
XNOR2_X1 U743 ( .A(KEYINPUT35), .B(KEYINPUT21), .ZN(n1043) );
NOR3_X1 U744 ( .A1(n1045), .A2(G953), .A3(G952), .ZN(n999) );
INV_X1 U745 ( .A(n1037), .ZN(n1045) );
NAND4_X1 U746 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1037) );
NOR4_X1 U747 ( .A1(n1050), .A2(n1012), .A3(n1051), .A4(n1052), .ZN(n1049) );
XOR2_X1 U748 ( .A(KEYINPUT20), .B(n1053), .Z(n1052) );
XNOR2_X1 U749 ( .A(G478), .B(n1054), .ZN(n1051) );
NOR3_X1 U750 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1048) );
NAND2_X1 U751 ( .A1(n1058), .A2(n1059), .ZN(n1047) );
XNOR2_X1 U752 ( .A(G469), .B(KEYINPUT12), .ZN(n1058) );
XOR2_X1 U753 ( .A(n1060), .B(n1061), .Z(n1046) );
NAND2_X1 U754 ( .A1(KEYINPUT28), .A2(n1062), .ZN(n1061) );
XOR2_X1 U755 ( .A(n1063), .B(n1064), .Z(G72) );
XOR2_X1 U756 ( .A(n1065), .B(n1066), .Z(n1064) );
NAND2_X1 U757 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U758 ( .A1(G900), .A2(G227), .ZN(n1068) );
NAND2_X1 U759 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NAND2_X1 U760 ( .A1(G953), .A2(n1071), .ZN(n1070) );
XOR2_X1 U761 ( .A(n1072), .B(n1073), .Z(n1069) );
XOR2_X1 U762 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U763 ( .A1(KEYINPUT4), .A2(n1076), .ZN(n1075) );
NAND2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
XOR2_X1 U765 ( .A(KEYINPUT30), .B(KEYINPUT25), .Z(n1078) );
NOR2_X1 U766 ( .A1(n1079), .A2(G953), .ZN(n1063) );
NOR2_X1 U767 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U768 ( .A(n1082), .B(n1083), .Z(G69) );
XOR2_X1 U769 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR2_X1 U770 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U771 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U772 ( .A1(n1090), .A2(KEYINPUT31), .ZN(n1088) );
XOR2_X1 U773 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U774 ( .A1(KEYINPUT3), .A2(n1093), .ZN(n1091) );
NAND2_X1 U775 ( .A1(n1067), .A2(n1094), .ZN(n1084) );
NAND2_X1 U776 ( .A1(G898), .A2(G224), .ZN(n1094) );
XNOR2_X1 U777 ( .A(G953), .B(KEYINPUT18), .ZN(n1067) );
NAND2_X1 U778 ( .A1(n1095), .A2(n1096), .ZN(n1082) );
NAND2_X1 U779 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XNOR2_X1 U780 ( .A(n1099), .B(KEYINPUT42), .ZN(n1097) );
XNOR2_X1 U781 ( .A(G953), .B(KEYINPUT45), .ZN(n1095) );
NOR2_X1 U782 ( .A1(n1100), .A2(n1101), .ZN(G66) );
XNOR2_X1 U783 ( .A(n1102), .B(n1103), .ZN(n1101) );
NOR2_X1 U784 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U785 ( .A1(n1100), .A2(n1106), .ZN(G63) );
XNOR2_X1 U786 ( .A(n1107), .B(n1108), .ZN(n1106) );
NOR2_X1 U787 ( .A1(n1109), .A2(n1105), .ZN(n1107) );
INV_X1 U788 ( .A(G478), .ZN(n1109) );
NOR2_X1 U789 ( .A1(n1100), .A2(n1110), .ZN(G60) );
XOR2_X1 U790 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U791 ( .A1(n1113), .A2(n1105), .ZN(n1111) );
XOR2_X1 U792 ( .A(G104), .B(n1114), .Z(G6) );
NOR2_X1 U793 ( .A1(n1100), .A2(n1115), .ZN(G57) );
XOR2_X1 U794 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U797 ( .A1(n1062), .A2(n1105), .ZN(n1120) );
NOR3_X1 U798 ( .A1(n1122), .A2(n1062), .A3(n1105), .ZN(n1118) );
XOR2_X1 U799 ( .A(KEYINPUT52), .B(n1121), .Z(n1122) );
XNOR2_X1 U800 ( .A(n1123), .B(n1124), .ZN(n1121) );
NAND2_X1 U801 ( .A1(KEYINPUT50), .A2(n1125), .ZN(n1116) );
NOR2_X1 U802 ( .A1(n1100), .A2(n1126), .ZN(G54) );
XOR2_X1 U803 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U804 ( .A(KEYINPUT32), .B(n1129), .Z(n1128) );
NOR2_X1 U805 ( .A1(n1105), .A2(n1130), .ZN(n1129) );
XOR2_X1 U806 ( .A(KEYINPUT58), .B(G469), .Z(n1130) );
NOR2_X1 U807 ( .A1(n1100), .A2(n1131), .ZN(G51) );
XOR2_X1 U808 ( .A(n1132), .B(n1133), .Z(n1131) );
XNOR2_X1 U809 ( .A(n1134), .B(n1135), .ZN(n1133) );
XOR2_X1 U810 ( .A(n1136), .B(n1137), .Z(n1132) );
NOR2_X1 U811 ( .A1(n1138), .A2(KEYINPUT39), .ZN(n1137) );
XNOR2_X1 U812 ( .A(G125), .B(n1139), .ZN(n1136) );
NOR2_X1 U813 ( .A1(n1140), .A2(n1105), .ZN(n1139) );
NAND2_X1 U814 ( .A1(G902), .A2(n1003), .ZN(n1105) );
NAND4_X1 U815 ( .A1(n1099), .A2(n1098), .A3(n1141), .A4(n1142), .ZN(n1003) );
XOR2_X1 U816 ( .A(KEYINPUT36), .B(n1080), .Z(n1142) );
INV_X1 U817 ( .A(n1081), .ZN(n1141) );
NAND4_X1 U818 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1081) );
NOR2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
INV_X1 U820 ( .A(n1149), .ZN(n1147) );
NAND3_X1 U821 ( .A1(n1035), .A2(n1150), .A3(n1151), .ZN(n1144) );
NAND2_X1 U822 ( .A1(n1036), .A2(n1034), .ZN(n1150) );
NAND2_X1 U823 ( .A1(n1030), .A2(n1152), .ZN(n1143) );
NAND2_X1 U824 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U825 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U826 ( .A1(n1034), .A2(n1157), .ZN(n1156) );
NAND2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
INV_X1 U828 ( .A(n1160), .ZN(n1155) );
OR2_X1 U829 ( .A1(n1159), .A2(n1161), .ZN(n1153) );
INV_X1 U830 ( .A(KEYINPUT24), .ZN(n1159) );
NOR4_X1 U831 ( .A1(n1162), .A2(n1114), .A3(n1163), .A4(n998), .ZN(n1098) );
AND3_X1 U832 ( .A1(n1164), .A2(n1165), .A3(n1016), .ZN(n998) );
AND3_X1 U833 ( .A1(n1016), .A2(n1164), .A3(n1158), .ZN(n1114) );
AND4_X1 U834 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1099) );
NAND2_X1 U835 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
XNOR2_X1 U836 ( .A(KEYINPUT37), .B(n1024), .ZN(n1171) );
NOR2_X1 U837 ( .A1(n1038), .A2(G952), .ZN(n1100) );
XNOR2_X1 U838 ( .A(G146), .B(n1172), .ZN(G48) );
NAND2_X1 U839 ( .A1(n1161), .A2(n1030), .ZN(n1172) );
NOR2_X1 U840 ( .A1(n1160), .A2(n1036), .ZN(n1161) );
INV_X1 U841 ( .A(n1158), .ZN(n1036) );
XNOR2_X1 U842 ( .A(G143), .B(n1146), .ZN(G45) );
NAND4_X1 U843 ( .A1(n1173), .A2(n1151), .A3(n1030), .A4(n1050), .ZN(n1146) );
XOR2_X1 U844 ( .A(G140), .B(n1148), .Z(G42) );
AND3_X1 U845 ( .A1(n1035), .A2(n1016), .A3(n1174), .ZN(n1148) );
XOR2_X1 U846 ( .A(G137), .B(n1080), .Z(G39) );
NOR3_X1 U847 ( .A1(n1011), .A2(n1010), .A3(n1160), .ZN(n1080) );
INV_X1 U848 ( .A(n1175), .ZN(n1010) );
XOR2_X1 U849 ( .A(G134), .B(n1176), .Z(G36) );
NOR4_X1 U850 ( .A1(KEYINPUT13), .A2(n1034), .A3(n1011), .A4(n1177), .ZN(n1176) );
NAND3_X1 U851 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(G33) );
NAND2_X1 U852 ( .A1(G131), .A2(n1181), .ZN(n1180) );
NAND2_X1 U853 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
INV_X1 U854 ( .A(KEYINPUT23), .ZN(n1183) );
NAND2_X1 U855 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
XNOR2_X1 U856 ( .A(KEYINPUT0), .B(n1186), .ZN(n1185) );
NAND2_X1 U857 ( .A1(KEYINPUT23), .A2(n1187), .ZN(n1178) );
NAND2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NAND3_X1 U859 ( .A1(KEYINPUT0), .A2(n1184), .A3(n1186), .ZN(n1189) );
INV_X1 U860 ( .A(n1181), .ZN(n1184) );
NAND3_X1 U861 ( .A1(n1158), .A2(n1190), .A3(n1151), .ZN(n1181) );
INV_X1 U862 ( .A(n1177), .ZN(n1151) );
NAND4_X1 U863 ( .A1(n1021), .A2(n1016), .A3(n1017), .A4(n1191), .ZN(n1177) );
XNOR2_X1 U864 ( .A(KEYINPUT40), .B(n1011), .ZN(n1190) );
INV_X1 U865 ( .A(n1035), .ZN(n1011) );
NOR2_X1 U866 ( .A1(n1031), .A2(n1055), .ZN(n1035) );
INV_X1 U867 ( .A(n1032), .ZN(n1055) );
OR2_X1 U868 ( .A1(n1186), .A2(KEYINPUT0), .ZN(n1188) );
XNOR2_X1 U869 ( .A(n1192), .B(n1193), .ZN(G30) );
NOR4_X1 U870 ( .A1(KEYINPUT16), .A2(n1194), .A3(n1034), .A4(n1160), .ZN(n1193) );
NAND4_X1 U871 ( .A1(n1016), .A2(n1017), .A3(n1012), .A4(n1191), .ZN(n1160) );
XNOR2_X1 U872 ( .A(n1195), .B(n1163), .ZN(G3) );
AND3_X1 U873 ( .A1(n1016), .A2(n1175), .A3(n1196), .ZN(n1163) );
XNOR2_X1 U874 ( .A(n1197), .B(n1198), .ZN(G27) );
NAND2_X1 U875 ( .A1(KEYINPUT1), .A2(n1149), .ZN(n1197) );
NAND3_X1 U876 ( .A1(n1018), .A2(n1030), .A3(n1174), .ZN(n1149) );
AND4_X1 U877 ( .A1(n1022), .A2(n1158), .A3(n1012), .A4(n1191), .ZN(n1174) );
NAND2_X1 U878 ( .A1(n1005), .A2(n1199), .ZN(n1191) );
NAND4_X1 U879 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1071), .ZN(n1199) );
INV_X1 U880 ( .A(G900), .ZN(n1071) );
XNOR2_X1 U881 ( .A(KEYINPUT63), .B(n1201), .ZN(n1200) );
XNOR2_X1 U882 ( .A(G122), .B(n1202), .ZN(G24) );
NAND2_X1 U883 ( .A1(n1170), .A2(n1018), .ZN(n1202) );
AND3_X1 U884 ( .A1(n1173), .A2(n1050), .A3(n1164), .ZN(n1170) );
AND2_X1 U885 ( .A1(n1203), .A2(n1019), .ZN(n1164) );
XOR2_X1 U886 ( .A(G119), .B(n1204), .Z(G21) );
NOR2_X1 U887 ( .A1(KEYINPUT27), .A2(n1167), .ZN(n1204) );
NAND4_X1 U888 ( .A1(n1030), .A2(n1175), .A3(n1018), .A4(n1205), .ZN(n1167) );
NOR3_X1 U889 ( .A1(n1019), .A2(n1206), .A3(n1021), .ZN(n1205) );
INV_X1 U890 ( .A(n1017), .ZN(n1019) );
XNOR2_X1 U891 ( .A(G116), .B(n1168), .ZN(G18) );
NAND3_X1 U892 ( .A1(n1018), .A2(n1165), .A3(n1196), .ZN(n1168) );
INV_X1 U893 ( .A(n1034), .ZN(n1165) );
NAND2_X1 U894 ( .A1(n1207), .A2(n1173), .ZN(n1034) );
XNOR2_X1 U895 ( .A(KEYINPUT54), .B(n1050), .ZN(n1207) );
NAND2_X1 U896 ( .A1(n1208), .A2(n1209), .ZN(G15) );
NAND2_X1 U897 ( .A1(G113), .A2(n1169), .ZN(n1209) );
XOR2_X1 U898 ( .A(n1210), .B(KEYINPUT41), .Z(n1208) );
OR2_X1 U899 ( .A1(n1169), .A2(G113), .ZN(n1210) );
NAND3_X1 U900 ( .A1(n1018), .A2(n1158), .A3(n1196), .ZN(n1169) );
AND2_X1 U901 ( .A1(n1203), .A2(n1017), .ZN(n1196) );
NOR3_X1 U902 ( .A1(n1012), .A2(n1206), .A3(n1194), .ZN(n1203) );
INV_X1 U903 ( .A(n1024), .ZN(n1018) );
NAND2_X1 U904 ( .A1(n1040), .A2(n1044), .ZN(n1024) );
XNOR2_X1 U905 ( .A(n1211), .B(n1212), .ZN(G12) );
NAND3_X1 U906 ( .A1(n1213), .A2(n1214), .A3(KEYINPUT11), .ZN(n1211) );
NAND2_X1 U907 ( .A1(n1162), .A2(n1215), .ZN(n1214) );
INV_X1 U908 ( .A(KEYINPUT5), .ZN(n1215) );
NOR2_X1 U909 ( .A1(n1216), .A2(n1194), .ZN(n1162) );
NAND3_X1 U910 ( .A1(n1030), .A2(n1216), .A3(KEYINPUT5), .ZN(n1213) );
NAND4_X1 U911 ( .A1(n1022), .A2(n1016), .A3(n1217), .A4(n1175), .ZN(n1216) );
NAND2_X1 U912 ( .A1(n1218), .A2(n1219), .ZN(n1175) );
OR3_X1 U913 ( .A1(n1173), .A2(n1050), .A3(KEYINPUT54), .ZN(n1219) );
NAND2_X1 U914 ( .A1(KEYINPUT54), .A2(n1158), .ZN(n1218) );
NOR2_X1 U915 ( .A1(n1220), .A2(n1173), .ZN(n1158) );
XOR2_X1 U916 ( .A(n1221), .B(G478), .Z(n1173) );
NAND2_X1 U917 ( .A1(KEYINPUT29), .A2(n1054), .ZN(n1221) );
NAND2_X1 U918 ( .A1(n1108), .A2(n1222), .ZN(n1054) );
XNOR2_X1 U919 ( .A(KEYINPUT61), .B(n1223), .ZN(n1222) );
XOR2_X1 U920 ( .A(n1224), .B(n1225), .Z(n1108) );
XOR2_X1 U921 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U922 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
INV_X1 U923 ( .A(G217), .ZN(n1228) );
NOR2_X1 U924 ( .A1(G134), .A2(KEYINPUT47), .ZN(n1226) );
XOR2_X1 U925 ( .A(n1230), .B(n1231), .Z(n1224) );
XNOR2_X1 U926 ( .A(G143), .B(n1192), .ZN(n1231) );
NAND2_X1 U927 ( .A1(n1232), .A2(n1233), .ZN(n1230) );
OR2_X1 U928 ( .A1(n1234), .A2(G107), .ZN(n1233) );
XOR2_X1 U929 ( .A(n1235), .B(KEYINPUT22), .Z(n1232) );
NAND2_X1 U930 ( .A1(G107), .A2(n1234), .ZN(n1235) );
XOR2_X1 U931 ( .A(G116), .B(G122), .Z(n1234) );
INV_X1 U932 ( .A(n1050), .ZN(n1220) );
XOR2_X1 U933 ( .A(n1236), .B(n1113), .Z(n1050) );
INV_X1 U934 ( .A(G475), .ZN(n1113) );
OR2_X1 U935 ( .A1(n1112), .A2(G902), .ZN(n1236) );
XNOR2_X1 U936 ( .A(n1237), .B(n1238), .ZN(n1112) );
XOR2_X1 U937 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U938 ( .A(G122), .B(G104), .Z(n1240) );
XNOR2_X1 U939 ( .A(G143), .B(n1186), .ZN(n1239) );
INV_X1 U940 ( .A(G131), .ZN(n1186) );
XOR2_X1 U941 ( .A(n1241), .B(n1242), .Z(n1237) );
AND2_X1 U942 ( .A1(G214), .A2(n1243), .ZN(n1242) );
XOR2_X1 U943 ( .A(n1244), .B(n1245), .Z(n1241) );
NOR2_X1 U944 ( .A1(KEYINPUT2), .A2(G113), .ZN(n1245) );
NAND2_X1 U945 ( .A1(n1246), .A2(n1247), .ZN(n1244) );
NAND2_X1 U946 ( .A1(G146), .A2(n1248), .ZN(n1247) );
XOR2_X1 U947 ( .A(KEYINPUT55), .B(n1249), .Z(n1246) );
NOR2_X1 U948 ( .A1(G146), .A2(n1248), .ZN(n1249) );
INV_X1 U949 ( .A(n1076), .ZN(n1248) );
XOR2_X1 U950 ( .A(G140), .B(n1198), .Z(n1076) );
NOR2_X1 U951 ( .A1(n1206), .A2(n1021), .ZN(n1217) );
INV_X1 U952 ( .A(n1012), .ZN(n1021) );
XOR2_X1 U953 ( .A(n1250), .B(n1104), .Z(n1012) );
NAND2_X1 U954 ( .A1(G217), .A2(n1251), .ZN(n1104) );
NAND2_X1 U955 ( .A1(n1102), .A2(n1223), .ZN(n1250) );
XNOR2_X1 U956 ( .A(n1252), .B(n1253), .ZN(n1102) );
XOR2_X1 U957 ( .A(n1254), .B(n1255), .Z(n1253) );
NOR2_X1 U958 ( .A1(G125), .A2(KEYINPUT49), .ZN(n1254) );
XOR2_X1 U959 ( .A(n1256), .B(n1257), .Z(n1252) );
NOR2_X1 U960 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U961 ( .A(n1260), .B(KEYINPUT34), .Z(n1259) );
NAND2_X1 U962 ( .A1(G119), .A2(n1192), .ZN(n1260) );
NOR2_X1 U963 ( .A1(G119), .A2(n1192), .ZN(n1258) );
INV_X1 U964 ( .A(G128), .ZN(n1192) );
XNOR2_X1 U965 ( .A(n1261), .B(n1262), .ZN(n1256) );
NOR2_X1 U966 ( .A1(KEYINPUT33), .A2(n1263), .ZN(n1262) );
XOR2_X1 U967 ( .A(KEYINPUT7), .B(G146), .Z(n1263) );
NOR2_X1 U968 ( .A1(KEYINPUT43), .A2(n1264), .ZN(n1261) );
XNOR2_X1 U969 ( .A(G137), .B(n1265), .ZN(n1264) );
NOR2_X1 U970 ( .A1(n1266), .A2(n1229), .ZN(n1265) );
NAND2_X1 U971 ( .A1(G234), .A2(n1267), .ZN(n1229) );
INV_X1 U972 ( .A(G221), .ZN(n1266) );
AND2_X1 U973 ( .A1(n1005), .A2(n1268), .ZN(n1206) );
NAND3_X1 U974 ( .A1(n1086), .A2(n1201), .A3(G902), .ZN(n1268) );
AND2_X1 U975 ( .A1(n1269), .A2(G953), .ZN(n1086) );
XNOR2_X1 U976 ( .A(G898), .B(KEYINPUT48), .ZN(n1269) );
NAND3_X1 U977 ( .A1(n1201), .A2(n1038), .A3(G952), .ZN(n1005) );
NAND2_X1 U978 ( .A1(G237), .A2(G234), .ZN(n1201) );
NOR2_X1 U979 ( .A1(n1056), .A2(n1040), .ZN(n1016) );
NOR2_X1 U980 ( .A1(n1270), .A2(n1057), .ZN(n1040) );
NOR2_X1 U981 ( .A1(n1059), .A2(G469), .ZN(n1057) );
AND2_X1 U982 ( .A1(G469), .A2(n1059), .ZN(n1270) );
NAND2_X1 U983 ( .A1(n1271), .A2(n1223), .ZN(n1059) );
XNOR2_X1 U984 ( .A(n1127), .B(KEYINPUT19), .ZN(n1271) );
XNOR2_X1 U985 ( .A(n1272), .B(n1273), .ZN(n1127) );
XOR2_X1 U986 ( .A(n1072), .B(n1274), .Z(n1273) );
XOR2_X1 U987 ( .A(n1275), .B(n1255), .Z(n1274) );
XNOR2_X1 U988 ( .A(n1212), .B(G140), .ZN(n1255) );
INV_X1 U989 ( .A(G110), .ZN(n1212) );
XOR2_X1 U990 ( .A(n1276), .B(n1277), .Z(n1072) );
NAND2_X1 U991 ( .A1(KEYINPUT57), .A2(G128), .ZN(n1276) );
XNOR2_X1 U992 ( .A(n1278), .B(n1077), .ZN(n1272) );
XNOR2_X1 U993 ( .A(n1279), .B(n1195), .ZN(n1278) );
NAND2_X1 U994 ( .A1(G227), .A2(n1267), .ZN(n1279) );
INV_X1 U995 ( .A(n1044), .ZN(n1056) );
NAND2_X1 U996 ( .A1(G221), .A2(n1251), .ZN(n1044) );
NAND2_X1 U997 ( .A1(G234), .A2(n1223), .ZN(n1251) );
XNOR2_X1 U998 ( .A(n1017), .B(KEYINPUT9), .ZN(n1022) );
XOR2_X1 U999 ( .A(n1060), .B(n1062), .Z(n1017) );
INV_X1 U1000 ( .A(G472), .ZN(n1062) );
NAND2_X1 U1001 ( .A1(n1280), .A2(n1223), .ZN(n1060) );
XOR2_X1 U1002 ( .A(n1281), .B(n1125), .Z(n1280) );
AND2_X1 U1003 ( .A1(n1282), .A2(n1283), .ZN(n1125) );
NAND2_X1 U1004 ( .A1(n1284), .A2(n1195), .ZN(n1283) );
NAND2_X1 U1005 ( .A1(n1243), .A2(n1285), .ZN(n1284) );
NAND3_X1 U1006 ( .A1(n1243), .A2(n1285), .A3(G101), .ZN(n1282) );
XNOR2_X1 U1007 ( .A(G210), .B(KEYINPUT62), .ZN(n1285) );
AND2_X1 U1008 ( .A1(n1267), .A2(n1286), .ZN(n1243) );
XNOR2_X1 U1009 ( .A(n1287), .B(n1123), .ZN(n1281) );
XOR2_X1 U1010 ( .A(n1288), .B(n1289), .Z(n1123) );
XNOR2_X1 U1011 ( .A(KEYINPUT10), .B(n1290), .ZN(n1289) );
XOR2_X1 U1012 ( .A(n1077), .B(n1291), .Z(n1288) );
XNOR2_X1 U1013 ( .A(G131), .B(n1292), .ZN(n1077) );
XOR2_X1 U1014 ( .A(G137), .B(G134), .Z(n1292) );
NAND2_X1 U1015 ( .A1(KEYINPUT60), .A2(n1134), .ZN(n1287) );
INV_X1 U1016 ( .A(n1194), .ZN(n1030) );
NAND2_X1 U1017 ( .A1(n1031), .A2(n1032), .ZN(n1194) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1293), .ZN(n1032) );
XNOR2_X1 U1019 ( .A(n1053), .B(KEYINPUT56), .ZN(n1031) );
XOR2_X1 U1020 ( .A(n1294), .B(n1140), .Z(n1053) );
NAND2_X1 U1021 ( .A1(G210), .A2(n1293), .ZN(n1140) );
NAND2_X1 U1022 ( .A1(n1286), .A2(n1223), .ZN(n1293) );
INV_X1 U1023 ( .A(G237), .ZN(n1286) );
NAND2_X1 U1024 ( .A1(n1295), .A2(n1223), .ZN(n1294) );
INV_X1 U1025 ( .A(G902), .ZN(n1223) );
XNOR2_X1 U1026 ( .A(n1135), .B(n1296), .ZN(n1295) );
XNOR2_X1 U1027 ( .A(n1297), .B(n1138), .ZN(n1296) );
AND2_X1 U1028 ( .A1(G224), .A2(n1267), .ZN(n1138) );
XNOR2_X1 U1029 ( .A(n1038), .B(KEYINPUT46), .ZN(n1267) );
INV_X1 U1030 ( .A(G953), .ZN(n1038) );
NAND3_X1 U1031 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1297) );
NAND2_X1 U1032 ( .A1(n1124), .A2(n1301), .ZN(n1300) );
NAND3_X1 U1033 ( .A1(n1302), .A2(n1134), .A3(KEYINPUT17), .ZN(n1299) );
INV_X1 U1034 ( .A(n1124), .ZN(n1134) );
XOR2_X1 U1035 ( .A(G128), .B(n1277), .Z(n1124) );
XOR2_X1 U1036 ( .A(G143), .B(G146), .Z(n1277) );
INV_X1 U1037 ( .A(n1301), .ZN(n1302) );
NAND2_X1 U1038 ( .A1(n1303), .A2(n1198), .ZN(n1301) );
XOR2_X1 U1039 ( .A(KEYINPUT53), .B(KEYINPUT51), .Z(n1303) );
OR2_X1 U1040 ( .A1(n1198), .A2(KEYINPUT17), .ZN(n1298) );
INV_X1 U1041 ( .A(G125), .ZN(n1198) );
XNOR2_X1 U1042 ( .A(n1093), .B(n1304), .ZN(n1135) );
XNOR2_X1 U1043 ( .A(n1305), .B(n1092), .ZN(n1304) );
XNOR2_X1 U1044 ( .A(n1306), .B(KEYINPUT44), .ZN(n1092) );
NAND2_X1 U1045 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1046 ( .A1(n1275), .A2(n1309), .ZN(n1308) );
NAND2_X1 U1047 ( .A1(G101), .A2(n1310), .ZN(n1309) );
NAND2_X1 U1048 ( .A1(KEYINPUT6), .A2(KEYINPUT15), .ZN(n1310) );
NAND3_X1 U1049 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1307) );
INV_X1 U1050 ( .A(KEYINPUT6), .ZN(n1313) );
OR2_X1 U1051 ( .A1(n1195), .A2(KEYINPUT15), .ZN(n1312) );
NAND2_X1 U1052 ( .A1(KEYINPUT15), .A2(n1314), .ZN(n1311) );
OR2_X1 U1053 ( .A1(n1195), .A2(n1275), .ZN(n1314) );
XNOR2_X1 U1054 ( .A(G104), .B(G107), .ZN(n1275) );
INV_X1 U1055 ( .A(G101), .ZN(n1195) );
NAND2_X1 U1056 ( .A1(KEYINPUT8), .A2(n1089), .ZN(n1305) );
XNOR2_X1 U1057 ( .A(G110), .B(n1315), .ZN(n1089) );
XOR2_X1 U1058 ( .A(KEYINPUT38), .B(G122), .Z(n1315) );
XOR2_X1 U1059 ( .A(n1316), .B(n1291), .Z(n1093) );
XOR2_X1 U1060 ( .A(G113), .B(KEYINPUT14), .Z(n1291) );
NAND2_X1 U1061 ( .A1(KEYINPUT26), .A2(n1290), .ZN(n1316) );
XNOR2_X1 U1062 ( .A(G116), .B(G119), .ZN(n1290) );
endmodule


