//Key = 0010101000100001101101111011010111110111011001000100011011011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;

XNOR2_X1 U759 ( .A(n1051), .B(n1052), .ZN(G9) );
NOR2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(G75) );
NOR4_X1 U761 ( .A1(n1055), .A2(n1056), .A3(G953), .A4(n1057), .ZN(n1054) );
NOR3_X1 U762 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
INV_X1 U763 ( .A(n1061), .ZN(n1060) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NOR2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U767 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U769 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR3_X1 U770 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1066) );
NOR3_X1 U771 ( .A1(n1075), .A2(n1077), .A3(n1069), .ZN(n1062) );
NAND3_X1 U772 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1055) );
NAND2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND3_X1 U775 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NAND2_X1 U776 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NAND2_X1 U777 ( .A1(n1061), .A2(n1090), .ZN(n1089) );
XNOR2_X1 U778 ( .A(KEYINPUT5), .B(n1091), .ZN(n1090) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NAND2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XOR2_X1 U781 ( .A(n1096), .B(KEYINPUT55), .Z(n1083) );
NAND4_X1 U782 ( .A1(n1087), .A2(n1097), .A3(n1092), .A4(n1061), .ZN(n1096) );
INV_X1 U783 ( .A(n1058), .ZN(n1087) );
NOR3_X1 U784 ( .A1(n1057), .A2(G953), .A3(G952), .ZN(n1053) );
AND4_X1 U785 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1057) );
NOR3_X1 U786 ( .A1(n1102), .A2(n1069), .A3(n1103), .ZN(n1101) );
INV_X1 U787 ( .A(n1092), .ZN(n1069) );
NAND3_X1 U788 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1102) );
XNOR2_X1 U789 ( .A(n1107), .B(n1108), .ZN(n1106) );
NAND2_X1 U790 ( .A1(KEYINPUT48), .A2(n1109), .ZN(n1105) );
OR2_X1 U791 ( .A1(n1110), .A2(KEYINPUT48), .ZN(n1104) );
NOR3_X1 U792 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1100) );
XNOR2_X1 U793 ( .A(n1114), .B(n1115), .ZN(n1098) );
NOR2_X1 U794 ( .A1(n1116), .A2(KEYINPUT46), .ZN(n1115) );
XOR2_X1 U795 ( .A(n1117), .B(n1118), .Z(G72) );
XOR2_X1 U796 ( .A(n1119), .B(n1120), .Z(n1118) );
NAND2_X1 U797 ( .A1(G953), .A2(n1121), .ZN(n1120) );
NAND2_X1 U798 ( .A1(G900), .A2(G227), .ZN(n1121) );
NAND2_X1 U799 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
NAND2_X1 U800 ( .A1(G953), .A2(n1124), .ZN(n1123) );
XOR2_X1 U801 ( .A(n1125), .B(n1126), .Z(n1122) );
XNOR2_X1 U802 ( .A(n1127), .B(n1128), .ZN(n1126) );
XNOR2_X1 U803 ( .A(n1129), .B(G134), .ZN(n1128) );
INV_X1 U804 ( .A(G131), .ZN(n1127) );
XOR2_X1 U805 ( .A(n1130), .B(n1131), .Z(n1125) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1130) );
NOR2_X1 U807 ( .A1(KEYINPUT30), .A2(n1134), .ZN(n1133) );
NOR2_X1 U808 ( .A1(n1080), .A2(G953), .ZN(n1117) );
NAND2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(G69) );
NAND2_X1 U810 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U811 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
OR2_X1 U812 ( .A1(n1141), .A2(KEYINPUT62), .ZN(n1140) );
INV_X1 U813 ( .A(n1142), .ZN(n1137) );
NAND3_X1 U814 ( .A1(n1143), .A2(n1144), .A3(KEYINPUT62), .ZN(n1135) );
NAND2_X1 U815 ( .A1(n1139), .A2(n1141), .ZN(n1144) );
INV_X1 U816 ( .A(KEYINPUT34), .ZN(n1141) );
NAND2_X1 U817 ( .A1(KEYINPUT34), .A2(n1145), .ZN(n1143) );
NAND2_X1 U818 ( .A1(n1142), .A2(n1139), .ZN(n1145) );
NAND2_X1 U819 ( .A1(G953), .A2(n1146), .ZN(n1139) );
NAND2_X1 U820 ( .A1(G898), .A2(G224), .ZN(n1146) );
NAND2_X1 U821 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
NAND2_X1 U822 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XNOR2_X1 U823 ( .A(n1151), .B(n1078), .ZN(n1149) );
NAND3_X1 U824 ( .A1(n1151), .A2(n1152), .A3(G953), .ZN(n1147) );
XNOR2_X1 U825 ( .A(G898), .B(KEYINPUT45), .ZN(n1152) );
XNOR2_X1 U826 ( .A(n1153), .B(n1154), .ZN(n1151) );
XOR2_X1 U827 ( .A(KEYINPUT57), .B(KEYINPUT41), .Z(n1154) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U830 ( .A(KEYINPUT17), .B(n1159), .ZN(n1158) );
NOR2_X1 U831 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NOR2_X1 U832 ( .A1(n1155), .A2(n1162), .ZN(G63) );
XNOR2_X1 U833 ( .A(n1163), .B(n1164), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1109), .A2(n1161), .ZN(n1163) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1165), .ZN(G60) );
NOR3_X1 U836 ( .A1(n1116), .A2(n1166), .A3(n1167), .ZN(n1165) );
NOR3_X1 U837 ( .A1(n1168), .A2(n1114), .A3(n1161), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
AND2_X1 U839 ( .A1(n1171), .A2(G475), .ZN(n1169) );
XNOR2_X1 U840 ( .A(n1172), .B(n1173), .ZN(G6) );
NOR2_X1 U841 ( .A1(KEYINPUT25), .A2(n1174), .ZN(n1173) );
NOR2_X1 U842 ( .A1(n1155), .A2(n1175), .ZN(G57) );
XOR2_X1 U843 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U844 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1176) );
NOR2_X1 U846 ( .A1(n1182), .A2(n1161), .ZN(n1181) );
XOR2_X1 U847 ( .A(n1183), .B(KEYINPUT63), .Z(n1180) );
NAND2_X1 U848 ( .A1(KEYINPUT31), .A2(n1184), .ZN(n1183) );
NOR2_X1 U849 ( .A1(n1155), .A2(n1185), .ZN(G54) );
XOR2_X1 U850 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U851 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR2_X1 U852 ( .A1(KEYINPUT50), .A2(n1190), .ZN(n1189) );
NOR2_X1 U853 ( .A1(KEYINPUT58), .A2(n1191), .ZN(n1188) );
XNOR2_X1 U854 ( .A(n1192), .B(n1193), .ZN(n1191) );
XNOR2_X1 U855 ( .A(n1194), .B(KEYINPUT44), .ZN(n1193) );
XOR2_X1 U856 ( .A(n1195), .B(n1196), .Z(n1186) );
NOR2_X1 U857 ( .A1(n1197), .A2(n1161), .ZN(n1196) );
NOR2_X1 U858 ( .A1(n1155), .A2(n1198), .ZN(G51) );
XOR2_X1 U859 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U860 ( .A1(n1108), .A2(n1161), .ZN(n1200) );
NAND2_X1 U861 ( .A1(G902), .A2(n1171), .ZN(n1161) );
NAND2_X1 U862 ( .A1(n1201), .A2(n1078), .ZN(n1171) );
AND4_X1 U863 ( .A1(n1202), .A2(n1172), .A3(n1203), .A4(n1204), .ZN(n1078) );
NOR4_X1 U864 ( .A1(n1052), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1204) );
AND3_X1 U865 ( .A1(n1208), .A2(n1061), .A3(n1209), .ZN(n1052) );
OR2_X1 U866 ( .A1(n1210), .A2(n1211), .ZN(n1203) );
NAND3_X1 U867 ( .A1(n1209), .A2(n1061), .A3(n1097), .ZN(n1172) );
NAND2_X1 U868 ( .A1(n1212), .A2(n1213), .ZN(n1202) );
NAND2_X1 U869 ( .A1(n1214), .A2(n1095), .ZN(n1213) );
XNOR2_X1 U870 ( .A(n1215), .B(KEYINPUT9), .ZN(n1214) );
XNOR2_X1 U871 ( .A(n1080), .B(KEYINPUT33), .ZN(n1201) );
AND2_X1 U872 ( .A1(n1216), .A2(n1217), .ZN(n1080) );
NOR4_X1 U873 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
NOR3_X1 U874 ( .A1(n1222), .A2(n1223), .A3(n1075), .ZN(n1219) );
INV_X1 U875 ( .A(n1081), .ZN(n1075) );
XNOR2_X1 U876 ( .A(KEYINPUT49), .B(n1091), .ZN(n1222) );
INV_X1 U877 ( .A(n1224), .ZN(n1218) );
AND4_X1 U878 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1216) );
NAND2_X1 U879 ( .A1(n1229), .A2(KEYINPUT27), .ZN(n1199) );
XOR2_X1 U880 ( .A(n1230), .B(n1153), .Z(n1229) );
NAND2_X1 U881 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NOR2_X1 U882 ( .A1(n1150), .A2(G952), .ZN(n1155) );
XNOR2_X1 U883 ( .A(G146), .B(n1224), .ZN(G48) );
NAND3_X1 U884 ( .A1(n1097), .A2(n1233), .A3(n1234), .ZN(n1224) );
NOR3_X1 U885 ( .A1(n1211), .A2(n1235), .A3(n1091), .ZN(n1234) );
XOR2_X1 U886 ( .A(n1228), .B(n1236), .Z(G45) );
NAND2_X1 U887 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1236) );
NAND2_X1 U888 ( .A1(n1237), .A2(n1238), .ZN(n1228) );
XNOR2_X1 U889 ( .A(G140), .B(n1239), .ZN(G42) );
NOR2_X1 U890 ( .A1(n1240), .A2(KEYINPUT36), .ZN(n1239) );
INV_X1 U891 ( .A(n1227), .ZN(n1240) );
NAND4_X1 U892 ( .A1(n1215), .A2(n1081), .A3(n1241), .A4(n1097), .ZN(n1227) );
NOR2_X1 U893 ( .A1(n1235), .A2(n1091), .ZN(n1241) );
XOR2_X1 U894 ( .A(n1242), .B(n1243), .Z(G39) );
NOR3_X1 U895 ( .A1(n1223), .A2(n1244), .A3(n1091), .ZN(n1243) );
XNOR2_X1 U896 ( .A(n1081), .B(KEYINPUT47), .ZN(n1244) );
NAND3_X1 U897 ( .A1(n1233), .A2(n1245), .A3(n1085), .ZN(n1223) );
NAND2_X1 U898 ( .A1(KEYINPUT21), .A2(n1129), .ZN(n1242) );
XOR2_X1 U899 ( .A(n1246), .B(G134), .Z(G36) );
NAND2_X1 U900 ( .A1(KEYINPUT54), .A2(n1226), .ZN(n1246) );
NAND3_X1 U901 ( .A1(n1081), .A2(n1208), .A3(n1238), .ZN(n1226) );
XNOR2_X1 U902 ( .A(G131), .B(n1225), .ZN(G33) );
NAND3_X1 U903 ( .A1(n1081), .A2(n1097), .A3(n1238), .ZN(n1225) );
NOR3_X1 U904 ( .A1(n1091), .A2(n1235), .A3(n1095), .ZN(n1238) );
INV_X1 U905 ( .A(n1245), .ZN(n1235) );
NOR2_X1 U906 ( .A1(n1072), .A2(n1113), .ZN(n1081) );
INV_X1 U907 ( .A(n1073), .ZN(n1113) );
XOR2_X1 U908 ( .A(G128), .B(n1221), .Z(G30) );
AND4_X1 U909 ( .A1(n1247), .A2(n1245), .A3(n1071), .A4(n1248), .ZN(n1221) );
NOR2_X1 U910 ( .A1(n1077), .A2(n1249), .ZN(n1248) );
XNOR2_X1 U911 ( .A(G101), .B(n1250), .ZN(G3) );
NAND2_X1 U912 ( .A1(n1212), .A2(n1251), .ZN(n1250) );
INV_X1 U913 ( .A(n1252), .ZN(n1212) );
XNOR2_X1 U914 ( .A(n1253), .B(n1134), .ZN(G27) );
INV_X1 U915 ( .A(G125), .ZN(n1134) );
NAND2_X1 U916 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND3_X1 U917 ( .A1(n1256), .A2(n1211), .A3(n1257), .ZN(n1255) );
INV_X1 U918 ( .A(KEYINPUT35), .ZN(n1257) );
NAND2_X1 U919 ( .A1(n1220), .A2(KEYINPUT35), .ZN(n1254) );
AND2_X1 U920 ( .A1(n1256), .A2(n1071), .ZN(n1220) );
AND4_X1 U921 ( .A1(n1215), .A2(n1097), .A3(n1092), .A4(n1245), .ZN(n1256) );
NAND2_X1 U922 ( .A1(n1058), .A2(n1258), .ZN(n1245) );
NAND4_X1 U923 ( .A1(G902), .A2(G953), .A3(n1259), .A4(n1124), .ZN(n1258) );
INV_X1 U924 ( .A(G900), .ZN(n1124) );
XOR2_X1 U925 ( .A(G122), .B(n1207), .Z(G24) );
AND3_X1 U926 ( .A1(n1237), .A2(n1061), .A3(n1260), .ZN(n1207) );
NOR2_X1 U927 ( .A1(n1261), .A2(n1103), .ZN(n1061) );
AND3_X1 U928 ( .A1(n1262), .A2(n1071), .A3(n1263), .ZN(n1237) );
XNOR2_X1 U929 ( .A(G119), .B(n1264), .ZN(G21) );
NAND2_X1 U930 ( .A1(n1265), .A2(n1071), .ZN(n1264) );
XOR2_X1 U931 ( .A(n1210), .B(KEYINPUT37), .Z(n1265) );
NAND3_X1 U932 ( .A1(n1085), .A2(n1233), .A3(n1260), .ZN(n1210) );
INV_X1 U933 ( .A(n1249), .ZN(n1233) );
NAND2_X1 U934 ( .A1(n1103), .A2(n1261), .ZN(n1249) );
XOR2_X1 U935 ( .A(G116), .B(n1206), .Z(G18) );
AND2_X1 U936 ( .A1(n1266), .A2(n1208), .ZN(n1206) );
INV_X1 U937 ( .A(n1077), .ZN(n1208) );
NAND2_X1 U938 ( .A1(n1262), .A2(n1267), .ZN(n1077) );
XNOR2_X1 U939 ( .A(n1268), .B(KEYINPUT51), .ZN(n1262) );
NAND2_X1 U940 ( .A1(n1269), .A2(n1270), .ZN(G15) );
NAND2_X1 U941 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND2_X1 U942 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
OR2_X1 U943 ( .A1(n1205), .A2(KEYINPUT4), .ZN(n1274) );
INV_X1 U944 ( .A(n1275), .ZN(n1205) );
NAND2_X1 U945 ( .A1(KEYINPUT4), .A2(n1276), .ZN(n1273) );
OR2_X1 U946 ( .A1(n1272), .A2(n1276), .ZN(n1269) );
NAND2_X1 U947 ( .A1(KEYINPUT15), .A2(n1275), .ZN(n1276) );
NAND2_X1 U948 ( .A1(n1266), .A2(n1097), .ZN(n1275) );
AND2_X1 U949 ( .A1(n1263), .A2(n1268), .ZN(n1097) );
XNOR2_X1 U950 ( .A(n1267), .B(KEYINPUT40), .ZN(n1263) );
AND3_X1 U951 ( .A1(n1251), .A2(n1071), .A3(n1260), .ZN(n1266) );
AND2_X1 U952 ( .A1(n1092), .A2(n1277), .ZN(n1260) );
NOR2_X1 U953 ( .A1(n1076), .A2(n1278), .ZN(n1092) );
INV_X1 U954 ( .A(n1074), .ZN(n1278) );
INV_X1 U955 ( .A(n1095), .ZN(n1251) );
NAND2_X1 U956 ( .A1(n1279), .A2(n1103), .ZN(n1095) );
XOR2_X1 U957 ( .A(n1280), .B(n1281), .Z(G12) );
NOR2_X1 U958 ( .A1(n1094), .A2(n1252), .ZN(n1281) );
NAND2_X1 U959 ( .A1(n1085), .A2(n1209), .ZN(n1252) );
AND3_X1 U960 ( .A1(n1247), .A2(n1277), .A3(n1071), .ZN(n1209) );
INV_X1 U961 ( .A(n1211), .ZN(n1071) );
NAND2_X1 U962 ( .A1(n1282), .A2(n1073), .ZN(n1211) );
NAND2_X1 U963 ( .A1(G214), .A2(n1283), .ZN(n1073) );
XNOR2_X1 U964 ( .A(KEYINPUT24), .B(n1072), .ZN(n1282) );
XNOR2_X1 U965 ( .A(n1284), .B(n1107), .ZN(n1072) );
NAND2_X1 U966 ( .A1(n1285), .A2(n1286), .ZN(n1107) );
XOR2_X1 U967 ( .A(n1287), .B(n1153), .Z(n1285) );
XOR2_X1 U968 ( .A(n1288), .B(n1289), .Z(n1153) );
XNOR2_X1 U969 ( .A(n1272), .B(n1290), .ZN(n1289) );
XOR2_X1 U970 ( .A(KEYINPUT28), .B(G119), .Z(n1290) );
XOR2_X1 U971 ( .A(n1291), .B(n1292), .Z(n1288) );
NOR2_X1 U972 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NOR3_X1 U973 ( .A1(KEYINPUT26), .A2(G107), .A3(n1174), .ZN(n1294) );
NOR2_X1 U974 ( .A1(n1295), .A2(n1296), .ZN(n1293) );
INV_X1 U975 ( .A(KEYINPUT26), .ZN(n1296) );
XNOR2_X1 U976 ( .A(n1297), .B(n1298), .ZN(n1291) );
NAND2_X1 U977 ( .A1(n1299), .A2(n1231), .ZN(n1287) );
NAND3_X1 U978 ( .A1(n1300), .A2(G224), .A3(n1301), .ZN(n1231) );
XNOR2_X1 U979 ( .A(n1302), .B(G125), .ZN(n1301) );
XNOR2_X1 U980 ( .A(KEYINPUT10), .B(n1232), .ZN(n1299) );
NAND2_X1 U981 ( .A1(n1303), .A2(n1304), .ZN(n1232) );
NAND2_X1 U982 ( .A1(G224), .A2(n1300), .ZN(n1304) );
XNOR2_X1 U983 ( .A(G125), .B(n1305), .ZN(n1303) );
NAND2_X1 U984 ( .A1(KEYINPUT6), .A2(n1108), .ZN(n1284) );
NAND2_X1 U985 ( .A1(G210), .A2(n1283), .ZN(n1108) );
NAND2_X1 U986 ( .A1(n1306), .A2(n1286), .ZN(n1283) );
INV_X1 U987 ( .A(G237), .ZN(n1306) );
NAND2_X1 U988 ( .A1(n1307), .A2(n1058), .ZN(n1277) );
NAND3_X1 U989 ( .A1(n1259), .A2(n1150), .A3(G952), .ZN(n1058) );
XOR2_X1 U990 ( .A(KEYINPUT38), .B(n1308), .Z(n1307) );
NOR4_X1 U991 ( .A1(G898), .A2(n1309), .A3(n1150), .A4(n1286), .ZN(n1308) );
INV_X1 U992 ( .A(n1259), .ZN(n1309) );
NAND2_X1 U993 ( .A1(G237), .A2(G234), .ZN(n1259) );
XOR2_X1 U994 ( .A(n1091), .B(KEYINPUT16), .Z(n1247) );
NAND2_X1 U995 ( .A1(n1076), .A2(n1074), .ZN(n1091) );
NAND2_X1 U996 ( .A1(G221), .A2(n1310), .ZN(n1074) );
XOR2_X1 U997 ( .A(n1311), .B(n1197), .Z(n1076) );
INV_X1 U998 ( .A(G469), .ZN(n1197) );
NAND2_X1 U999 ( .A1(n1312), .A2(n1286), .ZN(n1311) );
XNOR2_X1 U1000 ( .A(n1313), .B(n1314), .ZN(n1312) );
INV_X1 U1001 ( .A(n1192), .ZN(n1314) );
XNOR2_X1 U1002 ( .A(n1315), .B(n1295), .ZN(n1192) );
XNOR2_X1 U1003 ( .A(n1174), .B(G107), .ZN(n1295) );
INV_X1 U1004 ( .A(G104), .ZN(n1174) );
XOR2_X1 U1005 ( .A(n1132), .B(KEYINPUT43), .Z(n1315) );
NAND2_X1 U1006 ( .A1(n1316), .A2(n1317), .ZN(n1132) );
OR2_X1 U1007 ( .A1(n1318), .A2(G128), .ZN(n1317) );
XOR2_X1 U1008 ( .A(n1319), .B(KEYINPUT13), .Z(n1316) );
NAND2_X1 U1009 ( .A1(G128), .A2(n1318), .ZN(n1319) );
XOR2_X1 U1010 ( .A(n1195), .B(n1297), .Z(n1313) );
XOR2_X1 U1011 ( .A(G110), .B(n1194), .Z(n1297) );
XOR2_X1 U1012 ( .A(G101), .B(KEYINPUT29), .Z(n1194) );
XOR2_X1 U1013 ( .A(n1320), .B(n1131), .Z(n1195) );
XOR2_X1 U1014 ( .A(n1321), .B(n1322), .Z(n1320) );
NOR2_X1 U1015 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XNOR2_X1 U1016 ( .A(KEYINPUT12), .B(n1300), .ZN(n1324) );
INV_X1 U1017 ( .A(G227), .ZN(n1323) );
INV_X1 U1018 ( .A(n1065), .ZN(n1085) );
NAND2_X1 U1019 ( .A1(n1268), .A2(n1267), .ZN(n1065) );
XNOR2_X1 U1020 ( .A(n1325), .B(n1116), .ZN(n1267) );
NOR2_X1 U1021 ( .A1(n1170), .A2(G902), .ZN(n1116) );
INV_X1 U1022 ( .A(n1168), .ZN(n1170) );
XNOR2_X1 U1023 ( .A(n1326), .B(n1327), .ZN(n1168) );
XNOR2_X1 U1024 ( .A(G122), .B(n1272), .ZN(n1327) );
INV_X1 U1025 ( .A(G113), .ZN(n1272) );
XNOR2_X1 U1026 ( .A(G104), .B(n1328), .ZN(n1326) );
NOR2_X1 U1027 ( .A1(KEYINPUT11), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1028 ( .A(n1330), .B(n1331), .Z(n1329) );
XOR2_X1 U1029 ( .A(n1332), .B(n1333), .Z(n1331) );
NOR2_X1 U1030 ( .A1(KEYINPUT20), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1031 ( .A(G146), .B(n1335), .ZN(n1334) );
NAND2_X1 U1032 ( .A1(n1336), .A2(G214), .ZN(n1332) );
XNOR2_X1 U1033 ( .A(G131), .B(G143), .ZN(n1330) );
NAND2_X1 U1034 ( .A1(KEYINPUT2), .A2(n1114), .ZN(n1325) );
INV_X1 U1035 ( .A(G475), .ZN(n1114) );
NOR2_X1 U1036 ( .A1(n1337), .A2(n1112), .ZN(n1268) );
AND3_X1 U1037 ( .A1(n1109), .A2(n1286), .A3(n1164), .ZN(n1112) );
INV_X1 U1038 ( .A(G478), .ZN(n1109) );
INV_X1 U1039 ( .A(n1110), .ZN(n1337) );
NAND2_X1 U1040 ( .A1(G478), .A2(n1338), .ZN(n1110) );
NAND2_X1 U1041 ( .A1(n1164), .A2(n1286), .ZN(n1338) );
XOR2_X1 U1042 ( .A(n1339), .B(n1340), .Z(n1164) );
XOR2_X1 U1043 ( .A(n1341), .B(n1342), .Z(n1340) );
XOR2_X1 U1044 ( .A(G134), .B(G128), .Z(n1342) );
XOR2_X1 U1045 ( .A(KEYINPUT0), .B(G143), .Z(n1341) );
XNOR2_X1 U1046 ( .A(n1298), .B(n1343), .ZN(n1339) );
XOR2_X1 U1047 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1048 ( .A1(KEYINPUT53), .A2(n1051), .ZN(n1345) );
INV_X1 U1049 ( .A(G107), .ZN(n1051) );
NAND2_X1 U1050 ( .A1(G217), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1051 ( .A(G116), .B(G122), .Z(n1298) );
INV_X1 U1052 ( .A(n1215), .ZN(n1094) );
NOR2_X1 U1053 ( .A1(n1103), .A2(n1279), .ZN(n1215) );
INV_X1 U1054 ( .A(n1261), .ZN(n1279) );
NAND3_X1 U1055 ( .A1(n1347), .A2(n1348), .A3(n1099), .ZN(n1261) );
NAND3_X1 U1056 ( .A1(n1160), .A2(n1286), .A3(n1159), .ZN(n1099) );
NAND2_X1 U1057 ( .A1(n1160), .A2(n1349), .ZN(n1348) );
INV_X1 U1058 ( .A(KEYINPUT19), .ZN(n1349) );
NAND2_X1 U1059 ( .A1(n1111), .A2(KEYINPUT19), .ZN(n1347) );
NOR2_X1 U1060 ( .A1(n1160), .A2(n1350), .ZN(n1111) );
AND2_X1 U1061 ( .A1(n1159), .A2(n1286), .ZN(n1350) );
NAND2_X1 U1062 ( .A1(n1351), .A2(n1352), .ZN(n1159) );
OR2_X1 U1063 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
XOR2_X1 U1064 ( .A(n1355), .B(KEYINPUT7), .Z(n1351) );
NAND2_X1 U1065 ( .A1(n1354), .A2(n1353), .ZN(n1355) );
XOR2_X1 U1066 ( .A(n1356), .B(n1129), .Z(n1353) );
INV_X1 U1067 ( .A(G137), .ZN(n1129) );
NAND2_X1 U1068 ( .A1(n1346), .A2(G221), .ZN(n1356) );
AND2_X1 U1069 ( .A1(G234), .A2(n1300), .ZN(n1346) );
XNOR2_X1 U1070 ( .A(n1357), .B(n1358), .ZN(n1354) );
XNOR2_X1 U1071 ( .A(n1190), .B(n1359), .ZN(n1358) );
XNOR2_X1 U1072 ( .A(n1360), .B(G128), .ZN(n1359) );
XNOR2_X1 U1073 ( .A(n1361), .B(n1362), .ZN(n1357) );
NAND2_X1 U1074 ( .A1(KEYINPUT32), .A2(G119), .ZN(n1362) );
NAND2_X1 U1075 ( .A1(KEYINPUT18), .A2(n1335), .ZN(n1361) );
XNOR2_X1 U1076 ( .A(G125), .B(n1131), .ZN(n1335) );
XOR2_X1 U1077 ( .A(G140), .B(KEYINPUT1), .Z(n1131) );
NAND2_X1 U1078 ( .A1(G217), .A2(n1310), .ZN(n1160) );
NAND2_X1 U1079 ( .A1(G234), .A2(n1286), .ZN(n1310) );
XOR2_X1 U1080 ( .A(n1363), .B(n1182), .Z(n1103) );
INV_X1 U1081 ( .A(G472), .ZN(n1182) );
NAND2_X1 U1082 ( .A1(n1364), .A2(n1286), .ZN(n1363) );
INV_X1 U1083 ( .A(G902), .ZN(n1286) );
XOR2_X1 U1084 ( .A(n1178), .B(n1365), .Z(n1364) );
XNOR2_X1 U1085 ( .A(n1366), .B(n1184), .ZN(n1365) );
XNOR2_X1 U1086 ( .A(n1367), .B(n1368), .ZN(n1184) );
XNOR2_X1 U1087 ( .A(G113), .B(n1369), .ZN(n1368) );
NAND2_X1 U1088 ( .A1(KEYINPUT60), .A2(n1370), .ZN(n1369) );
XOR2_X1 U1089 ( .A(KEYINPUT22), .B(G119), .Z(n1370) );
XNOR2_X1 U1090 ( .A(G116), .B(KEYINPUT52), .ZN(n1367) );
NAND2_X1 U1091 ( .A1(KEYINPUT39), .A2(n1371), .ZN(n1366) );
XOR2_X1 U1092 ( .A(KEYINPUT3), .B(n1179), .Z(n1371) );
XNOR2_X1 U1093 ( .A(n1372), .B(G101), .ZN(n1179) );
NAND2_X1 U1094 ( .A1(n1336), .A2(G210), .ZN(n1372) );
AND2_X1 U1095 ( .A1(n1373), .A2(n1300), .ZN(n1336) );
XOR2_X1 U1096 ( .A(n1150), .B(KEYINPUT14), .Z(n1300) );
INV_X1 U1097 ( .A(G953), .ZN(n1150) );
XNOR2_X1 U1098 ( .A(G237), .B(KEYINPUT61), .ZN(n1373) );
XNOR2_X1 U1099 ( .A(n1321), .B(n1305), .ZN(n1178) );
INV_X1 U1100 ( .A(n1302), .ZN(n1305) );
XNOR2_X1 U1101 ( .A(n1374), .B(G128), .ZN(n1302) );
NAND2_X1 U1102 ( .A1(KEYINPUT23), .A2(n1318), .ZN(n1374) );
XNOR2_X1 U1103 ( .A(G143), .B(n1360), .ZN(n1318) );
INV_X1 U1104 ( .A(G146), .ZN(n1360) );
NAND2_X1 U1105 ( .A1(n1375), .A2(n1376), .ZN(n1321) );
NAND2_X1 U1106 ( .A1(G131), .A2(n1377), .ZN(n1376) );
XOR2_X1 U1107 ( .A(KEYINPUT59), .B(n1378), .Z(n1375) );
NOR2_X1 U1108 ( .A1(G131), .A2(n1377), .ZN(n1378) );
XNOR2_X1 U1109 ( .A(n1379), .B(G137), .ZN(n1377) );
NAND2_X1 U1110 ( .A1(KEYINPUT42), .A2(G134), .ZN(n1379) );
NOR2_X1 U1111 ( .A1(KEYINPUT8), .A2(n1190), .ZN(n1280) );
INV_X1 U1112 ( .A(G110), .ZN(n1190) );
endmodule


