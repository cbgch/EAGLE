//Key = 0010000101010000001011011101010110010001010000010100110111100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329;

XOR2_X1 U742 ( .A(n1028), .B(n1029), .Z(G9) );
NAND2_X1 U743 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
XOR2_X1 U744 ( .A(KEYINPUT61), .B(G107), .Z(n1031) );
XNOR2_X1 U745 ( .A(KEYINPUT34), .B(KEYINPUT12), .ZN(n1030) );
NAND4_X1 U746 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1028) );
XNOR2_X1 U747 ( .A(n1036), .B(KEYINPUT57), .ZN(n1032) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR4_X1 U749 ( .A1(n1039), .A2(n1040), .A3(G953), .A4(n1041), .ZN(n1038) );
NOR2_X1 U750 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR3_X1 U751 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1042) );
AND2_X1 U752 ( .A1(n1034), .A2(n1047), .ZN(n1046) );
NOR3_X1 U753 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1045) );
NOR4_X1 U754 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1050) );
NOR2_X1 U755 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U756 ( .A1(KEYINPUT42), .A2(n1057), .ZN(n1053) );
AND2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1052) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1049) );
AND2_X1 U759 ( .A1(n1033), .A2(KEYINPUT42), .ZN(n1061) );
XOR2_X1 U760 ( .A(KEYINPUT30), .B(n1062), .Z(n1044) );
AND4_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1060), .A4(n1065), .ZN(n1062) );
NAND3_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1039) );
NAND2_X1 U763 ( .A1(n1047), .A2(n1069), .ZN(n1067) );
NAND3_X1 U764 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND3_X1 U765 ( .A1(n1073), .A2(n1074), .A3(n1060), .ZN(n1072) );
OR2_X1 U766 ( .A1(n1075), .A2(KEYINPUT23), .ZN(n1074) );
NAND2_X1 U767 ( .A1(KEYINPUT23), .A2(n1076), .ZN(n1073) );
NAND2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
INV_X1 U769 ( .A(n1079), .ZN(n1071) );
NAND3_X1 U770 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1070) );
XNOR2_X1 U771 ( .A(KEYINPUT1), .B(n1043), .ZN(n1081) );
AND3_X1 U772 ( .A1(n1064), .A2(n1063), .A3(n1059), .ZN(n1047) );
NOR3_X1 U773 ( .A1(n1041), .A2(G953), .A3(G952), .ZN(n1037) );
AND4_X1 U774 ( .A1(n1083), .A2(n1075), .A3(n1084), .A4(n1085), .ZN(n1041) );
NOR3_X1 U775 ( .A1(n1051), .A2(n1086), .A3(n1087), .ZN(n1085) );
XOR2_X1 U776 ( .A(n1088), .B(n1089), .Z(n1086) );
NAND2_X1 U777 ( .A1(KEYINPUT31), .A2(n1090), .ZN(n1088) );
XNOR2_X1 U778 ( .A(n1091), .B(KEYINPUT8), .ZN(n1084) );
XNOR2_X1 U779 ( .A(n1092), .B(n1093), .ZN(n1083) );
XOR2_X1 U780 ( .A(n1094), .B(n1095), .Z(G72) );
NAND2_X1 U781 ( .A1(G953), .A2(n1096), .ZN(n1095) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1096) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
XOR2_X1 U784 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U785 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(n1099) );
NAND2_X1 U787 ( .A1(G953), .A2(n1105), .ZN(n1104) );
XOR2_X1 U788 ( .A(n1106), .B(n1107), .Z(n1103) );
NAND2_X1 U789 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
OR2_X1 U790 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U791 ( .A(n1112), .B(KEYINPUT26), .Z(n1108) );
NAND2_X1 U792 ( .A1(n1110), .A2(n1111), .ZN(n1112) );
XNOR2_X1 U793 ( .A(KEYINPUT53), .B(KEYINPUT29), .ZN(n1097) );
XOR2_X1 U794 ( .A(n1113), .B(n1114), .Z(G69) );
XOR2_X1 U795 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U796 ( .A1(n1066), .A2(n1117), .ZN(n1116) );
XNOR2_X1 U797 ( .A(KEYINPUT13), .B(n1101), .ZN(n1117) );
NAND3_X1 U798 ( .A1(n1118), .A2(n1119), .A3(KEYINPUT35), .ZN(n1115) );
NAND2_X1 U799 ( .A1(G953), .A2(n1120), .ZN(n1119) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(n1118) );
XNOR2_X1 U801 ( .A(KEYINPUT58), .B(KEYINPUT36), .ZN(n1122) );
NAND2_X1 U802 ( .A1(G953), .A2(n1123), .ZN(n1113) );
NAND2_X1 U803 ( .A1(G224), .A2(G898), .ZN(n1123) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1124), .A2(n1130), .ZN(G63) );
XOR2_X1 U808 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U809 ( .A(KEYINPUT48), .B(n1133), .ZN(n1132) );
NOR3_X1 U810 ( .A1(n1129), .A2(KEYINPUT14), .A3(n1090), .ZN(n1133) );
INV_X1 U811 ( .A(G478), .ZN(n1090) );
NOR2_X1 U812 ( .A1(n1124), .A2(n1134), .ZN(G60) );
XOR2_X1 U813 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U814 ( .A1(n1137), .A2(n1129), .ZN(n1135) );
XOR2_X1 U815 ( .A(G104), .B(n1138), .Z(G6) );
NOR2_X1 U816 ( .A1(n1124), .A2(n1139), .ZN(G57) );
XOR2_X1 U817 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U818 ( .A(n1142), .B(n1143), .ZN(n1141) );
XNOR2_X1 U819 ( .A(n1144), .B(n1145), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1093), .A2(n1129), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1124), .A2(n1146), .ZN(G54) );
XOR2_X1 U822 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U823 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U824 ( .A1(n1151), .A2(n1129), .ZN(n1150) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(n1147) );
NOR2_X1 U826 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U827 ( .A(KEYINPUT0), .B(n1156), .Z(n1155) );
NOR2_X1 U828 ( .A1(n1157), .A2(n1110), .ZN(n1156) );
AND2_X1 U829 ( .A1(n1157), .A2(n1110), .ZN(n1154) );
NAND2_X1 U830 ( .A1(KEYINPUT39), .A2(n1158), .ZN(n1152) );
XNOR2_X1 U831 ( .A(G110), .B(n1159), .ZN(n1158) );
NOR2_X1 U832 ( .A1(n1124), .A2(n1160), .ZN(G51) );
XOR2_X1 U833 ( .A(n1121), .B(n1161), .Z(n1160) );
XOR2_X1 U834 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U835 ( .A1(n1164), .A2(n1129), .ZN(n1163) );
NAND2_X1 U836 ( .A1(G902), .A2(n1165), .ZN(n1129) );
NAND2_X1 U837 ( .A1(n1166), .A2(n1066), .ZN(n1165) );
AND4_X1 U838 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1066) );
NOR4_X1 U839 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1138), .A2(n1175), .ZN(n1169) );
AND4_X1 U841 ( .A1(n1035), .A2(n1079), .A3(n1176), .A4(n1055), .ZN(n1175) );
AND3_X1 U842 ( .A1(n1065), .A2(n1064), .A3(n1177), .ZN(n1138) );
NAND2_X1 U843 ( .A1(n1178), .A2(n1179), .ZN(n1168) );
XOR2_X1 U844 ( .A(n1180), .B(KEYINPUT20), .Z(n1178) );
NAND2_X1 U845 ( .A1(n1177), .A2(n1033), .ZN(n1167) );
INV_X1 U846 ( .A(n1057), .ZN(n1033) );
NAND2_X1 U847 ( .A1(n1064), .A2(n1181), .ZN(n1057) );
XNOR2_X1 U848 ( .A(n1068), .B(KEYINPUT32), .ZN(n1166) );
INV_X1 U849 ( .A(n1102), .ZN(n1068) );
NAND4_X1 U850 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1102) );
AND4_X1 U851 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
NAND2_X1 U852 ( .A1(n1190), .A2(n1191), .ZN(n1184) );
NAND2_X1 U853 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XNOR2_X1 U854 ( .A(n1065), .B(KEYINPUT28), .ZN(n1192) );
NOR2_X1 U855 ( .A1(KEYINPUT44), .A2(n1194), .ZN(n1162) );
XOR2_X1 U856 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U857 ( .A(G125), .B(n1197), .Z(n1196) );
NOR2_X1 U858 ( .A1(KEYINPUT62), .A2(n1198), .ZN(n1195) );
NOR2_X1 U859 ( .A1(n1101), .A2(G952), .ZN(n1124) );
XNOR2_X1 U860 ( .A(G146), .B(n1199), .ZN(G48) );
NAND2_X1 U861 ( .A1(n1190), .A2(n1065), .ZN(n1199) );
XNOR2_X1 U862 ( .A(G143), .B(n1182), .ZN(G45) );
NAND4_X1 U863 ( .A1(n1200), .A2(n1058), .A3(n1201), .A4(n1087), .ZN(n1182) );
XNOR2_X1 U864 ( .A(G140), .B(n1183), .ZN(G42) );
NAND2_X1 U865 ( .A1(n1202), .A2(n1203), .ZN(n1183) );
XNOR2_X1 U866 ( .A(G137), .B(n1189), .ZN(G39) );
NAND3_X1 U867 ( .A1(n1055), .A2(n1202), .A3(n1176), .ZN(n1189) );
XNOR2_X1 U868 ( .A(G134), .B(n1188), .ZN(G36) );
NAND3_X1 U869 ( .A1(n1202), .A2(n1181), .A3(n1058), .ZN(n1188) );
XNOR2_X1 U870 ( .A(G131), .B(n1187), .ZN(G33) );
NAND3_X1 U871 ( .A1(n1202), .A2(n1065), .A3(n1058), .ZN(n1187) );
AND3_X1 U872 ( .A1(n1034), .A2(n1204), .A3(n1075), .ZN(n1202) );
INV_X1 U873 ( .A(n1043), .ZN(n1075) );
NAND2_X1 U874 ( .A1(n1078), .A2(n1205), .ZN(n1043) );
XNOR2_X1 U875 ( .A(G128), .B(n1206), .ZN(G30) );
NAND2_X1 U876 ( .A1(n1190), .A2(n1181), .ZN(n1206) );
AND3_X1 U877 ( .A1(n1055), .A2(n1091), .A3(n1200), .ZN(n1190) );
AND3_X1 U878 ( .A1(n1034), .A2(n1204), .A3(n1179), .ZN(n1200) );
INV_X1 U879 ( .A(n1207), .ZN(n1179) );
XOR2_X1 U880 ( .A(G101), .B(n1171), .Z(G3) );
AND3_X1 U881 ( .A1(n1059), .A2(n1058), .A3(n1177), .ZN(n1171) );
XNOR2_X1 U882 ( .A(G125), .B(n1186), .ZN(G27) );
NAND3_X1 U883 ( .A1(n1203), .A2(n1204), .A3(n1079), .ZN(n1186) );
NAND2_X1 U884 ( .A1(n1208), .A2(n1209), .ZN(n1204) );
NAND2_X1 U885 ( .A1(n1210), .A2(n1105), .ZN(n1209) );
INV_X1 U886 ( .A(G900), .ZN(n1105) );
XOR2_X1 U887 ( .A(n1211), .B(KEYINPUT10), .Z(n1208) );
AND3_X1 U888 ( .A1(n1091), .A2(n1212), .A3(n1065), .ZN(n1203) );
XOR2_X1 U889 ( .A(G122), .B(n1174), .Z(G24) );
AND3_X1 U890 ( .A1(n1079), .A2(n1064), .A3(n1213), .ZN(n1174) );
AND3_X1 U891 ( .A1(n1201), .A2(n1035), .A3(n1087), .ZN(n1213) );
NOR2_X1 U892 ( .A1(n1091), .A2(n1055), .ZN(n1064) );
XOR2_X1 U893 ( .A(n1214), .B(n1215), .Z(G21) );
NAND2_X1 U894 ( .A1(KEYINPUT18), .A2(G119), .ZN(n1215) );
NAND4_X1 U895 ( .A1(n1055), .A2(n1176), .A3(n1079), .A4(n1216), .ZN(n1214) );
XNOR2_X1 U896 ( .A(KEYINPUT49), .B(n1035), .ZN(n1216) );
NOR2_X1 U897 ( .A1(n1207), .A2(n1051), .ZN(n1079) );
INV_X1 U898 ( .A(n1212), .ZN(n1055) );
XNOR2_X1 U899 ( .A(n1217), .B(n1218), .ZN(G18) );
NOR2_X1 U900 ( .A1(n1207), .A2(n1180), .ZN(n1218) );
NAND4_X1 U901 ( .A1(n1058), .A2(n1060), .A3(n1181), .A4(n1035), .ZN(n1180) );
INV_X1 U902 ( .A(n1193), .ZN(n1181) );
NAND2_X1 U903 ( .A1(n1201), .A2(n1219), .ZN(n1193) );
XOR2_X1 U904 ( .A(n1036), .B(KEYINPUT2), .Z(n1207) );
XOR2_X1 U905 ( .A(G113), .B(n1173), .Z(G15) );
AND4_X1 U906 ( .A1(n1058), .A2(n1065), .A3(n1220), .A4(n1060), .ZN(n1173) );
AND2_X1 U907 ( .A1(n1035), .A2(n1036), .ZN(n1220) );
NOR2_X1 U908 ( .A1(n1219), .A2(n1201), .ZN(n1065) );
INV_X1 U909 ( .A(n1087), .ZN(n1219) );
NOR2_X1 U910 ( .A1(n1212), .A2(n1091), .ZN(n1058) );
XNOR2_X1 U911 ( .A(n1221), .B(n1172), .ZN(G12) );
AND3_X1 U912 ( .A1(n1176), .A2(n1212), .A3(n1177), .ZN(n1172) );
AND3_X1 U913 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1177) );
NOR2_X1 U914 ( .A1(n1078), .A2(n1077), .ZN(n1036) );
INV_X1 U915 ( .A(n1205), .ZN(n1077) );
NAND2_X1 U916 ( .A1(G214), .A2(n1222), .ZN(n1205) );
XNOR2_X1 U917 ( .A(n1223), .B(n1164), .ZN(n1078) );
NAND2_X1 U918 ( .A1(G210), .A2(n1222), .ZN(n1164) );
NAND2_X1 U919 ( .A1(n1224), .A2(n1225), .ZN(n1222) );
INV_X1 U920 ( .A(G237), .ZN(n1225) );
NAND3_X1 U921 ( .A1(n1226), .A2(n1224), .A3(n1227), .ZN(n1223) );
XOR2_X1 U922 ( .A(n1228), .B(KEYINPUT5), .Z(n1227) );
OR2_X1 U923 ( .A1(n1229), .A2(n1121), .ZN(n1228) );
NAND2_X1 U924 ( .A1(n1121), .A2(n1229), .ZN(n1226) );
XNOR2_X1 U925 ( .A(n1230), .B(n1197), .ZN(n1229) );
AND2_X1 U926 ( .A1(G224), .A2(n1101), .ZN(n1197) );
NAND2_X1 U927 ( .A1(n1231), .A2(KEYINPUT41), .ZN(n1230) );
XNOR2_X1 U928 ( .A(G125), .B(n1198), .ZN(n1231) );
XOR2_X1 U929 ( .A(n1232), .B(n1233), .Z(n1121) );
XOR2_X1 U930 ( .A(n1234), .B(n1235), .Z(n1233) );
XNOR2_X1 U931 ( .A(G110), .B(G119), .ZN(n1235) );
NAND3_X1 U932 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1234) );
NAND2_X1 U933 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
OR3_X1 U934 ( .A1(n1240), .A2(n1239), .A3(KEYINPUT63), .ZN(n1237) );
XNOR2_X1 U935 ( .A(n1241), .B(KEYINPUT27), .ZN(n1239) );
NAND2_X1 U936 ( .A1(KEYINPUT25), .A2(n1142), .ZN(n1240) );
NAND2_X1 U937 ( .A1(n1242), .A2(KEYINPUT63), .ZN(n1236) );
XNOR2_X1 U938 ( .A(n1243), .B(n1244), .ZN(n1232) );
NOR2_X1 U939 ( .A1(G113), .A2(KEYINPUT40), .ZN(n1244) );
NAND2_X1 U940 ( .A1(n1211), .A2(n1245), .ZN(n1035) );
NAND2_X1 U941 ( .A1(n1210), .A2(n1120), .ZN(n1245) );
XOR2_X1 U942 ( .A(G898), .B(KEYINPUT55), .Z(n1120) );
NOR3_X1 U943 ( .A1(n1101), .A2(n1048), .A3(n1224), .ZN(n1210) );
INV_X1 U944 ( .A(n1063), .ZN(n1048) );
NAND3_X1 U945 ( .A1(G952), .A2(n1063), .A3(n1246), .ZN(n1211) );
XNOR2_X1 U946 ( .A(G953), .B(KEYINPUT43), .ZN(n1246) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1063) );
NAND2_X1 U948 ( .A1(n1247), .A2(n1248), .ZN(n1034) );
OR3_X1 U949 ( .A1(n1080), .A2(n1082), .A3(KEYINPUT51), .ZN(n1248) );
INV_X1 U950 ( .A(n1249), .ZN(n1082) );
NAND2_X1 U951 ( .A1(KEYINPUT51), .A2(n1060), .ZN(n1247) );
INV_X1 U952 ( .A(n1051), .ZN(n1060) );
NAND2_X1 U953 ( .A1(n1080), .A2(n1249), .ZN(n1051) );
NAND2_X1 U954 ( .A1(G221), .A2(n1250), .ZN(n1249) );
XNOR2_X1 U955 ( .A(n1251), .B(n1151), .ZN(n1080) );
INV_X1 U956 ( .A(G469), .ZN(n1151) );
NAND2_X1 U957 ( .A1(n1252), .A2(n1224), .ZN(n1251) );
XOR2_X1 U958 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U959 ( .A(n1149), .B(n1110), .ZN(n1254) );
XOR2_X1 U960 ( .A(G128), .B(n1255), .Z(n1110) );
NOR2_X1 U961 ( .A1(KEYINPUT38), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U962 ( .A(G143), .B(G146), .ZN(n1256) );
XNOR2_X1 U963 ( .A(n1111), .B(KEYINPUT11), .ZN(n1149) );
XNOR2_X1 U964 ( .A(n1157), .B(n1257), .ZN(n1253) );
XNOR2_X1 U965 ( .A(KEYINPUT52), .B(n1258), .ZN(n1257) );
NOR2_X1 U966 ( .A1(KEYINPUT16), .A2(n1259), .ZN(n1258) );
XOR2_X1 U967 ( .A(n1260), .B(n1159), .Z(n1259) );
XNOR2_X1 U968 ( .A(G140), .B(n1261), .ZN(n1159) );
AND2_X1 U969 ( .A1(n1101), .A2(G227), .ZN(n1261) );
NAND2_X1 U970 ( .A1(KEYINPUT24), .A2(n1221), .ZN(n1260) );
XNOR2_X1 U971 ( .A(n1241), .B(n1262), .ZN(n1157) );
XNOR2_X1 U972 ( .A(KEYINPUT33), .B(n1142), .ZN(n1262) );
INV_X1 U973 ( .A(n1242), .ZN(n1142) );
XNOR2_X1 U974 ( .A(G104), .B(G107), .ZN(n1241) );
XOR2_X1 U975 ( .A(n1263), .B(n1092), .Z(n1212) );
NAND2_X1 U976 ( .A1(n1264), .A2(n1224), .ZN(n1092) );
XNOR2_X1 U977 ( .A(n1143), .B(n1265), .ZN(n1264) );
NOR2_X1 U978 ( .A1(KEYINPUT17), .A2(n1266), .ZN(n1265) );
XNOR2_X1 U979 ( .A(n1242), .B(n1267), .ZN(n1266) );
NOR2_X1 U980 ( .A1(KEYINPUT50), .A2(n1144), .ZN(n1267) );
NAND2_X1 U981 ( .A1(G210), .A2(n1268), .ZN(n1144) );
XOR2_X1 U982 ( .A(G101), .B(KEYINPUT59), .Z(n1242) );
XNOR2_X1 U983 ( .A(n1269), .B(n1270), .ZN(n1143) );
XNOR2_X1 U984 ( .A(n1198), .B(n1271), .ZN(n1270) );
INV_X1 U985 ( .A(n1111), .ZN(n1271) );
XOR2_X1 U986 ( .A(G131), .B(n1272), .Z(n1111) );
XNOR2_X1 U987 ( .A(n1273), .B(G134), .ZN(n1272) );
XNOR2_X1 U988 ( .A(n1274), .B(n1275), .ZN(n1198) );
NOR2_X1 U989 ( .A1(G146), .A2(KEYINPUT45), .ZN(n1275) );
XNOR2_X1 U990 ( .A(G143), .B(n1276), .ZN(n1274) );
NOR2_X1 U991 ( .A1(G128), .A2(KEYINPUT22), .ZN(n1276) );
XOR2_X1 U992 ( .A(n1277), .B(n1278), .Z(n1269) );
XOR2_X1 U993 ( .A(G119), .B(G113), .Z(n1278) );
NAND2_X1 U994 ( .A1(KEYINPUT47), .A2(n1217), .ZN(n1277) );
NAND2_X1 U995 ( .A1(KEYINPUT21), .A2(n1093), .ZN(n1263) );
INV_X1 U996 ( .A(G472), .ZN(n1093) );
INV_X1 U997 ( .A(n1056), .ZN(n1176) );
NAND2_X1 U998 ( .A1(n1059), .A2(n1091), .ZN(n1056) );
XOR2_X1 U999 ( .A(n1279), .B(n1128), .Z(n1091) );
NAND2_X1 U1000 ( .A1(G217), .A2(n1250), .ZN(n1128) );
NAND2_X1 U1001 ( .A1(n1280), .A2(n1224), .ZN(n1250) );
XOR2_X1 U1002 ( .A(KEYINPUT60), .B(G234), .Z(n1280) );
OR2_X1 U1003 ( .A1(n1127), .A2(G902), .ZN(n1279) );
XNOR2_X1 U1004 ( .A(n1281), .B(n1282), .ZN(n1127) );
XOR2_X1 U1005 ( .A(n1283), .B(n1284), .Z(n1282) );
NAND2_X1 U1006 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U1007 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U1008 ( .A(KEYINPUT3), .B(G125), .Z(n1288) );
XNOR2_X1 U1009 ( .A(KEYINPUT54), .B(n1289), .ZN(n1287) );
NAND2_X1 U1010 ( .A1(n1290), .A2(n1291), .ZN(n1285) );
XNOR2_X1 U1011 ( .A(KEYINPUT3), .B(G125), .ZN(n1291) );
XNOR2_X1 U1012 ( .A(G140), .B(KEYINPUT19), .ZN(n1290) );
NAND3_X1 U1013 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1283) );
OR2_X1 U1014 ( .A1(n1295), .A2(G119), .ZN(n1294) );
NAND2_X1 U1015 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
INV_X1 U1016 ( .A(KEYINPUT56), .ZN(n1297) );
NAND2_X1 U1017 ( .A1(n1298), .A2(n1295), .ZN(n1296) );
XNOR2_X1 U1018 ( .A(KEYINPUT9), .B(G119), .ZN(n1298) );
NAND2_X1 U1019 ( .A1(KEYINPUT56), .A2(n1299), .ZN(n1292) );
NAND2_X1 U1020 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
OR2_X1 U1021 ( .A1(G119), .A2(KEYINPUT9), .ZN(n1301) );
NAND3_X1 U1022 ( .A1(G119), .A2(n1295), .A3(KEYINPUT9), .ZN(n1300) );
INV_X1 U1023 ( .A(G128), .ZN(n1295) );
XOR2_X1 U1024 ( .A(n1302), .B(n1303), .Z(n1281) );
XNOR2_X1 U1025 ( .A(G146), .B(n1221), .ZN(n1303) );
NAND2_X1 U1026 ( .A1(n1304), .A2(n1305), .ZN(n1302) );
NAND4_X1 U1027 ( .A1(G221), .A2(G234), .A3(G137), .A4(n1306), .ZN(n1305) );
XOR2_X1 U1028 ( .A(n1307), .B(KEYINPUT15), .Z(n1304) );
NAND2_X1 U1029 ( .A1(n1273), .A2(n1308), .ZN(n1307) );
NAND3_X1 U1030 ( .A1(G234), .A2(n1306), .A3(G221), .ZN(n1308) );
XNOR2_X1 U1031 ( .A(n1101), .B(KEYINPUT7), .ZN(n1306) );
INV_X1 U1032 ( .A(G137), .ZN(n1273) );
NOR2_X1 U1033 ( .A1(n1087), .A2(n1201), .ZN(n1059) );
XNOR2_X1 U1034 ( .A(G478), .B(n1309), .ZN(n1201) );
NOR2_X1 U1035 ( .A1(n1089), .A2(KEYINPUT4), .ZN(n1309) );
AND2_X1 U1036 ( .A1(n1131), .A2(n1224), .ZN(n1089) );
INV_X1 U1037 ( .A(G902), .ZN(n1224) );
XOR2_X1 U1038 ( .A(n1310), .B(n1311), .Z(n1131) );
XOR2_X1 U1039 ( .A(G107), .B(n1312), .Z(n1311) );
NOR2_X1 U1040 ( .A1(KEYINPUT6), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1041 ( .A(n1314), .B(n1315), .Z(n1313) );
NOR2_X1 U1042 ( .A1(KEYINPUT46), .A2(G128), .ZN(n1315) );
XNOR2_X1 U1043 ( .A(G134), .B(G143), .ZN(n1314) );
XOR2_X1 U1044 ( .A(n1316), .B(n1243), .Z(n1310) );
XNOR2_X1 U1045 ( .A(n1217), .B(G122), .ZN(n1243) );
INV_X1 U1046 ( .A(G116), .ZN(n1217) );
NAND3_X1 U1047 ( .A1(G234), .A2(n1101), .A3(G217), .ZN(n1316) );
INV_X1 U1048 ( .A(G953), .ZN(n1101) );
XOR2_X1 U1049 ( .A(n1317), .B(n1137), .Z(n1087) );
INV_X1 U1050 ( .A(G475), .ZN(n1137) );
OR2_X1 U1051 ( .A1(n1136), .A2(G902), .ZN(n1317) );
XNOR2_X1 U1052 ( .A(n1318), .B(n1319), .ZN(n1136) );
XOR2_X1 U1053 ( .A(G113), .B(n1320), .Z(n1319) );
XOR2_X1 U1054 ( .A(G146), .B(G122), .Z(n1320) );
XOR2_X1 U1055 ( .A(n1321), .B(n1107), .Z(n1318) );
XNOR2_X1 U1056 ( .A(n1289), .B(G125), .ZN(n1107) );
INV_X1 U1057 ( .A(G140), .ZN(n1289) );
XOR2_X1 U1058 ( .A(n1322), .B(G104), .Z(n1321) );
NAND2_X1 U1059 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
OR2_X1 U1060 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1061 ( .A(n1327), .B(KEYINPUT37), .Z(n1323) );
NAND2_X1 U1062 ( .A1(n1325), .A2(n1326), .ZN(n1327) );
INV_X1 U1063 ( .A(G131), .ZN(n1326) );
XOR2_X1 U1064 ( .A(n1328), .B(n1329), .Z(n1325) );
INV_X1 U1065 ( .A(G143), .ZN(n1329) );
NAND2_X1 U1066 ( .A1(G214), .A2(n1268), .ZN(n1328) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1268) );
INV_X1 U1068 ( .A(G110), .ZN(n1221) );
endmodule


