//Key = 0010101101010000011001010110111101100100101010000000010001001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368;

NAND3_X1 U746 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(G9) );
OR2_X1 U747 ( .A1(n1036), .A2(KEYINPUT11), .ZN(n1035) );
NAND3_X1 U748 ( .A1(KEYINPUT11), .A2(n1036), .A3(n1037), .ZN(n1034) );
NAND2_X1 U749 ( .A1(G107), .A2(n1038), .ZN(n1033) );
NAND2_X1 U750 ( .A1(n1039), .A2(KEYINPUT11), .ZN(n1038) );
XNOR2_X1 U751 ( .A(n1036), .B(KEYINPUT61), .ZN(n1039) );
INV_X1 U752 ( .A(n1040), .ZN(n1036) );
NOR2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1049) );
XOR2_X1 U759 ( .A(KEYINPUT19), .B(n1055), .Z(n1044) );
NOR3_X1 U760 ( .A1(n1056), .A2(n1048), .A3(n1057), .ZN(n1055) );
NAND3_X1 U761 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1048) );
NAND3_X1 U762 ( .A1(G214), .A2(n1061), .A3(n1062), .ZN(n1056) );
NAND3_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1043) );
NAND4_X1 U764 ( .A1(n1060), .A2(n1066), .A3(n1062), .A4(n1067), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U766 ( .A1(n1059), .A2(n1070), .ZN(n1069) );
OR2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U768 ( .A1(n1058), .A2(n1073), .ZN(n1068) );
NAND3_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
OR3_X1 U770 ( .A1(n1077), .A2(n1078), .A3(KEYINPUT38), .ZN(n1075) );
NAND2_X1 U771 ( .A1(KEYINPUT38), .A2(n1059), .ZN(n1074) );
INV_X1 U772 ( .A(n1079), .ZN(n1060) );
NOR3_X1 U773 ( .A1(n1080), .A2(G953), .A3(G952), .ZN(n1041) );
INV_X1 U774 ( .A(n1063), .ZN(n1080) );
NAND4_X1 U775 ( .A1(n1059), .A2(n1066), .A3(n1081), .A4(n1082), .ZN(n1063) );
NOR3_X1 U776 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
XNOR2_X1 U777 ( .A(n1086), .B(KEYINPUT44), .ZN(n1085) );
XOR2_X1 U778 ( .A(n1087), .B(n1088), .Z(n1084) );
NOR2_X1 U779 ( .A1(n1089), .A2(KEYINPUT36), .ZN(n1088) );
XNOR2_X1 U780 ( .A(G478), .B(n1090), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1091), .B(n1092), .Z(G72) );
XOR2_X1 U782 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U783 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U784 ( .A(n1097), .B(n1098), .Z(n1096) );
XNOR2_X1 U785 ( .A(n1099), .B(n1100), .ZN(n1098) );
NOR2_X1 U786 ( .A1(KEYINPUT46), .A2(n1101), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
XOR2_X1 U788 ( .A(n1104), .B(G140), .Z(n1097) );
XNOR2_X1 U789 ( .A(KEYINPUT63), .B(KEYINPUT60), .ZN(n1104) );
NOR2_X1 U790 ( .A1(G900), .A2(n1105), .ZN(n1095) );
NOR2_X1 U791 ( .A1(G953), .A2(n1106), .ZN(n1093) );
NOR3_X1 U792 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
XNOR2_X1 U793 ( .A(n1110), .B(KEYINPUT1), .ZN(n1108) );
XNOR2_X1 U794 ( .A(KEYINPUT51), .B(n1111), .ZN(n1107) );
NOR2_X1 U795 ( .A1(n1112), .A2(n1064), .ZN(n1091) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1115), .B(n1116), .Z(G69) );
XOR2_X1 U798 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U799 ( .A1(n1119), .A2(G953), .ZN(n1118) );
NOR2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
NOR2_X1 U801 ( .A1(G898), .A2(n1105), .ZN(n1120) );
NOR2_X1 U802 ( .A1(n1122), .A2(n1064), .ZN(n1115) );
NOR2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR3_X1 U804 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(G66) );
NOR3_X1 U805 ( .A1(n1128), .A2(G953), .A3(G952), .ZN(n1127) );
AND2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
INV_X1 U807 ( .A(KEYINPUT13), .ZN(n1128) );
NOR2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1125) );
XOR2_X1 U809 ( .A(KEYINPUT55), .B(n1132), .Z(n1131) );
NOR2_X1 U810 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
AND2_X1 U811 ( .A1(n1134), .A2(n1133), .ZN(n1130) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1089), .ZN(n1134) );
NOR2_X1 U813 ( .A1(n1129), .A2(n1136), .ZN(G63) );
NOR3_X1 U814 ( .A1(n1090), .A2(n1137), .A3(n1138), .ZN(n1136) );
AND2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR3_X1 U816 ( .A1(n1140), .A2(n1141), .A3(n1139), .ZN(n1137) );
NAND2_X1 U817 ( .A1(n1142), .A2(G478), .ZN(n1139) );
XOR2_X1 U818 ( .A(n1046), .B(KEYINPUT47), .Z(n1142) );
NOR2_X1 U819 ( .A1(n1129), .A2(n1143), .ZN(G60) );
XOR2_X1 U820 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U821 ( .A(KEYINPUT7), .B(n1146), .Z(n1145) );
AND2_X1 U822 ( .A1(G475), .A2(n1135), .ZN(n1146) );
XNOR2_X1 U823 ( .A(n1147), .B(n1148), .ZN(G6) );
NOR2_X1 U824 ( .A1(KEYINPUT41), .A2(n1149), .ZN(n1148) );
INV_X1 U825 ( .A(G104), .ZN(n1149) );
NOR2_X1 U826 ( .A1(n1129), .A2(n1150), .ZN(G57) );
XOR2_X1 U827 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U828 ( .A(KEYINPUT57), .B(n1153), .Z(n1152) );
AND2_X1 U829 ( .A1(G472), .A2(n1135), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1129), .A2(n1154), .ZN(G54) );
XOR2_X1 U831 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U832 ( .A(n1157), .B(n1158), .ZN(n1156) );
XOR2_X1 U833 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U834 ( .A(n1161), .B(n1162), .Z(n1155) );
XOR2_X1 U835 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U836 ( .A1(KEYINPUT43), .A2(n1102), .ZN(n1163) );
XOR2_X1 U837 ( .A(KEYINPUT33), .B(n1165), .Z(n1161) );
AND2_X1 U838 ( .A1(G469), .A2(n1135), .ZN(n1165) );
NOR2_X1 U839 ( .A1(n1129), .A2(n1166), .ZN(G51) );
XOR2_X1 U840 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND3_X1 U841 ( .A1(n1135), .A2(n1169), .A3(KEYINPUT9), .ZN(n1167) );
AND2_X1 U842 ( .A1(G902), .A2(n1046), .ZN(n1135) );
NAND4_X1 U843 ( .A1(n1110), .A2(n1119), .A3(n1170), .A4(n1111), .ZN(n1046) );
NAND3_X1 U844 ( .A1(n1171), .A2(n1172), .A3(n1071), .ZN(n1111) );
INV_X1 U845 ( .A(n1109), .ZN(n1170) );
NAND3_X1 U846 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1109) );
NAND2_X1 U847 ( .A1(n1176), .A2(n1171), .ZN(n1175) );
AND4_X1 U848 ( .A1(n1177), .A2(n1178), .A3(n1040), .A4(n1179), .ZN(n1119) );
NOR4_X1 U849 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
NOR2_X1 U850 ( .A1(n1147), .A2(n1184), .ZN(n1183) );
INV_X1 U851 ( .A(KEYINPUT53), .ZN(n1184) );
NAND2_X1 U852 ( .A1(n1185), .A2(n1186), .ZN(n1147) );
NOR2_X1 U853 ( .A1(n1053), .A2(n1187), .ZN(n1182) );
NOR2_X1 U854 ( .A1(n1172), .A2(n1188), .ZN(n1053) );
NOR3_X1 U855 ( .A1(n1186), .A2(KEYINPUT34), .A3(n1189), .ZN(n1181) );
NOR2_X1 U856 ( .A1(n1190), .A2(n1051), .ZN(n1180) );
NOR3_X1 U857 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
NOR2_X1 U858 ( .A1(KEYINPUT53), .A2(n1185), .ZN(n1193) );
NOR4_X1 U859 ( .A1(n1194), .A2(n1052), .A3(n1076), .A4(n1195), .ZN(n1185) );
NOR3_X1 U860 ( .A1(n1196), .A2(n1195), .A3(n1197), .ZN(n1192) );
NOR2_X1 U861 ( .A1(n1189), .A2(n1198), .ZN(n1191) );
INV_X1 U862 ( .A(KEYINPUT34), .ZN(n1198) );
NAND4_X1 U863 ( .A1(n1062), .A2(n1072), .A3(n1199), .A4(n1200), .ZN(n1040) );
NOR2_X1 U864 ( .A1(n1195), .A2(n1051), .ZN(n1199) );
NOR4_X1 U865 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1110) );
NOR2_X1 U866 ( .A1(n1064), .A2(G952), .ZN(n1129) );
XNOR2_X1 U867 ( .A(n1205), .B(n1173), .ZN(G48) );
NAND3_X1 U868 ( .A1(n1071), .A2(n1206), .A3(n1207), .ZN(n1173) );
NAND2_X1 U869 ( .A1(KEYINPUT18), .A2(n1208), .ZN(n1205) );
XNOR2_X1 U870 ( .A(G143), .B(n1174), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1207), .A2(n1188), .A3(n1209), .A4(n1083), .ZN(n1174) );
XOR2_X1 U872 ( .A(G140), .B(n1210), .Z(G42) );
NOR3_X1 U873 ( .A1(n1211), .A2(n1212), .A3(n1054), .ZN(n1210) );
INV_X1 U874 ( .A(n1066), .ZN(n1054) );
XNOR2_X1 U875 ( .A(n1200), .B(KEYINPUT10), .ZN(n1212) );
NAND2_X1 U876 ( .A1(n1213), .A2(n1214), .ZN(G39) );
NAND4_X1 U877 ( .A1(n1176), .A2(n1171), .A3(n1215), .A4(n1216), .ZN(n1214) );
NAND2_X1 U878 ( .A1(G137), .A2(n1217), .ZN(n1216) );
NAND2_X1 U879 ( .A1(KEYINPUT24), .A2(n1218), .ZN(n1215) );
NAND3_X1 U880 ( .A1(n1219), .A2(n1217), .A3(G137), .ZN(n1213) );
INV_X1 U881 ( .A(KEYINPUT15), .ZN(n1217) );
NAND3_X1 U882 ( .A1(n1171), .A2(n1220), .A3(n1176), .ZN(n1219) );
INV_X1 U883 ( .A(n1196), .ZN(n1176) );
INV_X1 U884 ( .A(KEYINPUT24), .ZN(n1220) );
XOR2_X1 U885 ( .A(G134), .B(n1201), .Z(G36) );
AND3_X1 U886 ( .A1(n1171), .A2(n1072), .A3(n1188), .ZN(n1201) );
XOR2_X1 U887 ( .A(G131), .B(n1202), .Z(G33) );
AND3_X1 U888 ( .A1(n1071), .A2(n1171), .A3(n1188), .ZN(n1202) );
AND3_X1 U889 ( .A1(n1200), .A2(n1221), .A3(n1066), .ZN(n1171) );
NOR2_X1 U890 ( .A1(n1057), .A2(n1222), .ZN(n1066) );
AND2_X1 U891 ( .A1(G214), .A2(n1061), .ZN(n1222) );
XNOR2_X1 U892 ( .A(G128), .B(n1223), .ZN(G30) );
NOR2_X1 U893 ( .A1(n1203), .A2(KEYINPUT52), .ZN(n1223) );
AND3_X1 U894 ( .A1(n1072), .A2(n1206), .A3(n1207), .ZN(n1203) );
AND3_X1 U895 ( .A1(n1186), .A2(n1221), .A3(n1200), .ZN(n1207) );
XOR2_X1 U896 ( .A(G101), .B(n1224), .Z(G3) );
NOR2_X1 U897 ( .A1(n1225), .A2(n1187), .ZN(n1224) );
XNOR2_X1 U898 ( .A(n1099), .B(n1204), .ZN(G27) );
NOR3_X1 U899 ( .A1(n1197), .A2(n1051), .A3(n1211), .ZN(n1204) );
NAND3_X1 U900 ( .A1(n1172), .A2(n1221), .A3(n1071), .ZN(n1211) );
NAND2_X1 U901 ( .A1(n1079), .A2(n1226), .ZN(n1221) );
NAND2_X1 U902 ( .A1(n1227), .A2(n1114), .ZN(n1226) );
INV_X1 U903 ( .A(G900), .ZN(n1114) );
XOR2_X1 U904 ( .A(G122), .B(n1228), .Z(G24) );
NOR2_X1 U905 ( .A1(n1229), .A2(n1051), .ZN(n1228) );
XOR2_X1 U906 ( .A(n1189), .B(KEYINPUT62), .Z(n1229) );
NAND4_X1 U907 ( .A1(n1083), .A2(n1230), .A3(n1209), .A4(n1231), .ZN(n1189) );
NOR2_X1 U908 ( .A1(n1052), .A2(n1197), .ZN(n1231) );
INV_X1 U909 ( .A(n1062), .ZN(n1052) );
XNOR2_X1 U910 ( .A(G119), .B(n1232), .ZN(G21) );
NAND2_X1 U911 ( .A1(n1186), .A2(n1233), .ZN(n1232) );
XOR2_X1 U912 ( .A(KEYINPUT50), .B(n1234), .Z(n1233) );
NOR3_X1 U913 ( .A1(n1196), .A2(n1195), .A3(n1235), .ZN(n1234) );
XNOR2_X1 U914 ( .A(n1059), .B(KEYINPUT16), .ZN(n1235) );
INV_X1 U915 ( .A(n1197), .ZN(n1059) );
NAND2_X1 U916 ( .A1(n1058), .A2(n1206), .ZN(n1196) );
NAND2_X1 U917 ( .A1(n1236), .A2(n1237), .ZN(n1206) );
NAND3_X1 U918 ( .A1(n1238), .A2(n1086), .A3(n1239), .ZN(n1237) );
INV_X1 U919 ( .A(KEYINPUT12), .ZN(n1239) );
NAND2_X1 U920 ( .A1(KEYINPUT12), .A2(n1188), .ZN(n1236) );
INV_X1 U921 ( .A(n1225), .ZN(n1188) );
XNOR2_X1 U922 ( .A(G116), .B(n1177), .ZN(G18) );
NAND2_X1 U923 ( .A1(n1240), .A2(n1072), .ZN(n1177) );
NOR2_X1 U924 ( .A1(n1083), .A2(n1241), .ZN(n1072) );
NAND3_X1 U925 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(G15) );
NAND2_X1 U926 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U927 ( .A1(KEYINPUT54), .A2(n1247), .ZN(n1243) );
NAND2_X1 U928 ( .A1(n1248), .A2(G113), .ZN(n1247) );
XNOR2_X1 U929 ( .A(KEYINPUT5), .B(n1245), .ZN(n1248) );
NAND2_X1 U930 ( .A1(n1249), .A2(n1250), .ZN(n1242) );
INV_X1 U931 ( .A(KEYINPUT54), .ZN(n1250) );
NAND2_X1 U932 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
OR3_X1 U933 ( .A1(n1246), .A2(n1245), .A3(KEYINPUT5), .ZN(n1252) );
NAND2_X1 U934 ( .A1(KEYINPUT5), .A2(n1245), .ZN(n1251) );
INV_X1 U935 ( .A(n1178), .ZN(n1245) );
NAND2_X1 U936 ( .A1(n1240), .A2(n1071), .ZN(n1178) );
INV_X1 U937 ( .A(n1194), .ZN(n1071) );
NAND2_X1 U938 ( .A1(n1241), .A2(n1083), .ZN(n1194) );
NOR4_X1 U939 ( .A1(n1225), .A2(n1197), .A3(n1051), .A4(n1195), .ZN(n1240) );
INV_X1 U940 ( .A(n1230), .ZN(n1195) );
NAND2_X1 U941 ( .A1(n1253), .A2(n1077), .ZN(n1197) );
NAND2_X1 U942 ( .A1(n1254), .A2(n1086), .ZN(n1225) );
XNOR2_X1 U943 ( .A(n1255), .B(n1256), .ZN(G12) );
NOR2_X1 U944 ( .A1(n1257), .A2(n1187), .ZN(n1256) );
NAND4_X1 U945 ( .A1(n1058), .A2(n1200), .A3(n1186), .A4(n1230), .ZN(n1187) );
NAND2_X1 U946 ( .A1(n1079), .A2(n1258), .ZN(n1230) );
NAND2_X1 U947 ( .A1(n1227), .A2(n1124), .ZN(n1258) );
INV_X1 U948 ( .A(G898), .ZN(n1124) );
NOR3_X1 U949 ( .A1(n1105), .A2(n1259), .A3(n1141), .ZN(n1227) );
INV_X1 U950 ( .A(n1260), .ZN(n1259) );
XOR2_X1 U951 ( .A(G953), .B(KEYINPUT6), .Z(n1105) );
NAND3_X1 U952 ( .A1(n1260), .A2(n1064), .A3(n1261), .ZN(n1079) );
XNOR2_X1 U953 ( .A(G952), .B(KEYINPUT37), .ZN(n1261) );
NAND2_X1 U954 ( .A1(G237), .A2(G234), .ZN(n1260) );
INV_X1 U955 ( .A(n1051), .ZN(n1186) );
NAND2_X1 U956 ( .A1(n1057), .A2(n1262), .ZN(n1051) );
NAND2_X1 U957 ( .A1(G214), .A2(n1061), .ZN(n1262) );
XNOR2_X1 U958 ( .A(n1263), .B(n1169), .ZN(n1057) );
AND2_X1 U959 ( .A1(G210), .A2(n1061), .ZN(n1169) );
NAND2_X1 U960 ( .A1(n1264), .A2(n1141), .ZN(n1061) );
XOR2_X1 U961 ( .A(KEYINPUT2), .B(G237), .Z(n1264) );
NAND2_X1 U962 ( .A1(n1168), .A2(n1141), .ZN(n1263) );
XNOR2_X1 U963 ( .A(n1265), .B(n1266), .ZN(n1168) );
XNOR2_X1 U964 ( .A(G125), .B(n1267), .ZN(n1266) );
XNOR2_X1 U965 ( .A(n1121), .B(n1268), .ZN(n1265) );
NOR2_X1 U966 ( .A1(G953), .A2(n1123), .ZN(n1268) );
INV_X1 U967 ( .A(G224), .ZN(n1123) );
XNOR2_X1 U968 ( .A(n1269), .B(n1270), .ZN(n1121) );
XOR2_X1 U969 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U970 ( .A(n1273), .B(G116), .Z(n1272) );
NAND2_X1 U971 ( .A1(KEYINPUT42), .A2(n1246), .ZN(n1273) );
XNOR2_X1 U972 ( .A(G119), .B(KEYINPUT29), .ZN(n1271) );
XOR2_X1 U973 ( .A(n1274), .B(n1164), .Z(n1269) );
XNOR2_X1 U974 ( .A(n1255), .B(n1275), .ZN(n1164) );
XOR2_X1 U975 ( .A(n1276), .B(n1277), .Z(n1274) );
NAND2_X1 U976 ( .A1(KEYINPUT25), .A2(n1160), .ZN(n1276) );
INV_X1 U977 ( .A(n1076), .ZN(n1200) );
NAND2_X1 U978 ( .A1(n1078), .A2(n1077), .ZN(n1076) );
NAND2_X1 U979 ( .A1(G221), .A2(n1278), .ZN(n1077) );
INV_X1 U980 ( .A(n1253), .ZN(n1078) );
XOR2_X1 U981 ( .A(n1279), .B(G469), .Z(n1253) );
NAND2_X1 U982 ( .A1(n1280), .A2(n1141), .ZN(n1279) );
XOR2_X1 U983 ( .A(n1159), .B(n1281), .Z(n1280) );
XOR2_X1 U984 ( .A(n1282), .B(n1283), .Z(n1281) );
NOR2_X1 U985 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U986 ( .A(n1286), .B(KEYINPUT4), .Z(n1285) );
NAND2_X1 U987 ( .A1(n1287), .A2(n1102), .ZN(n1286) );
NOR2_X1 U988 ( .A1(n1287), .A2(n1102), .ZN(n1284) );
NAND2_X1 U989 ( .A1(n1288), .A2(n1289), .ZN(n1102) );
NAND2_X1 U990 ( .A1(n1290), .A2(n1208), .ZN(n1289) );
XOR2_X1 U991 ( .A(KEYINPUT30), .B(n1291), .Z(n1290) );
XOR2_X1 U992 ( .A(n1275), .B(n1160), .Z(n1287) );
XNOR2_X1 U993 ( .A(G104), .B(KEYINPUT35), .ZN(n1160) );
XNOR2_X1 U994 ( .A(G101), .B(n1037), .ZN(n1275) );
INV_X1 U995 ( .A(G107), .ZN(n1037) );
NOR2_X1 U996 ( .A1(KEYINPUT27), .A2(n1292), .ZN(n1282) );
XOR2_X1 U997 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U998 ( .A(G110), .B(n1157), .ZN(n1294) );
XOR2_X1 U999 ( .A(G140), .B(n1295), .Z(n1157) );
NOR2_X1 U1000 ( .A1(G953), .A2(n1113), .ZN(n1295) );
INV_X1 U1001 ( .A(G227), .ZN(n1113) );
XNOR2_X1 U1002 ( .A(KEYINPUT48), .B(KEYINPUT23), .ZN(n1293) );
NOR2_X1 U1003 ( .A1(n1083), .A2(n1209), .ZN(n1058) );
INV_X1 U1004 ( .A(n1241), .ZN(n1209) );
XNOR2_X1 U1005 ( .A(n1296), .B(n1090), .ZN(n1241) );
AND2_X1 U1006 ( .A1(n1140), .A2(n1141), .ZN(n1090) );
XNOR2_X1 U1007 ( .A(n1297), .B(n1298), .ZN(n1140) );
XOR2_X1 U1008 ( .A(n1299), .B(n1300), .Z(n1298) );
XOR2_X1 U1009 ( .A(n1301), .B(n1302), .Z(n1300) );
AND3_X1 U1010 ( .A1(G217), .A2(n1064), .A3(G234), .ZN(n1302) );
INV_X1 U1011 ( .A(G953), .ZN(n1064) );
NOR2_X1 U1012 ( .A1(KEYINPUT39), .A2(n1303), .ZN(n1301) );
XNOR2_X1 U1013 ( .A(n1304), .B(G107), .ZN(n1299) );
XNOR2_X1 U1014 ( .A(n1277), .B(n1305), .ZN(n1297) );
XNOR2_X1 U1015 ( .A(n1306), .B(n1307), .ZN(n1305) );
NOR2_X1 U1016 ( .A1(G116), .A2(KEYINPUT58), .ZN(n1307) );
NAND2_X1 U1017 ( .A1(KEYINPUT26), .A2(G134), .ZN(n1306) );
NAND2_X1 U1018 ( .A1(KEYINPUT21), .A2(n1308), .ZN(n1296) );
INV_X1 U1019 ( .A(G478), .ZN(n1308) );
XNOR2_X1 U1020 ( .A(n1309), .B(G475), .ZN(n1083) );
NAND2_X1 U1021 ( .A1(n1144), .A2(n1141), .ZN(n1309) );
XOR2_X1 U1022 ( .A(n1310), .B(n1311), .Z(n1144) );
XNOR2_X1 U1023 ( .A(n1246), .B(G104), .ZN(n1311) );
XNOR2_X1 U1024 ( .A(n1277), .B(n1312), .ZN(n1310) );
NOR2_X1 U1025 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1026 ( .A(KEYINPUT8), .B(n1315), .Z(n1314) );
NOR2_X1 U1027 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
AND2_X1 U1028 ( .A1(n1317), .A2(n1316), .ZN(n1313) );
NAND2_X1 U1029 ( .A1(n1318), .A2(n1319), .ZN(n1316) );
NAND2_X1 U1030 ( .A1(n1320), .A2(n1099), .ZN(n1319) );
INV_X1 U1031 ( .A(G125), .ZN(n1099) );
NAND2_X1 U1032 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NAND2_X1 U1033 ( .A1(n1323), .A2(G125), .ZN(n1318) );
XNOR2_X1 U1034 ( .A(G146), .B(n1324), .ZN(n1323) );
XNOR2_X1 U1035 ( .A(n1325), .B(n1326), .ZN(n1317) );
XNOR2_X1 U1036 ( .A(n1304), .B(G131), .ZN(n1326) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1327), .ZN(n1325) );
XOR2_X1 U1038 ( .A(G122), .B(KEYINPUT40), .Z(n1277) );
XNOR2_X1 U1039 ( .A(KEYINPUT14), .B(n1172), .ZN(n1257) );
NAND2_X1 U1040 ( .A1(n1328), .A2(n1329), .ZN(n1172) );
OR3_X1 U1041 ( .A1(n1254), .A2(n1086), .A3(KEYINPUT12), .ZN(n1329) );
INV_X1 U1042 ( .A(n1238), .ZN(n1254) );
NAND2_X1 U1043 ( .A1(KEYINPUT12), .A2(n1062), .ZN(n1328) );
NOR2_X1 U1044 ( .A1(n1086), .A2(n1238), .ZN(n1062) );
XNOR2_X1 U1045 ( .A(n1087), .B(n1089), .ZN(n1238) );
AND2_X1 U1046 ( .A1(G217), .A2(n1278), .ZN(n1089) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1141), .ZN(n1278) );
NAND2_X1 U1048 ( .A1(n1133), .A2(n1141), .ZN(n1087) );
XNOR2_X1 U1049 ( .A(n1330), .B(n1331), .ZN(n1133) );
XNOR2_X1 U1050 ( .A(n1255), .B(n1332), .ZN(n1331) );
XNOR2_X1 U1051 ( .A(n1303), .B(G119), .ZN(n1332) );
INV_X1 U1052 ( .A(G128), .ZN(n1303) );
XOR2_X1 U1053 ( .A(n1333), .B(n1334), .Z(n1330) );
NOR3_X1 U1054 ( .A1(n1335), .A2(KEYINPUT0), .A3(n1336), .ZN(n1334) );
NOR4_X1 U1055 ( .A1(G953), .A2(n1337), .A3(n1338), .A4(n1339), .ZN(n1336) );
XNOR2_X1 U1056 ( .A(G137), .B(KEYINPUT32), .ZN(n1337) );
NOR2_X1 U1057 ( .A1(n1340), .A2(G137), .ZN(n1335) );
NOR3_X1 U1058 ( .A1(n1339), .A2(G953), .A3(n1338), .ZN(n1340) );
INV_X1 U1059 ( .A(G234), .ZN(n1338) );
INV_X1 U1060 ( .A(G221), .ZN(n1339) );
NAND3_X1 U1061 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1333) );
XNOR2_X1 U1062 ( .A(KEYINPUT31), .B(KEYINPUT28), .ZN(n1343) );
NAND4_X1 U1063 ( .A1(n1344), .A2(n1321), .A3(n1345), .A4(n1346), .ZN(n1342) );
NAND2_X1 U1064 ( .A1(G146), .A2(n1347), .ZN(n1346) );
OR2_X1 U1065 ( .A1(n1322), .A2(n1347), .ZN(n1345) );
INV_X1 U1066 ( .A(n1348), .ZN(n1321) );
NAND2_X1 U1067 ( .A1(G125), .A2(n1349), .ZN(n1344) );
NAND3_X1 U1068 ( .A1(n1350), .A2(n1349), .A3(G125), .ZN(n1341) );
INV_X1 U1069 ( .A(KEYINPUT59), .ZN(n1349) );
NAND3_X1 U1070 ( .A1(n1351), .A2(n1352), .A3(n1322), .ZN(n1350) );
NAND2_X1 U1071 ( .A1(n1324), .A2(n1208), .ZN(n1322) );
NAND2_X1 U1072 ( .A1(n1208), .A2(n1347), .ZN(n1352) );
INV_X1 U1073 ( .A(KEYINPUT17), .ZN(n1347) );
NAND2_X1 U1074 ( .A1(n1348), .A2(KEYINPUT17), .ZN(n1351) );
NOR2_X1 U1075 ( .A1(n1324), .A2(n1208), .ZN(n1348) );
XOR2_X1 U1076 ( .A(G140), .B(KEYINPUT20), .Z(n1324) );
XNOR2_X1 U1077 ( .A(n1353), .B(G472), .ZN(n1086) );
NAND2_X1 U1078 ( .A1(n1151), .A2(n1141), .ZN(n1353) );
INV_X1 U1079 ( .A(G902), .ZN(n1141) );
XNOR2_X1 U1080 ( .A(n1354), .B(n1355), .ZN(n1151) );
XNOR2_X1 U1081 ( .A(n1356), .B(n1159), .ZN(n1355) );
XOR2_X1 U1082 ( .A(n1103), .B(KEYINPUT56), .Z(n1159) );
XOR2_X1 U1083 ( .A(G131), .B(n1357), .Z(n1103) );
XNOR2_X1 U1084 ( .A(n1218), .B(G134), .ZN(n1357) );
INV_X1 U1085 ( .A(G137), .ZN(n1218) );
NAND2_X1 U1086 ( .A1(n1358), .A2(n1359), .ZN(n1356) );
NAND2_X1 U1087 ( .A1(n1360), .A2(n1361), .ZN(n1359) );
XNOR2_X1 U1088 ( .A(KEYINPUT22), .B(n1246), .ZN(n1361) );
XNOR2_X1 U1089 ( .A(G119), .B(n1362), .ZN(n1360) );
XOR2_X1 U1090 ( .A(n1363), .B(KEYINPUT49), .Z(n1358) );
NAND2_X1 U1091 ( .A1(n1364), .A2(n1246), .ZN(n1363) );
INV_X1 U1092 ( .A(G113), .ZN(n1246) );
XOR2_X1 U1093 ( .A(G119), .B(n1362), .Z(n1364) );
NOR2_X1 U1094 ( .A1(G116), .A2(KEYINPUT3), .ZN(n1362) );
XOR2_X1 U1095 ( .A(n1365), .B(n1366), .Z(n1354) );
XNOR2_X1 U1096 ( .A(G101), .B(n1267), .ZN(n1366) );
NAND2_X1 U1097 ( .A1(n1367), .A2(n1288), .ZN(n1267) );
NAND2_X1 U1098 ( .A1(G146), .A2(n1291), .ZN(n1288) );
NAND2_X1 U1099 ( .A1(n1368), .A2(n1208), .ZN(n1367) );
INV_X1 U1100 ( .A(G146), .ZN(n1208) );
XNOR2_X1 U1101 ( .A(n1291), .B(KEYINPUT45), .ZN(n1368) );
XNOR2_X1 U1102 ( .A(G128), .B(n1304), .ZN(n1291) );
INV_X1 U1103 ( .A(G143), .ZN(n1304) );
NAND2_X1 U1104 ( .A1(G210), .A2(n1327), .ZN(n1365) );
NOR2_X1 U1105 ( .A1(G953), .A2(G237), .ZN(n1327) );
INV_X1 U1106 ( .A(G110), .ZN(n1255) );
endmodule


