//Key = 1011010001010011011011000100011011110101011011010010011001011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;

XOR2_X1 U734 ( .A(G107), .B(n1010), .Z(G9) );
NOR2_X1 U735 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U736 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR3_X1 U737 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NOR2_X1 U738 ( .A1(KEYINPUT18), .A2(n1018), .ZN(n1016) );
AND4_X1 U739 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NAND3_X1 U740 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1015) );
NAND2_X1 U741 ( .A1(n1022), .A2(n1026), .ZN(n1025) );
NAND2_X1 U742 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U743 ( .A1(n1019), .A2(n1029), .A3(n1030), .ZN(n1028) );
NAND2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NAND2_X1 U745 ( .A1(n1021), .A2(n1033), .ZN(n1032) );
NAND2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U747 ( .A1(KEYINPUT18), .A2(n1036), .ZN(n1035) );
INV_X1 U748 ( .A(n1037), .ZN(n1036) );
INV_X1 U749 ( .A(n1038), .ZN(n1034) );
NAND2_X1 U750 ( .A1(n1039), .A2(n1040), .ZN(n1031) );
NAND2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U753 ( .A1(n1039), .A2(n1045), .A3(n1021), .ZN(n1027) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1019), .A2(n1048), .ZN(n1047) );
NAND2_X1 U756 ( .A1(n1049), .A2(n1012), .ZN(n1048) );
NAND2_X1 U757 ( .A1(n1030), .A2(n1050), .ZN(n1046) );
NAND2_X1 U758 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U759 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
XNOR2_X1 U760 ( .A(n1055), .B(KEYINPUT36), .ZN(n1053) );
INV_X1 U761 ( .A(n1056), .ZN(n1022) );
NOR3_X1 U762 ( .A1(n1057), .A2(G953), .A3(G952), .ZN(n1013) );
INV_X1 U763 ( .A(n1023), .ZN(n1057) );
NAND4_X1 U764 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1023) );
NOR4_X1 U765 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061) );
XOR2_X1 U766 ( .A(KEYINPUT8), .B(n1066), .Z(n1065) );
NOR2_X1 U767 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XNOR2_X1 U768 ( .A(n1069), .B(KEYINPUT62), .ZN(n1063) );
XNOR2_X1 U769 ( .A(n1070), .B(n1071), .ZN(n1062) );
NAND2_X1 U770 ( .A1(KEYINPUT34), .A2(n1072), .ZN(n1070) );
NOR2_X1 U771 ( .A1(n1043), .A2(n1054), .ZN(n1060) );
NAND2_X1 U772 ( .A1(n1068), .A2(n1067), .ZN(n1059) );
XNOR2_X1 U773 ( .A(n1073), .B(KEYINPUT6), .ZN(n1068) );
XOR2_X1 U774 ( .A(n1074), .B(n1075), .Z(n1058) );
NOR2_X1 U775 ( .A1(n1076), .A2(KEYINPUT23), .ZN(n1074) );
XOR2_X1 U776 ( .A(n1077), .B(n1078), .Z(G72) );
NOR2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U778 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND3_X1 U779 ( .A1(n1083), .A2(n1084), .A3(KEYINPUT39), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U781 ( .A(KEYINPUT15), .B(n1087), .Z(n1085) );
NAND2_X1 U782 ( .A1(n1088), .A2(n1089), .ZN(n1083) );
XNOR2_X1 U783 ( .A(n1087), .B(KEYINPUT25), .ZN(n1089) );
XNOR2_X1 U784 ( .A(n1090), .B(n1091), .ZN(n1087) );
NAND3_X1 U785 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1077) );
INV_X1 U786 ( .A(n1079), .ZN(n1094) );
OR2_X1 U787 ( .A1(n1024), .A2(G227), .ZN(n1093) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1024), .ZN(n1092) );
NAND2_X1 U789 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U790 ( .A(n1098), .B(KEYINPUT43), .Z(n1096) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(G69) );
NOR2_X1 U792 ( .A1(n1101), .A2(G953), .ZN(n1100) );
XOR2_X1 U793 ( .A(n1102), .B(n1103), .Z(n1099) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND3_X1 U795 ( .A1(n1106), .A2(n1107), .A3(KEYINPUT11), .ZN(n1102) );
INV_X1 U796 ( .A(n1104), .ZN(n1107) );
OR2_X1 U797 ( .A1(n1024), .A2(G224), .ZN(n1106) );
NOR2_X1 U798 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XOR2_X1 U799 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND3_X1 U800 ( .A1(n1112), .A2(n1017), .A3(n1073), .ZN(n1110) );
INV_X1 U801 ( .A(n1113), .ZN(n1073) );
XNOR2_X1 U802 ( .A(KEYINPUT40), .B(n1114), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1108), .A2(n1115), .ZN(G63) );
XOR2_X1 U804 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U805 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NOR2_X1 U806 ( .A1(n1108), .A2(n1120), .ZN(G60) );
XOR2_X1 U807 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1119), .ZN(n1121) );
XOR2_X1 U809 ( .A(G104), .B(n1124), .Z(G6) );
NOR2_X1 U810 ( .A1(KEYINPUT22), .A2(n1125), .ZN(n1124) );
INV_X1 U811 ( .A(n1126), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1108), .A2(n1127), .ZN(G57) );
XOR2_X1 U813 ( .A(n1128), .B(n1129), .Z(n1127) );
XNOR2_X1 U814 ( .A(n1130), .B(n1131), .ZN(n1129) );
NAND2_X1 U815 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NAND2_X1 U816 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND2_X1 U817 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U818 ( .A1(KEYINPUT45), .A2(n1138), .ZN(n1137) );
INV_X1 U819 ( .A(KEYINPUT46), .ZN(n1136) );
NAND2_X1 U820 ( .A1(n1139), .A2(n1140), .ZN(n1132) );
NAND2_X1 U821 ( .A1(KEYINPUT45), .A2(n1141), .ZN(n1140) );
OR2_X1 U822 ( .A1(n1134), .A2(KEYINPUT46), .ZN(n1141) );
XOR2_X1 U823 ( .A(n1142), .B(n1143), .Z(n1134) );
NAND2_X1 U824 ( .A1(KEYINPUT60), .A2(n1144), .ZN(n1142) );
XOR2_X1 U825 ( .A(n1145), .B(n1146), .Z(n1128) );
NOR2_X1 U826 ( .A1(n1147), .A2(n1119), .ZN(n1146) );
NOR2_X1 U827 ( .A1(n1108), .A2(n1148), .ZN(G54) );
XOR2_X1 U828 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U829 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U830 ( .A(n1153), .B(n1086), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1154), .A2(n1119), .ZN(n1153) );
XOR2_X1 U832 ( .A(n1155), .B(n1156), .Z(n1149) );
XOR2_X1 U833 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U834 ( .A1(KEYINPUT33), .A2(n1159), .ZN(n1158) );
XNOR2_X1 U835 ( .A(n1144), .B(KEYINPUT49), .ZN(n1155) );
NOR2_X1 U836 ( .A1(n1108), .A2(n1160), .ZN(G51) );
XOR2_X1 U837 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U838 ( .A(n1163), .B(n1164), .ZN(n1162) );
XOR2_X1 U839 ( .A(n1165), .B(KEYINPUT48), .Z(n1164) );
XOR2_X1 U840 ( .A(n1105), .B(n1166), .Z(n1161) );
XOR2_X1 U841 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U842 ( .A1(KEYINPUT12), .A2(n1169), .ZN(n1168) );
NOR2_X1 U843 ( .A1(n1071), .A2(n1119), .ZN(n1167) );
NAND2_X1 U844 ( .A1(G902), .A2(n1017), .ZN(n1119) );
NAND3_X1 U845 ( .A1(n1097), .A2(n1098), .A3(n1101), .ZN(n1017) );
AND4_X1 U846 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1101) );
NOR4_X1 U847 ( .A1(n1174), .A2(n1126), .A3(n1175), .A4(n1176), .ZN(n1173) );
NOR4_X1 U848 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
XNOR2_X1 U849 ( .A(n1181), .B(KEYINPUT27), .ZN(n1178) );
NAND2_X1 U850 ( .A1(n1182), .A2(n1039), .ZN(n1177) );
NOR2_X1 U851 ( .A1(n1183), .A2(n1184), .ZN(n1175) );
XNOR2_X1 U852 ( .A(KEYINPUT57), .B(n1041), .ZN(n1184) );
NOR2_X1 U853 ( .A1(n1049), .A2(n1011), .ZN(n1126) );
NAND2_X1 U854 ( .A1(n1185), .A2(n1039), .ZN(n1011) );
AND2_X1 U855 ( .A1(n1186), .A2(n1187), .ZN(n1172) );
NAND2_X1 U856 ( .A1(n1188), .A2(n1021), .ZN(n1098) );
AND4_X1 U857 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1097) );
NOR4_X1 U858 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
INV_X1 U859 ( .A(n1197), .ZN(n1196) );
NAND2_X1 U860 ( .A1(n1198), .A2(n1199), .ZN(n1191) );
NOR2_X1 U861 ( .A1(n1024), .A2(G952), .ZN(n1108) );
XNOR2_X1 U862 ( .A(G146), .B(n1189), .ZN(G48) );
NAND3_X1 U863 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1189) );
XNOR2_X1 U864 ( .A(G143), .B(n1190), .ZN(G45) );
NAND2_X1 U865 ( .A1(n1203), .A2(n1204), .ZN(n1190) );
NAND2_X1 U866 ( .A1(n1205), .A2(n1206), .ZN(G42) );
NAND3_X1 U867 ( .A1(n1198), .A2(n1207), .A3(n1208), .ZN(n1206) );
XOR2_X1 U868 ( .A(n1209), .B(KEYINPUT1), .Z(n1205) );
NAND2_X1 U869 ( .A1(G140), .A2(n1210), .ZN(n1209) );
NAND2_X1 U870 ( .A1(n1208), .A2(n1198), .ZN(n1210) );
NOR4_X1 U871 ( .A1(n1211), .A2(n1049), .A3(n1037), .A4(n1051), .ZN(n1198) );
XOR2_X1 U872 ( .A(n1199), .B(KEYINPUT7), .Z(n1208) );
XNOR2_X1 U873 ( .A(G137), .B(n1212), .ZN(G39) );
NAND2_X1 U874 ( .A1(KEYINPUT37), .A2(n1195), .ZN(n1212) );
AND3_X1 U875 ( .A1(n1202), .A2(n1030), .A3(n1021), .ZN(n1195) );
XNOR2_X1 U876 ( .A(G134), .B(n1213), .ZN(G36) );
NAND2_X1 U877 ( .A1(n1214), .A2(n1021), .ZN(n1213) );
XNOR2_X1 U878 ( .A(n1188), .B(KEYINPUT54), .ZN(n1214) );
AND2_X1 U879 ( .A1(n1203), .A2(n1182), .ZN(n1188) );
XNOR2_X1 U880 ( .A(G131), .B(n1197), .ZN(G33) );
NAND3_X1 U881 ( .A1(n1021), .A2(n1200), .A3(n1203), .ZN(n1197) );
AND3_X1 U882 ( .A1(n1181), .A2(n1199), .A3(n1038), .ZN(n1203) );
INV_X1 U883 ( .A(n1211), .ZN(n1021) );
NAND2_X1 U884 ( .A1(n1044), .A2(n1215), .ZN(n1211) );
NAND2_X1 U885 ( .A1(n1216), .A2(n1217), .ZN(G30) );
NAND2_X1 U886 ( .A1(n1194), .A2(n1218), .ZN(n1217) );
XOR2_X1 U887 ( .A(KEYINPUT29), .B(n1219), .Z(n1216) );
NOR2_X1 U888 ( .A1(n1194), .A2(n1218), .ZN(n1219) );
AND3_X1 U889 ( .A1(n1182), .A2(n1201), .A3(n1202), .ZN(n1194) );
AND4_X1 U890 ( .A1(n1181), .A2(n1220), .A3(n1069), .A4(n1199), .ZN(n1202) );
XOR2_X1 U891 ( .A(G101), .B(n1174), .Z(G3) );
AND3_X1 U892 ( .A1(n1030), .A2(n1185), .A3(n1038), .ZN(n1174) );
XNOR2_X1 U893 ( .A(G125), .B(n1221), .ZN(G27) );
NAND2_X1 U894 ( .A1(KEYINPUT2), .A2(n1193), .ZN(n1221) );
AND4_X1 U895 ( .A1(n1019), .A2(n1199), .A3(n1201), .A4(n1222), .ZN(n1193) );
NOR2_X1 U896 ( .A1(n1037), .A2(n1049), .ZN(n1222) );
INV_X1 U897 ( .A(n1200), .ZN(n1049) );
NAND2_X1 U898 ( .A1(n1056), .A2(n1223), .ZN(n1199) );
NAND2_X1 U899 ( .A1(n1079), .A2(n1224), .ZN(n1223) );
NOR2_X1 U900 ( .A1(G900), .A2(n1024), .ZN(n1079) );
XNOR2_X1 U901 ( .A(G122), .B(n1170), .ZN(G24) );
NAND3_X1 U902 ( .A1(n1225), .A2(n1039), .A3(n1204), .ZN(n1170) );
AND3_X1 U903 ( .A1(n1226), .A2(n1227), .A3(n1201), .ZN(n1204) );
NOR2_X1 U904 ( .A1(n1069), .A2(n1220), .ZN(n1039) );
XOR2_X1 U905 ( .A(G119), .B(n1228), .Z(G21) );
NOR2_X1 U906 ( .A1(n1041), .A2(n1183), .ZN(n1228) );
NAND4_X1 U907 ( .A1(n1225), .A2(n1030), .A3(n1220), .A4(n1069), .ZN(n1183) );
INV_X1 U908 ( .A(n1201), .ZN(n1041) );
XNOR2_X1 U909 ( .A(G116), .B(n1171), .ZN(G18) );
NAND4_X1 U910 ( .A1(n1225), .A2(n1038), .A3(n1182), .A4(n1201), .ZN(n1171) );
INV_X1 U911 ( .A(n1012), .ZN(n1182) );
NAND2_X1 U912 ( .A1(n1229), .A2(n1227), .ZN(n1012) );
XNOR2_X1 U913 ( .A(n1226), .B(KEYINPUT56), .ZN(n1229) );
XNOR2_X1 U914 ( .A(G113), .B(n1187), .ZN(G15) );
NAND4_X1 U915 ( .A1(n1200), .A2(n1225), .A3(n1038), .A4(n1230), .ZN(n1187) );
NOR2_X1 U916 ( .A1(n1220), .A2(n1231), .ZN(n1038) );
AND2_X1 U917 ( .A1(n1019), .A2(n1232), .ZN(n1225) );
NAND2_X1 U918 ( .A1(n1233), .A2(n1234), .ZN(n1019) );
OR3_X1 U919 ( .A1(n1055), .A2(n1054), .A3(KEYINPUT36), .ZN(n1234) );
NAND2_X1 U920 ( .A1(KEYINPUT36), .A2(n1181), .ZN(n1233) );
NOR2_X1 U921 ( .A1(n1227), .A2(n1235), .ZN(n1200) );
INV_X1 U922 ( .A(n1226), .ZN(n1235) );
XNOR2_X1 U923 ( .A(G110), .B(n1186), .ZN(G12) );
NAND2_X1 U924 ( .A1(n1020), .A2(n1185), .ZN(n1186) );
NOR3_X1 U925 ( .A1(n1180), .A2(n1179), .A3(n1051), .ZN(n1185) );
INV_X1 U926 ( .A(n1181), .ZN(n1051) );
NOR2_X1 U927 ( .A1(n1236), .A2(n1054), .ZN(n1181) );
AND2_X1 U928 ( .A1(G221), .A2(n1237), .ZN(n1054) );
INV_X1 U929 ( .A(n1055), .ZN(n1236) );
XOR2_X1 U930 ( .A(n1076), .B(n1075), .Z(n1055) );
XNOR2_X1 U931 ( .A(n1154), .B(KEYINPUT52), .ZN(n1075) );
INV_X1 U932 ( .A(G469), .ZN(n1154) );
AND2_X1 U933 ( .A1(n1238), .A2(n1114), .ZN(n1076) );
XOR2_X1 U934 ( .A(n1239), .B(n1240), .Z(n1238) );
XNOR2_X1 U935 ( .A(n1241), .B(n1157), .ZN(n1240) );
NAND2_X1 U936 ( .A1(G227), .A2(n1024), .ZN(n1157) );
NOR2_X1 U937 ( .A1(KEYINPUT63), .A2(n1242), .ZN(n1241) );
XOR2_X1 U938 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U939 ( .A(n1086), .B(n1159), .ZN(n1244) );
XOR2_X1 U940 ( .A(n1245), .B(G104), .Z(n1159) );
INV_X1 U941 ( .A(n1088), .ZN(n1086) );
XOR2_X1 U942 ( .A(G143), .B(n1246), .Z(n1088) );
XNOR2_X1 U943 ( .A(n1144), .B(KEYINPUT3), .ZN(n1243) );
NOR2_X1 U944 ( .A1(KEYINPUT31), .A2(n1151), .ZN(n1239) );
XNOR2_X1 U945 ( .A(G110), .B(G140), .ZN(n1151) );
INV_X1 U946 ( .A(n1232), .ZN(n1179) );
NAND2_X1 U947 ( .A1(n1056), .A2(n1247), .ZN(n1232) );
NAND2_X1 U948 ( .A1(n1224), .A2(n1104), .ZN(n1247) );
NOR2_X1 U949 ( .A1(G898), .A2(n1024), .ZN(n1104) );
AND2_X1 U950 ( .A1(n1248), .A2(n1249), .ZN(n1224) );
XNOR2_X1 U951 ( .A(G902), .B(KEYINPUT0), .ZN(n1248) );
NAND3_X1 U952 ( .A1(n1249), .A2(n1024), .A3(G952), .ZN(n1056) );
NAND2_X1 U953 ( .A1(G237), .A2(G234), .ZN(n1249) );
INV_X1 U954 ( .A(n1230), .ZN(n1180) );
XOR2_X1 U955 ( .A(n1201), .B(KEYINPUT13), .Z(n1230) );
NOR2_X1 U956 ( .A1(n1044), .A2(n1043), .ZN(n1201) );
INV_X1 U957 ( .A(n1215), .ZN(n1043) );
NAND2_X1 U958 ( .A1(G214), .A2(n1250), .ZN(n1215) );
XOR2_X1 U959 ( .A(n1251), .B(n1071), .Z(n1044) );
NAND2_X1 U960 ( .A1(G210), .A2(n1250), .ZN(n1071) );
NAND2_X1 U961 ( .A1(n1252), .A2(n1114), .ZN(n1250) );
INV_X1 U962 ( .A(G237), .ZN(n1252) );
NAND2_X1 U963 ( .A1(KEYINPUT20), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U964 ( .A(KEYINPUT41), .B(n1072), .ZN(n1253) );
NAND2_X1 U965 ( .A1(n1254), .A2(n1114), .ZN(n1072) );
XOR2_X1 U966 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U967 ( .A(n1165), .B(n1257), .Z(n1256) );
NOR2_X1 U968 ( .A1(KEYINPUT55), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U969 ( .A(n1163), .B(n1169), .ZN(n1258) );
INV_X1 U970 ( .A(n1143), .ZN(n1163) );
NAND2_X1 U971 ( .A1(G224), .A2(n1024), .ZN(n1165) );
NAND2_X1 U972 ( .A1(KEYINPUT42), .A2(n1105), .ZN(n1255) );
XOR2_X1 U973 ( .A(n1259), .B(n1260), .Z(n1105) );
XOR2_X1 U974 ( .A(n1245), .B(n1261), .Z(n1260) );
XNOR2_X1 U975 ( .A(G107), .B(n1262), .ZN(n1245) );
XNOR2_X1 U976 ( .A(n1263), .B(n1264), .ZN(n1259) );
NAND3_X1 U977 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1263) );
OR2_X1 U978 ( .A1(n1268), .A2(KEYINPUT14), .ZN(n1267) );
NAND3_X1 U979 ( .A1(KEYINPUT14), .A2(n1268), .A3(n1269), .ZN(n1266) );
NAND2_X1 U980 ( .A1(n1270), .A2(n1271), .ZN(n1265) );
NAND2_X1 U981 ( .A1(n1272), .A2(KEYINPUT14), .ZN(n1271) );
XNOR2_X1 U982 ( .A(n1268), .B(KEYINPUT17), .ZN(n1272) );
XNOR2_X1 U983 ( .A(n1273), .B(KEYINPUT4), .ZN(n1268) );
INV_X1 U984 ( .A(n1269), .ZN(n1270) );
XOR2_X1 U985 ( .A(G113), .B(KEYINPUT24), .Z(n1269) );
NOR2_X1 U986 ( .A1(n1037), .A2(n1064), .ZN(n1020) );
INV_X1 U987 ( .A(n1030), .ZN(n1064) );
NOR2_X1 U988 ( .A1(n1227), .A2(n1226), .ZN(n1030) );
XOR2_X1 U989 ( .A(n1274), .B(n1123), .Z(n1226) );
INV_X1 U990 ( .A(G475), .ZN(n1123) );
OR2_X1 U991 ( .A1(n1122), .A2(G902), .ZN(n1274) );
XOR2_X1 U992 ( .A(n1261), .B(n1275), .Z(n1122) );
XNOR2_X1 U993 ( .A(n1276), .B(n1277), .ZN(n1275) );
NOR4_X1 U994 ( .A1(n1278), .A2(n1279), .A3(KEYINPUT61), .A4(n1280), .ZN(n1277) );
AND2_X1 U995 ( .A1(n1281), .A2(KEYINPUT10), .ZN(n1280) );
NOR2_X1 U996 ( .A1(n1282), .A2(n1283), .ZN(n1279) );
INV_X1 U997 ( .A(n1284), .ZN(n1283) );
NOR2_X1 U998 ( .A1(n1281), .A2(n1285), .ZN(n1282) );
NOR4_X1 U999 ( .A1(n1284), .A2(n1285), .A3(KEYINPUT10), .A4(n1281), .ZN(n1278) );
XOR2_X1 U1000 ( .A(n1286), .B(n1287), .Z(n1281) );
XNOR2_X1 U1001 ( .A(n1288), .B(G131), .ZN(n1287) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1289), .ZN(n1286) );
INV_X1 U1003 ( .A(KEYINPUT59), .ZN(n1285) );
XOR2_X1 U1004 ( .A(G146), .B(n1082), .Z(n1284) );
XNOR2_X1 U1005 ( .A(n1207), .B(n1169), .ZN(n1082) );
XOR2_X1 U1006 ( .A(G104), .B(G122), .Z(n1261) );
XOR2_X1 U1007 ( .A(n1290), .B(n1118), .Z(n1227) );
INV_X1 U1008 ( .A(G478), .ZN(n1118) );
OR2_X1 U1009 ( .A1(n1117), .A2(G902), .ZN(n1290) );
XNOR2_X1 U1010 ( .A(n1291), .B(n1292), .ZN(n1117) );
XNOR2_X1 U1011 ( .A(n1293), .B(n1294), .ZN(n1292) );
XOR2_X1 U1012 ( .A(KEYINPUT28), .B(G122), .Z(n1294) );
INV_X1 U1013 ( .A(G116), .ZN(n1293) );
XOR2_X1 U1014 ( .A(n1295), .B(n1296), .Z(n1291) );
NOR2_X1 U1015 ( .A1(KEYINPUT19), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U1016 ( .A(n1218), .B(n1298), .ZN(n1297) );
XNOR2_X1 U1017 ( .A(n1288), .B(G134), .ZN(n1298) );
XOR2_X1 U1018 ( .A(n1299), .B(G107), .Z(n1295) );
NAND3_X1 U1019 ( .A1(n1300), .A2(n1024), .A3(G217), .ZN(n1299) );
NAND2_X1 U1020 ( .A1(n1231), .A2(n1220), .ZN(n1037) );
XNOR2_X1 U1021 ( .A(n1067), .B(n1113), .ZN(n1220) );
NAND2_X1 U1022 ( .A1(G217), .A2(n1237), .ZN(n1113) );
NAND2_X1 U1023 ( .A1(G234), .A2(n1114), .ZN(n1237) );
AND2_X1 U1024 ( .A1(n1111), .A2(n1114), .ZN(n1067) );
XNOR2_X1 U1025 ( .A(n1301), .B(n1302), .ZN(n1111) );
XOR2_X1 U1026 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U1027 ( .A(n1305), .B(n1246), .ZN(n1304) );
XNOR2_X1 U1028 ( .A(G146), .B(n1218), .ZN(n1246) );
NAND3_X1 U1029 ( .A1(n1300), .A2(n1024), .A3(G221), .ZN(n1305) );
INV_X1 U1030 ( .A(G953), .ZN(n1024) );
XNOR2_X1 U1031 ( .A(G234), .B(KEYINPUT21), .ZN(n1300) );
XOR2_X1 U1032 ( .A(n1306), .B(n1307), .Z(n1301) );
XNOR2_X1 U1033 ( .A(G119), .B(n1264), .ZN(n1307) );
INV_X1 U1034 ( .A(G110), .ZN(n1264) );
NAND3_X1 U1035 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1306) );
OR2_X1 U1036 ( .A1(n1207), .A2(n1169), .ZN(n1310) );
NAND2_X1 U1037 ( .A1(KEYINPUT16), .A2(n1311), .ZN(n1309) );
NAND2_X1 U1038 ( .A1(n1312), .A2(n1207), .ZN(n1311) );
XNOR2_X1 U1039 ( .A(KEYINPUT35), .B(n1169), .ZN(n1312) );
NAND2_X1 U1040 ( .A1(n1313), .A2(n1314), .ZN(n1308) );
INV_X1 U1041 ( .A(KEYINPUT16), .ZN(n1314) );
NAND2_X1 U1042 ( .A1(n1315), .A2(n1316), .ZN(n1313) );
OR2_X1 U1043 ( .A1(n1169), .A2(KEYINPUT35), .ZN(n1316) );
NAND3_X1 U1044 ( .A1(n1169), .A2(n1207), .A3(KEYINPUT35), .ZN(n1315) );
INV_X1 U1045 ( .A(G140), .ZN(n1207) );
XOR2_X1 U1046 ( .A(G125), .B(KEYINPUT26), .Z(n1169) );
INV_X1 U1047 ( .A(n1069), .ZN(n1231) );
XOR2_X1 U1048 ( .A(n1317), .B(n1147), .Z(n1069) );
INV_X1 U1049 ( .A(G472), .ZN(n1147) );
NAND2_X1 U1050 ( .A1(n1318), .A2(n1114), .ZN(n1317) );
INV_X1 U1051 ( .A(G902), .ZN(n1114) );
XOR2_X1 U1052 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1053 ( .A(n1139), .B(n1145), .ZN(n1320) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1289), .ZN(n1145) );
NOR2_X1 U1055 ( .A1(G953), .A2(G237), .ZN(n1289) );
INV_X1 U1056 ( .A(n1138), .ZN(n1139) );
XOR2_X1 U1057 ( .A(n1321), .B(n1276), .Z(n1138) );
INV_X1 U1058 ( .A(G113), .ZN(n1276) );
NAND2_X1 U1059 ( .A1(KEYINPUT44), .A2(n1273), .ZN(n1321) );
XNOR2_X1 U1060 ( .A(G116), .B(G119), .ZN(n1273) );
XNOR2_X1 U1061 ( .A(n1322), .B(n1143), .ZN(n1319) );
NAND2_X1 U1062 ( .A1(n1323), .A2(n1324), .ZN(n1143) );
NAND2_X1 U1063 ( .A1(n1325), .A2(n1218), .ZN(n1324) );
XOR2_X1 U1064 ( .A(KEYINPUT30), .B(n1326), .Z(n1325) );
XOR2_X1 U1065 ( .A(KEYINPUT50), .B(n1327), .Z(n1323) );
NOR2_X1 U1066 ( .A1(n1328), .A2(n1218), .ZN(n1327) );
INV_X1 U1067 ( .A(G128), .ZN(n1218) );
XNOR2_X1 U1068 ( .A(n1326), .B(KEYINPUT38), .ZN(n1328) );
XNOR2_X1 U1069 ( .A(n1288), .B(G146), .ZN(n1326) );
INV_X1 U1070 ( .A(G143), .ZN(n1288) );
XNOR2_X1 U1071 ( .A(n1144), .B(n1329), .ZN(n1322) );
NOR2_X1 U1072 ( .A1(n1262), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1073 ( .A(KEYINPUT9), .B(KEYINPUT58), .ZN(n1330) );
INV_X1 U1074 ( .A(n1131), .ZN(n1262) );
XOR2_X1 U1075 ( .A(G101), .B(KEYINPUT47), .Z(n1131) );
AND2_X1 U1076 ( .A1(n1331), .A2(n1332), .ZN(n1144) );
NAND2_X1 U1077 ( .A1(n1333), .A2(G131), .ZN(n1332) );
XOR2_X1 U1078 ( .A(n1334), .B(KEYINPUT51), .Z(n1331) );
NAND2_X1 U1079 ( .A1(n1335), .A2(n1091), .ZN(n1334) );
INV_X1 U1080 ( .A(G131), .ZN(n1091) );
XOR2_X1 U1081 ( .A(KEYINPUT32), .B(n1333), .Z(n1335) );
AND2_X1 U1082 ( .A1(n1336), .A2(n1337), .ZN(n1333) );
NAND3_X1 U1083 ( .A1(G134), .A2(n1303), .A3(n1338), .ZN(n1337) );
INV_X1 U1084 ( .A(KEYINPUT5), .ZN(n1338) );
NAND2_X1 U1085 ( .A1(n1090), .A2(KEYINPUT5), .ZN(n1336) );
XOR2_X1 U1086 ( .A(G134), .B(n1303), .Z(n1090) );
XOR2_X1 U1087 ( .A(G137), .B(KEYINPUT53), .Z(n1303) );
endmodule


