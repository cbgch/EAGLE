//Key = 0010010110000011100110011000000000100101110111101111110011011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353;

NAND2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(G9) );
NAND2_X1 U746 ( .A1(G107), .A2(n1034), .ZN(n1033) );
XOR2_X1 U747 ( .A(n1035), .B(KEYINPUT30), .Z(n1032) );
OR2_X1 U748 ( .A1(n1034), .A2(G107), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1036), .A2(n1037), .ZN(G75) );
AND4_X1 U750 ( .A1(n1038), .A2(n1039), .A3(KEYINPUT41), .A4(n1040), .ZN(n1037) );
NOR4_X1 U751 ( .A1(G953), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1040) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1044) );
NOR4_X1 U754 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1049) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U757 ( .A1(n1057), .A2(n1058), .ZN(n1047) );
NOR2_X1 U758 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
AND2_X1 U759 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U760 ( .A1(n1063), .A2(n1051), .ZN(n1059) );
NOR2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
AND2_X1 U762 ( .A1(n1066), .A2(KEYINPUT19), .ZN(n1064) );
NOR2_X1 U763 ( .A1(n1067), .A2(KEYINPUT19), .ZN(n1046) );
NOR3_X1 U764 ( .A1(n1058), .A2(n1068), .A3(n1051), .ZN(n1067) );
NOR3_X1 U765 ( .A1(n1058), .A2(n1069), .A3(n1050), .ZN(n1042) );
INV_X1 U766 ( .A(n1061), .ZN(n1050) );
NOR2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U768 ( .A1(n1072), .A2(n1051), .ZN(n1071) );
NOR2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR2_X1 U770 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
AND3_X1 U771 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1070) );
NAND2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1058) );
INV_X1 U773 ( .A(n1082), .ZN(n1039) );
NOR3_X1 U774 ( .A1(n1041), .A2(G953), .A3(G952), .ZN(n1036) );
AND4_X1 U775 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1041) );
NOR4_X1 U776 ( .A1(n1087), .A2(n1088), .A3(n1045), .A4(n1089), .ZN(n1086) );
XOR2_X1 U777 ( .A(G469), .B(n1090), .Z(n1089) );
NOR3_X1 U778 ( .A1(n1077), .A2(n1091), .A3(n1092), .ZN(n1085) );
NAND2_X1 U779 ( .A1(G472), .A2(n1093), .ZN(n1084) );
NAND2_X1 U780 ( .A1(n1094), .A2(G478), .ZN(n1083) );
XOR2_X1 U781 ( .A(n1095), .B(KEYINPUT13), .Z(n1094) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(G72) );
NOR2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U784 ( .A1(KEYINPUT45), .A2(n1100), .ZN(n1099) );
INV_X1 U785 ( .A(n1101), .ZN(n1100) );
NOR2_X1 U786 ( .A1(KEYINPUT9), .A2(n1101), .ZN(n1098) );
NAND3_X1 U787 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NAND2_X1 U788 ( .A1(G953), .A2(n1105), .ZN(n1104) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(n1106) );
OR2_X1 U792 ( .A1(n1112), .A2(KEYINPUT12), .ZN(n1110) );
NAND3_X1 U793 ( .A1(n1113), .A2(n1109), .A3(n1108), .ZN(n1102) );
INV_X1 U794 ( .A(KEYINPUT25), .ZN(n1109) );
XOR2_X1 U795 ( .A(n1114), .B(n1111), .Z(n1113) );
XNOR2_X1 U796 ( .A(n1115), .B(KEYINPUT5), .ZN(n1111) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1116), .ZN(n1114) );
INV_X1 U798 ( .A(KEYINPUT12), .ZN(n1116) );
XOR2_X1 U799 ( .A(n1117), .B(n1118), .Z(n1096) );
NOR2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1105), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(n1117) );
NAND4_X1 U803 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1123) );
XNOR2_X1 U804 ( .A(G953), .B(KEYINPUT11), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1128), .A2(n1129), .ZN(G69) );
NAND2_X1 U806 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
OR2_X1 U807 ( .A1(n1120), .A2(G224), .ZN(n1131) );
NAND3_X1 U808 ( .A1(n1132), .A2(n1133), .A3(G953), .ZN(n1128) );
NAND2_X1 U809 ( .A1(G898), .A2(G224), .ZN(n1133) );
XOR2_X1 U810 ( .A(KEYINPUT39), .B(n1130), .Z(n1132) );
XNOR2_X1 U811 ( .A(n1134), .B(n1135), .ZN(n1130) );
NOR2_X1 U812 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U813 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U814 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U815 ( .A(KEYINPUT42), .B(n1142), .ZN(n1138) );
NOR2_X1 U816 ( .A1(KEYINPUT6), .A2(n1143), .ZN(n1142) );
XNOR2_X1 U817 ( .A(G101), .B(n1144), .ZN(n1143) );
NOR2_X1 U818 ( .A1(G898), .A2(n1120), .ZN(n1136) );
NAND2_X1 U819 ( .A1(n1120), .A2(n1082), .ZN(n1134) );
NOR2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XNOR2_X1 U821 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U822 ( .A(n1149), .B(KEYINPUT26), .Z(n1147) );
NAND2_X1 U823 ( .A1(n1150), .A2(G217), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1145), .A2(n1151), .ZN(G63) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U826 ( .A1(n1150), .A2(G478), .ZN(n1152) );
NOR2_X1 U827 ( .A1(n1145), .A2(n1154), .ZN(G60) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U829 ( .A1(n1157), .A2(KEYINPUT62), .ZN(n1155) );
AND2_X1 U830 ( .A1(G475), .A2(n1150), .ZN(n1157) );
XNOR2_X1 U831 ( .A(G104), .B(n1158), .ZN(G6) );
NOR2_X1 U832 ( .A1(n1145), .A2(n1159), .ZN(G57) );
XOR2_X1 U833 ( .A(n1160), .B(n1161), .Z(n1159) );
XNOR2_X1 U834 ( .A(n1162), .B(n1163), .ZN(n1161) );
XNOR2_X1 U835 ( .A(n1164), .B(n1165), .ZN(n1160) );
NAND2_X1 U836 ( .A1(n1150), .A2(G472), .ZN(n1164) );
NOR2_X1 U837 ( .A1(n1145), .A2(n1166), .ZN(G54) );
XOR2_X1 U838 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U839 ( .A(n1169), .B(n1170), .ZN(n1168) );
XOR2_X1 U840 ( .A(n1171), .B(n1108), .Z(n1170) );
XOR2_X1 U841 ( .A(n1172), .B(n1173), .Z(n1167) );
XOR2_X1 U842 ( .A(KEYINPUT4), .B(G140), .Z(n1173) );
XNOR2_X1 U843 ( .A(n1174), .B(n1175), .ZN(n1172) );
NAND2_X1 U844 ( .A1(KEYINPUT15), .A2(n1176), .ZN(n1175) );
NAND3_X1 U845 ( .A1(n1150), .A2(G469), .A3(KEYINPUT60), .ZN(n1174) );
NOR2_X1 U846 ( .A1(n1145), .A2(n1177), .ZN(G51) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U848 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U849 ( .A1(KEYINPUT49), .A2(n1182), .ZN(n1181) );
NAND2_X1 U850 ( .A1(n1150), .A2(G210), .ZN(n1180) );
AND2_X1 U851 ( .A1(G902), .A2(n1183), .ZN(n1150) );
NAND2_X1 U852 ( .A1(n1038), .A2(n1184), .ZN(n1183) );
XNOR2_X1 U853 ( .A(KEYINPUT31), .B(n1082), .ZN(n1184) );
NAND4_X1 U854 ( .A1(n1158), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1082) );
AND4_X1 U855 ( .A1(n1034), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1187) );
NAND3_X1 U856 ( .A1(n1065), .A2(n1191), .A3(n1081), .ZN(n1034) );
NAND2_X1 U857 ( .A1(n1074), .A2(n1192), .ZN(n1186) );
NAND2_X1 U858 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XOR2_X1 U859 ( .A(n1195), .B(KEYINPUT35), .Z(n1193) );
NAND3_X1 U860 ( .A1(n1081), .A2(n1191), .A3(n1066), .ZN(n1158) );
AND4_X1 U861 ( .A1(n1124), .A2(n1196), .A3(n1125), .A4(n1126), .ZN(n1038) );
NAND2_X1 U862 ( .A1(n1197), .A2(n1198), .ZN(n1126) );
XNOR2_X1 U863 ( .A(n1199), .B(KEYINPUT14), .ZN(n1197) );
NAND3_X1 U864 ( .A1(n1199), .A2(n1061), .A3(n1200), .ZN(n1125) );
XNOR2_X1 U865 ( .A(KEYINPUT34), .B(n1127), .ZN(n1196) );
AND4_X1 U866 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1124) );
NOR2_X1 U867 ( .A1(n1205), .A2(n1206), .ZN(n1203) );
INV_X1 U868 ( .A(n1207), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1120), .A2(G952), .ZN(n1145) );
XNOR2_X1 U870 ( .A(G146), .B(n1208), .ZN(G48) );
NAND2_X1 U871 ( .A1(n1198), .A2(n1199), .ZN(n1208) );
AND2_X1 U872 ( .A1(n1066), .A2(n1209), .ZN(n1198) );
XNOR2_X1 U873 ( .A(G143), .B(n1201), .ZN(G45) );
NAND4_X1 U874 ( .A1(n1209), .A2(n1054), .A3(n1088), .A4(n1210), .ZN(n1201) );
XNOR2_X1 U875 ( .A(n1202), .B(n1211), .ZN(G42) );
XOR2_X1 U876 ( .A(KEYINPUT3), .B(G140), .Z(n1211) );
NAND2_X1 U877 ( .A1(n1212), .A2(n1200), .ZN(n1202) );
XNOR2_X1 U878 ( .A(G137), .B(n1213), .ZN(G39) );
NAND4_X1 U879 ( .A1(n1214), .A2(KEYINPUT57), .A3(n1200), .A4(n1061), .ZN(n1213) );
XNOR2_X1 U880 ( .A(n1199), .B(KEYINPUT7), .ZN(n1214) );
XNOR2_X1 U881 ( .A(G134), .B(n1204), .ZN(G36) );
NAND3_X1 U882 ( .A1(n1065), .A2(n1054), .A3(n1200), .ZN(n1204) );
XOR2_X1 U883 ( .A(n1206), .B(n1215), .Z(G33) );
NOR2_X1 U884 ( .A1(KEYINPUT29), .A2(n1216), .ZN(n1215) );
INV_X1 U885 ( .A(G131), .ZN(n1216) );
AND3_X1 U886 ( .A1(n1066), .A2(n1054), .A3(n1200), .ZN(n1206) );
AND3_X1 U887 ( .A1(n1062), .A2(n1217), .A3(n1079), .ZN(n1200) );
INV_X1 U888 ( .A(n1045), .ZN(n1079) );
NAND2_X1 U889 ( .A1(n1218), .A2(n1076), .ZN(n1045) );
INV_X1 U890 ( .A(n1075), .ZN(n1218) );
XNOR2_X1 U891 ( .A(G128), .B(n1207), .ZN(G30) );
NAND3_X1 U892 ( .A1(n1209), .A2(n1065), .A3(n1199), .ZN(n1207) );
AND3_X1 U893 ( .A1(n1074), .A2(n1217), .A3(n1062), .ZN(n1209) );
XNOR2_X1 U894 ( .A(G101), .B(n1185), .ZN(G3) );
NAND3_X1 U895 ( .A1(n1054), .A2(n1061), .A3(n1191), .ZN(n1185) );
AND2_X1 U896 ( .A1(n1062), .A2(n1219), .ZN(n1191) );
NAND3_X1 U897 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(G27) );
NAND2_X1 U898 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NAND2_X1 U899 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
INV_X1 U900 ( .A(KEYINPUT2), .ZN(n1226) );
NAND2_X1 U901 ( .A1(n1227), .A2(n1127), .ZN(n1225) );
XNOR2_X1 U902 ( .A(KEYINPUT33), .B(n1224), .ZN(n1227) );
NAND2_X1 U903 ( .A1(KEYINPUT2), .A2(n1228), .ZN(n1220) );
NAND2_X1 U904 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
OR3_X1 U905 ( .A1(n1224), .A2(n1223), .A3(KEYINPUT33), .ZN(n1230) );
INV_X1 U906 ( .A(n1127), .ZN(n1223) );
NAND4_X1 U907 ( .A1(n1231), .A2(n1212), .A3(n1074), .A4(n1217), .ZN(n1127) );
NAND2_X1 U908 ( .A1(n1052), .A2(n1232), .ZN(n1217) );
NAND4_X1 U909 ( .A1(G902), .A2(G953), .A3(n1233), .A4(n1105), .ZN(n1232) );
INV_X1 U910 ( .A(G900), .ZN(n1105) );
XNOR2_X1 U911 ( .A(KEYINPUT52), .B(n1234), .ZN(n1233) );
NOR3_X1 U912 ( .A1(n1056), .A2(n1055), .A3(n1068), .ZN(n1212) );
NAND2_X1 U913 ( .A1(KEYINPUT33), .A2(n1224), .ZN(n1229) );
XNOR2_X1 U914 ( .A(G122), .B(n1190), .ZN(G24) );
NAND4_X1 U915 ( .A1(n1235), .A2(n1081), .A3(n1088), .A4(n1210), .ZN(n1190) );
XNOR2_X1 U916 ( .A(G119), .B(n1189), .ZN(G21) );
NAND3_X1 U917 ( .A1(n1199), .A2(n1061), .A3(n1235), .ZN(n1189) );
NOR2_X1 U918 ( .A1(n1055), .A2(n1236), .ZN(n1199) );
NAND2_X1 U919 ( .A1(n1237), .A2(n1238), .ZN(G18) );
NAND2_X1 U920 ( .A1(KEYINPUT54), .A2(n1239), .ZN(n1238) );
XOR2_X1 U921 ( .A(n1240), .B(n1241), .Z(n1237) );
NOR2_X1 U922 ( .A1(n1242), .A2(n1195), .ZN(n1241) );
NAND4_X1 U923 ( .A1(n1231), .A2(n1065), .A3(n1054), .A4(n1243), .ZN(n1195) );
OR2_X1 U924 ( .A1(n1239), .A2(KEYINPUT54), .ZN(n1240) );
XNOR2_X1 U925 ( .A(G113), .B(n1188), .ZN(G15) );
NAND3_X1 U926 ( .A1(n1066), .A2(n1054), .A3(n1235), .ZN(n1188) );
AND2_X1 U927 ( .A1(n1231), .A2(n1219), .ZN(n1235) );
AND2_X1 U928 ( .A1(n1074), .A2(n1243), .ZN(n1219) );
NAND2_X1 U929 ( .A1(n1244), .A2(n1052), .ZN(n1243) );
INV_X1 U930 ( .A(n1245), .ZN(n1244) );
INV_X1 U931 ( .A(n1242), .ZN(n1074) );
INV_X1 U932 ( .A(n1051), .ZN(n1231) );
NAND2_X1 U933 ( .A1(n1078), .A2(n1246), .ZN(n1051) );
NAND2_X1 U934 ( .A1(n1247), .A2(n1248), .ZN(n1054) );
NAND2_X1 U935 ( .A1(n1081), .A2(n1249), .ZN(n1248) );
INV_X1 U936 ( .A(KEYINPUT56), .ZN(n1249) );
NOR2_X1 U937 ( .A1(n1056), .A2(n1087), .ZN(n1081) );
NAND3_X1 U938 ( .A1(n1055), .A2(n1056), .A3(KEYINPUT56), .ZN(n1247) );
INV_X1 U939 ( .A(n1236), .ZN(n1056) );
INV_X1 U940 ( .A(n1068), .ZN(n1066) );
NAND2_X1 U941 ( .A1(n1250), .A2(n1088), .ZN(n1068) );
XNOR2_X1 U942 ( .A(n1251), .B(KEYINPUT44), .ZN(n1250) );
XNOR2_X1 U943 ( .A(n1176), .B(n1252), .ZN(G12) );
NOR2_X1 U944 ( .A1(n1253), .A2(n1242), .ZN(n1252) );
NAND2_X1 U945 ( .A1(n1075), .A2(n1076), .ZN(n1242) );
NAND2_X1 U946 ( .A1(G214), .A2(n1254), .ZN(n1076) );
XNOR2_X1 U947 ( .A(n1255), .B(n1256), .ZN(n1075) );
AND2_X1 U948 ( .A1(n1254), .A2(G210), .ZN(n1256) );
OR2_X1 U949 ( .A1(G902), .A2(G237), .ZN(n1254) );
NAND2_X1 U950 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
XOR2_X1 U951 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U952 ( .A(n1178), .B(n1182), .Z(n1260) );
XNOR2_X1 U953 ( .A(n1261), .B(n1262), .ZN(n1178) );
XOR2_X1 U954 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U955 ( .A(n1224), .B(n1144), .ZN(n1264) );
NOR2_X1 U956 ( .A1(KEYINPUT28), .A2(n1265), .ZN(n1144) );
XOR2_X1 U957 ( .A(KEYINPUT37), .B(KEYINPUT32), .Z(n1263) );
XOR2_X1 U958 ( .A(n1162), .B(n1266), .Z(n1261) );
XOR2_X1 U959 ( .A(n1267), .B(n1140), .Z(n1266) );
NAND2_X1 U960 ( .A1(n1268), .A2(n1269), .ZN(n1140) );
NAND2_X1 U961 ( .A1(G110), .A2(n1270), .ZN(n1269) );
XOR2_X1 U962 ( .A(n1271), .B(KEYINPUT1), .Z(n1268) );
NAND2_X1 U963 ( .A1(G122), .A2(n1176), .ZN(n1271) );
NAND2_X1 U964 ( .A1(G224), .A2(n1272), .ZN(n1267) );
XNOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT40), .ZN(n1259) );
XNOR2_X1 U966 ( .A(KEYINPUT24), .B(n1273), .ZN(n1257) );
XOR2_X1 U967 ( .A(n1194), .B(KEYINPUT0), .Z(n1253) );
NAND4_X1 U968 ( .A1(n1062), .A2(n1236), .A3(n1274), .A4(n1061), .ZN(n1194) );
NAND2_X1 U969 ( .A1(n1275), .A2(n1276), .ZN(n1061) );
NAND2_X1 U970 ( .A1(n1065), .A2(n1277), .ZN(n1276) );
NOR2_X1 U971 ( .A1(n1088), .A2(n1251), .ZN(n1065) );
OR3_X1 U972 ( .A1(n1210), .A2(n1088), .A3(n1277), .ZN(n1275) );
INV_X1 U973 ( .A(KEYINPUT44), .ZN(n1277) );
XNOR2_X1 U974 ( .A(n1278), .B(G475), .ZN(n1088) );
NAND2_X1 U975 ( .A1(n1156), .A2(n1273), .ZN(n1278) );
XNOR2_X1 U976 ( .A(n1279), .B(n1280), .ZN(n1156) );
XNOR2_X1 U977 ( .A(G104), .B(n1281), .ZN(n1280) );
NAND2_X1 U978 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
OR2_X1 U979 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U980 ( .A(n1286), .B(KEYINPUT58), .Z(n1282) );
NAND2_X1 U981 ( .A1(n1284), .A2(n1285), .ZN(n1286) );
XNOR2_X1 U982 ( .A(n1287), .B(n1288), .ZN(n1284) );
AND2_X1 U983 ( .A1(n1289), .A2(G214), .ZN(n1288) );
XNOR2_X1 U984 ( .A(G131), .B(G143), .ZN(n1287) );
NAND2_X1 U985 ( .A1(KEYINPUT53), .A2(n1290), .ZN(n1279) );
XNOR2_X1 U986 ( .A(n1270), .B(G113), .ZN(n1290) );
INV_X1 U987 ( .A(G122), .ZN(n1270) );
INV_X1 U988 ( .A(n1251), .ZN(n1210) );
NOR2_X1 U989 ( .A1(n1092), .A2(n1291), .ZN(n1251) );
AND2_X1 U990 ( .A1(G478), .A2(n1095), .ZN(n1291) );
NOR2_X1 U991 ( .A1(n1095), .A2(G478), .ZN(n1092) );
NAND2_X1 U992 ( .A1(n1153), .A2(n1273), .ZN(n1095) );
XNOR2_X1 U993 ( .A(n1292), .B(n1293), .ZN(n1153) );
XOR2_X1 U994 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U995 ( .A(n1296), .B(n1297), .Z(n1295) );
NOR2_X1 U996 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NOR2_X1 U997 ( .A1(KEYINPUT22), .A2(G128), .ZN(n1296) );
XNOR2_X1 U998 ( .A(n1239), .B(G107), .ZN(n1294) );
XOR2_X1 U999 ( .A(n1300), .B(n1301), .Z(n1292) );
XNOR2_X1 U1000 ( .A(KEYINPUT59), .B(n1302), .ZN(n1301) );
XNOR2_X1 U1001 ( .A(G134), .B(G122), .ZN(n1300) );
NOR2_X1 U1002 ( .A1(n1055), .A2(n1303), .ZN(n1274) );
NOR2_X1 U1003 ( .A1(n1080), .A2(n1245), .ZN(n1303) );
NOR4_X1 U1004 ( .A1(n1304), .A2(n1273), .A3(n1305), .A4(G898), .ZN(n1245) );
INV_X1 U1005 ( .A(n1234), .ZN(n1305) );
XNOR2_X1 U1006 ( .A(n1120), .B(KEYINPUT20), .ZN(n1304) );
INV_X1 U1007 ( .A(n1052), .ZN(n1080) );
NAND3_X1 U1008 ( .A1(n1234), .A2(n1120), .A3(G952), .ZN(n1052) );
INV_X1 U1009 ( .A(G953), .ZN(n1120) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1234) );
INV_X1 U1011 ( .A(n1087), .ZN(n1055) );
NAND3_X1 U1012 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1087) );
NAND2_X1 U1013 ( .A1(n1309), .A2(n1148), .ZN(n1308) );
OR3_X1 U1014 ( .A1(n1148), .A2(n1309), .A3(G902), .ZN(n1307) );
NOR2_X1 U1015 ( .A1(n1298), .A2(G234), .ZN(n1309) );
INV_X1 U1016 ( .A(G217), .ZN(n1298) );
XOR2_X1 U1017 ( .A(n1310), .B(n1311), .Z(n1148) );
XOR2_X1 U1018 ( .A(n1312), .B(n1285), .Z(n1311) );
XNOR2_X1 U1019 ( .A(n1313), .B(n1115), .ZN(n1285) );
XNOR2_X1 U1020 ( .A(G140), .B(n1224), .ZN(n1115) );
INV_X1 U1021 ( .A(G125), .ZN(n1224) );
NOR2_X1 U1022 ( .A1(n1299), .A2(n1314), .ZN(n1312) );
INV_X1 U1023 ( .A(G221), .ZN(n1314) );
NAND2_X1 U1024 ( .A1(G234), .A2(n1272), .ZN(n1299) );
XNOR2_X1 U1025 ( .A(G137), .B(n1315), .ZN(n1310) );
NOR2_X1 U1026 ( .A1(KEYINPUT21), .A2(n1316), .ZN(n1315) );
XNOR2_X1 U1027 ( .A(G110), .B(n1317), .ZN(n1316) );
NOR2_X1 U1028 ( .A1(KEYINPUT38), .A2(n1318), .ZN(n1317) );
XNOR2_X1 U1029 ( .A(G119), .B(n1319), .ZN(n1318) );
NAND2_X1 U1030 ( .A1(KEYINPUT50), .A2(n1320), .ZN(n1319) );
NAND2_X1 U1031 ( .A1(G902), .A2(G217), .ZN(n1306) );
NOR2_X1 U1032 ( .A1(n1321), .A2(n1091), .ZN(n1236) );
NOR2_X1 U1033 ( .A1(n1093), .A2(G472), .ZN(n1091) );
AND2_X1 U1034 ( .A1(n1322), .A2(n1093), .ZN(n1321) );
NAND2_X1 U1035 ( .A1(n1323), .A2(n1273), .ZN(n1093) );
XOR2_X1 U1036 ( .A(n1162), .B(n1324), .Z(n1323) );
XNOR2_X1 U1037 ( .A(n1325), .B(n1326), .ZN(n1324) );
NOR2_X1 U1038 ( .A1(KEYINPUT17), .A2(n1163), .ZN(n1326) );
XOR2_X1 U1039 ( .A(n1327), .B(n1182), .Z(n1163) );
XOR2_X1 U1040 ( .A(n1328), .B(n1329), .Z(n1182) );
NOR2_X1 U1041 ( .A1(KEYINPUT55), .A2(n1302), .ZN(n1329) );
INV_X1 U1042 ( .A(G143), .ZN(n1302) );
XNOR2_X1 U1043 ( .A(G128), .B(G146), .ZN(n1328) );
NAND2_X1 U1044 ( .A1(n1330), .A2(KEYINPUT16), .ZN(n1325) );
XOR2_X1 U1045 ( .A(n1165), .B(KEYINPUT23), .Z(n1330) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1289), .ZN(n1165) );
NOR2_X1 U1047 ( .A1(n1331), .A2(G237), .ZN(n1289) );
XOR2_X1 U1048 ( .A(n1141), .B(G101), .Z(n1162) );
XNOR2_X1 U1049 ( .A(G113), .B(n1332), .ZN(n1141) );
XNOR2_X1 U1050 ( .A(G119), .B(n1239), .ZN(n1332) );
INV_X1 U1051 ( .A(G116), .ZN(n1239) );
XOR2_X1 U1052 ( .A(KEYINPUT27), .B(G472), .Z(n1322) );
NOR2_X1 U1053 ( .A1(n1078), .A2(n1077), .ZN(n1062) );
INV_X1 U1054 ( .A(n1246), .ZN(n1077) );
NAND2_X1 U1055 ( .A1(G221), .A2(n1333), .ZN(n1246) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1273), .ZN(n1333) );
NAND3_X1 U1057 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1078) );
NAND2_X1 U1058 ( .A1(G469), .A2(n1337), .ZN(n1336) );
OR3_X1 U1059 ( .A1(n1337), .A2(G469), .A3(KEYINPUT18), .ZN(n1335) );
OR2_X1 U1060 ( .A1(n1090), .A2(KEYINPUT63), .ZN(n1337) );
NAND2_X1 U1061 ( .A1(n1090), .A2(KEYINPUT18), .ZN(n1334) );
AND2_X1 U1062 ( .A1(n1338), .A2(n1273), .ZN(n1090) );
INV_X1 U1063 ( .A(G902), .ZN(n1273) );
XOR2_X1 U1064 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1065 ( .A(n1171), .B(n1341), .Z(n1340) );
NOR2_X1 U1066 ( .A1(KEYINPUT47), .A2(n1342), .ZN(n1341) );
XOR2_X1 U1067 ( .A(n1343), .B(n1108), .Z(n1342) );
XNOR2_X1 U1068 ( .A(n1344), .B(n1320), .ZN(n1108) );
INV_X1 U1069 ( .A(G128), .ZN(n1320) );
NAND3_X1 U1070 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1344) );
NAND2_X1 U1071 ( .A1(G146), .A2(n1348), .ZN(n1347) );
NAND2_X1 U1072 ( .A1(n1349), .A2(KEYINPUT61), .ZN(n1348) );
XNOR2_X1 U1073 ( .A(G143), .B(KEYINPUT48), .ZN(n1349) );
NAND3_X1 U1074 ( .A1(KEYINPUT61), .A2(n1313), .A3(G143), .ZN(n1346) );
INV_X1 U1075 ( .A(G146), .ZN(n1313) );
OR2_X1 U1076 ( .A1(G143), .A2(KEYINPUT61), .ZN(n1345) );
NAND2_X1 U1077 ( .A1(n1169), .A2(n1350), .ZN(n1343) );
XOR2_X1 U1078 ( .A(KEYINPUT43), .B(KEYINPUT36), .Z(n1350) );
XOR2_X1 U1079 ( .A(G101), .B(n1265), .Z(n1169) );
XNOR2_X1 U1080 ( .A(G104), .B(G107), .ZN(n1265) );
XOR2_X1 U1081 ( .A(n1327), .B(n1351), .Z(n1171) );
NOR2_X1 U1082 ( .A1(n1331), .A2(n1121), .ZN(n1351) );
INV_X1 U1083 ( .A(G227), .ZN(n1121) );
INV_X1 U1084 ( .A(n1272), .ZN(n1331) );
XOR2_X1 U1085 ( .A(G953), .B(KEYINPUT51), .Z(n1272) );
XNOR2_X1 U1086 ( .A(n1112), .B(KEYINPUT10), .ZN(n1327) );
XOR2_X1 U1087 ( .A(G131), .B(n1352), .Z(n1112) );
XOR2_X1 U1088 ( .A(G137), .B(G134), .Z(n1352) );
XNOR2_X1 U1089 ( .A(G110), .B(n1353), .ZN(n1339) );
XOR2_X1 U1090 ( .A(KEYINPUT8), .B(G140), .Z(n1353) );
INV_X1 U1091 ( .A(G110), .ZN(n1176) );
endmodule


