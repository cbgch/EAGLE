//Key = 1111101000010100101110011100111111011011111110100101111010010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300;

XNOR2_X1 U716 ( .A(G107), .B(n987), .ZN(G9) );
NOR2_X1 U717 ( .A1(n988), .A2(n989), .ZN(G75) );
XOR2_X1 U718 ( .A(KEYINPUT26), .B(n990), .Z(n989) );
NOR4_X1 U719 ( .A1(n991), .A2(n992), .A3(n993), .A4(n994), .ZN(n990) );
NOR2_X1 U720 ( .A1(n995), .A2(n996), .ZN(n993) );
INV_X1 U721 ( .A(n997), .ZN(n996) );
NOR2_X1 U722 ( .A1(n998), .A2(n999), .ZN(n995) );
NOR2_X1 U723 ( .A1(n1000), .A2(n1001), .ZN(n999) );
INV_X1 U724 ( .A(n1002), .ZN(n1001) );
NOR3_X1 U725 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1000) );
NOR2_X1 U726 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NOR3_X1 U727 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1006) );
NOR2_X1 U728 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
AND2_X1 U729 ( .A1(n1013), .A2(n1014), .ZN(n1009) );
NOR2_X1 U730 ( .A1(n1015), .A2(n1016), .ZN(n1008) );
NOR4_X1 U731 ( .A1(n1017), .A2(n1012), .A3(n1018), .A4(n1019), .ZN(n1004) );
XOR2_X1 U732 ( .A(n1007), .B(KEYINPUT60), .Z(n1017) );
NOR2_X1 U733 ( .A1(KEYINPUT28), .A2(n1020), .ZN(n1003) );
NOR2_X1 U734 ( .A1(n1021), .A2(n1020), .ZN(n998) );
INV_X1 U735 ( .A(n1022), .ZN(n1020) );
NOR2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR3_X1 U737 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1023) );
INV_X1 U738 ( .A(KEYINPUT28), .ZN(n1025) );
NAND4_X1 U739 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n991) );
NAND3_X1 U740 ( .A1(n1002), .A2(n1032), .A3(n1022), .ZN(n1028) );
NOR3_X1 U741 ( .A1(n1016), .A2(n1012), .A3(n1007), .ZN(n1022) );
INV_X1 U742 ( .A(n1033), .ZN(n1012) );
INV_X1 U743 ( .A(n1014), .ZN(n1016) );
NAND2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NAND2_X1 U745 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
INV_X1 U746 ( .A(n1038), .ZN(n1034) );
NOR3_X1 U747 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n988) );
INV_X1 U748 ( .A(n1030), .ZN(n1039) );
NAND4_X1 U749 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1030) );
NOR4_X1 U750 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
XOR2_X1 U751 ( .A(n1048), .B(G469), .Z(n1045) );
NAND2_X1 U752 ( .A1(KEYINPUT13), .A2(n1049), .ZN(n1048) );
XOR2_X1 U753 ( .A(n1050), .B(n1051), .Z(n1044) );
NAND2_X1 U754 ( .A1(n1052), .A2(KEYINPUT35), .ZN(n1050) );
XOR2_X1 U755 ( .A(n1053), .B(KEYINPUT12), .Z(n1052) );
AND3_X1 U756 ( .A1(n1027), .A2(n1019), .A3(n1054), .ZN(n1042) );
NAND2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1041) );
INV_X1 U758 ( .A(n1057), .ZN(n1056) );
XOR2_X1 U759 ( .A(n1058), .B(KEYINPUT39), .Z(n1055) );
XOR2_X1 U760 ( .A(n1059), .B(n1060), .Z(n1040) );
XNOR2_X1 U761 ( .A(G475), .B(KEYINPUT11), .ZN(n1060) );
XOR2_X1 U762 ( .A(n1061), .B(n1062), .Z(G72) );
NOR2_X1 U763 ( .A1(n1063), .A2(n1031), .ZN(n1062) );
AND2_X1 U764 ( .A1(G227), .A2(G900), .ZN(n1063) );
NAND2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NAND3_X1 U766 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NAND2_X1 U767 ( .A1(G953), .A2(n1069), .ZN(n1067) );
OR2_X1 U768 ( .A1(n1066), .A2(n1068), .ZN(n1064) );
NAND2_X1 U769 ( .A1(n1031), .A2(n1070), .ZN(n1068) );
NAND4_X1 U770 ( .A1(n1071), .A2(n1029), .A3(n1072), .A4(n1073), .ZN(n1070) );
NOR2_X1 U771 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
INV_X1 U772 ( .A(n1076), .ZN(n1074) );
XOR2_X1 U773 ( .A(n1077), .B(KEYINPUT43), .Z(n1066) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U776 ( .A(n1082), .B(KEYINPUT21), .Z(n1078) );
OR2_X1 U777 ( .A1(n1081), .A2(n1080), .ZN(n1082) );
NAND2_X1 U778 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NAND2_X1 U779 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U780 ( .A(n1087), .B(KEYINPUT37), .Z(n1083) );
OR2_X1 U781 ( .A1(n1086), .A2(n1085), .ZN(n1087) );
XNOR2_X1 U782 ( .A(n1088), .B(n1089), .ZN(n1086) );
NAND2_X1 U783 ( .A1(KEYINPUT46), .A2(n1090), .ZN(n1088) );
XOR2_X1 U784 ( .A(KEYINPUT23), .B(n1091), .Z(n1090) );
XOR2_X1 U785 ( .A(n1092), .B(n1093), .Z(G69) );
NOR2_X1 U786 ( .A1(n1094), .A2(n1031), .ZN(n1093) );
AND2_X1 U787 ( .A1(G224), .A2(G898), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NAND3_X1 U789 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NAND2_X1 U790 ( .A1(G953), .A2(n1100), .ZN(n1098) );
OR2_X1 U791 ( .A1(n1099), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U792 ( .A(n1101), .B(n1102), .ZN(n1097) );
NAND2_X1 U793 ( .A1(n1031), .A2(n1103), .ZN(n1099) );
NAND4_X1 U794 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1103) );
NOR2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U796 ( .A(KEYINPUT5), .B(n987), .ZN(n1109) );
NOR2_X1 U797 ( .A1(n1110), .A2(n1111), .ZN(G66) );
XNOR2_X1 U798 ( .A(n1112), .B(n1113), .ZN(n1111) );
NAND2_X1 U799 ( .A1(KEYINPUT38), .A2(n1114), .ZN(n1112) );
NAND2_X1 U800 ( .A1(n1115), .A2(n1051), .ZN(n1114) );
NOR2_X1 U801 ( .A1(n1110), .A2(n1116), .ZN(G63) );
XOR2_X1 U802 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U803 ( .A(KEYINPUT34), .B(n1119), .Z(n1118) );
AND2_X1 U804 ( .A1(G478), .A2(n1115), .ZN(n1119) );
NOR2_X1 U805 ( .A1(n1110), .A2(n1120), .ZN(G60) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U807 ( .A(KEYINPUT22), .B(n1123), .Z(n1122) );
AND2_X1 U808 ( .A1(G475), .A2(n1115), .ZN(n1123) );
NAND2_X1 U809 ( .A1(KEYINPUT49), .A2(n1124), .ZN(n1121) );
XOR2_X1 U810 ( .A(G104), .B(n1125), .Z(G6) );
NOR2_X1 U811 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1110), .A2(n1128), .ZN(G57) );
XOR2_X1 U813 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U814 ( .A(n1131), .B(n1132), .ZN(n1130) );
XNOR2_X1 U815 ( .A(n1133), .B(n1134), .ZN(n1129) );
XNOR2_X1 U816 ( .A(n1135), .B(n1136), .ZN(n1134) );
AND2_X1 U817 ( .A1(G472), .A2(n1115), .ZN(n1135) );
NOR2_X1 U818 ( .A1(n1110), .A2(n1137), .ZN(G54) );
XOR2_X1 U819 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U820 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U821 ( .A1(KEYINPUT58), .A2(n1133), .ZN(n1140) );
XOR2_X1 U822 ( .A(n1142), .B(n1143), .Z(n1138) );
AND2_X1 U823 ( .A1(G469), .A2(n1115), .ZN(n1143) );
INV_X1 U824 ( .A(n1144), .ZN(n1115) );
NAND2_X1 U825 ( .A1(n1145), .A2(KEYINPUT40), .ZN(n1142) );
XNOR2_X1 U826 ( .A(n1146), .B(n1147), .ZN(n1145) );
XNOR2_X1 U827 ( .A(n1148), .B(n1149), .ZN(n1147) );
NAND2_X1 U828 ( .A1(KEYINPUT4), .A2(n1150), .ZN(n1148) );
NOR2_X1 U829 ( .A1(n1110), .A2(n1151), .ZN(G51) );
XNOR2_X1 U830 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR2_X1 U831 ( .A1(n1058), .A2(n1144), .ZN(n1153) );
NAND2_X1 U832 ( .A1(G902), .A2(n1154), .ZN(n1144) );
NAND3_X1 U833 ( .A1(n1155), .A2(n1029), .A3(n1156), .ZN(n1154) );
XOR2_X1 U834 ( .A(n992), .B(KEYINPUT29), .Z(n1156) );
NAND3_X1 U835 ( .A1(n1157), .A2(n1106), .A3(n1158), .ZN(n992) );
AND3_X1 U836 ( .A1(n987), .A2(n1105), .A3(n1104), .ZN(n1158) );
NAND3_X1 U837 ( .A1(n1159), .A2(n1160), .A3(n997), .ZN(n987) );
NAND2_X1 U838 ( .A1(n1161), .A2(n1024), .ZN(n1106) );
XOR2_X1 U839 ( .A(n1127), .B(KEYINPUT44), .Z(n1161) );
NAND4_X1 U840 ( .A1(n1013), .A2(n997), .A3(n1162), .A4(n1160), .ZN(n1127) );
XOR2_X1 U841 ( .A(n1108), .B(KEYINPUT16), .Z(n1157) );
NAND4_X1 U842 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1108) );
NAND2_X1 U843 ( .A1(n1167), .A2(n1168), .ZN(n1029) );
XNOR2_X1 U844 ( .A(n1014), .B(KEYINPUT51), .ZN(n1167) );
INV_X1 U845 ( .A(n994), .ZN(n1155) );
NAND4_X1 U846 ( .A1(n1169), .A2(n1076), .A3(n1072), .A4(n1071), .ZN(n994) );
XNOR2_X1 U847 ( .A(KEYINPUT27), .B(n1075), .ZN(n1169) );
NAND4_X1 U848 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1075) );
NAND3_X1 U849 ( .A1(n1174), .A2(n1047), .A3(n1175), .ZN(n1170) );
INV_X1 U850 ( .A(n1176), .ZN(n1175) );
XNOR2_X1 U851 ( .A(KEYINPUT14), .B(n1011), .ZN(n1174) );
NOR2_X1 U852 ( .A1(n1031), .A2(G952), .ZN(n1110) );
XOR2_X1 U853 ( .A(G146), .B(n1177), .Z(G48) );
NOR3_X1 U854 ( .A1(n1176), .A2(n1036), .A3(n1011), .ZN(n1177) );
XNOR2_X1 U855 ( .A(G143), .B(n1171), .ZN(G45) );
NAND4_X1 U856 ( .A1(n1038), .A2(n1162), .A3(n1178), .A4(n1179), .ZN(n1171) );
AND3_X1 U857 ( .A1(n1024), .A2(n1180), .A3(n1046), .ZN(n1179) );
XNOR2_X1 U858 ( .A(n1172), .B(n1181), .ZN(G42) );
NOR2_X1 U859 ( .A1(KEYINPUT15), .A2(n1182), .ZN(n1181) );
INV_X1 U860 ( .A(G140), .ZN(n1182) );
NAND4_X1 U861 ( .A1(n1183), .A2(n1013), .A3(n1036), .A4(n1037), .ZN(n1172) );
XNOR2_X1 U862 ( .A(G137), .B(n1173), .ZN(G39) );
NAND3_X1 U863 ( .A1(n1184), .A2(n1033), .A3(n1183), .ZN(n1173) );
XNOR2_X1 U864 ( .A(G134), .B(n1076), .ZN(G36) );
NAND3_X1 U865 ( .A1(n1038), .A2(n1185), .A3(n1183), .ZN(n1076) );
XNOR2_X1 U866 ( .A(G131), .B(n1072), .ZN(G33) );
NAND3_X1 U867 ( .A1(n1013), .A2(n1038), .A3(n1183), .ZN(n1072) );
AND3_X1 U868 ( .A1(n1162), .A2(n1180), .A3(n1002), .ZN(n1183) );
NOR2_X1 U869 ( .A1(n1026), .A2(n1186), .ZN(n1002) );
INV_X1 U870 ( .A(n1027), .ZN(n1186) );
XNOR2_X1 U871 ( .A(G128), .B(n1071), .ZN(G30) );
NAND3_X1 U872 ( .A1(n1159), .A2(n1180), .A3(n1184), .ZN(n1071) );
NOR3_X1 U873 ( .A1(n1126), .A2(n1015), .A3(n1011), .ZN(n1159) );
INV_X1 U874 ( .A(n1185), .ZN(n1015) );
XNOR2_X1 U875 ( .A(G101), .B(n1104), .ZN(G3) );
NAND2_X1 U876 ( .A1(n1038), .A2(n1187), .ZN(n1104) );
XNOR2_X1 U877 ( .A(G125), .B(n1188), .ZN(G27) );
NAND2_X1 U878 ( .A1(n1168), .A2(n1014), .ZN(n1188) );
NOR2_X1 U879 ( .A1(n1176), .A2(n1047), .ZN(n1168) );
NAND4_X1 U880 ( .A1(n1013), .A2(n1024), .A3(n1037), .A4(n1180), .ZN(n1176) );
NAND2_X1 U881 ( .A1(n1007), .A2(n1189), .ZN(n1180) );
NAND4_X1 U882 ( .A1(G902), .A2(G953), .A3(n1190), .A4(n1069), .ZN(n1189) );
INV_X1 U883 ( .A(G900), .ZN(n1069) );
XNOR2_X1 U884 ( .A(G122), .B(n1191), .ZN(G24) );
NAND2_X1 U885 ( .A1(KEYINPUT6), .A2(n1192), .ZN(n1191) );
INV_X1 U886 ( .A(n1163), .ZN(n1192) );
NAND4_X1 U887 ( .A1(n1178), .A2(n1193), .A3(n997), .A4(n1046), .ZN(n1163) );
NOR2_X1 U888 ( .A1(n1037), .A2(n1047), .ZN(n997) );
XNOR2_X1 U889 ( .A(G119), .B(n1164), .ZN(G21) );
NAND3_X1 U890 ( .A1(n1193), .A2(n1033), .A3(n1184), .ZN(n1164) );
AND2_X1 U891 ( .A1(n1047), .A2(n1037), .ZN(n1184) );
XNOR2_X1 U892 ( .A(G116), .B(n1194), .ZN(G18) );
NAND2_X1 U893 ( .A1(KEYINPUT41), .A2(n1195), .ZN(n1194) );
INV_X1 U894 ( .A(n1165), .ZN(n1195) );
NAND3_X1 U895 ( .A1(n1038), .A2(n1185), .A3(n1193), .ZN(n1165) );
NOR2_X1 U896 ( .A1(n1178), .A2(n1196), .ZN(n1185) );
INV_X1 U897 ( .A(n1046), .ZN(n1196) );
XNOR2_X1 U898 ( .A(G113), .B(n1166), .ZN(G15) );
NAND3_X1 U899 ( .A1(n1013), .A2(n1038), .A3(n1193), .ZN(n1166) );
AND3_X1 U900 ( .A1(n1024), .A2(n1160), .A3(n1014), .ZN(n1193) );
NOR2_X1 U901 ( .A1(n1018), .A2(n1197), .ZN(n1014) );
INV_X1 U902 ( .A(n1019), .ZN(n1197) );
NOR2_X1 U903 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
NOR2_X1 U904 ( .A1(n1198), .A2(n1046), .ZN(n1013) );
XNOR2_X1 U905 ( .A(n1199), .B(n1105), .ZN(G12) );
NAND3_X1 U906 ( .A1(n1036), .A2(n1037), .A3(n1187), .ZN(n1105) );
AND4_X1 U907 ( .A1(n1033), .A2(n1162), .A3(n1024), .A4(n1160), .ZN(n1187) );
NAND2_X1 U908 ( .A1(n1007), .A2(n1200), .ZN(n1160) );
NAND4_X1 U909 ( .A1(G902), .A2(G953), .A3(n1190), .A4(n1100), .ZN(n1200) );
INV_X1 U910 ( .A(G898), .ZN(n1100) );
NAND3_X1 U911 ( .A1(n1190), .A2(n1031), .A3(G952), .ZN(n1007) );
INV_X1 U912 ( .A(G953), .ZN(n1031) );
NAND2_X1 U913 ( .A1(G237), .A2(G234), .ZN(n1190) );
INV_X1 U914 ( .A(n1126), .ZN(n1024) );
NAND2_X1 U915 ( .A1(n1027), .A2(n1026), .ZN(n1126) );
NAND2_X1 U916 ( .A1(n1201), .A2(n1054), .ZN(n1026) );
NAND2_X1 U917 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
OR2_X1 U918 ( .A1(n1058), .A2(n1057), .ZN(n1201) );
NOR2_X1 U919 ( .A1(n1202), .A2(G902), .ZN(n1057) );
INV_X1 U920 ( .A(n1152), .ZN(n1202) );
XNOR2_X1 U921 ( .A(n1203), .B(n1204), .ZN(n1152) );
XOR2_X1 U922 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U923 ( .A(n1207), .B(G125), .Z(n1206) );
NAND2_X1 U924 ( .A1(G224), .A2(n1208), .ZN(n1207) );
NAND2_X1 U925 ( .A1(KEYINPUT32), .A2(n1102), .ZN(n1205) );
XNOR2_X1 U926 ( .A(G122), .B(n1209), .ZN(n1102) );
XNOR2_X1 U927 ( .A(n1101), .B(n1136), .ZN(n1203) );
XNOR2_X1 U928 ( .A(n1210), .B(n1211), .ZN(n1101) );
XOR2_X1 U929 ( .A(n1212), .B(G113), .Z(n1210) );
NAND2_X1 U930 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XOR2_X1 U931 ( .A(KEYINPUT33), .B(n1215), .Z(n1213) );
NAND2_X1 U932 ( .A1(G210), .A2(n1216), .ZN(n1058) );
NAND2_X1 U933 ( .A1(G214), .A2(n1216), .ZN(n1027) );
NAND2_X1 U934 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
INV_X1 U935 ( .A(n1011), .ZN(n1162) );
NAND2_X1 U936 ( .A1(n1018), .A2(n1019), .ZN(n1011) );
NAND2_X1 U937 ( .A1(G221), .A2(n1219), .ZN(n1019) );
NAND2_X1 U938 ( .A1(n1220), .A2(n1221), .ZN(n1018) );
NAND2_X1 U939 ( .A1(G469), .A2(n1049), .ZN(n1221) );
XOR2_X1 U940 ( .A(n1222), .B(KEYINPUT48), .Z(n1220) );
OR2_X1 U941 ( .A1(n1049), .A2(G469), .ZN(n1222) );
NAND2_X1 U942 ( .A1(n1223), .A2(n1218), .ZN(n1049) );
XOR2_X1 U943 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U944 ( .A(n1226), .B(n1146), .ZN(n1225) );
NAND2_X1 U945 ( .A1(KEYINPUT19), .A2(n1149), .ZN(n1226) );
XOR2_X1 U946 ( .A(n1227), .B(n1150), .Z(n1224) );
NAND2_X1 U947 ( .A1(G227), .A2(n1208), .ZN(n1150) );
NAND2_X1 U948 ( .A1(KEYINPUT2), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U949 ( .A(n1141), .B(n1133), .ZN(n1228) );
INV_X1 U950 ( .A(n1229), .ZN(n1133) );
XNOR2_X1 U951 ( .A(n1085), .B(n1230), .ZN(n1141) );
NOR2_X1 U952 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XNOR2_X1 U953 ( .A(n1215), .B(KEYINPUT36), .ZN(n1232) );
NOR2_X1 U954 ( .A1(n1233), .A2(G101), .ZN(n1215) );
INV_X1 U955 ( .A(n1214), .ZN(n1231) );
NAND2_X1 U956 ( .A1(G101), .A2(n1233), .ZN(n1214) );
XOR2_X1 U957 ( .A(G104), .B(G107), .Z(n1233) );
XOR2_X1 U958 ( .A(n1234), .B(n1235), .Z(n1085) );
NAND2_X1 U959 ( .A1(KEYINPUT56), .A2(n1236), .ZN(n1234) );
NOR2_X1 U960 ( .A1(n1046), .A2(n1178), .ZN(n1033) );
INV_X1 U961 ( .A(n1198), .ZN(n1178) );
XOR2_X1 U962 ( .A(n1237), .B(n1059), .Z(n1198) );
NAND2_X1 U963 ( .A1(n1124), .A2(n1218), .ZN(n1059) );
XNOR2_X1 U964 ( .A(n1238), .B(n1239), .ZN(n1124) );
XOR2_X1 U965 ( .A(G122), .B(G113), .Z(n1239) );
XNOR2_X1 U966 ( .A(G104), .B(n1240), .ZN(n1238) );
NOR2_X1 U967 ( .A1(KEYINPUT10), .A2(n1241), .ZN(n1240) );
XOR2_X1 U968 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U969 ( .A(n1080), .B(n1244), .ZN(n1243) );
NOR2_X1 U970 ( .A1(G146), .A2(KEYINPUT7), .ZN(n1244) );
XOR2_X1 U971 ( .A(n1245), .B(n1246), .Z(n1242) );
AND4_X1 U972 ( .A1(n1247), .A2(n1217), .A3(n1208), .A4(G214), .ZN(n1246) );
INV_X1 U973 ( .A(KEYINPUT55), .ZN(n1247) );
XNOR2_X1 U974 ( .A(G131), .B(G143), .ZN(n1245) );
NAND2_X1 U975 ( .A1(n1248), .A2(KEYINPUT63), .ZN(n1237) );
XNOR2_X1 U976 ( .A(G475), .B(KEYINPUT8), .ZN(n1248) );
XNOR2_X1 U977 ( .A(n1249), .B(G478), .ZN(n1046) );
OR2_X1 U978 ( .A1(n1117), .A2(G902), .ZN(n1249) );
NAND2_X1 U979 ( .A1(n1250), .A2(n1251), .ZN(n1117) );
NAND2_X1 U980 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U981 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U982 ( .A1(KEYINPUT62), .A2(n1256), .ZN(n1255) );
INV_X1 U983 ( .A(n1257), .ZN(n1256) );
XOR2_X1 U984 ( .A(n1258), .B(KEYINPUT59), .Z(n1252) );
NAND2_X1 U985 ( .A1(n1257), .A2(n1259), .ZN(n1250) );
NAND2_X1 U986 ( .A1(KEYINPUT62), .A2(n1254), .ZN(n1259) );
XNOR2_X1 U987 ( .A(KEYINPUT61), .B(n1258), .ZN(n1254) );
NAND3_X1 U988 ( .A1(G234), .A2(n1208), .A3(G217), .ZN(n1258) );
XNOR2_X1 U989 ( .A(n1260), .B(n1261), .ZN(n1257) );
XOR2_X1 U990 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U991 ( .A(G116), .B(G107), .Z(n1263) );
XNOR2_X1 U992 ( .A(G122), .B(n1264), .ZN(n1260) );
XNOR2_X1 U993 ( .A(n1265), .B(G134), .ZN(n1264) );
XNOR2_X1 U994 ( .A(n1053), .B(n1051), .ZN(n1037) );
AND2_X1 U995 ( .A1(G217), .A2(n1219), .ZN(n1051) );
NAND2_X1 U996 ( .A1(G234), .A2(n1218), .ZN(n1219) );
NAND2_X1 U997 ( .A1(n1113), .A2(n1218), .ZN(n1053) );
XNOR2_X1 U998 ( .A(n1266), .B(n1267), .ZN(n1113) );
XNOR2_X1 U999 ( .A(G137), .B(n1268), .ZN(n1267) );
NAND3_X1 U1000 ( .A1(G234), .A2(n1208), .A3(G221), .ZN(n1268) );
NAND2_X1 U1001 ( .A1(n1269), .A2(KEYINPUT42), .ZN(n1266) );
XOR2_X1 U1002 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U1003 ( .A(n1272), .B(n1273), .ZN(n1271) );
XOR2_X1 U1004 ( .A(KEYINPUT25), .B(G146), .Z(n1273) );
INV_X1 U1005 ( .A(G119), .ZN(n1272) );
XNOR2_X1 U1006 ( .A(n1080), .B(n1274), .ZN(n1270) );
XOR2_X1 U1007 ( .A(n1275), .B(n1262), .Z(n1274) );
NOR2_X1 U1008 ( .A1(KEYINPUT47), .A2(n1209), .ZN(n1275) );
INV_X1 U1009 ( .A(n1146), .ZN(n1209) );
XOR2_X1 U1010 ( .A(G110), .B(KEYINPUT0), .Z(n1146) );
XNOR2_X1 U1011 ( .A(G125), .B(n1276), .ZN(n1080) );
INV_X1 U1012 ( .A(n1149), .ZN(n1276) );
XOR2_X1 U1013 ( .A(G140), .B(KEYINPUT9), .Z(n1149) );
INV_X1 U1014 ( .A(n1047), .ZN(n1036) );
XNOR2_X1 U1015 ( .A(n1277), .B(G472), .ZN(n1047) );
NAND2_X1 U1016 ( .A1(n1278), .A2(n1218), .ZN(n1277) );
INV_X1 U1017 ( .A(G902), .ZN(n1218) );
XNOR2_X1 U1018 ( .A(n1279), .B(n1280), .ZN(n1278) );
INV_X1 U1019 ( .A(n1131), .ZN(n1280) );
XNOR2_X1 U1020 ( .A(n1281), .B(G101), .ZN(n1131) );
NAND3_X1 U1021 ( .A1(n1208), .A2(n1217), .A3(G210), .ZN(n1281) );
INV_X1 U1022 ( .A(G237), .ZN(n1217) );
XOR2_X1 U1023 ( .A(G953), .B(KEYINPUT24), .Z(n1208) );
XNOR2_X1 U1024 ( .A(KEYINPUT3), .B(n1282), .ZN(n1279) );
NOR2_X1 U1025 ( .A1(KEYINPUT50), .A2(n1283), .ZN(n1282) );
XOR2_X1 U1026 ( .A(n1132), .B(n1284), .Z(n1283) );
XNOR2_X1 U1027 ( .A(n1285), .B(KEYINPUT1), .ZN(n1284) );
NAND2_X1 U1028 ( .A1(KEYINPUT31), .A2(n1286), .ZN(n1285) );
NAND3_X1 U1029 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1286) );
NAND2_X1 U1030 ( .A1(n1136), .A2(n1229), .ZN(n1289) );
NAND2_X1 U1031 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
INV_X1 U1032 ( .A(KEYINPUT52), .ZN(n1291) );
NAND2_X1 U1033 ( .A1(n1292), .A2(n1293), .ZN(n1290) );
XNOR2_X1 U1034 ( .A(n1229), .B(KEYINPUT45), .ZN(n1292) );
NAND2_X1 U1035 ( .A1(KEYINPUT52), .A2(n1294), .ZN(n1287) );
NAND2_X1 U1036 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
OR3_X1 U1037 ( .A1(n1136), .A2(n1229), .A3(KEYINPUT45), .ZN(n1296) );
INV_X1 U1038 ( .A(n1293), .ZN(n1136) );
XNOR2_X1 U1039 ( .A(n1297), .B(n1236), .ZN(n1293) );
XNOR2_X1 U1040 ( .A(n1265), .B(G146), .ZN(n1236) );
INV_X1 U1041 ( .A(G143), .ZN(n1265) );
NAND2_X1 U1042 ( .A1(KEYINPUT54), .A2(n1235), .ZN(n1297) );
XOR2_X1 U1043 ( .A(n1262), .B(KEYINPUT57), .Z(n1235) );
XOR2_X1 U1044 ( .A(G128), .B(KEYINPUT20), .Z(n1262) );
NAND2_X1 U1045 ( .A1(KEYINPUT45), .A2(n1229), .ZN(n1295) );
XOR2_X1 U1046 ( .A(n1091), .B(n1298), .Z(n1229) );
XOR2_X1 U1047 ( .A(KEYINPUT53), .B(n1089), .Z(n1298) );
XOR2_X1 U1048 ( .A(G134), .B(G137), .Z(n1089) );
XOR2_X1 U1049 ( .A(G131), .B(KEYINPUT30), .Z(n1091) );
XNOR2_X1 U1050 ( .A(G113), .B(n1299), .ZN(n1132) );
NOR2_X1 U1051 ( .A1(KEYINPUT17), .A2(n1211), .ZN(n1299) );
XNOR2_X1 U1052 ( .A(G116), .B(G119), .ZN(n1211) );
NAND2_X1 U1053 ( .A1(KEYINPUT18), .A2(n1300), .ZN(n1199) );
INV_X1 U1054 ( .A(G110), .ZN(n1300) );
endmodule


