//Key = 0101001000010101000100100001011110001100110100011010110101100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266;

XNOR2_X1 U692 ( .A(G107), .B(n962), .ZN(G9) );
OR2_X1 U693 ( .A1(n963), .A2(n964), .ZN(n962) );
NOR2_X1 U694 ( .A1(n965), .A2(n966), .ZN(G75) );
XOR2_X1 U695 ( .A(KEYINPUT63), .B(n967), .Z(n966) );
AND3_X1 U696 ( .A1(n968), .A2(n969), .A3(n970), .ZN(n967) );
NOR3_X1 U697 ( .A1(n971), .A2(n970), .A3(n972), .ZN(n965) );
INV_X1 U698 ( .A(G952), .ZN(n970) );
NAND3_X1 U699 ( .A1(n968), .A2(n969), .A3(n973), .ZN(n971) );
NAND2_X1 U700 ( .A1(n974), .A2(n975), .ZN(n973) );
NAND2_X1 U701 ( .A1(n976), .A2(n977), .ZN(n975) );
NAND3_X1 U702 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n977) );
NAND2_X1 U703 ( .A1(n981), .A2(n982), .ZN(n979) );
NAND2_X1 U704 ( .A1(n983), .A2(n984), .ZN(n982) );
OR2_X1 U705 ( .A1(n985), .A2(n986), .ZN(n984) );
NAND2_X1 U706 ( .A1(n987), .A2(n988), .ZN(n981) );
NAND2_X1 U707 ( .A1(n989), .A2(n990), .ZN(n988) );
NAND2_X1 U708 ( .A1(n991), .A2(n992), .ZN(n990) );
XNOR2_X1 U709 ( .A(KEYINPUT19), .B(n993), .ZN(n989) );
NAND3_X1 U710 ( .A1(n987), .A2(n994), .A3(n983), .ZN(n976) );
NAND2_X1 U711 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U712 ( .A1(n980), .A2(n997), .ZN(n996) );
NAND2_X1 U713 ( .A1(n963), .A2(n998), .ZN(n997) );
NAND2_X1 U714 ( .A1(n999), .A2(n1000), .ZN(n998) );
INV_X1 U715 ( .A(n1001), .ZN(n963) );
NAND2_X1 U716 ( .A1(n978), .A2(n1002), .ZN(n995) );
NAND2_X1 U717 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
INV_X1 U718 ( .A(n1005), .ZN(n1004) );
XOR2_X1 U719 ( .A(KEYINPUT36), .B(n1006), .Z(n1003) );
NAND4_X1 U720 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n968) );
NOR4_X1 U721 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
XOR2_X1 U722 ( .A(n1015), .B(n1016), .Z(n1014) );
NAND2_X1 U723 ( .A1(KEYINPUT15), .A2(G475), .ZN(n1016) );
XNOR2_X1 U724 ( .A(n1017), .B(n1018), .ZN(n1013) );
NOR2_X1 U725 ( .A1(n1019), .A2(n999), .ZN(n1009) );
NAND2_X1 U726 ( .A1(n1020), .A2(n1021), .ZN(n1008) );
XNOR2_X1 U727 ( .A(G478), .B(KEYINPUT30), .ZN(n1020) );
XOR2_X1 U728 ( .A(n1022), .B(n1023), .Z(G72) );
XOR2_X1 U729 ( .A(n1024), .B(n1025), .Z(n1023) );
NOR2_X1 U730 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
XNOR2_X1 U731 ( .A(KEYINPUT35), .B(n969), .ZN(n1027) );
NOR2_X1 U732 ( .A1(n1028), .A2(n1029), .ZN(n1024) );
XOR2_X1 U733 ( .A(n1030), .B(n1031), .Z(n1029) );
XOR2_X1 U734 ( .A(n1032), .B(n1033), .Z(n1031) );
XOR2_X1 U735 ( .A(n1034), .B(n1035), .Z(n1030) );
NOR2_X1 U736 ( .A1(G134), .A2(KEYINPUT24), .ZN(n1035) );
NAND2_X1 U737 ( .A1(n1036), .A2(KEYINPUT1), .ZN(n1034) );
XNOR2_X1 U738 ( .A(G125), .B(n1037), .ZN(n1036) );
NOR2_X1 U739 ( .A1(G140), .A2(KEYINPUT26), .ZN(n1037) );
NOR2_X1 U740 ( .A1(n1038), .A2(n969), .ZN(n1022) );
AND2_X1 U741 ( .A1(G227), .A2(G900), .ZN(n1038) );
NAND2_X1 U742 ( .A1(n1039), .A2(n1040), .ZN(G69) );
NAND2_X1 U743 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
XOR2_X1 U744 ( .A(KEYINPUT58), .B(n1043), .Z(n1039) );
NOR2_X1 U745 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
XOR2_X1 U746 ( .A(n1044), .B(n1045), .Z(n1041) );
NAND2_X1 U747 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U748 ( .A1(G953), .A2(n1048), .ZN(n1047) );
XNOR2_X1 U749 ( .A(KEYINPUT6), .B(n1049), .ZN(n1048) );
XOR2_X1 U750 ( .A(n1050), .B(n1051), .Z(n1046) );
NOR2_X1 U751 ( .A1(KEYINPUT7), .A2(n1052), .ZN(n1050) );
NAND2_X1 U752 ( .A1(n1053), .A2(n1054), .ZN(n1044) );
NAND3_X1 U753 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
XOR2_X1 U754 ( .A(KEYINPUT5), .B(n1058), .Z(n1055) );
XNOR2_X1 U755 ( .A(KEYINPUT57), .B(n969), .ZN(n1053) );
NAND2_X1 U756 ( .A1(G953), .A2(n1059), .ZN(n1042) );
NAND2_X1 U757 ( .A1(G898), .A2(G224), .ZN(n1059) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(G66) );
XNOR2_X1 U759 ( .A(n1062), .B(n1063), .ZN(n1061) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR2_X1 U761 ( .A1(n1060), .A2(n1066), .ZN(G63) );
XOR2_X1 U762 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U763 ( .A1(n1069), .A2(KEYINPUT46), .ZN(n1068) );
NAND2_X1 U764 ( .A1(n1070), .A2(G478), .ZN(n1067) );
NOR2_X1 U765 ( .A1(n1060), .A2(n1071), .ZN(G60) );
XNOR2_X1 U766 ( .A(n1072), .B(n1073), .ZN(n1071) );
AND2_X1 U767 ( .A1(G475), .A2(n1070), .ZN(n1073) );
XNOR2_X1 U768 ( .A(G104), .B(n1074), .ZN(G6) );
NOR2_X1 U769 ( .A1(n1075), .A2(n1076), .ZN(G57) );
XOR2_X1 U770 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U771 ( .A(n1079), .B(n1080), .Z(n1078) );
XNOR2_X1 U772 ( .A(n1081), .B(n1082), .ZN(n1080) );
NOR2_X1 U773 ( .A1(KEYINPUT25), .A2(n1083), .ZN(n1082) );
XNOR2_X1 U774 ( .A(n1084), .B(KEYINPUT17), .ZN(n1083) );
XOR2_X1 U775 ( .A(KEYINPUT32), .B(KEYINPUT13), .Z(n1079) );
XOR2_X1 U776 ( .A(n1085), .B(n1086), .Z(n1077) );
XOR2_X1 U777 ( .A(n1087), .B(n1088), .Z(n1086) );
XOR2_X1 U778 ( .A(n1089), .B(n1090), .Z(n1085) );
AND2_X1 U779 ( .A1(G472), .A2(n1070), .ZN(n1090) );
INV_X1 U780 ( .A(n1065), .ZN(n1070) );
NOR2_X1 U781 ( .A1(n1091), .A2(n969), .ZN(n1075) );
XNOR2_X1 U782 ( .A(G952), .B(KEYINPUT31), .ZN(n1091) );
NOR2_X1 U783 ( .A1(n1060), .A2(n1092), .ZN(G54) );
XOR2_X1 U784 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U785 ( .A1(n1095), .A2(n1065), .ZN(n1093) );
XNOR2_X1 U786 ( .A(G469), .B(KEYINPUT38), .ZN(n1095) );
NOR2_X1 U787 ( .A1(n1060), .A2(n1096), .ZN(G51) );
XOR2_X1 U788 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U789 ( .A1(n1099), .A2(n1065), .ZN(n1098) );
NAND2_X1 U790 ( .A1(n1100), .A2(n972), .ZN(n1065) );
NAND4_X1 U791 ( .A1(n1101), .A2(n1058), .A3(n1026), .A4(n1057), .ZN(n972) );
AND3_X1 U792 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1057) );
AND4_X1 U793 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1026) );
NOR4_X1 U794 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
INV_X1 U795 ( .A(n1113), .ZN(n1111) );
INV_X1 U796 ( .A(n1114), .ZN(n1109) );
AND2_X1 U797 ( .A1(n1115), .A2(n1116), .ZN(n1107) );
AND3_X1 U798 ( .A1(n1117), .A2(n1074), .A3(n1118), .ZN(n1058) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U801 ( .A(KEYINPUT37), .B(n985), .Z(n1121) );
NAND3_X1 U802 ( .A1(n1001), .A2(n1123), .A3(n1006), .ZN(n1074) );
NAND2_X1 U803 ( .A1(n1124), .A2(n1001), .ZN(n1117) );
XOR2_X1 U804 ( .A(n964), .B(KEYINPUT22), .Z(n1124) );
NAND2_X1 U805 ( .A1(n1005), .A2(n1123), .ZN(n964) );
AND3_X1 U806 ( .A1(n987), .A2(n1125), .A3(n1126), .ZN(n1123) );
XNOR2_X1 U807 ( .A(n1127), .B(KEYINPUT12), .ZN(n1101) );
XNOR2_X1 U808 ( .A(G902), .B(KEYINPUT48), .ZN(n1100) );
NOR2_X1 U809 ( .A1(KEYINPUT18), .A2(n1128), .ZN(n1097) );
XOR2_X1 U810 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U811 ( .A(n1131), .B(n1132), .ZN(n1130) );
NOR2_X1 U812 ( .A1(n969), .A2(G952), .ZN(n1060) );
XOR2_X1 U813 ( .A(n1112), .B(n1133), .Z(G48) );
XOR2_X1 U814 ( .A(KEYINPUT34), .B(G146), .Z(n1133) );
AND3_X1 U815 ( .A1(n1006), .A2(n1134), .A3(n1135), .ZN(n1112) );
XNOR2_X1 U816 ( .A(G143), .B(n1113), .ZN(G45) );
NAND3_X1 U817 ( .A1(n1136), .A2(n986), .A3(n1137), .ZN(n1113) );
NOR3_X1 U818 ( .A1(n993), .A2(n1138), .A3(n1139), .ZN(n1137) );
INV_X1 U819 ( .A(n1134), .ZN(n993) );
XNOR2_X1 U820 ( .A(G140), .B(n1105), .ZN(G42) );
NAND3_X1 U821 ( .A1(n985), .A2(n1006), .A3(n1140), .ZN(n1105) );
XNOR2_X1 U822 ( .A(G137), .B(n1106), .ZN(G39) );
NAND4_X1 U823 ( .A1(n1140), .A2(n980), .A3(n1141), .A4(n1012), .ZN(n1106) );
XNOR2_X1 U824 ( .A(G134), .B(n1116), .ZN(G36) );
NAND3_X1 U825 ( .A1(n1140), .A2(n1005), .A3(n986), .ZN(n1116) );
XNOR2_X1 U826 ( .A(G131), .B(n1115), .ZN(G33) );
NAND3_X1 U827 ( .A1(n1140), .A2(n1006), .A3(n986), .ZN(n1115) );
AND3_X1 U828 ( .A1(n1134), .A2(n1142), .A3(n978), .ZN(n1140) );
NOR2_X1 U829 ( .A1(n1143), .A2(n999), .ZN(n978) );
XOR2_X1 U830 ( .A(n1126), .B(KEYINPUT60), .Z(n1134) );
XNOR2_X1 U831 ( .A(n1144), .B(n1110), .ZN(G30) );
AND3_X1 U832 ( .A1(n1005), .A2(n1126), .A3(n1135), .ZN(n1110) );
AND3_X1 U833 ( .A1(n1141), .A2(n1012), .A3(n1136), .ZN(n1135) );
XNOR2_X1 U834 ( .A(n1081), .B(n1145), .ZN(G3) );
NOR4_X1 U835 ( .A1(n1146), .A2(n1147), .A3(KEYINPUT45), .A4(n1122), .ZN(n1145) );
INV_X1 U836 ( .A(n986), .ZN(n1122) );
NOR2_X1 U837 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
INV_X1 U838 ( .A(KEYINPUT42), .ZN(n1149) );
NOR2_X1 U839 ( .A1(n980), .A2(n1150), .ZN(n1148) );
NOR2_X1 U840 ( .A1(KEYINPUT42), .A2(n1119), .ZN(n1146) );
XNOR2_X1 U841 ( .A(G125), .B(n1114), .ZN(G27) );
NAND4_X1 U842 ( .A1(n1136), .A2(n985), .A3(n1006), .A4(n983), .ZN(n1114) );
AND2_X1 U843 ( .A1(n1001), .A2(n1142), .ZN(n1136) );
NAND2_X1 U844 ( .A1(n1151), .A2(n1152), .ZN(n1142) );
NAND3_X1 U845 ( .A1(G902), .A2(n1153), .A3(n1028), .ZN(n1152) );
AND2_X1 U846 ( .A1(n1154), .A2(G953), .ZN(n1028) );
XNOR2_X1 U847 ( .A(G900), .B(KEYINPUT56), .ZN(n1154) );
XNOR2_X1 U848 ( .A(n974), .B(KEYINPUT54), .ZN(n1151) );
INV_X1 U849 ( .A(n1155), .ZN(n974) );
NAND2_X1 U850 ( .A1(n1156), .A2(n1157), .ZN(G24) );
NAND2_X1 U851 ( .A1(n1127), .A2(n1158), .ZN(n1157) );
XOR2_X1 U852 ( .A(KEYINPUT47), .B(n1159), .Z(n1156) );
NOR2_X1 U853 ( .A1(n1127), .A2(n1158), .ZN(n1159) );
INV_X1 U854 ( .A(n1056), .ZN(n1127) );
NAND4_X1 U855 ( .A1(n1160), .A2(n987), .A3(n1161), .A4(n1162), .ZN(n1056) );
AND2_X1 U856 ( .A1(n1163), .A2(n1164), .ZN(n987) );
XNOR2_X1 U857 ( .A(KEYINPUT27), .B(n1007), .ZN(n1164) );
XOR2_X1 U858 ( .A(n1104), .B(n1165), .Z(G21) );
XNOR2_X1 U859 ( .A(G119), .B(KEYINPUT28), .ZN(n1165) );
NAND4_X1 U860 ( .A1(n1160), .A2(n980), .A3(n1141), .A4(n1012), .ZN(n1104) );
XOR2_X1 U861 ( .A(n1102), .B(n1166), .Z(G18) );
XOR2_X1 U862 ( .A(KEYINPUT53), .B(G116), .Z(n1166) );
NAND3_X1 U863 ( .A1(n986), .A2(n1005), .A3(n1160), .ZN(n1102) );
NOR2_X1 U864 ( .A1(n1161), .A2(n1138), .ZN(n1005) );
XNOR2_X1 U865 ( .A(G113), .B(n1103), .ZN(G15) );
NAND3_X1 U866 ( .A1(n986), .A2(n1006), .A3(n1160), .ZN(n1103) );
AND3_X1 U867 ( .A1(n1001), .A2(n1125), .A3(n983), .ZN(n1160) );
INV_X1 U868 ( .A(n1011), .ZN(n983) );
NAND2_X1 U869 ( .A1(n992), .A2(n1167), .ZN(n1011) );
NOR2_X1 U870 ( .A1(n1162), .A2(n1139), .ZN(n1006) );
INV_X1 U871 ( .A(n1161), .ZN(n1139) );
NOR2_X1 U872 ( .A1(n1012), .A2(n1007), .ZN(n986) );
INV_X1 U873 ( .A(n1141), .ZN(n1007) );
XNOR2_X1 U874 ( .A(n1168), .B(n1169), .ZN(G12) );
AND2_X1 U875 ( .A1(n985), .A2(n1119), .ZN(n1169) );
NOR2_X1 U876 ( .A1(n1150), .A2(n1170), .ZN(n1119) );
INV_X1 U877 ( .A(n980), .ZN(n1170) );
NOR2_X1 U878 ( .A1(n1162), .A2(n1161), .ZN(n980) );
XNOR2_X1 U879 ( .A(n1015), .B(G475), .ZN(n1161) );
NAND2_X1 U880 ( .A1(n1072), .A2(n1171), .ZN(n1015) );
XNOR2_X1 U881 ( .A(n1172), .B(G131), .ZN(n1072) );
XOR2_X1 U882 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U883 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U884 ( .A(n1158), .B(G113), .ZN(n1176) );
XNOR2_X1 U885 ( .A(KEYINPUT62), .B(n1131), .ZN(n1175) );
XOR2_X1 U886 ( .A(n1177), .B(n1178), .Z(n1173) );
XNOR2_X1 U887 ( .A(G104), .B(n1179), .ZN(n1178) );
NAND2_X1 U888 ( .A1(KEYINPUT11), .A2(n1180), .ZN(n1179) );
XOR2_X1 U889 ( .A(n1181), .B(n1182), .Z(n1177) );
NAND2_X1 U890 ( .A1(n1183), .A2(G214), .ZN(n1181) );
INV_X1 U891 ( .A(n1138), .ZN(n1162) );
NOR2_X1 U892 ( .A1(n1184), .A2(n1019), .ZN(n1138) );
NOR2_X1 U893 ( .A1(n1021), .A2(G478), .ZN(n1019) );
AND2_X1 U894 ( .A1(G478), .A2(n1021), .ZN(n1184) );
OR2_X1 U895 ( .A1(n1069), .A2(G902), .ZN(n1021) );
AND2_X1 U896 ( .A1(n1185), .A2(n1186), .ZN(n1069) );
NAND4_X1 U897 ( .A1(G234), .A2(G217), .A3(n1187), .A4(n969), .ZN(n1186) );
NAND2_X1 U898 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
NAND3_X1 U899 ( .A1(G217), .A2(n969), .A3(G234), .ZN(n1189) );
XNOR2_X1 U900 ( .A(n1187), .B(KEYINPUT49), .ZN(n1188) );
XNOR2_X1 U901 ( .A(n1190), .B(n1191), .ZN(n1187) );
XNOR2_X1 U902 ( .A(n1192), .B(G134), .ZN(n1191) );
INV_X1 U903 ( .A(G143), .ZN(n1192) );
XNOR2_X1 U904 ( .A(n1193), .B(n1144), .ZN(n1190) );
NAND2_X1 U905 ( .A1(n1194), .A2(KEYINPUT3), .ZN(n1193) );
XOR2_X1 U906 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U907 ( .A(KEYINPUT23), .B(n1158), .ZN(n1196) );
XNOR2_X1 U908 ( .A(G107), .B(G116), .ZN(n1195) );
NAND3_X1 U909 ( .A1(n1126), .A2(n1125), .A3(n1001), .ZN(n1150) );
NOR2_X1 U910 ( .A1(n1000), .A2(n999), .ZN(n1001) );
AND2_X1 U911 ( .A1(G214), .A2(n1197), .ZN(n999) );
INV_X1 U912 ( .A(n1143), .ZN(n1000) );
XNOR2_X1 U913 ( .A(n1017), .B(n1198), .ZN(n1143) );
XOR2_X1 U914 ( .A(KEYINPUT55), .B(n1199), .Z(n1198) );
NOR2_X1 U915 ( .A1(KEYINPUT21), .A2(n1018), .ZN(n1199) );
INV_X1 U916 ( .A(n1099), .ZN(n1018) );
NAND2_X1 U917 ( .A1(G210), .A2(n1197), .ZN(n1099) );
NAND2_X1 U918 ( .A1(n1200), .A2(n1171), .ZN(n1197) );
INV_X1 U919 ( .A(G237), .ZN(n1200) );
NAND3_X1 U920 ( .A1(n1201), .A2(n1202), .A3(n1171), .ZN(n1017) );
NAND3_X1 U921 ( .A1(n1132), .A2(n1203), .A3(n1204), .ZN(n1202) );
INV_X1 U922 ( .A(n1205), .ZN(n1204) );
NAND2_X1 U923 ( .A1(n1205), .A2(n1206), .ZN(n1201) );
NAND2_X1 U924 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U925 ( .A1(KEYINPUT29), .A2(n1209), .ZN(n1208) );
NAND2_X1 U926 ( .A1(n1132), .A2(n1203), .ZN(n1209) );
INV_X1 U927 ( .A(KEYINPUT20), .ZN(n1203) );
NAND2_X1 U928 ( .A1(n1132), .A2(n1210), .ZN(n1207) );
INV_X1 U929 ( .A(KEYINPUT29), .ZN(n1210) );
XOR2_X1 U930 ( .A(n1051), .B(n1211), .Z(n1132) );
NOR2_X1 U931 ( .A1(KEYINPUT14), .A2(n1212), .ZN(n1211) );
INV_X1 U932 ( .A(n1052), .ZN(n1212) );
XNOR2_X1 U933 ( .A(n1213), .B(n1214), .ZN(n1052) );
XOR2_X1 U934 ( .A(G116), .B(n1215), .Z(n1214) );
NOR2_X1 U935 ( .A1(KEYINPUT8), .A2(n1216), .ZN(n1215) );
XOR2_X1 U936 ( .A(KEYINPUT0), .B(G113), .Z(n1216) );
XNOR2_X1 U937 ( .A(G119), .B(KEYINPUT39), .ZN(n1213) );
XNOR2_X1 U938 ( .A(n1217), .B(n1218), .ZN(n1051) );
XNOR2_X1 U939 ( .A(KEYINPUT59), .B(n1081), .ZN(n1218) );
XOR2_X1 U940 ( .A(n1219), .B(n1220), .Z(n1217) );
NOR2_X1 U941 ( .A1(KEYINPUT16), .A2(n1221), .ZN(n1220) );
NAND2_X1 U942 ( .A1(n1222), .A2(n1223), .ZN(n1219) );
NAND2_X1 U943 ( .A1(G122), .A2(n1168), .ZN(n1223) );
XOR2_X1 U944 ( .A(n1224), .B(KEYINPUT9), .Z(n1222) );
NAND2_X1 U945 ( .A1(G110), .A2(n1158), .ZN(n1224) );
INV_X1 U946 ( .A(G122), .ZN(n1158) );
XNOR2_X1 U947 ( .A(n1225), .B(n1129), .ZN(n1205) );
XNOR2_X1 U948 ( .A(n1226), .B(n1088), .ZN(n1129) );
NAND2_X1 U949 ( .A1(G224), .A2(n969), .ZN(n1226) );
NAND2_X1 U950 ( .A1(KEYINPUT52), .A2(n1131), .ZN(n1225) );
INV_X1 U951 ( .A(G125), .ZN(n1131) );
NAND2_X1 U952 ( .A1(n1155), .A2(n1227), .ZN(n1125) );
NAND4_X1 U953 ( .A1(G953), .A2(G902), .A3(n1153), .A4(n1049), .ZN(n1227) );
INV_X1 U954 ( .A(G898), .ZN(n1049) );
NAND3_X1 U955 ( .A1(n1153), .A2(n969), .A3(G952), .ZN(n1155) );
NAND2_X1 U956 ( .A1(G237), .A2(G234), .ZN(n1153) );
NOR2_X1 U957 ( .A1(n992), .A2(n991), .ZN(n1126) );
INV_X1 U958 ( .A(n1167), .ZN(n991) );
NAND2_X1 U959 ( .A1(G221), .A2(n1228), .ZN(n1167) );
XOR2_X1 U960 ( .A(n1229), .B(G469), .Z(n992) );
NAND2_X1 U961 ( .A1(n1230), .A2(n1171), .ZN(n1229) );
XOR2_X1 U962 ( .A(KEYINPUT40), .B(n1094), .Z(n1230) );
XNOR2_X1 U963 ( .A(n1231), .B(n1232), .ZN(n1094) );
XOR2_X1 U964 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U965 ( .A(n1081), .B(n1235), .ZN(n1234) );
AND2_X1 U966 ( .A1(n969), .A2(G227), .ZN(n1235) );
XNOR2_X1 U967 ( .A(n1180), .B(G110), .ZN(n1233) );
XOR2_X1 U968 ( .A(n1032), .B(n1236), .Z(n1231) );
XNOR2_X1 U969 ( .A(n1084), .B(n1221), .ZN(n1236) );
XNOR2_X1 U970 ( .A(G104), .B(G107), .ZN(n1221) );
XNOR2_X1 U971 ( .A(n1237), .B(n1238), .ZN(n1032) );
NAND2_X1 U972 ( .A1(KEYINPUT41), .A2(n1144), .ZN(n1237) );
NOR2_X1 U973 ( .A1(n1141), .A2(n1163), .ZN(n985) );
INV_X1 U974 ( .A(n1012), .ZN(n1163) );
XOR2_X1 U975 ( .A(n1239), .B(n1064), .Z(n1012) );
NAND2_X1 U976 ( .A1(G217), .A2(n1228), .ZN(n1064) );
NAND2_X1 U977 ( .A1(G234), .A2(n1171), .ZN(n1228) );
NAND2_X1 U978 ( .A1(n1062), .A2(n1171), .ZN(n1239) );
XNOR2_X1 U979 ( .A(n1240), .B(n1241), .ZN(n1062) );
XOR2_X1 U980 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U981 ( .A(G110), .B(n1244), .ZN(n1243) );
NAND2_X1 U982 ( .A1(KEYINPUT43), .A2(n1245), .ZN(n1244) );
XOR2_X1 U983 ( .A(n1246), .B(n1247), .Z(n1245) );
XNOR2_X1 U984 ( .A(n1180), .B(G125), .ZN(n1247) );
INV_X1 U985 ( .A(G140), .ZN(n1180) );
XOR2_X1 U986 ( .A(G146), .B(n1248), .Z(n1246) );
XOR2_X1 U987 ( .A(KEYINPUT62), .B(KEYINPUT61), .Z(n1248) );
AND3_X1 U988 ( .A1(G221), .A2(n969), .A3(G234), .ZN(n1242) );
INV_X1 U989 ( .A(G953), .ZN(n969) );
XNOR2_X1 U990 ( .A(G119), .B(n1249), .ZN(n1240) );
XNOR2_X1 U991 ( .A(G137), .B(n1144), .ZN(n1249) );
INV_X1 U992 ( .A(G128), .ZN(n1144) );
XNOR2_X1 U993 ( .A(n1250), .B(G472), .ZN(n1141) );
NAND2_X1 U994 ( .A1(n1251), .A2(n1171), .ZN(n1250) );
INV_X1 U995 ( .A(G902), .ZN(n1171) );
XNOR2_X1 U996 ( .A(n1087), .B(n1252), .ZN(n1251) );
XOR2_X1 U997 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U998 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U999 ( .A(KEYINPUT33), .B(n1257), .Z(n1256) );
NOR2_X1 U1000 ( .A1(n1081), .A2(n1089), .ZN(n1257) );
AND2_X1 U1001 ( .A1(n1081), .A2(n1089), .ZN(n1255) );
NAND2_X1 U1002 ( .A1(n1183), .A2(G210), .ZN(n1089) );
NOR2_X1 U1003 ( .A1(G953), .A2(G237), .ZN(n1183) );
INV_X1 U1004 ( .A(G101), .ZN(n1081) );
NAND2_X1 U1005 ( .A1(n1258), .A2(n1259), .ZN(n1253) );
OR2_X1 U1006 ( .A1(n1084), .A2(n1088), .ZN(n1259) );
XOR2_X1 U1007 ( .A(n1260), .B(KEYINPUT44), .Z(n1258) );
NAND2_X1 U1008 ( .A1(n1084), .A2(n1088), .ZN(n1260) );
XOR2_X1 U1009 ( .A(G128), .B(n1261), .Z(n1088) );
NOR2_X1 U1010 ( .A1(KEYINPUT51), .A2(n1238), .ZN(n1261) );
XNOR2_X1 U1011 ( .A(n1182), .B(KEYINPUT2), .ZN(n1238) );
XOR2_X1 U1012 ( .A(G143), .B(G146), .Z(n1182) );
XNOR2_X1 U1013 ( .A(n1262), .B(n1033), .ZN(n1084) );
XOR2_X1 U1014 ( .A(G131), .B(G137), .Z(n1033) );
XNOR2_X1 U1015 ( .A(G134), .B(KEYINPUT4), .ZN(n1262) );
XNOR2_X1 U1016 ( .A(n1263), .B(n1264), .ZN(n1087) );
XOR2_X1 U1017 ( .A(G116), .B(n1265), .Z(n1264) );
NOR2_X1 U1018 ( .A1(G113), .A2(KEYINPUT10), .ZN(n1265) );
NAND2_X1 U1019 ( .A1(KEYINPUT50), .A2(n1266), .ZN(n1263) );
INV_X1 U1020 ( .A(G119), .ZN(n1266) );
INV_X1 U1021 ( .A(G110), .ZN(n1168) );
endmodule


