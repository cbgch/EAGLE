//Key = 0101101010011011101001010011010100100011000001011110101001101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335;

XNOR2_X1 U731 ( .A(G107), .B(n1004), .ZN(G9) );
NAND4_X1 U732 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
XNOR2_X1 U733 ( .A(n1009), .B(KEYINPUT47), .ZN(n1005) );
NOR2_X1 U734 ( .A1(n1010), .A2(n1011), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
XOR2_X1 U736 ( .A(KEYINPUT39), .B(n1016), .Z(n1013) );
NAND3_X1 U737 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1012) );
NAND2_X1 U738 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND3_X1 U739 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
XOR2_X1 U740 ( .A(KEYINPUT3), .B(n1025), .Z(n1024) );
NOR2_X1 U741 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND3_X1 U742 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1023) );
NAND2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NAND2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
OR2_X1 U745 ( .A1(n1035), .A2(n1007), .ZN(n1034) );
NAND2_X1 U746 ( .A1(n1036), .A2(n1006), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1022) );
INV_X1 U748 ( .A(n1027), .ZN(n1037) );
NAND3_X1 U749 ( .A1(n1036), .A2(n1033), .A3(n1030), .ZN(n1027) );
NAND4_X1 U750 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1017) );
AND3_X1 U751 ( .A1(n1030), .A2(n1028), .A3(n1036), .ZN(n1042) );
INV_X1 U752 ( .A(n1043), .ZN(n1030) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1040) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NAND2_X1 U755 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U756 ( .A1(n1050), .A2(n1051), .ZN(n1039) );
AND3_X1 U757 ( .A1(n1052), .A2(n1018), .A3(n1016), .ZN(n1010) );
NAND4_X1 U758 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1018) );
NOR4_X1 U759 ( .A1(n1050), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1056) );
NOR2_X1 U760 ( .A1(n1060), .A2(n1061), .ZN(n1055) );
XOR2_X1 U761 ( .A(n1062), .B(n1063), .Z(n1061) );
NAND2_X1 U762 ( .A1(KEYINPUT11), .A2(n1064), .ZN(n1063) );
XNOR2_X1 U763 ( .A(n1065), .B(KEYINPUT46), .ZN(n1054) );
XNOR2_X1 U764 ( .A(G478), .B(n1066), .ZN(n1053) );
XNOR2_X1 U765 ( .A(n1014), .B(KEYINPUT34), .ZN(n1052) );
XOR2_X1 U766 ( .A(n1067), .B(n1068), .Z(G72) );
XOR2_X1 U767 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U769 ( .A(n1073), .B(n1074), .Z(n1072) );
XNOR2_X1 U770 ( .A(n1075), .B(n1076), .ZN(n1074) );
NOR3_X1 U771 ( .A1(n1077), .A2(KEYINPUT32), .A3(n1078), .ZN(n1076) );
NOR2_X1 U772 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U773 ( .A(KEYINPUT19), .B(n1081), .Z(n1080) );
XOR2_X1 U774 ( .A(KEYINPUT5), .B(n1082), .Z(n1077) );
NOR2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U776 ( .A(KEYINPUT19), .B(n1081), .ZN(n1084) );
XNOR2_X1 U777 ( .A(n1085), .B(n1086), .ZN(n1073) );
NAND2_X1 U778 ( .A1(KEYINPUT38), .A2(n1087), .ZN(n1085) );
NOR2_X1 U779 ( .A1(G900), .A2(n1088), .ZN(n1071) );
NAND3_X1 U780 ( .A1(n1089), .A2(n1088), .A3(KEYINPUT26), .ZN(n1069) );
NAND2_X1 U781 ( .A1(G953), .A2(n1090), .ZN(n1067) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1090) );
NAND2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(G69) );
NAND2_X1 U784 ( .A1(G953), .A2(n1093), .ZN(n1092) );
NAND2_X1 U785 ( .A1(G898), .A2(n1094), .ZN(n1093) );
NAND2_X1 U786 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U787 ( .A(KEYINPUT14), .B(n1097), .Z(n1091) );
NOR2_X1 U788 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U789 ( .A(KEYINPUT22), .B(n1095), .Z(n1099) );
XNOR2_X1 U790 ( .A(n1100), .B(n1101), .ZN(n1095) );
XNOR2_X1 U791 ( .A(n1102), .B(n1103), .ZN(n1101) );
XOR2_X1 U792 ( .A(n1104), .B(KEYINPUT25), .Z(n1100) );
NAND2_X1 U793 ( .A1(n1088), .A2(n1105), .ZN(n1104) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U795 ( .A(n1108), .B(KEYINPUT59), .Z(n1106) );
NOR2_X1 U796 ( .A1(G224), .A2(n1088), .ZN(n1098) );
NOR3_X1 U797 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(G66) );
NOR3_X1 U798 ( .A1(n1112), .A2(G953), .A3(G952), .ZN(n1111) );
AND2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
INV_X1 U800 ( .A(KEYINPUT37), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(n1109) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U803 ( .A(G217), .B(KEYINPUT42), .ZN(n1116) );
NOR2_X1 U804 ( .A1(n1113), .A2(n1118), .ZN(G63) );
NOR3_X1 U805 ( .A1(n1066), .A2(n1119), .A3(n1120), .ZN(n1118) );
NOR3_X1 U806 ( .A1(n1121), .A2(n1122), .A3(n1117), .ZN(n1120) );
NOR2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1119) );
AND2_X1 U808 ( .A1(n1015), .A2(G478), .ZN(n1123) );
NOR2_X1 U809 ( .A1(n1113), .A2(n1125), .ZN(G60) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U811 ( .A(KEYINPUT1), .B(n1128), .Z(n1127) );
NOR2_X1 U812 ( .A1(n1129), .A2(n1117), .ZN(n1128) );
XNOR2_X1 U813 ( .A(G475), .B(KEYINPUT43), .ZN(n1129) );
XNOR2_X1 U814 ( .A(G104), .B(n1130), .ZN(G6) );
NAND3_X1 U815 ( .A1(n1008), .A2(n1131), .A3(n1132), .ZN(n1130) );
XOR2_X1 U816 ( .A(KEYINPUT36), .B(n1035), .Z(n1131) );
NOR2_X1 U817 ( .A1(n1113), .A2(n1133), .ZN(G57) );
XOR2_X1 U818 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U819 ( .A1(n1136), .A2(n1137), .ZN(n1134) );
NOR2_X1 U820 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U821 ( .A1(n1140), .A2(n1117), .ZN(n1139) );
NOR2_X1 U822 ( .A1(n1141), .A2(n1142), .ZN(n1138) );
NOR2_X1 U823 ( .A1(KEYINPUT41), .A2(n1143), .ZN(n1141) );
NOR2_X1 U824 ( .A1(n1144), .A2(n1145), .ZN(n1136) );
INV_X1 U825 ( .A(n1143), .ZN(n1145) );
XOR2_X1 U826 ( .A(n1146), .B(n1086), .Z(n1143) );
NOR2_X1 U827 ( .A1(n1147), .A2(KEYINPUT41), .ZN(n1144) );
NOR3_X1 U828 ( .A1(n1142), .A2(n1140), .A3(n1117), .ZN(n1147) );
INV_X1 U829 ( .A(KEYINPUT49), .ZN(n1142) );
NOR2_X1 U830 ( .A1(n1113), .A2(n1148), .ZN(G54) );
XOR2_X1 U831 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U832 ( .A1(n1151), .A2(n1117), .ZN(n1150) );
NOR3_X1 U833 ( .A1(n1152), .A2(KEYINPUT55), .A3(n1153), .ZN(n1149) );
NOR3_X1 U834 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
XNOR2_X1 U835 ( .A(n1157), .B(KEYINPUT62), .ZN(n1154) );
NOR2_X1 U836 ( .A1(n1158), .A2(n1157), .ZN(n1152) );
AND2_X1 U837 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U838 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U839 ( .A(n1163), .B(KEYINPUT0), .Z(n1159) );
NAND2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
INV_X1 U841 ( .A(n1161), .ZN(n1165) );
XNOR2_X1 U842 ( .A(n1162), .B(n1166), .ZN(n1164) );
XNOR2_X1 U843 ( .A(KEYINPUT33), .B(KEYINPUT15), .ZN(n1166) );
XNOR2_X1 U844 ( .A(n1167), .B(n1086), .ZN(n1162) );
NOR2_X1 U845 ( .A1(n1155), .A2(n1156), .ZN(n1158) );
AND2_X1 U846 ( .A1(n1168), .A2(n1169), .ZN(n1156) );
NOR2_X1 U847 ( .A1(n1113), .A2(n1170), .ZN(G51) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U849 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U850 ( .A1(n1175), .A2(n1117), .ZN(n1174) );
NAND2_X1 U851 ( .A1(G902), .A2(n1015), .ZN(n1117) );
NAND3_X1 U852 ( .A1(n1107), .A2(n1108), .A3(n1176), .ZN(n1015) );
INV_X1 U853 ( .A(n1089), .ZN(n1176) );
NAND4_X1 U854 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1089) );
AND4_X1 U855 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
NOR2_X1 U856 ( .A1(n1185), .A2(n1186), .ZN(n1179) );
AND3_X1 U857 ( .A1(n1036), .A2(n1187), .A3(n1188), .ZN(n1186) );
AND4_X1 U858 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1107) );
NOR3_X1 U859 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1192) );
INV_X1 U860 ( .A(n1196), .ZN(n1195) );
NAND2_X1 U861 ( .A1(n1132), .A2(n1197), .ZN(n1191) );
NAND2_X1 U862 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND3_X1 U863 ( .A1(n1038), .A2(n1200), .A3(n1036), .ZN(n1199) );
NAND2_X1 U864 ( .A1(n1007), .A2(n1008), .ZN(n1198) );
NAND4_X1 U865 ( .A1(n1035), .A2(n1006), .A3(n1008), .A4(n1201), .ZN(n1189) );
XNOR2_X1 U866 ( .A(KEYINPUT17), .B(n1045), .ZN(n1201) );
AND2_X1 U867 ( .A1(n1028), .A2(n1200), .ZN(n1008) );
NAND2_X1 U868 ( .A1(KEYINPUT63), .A2(n1202), .ZN(n1173) );
XNOR2_X1 U869 ( .A(n1203), .B(n1204), .ZN(n1202) );
NOR2_X1 U870 ( .A1(n1088), .A2(G952), .ZN(n1113) );
XOR2_X1 U871 ( .A(G146), .B(n1185), .Z(G48) );
AND3_X1 U872 ( .A1(n1205), .A2(n1035), .A3(n1187), .ZN(n1185) );
XNOR2_X1 U873 ( .A(G143), .B(n1177), .ZN(G45) );
NAND4_X1 U874 ( .A1(n1206), .A2(n1205), .A3(n1207), .A4(n1058), .ZN(n1177) );
XNOR2_X1 U875 ( .A(G140), .B(n1178), .ZN(G42) );
NAND3_X1 U876 ( .A1(n1038), .A2(n1035), .A3(n1188), .ZN(n1178) );
XOR2_X1 U877 ( .A(G137), .B(n1208), .Z(G39) );
NOR2_X1 U878 ( .A1(n1051), .A2(n1209), .ZN(n1208) );
XOR2_X1 U879 ( .A(KEYINPUT58), .B(n1210), .Z(n1209) );
NOR4_X1 U880 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
XNOR2_X1 U881 ( .A(KEYINPUT56), .B(n1215), .ZN(n1214) );
INV_X1 U882 ( .A(n1036), .ZN(n1213) );
XOR2_X1 U883 ( .A(n1184), .B(n1216), .Z(G36) );
NAND2_X1 U884 ( .A1(KEYINPUT50), .A2(G134), .ZN(n1216) );
NAND3_X1 U885 ( .A1(n1188), .A2(n1007), .A3(n1206), .ZN(n1184) );
XNOR2_X1 U886 ( .A(G131), .B(n1183), .ZN(G33) );
NAND3_X1 U887 ( .A1(n1188), .A2(n1035), .A3(n1206), .ZN(n1183) );
NOR3_X1 U888 ( .A1(n1211), .A2(n1217), .A3(n1051), .ZN(n1188) );
INV_X1 U889 ( .A(n1020), .ZN(n1051) );
NOR2_X1 U890 ( .A1(n1065), .A2(n1057), .ZN(n1020) );
XNOR2_X1 U891 ( .A(G128), .B(n1182), .ZN(G30) );
NAND3_X1 U892 ( .A1(n1205), .A2(n1007), .A3(n1187), .ZN(n1182) );
AND2_X1 U893 ( .A1(n1132), .A2(n1215), .ZN(n1205) );
XNOR2_X1 U894 ( .A(G101), .B(n1190), .ZN(G3) );
NAND4_X1 U895 ( .A1(n1036), .A2(n1206), .A3(n1132), .A4(n1200), .ZN(n1190) );
XNOR2_X1 U896 ( .A(G125), .B(n1181), .ZN(G27) );
NAND4_X1 U897 ( .A1(n1038), .A2(n1035), .A3(n1218), .A4(n1033), .ZN(n1181) );
NOR2_X1 U898 ( .A1(n1217), .A2(n1045), .ZN(n1218) );
INV_X1 U899 ( .A(n1215), .ZN(n1217) );
NAND2_X1 U900 ( .A1(n1043), .A2(n1219), .ZN(n1215) );
NAND4_X1 U901 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1221), .ZN(n1219) );
INV_X1 U902 ( .A(G900), .ZN(n1221) );
XNOR2_X1 U903 ( .A(G122), .B(n1108), .ZN(G24) );
NAND4_X1 U904 ( .A1(n1222), .A2(n1028), .A3(n1207), .A4(n1058), .ZN(n1108) );
NOR2_X1 U905 ( .A1(n1060), .A2(n1223), .ZN(n1028) );
XNOR2_X1 U906 ( .A(G119), .B(n1196), .ZN(G21) );
NAND3_X1 U907 ( .A1(n1187), .A2(n1222), .A3(n1036), .ZN(n1196) );
INV_X1 U908 ( .A(n1212), .ZN(n1187) );
NAND2_X1 U909 ( .A1(n1223), .A2(n1060), .ZN(n1212) );
INV_X1 U910 ( .A(n1224), .ZN(n1223) );
NAND2_X1 U911 ( .A1(n1225), .A2(n1226), .ZN(G18) );
NAND2_X1 U912 ( .A1(G116), .A2(n1227), .ZN(n1226) );
XOR2_X1 U913 ( .A(n1228), .B(KEYINPUT53), .Z(n1225) );
NAND2_X1 U914 ( .A1(n1193), .A2(n1229), .ZN(n1228) );
INV_X1 U915 ( .A(n1227), .ZN(n1193) );
NAND3_X1 U916 ( .A1(n1222), .A2(n1007), .A3(n1206), .ZN(n1227) );
NOR2_X1 U917 ( .A1(n1058), .A2(n1230), .ZN(n1007) );
XOR2_X1 U918 ( .A(n1194), .B(n1231), .Z(G15) );
NOR2_X1 U919 ( .A1(KEYINPUT7), .A2(n1232), .ZN(n1231) );
AND3_X1 U920 ( .A1(n1035), .A2(n1222), .A3(n1206), .ZN(n1194) );
INV_X1 U921 ( .A(n1026), .ZN(n1206) );
NAND2_X1 U922 ( .A1(n1060), .A2(n1224), .ZN(n1026) );
AND3_X1 U923 ( .A1(n1009), .A2(n1200), .A3(n1033), .ZN(n1222) );
AND2_X1 U924 ( .A1(n1041), .A2(n1049), .ZN(n1033) );
AND2_X1 U925 ( .A1(n1230), .A2(n1058), .ZN(n1035) );
XNOR2_X1 U926 ( .A(G110), .B(n1233), .ZN(G12) );
NAND4_X1 U927 ( .A1(n1036), .A2(n1132), .A3(n1038), .A4(n1234), .ZN(n1233) );
XNOR2_X1 U928 ( .A(KEYINPUT54), .B(n1200), .ZN(n1234) );
NAND2_X1 U929 ( .A1(n1043), .A2(n1235), .ZN(n1200) );
NAND4_X1 U930 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1236), .ZN(n1235) );
INV_X1 U931 ( .A(G898), .ZN(n1236) );
NAND3_X1 U932 ( .A1(n1237), .A2(n1220), .A3(n1016), .ZN(n1043) );
XOR2_X1 U933 ( .A(G953), .B(KEYINPUT57), .Z(n1016) );
NAND2_X1 U934 ( .A1(G237), .A2(G234), .ZN(n1220) );
XNOR2_X1 U935 ( .A(KEYINPUT24), .B(n1014), .ZN(n1237) );
INV_X1 U936 ( .A(G952), .ZN(n1014) );
NOR2_X1 U937 ( .A1(n1224), .A2(n1060), .ZN(n1038) );
XOR2_X1 U938 ( .A(n1238), .B(n1140), .Z(n1060) );
INV_X1 U939 ( .A(G472), .ZN(n1140) );
NAND2_X1 U940 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XOR2_X1 U941 ( .A(n1146), .B(n1241), .Z(n1240) );
XOR2_X1 U942 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR2_X1 U943 ( .A1(KEYINPUT51), .A2(n1204), .ZN(n1243) );
NAND2_X1 U944 ( .A1(KEYINPUT4), .A2(n1135), .ZN(n1242) );
AND2_X1 U945 ( .A1(n1244), .A2(n1245), .ZN(n1135) );
NAND2_X1 U946 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U947 ( .A1(G210), .A2(n1248), .ZN(n1246) );
NAND3_X1 U948 ( .A1(G210), .A2(n1248), .A3(G101), .ZN(n1244) );
XNOR2_X1 U949 ( .A(n1249), .B(n1161), .ZN(n1146) );
XNOR2_X1 U950 ( .A(n1250), .B(n1251), .ZN(n1249) );
NAND2_X1 U951 ( .A1(n1252), .A2(KEYINPUT52), .ZN(n1250) );
XNOR2_X1 U952 ( .A(n1253), .B(KEYINPUT18), .ZN(n1252) );
XNOR2_X1 U953 ( .A(G902), .B(KEYINPUT9), .ZN(n1239) );
XNOR2_X1 U954 ( .A(n1062), .B(n1254), .ZN(n1224) );
NOR2_X1 U955 ( .A1(n1064), .A2(KEYINPUT35), .ZN(n1254) );
NOR2_X1 U956 ( .A1(n1114), .A2(G902), .ZN(n1064) );
XOR2_X1 U957 ( .A(n1255), .B(n1256), .Z(n1114) );
XNOR2_X1 U958 ( .A(n1257), .B(n1258), .ZN(n1256) );
XNOR2_X1 U959 ( .A(G137), .B(n1259), .ZN(n1258) );
INV_X1 U960 ( .A(G119), .ZN(n1259) );
INV_X1 U961 ( .A(G110), .ZN(n1257) );
XOR2_X1 U962 ( .A(n1260), .B(n1261), .Z(n1255) );
NOR2_X1 U963 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NOR3_X1 U964 ( .A1(KEYINPUT8), .A2(G125), .A3(n1087), .ZN(n1263) );
NOR2_X1 U965 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
INV_X1 U966 ( .A(KEYINPUT8), .ZN(n1265) );
XOR2_X1 U967 ( .A(n1266), .B(n1267), .Z(n1260) );
NAND3_X1 U968 ( .A1(n1268), .A2(G221), .A3(KEYINPUT23), .ZN(n1266) );
NAND2_X1 U969 ( .A1(G217), .A2(n1269), .ZN(n1062) );
NOR2_X1 U970 ( .A1(n1211), .A2(n1045), .ZN(n1132) );
INV_X1 U971 ( .A(n1009), .ZN(n1045) );
NOR2_X1 U972 ( .A1(n1046), .A2(n1057), .ZN(n1009) );
INV_X1 U973 ( .A(n1048), .ZN(n1057) );
NAND2_X1 U974 ( .A1(G214), .A2(n1270), .ZN(n1048) );
INV_X1 U975 ( .A(n1065), .ZN(n1046) );
XOR2_X1 U976 ( .A(n1271), .B(n1175), .Z(n1065) );
NAND2_X1 U977 ( .A1(G210), .A2(n1270), .ZN(n1175) );
NAND2_X1 U978 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
INV_X1 U979 ( .A(G237), .ZN(n1272) );
NAND3_X1 U980 ( .A1(n1274), .A2(n1273), .A3(n1275), .ZN(n1271) );
NAND2_X1 U981 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U982 ( .A(KEYINPUT12), .B(n1204), .ZN(n1276) );
NAND2_X1 U983 ( .A1(n1278), .A2(n1279), .ZN(n1274) );
XNOR2_X1 U984 ( .A(KEYINPUT40), .B(n1277), .ZN(n1279) );
XNOR2_X1 U985 ( .A(n1171), .B(n1203), .ZN(n1277) );
XNOR2_X1 U986 ( .A(G125), .B(KEYINPUT30), .ZN(n1203) );
XOR2_X1 U987 ( .A(n1280), .B(n1102), .Z(n1171) );
XOR2_X1 U988 ( .A(G110), .B(G122), .Z(n1102) );
XOR2_X1 U989 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U990 ( .A1(G953), .A2(n1096), .ZN(n1282) );
INV_X1 U991 ( .A(G224), .ZN(n1096) );
NAND2_X1 U992 ( .A1(KEYINPUT6), .A2(n1103), .ZN(n1281) );
XOR2_X1 U993 ( .A(n1283), .B(n1284), .Z(n1103) );
NOR3_X1 U994 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1284) );
NOR2_X1 U995 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NOR3_X1 U996 ( .A1(G107), .A2(KEYINPUT10), .A3(n1290), .ZN(n1286) );
INV_X1 U997 ( .A(n1288), .ZN(n1290) );
NOR2_X1 U998 ( .A1(KEYINPUT2), .A2(n1291), .ZN(n1288) );
AND2_X1 U999 ( .A1(n1291), .A2(KEYINPUT10), .ZN(n1285) );
XNOR2_X1 U1000 ( .A(n1292), .B(n1247), .ZN(n1283) );
NAND2_X1 U1001 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NAND2_X1 U1002 ( .A1(n1251), .A2(n1253), .ZN(n1294) );
XOR2_X1 U1003 ( .A(KEYINPUT31), .B(n1295), .Z(n1293) );
NOR2_X1 U1004 ( .A1(n1251), .A2(n1253), .ZN(n1295) );
XNOR2_X1 U1005 ( .A(G119), .B(n1229), .ZN(n1253) );
XNOR2_X1 U1006 ( .A(KEYINPUT12), .B(n1086), .ZN(n1278) );
INV_X1 U1007 ( .A(n1006), .ZN(n1211) );
NOR2_X1 U1008 ( .A1(n1041), .A2(n1050), .ZN(n1006) );
INV_X1 U1009 ( .A(n1049), .ZN(n1050) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1269), .ZN(n1049) );
NAND2_X1 U1011 ( .A1(G234), .A2(n1273), .ZN(n1269) );
XOR2_X1 U1012 ( .A(n1059), .B(KEYINPUT21), .Z(n1041) );
XOR2_X1 U1013 ( .A(n1296), .B(n1151), .Z(n1059) );
INV_X1 U1014 ( .A(G469), .ZN(n1151) );
NAND2_X1 U1015 ( .A1(n1297), .A2(n1273), .ZN(n1296) );
XNOR2_X1 U1016 ( .A(n1298), .B(n1161), .ZN(n1297) );
XOR2_X1 U1017 ( .A(n1081), .B(n1083), .Z(n1161) );
INV_X1 U1018 ( .A(n1079), .ZN(n1083) );
XOR2_X1 U1019 ( .A(G131), .B(KEYINPUT20), .Z(n1079) );
XOR2_X1 U1020 ( .A(G134), .B(G137), .Z(n1081) );
XOR2_X1 U1021 ( .A(n1299), .B(n1300), .Z(n1298) );
NOR2_X1 U1022 ( .A1(n1155), .A2(n1301), .ZN(n1300) );
NOR2_X1 U1023 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XOR2_X1 U1024 ( .A(n1169), .B(KEYINPUT61), .Z(n1303) );
INV_X1 U1025 ( .A(n1168), .ZN(n1302) );
NOR2_X1 U1026 ( .A1(n1169), .A2(n1168), .ZN(n1155) );
XNOR2_X1 U1027 ( .A(G110), .B(n1087), .ZN(n1168) );
INV_X1 U1028 ( .A(G140), .ZN(n1087) );
NAND2_X1 U1029 ( .A1(G227), .A2(n1088), .ZN(n1169) );
NAND2_X1 U1030 ( .A1(n1304), .A2(n1305), .ZN(n1299) );
NAND2_X1 U1031 ( .A1(n1204), .A2(n1306), .ZN(n1305) );
NAND2_X1 U1032 ( .A1(n1167), .A2(n1307), .ZN(n1306) );
NAND2_X1 U1033 ( .A1(KEYINPUT44), .A2(KEYINPUT29), .ZN(n1307) );
NAND3_X1 U1034 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1304) );
INV_X1 U1035 ( .A(KEYINPUT44), .ZN(n1310) );
NAND2_X1 U1036 ( .A1(KEYINPUT29), .A2(n1311), .ZN(n1309) );
NAND2_X1 U1037 ( .A1(n1086), .A2(n1167), .ZN(n1311) );
INV_X1 U1038 ( .A(n1204), .ZN(n1086) );
XOR2_X1 U1039 ( .A(G143), .B(n1267), .Z(n1204) );
XOR2_X1 U1040 ( .A(G128), .B(G146), .Z(n1267) );
OR2_X1 U1041 ( .A1(n1312), .A2(KEYINPUT29), .ZN(n1308) );
INV_X1 U1042 ( .A(n1167), .ZN(n1312) );
XNOR2_X1 U1043 ( .A(n1313), .B(n1314), .ZN(n1167) );
XNOR2_X1 U1044 ( .A(KEYINPUT28), .B(n1289), .ZN(n1314) );
XNOR2_X1 U1045 ( .A(n1315), .B(n1247), .ZN(n1313) );
INV_X1 U1046 ( .A(G101), .ZN(n1247) );
NAND2_X1 U1047 ( .A1(KEYINPUT60), .A2(n1316), .ZN(n1315) );
NOR2_X1 U1048 ( .A1(n1058), .A2(n1207), .ZN(n1036) );
INV_X1 U1049 ( .A(n1230), .ZN(n1207) );
XNOR2_X1 U1050 ( .A(n1317), .B(n1066), .ZN(n1230) );
NOR2_X1 U1051 ( .A1(n1124), .A2(G902), .ZN(n1066) );
INV_X1 U1052 ( .A(n1121), .ZN(n1124) );
XNOR2_X1 U1053 ( .A(n1318), .B(n1319), .ZN(n1121) );
XOR2_X1 U1054 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1055 ( .A(n1289), .B(n1322), .ZN(n1321) );
NOR2_X1 U1056 ( .A1(KEYINPUT13), .A2(n1323), .ZN(n1322) );
XNOR2_X1 U1057 ( .A(G122), .B(n1324), .ZN(n1323) );
NAND2_X1 U1058 ( .A1(KEYINPUT27), .A2(n1229), .ZN(n1324) );
INV_X1 U1059 ( .A(G116), .ZN(n1229) );
INV_X1 U1060 ( .A(G107), .ZN(n1289) );
AND2_X1 U1061 ( .A1(n1268), .A2(G217), .ZN(n1320) );
AND2_X1 U1062 ( .A1(G234), .A2(n1088), .ZN(n1268) );
INV_X1 U1063 ( .A(G953), .ZN(n1088) );
XNOR2_X1 U1064 ( .A(G128), .B(n1325), .ZN(n1318) );
XNOR2_X1 U1065 ( .A(n1326), .B(G134), .ZN(n1325) );
NAND2_X1 U1066 ( .A1(KEYINPUT45), .A2(n1122), .ZN(n1317) );
INV_X1 U1067 ( .A(G478), .ZN(n1122) );
XNOR2_X1 U1068 ( .A(n1327), .B(G475), .ZN(n1058) );
NAND2_X1 U1069 ( .A1(n1126), .A2(n1273), .ZN(n1327) );
INV_X1 U1070 ( .A(G902), .ZN(n1273) );
XNOR2_X1 U1071 ( .A(n1328), .B(n1329), .ZN(n1126) );
XOR2_X1 U1072 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1073 ( .A(n1332), .B(G122), .ZN(n1331) );
INV_X1 U1074 ( .A(G131), .ZN(n1332) );
XNOR2_X1 U1075 ( .A(G146), .B(n1326), .ZN(n1330) );
INV_X1 U1076 ( .A(G143), .ZN(n1326) );
XOR2_X1 U1077 ( .A(n1333), .B(n1334), .Z(n1328) );
XNOR2_X1 U1078 ( .A(n1291), .B(n1264), .ZN(n1334) );
XNOR2_X1 U1079 ( .A(n1075), .B(G140), .ZN(n1264) );
INV_X1 U1080 ( .A(G125), .ZN(n1075) );
INV_X1 U1081 ( .A(n1316), .ZN(n1291) );
XOR2_X1 U1082 ( .A(G104), .B(KEYINPUT48), .Z(n1316) );
XNOR2_X1 U1083 ( .A(n1335), .B(n1251), .ZN(n1333) );
XOR2_X1 U1084 ( .A(n1232), .B(KEYINPUT16), .Z(n1251) );
INV_X1 U1085 ( .A(G113), .ZN(n1232) );
NAND2_X1 U1086 ( .A1(G214), .A2(n1248), .ZN(n1335) );
NOR2_X1 U1087 ( .A1(G953), .A2(G237), .ZN(n1248) );
endmodule


