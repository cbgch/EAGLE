//Key = 1010111010100000111010010000000111000101001100000100011010001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;

XNOR2_X1 U769 ( .A(n1059), .B(n1060), .ZN(G9) );
NOR2_X1 U770 ( .A1(n1061), .A2(n1062), .ZN(G75) );
NOR4_X1 U771 ( .A1(G953), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1062) );
NOR2_X1 U772 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U773 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR3_X1 U774 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NOR2_X1 U775 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U776 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U778 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(n1073) );
NOR2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR3_X1 U781 ( .A1(n1082), .A2(n1085), .A3(n1086), .ZN(n1068) );
NOR3_X1 U782 ( .A1(n1076), .A2(n1087), .A3(n1088), .ZN(n1086) );
NOR2_X1 U783 ( .A1(n1089), .A2(n1072), .ZN(n1088) );
NOR2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U786 ( .A1(n1094), .A2(n1070), .ZN(n1087) );
NOR2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U788 ( .A(KEYINPUT34), .B(n1097), .Z(n1096) );
NOR2_X1 U789 ( .A1(KEYINPUT3), .A2(n1098), .ZN(n1095) );
NOR2_X1 U790 ( .A1(n1099), .A2(n1100), .ZN(n1085) );
AND3_X1 U791 ( .A1(KEYINPUT3), .A2(n1101), .A3(n1102), .ZN(n1100) );
INV_X1 U792 ( .A(n1103), .ZN(n1082) );
NOR3_X1 U793 ( .A1(n1063), .A2(G953), .A3(G952), .ZN(n1061) );
AND4_X1 U794 ( .A1(n1099), .A2(n1104), .A3(n1103), .A4(n1105), .ZN(n1063) );
NOR4_X1 U795 ( .A1(n1106), .A2(n1107), .A3(n1070), .A4(n1108), .ZN(n1105) );
XNOR2_X1 U796 ( .A(G475), .B(n1109), .ZN(n1108) );
NOR3_X1 U797 ( .A1(n1110), .A2(KEYINPUT50), .A3(n1111), .ZN(n1107) );
AND2_X1 U798 ( .A1(n1110), .A2(KEYINPUT50), .ZN(n1106) );
XOR2_X1 U799 ( .A(n1112), .B(n1113), .Z(G72) );
NOR2_X1 U800 ( .A1(KEYINPUT59), .A2(n1114), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U804 ( .A(KEYINPUT4), .B(n1121), .ZN(n1120) );
NAND2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1115) );
NAND2_X1 U806 ( .A1(G953), .A2(n1124), .ZN(n1123) );
XNOR2_X1 U807 ( .A(n1125), .B(n1126), .ZN(n1122) );
XOR2_X1 U808 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U810 ( .A(KEYINPUT25), .B(n1131), .Z(n1130) );
NOR2_X1 U811 ( .A1(G131), .A2(n1132), .ZN(n1131) );
AND2_X1 U812 ( .A1(n1132), .A2(G131), .ZN(n1129) );
NAND2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
OR2_X1 U814 ( .A1(n1135), .A2(G137), .ZN(n1134) );
XOR2_X1 U815 ( .A(n1136), .B(KEYINPUT13), .Z(n1133) );
NAND2_X1 U816 ( .A1(G137), .A2(n1135), .ZN(n1136) );
NOR2_X1 U817 ( .A1(KEYINPUT30), .A2(n1137), .ZN(n1127) );
NAND2_X1 U818 ( .A1(G953), .A2(n1138), .ZN(n1112) );
NAND2_X1 U819 ( .A1(G900), .A2(G227), .ZN(n1138) );
XOR2_X1 U820 ( .A(n1139), .B(n1140), .Z(G69) );
NAND2_X1 U821 ( .A1(G953), .A2(n1141), .ZN(n1140) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1141) );
NAND2_X1 U823 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
NAND2_X1 U824 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U825 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
OR2_X1 U826 ( .A1(n1148), .A2(KEYINPUT27), .ZN(n1147) );
NAND2_X1 U827 ( .A1(G953), .A2(n1149), .ZN(n1146) );
NAND2_X1 U828 ( .A1(n1150), .A2(n1148), .ZN(n1142) );
NAND2_X1 U829 ( .A1(n1117), .A2(n1151), .ZN(n1148) );
NAND2_X1 U830 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XNOR2_X1 U831 ( .A(KEYINPUT0), .B(n1154), .ZN(n1153) );
NAND2_X1 U832 ( .A1(n1144), .A2(n1155), .ZN(n1150) );
INV_X1 U833 ( .A(KEYINPUT27), .ZN(n1155) );
XOR2_X1 U834 ( .A(KEYINPUT60), .B(n1156), .Z(n1144) );
NOR2_X1 U835 ( .A1(n1157), .A2(n1158), .ZN(G66) );
XOR2_X1 U836 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR3_X1 U837 ( .A1(n1161), .A2(KEYINPUT52), .A3(n1162), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1157), .A2(n1163), .ZN(G63) );
XOR2_X1 U839 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U840 ( .A(n1166), .B(KEYINPUT36), .Z(n1164) );
NAND2_X1 U841 ( .A1(n1167), .A2(G478), .ZN(n1166) );
NOR3_X1 U842 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(G60) );
AND3_X1 U843 ( .A1(KEYINPUT7), .A2(n1171), .A3(G952), .ZN(n1170) );
NOR2_X1 U844 ( .A1(KEYINPUT7), .A2(n1172), .ZN(n1169) );
XOR2_X1 U845 ( .A(n1173), .B(n1174), .Z(n1168) );
NAND2_X1 U846 ( .A1(n1167), .A2(G475), .ZN(n1173) );
NAND2_X1 U847 ( .A1(n1175), .A2(n1176), .ZN(G6) );
OR2_X1 U848 ( .A1(G104), .A2(KEYINPUT17), .ZN(n1176) );
XOR2_X1 U849 ( .A(n1177), .B(n1178), .Z(n1175) );
NOR2_X1 U850 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND2_X1 U851 ( .A1(KEYINPUT17), .A2(G104), .ZN(n1177) );
NOR2_X1 U852 ( .A1(n1157), .A2(n1181), .ZN(G57) );
XOR2_X1 U853 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U854 ( .A(n1184), .B(n1185), .ZN(n1183) );
XOR2_X1 U855 ( .A(n1186), .B(n1187), .Z(n1182) );
XOR2_X1 U856 ( .A(n1188), .B(n1189), .Z(n1186) );
NAND2_X1 U857 ( .A1(n1167), .A2(G472), .ZN(n1188) );
NOR2_X1 U858 ( .A1(n1157), .A2(n1190), .ZN(G54) );
XOR2_X1 U859 ( .A(n1191), .B(n1192), .Z(n1190) );
AND2_X1 U860 ( .A1(G469), .A2(n1167), .ZN(n1192) );
NAND2_X1 U861 ( .A1(KEYINPUT33), .A2(n1193), .ZN(n1191) );
NAND2_X1 U862 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U863 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U864 ( .A(n1198), .B(KEYINPUT38), .Z(n1194) );
OR2_X1 U865 ( .A1(n1197), .A2(n1196), .ZN(n1198) );
XOR2_X1 U866 ( .A(n1199), .B(n1200), .Z(n1196) );
XNOR2_X1 U867 ( .A(KEYINPUT18), .B(n1201), .ZN(n1200) );
XOR2_X1 U868 ( .A(n1202), .B(n1203), .Z(n1199) );
NAND2_X1 U869 ( .A1(KEYINPUT42), .A2(n1204), .ZN(n1202) );
XNOR2_X1 U870 ( .A(n1205), .B(n1187), .ZN(n1197) );
NAND2_X1 U871 ( .A1(n1206), .A2(KEYINPUT6), .ZN(n1205) );
XNOR2_X1 U872 ( .A(n1207), .B(n1125), .ZN(n1206) );
INV_X1 U873 ( .A(n1172), .ZN(n1157) );
NOR3_X1 U874 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(G51) );
AND3_X1 U875 ( .A1(KEYINPUT61), .A2(n1171), .A3(G952), .ZN(n1210) );
NOR2_X1 U876 ( .A1(KEYINPUT61), .A2(n1172), .ZN(n1209) );
NAND2_X1 U877 ( .A1(n1171), .A2(n1211), .ZN(n1172) );
INV_X1 U878 ( .A(G952), .ZN(n1211) );
XOR2_X1 U879 ( .A(G953), .B(KEYINPUT14), .Z(n1171) );
XOR2_X1 U880 ( .A(n1212), .B(n1213), .Z(n1208) );
XOR2_X1 U881 ( .A(n1214), .B(n1215), .Z(n1213) );
NAND2_X1 U882 ( .A1(KEYINPUT23), .A2(n1156), .ZN(n1215) );
NAND2_X1 U883 ( .A1(n1167), .A2(G210), .ZN(n1214) );
INV_X1 U884 ( .A(n1161), .ZN(n1167) );
NAND2_X1 U885 ( .A1(G902), .A2(n1065), .ZN(n1161) );
NAND4_X1 U886 ( .A1(n1152), .A2(n1119), .A3(n1154), .A4(n1121), .ZN(n1065) );
NAND2_X1 U887 ( .A1(n1078), .A2(n1216), .ZN(n1154) );
XNOR2_X1 U888 ( .A(KEYINPUT35), .B(n1180), .ZN(n1216) );
NAND4_X1 U889 ( .A1(n1097), .A2(n1099), .A3(n1090), .A4(n1217), .ZN(n1180) );
INV_X1 U890 ( .A(n1076), .ZN(n1099) );
AND4_X1 U891 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1119) );
AND4_X1 U892 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
NAND2_X1 U893 ( .A1(n1226), .A2(n1227), .ZN(n1220) );
XNOR2_X1 U894 ( .A(n1103), .B(KEYINPUT10), .ZN(n1226) );
AND4_X1 U895 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1152) );
NOR4_X1 U896 ( .A1(n1232), .A2(n1233), .A3(n1060), .A4(n1234), .ZN(n1231) );
INV_X1 U897 ( .A(n1235), .ZN(n1234) );
NOR3_X1 U898 ( .A1(n1076), .A2(n1098), .A3(n1236), .ZN(n1060) );
INV_X1 U899 ( .A(n1101), .ZN(n1098) );
NAND2_X1 U900 ( .A1(n1237), .A2(n1078), .ZN(n1230) );
XOR2_X1 U901 ( .A(n1238), .B(KEYINPUT16), .Z(n1237) );
NAND4_X1 U902 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1217), .ZN(n1229) );
INV_X1 U903 ( .A(n1242), .ZN(n1241) );
XNOR2_X1 U904 ( .A(n1090), .B(KEYINPUT49), .ZN(n1240) );
XNOR2_X1 U905 ( .A(n1078), .B(KEYINPUT54), .ZN(n1239) );
NAND3_X1 U906 ( .A1(n1243), .A2(n1244), .A3(n1084), .ZN(n1228) );
XNOR2_X1 U907 ( .A(G146), .B(n1223), .ZN(G48) );
NAND3_X1 U908 ( .A1(n1245), .A2(n1078), .A3(n1097), .ZN(n1223) );
XNOR2_X1 U909 ( .A(G143), .B(n1222), .ZN(G45) );
NAND4_X1 U910 ( .A1(n1246), .A2(n1247), .A3(n1078), .A4(n1248), .ZN(n1222) );
XNOR2_X1 U911 ( .A(G140), .B(n1218), .ZN(G42) );
NAND3_X1 U912 ( .A1(n1103), .A2(n1090), .A3(n1249), .ZN(n1218) );
XNOR2_X1 U913 ( .A(G137), .B(n1219), .ZN(G39) );
NAND3_X1 U914 ( .A1(n1103), .A2(n1244), .A3(n1245), .ZN(n1219) );
XNOR2_X1 U915 ( .A(G134), .B(n1250), .ZN(G36) );
NAND2_X1 U916 ( .A1(n1227), .A2(n1103), .ZN(n1250) );
AND2_X1 U917 ( .A1(n1247), .A2(n1101), .ZN(n1227) );
XNOR2_X1 U918 ( .A(G131), .B(n1225), .ZN(G33) );
NAND3_X1 U919 ( .A1(n1097), .A2(n1103), .A3(n1247), .ZN(n1225) );
AND3_X1 U920 ( .A1(n1090), .A2(n1251), .A3(n1084), .ZN(n1247) );
NOR2_X1 U921 ( .A1(n1079), .A2(n1252), .ZN(n1103) );
XNOR2_X1 U922 ( .A(G128), .B(n1121), .ZN(G30) );
NAND3_X1 U923 ( .A1(n1078), .A2(n1101), .A3(n1245), .ZN(n1121) );
AND4_X1 U924 ( .A1(n1253), .A2(n1090), .A3(n1254), .A4(n1251), .ZN(n1245) );
INV_X1 U925 ( .A(n1255), .ZN(n1090) );
XNOR2_X1 U926 ( .A(G101), .B(n1256), .ZN(G3) );
NAND3_X1 U927 ( .A1(n1243), .A2(n1257), .A3(n1084), .ZN(n1256) );
XNOR2_X1 U928 ( .A(KEYINPUT55), .B(n1072), .ZN(n1257) );
XNOR2_X1 U929 ( .A(G125), .B(n1224), .ZN(G27) );
NAND3_X1 U930 ( .A1(n1102), .A2(n1078), .A3(n1249), .ZN(n1224) );
AND3_X1 U931 ( .A1(n1097), .A2(n1251), .A3(n1083), .ZN(n1249) );
NAND2_X1 U932 ( .A1(n1067), .A2(n1258), .ZN(n1251) );
NAND4_X1 U933 ( .A1(G953), .A2(G902), .A3(n1259), .A4(n1124), .ZN(n1258) );
INV_X1 U934 ( .A(G900), .ZN(n1124) );
INV_X1 U935 ( .A(n1179), .ZN(n1078) );
XOR2_X1 U936 ( .A(G122), .B(n1260), .Z(G24) );
NOR3_X1 U937 ( .A1(KEYINPUT47), .A2(n1261), .A3(n1262), .ZN(n1260) );
NOR2_X1 U938 ( .A1(KEYINPUT19), .A2(n1263), .ZN(n1262) );
NOR2_X1 U939 ( .A1(n1179), .A2(n1238), .ZN(n1263) );
NAND3_X1 U940 ( .A1(n1246), .A2(n1102), .A3(n1264), .ZN(n1238) );
NOR3_X1 U941 ( .A1(n1076), .A2(n1265), .A3(n1266), .ZN(n1264) );
INV_X1 U942 ( .A(n1070), .ZN(n1102) );
NOR2_X1 U943 ( .A1(n1267), .A2(n1268), .ZN(n1261) );
INV_X1 U944 ( .A(KEYINPUT19), .ZN(n1268) );
NOR3_X1 U945 ( .A1(n1269), .A2(n1270), .A3(n1076), .ZN(n1267) );
NAND2_X1 U946 ( .A1(n1271), .A2(n1272), .ZN(n1076) );
NOR2_X1 U947 ( .A1(n1265), .A2(n1273), .ZN(n1270) );
INV_X1 U948 ( .A(n1248), .ZN(n1265) );
INV_X1 U949 ( .A(n1274), .ZN(n1269) );
XOR2_X1 U950 ( .A(G119), .B(n1233), .Z(G21) );
AND4_X1 U951 ( .A1(n1253), .A2(n1274), .A3(n1244), .A4(n1254), .ZN(n1233) );
XOR2_X1 U952 ( .A(n1275), .B(KEYINPUT28), .Z(n1253) );
NAND2_X1 U953 ( .A1(n1276), .A2(n1277), .ZN(G18) );
OR2_X1 U954 ( .A1(n1278), .A2(G116), .ZN(n1277) );
NAND2_X1 U955 ( .A1(G116), .A2(n1279), .ZN(n1276) );
NAND2_X1 U956 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NAND2_X1 U957 ( .A1(KEYINPUT29), .A2(n1232), .ZN(n1281) );
NAND2_X1 U958 ( .A1(n1278), .A2(n1282), .ZN(n1280) );
INV_X1 U959 ( .A(KEYINPUT29), .ZN(n1282) );
NAND2_X1 U960 ( .A1(KEYINPUT32), .A2(n1232), .ZN(n1278) );
AND3_X1 U961 ( .A1(n1274), .A2(n1101), .A3(n1084), .ZN(n1232) );
NAND2_X1 U962 ( .A1(n1283), .A2(n1284), .ZN(n1101) );
OR2_X1 U963 ( .A1(n1072), .A2(KEYINPUT8), .ZN(n1284) );
INV_X1 U964 ( .A(n1244), .ZN(n1072) );
NAND3_X1 U965 ( .A1(n1273), .A2(n1248), .A3(KEYINPUT8), .ZN(n1283) );
XNOR2_X1 U966 ( .A(G113), .B(n1235), .ZN(G15) );
NAND3_X1 U967 ( .A1(n1274), .A2(n1097), .A3(n1084), .ZN(n1235) );
AND2_X1 U968 ( .A1(n1272), .A2(n1254), .ZN(n1084) );
NOR2_X1 U969 ( .A1(n1273), .A2(n1248), .ZN(n1097) );
NOR3_X1 U970 ( .A1(n1179), .A2(n1266), .A3(n1070), .ZN(n1274) );
NAND2_X1 U971 ( .A1(n1285), .A2(n1093), .ZN(n1070) );
INV_X1 U972 ( .A(n1092), .ZN(n1285) );
XOR2_X1 U973 ( .A(n1286), .B(n1287), .Z(G12) );
NOR2_X1 U974 ( .A1(n1236), .A2(n1242), .ZN(n1287) );
NAND2_X1 U975 ( .A1(n1083), .A2(n1244), .ZN(n1242) );
NOR2_X1 U976 ( .A1(n1248), .A2(n1246), .ZN(n1244) );
INV_X1 U977 ( .A(n1273), .ZN(n1246) );
XNOR2_X1 U978 ( .A(n1109), .B(n1288), .ZN(n1273) );
NOR2_X1 U979 ( .A1(G475), .A2(KEYINPUT1), .ZN(n1288) );
NAND2_X1 U980 ( .A1(n1174), .A2(n1289), .ZN(n1109) );
XNOR2_X1 U981 ( .A(n1290), .B(n1291), .ZN(n1174) );
XNOR2_X1 U982 ( .A(n1292), .B(n1293), .ZN(n1291) );
NOR2_X1 U983 ( .A1(KEYINPUT26), .A2(n1294), .ZN(n1293) );
XNOR2_X1 U984 ( .A(n1137), .B(n1295), .ZN(n1294) );
NOR2_X1 U985 ( .A1(G146), .A2(KEYINPUT40), .ZN(n1295) );
XNOR2_X1 U986 ( .A(G125), .B(n1201), .ZN(n1137) );
XOR2_X1 U987 ( .A(n1296), .B(n1297), .Z(n1290) );
NAND3_X1 U988 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1296) );
NAND2_X1 U989 ( .A1(KEYINPUT51), .A2(G131), .ZN(n1300) );
OR3_X1 U990 ( .A1(G131), .A2(KEYINPUT51), .A3(n1301), .ZN(n1299) );
NAND2_X1 U991 ( .A1(n1302), .A2(n1301), .ZN(n1298) );
NAND2_X1 U992 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
NAND2_X1 U993 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U994 ( .A(n1307), .B(KEYINPUT24), .Z(n1303) );
OR2_X1 U995 ( .A1(n1305), .A2(n1306), .ZN(n1307) );
NAND3_X1 U996 ( .A1(n1308), .A2(n1117), .A3(G214), .ZN(n1305) );
NAND2_X1 U997 ( .A1(n1309), .A2(n1310), .ZN(n1302) );
INV_X1 U998 ( .A(KEYINPUT51), .ZN(n1310) );
XNOR2_X1 U999 ( .A(G131), .B(KEYINPUT45), .ZN(n1309) );
NAND2_X1 U1000 ( .A1(n1311), .A2(n1104), .ZN(n1248) );
NAND2_X1 U1001 ( .A1(n1111), .A2(n1110), .ZN(n1104) );
INV_X1 U1002 ( .A(G478), .ZN(n1110) );
INV_X1 U1003 ( .A(n1312), .ZN(n1111) );
NAND2_X1 U1004 ( .A1(G478), .A2(n1312), .ZN(n1311) );
NAND2_X1 U1005 ( .A1(n1165), .A2(n1289), .ZN(n1312) );
XNOR2_X1 U1006 ( .A(n1313), .B(n1314), .ZN(n1165) );
NOR2_X1 U1007 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
INV_X1 U1008 ( .A(G217), .ZN(n1315) );
NAND2_X1 U1009 ( .A1(n1317), .A2(KEYINPUT53), .ZN(n1313) );
XNOR2_X1 U1010 ( .A(n1318), .B(n1319), .ZN(n1317) );
XNOR2_X1 U1011 ( .A(n1135), .B(n1320), .ZN(n1319) );
NOR2_X1 U1012 ( .A1(KEYINPUT22), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1013 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1014 ( .A(KEYINPUT62), .B(G122), .Z(n1323) );
INV_X1 U1015 ( .A(G134), .ZN(n1135) );
AND2_X1 U1016 ( .A1(n1275), .A2(n1271), .ZN(n1083) );
INV_X1 U1017 ( .A(n1254), .ZN(n1271) );
XNOR2_X1 U1018 ( .A(n1324), .B(G472), .ZN(n1254) );
NAND2_X1 U1019 ( .A1(n1325), .A2(n1289), .ZN(n1324) );
XOR2_X1 U1020 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1021 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U1022 ( .A1(KEYINPUT11), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1023 ( .A(n1187), .B(KEYINPUT2), .ZN(n1330) );
NAND2_X1 U1024 ( .A1(KEYINPUT43), .A2(n1189), .ZN(n1328) );
AND3_X1 U1025 ( .A1(n1308), .A2(n1117), .A3(G210), .ZN(n1189) );
INV_X1 U1026 ( .A(G237), .ZN(n1308) );
XNOR2_X1 U1027 ( .A(n1331), .B(n1184), .ZN(n1326) );
XOR2_X1 U1028 ( .A(n1332), .B(G101), .Z(n1184) );
NAND2_X1 U1029 ( .A1(KEYINPUT39), .A2(n1185), .ZN(n1331) );
XNOR2_X1 U1030 ( .A(n1333), .B(n1334), .ZN(n1185) );
XOR2_X1 U1031 ( .A(G119), .B(G116), .Z(n1334) );
NAND2_X1 U1032 ( .A1(KEYINPUT31), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1033 ( .A(n1272), .B(KEYINPUT20), .Z(n1275) );
XNOR2_X1 U1034 ( .A(n1336), .B(n1162), .ZN(n1272) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1337), .ZN(n1162) );
OR2_X1 U1036 ( .A1(n1160), .A2(G902), .ZN(n1336) );
XNOR2_X1 U1037 ( .A(n1338), .B(n1339), .ZN(n1160) );
XOR2_X1 U1038 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1039 ( .A(n1342), .B(G137), .ZN(n1341) );
NOR2_X1 U1040 ( .A1(KEYINPUT48), .A2(G128), .ZN(n1340) );
XNOR2_X1 U1041 ( .A(n1343), .B(n1344), .ZN(n1338) );
XOR2_X1 U1042 ( .A(n1345), .B(n1346), .Z(n1344) );
NOR2_X1 U1043 ( .A1(n1347), .A2(n1316), .ZN(n1346) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1117), .ZN(n1316) );
INV_X1 U1045 ( .A(G221), .ZN(n1347) );
NOR2_X1 U1046 ( .A1(KEYINPUT12), .A2(n1348), .ZN(n1345) );
XOR2_X1 U1047 ( .A(n1349), .B(n1350), .Z(n1348) );
NOR2_X1 U1048 ( .A1(KEYINPUT21), .A2(n1351), .ZN(n1350) );
XNOR2_X1 U1049 ( .A(KEYINPUT58), .B(n1201), .ZN(n1351) );
XNOR2_X1 U1050 ( .A(G125), .B(KEYINPUT56), .ZN(n1349) );
INV_X1 U1051 ( .A(n1243), .ZN(n1236) );
NOR3_X1 U1052 ( .A1(n1179), .A2(n1266), .A3(n1255), .ZN(n1243) );
NAND2_X1 U1053 ( .A1(n1092), .A2(n1093), .ZN(n1255) );
NAND2_X1 U1054 ( .A1(G221), .A2(n1337), .ZN(n1093) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1289), .ZN(n1337) );
XNOR2_X1 U1056 ( .A(n1352), .B(G469), .ZN(n1092) );
NAND2_X1 U1057 ( .A1(n1353), .A2(n1289), .ZN(n1352) );
XOR2_X1 U1058 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1059 ( .A(n1204), .B(n1356), .ZN(n1355) );
XNOR2_X1 U1060 ( .A(KEYINPUT37), .B(n1201), .ZN(n1356) );
INV_X1 U1061 ( .A(G140), .ZN(n1201) );
XOR2_X1 U1062 ( .A(n1357), .B(n1187), .Z(n1354) );
XNOR2_X1 U1063 ( .A(n1358), .B(n1359), .ZN(n1187) );
XOR2_X1 U1064 ( .A(KEYINPUT44), .B(G137), .Z(n1359) );
XNOR2_X1 U1065 ( .A(G134), .B(G131), .ZN(n1358) );
XOR2_X1 U1066 ( .A(n1360), .B(n1203), .Z(n1357) );
AND2_X1 U1067 ( .A1(G227), .A2(n1117), .ZN(n1203) );
NAND2_X1 U1068 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
NAND2_X1 U1069 ( .A1(n1207), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1070 ( .A(n1364), .B(KEYINPUT46), .Z(n1361) );
OR2_X1 U1071 ( .A1(n1363), .A2(n1207), .ZN(n1364) );
AND2_X1 U1072 ( .A1(n1365), .A2(n1366), .ZN(n1207) );
NAND2_X1 U1073 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
INV_X1 U1074 ( .A(G101), .ZN(n1368) );
XNOR2_X1 U1075 ( .A(G107), .B(n1369), .ZN(n1367) );
NAND2_X1 U1076 ( .A1(n1370), .A2(G101), .ZN(n1365) );
XNOR2_X1 U1077 ( .A(n1059), .B(n1369), .ZN(n1370) );
NOR2_X1 U1078 ( .A1(KEYINPUT57), .A2(n1292), .ZN(n1369) );
INV_X1 U1079 ( .A(G104), .ZN(n1292) );
XNOR2_X1 U1080 ( .A(n1125), .B(KEYINPUT9), .ZN(n1363) );
XNOR2_X1 U1081 ( .A(G146), .B(n1318), .ZN(n1125) );
XNOR2_X1 U1082 ( .A(G128), .B(n1306), .ZN(n1318) );
INV_X1 U1083 ( .A(G143), .ZN(n1306) );
INV_X1 U1084 ( .A(n1217), .ZN(n1266) );
NAND2_X1 U1085 ( .A1(n1371), .A2(n1067), .ZN(n1217) );
NAND3_X1 U1086 ( .A1(n1259), .A2(n1117), .A3(G952), .ZN(n1067) );
XOR2_X1 U1087 ( .A(n1372), .B(KEYINPUT15), .Z(n1371) );
NAND4_X1 U1088 ( .A1(G953), .A2(G902), .A3(n1259), .A4(n1149), .ZN(n1372) );
INV_X1 U1089 ( .A(G898), .ZN(n1149) );
NAND2_X1 U1090 ( .A1(G237), .A2(G234), .ZN(n1259) );
NAND2_X1 U1091 ( .A1(n1079), .A2(n1080), .ZN(n1179) );
INV_X1 U1092 ( .A(n1252), .ZN(n1080) );
NOR2_X1 U1093 ( .A1(n1373), .A2(n1374), .ZN(n1252) );
INV_X1 U1094 ( .A(G214), .ZN(n1373) );
XNOR2_X1 U1095 ( .A(n1375), .B(n1376), .ZN(n1079) );
NOR2_X1 U1096 ( .A1(n1374), .A2(n1377), .ZN(n1376) );
XOR2_X1 U1097 ( .A(KEYINPUT5), .B(G210), .Z(n1377) );
NOR2_X1 U1098 ( .A1(G902), .A2(G237), .ZN(n1374) );
NAND2_X1 U1099 ( .A1(n1378), .A2(n1289), .ZN(n1375) );
INV_X1 U1100 ( .A(G902), .ZN(n1289) );
XNOR2_X1 U1101 ( .A(n1212), .B(n1156), .ZN(n1378) );
XNOR2_X1 U1102 ( .A(n1379), .B(n1380), .ZN(n1156) );
XOR2_X1 U1103 ( .A(n1297), .B(n1343), .Z(n1380) );
XNOR2_X1 U1104 ( .A(G119), .B(n1204), .ZN(n1343) );
XNOR2_X1 U1105 ( .A(n1335), .B(G122), .ZN(n1297) );
INV_X1 U1106 ( .A(G113), .ZN(n1335) );
XOR2_X1 U1107 ( .A(n1381), .B(n1322), .Z(n1379) );
XNOR2_X1 U1108 ( .A(n1059), .B(G116), .ZN(n1322) );
INV_X1 U1109 ( .A(G107), .ZN(n1059) );
XNOR2_X1 U1110 ( .A(G101), .B(G104), .ZN(n1381) );
XNOR2_X1 U1111 ( .A(n1332), .B(n1382), .ZN(n1212) );
XNOR2_X1 U1112 ( .A(n1383), .B(n1384), .ZN(n1382) );
AND2_X1 U1113 ( .A1(n1117), .A2(G224), .ZN(n1384) );
INV_X1 U1114 ( .A(G953), .ZN(n1117) );
INV_X1 U1115 ( .A(G125), .ZN(n1383) );
XOR2_X1 U1116 ( .A(n1385), .B(G128), .Z(n1332) );
NAND2_X1 U1117 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
NAND2_X1 U1118 ( .A1(G143), .A2(n1342), .ZN(n1387) );
XOR2_X1 U1119 ( .A(KEYINPUT63), .B(n1388), .Z(n1386) );
NOR2_X1 U1120 ( .A1(G143), .A2(n1342), .ZN(n1388) );
INV_X1 U1121 ( .A(G146), .ZN(n1342) );
NOR2_X1 U1122 ( .A1(KEYINPUT41), .A2(n1204), .ZN(n1286) );
INV_X1 U1123 ( .A(G110), .ZN(n1204) );
endmodule


