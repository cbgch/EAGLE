//Key = 0000001101011100011110001110111100100001011011110100101110101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317;

XOR2_X1 U721 ( .A(G107), .B(n1003), .Z(G9) );
NOR2_X1 U722 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR4_X1 U723 ( .A1(G953), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1005) );
NOR3_X1 U724 ( .A1(n1009), .A2(KEYINPUT36), .A3(n1010), .ZN(n1007) );
NOR2_X1 U725 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR2_X1 U726 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U727 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U728 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR2_X1 U729 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U730 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U731 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U732 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U733 ( .A1(n1027), .A2(n1028), .ZN(n1019) );
NOR2_X1 U734 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR3_X1 U735 ( .A1(n1028), .A2(n1031), .A3(n1022), .ZN(n1015) );
NOR3_X1 U736 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
AND3_X1 U737 ( .A1(KEYINPUT20), .A2(n1035), .A3(n1036), .ZN(n1034) );
NOR2_X1 U738 ( .A1(KEYINPUT20), .A2(n1018), .ZN(n1033) );
NOR4_X1 U739 ( .A1(n1037), .A2(n1022), .A3(n1028), .A4(n1018), .ZN(n1011) );
NOR2_X1 U740 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR3_X1 U741 ( .A1(n1006), .A2(G953), .A3(G952), .ZN(n1004) );
AND4_X1 U742 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1006) );
NOR4_X1 U743 ( .A1(n1044), .A2(n1045), .A3(n1036), .A4(n1046), .ZN(n1043) );
NOR2_X1 U744 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
INV_X1 U745 ( .A(n1049), .ZN(n1044) );
NOR2_X1 U746 ( .A1(n1050), .A2(n1051), .ZN(n1042) );
XOR2_X1 U747 ( .A(n1052), .B(n1053), .Z(n1051) );
XOR2_X1 U748 ( .A(n1054), .B(n1055), .Z(n1050) );
NAND2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
INV_X1 U750 ( .A(n1058), .ZN(n1056) );
XOR2_X1 U751 ( .A(n1059), .B(n1060), .Z(G72) );
XOR2_X1 U752 ( .A(n1061), .B(n1062), .Z(n1060) );
NAND2_X1 U753 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U754 ( .A1(G953), .A2(n1065), .ZN(n1064) );
XOR2_X1 U755 ( .A(n1066), .B(n1067), .Z(n1063) );
XOR2_X1 U756 ( .A(G140), .B(G131), .Z(n1067) );
XOR2_X1 U757 ( .A(n1068), .B(n1069), .Z(n1066) );
NAND2_X1 U758 ( .A1(G953), .A2(n1070), .ZN(n1061) );
NAND2_X1 U759 ( .A1(n1071), .A2(G227), .ZN(n1070) );
XOR2_X1 U760 ( .A(n1065), .B(KEYINPUT42), .Z(n1071) );
NOR2_X1 U761 ( .A1(n1072), .A2(G953), .ZN(n1059) );
XOR2_X1 U762 ( .A(n1073), .B(n1074), .Z(G69) );
NOR2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
AND4_X1 U764 ( .A1(KEYINPUT10), .A2(G898), .A3(G953), .A4(G224), .ZN(n1076) );
NOR2_X1 U765 ( .A1(KEYINPUT10), .A2(n1077), .ZN(n1075) );
NOR2_X1 U766 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U767 ( .A1(G224), .A2(n1080), .ZN(n1078) );
XOR2_X1 U768 ( .A(n1081), .B(n1082), .Z(n1073) );
NOR2_X1 U769 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U770 ( .A(n1080), .B(KEYINPUT30), .Z(n1084) );
NAND2_X1 U771 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
XOR2_X1 U772 ( .A(n1087), .B(n1088), .Z(n1085) );
XOR2_X1 U773 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U774 ( .A1(KEYINPUT50), .A2(n1091), .ZN(n1089) );
NOR2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(G66) );
XNOR2_X1 U776 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U777 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U778 ( .A(KEYINPUT11), .B(G217), .Z(n1097) );
NOR2_X1 U779 ( .A1(n1092), .A2(n1098), .ZN(G63) );
XOR2_X1 U780 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U781 ( .A1(n1048), .A2(n1096), .ZN(n1100) );
NOR2_X1 U782 ( .A1(n1092), .A2(n1101), .ZN(G60) );
XOR2_X1 U783 ( .A(n1058), .B(n1102), .Z(n1101) );
NOR2_X1 U784 ( .A1(n1054), .A2(n1096), .ZN(n1102) );
XOR2_X1 U785 ( .A(n1103), .B(n1104), .Z(G6) );
NAND2_X1 U786 ( .A1(n1105), .A2(n1032), .ZN(n1104) );
XOR2_X1 U787 ( .A(n1106), .B(KEYINPUT25), .Z(n1105) );
NAND4_X1 U788 ( .A1(n1041), .A2(n1024), .A3(n1107), .A4(n1108), .ZN(n1106) );
XOR2_X1 U789 ( .A(KEYINPUT2), .B(n1030), .Z(n1107) );
INV_X1 U790 ( .A(n1109), .ZN(n1024) );
NOR2_X1 U791 ( .A1(n1092), .A2(n1110), .ZN(G57) );
XOR2_X1 U792 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U793 ( .A(KEYINPUT33), .B(n1113), .Z(n1112) );
NOR2_X1 U794 ( .A1(n1114), .A2(n1096), .ZN(n1113) );
INV_X1 U795 ( .A(G472), .ZN(n1114) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1111) );
NAND2_X1 U797 ( .A1(KEYINPUT62), .A2(n1117), .ZN(n1115) );
INV_X1 U798 ( .A(n1118), .ZN(n1117) );
NOR2_X1 U799 ( .A1(n1092), .A2(n1119), .ZN(G54) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U801 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U802 ( .A(n1124), .B(n1125), .Z(n1120) );
NOR3_X1 U803 ( .A1(n1052), .A2(n1126), .A3(n1057), .ZN(n1125) );
XOR2_X1 U804 ( .A(n1008), .B(KEYINPUT6), .Z(n1126) );
NAND2_X1 U805 ( .A1(KEYINPUT58), .A2(n1127), .ZN(n1124) );
XOR2_X1 U806 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U807 ( .A1(KEYINPUT59), .A2(n1130), .ZN(n1128) );
NOR2_X1 U808 ( .A1(n1092), .A2(n1131), .ZN(G51) );
XOR2_X1 U809 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U810 ( .A1(n1134), .A2(KEYINPUT8), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1135), .A2(n1096), .ZN(n1134) );
NAND2_X1 U812 ( .A1(G902), .A2(n1008), .ZN(n1096) );
NAND2_X1 U813 ( .A1(n1083), .A2(n1072), .ZN(n1008) );
AND4_X1 U814 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1072) );
AND4_X1 U815 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1145), .ZN(n1138) );
NAND2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U818 ( .A(KEYINPUT34), .B(n1029), .Z(n1146) );
NAND2_X1 U819 ( .A1(n1148), .A2(n1149), .ZN(n1137) );
NAND3_X1 U820 ( .A1(n1038), .A2(n1029), .A3(n1150), .ZN(n1136) );
AND4_X1 U821 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1083) );
NOR4_X1 U822 ( .A1(n1155), .A2(n1156), .A3(n1003), .A4(n1157), .ZN(n1154) );
NOR3_X1 U823 ( .A1(n1158), .A2(n1159), .A3(n1014), .ZN(n1003) );
NOR2_X1 U824 ( .A1(n1160), .A2(n1161), .ZN(n1153) );
NOR2_X1 U825 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NOR3_X1 U826 ( .A1(n1147), .A2(n1158), .A3(n1014), .ZN(n1160) );
NOR3_X1 U827 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1132) );
NOR2_X1 U828 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
AND2_X1 U829 ( .A1(n1169), .A2(KEYINPUT12), .ZN(n1167) );
AND4_X1 U830 ( .A1(n1168), .A2(KEYINPUT31), .A3(n1169), .A4(KEYINPUT12), .ZN(n1165) );
NOR2_X1 U831 ( .A1(KEYINPUT31), .A2(n1169), .ZN(n1164) );
XNOR2_X1 U832 ( .A(n1170), .B(n1069), .ZN(n1169) );
XOR2_X1 U833 ( .A(G125), .B(n1171), .Z(n1069) );
NOR2_X1 U834 ( .A1(n1080), .A2(G952), .ZN(n1092) );
XOR2_X1 U835 ( .A(n1172), .B(n1173), .Z(G48) );
NAND3_X1 U836 ( .A1(n1144), .A2(n1030), .A3(KEYINPUT39), .ZN(n1173) );
INV_X1 U837 ( .A(n1174), .ZN(n1144) );
NAND2_X1 U838 ( .A1(n1175), .A2(n1176), .ZN(G45) );
NAND2_X1 U839 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
INV_X1 U840 ( .A(G143), .ZN(n1178) );
NAND2_X1 U841 ( .A1(G143), .A2(n1179), .ZN(n1175) );
NAND2_X1 U842 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND2_X1 U843 ( .A1(KEYINPUT27), .A2(n1182), .ZN(n1181) );
INV_X1 U844 ( .A(n1143), .ZN(n1182) );
OR2_X1 U845 ( .A1(n1177), .A2(KEYINPUT27), .ZN(n1180) );
NOR2_X1 U846 ( .A1(KEYINPUT21), .A2(n1143), .ZN(n1177) );
NAND4_X1 U847 ( .A1(n1183), .A2(n1038), .A3(n1184), .A4(n1185), .ZN(n1143) );
NOR2_X1 U848 ( .A1(n1186), .A2(n1187), .ZN(n1184) );
XOR2_X1 U849 ( .A(n1188), .B(n1142), .Z(G42) );
NAND3_X1 U850 ( .A1(n1030), .A2(n1039), .A3(n1150), .ZN(n1142) );
XOR2_X1 U851 ( .A(n1189), .B(n1141), .Z(G39) );
NAND4_X1 U852 ( .A1(n1150), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1141) );
XOR2_X1 U853 ( .A(n1193), .B(n1194), .Z(G36) );
NAND3_X1 U854 ( .A1(n1195), .A2(n1183), .A3(n1196), .ZN(n1194) );
NOR3_X1 U855 ( .A1(n1018), .A2(n1159), .A3(n1197), .ZN(n1196) );
XOR2_X1 U856 ( .A(n1109), .B(KEYINPUT41), .Z(n1195) );
XNOR2_X1 U857 ( .A(G131), .B(n1198), .ZN(G33) );
NAND2_X1 U858 ( .A1(KEYINPUT55), .A2(n1199), .ZN(n1198) );
INV_X1 U859 ( .A(n1140), .ZN(n1199) );
NAND3_X1 U860 ( .A1(n1030), .A2(n1038), .A3(n1150), .ZN(n1140) );
NOR3_X1 U861 ( .A1(n1018), .A2(n1109), .A3(n1200), .ZN(n1150) );
NAND2_X1 U862 ( .A1(n1035), .A2(n1201), .ZN(n1018) );
XNOR2_X1 U863 ( .A(n1040), .B(KEYINPUT54), .ZN(n1035) );
XOR2_X1 U864 ( .A(n1202), .B(n1203), .Z(G30) );
NOR2_X1 U865 ( .A1(KEYINPUT35), .A2(n1204), .ZN(n1203) );
NOR2_X1 U866 ( .A1(n1159), .A2(n1174), .ZN(n1202) );
NAND4_X1 U867 ( .A1(n1183), .A2(n1185), .A3(n1191), .A4(n1192), .ZN(n1174) );
INV_X1 U868 ( .A(n1200), .ZN(n1183) );
XNOR2_X1 U869 ( .A(G101), .B(n1205), .ZN(G3) );
NAND2_X1 U870 ( .A1(KEYINPUT46), .A2(n1156), .ZN(n1205) );
NOR3_X1 U871 ( .A1(n1022), .A2(n1158), .A3(n1197), .ZN(n1156) );
INV_X1 U872 ( .A(n1038), .ZN(n1197) );
XOR2_X1 U873 ( .A(n1206), .B(n1207), .Z(G27) );
NAND2_X1 U874 ( .A1(n1208), .A2(n1148), .ZN(n1207) );
NOR4_X1 U875 ( .A1(n1200), .A2(n1147), .A3(n1162), .A4(n1209), .ZN(n1148) );
INV_X1 U876 ( .A(n1030), .ZN(n1147) );
NAND3_X1 U877 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1200) );
OR2_X1 U878 ( .A1(G952), .A2(G953), .ZN(n1211) );
NAND2_X1 U879 ( .A1(G953), .A2(n1213), .ZN(n1210) );
NAND2_X1 U880 ( .A1(G902), .A2(n1065), .ZN(n1213) );
INV_X1 U881 ( .A(G900), .ZN(n1065) );
XOR2_X1 U882 ( .A(n1028), .B(KEYINPUT60), .Z(n1208) );
XOR2_X1 U883 ( .A(n1214), .B(G122), .Z(G24) );
NAND2_X1 U884 ( .A1(KEYINPUT18), .A2(n1215), .ZN(n1214) );
NAND2_X1 U885 ( .A1(n1032), .A2(n1216), .ZN(n1215) );
XNOR2_X1 U886 ( .A(KEYINPUT51), .B(n1163), .ZN(n1216) );
NAND4_X1 U887 ( .A1(n1217), .A2(n1108), .A3(n1218), .A4(n1219), .ZN(n1163) );
NOR2_X1 U888 ( .A1(n1014), .A2(n1028), .ZN(n1219) );
INV_X1 U889 ( .A(n1149), .ZN(n1028) );
INV_X1 U890 ( .A(n1187), .ZN(n1218) );
XOR2_X1 U891 ( .A(n1151), .B(n1220), .Z(G21) );
XNOR2_X1 U892 ( .A(G119), .B(KEYINPUT57), .ZN(n1220) );
NAND4_X1 U893 ( .A1(n1221), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1151) );
INV_X1 U894 ( .A(n1022), .ZN(n1190) );
XNOR2_X1 U895 ( .A(G116), .B(n1152), .ZN(G18) );
NAND3_X1 U896 ( .A1(n1038), .A2(n1029), .A3(n1221), .ZN(n1152) );
INV_X1 U897 ( .A(n1159), .ZN(n1029) );
NAND2_X1 U898 ( .A1(n1187), .A2(n1217), .ZN(n1159) );
INV_X1 U899 ( .A(n1186), .ZN(n1217) );
XOR2_X1 U900 ( .A(n1222), .B(KEYINPUT26), .Z(n1186) );
XOR2_X1 U901 ( .A(G113), .B(n1157), .Z(G15) );
AND3_X1 U902 ( .A1(n1221), .A2(n1038), .A3(n1030), .ZN(n1157) );
NOR2_X1 U903 ( .A1(n1222), .A2(n1187), .ZN(n1030) );
NOR2_X1 U904 ( .A1(n1192), .A2(n1223), .ZN(n1038) );
AND3_X1 U905 ( .A1(n1032), .A2(n1108), .A3(n1149), .ZN(n1221) );
NOR2_X1 U906 ( .A1(n1025), .A2(n1045), .ZN(n1149) );
INV_X1 U907 ( .A(n1026), .ZN(n1045) );
XOR2_X1 U908 ( .A(G110), .B(n1155), .Z(G12) );
NOR3_X1 U909 ( .A1(n1158), .A2(n1209), .A3(n1022), .ZN(n1155) );
NAND2_X1 U910 ( .A1(n1224), .A2(n1187), .ZN(n1022) );
XOR2_X1 U911 ( .A(n1225), .B(n1226), .Z(n1187) );
NOR3_X1 U912 ( .A1(n1058), .A2(KEYINPUT16), .A3(G902), .ZN(n1226) );
XOR2_X1 U913 ( .A(n1227), .B(n1228), .Z(n1058) );
XOR2_X1 U914 ( .A(G104), .B(n1229), .Z(n1228) );
NOR2_X1 U915 ( .A1(KEYINPUT4), .A2(n1230), .ZN(n1229) );
XOR2_X1 U916 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U917 ( .A(n1233), .B(n1234), .Z(n1232) );
XNOR2_X1 U918 ( .A(G131), .B(n1235), .ZN(n1234) );
NOR2_X1 U919 ( .A1(KEYINPUT23), .A2(G125), .ZN(n1235) );
NAND2_X1 U920 ( .A1(n1236), .A2(KEYINPUT47), .ZN(n1233) );
XOR2_X1 U921 ( .A(n1237), .B(G143), .Z(n1236) );
NAND2_X1 U922 ( .A1(G214), .A2(n1238), .ZN(n1237) );
XOR2_X1 U923 ( .A(n1188), .B(n1239), .Z(n1231) );
XOR2_X1 U924 ( .A(KEYINPUT37), .B(G146), .Z(n1239) );
XNOR2_X1 U925 ( .A(G113), .B(G122), .ZN(n1227) );
XOR2_X1 U926 ( .A(n1054), .B(KEYINPUT38), .Z(n1225) );
INV_X1 U927 ( .A(G475), .ZN(n1054) );
XOR2_X1 U928 ( .A(n1222), .B(KEYINPUT45), .Z(n1224) );
NAND3_X1 U929 ( .A1(n1240), .A2(n1241), .A3(n1049), .ZN(n1222) );
NAND2_X1 U930 ( .A1(n1047), .A2(n1048), .ZN(n1049) );
OR3_X1 U931 ( .A1(n1048), .A2(n1047), .A3(KEYINPUT14), .ZN(n1241) );
INV_X1 U932 ( .A(G478), .ZN(n1048) );
NAND2_X1 U933 ( .A1(KEYINPUT14), .A2(n1047), .ZN(n1240) );
NOR2_X1 U934 ( .A1(n1099), .A2(G902), .ZN(n1047) );
XOR2_X1 U935 ( .A(n1242), .B(n1243), .Z(n1099) );
XNOR2_X1 U936 ( .A(n1244), .B(n1245), .ZN(n1243) );
NAND2_X1 U937 ( .A1(KEYINPUT28), .A2(n1246), .ZN(n1244) );
XOR2_X1 U938 ( .A(G122), .B(G116), .Z(n1246) );
XOR2_X1 U939 ( .A(n1247), .B(n1248), .Z(n1242) );
XOR2_X1 U940 ( .A(G134), .B(G107), .Z(n1248) );
NAND3_X1 U941 ( .A1(n1249), .A2(G217), .A3(KEYINPUT49), .ZN(n1247) );
INV_X1 U942 ( .A(n1039), .ZN(n1209) );
NAND2_X1 U943 ( .A1(n1250), .A2(n1251), .ZN(n1039) );
OR2_X1 U944 ( .A1(n1014), .A2(KEYINPUT29), .ZN(n1251) );
INV_X1 U945 ( .A(n1041), .ZN(n1014) );
NOR2_X1 U946 ( .A1(n1192), .A2(n1191), .ZN(n1041) );
INV_X1 U947 ( .A(n1223), .ZN(n1191) );
NAND3_X1 U948 ( .A1(n1223), .A2(n1192), .A3(KEYINPUT29), .ZN(n1250) );
NAND3_X1 U949 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1192) );
OR2_X1 U950 ( .A1(n1255), .A2(n1094), .ZN(n1254) );
NAND3_X1 U951 ( .A1(n1094), .A2(n1255), .A3(n1057), .ZN(n1253) );
NAND2_X1 U952 ( .A1(G217), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U953 ( .A(n1257), .B(n1258), .ZN(n1094) );
XOR2_X1 U954 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U955 ( .A(G125), .B(G119), .Z(n1260) );
XOR2_X1 U956 ( .A(KEYINPUT48), .B(G128), .Z(n1259) );
XOR2_X1 U957 ( .A(n1261), .B(n1262), .Z(n1257) );
XOR2_X1 U958 ( .A(n1263), .B(n1264), .Z(n1262) );
NAND2_X1 U959 ( .A1(KEYINPUT13), .A2(n1189), .ZN(n1264) );
INV_X1 U960 ( .A(G137), .ZN(n1189) );
NAND2_X1 U961 ( .A1(KEYINPUT9), .A2(n1172), .ZN(n1263) );
XOR2_X1 U962 ( .A(n1265), .B(n1266), .Z(n1261) );
AND2_X1 U963 ( .A1(n1249), .A2(G221), .ZN(n1266) );
NOR2_X1 U964 ( .A1(n1256), .A2(G953), .ZN(n1249) );
INV_X1 U965 ( .A(G234), .ZN(n1256) );
NAND2_X1 U966 ( .A1(G902), .A2(G217), .ZN(n1252) );
XOR2_X1 U967 ( .A(n1267), .B(G472), .Z(n1223) );
NAND2_X1 U968 ( .A1(n1268), .A2(n1057), .ZN(n1267) );
XNOR2_X1 U969 ( .A(n1116), .B(n1269), .ZN(n1268) );
XNOR2_X1 U970 ( .A(KEYINPUT15), .B(n1270), .ZN(n1269) );
NOR2_X1 U971 ( .A1(KEYINPUT22), .A2(n1118), .ZN(n1270) );
XOR2_X1 U972 ( .A(n1122), .B(KEYINPUT56), .Z(n1118) );
XOR2_X1 U973 ( .A(n1271), .B(n1272), .Z(n1122) );
XNOR2_X1 U974 ( .A(n1273), .B(n1090), .ZN(n1116) );
XOR2_X1 U975 ( .A(n1274), .B(n1275), .Z(n1273) );
NAND2_X1 U976 ( .A1(G210), .A2(n1238), .ZN(n1274) );
NOR2_X1 U977 ( .A1(G953), .A2(G237), .ZN(n1238) );
NAND2_X1 U978 ( .A1(n1185), .A2(n1108), .ZN(n1158) );
NAND2_X1 U979 ( .A1(n1276), .A2(n1277), .ZN(n1108) );
NAND3_X1 U980 ( .A1(n1212), .A2(n1080), .A3(G952), .ZN(n1277) );
XOR2_X1 U981 ( .A(KEYINPUT19), .B(n1278), .Z(n1276) );
NOR3_X1 U982 ( .A1(n1086), .A2(n1010), .A3(n1057), .ZN(n1278) );
INV_X1 U983 ( .A(n1212), .ZN(n1010) );
NAND2_X1 U984 ( .A1(G237), .A2(G234), .ZN(n1212) );
INV_X1 U985 ( .A(n1079), .ZN(n1086) );
NOR2_X1 U986 ( .A1(n1080), .A2(G898), .ZN(n1079) );
NOR2_X1 U987 ( .A1(n1162), .A2(n1109), .ZN(n1185) );
NAND2_X1 U988 ( .A1(n1025), .A2(n1026), .ZN(n1109) );
NAND2_X1 U989 ( .A1(G221), .A2(n1279), .ZN(n1026) );
NAND2_X1 U990 ( .A1(G234), .A2(n1057), .ZN(n1279) );
XOR2_X1 U991 ( .A(n1052), .B(n1280), .Z(n1025) );
NOR2_X1 U992 ( .A1(KEYINPUT61), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U993 ( .A(KEYINPUT32), .B(n1053), .ZN(n1281) );
NAND2_X1 U994 ( .A1(n1282), .A2(n1057), .ZN(n1053) );
XOR2_X1 U995 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U996 ( .A(n1129), .B(n1272), .Z(n1284) );
XOR2_X1 U997 ( .A(G131), .B(n1285), .Z(n1272) );
NOR2_X1 U998 ( .A1(KEYINPUT63), .A2(n1068), .ZN(n1285) );
XOR2_X1 U999 ( .A(n1193), .B(G137), .Z(n1068) );
INV_X1 U1000 ( .A(G134), .ZN(n1193) );
INV_X1 U1001 ( .A(n1265), .ZN(n1129) );
XOR2_X1 U1002 ( .A(n1188), .B(n1286), .Z(n1265) );
INV_X1 U1003 ( .A(G140), .ZN(n1188) );
XNOR2_X1 U1004 ( .A(n1287), .B(n1130), .ZN(n1283) );
NAND2_X1 U1005 ( .A1(G227), .A2(n1080), .ZN(n1130) );
XOR2_X1 U1006 ( .A(n1288), .B(KEYINPUT7), .Z(n1287) );
NAND3_X1 U1007 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1288) );
OR2_X1 U1008 ( .A1(n1123), .A2(n1271), .ZN(n1291) );
NAND2_X1 U1009 ( .A1(KEYINPUT3), .A2(n1292), .ZN(n1290) );
NAND2_X1 U1010 ( .A1(n1293), .A2(n1123), .ZN(n1292) );
XOR2_X1 U1011 ( .A(n1294), .B(n1171), .Z(n1293) );
NAND2_X1 U1012 ( .A1(n1295), .A2(n1296), .ZN(n1289) );
INV_X1 U1013 ( .A(KEYINPUT3), .ZN(n1296) );
NAND2_X1 U1014 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
NAND3_X1 U1015 ( .A1(n1123), .A2(n1271), .A3(n1294), .ZN(n1298) );
INV_X1 U1016 ( .A(KEYINPUT0), .ZN(n1294) );
XNOR2_X1 U1017 ( .A(n1299), .B(n1275), .ZN(n1123) );
NAND2_X1 U1018 ( .A1(KEYINPUT0), .A2(n1171), .ZN(n1297) );
INV_X1 U1019 ( .A(G469), .ZN(n1052) );
INV_X1 U1020 ( .A(n1032), .ZN(n1162) );
NOR2_X1 U1021 ( .A1(n1040), .A2(n1036), .ZN(n1032) );
INV_X1 U1022 ( .A(n1201), .ZN(n1036) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1300), .ZN(n1201) );
XNOR2_X1 U1024 ( .A(n1301), .B(n1135), .ZN(n1040) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1300), .ZN(n1135) );
NAND2_X1 U1026 ( .A1(n1302), .A2(n1057), .ZN(n1300) );
INV_X1 U1027 ( .A(G237), .ZN(n1302) );
NAND2_X1 U1028 ( .A1(n1303), .A2(n1057), .ZN(n1301) );
INV_X1 U1029 ( .A(G902), .ZN(n1057) );
XNOR2_X1 U1030 ( .A(n1304), .B(n1168), .ZN(n1303) );
XNOR2_X1 U1031 ( .A(n1090), .B(n1305), .ZN(n1168) );
XOR2_X1 U1032 ( .A(n1091), .B(n1306), .Z(n1305) );
NAND2_X1 U1033 ( .A1(KEYINPUT24), .A2(n1087), .ZN(n1306) );
XNOR2_X1 U1034 ( .A(G122), .B(n1286), .ZN(n1087) );
XOR2_X1 U1035 ( .A(G110), .B(KEYINPUT5), .Z(n1286) );
NAND2_X1 U1036 ( .A1(n1307), .A2(n1308), .ZN(n1091) );
NAND2_X1 U1037 ( .A1(n1299), .A2(n1275), .ZN(n1308) );
XOR2_X1 U1038 ( .A(n1309), .B(KEYINPUT53), .Z(n1307) );
NAND2_X1 U1039 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
INV_X1 U1040 ( .A(n1299), .ZN(n1311) );
XOR2_X1 U1041 ( .A(n1103), .B(G107), .Z(n1299) );
INV_X1 U1042 ( .A(G104), .ZN(n1103) );
XNOR2_X1 U1043 ( .A(n1275), .B(KEYINPUT1), .ZN(n1310) );
XOR2_X1 U1044 ( .A(G101), .B(KEYINPUT52), .Z(n1275) );
XOR2_X1 U1045 ( .A(G113), .B(n1312), .Z(n1090) );
XOR2_X1 U1046 ( .A(G119), .B(G116), .Z(n1312) );
NOR2_X1 U1047 ( .A1(KEYINPUT40), .A2(n1313), .ZN(n1304) );
XOR2_X1 U1048 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1049 ( .A(n1206), .B(n1316), .Z(n1315) );
NOR2_X1 U1050 ( .A1(KEYINPUT43), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1051 ( .A(KEYINPUT44), .B(n1170), .ZN(n1317) );
NAND2_X1 U1052 ( .A1(G224), .A2(n1080), .ZN(n1170) );
INV_X1 U1053 ( .A(G953), .ZN(n1080) );
INV_X1 U1054 ( .A(G125), .ZN(n1206) );
NAND2_X1 U1055 ( .A1(KEYINPUT17), .A2(n1171), .ZN(n1314) );
INV_X1 U1056 ( .A(n1271), .ZN(n1171) );
XOR2_X1 U1057 ( .A(n1172), .B(n1245), .Z(n1271) );
XNOR2_X1 U1058 ( .A(n1204), .B(G143), .ZN(n1245) );
INV_X1 U1059 ( .A(G128), .ZN(n1204) );
INV_X1 U1060 ( .A(G146), .ZN(n1172) );
endmodule


