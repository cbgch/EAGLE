//Key = 0010000011011011001001111100101010000111001100110001101100101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348;

XOR2_X1 U744 ( .A(n1022), .B(n1023), .Z(G9) );
NAND2_X1 U745 ( .A1(KEYINPUT23), .A2(n1024), .ZN(n1023) );
INV_X1 U746 ( .A(n1025), .ZN(n1024) );
NOR2_X1 U747 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR4_X1 U748 ( .A1(G953), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1027) );
NOR2_X1 U749 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U750 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U751 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U752 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U753 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U754 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U755 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1041) );
NOR2_X1 U759 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR3_X1 U761 ( .A1(n1050), .A2(n1055), .A3(n1044), .ZN(n1037) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR4_X1 U764 ( .A1(n1060), .A2(n1044), .A3(n1040), .A4(n1050), .ZN(n1033) );
INV_X1 U765 ( .A(n1061), .ZN(n1050) );
NOR3_X1 U766 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n1026) );
AND4_X1 U767 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1028) );
NOR4_X1 U768 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1065) );
XOR2_X1 U769 ( .A(n1070), .B(KEYINPUT25), .Z(n1069) );
XNOR2_X1 U770 ( .A(n1071), .B(n1072), .ZN(n1068) );
NAND2_X1 U771 ( .A1(KEYINPUT54), .A2(n1073), .ZN(n1071) );
XOR2_X1 U772 ( .A(n1074), .B(n1075), .Z(n1067) );
NAND2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U774 ( .A1(KEYINPUT51), .A2(n1078), .ZN(n1077) );
NAND2_X1 U775 ( .A1(KEYINPUT45), .A2(n1079), .ZN(n1076) );
XOR2_X1 U776 ( .A(n1080), .B(G472), .Z(n1064) );
XOR2_X1 U777 ( .A(n1081), .B(n1082), .Z(G72) );
NOR2_X1 U778 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U779 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND2_X1 U780 ( .A1(n1087), .A2(n1088), .ZN(n1081) );
NAND2_X1 U781 ( .A1(n1089), .A2(n1084), .ZN(n1088) );
XNOR2_X1 U782 ( .A(n1090), .B(n1091), .ZN(n1089) );
NOR3_X1 U783 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
XNOR2_X1 U784 ( .A(KEYINPUT4), .B(n1095), .ZN(n1092) );
NAND3_X1 U785 ( .A1(n1090), .A2(G900), .A3(G953), .ZN(n1087) );
NOR2_X1 U786 ( .A1(KEYINPUT13), .A2(n1096), .ZN(n1090) );
XOR2_X1 U787 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U788 ( .A1(n1099), .A2(KEYINPUT22), .ZN(n1098) );
XOR2_X1 U789 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U790 ( .A(n1102), .B(G131), .Z(n1100) );
NAND2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U792 ( .A(KEYINPUT47), .B(KEYINPUT37), .ZN(n1103) );
XOR2_X1 U793 ( .A(n1105), .B(n1106), .Z(G69) );
XOR2_X1 U794 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U795 ( .A1(n1109), .A2(G953), .ZN(n1108) );
NOR2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
XOR2_X1 U797 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U798 ( .A(G122), .B(G110), .Z(n1113) );
NAND2_X1 U799 ( .A1(n1114), .A2(KEYINPUT24), .ZN(n1112) );
XOR2_X1 U800 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U801 ( .A(KEYINPUT14), .B(G116), .Z(n1116) );
NOR2_X1 U802 ( .A1(G898), .A2(n1084), .ZN(n1110) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1084), .ZN(n1105) );
AND2_X1 U804 ( .A1(G224), .A2(G898), .ZN(n1117) );
NOR3_X1 U805 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(G66) );
AND3_X1 U806 ( .A1(KEYINPUT63), .A2(G953), .A3(G952), .ZN(n1120) );
NOR2_X1 U807 ( .A1(KEYINPUT63), .A2(n1121), .ZN(n1119) );
INV_X1 U808 ( .A(n1122), .ZN(n1121) );
XNOR2_X1 U809 ( .A(n1123), .B(n1124), .ZN(n1118) );
NOR2_X1 U810 ( .A1(n1078), .A2(n1125), .ZN(n1123) );
NOR2_X1 U811 ( .A1(n1122), .A2(n1126), .ZN(G63) );
XNOR2_X1 U812 ( .A(n1127), .B(n1128), .ZN(n1126) );
AND2_X1 U813 ( .A1(G478), .A2(n1129), .ZN(n1128) );
NOR2_X1 U814 ( .A1(n1122), .A2(n1130), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1131), .B(n1132), .ZN(n1130) );
NAND2_X1 U816 ( .A1(KEYINPUT11), .A2(n1133), .ZN(n1131) );
NAND2_X1 U817 ( .A1(n1129), .A2(G475), .ZN(n1133) );
XOR2_X1 U818 ( .A(n1134), .B(n1135), .Z(G6) );
NOR2_X1 U819 ( .A1(n1136), .A2(n1137), .ZN(G57) );
XOR2_X1 U820 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U821 ( .A(KEYINPUT6), .B(KEYINPUT12), .Z(n1139) );
XOR2_X1 U822 ( .A(n1140), .B(n1141), .Z(n1138) );
NOR2_X1 U823 ( .A1(KEYINPUT3), .A2(n1142), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U825 ( .A1(n1145), .A2(n1125), .ZN(n1144) );
NOR2_X1 U826 ( .A1(n1146), .A2(n1147), .ZN(n1143) );
XOR2_X1 U827 ( .A(KEYINPUT10), .B(n1148), .Z(n1147) );
NOR2_X1 U828 ( .A1(n1084), .A2(n1149), .ZN(n1136) );
XOR2_X1 U829 ( .A(KEYINPUT7), .B(G952), .Z(n1149) );
NOR2_X1 U830 ( .A1(n1122), .A2(n1150), .ZN(G54) );
XOR2_X1 U831 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U832 ( .A1(G469), .A2(n1129), .ZN(n1152) );
INV_X1 U833 ( .A(n1125), .ZN(n1129) );
NOR2_X1 U834 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
XOR2_X1 U835 ( .A(KEYINPUT29), .B(n1155), .Z(n1154) );
NOR2_X1 U836 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XNOR2_X1 U837 ( .A(n1158), .B(KEYINPUT31), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
XOR2_X1 U839 ( .A(n1156), .B(KEYINPUT28), .Z(n1159) );
XOR2_X1 U840 ( .A(n1160), .B(n1161), .Z(n1156) );
XNOR2_X1 U841 ( .A(KEYINPUT40), .B(n1162), .ZN(n1160) );
NOR2_X1 U842 ( .A1(KEYINPUT49), .A2(n1163), .ZN(n1162) );
AND2_X1 U843 ( .A1(n1164), .A2(n1165), .ZN(n1158) );
NAND3_X1 U844 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
XNOR2_X1 U845 ( .A(KEYINPUT56), .B(n1169), .ZN(n1166) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1170), .ZN(n1164) );
NAND2_X1 U847 ( .A1(n1168), .A2(n1167), .ZN(n1170) );
XNOR2_X1 U848 ( .A(n1171), .B(KEYINPUT60), .ZN(n1168) );
XOR2_X1 U849 ( .A(n1172), .B(KEYINPUT19), .Z(n1169) );
NOR2_X1 U850 ( .A1(n1122), .A2(n1173), .ZN(G51) );
XOR2_X1 U851 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U852 ( .A(n1176), .B(n1177), .ZN(n1175) );
NAND2_X1 U853 ( .A1(KEYINPUT58), .A2(n1178), .ZN(n1177) );
NAND2_X1 U854 ( .A1(KEYINPUT18), .A2(n1179), .ZN(n1176) );
XOR2_X1 U855 ( .A(n1180), .B(n1181), .Z(n1174) );
NAND3_X1 U856 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1180) );
NAND2_X1 U857 ( .A1(KEYINPUT52), .A2(n1125), .ZN(n1183) );
NAND2_X1 U858 ( .A1(G902), .A2(n1030), .ZN(n1125) );
NAND2_X1 U859 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
INV_X1 U860 ( .A(KEYINPUT52), .ZN(n1186) );
OR2_X1 U861 ( .A1(n1030), .A2(n1187), .ZN(n1185) );
NAND4_X1 U862 ( .A1(n1188), .A2(n1109), .A3(n1189), .A4(n1095), .ZN(n1030) );
INV_X1 U863 ( .A(n1094), .ZN(n1189) );
NAND4_X1 U864 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1094) );
NOR4_X1 U865 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NAND2_X1 U866 ( .A1(KEYINPUT21), .A2(n1198), .ZN(n1192) );
INV_X1 U867 ( .A(n1199), .ZN(n1198) );
NAND3_X1 U868 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1191) );
NAND2_X1 U869 ( .A1(n1046), .A2(n1203), .ZN(n1201) );
OR4_X1 U870 ( .A1(n1040), .A2(n1204), .A3(n1052), .A4(KEYINPUT21), .ZN(n1203) );
NAND2_X1 U871 ( .A1(n1205), .A2(n1206), .ZN(n1200) );
NAND2_X1 U872 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
INV_X1 U873 ( .A(KEYINPUT38), .ZN(n1208) );
NAND2_X1 U874 ( .A1(KEYINPUT38), .A2(n1209), .ZN(n1190) );
AND4_X1 U875 ( .A1(n1135), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1109) );
AND4_X1 U876 ( .A1(n1213), .A2(n1214), .A3(n1025), .A4(n1215), .ZN(n1212) );
NAND3_X1 U877 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1025) );
NAND2_X1 U878 ( .A1(n1219), .A2(n1220), .ZN(n1211) );
INV_X1 U879 ( .A(n1060), .ZN(n1220) );
NOR2_X1 U880 ( .A1(n1202), .A2(n1216), .ZN(n1060) );
NAND3_X1 U881 ( .A1(n1221), .A2(n1046), .A3(n1222), .ZN(n1210) );
XOR2_X1 U882 ( .A(n1223), .B(KEYINPUT50), .Z(n1222) );
NAND3_X1 U883 ( .A1(n1218), .A2(n1217), .A3(n1202), .ZN(n1135) );
INV_X1 U884 ( .A(n1044), .ZN(n1217) );
XOR2_X1 U885 ( .A(n1224), .B(KEYINPUT35), .Z(n1188) );
NOR2_X1 U886 ( .A1(n1084), .A2(G952), .ZN(n1122) );
XOR2_X1 U887 ( .A(n1209), .B(n1225), .Z(G48) );
NOR2_X1 U888 ( .A1(KEYINPUT62), .A2(n1226), .ZN(n1225) );
AND3_X1 U889 ( .A1(n1202), .A2(n1046), .A3(n1207), .ZN(n1209) );
XOR2_X1 U890 ( .A(G143), .B(n1093), .Z(G45) );
INV_X1 U891 ( .A(n1224), .ZN(n1093) );
NAND4_X1 U892 ( .A1(n1227), .A2(n1046), .A3(n1228), .A4(n1229), .ZN(n1224) );
XOR2_X1 U893 ( .A(G140), .B(n1197), .Z(G42) );
AND4_X1 U894 ( .A1(n1061), .A2(n1202), .A3(n1230), .A4(n1052), .ZN(n1197) );
NOR2_X1 U895 ( .A1(n1204), .A2(n1231), .ZN(n1230) );
XOR2_X1 U896 ( .A(n1196), .B(n1232), .Z(G39) );
NOR2_X1 U897 ( .A1(KEYINPUT59), .A2(n1233), .ZN(n1232) );
AND3_X1 U898 ( .A1(n1061), .A2(n1234), .A3(n1207), .ZN(n1196) );
XOR2_X1 U899 ( .A(n1095), .B(n1235), .Z(G36) );
NAND2_X1 U900 ( .A1(KEYINPUT8), .A2(G134), .ZN(n1235) );
NAND3_X1 U901 ( .A1(n1227), .A2(n1216), .A3(n1061), .ZN(n1095) );
XOR2_X1 U902 ( .A(n1236), .B(n1237), .Z(G33) );
NAND2_X1 U903 ( .A1(KEYINPUT30), .A2(n1195), .ZN(n1237) );
AND3_X1 U904 ( .A1(n1227), .A2(n1202), .A3(n1061), .ZN(n1195) );
NOR2_X1 U905 ( .A1(n1047), .A2(n1066), .ZN(n1061) );
INV_X1 U906 ( .A(n1048), .ZN(n1066) );
NOR4_X1 U907 ( .A1(n1054), .A2(n1231), .A3(n1053), .A4(n1204), .ZN(n1227) );
INV_X1 U908 ( .A(n1238), .ZN(n1054) );
XOR2_X1 U909 ( .A(G128), .B(n1194), .Z(G30) );
AND3_X1 U910 ( .A1(n1216), .A2(n1046), .A3(n1207), .ZN(n1194) );
AND4_X1 U911 ( .A1(n1239), .A2(n1057), .A3(n1240), .A4(n1241), .ZN(n1207) );
XNOR2_X1 U912 ( .A(G101), .B(n1215), .ZN(G3) );
NAND4_X1 U913 ( .A1(n1234), .A2(n1218), .A3(n1238), .A4(n1240), .ZN(n1215) );
XOR2_X1 U914 ( .A(n1242), .B(n1199), .Z(G27) );
NAND4_X1 U915 ( .A1(n1202), .A2(n1052), .A3(n1243), .A4(n1063), .ZN(n1199) );
NOR2_X1 U916 ( .A1(n1204), .A2(n1206), .ZN(n1243) );
INV_X1 U917 ( .A(n1241), .ZN(n1204) );
NAND2_X1 U918 ( .A1(n1032), .A2(n1244), .ZN(n1241) );
NAND4_X1 U919 ( .A1(G953), .A2(G902), .A3(n1245), .A4(n1086), .ZN(n1244) );
INV_X1 U920 ( .A(G900), .ZN(n1086) );
NAND2_X1 U921 ( .A1(n1246), .A2(n1247), .ZN(G24) );
NAND4_X1 U922 ( .A1(n1248), .A2(n1221), .A3(n1223), .A4(n1249), .ZN(n1247) );
XOR2_X1 U923 ( .A(n1250), .B(KEYINPUT36), .Z(n1246) );
NAND2_X1 U924 ( .A1(G122), .A2(n1251), .ZN(n1250) );
NAND3_X1 U925 ( .A1(n1221), .A2(n1223), .A3(n1248), .ZN(n1251) );
XOR2_X1 U926 ( .A(n1206), .B(KEYINPUT2), .Z(n1248) );
NOR4_X1 U927 ( .A1(n1040), .A2(n1044), .A3(n1070), .A4(n1062), .ZN(n1221) );
NAND2_X1 U928 ( .A1(n1252), .A2(n1238), .ZN(n1044) );
XOR2_X1 U929 ( .A(n1214), .B(n1253), .Z(G21) );
NOR2_X1 U930 ( .A1(G119), .A2(KEYINPUT17), .ZN(n1253) );
NAND3_X1 U931 ( .A1(n1239), .A2(n1234), .A3(n1254), .ZN(n1214) );
XOR2_X1 U932 ( .A(n1255), .B(n1256), .Z(G18) );
NAND2_X1 U933 ( .A1(n1219), .A2(n1216), .ZN(n1256) );
NOR2_X1 U934 ( .A1(n1228), .A2(n1062), .ZN(n1216) );
INV_X1 U935 ( .A(n1070), .ZN(n1228) );
XNOR2_X1 U936 ( .A(G113), .B(n1257), .ZN(G15) );
NAND2_X1 U937 ( .A1(n1258), .A2(n1219), .ZN(n1257) );
AND2_X1 U938 ( .A1(n1254), .A2(n1238), .ZN(n1219) );
AND4_X1 U939 ( .A1(n1063), .A2(n1046), .A3(n1240), .A4(n1223), .ZN(n1254) );
INV_X1 U940 ( .A(n1053), .ZN(n1240) );
INV_X1 U941 ( .A(n1040), .ZN(n1063) );
NAND2_X1 U942 ( .A1(n1259), .A2(n1059), .ZN(n1040) );
XNOR2_X1 U943 ( .A(n1202), .B(KEYINPUT42), .ZN(n1258) );
NOR2_X1 U944 ( .A1(n1229), .A2(n1070), .ZN(n1202) );
INV_X1 U945 ( .A(n1062), .ZN(n1229) );
XNOR2_X1 U946 ( .A(G110), .B(n1213), .ZN(G12) );
NAND3_X1 U947 ( .A1(n1234), .A2(n1218), .A3(n1052), .ZN(n1213) );
AND2_X1 U948 ( .A1(n1252), .A2(n1239), .ZN(n1052) );
XOR2_X1 U949 ( .A(n1238), .B(KEYINPUT46), .Z(n1239) );
XOR2_X1 U950 ( .A(n1074), .B(n1079), .Z(n1238) );
INV_X1 U951 ( .A(n1078), .ZN(n1079) );
NAND2_X1 U952 ( .A1(G217), .A2(n1260), .ZN(n1078) );
NAND2_X1 U953 ( .A1(n1124), .A2(n1261), .ZN(n1074) );
XOR2_X1 U954 ( .A(n1262), .B(n1263), .Z(n1124) );
XOR2_X1 U955 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U956 ( .A(G146), .B(G110), .Z(n1265) );
NOR2_X1 U957 ( .A1(KEYINPUT16), .A2(G137), .ZN(n1264) );
XOR2_X1 U958 ( .A(n1266), .B(n1267), .Z(n1262) );
NOR2_X1 U959 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U960 ( .A(n1270), .B(KEYINPUT32), .Z(n1269) );
NAND2_X1 U961 ( .A1(G128), .A2(n1271), .ZN(n1270) );
NOR2_X1 U962 ( .A1(G128), .A2(n1271), .ZN(n1268) );
XOR2_X1 U963 ( .A(n1272), .B(n1273), .Z(n1266) );
NAND2_X1 U964 ( .A1(n1274), .A2(G221), .ZN(n1272) );
XOR2_X1 U965 ( .A(n1053), .B(KEYINPUT48), .Z(n1252) );
XOR2_X1 U966 ( .A(n1080), .B(n1275), .Z(n1053) );
NOR2_X1 U967 ( .A1(KEYINPUT26), .A2(n1145), .ZN(n1275) );
INV_X1 U968 ( .A(G472), .ZN(n1145) );
NAND2_X1 U969 ( .A1(n1261), .A2(n1276), .ZN(n1080) );
XOR2_X1 U970 ( .A(n1277), .B(n1140), .Z(n1276) );
XOR2_X1 U971 ( .A(n1278), .B(G101), .Z(n1140) );
NAND2_X1 U972 ( .A1(n1279), .A2(G210), .ZN(n1278) );
OR2_X1 U973 ( .A1(n1148), .A2(n1146), .ZN(n1277) );
AND2_X1 U974 ( .A1(n1280), .A2(n1281), .ZN(n1146) );
NOR2_X1 U975 ( .A1(n1281), .A2(n1280), .ZN(n1148) );
XOR2_X1 U976 ( .A(n1172), .B(n1282), .Z(n1280) );
XOR2_X1 U977 ( .A(n1283), .B(n1284), .Z(n1281) );
XNOR2_X1 U978 ( .A(n1285), .B(KEYINPUT55), .ZN(n1284) );
NAND2_X1 U979 ( .A1(n1286), .A2(KEYINPUT39), .ZN(n1285) );
XOR2_X1 U980 ( .A(n1255), .B(KEYINPUT44), .Z(n1286) );
INV_X1 U981 ( .A(G116), .ZN(n1255) );
AND3_X1 U982 ( .A1(n1057), .A2(n1223), .A3(n1046), .ZN(n1218) );
INV_X1 U983 ( .A(n1206), .ZN(n1046) );
NAND2_X1 U984 ( .A1(n1047), .A2(n1048), .ZN(n1206) );
NAND2_X1 U985 ( .A1(G214), .A2(n1287), .ZN(n1048) );
XNOR2_X1 U986 ( .A(n1072), .B(n1184), .ZN(n1047) );
INV_X1 U987 ( .A(n1073), .ZN(n1184) );
NAND2_X1 U988 ( .A1(G210), .A2(n1287), .ZN(n1073) );
NAND2_X1 U989 ( .A1(n1288), .A2(n1187), .ZN(n1287) );
INV_X1 U990 ( .A(G237), .ZN(n1288) );
NAND4_X1 U991 ( .A1(n1289), .A2(n1290), .A3(n1291), .A4(n1292), .ZN(n1072) );
NAND2_X1 U992 ( .A1(KEYINPUT57), .A2(n1293), .ZN(n1292) );
NAND2_X1 U993 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XOR2_X1 U994 ( .A(n1178), .B(KEYINPUT43), .Z(n1294) );
NAND2_X1 U995 ( .A1(n1296), .A2(n1297), .ZN(n1291) );
INV_X1 U996 ( .A(KEYINPUT57), .ZN(n1297) );
NAND2_X1 U997 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
OR2_X1 U998 ( .A1(n1300), .A2(KEYINPUT43), .ZN(n1299) );
NAND3_X1 U999 ( .A1(n1300), .A2(n1295), .A3(KEYINPUT43), .ZN(n1298) );
OR2_X1 U1000 ( .A1(n1300), .A2(n1295), .ZN(n1290) );
XOR2_X1 U1001 ( .A(n1181), .B(n1179), .Z(n1295) );
XNOR2_X1 U1002 ( .A(G125), .B(n1282), .ZN(n1179) );
XOR2_X1 U1003 ( .A(G128), .B(n1301), .Z(n1282) );
NOR2_X1 U1004 ( .A1(KEYINPUT53), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1005 ( .A(G143), .B(n1226), .Z(n1302) );
AND2_X1 U1006 ( .A1(G224), .A2(n1084), .ZN(n1181) );
INV_X1 U1007 ( .A(n1178), .ZN(n1300) );
XOR2_X1 U1008 ( .A(n1303), .B(n1304), .Z(n1178) );
INV_X1 U1009 ( .A(n1115), .ZN(n1304) );
XOR2_X1 U1010 ( .A(n1283), .B(n1305), .Z(n1115) );
XNOR2_X1 U1011 ( .A(G101), .B(n1306), .ZN(n1305) );
NAND2_X1 U1012 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1013 ( .A1(G104), .A2(n1022), .ZN(n1308) );
XOR2_X1 U1014 ( .A(n1309), .B(KEYINPUT27), .Z(n1307) );
NAND2_X1 U1015 ( .A1(G107), .A2(n1134), .ZN(n1309) );
XOR2_X1 U1016 ( .A(G113), .B(n1271), .Z(n1283) );
INV_X1 U1017 ( .A(G119), .ZN(n1271) );
XNOR2_X1 U1018 ( .A(G110), .B(n1310), .ZN(n1303) );
XOR2_X1 U1019 ( .A(n1261), .B(KEYINPUT1), .Z(n1289) );
NAND2_X1 U1020 ( .A1(n1032), .A2(n1311), .ZN(n1223) );
NAND4_X1 U1021 ( .A1(n1312), .A2(G953), .A3(G902), .A4(n1245), .ZN(n1311) );
XNOR2_X1 U1022 ( .A(G898), .B(KEYINPUT33), .ZN(n1312) );
NAND3_X1 U1023 ( .A1(n1245), .A2(n1084), .A3(G952), .ZN(n1032) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1245) );
INV_X1 U1025 ( .A(n1231), .ZN(n1057) );
NAND2_X1 U1026 ( .A1(n1058), .A2(n1059), .ZN(n1231) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1260), .ZN(n1059) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1187), .ZN(n1260) );
INV_X1 U1029 ( .A(n1259), .ZN(n1058) );
XOR2_X1 U1030 ( .A(n1313), .B(G469), .Z(n1259) );
NAND2_X1 U1031 ( .A1(n1314), .A2(n1261), .ZN(n1313) );
XOR2_X1 U1032 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1033 ( .A(n1161), .B(n1163), .Z(n1316) );
XOR2_X1 U1034 ( .A(G140), .B(KEYINPUT34), .Z(n1163) );
XOR2_X1 U1035 ( .A(G110), .B(n1317), .Z(n1161) );
NOR2_X1 U1036 ( .A1(G953), .A2(n1085), .ZN(n1317) );
INV_X1 U1037 ( .A(G227), .ZN(n1085) );
XOR2_X1 U1038 ( .A(n1318), .B(n1319), .Z(n1315) );
AND2_X1 U1039 ( .A1(n1167), .A2(n1171), .ZN(n1319) );
NAND2_X1 U1040 ( .A1(n1320), .A2(n1101), .ZN(n1171) );
OR2_X1 U1041 ( .A1(n1101), .A2(n1320), .ZN(n1167) );
XOR2_X1 U1042 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1043 ( .A(G104), .B(G101), .Z(n1322) );
NAND2_X1 U1044 ( .A1(KEYINPUT15), .A2(n1022), .ZN(n1321) );
INV_X1 U1045 ( .A(G107), .ZN(n1022) );
XNOR2_X1 U1046 ( .A(n1226), .B(n1323), .ZN(n1101) );
NAND2_X1 U1047 ( .A1(KEYINPUT9), .A2(n1172), .ZN(n1318) );
XOR2_X1 U1048 ( .A(n1104), .B(n1236), .Z(n1172) );
INV_X1 U1049 ( .A(G131), .ZN(n1236) );
XNOR2_X1 U1050 ( .A(n1233), .B(n1324), .ZN(n1104) );
INV_X1 U1051 ( .A(G137), .ZN(n1233) );
INV_X1 U1052 ( .A(n1036), .ZN(n1234) );
NAND2_X1 U1053 ( .A1(n1062), .A2(n1070), .ZN(n1036) );
XOR2_X1 U1054 ( .A(n1325), .B(G475), .Z(n1070) );
NAND2_X1 U1055 ( .A1(n1261), .A2(n1132), .ZN(n1325) );
XOR2_X1 U1056 ( .A(n1326), .B(n1327), .Z(n1132) );
XOR2_X1 U1057 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1058 ( .A(n1330), .B(n1331), .Z(n1329) );
NOR2_X1 U1059 ( .A1(KEYINPUT20), .A2(G143), .ZN(n1331) );
NAND2_X1 U1060 ( .A1(n1279), .A2(G214), .ZN(n1330) );
NOR2_X1 U1061 ( .A1(G953), .A2(G237), .ZN(n1279) );
NAND2_X1 U1062 ( .A1(n1332), .A2(n1333), .ZN(n1328) );
NAND2_X1 U1063 ( .A1(G146), .A2(n1334), .ZN(n1333) );
NAND2_X1 U1064 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
XNOR2_X1 U1065 ( .A(KEYINPUT61), .B(n1337), .ZN(n1335) );
NAND2_X1 U1066 ( .A1(n1338), .A2(n1226), .ZN(n1332) );
INV_X1 U1067 ( .A(G146), .ZN(n1226) );
NAND2_X1 U1068 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
OR2_X1 U1069 ( .A1(n1337), .A2(KEYINPUT61), .ZN(n1340) );
NAND2_X1 U1070 ( .A1(n1273), .A2(KEYINPUT61), .ZN(n1339) );
INV_X1 U1071 ( .A(n1097), .ZN(n1273) );
NAND2_X1 U1072 ( .A1(n1337), .A2(n1336), .ZN(n1097) );
NAND2_X1 U1073 ( .A1(G140), .A2(n1242), .ZN(n1336) );
OR2_X1 U1074 ( .A1(n1242), .A2(G140), .ZN(n1337) );
INV_X1 U1075 ( .A(G125), .ZN(n1242) );
XOR2_X1 U1076 ( .A(n1341), .B(n1342), .Z(n1326) );
NOR2_X1 U1077 ( .A1(KEYINPUT5), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1078 ( .A(G113), .B(n1249), .Z(n1343) );
INV_X1 U1079 ( .A(G122), .ZN(n1249) );
XOR2_X1 U1080 ( .A(n1134), .B(G131), .Z(n1341) );
INV_X1 U1081 ( .A(G104), .ZN(n1134) );
XOR2_X1 U1082 ( .A(n1344), .B(G478), .Z(n1062) );
NAND2_X1 U1083 ( .A1(n1261), .A2(n1127), .ZN(n1344) );
XNOR2_X1 U1084 ( .A(n1345), .B(n1346), .ZN(n1127) );
XOR2_X1 U1085 ( .A(n1323), .B(n1310), .Z(n1346) );
XOR2_X1 U1086 ( .A(G116), .B(G122), .Z(n1310) );
XOR2_X1 U1087 ( .A(G128), .B(G143), .Z(n1323) );
XOR2_X1 U1088 ( .A(n1347), .B(n1324), .Z(n1345) );
XOR2_X1 U1089 ( .A(G134), .B(KEYINPUT41), .Z(n1324) );
XOR2_X1 U1090 ( .A(n1348), .B(G107), .Z(n1347) );
NAND2_X1 U1091 ( .A1(G217), .A2(n1274), .ZN(n1348) );
AND2_X1 U1092 ( .A1(G234), .A2(n1084), .ZN(n1274) );
INV_X1 U1093 ( .A(G953), .ZN(n1084) );
XOR2_X1 U1094 ( .A(n1187), .B(KEYINPUT0), .Z(n1261) );
INV_X1 U1095 ( .A(G902), .ZN(n1187) );
endmodule


