//Key = 0100001110111101000011001000011111110010001000100111111111011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369;

XNOR2_X1 U741 ( .A(G107), .B(n1035), .ZN(G9) );
NOR2_X1 U742 ( .A1(n1036), .A2(n1037), .ZN(G75) );
XOR2_X1 U743 ( .A(n1038), .B(KEYINPUT10), .Z(n1037) );
OR3_X1 U744 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
OR3_X1 U745 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NOR3_X1 U746 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
INV_X1 U747 ( .A(n1048), .ZN(n1047) );
NOR2_X1 U748 ( .A1(n1049), .A2(n1050), .ZN(n1046) );
NOR2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U751 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
XNOR2_X1 U753 ( .A(n1059), .B(n1060), .ZN(n1058) );
NOR2_X1 U754 ( .A1(KEYINPUT38), .A2(n1061), .ZN(n1057) );
NOR2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1053) );
NOR2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
AND3_X1 U757 ( .A1(KEYINPUT38), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR3_X1 U758 ( .A1(n1068), .A2(n1061), .A3(n1056), .ZN(n1049) );
XOR2_X1 U759 ( .A(KEYINPUT6), .B(n1069), .Z(n1068) );
NOR3_X1 U760 ( .A1(n1056), .A2(n1061), .A3(n1070), .ZN(n1043) );
NOR2_X1 U761 ( .A1(n1071), .A2(n1063), .ZN(n1070) );
NOR3_X1 U762 ( .A1(n1052), .A2(n1072), .A3(n1073), .ZN(n1071) );
NOR3_X1 U763 ( .A1(n1045), .A2(n1074), .A3(n1075), .ZN(n1073) );
NOR2_X1 U764 ( .A1(KEYINPUT25), .A2(n1076), .ZN(n1075) );
NOR2_X1 U765 ( .A1(KEYINPUT19), .A2(n1077), .ZN(n1074) );
INV_X1 U766 ( .A(n1078), .ZN(n1077) );
NOR2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1072) );
AND2_X1 U768 ( .A1(n1078), .A2(KEYINPUT19), .ZN(n1080) );
AND2_X1 U769 ( .A1(n1081), .A2(n1063), .ZN(n1061) );
INV_X1 U770 ( .A(n1082), .ZN(n1063) );
NAND4_X1 U771 ( .A1(KEYINPUT25), .A2(n1079), .A3(n1083), .A4(n1084), .ZN(n1081) );
INV_X1 U772 ( .A(n1045), .ZN(n1079) );
XOR2_X1 U773 ( .A(n1085), .B(KEYINPUT42), .Z(n1042) );
NAND4_X1 U774 ( .A1(n1082), .A2(n1086), .A3(n1048), .A4(n1087), .ZN(n1085) );
NOR3_X1 U775 ( .A1(n1088), .A2(n1056), .A3(n1045), .ZN(n1087) );
INV_X1 U776 ( .A(n1089), .ZN(n1056) );
NOR2_X1 U777 ( .A1(G952), .A2(n1040), .ZN(n1036) );
NAND2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1040) );
NAND4_X1 U779 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
NOR3_X1 U780 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
XOR2_X1 U781 ( .A(n1099), .B(KEYINPUT15), .Z(n1097) );
NAND3_X1 U782 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1096) );
XNOR2_X1 U783 ( .A(G472), .B(n1103), .ZN(n1102) );
NOR2_X1 U784 ( .A1(KEYINPUT4), .A2(n1104), .ZN(n1103) );
NAND2_X1 U785 ( .A1(n1105), .A2(n1106), .ZN(n1101) );
XOR2_X1 U786 ( .A(KEYINPUT23), .B(n1107), .Z(n1105) );
NAND2_X1 U787 ( .A1(n1108), .A2(G478), .ZN(n1100) );
XOR2_X1 U788 ( .A(KEYINPUT13), .B(n1107), .Z(n1108) );
NOR3_X1 U789 ( .A1(n1067), .A2(n1109), .A3(n1110), .ZN(n1094) );
NAND2_X1 U790 ( .A1(G475), .A2(n1111), .ZN(n1093) );
XNOR2_X1 U791 ( .A(KEYINPUT5), .B(n1112), .ZN(n1092) );
XOR2_X1 U792 ( .A(n1113), .B(n1114), .Z(G72) );
NOR2_X1 U793 ( .A1(n1115), .A2(n1090), .ZN(n1114) );
NOR2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1113) );
NAND2_X1 U796 ( .A1(n1120), .A2(n1090), .ZN(n1119) );
XOR2_X1 U797 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U798 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
OR3_X1 U799 ( .A1(n1117), .A2(n1122), .A3(n1090), .ZN(n1118) );
XNOR2_X1 U800 ( .A(n1125), .B(n1126), .ZN(n1122) );
XOR2_X1 U801 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1125) );
XOR2_X1 U803 ( .A(KEYINPUT9), .B(G131), .Z(n1130) );
NAND2_X1 U804 ( .A1(KEYINPUT21), .A2(n1131), .ZN(n1129) );
NAND2_X1 U805 ( .A1(n1132), .A2(n1133), .ZN(G69) );
NAND2_X1 U806 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U807 ( .A(KEYINPUT60), .B(n1136), .Z(n1132) );
NOR2_X1 U808 ( .A1(n1134), .A2(n1137), .ZN(n1136) );
XOR2_X1 U809 ( .A(n1135), .B(KEYINPUT16), .Z(n1137) );
NAND2_X1 U810 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
NAND2_X1 U811 ( .A1(G953), .A2(n1140), .ZN(n1139) );
AND2_X1 U812 ( .A1(n1141), .A2(n1142), .ZN(n1134) );
NAND2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U814 ( .A1(n1145), .A2(n1138), .ZN(n1144) );
INV_X1 U815 ( .A(n1146), .ZN(n1143) );
NAND3_X1 U816 ( .A1(n1145), .A2(n1138), .A3(n1146), .ZN(n1141) );
NAND2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U818 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XNOR2_X1 U819 ( .A(KEYINPUT8), .B(n1090), .ZN(n1147) );
INV_X1 U820 ( .A(n1151), .ZN(n1138) );
XOR2_X1 U821 ( .A(n1152), .B(n1153), .Z(n1145) );
NOR2_X1 U822 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U823 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND3_X1 U824 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1156) );
XNOR2_X1 U825 ( .A(G217), .B(KEYINPUT20), .ZN(n1160) );
NOR3_X1 U826 ( .A1(n1154), .A2(n1161), .A3(n1162), .ZN(G63) );
NOR2_X1 U827 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U828 ( .A(n1165), .B(KEYINPUT40), .Z(n1164) );
NOR2_X1 U829 ( .A1(n1166), .A2(n1167), .ZN(n1161) );
XOR2_X1 U830 ( .A(n1165), .B(KEYINPUT35), .Z(n1167) );
NAND2_X1 U831 ( .A1(n1158), .A2(G478), .ZN(n1165) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1168), .ZN(G60) );
XOR2_X1 U833 ( .A(n1169), .B(n1170), .Z(n1168) );
NAND2_X1 U834 ( .A1(n1158), .A2(G475), .ZN(n1169) );
XNOR2_X1 U835 ( .A(G104), .B(n1171), .ZN(G6) );
NOR2_X1 U836 ( .A1(n1154), .A2(n1172), .ZN(G57) );
XOR2_X1 U837 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U838 ( .A(n1175), .B(n1176), .ZN(n1174) );
NAND2_X1 U839 ( .A1(n1158), .A2(G472), .ZN(n1175) );
XNOR2_X1 U840 ( .A(n1177), .B(n1178), .ZN(n1173) );
NAND2_X1 U841 ( .A1(n1179), .A2(KEYINPUT24), .ZN(n1178) );
XOR2_X1 U842 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U843 ( .A(KEYINPUT26), .B(n1182), .ZN(n1181) );
NAND2_X1 U844 ( .A1(KEYINPUT54), .A2(n1183), .ZN(n1180) );
NAND2_X1 U845 ( .A1(KEYINPUT1), .A2(n1184), .ZN(n1177) );
NOR2_X1 U846 ( .A1(n1154), .A2(n1185), .ZN(G54) );
XNOR2_X1 U847 ( .A(n1186), .B(n1187), .ZN(n1185) );
XOR2_X1 U848 ( .A(n1188), .B(n1189), .Z(n1187) );
NAND2_X1 U849 ( .A1(n1158), .A2(G469), .ZN(n1189) );
NAND2_X1 U850 ( .A1(n1190), .A2(KEYINPUT62), .ZN(n1188) );
XNOR2_X1 U851 ( .A(G140), .B(n1191), .ZN(n1190) );
NOR2_X1 U852 ( .A1(n1154), .A2(n1192), .ZN(G51) );
XOR2_X1 U853 ( .A(n1193), .B(n1194), .Z(n1192) );
XNOR2_X1 U854 ( .A(n1195), .B(n1196), .ZN(n1194) );
XNOR2_X1 U855 ( .A(G125), .B(n1197), .ZN(n1193) );
NAND3_X1 U856 ( .A1(G210), .A2(n1198), .A3(n1158), .ZN(n1197) );
AND2_X1 U857 ( .A1(n1199), .A2(n1039), .ZN(n1158) );
NAND4_X1 U858 ( .A1(n1149), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1039) );
XNOR2_X1 U859 ( .A(KEYINPUT47), .B(n1123), .ZN(n1202) );
NAND4_X1 U860 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1123) );
NAND3_X1 U861 ( .A1(n1207), .A2(n1048), .A3(n1089), .ZN(n1203) );
XNOR2_X1 U862 ( .A(KEYINPUT12), .B(n1150), .ZN(n1201) );
INV_X1 U863 ( .A(n1124), .ZN(n1200) );
NAND4_X1 U864 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1124) );
NAND3_X1 U865 ( .A1(n1212), .A2(n1078), .A3(n1213), .ZN(n1208) );
XNOR2_X1 U866 ( .A(n1089), .B(KEYINPUT51), .ZN(n1213) );
AND4_X1 U867 ( .A1(n1214), .A2(n1215), .A3(n1171), .A4(n1216), .ZN(n1149) );
AND4_X1 U868 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1035), .ZN(n1216) );
NAND4_X1 U869 ( .A1(n1069), .A2(n1078), .A3(n1220), .A4(n1082), .ZN(n1035) );
NAND4_X1 U870 ( .A1(n1083), .A2(n1069), .A3(n1220), .A4(n1082), .ZN(n1171) );
XNOR2_X1 U871 ( .A(G902), .B(KEYINPUT61), .ZN(n1199) );
NOR2_X1 U872 ( .A1(n1090), .A2(G952), .ZN(n1154) );
XNOR2_X1 U873 ( .A(G146), .B(n1204), .ZN(G48) );
NAND3_X1 U874 ( .A1(n1083), .A2(n1065), .A3(n1207), .ZN(n1204) );
XNOR2_X1 U875 ( .A(G143), .B(n1205), .ZN(G45) );
NAND4_X1 U876 ( .A1(n1212), .A2(n1065), .A3(n1221), .A4(n1222), .ZN(n1205) );
XNOR2_X1 U877 ( .A(G140), .B(n1206), .ZN(G42) );
NAND3_X1 U878 ( .A1(n1223), .A2(n1069), .A3(n1089), .ZN(n1206) );
XNOR2_X1 U879 ( .A(G137), .B(n1224), .ZN(G39) );
NAND4_X1 U880 ( .A1(n1225), .A2(n1226), .A3(n1089), .A4(n1060), .ZN(n1224) );
XOR2_X1 U881 ( .A(n1227), .B(KEYINPUT36), .Z(n1225) );
XNOR2_X1 U882 ( .A(G134), .B(n1228), .ZN(G36) );
NAND2_X1 U883 ( .A1(n1229), .A2(n1078), .ZN(n1228) );
XNOR2_X1 U884 ( .A(G131), .B(n1209), .ZN(G33) );
NAND2_X1 U885 ( .A1(n1229), .A2(n1083), .ZN(n1209) );
AND2_X1 U886 ( .A1(n1212), .A2(n1089), .ZN(n1229) );
NOR2_X1 U887 ( .A1(n1112), .A2(n1067), .ZN(n1089) );
AND2_X1 U888 ( .A1(n1230), .A2(n1059), .ZN(n1212) );
XNOR2_X1 U889 ( .A(G128), .B(n1210), .ZN(G30) );
NAND3_X1 U890 ( .A1(n1078), .A2(n1065), .A3(n1207), .ZN(n1210) );
AND2_X1 U891 ( .A1(n1230), .A2(n1231), .ZN(n1207) );
AND3_X1 U892 ( .A1(n1060), .A2(n1227), .A3(n1069), .ZN(n1230) );
XNOR2_X1 U893 ( .A(n1232), .B(n1214), .ZN(G3) );
NAND3_X1 U894 ( .A1(n1048), .A2(n1069), .A3(n1233), .ZN(n1214) );
NOR3_X1 U895 ( .A1(n1234), .A2(n1235), .A3(n1231), .ZN(n1233) );
NAND2_X1 U896 ( .A1(KEYINPUT11), .A2(n1182), .ZN(n1232) );
XNOR2_X1 U897 ( .A(G125), .B(n1211), .ZN(G27) );
NAND3_X1 U898 ( .A1(n1084), .A2(n1065), .A3(n1223), .ZN(n1211) );
AND4_X1 U899 ( .A1(n1235), .A2(n1083), .A3(n1231), .A4(n1227), .ZN(n1223) );
NAND2_X1 U900 ( .A1(n1045), .A2(n1236), .ZN(n1227) );
NAND4_X1 U901 ( .A1(G902), .A2(G953), .A3(n1237), .A4(n1117), .ZN(n1236) );
INV_X1 U902 ( .A(G900), .ZN(n1117) );
XOR2_X1 U903 ( .A(n1215), .B(n1238), .Z(G24) );
NAND2_X1 U904 ( .A1(n1239), .A2(KEYINPUT29), .ZN(n1238) );
XNOR2_X1 U905 ( .A(G122), .B(KEYINPUT46), .ZN(n1239) );
NAND3_X1 U906 ( .A1(n1084), .A2(n1220), .A3(n1240), .ZN(n1215) );
AND3_X1 U907 ( .A1(n1082), .A2(n1222), .A3(n1221), .ZN(n1240) );
NOR2_X1 U908 ( .A1(n1060), .A2(n1231), .ZN(n1082) );
INV_X1 U909 ( .A(n1052), .ZN(n1084) );
XNOR2_X1 U910 ( .A(G119), .B(n1219), .ZN(G21) );
NAND3_X1 U911 ( .A1(n1241), .A2(n1231), .A3(n1048), .ZN(n1219) );
XNOR2_X1 U912 ( .A(G116), .B(n1218), .ZN(G18) );
NAND3_X1 U913 ( .A1(n1059), .A2(n1078), .A3(n1241), .ZN(n1218) );
NOR2_X1 U914 ( .A1(n1222), .A2(n1242), .ZN(n1078) );
XNOR2_X1 U915 ( .A(G113), .B(n1217), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1059), .A2(n1083), .A3(n1241), .ZN(n1217) );
NOR3_X1 U917 ( .A1(n1234), .A2(n1235), .A3(n1052), .ZN(n1241) );
NAND2_X1 U918 ( .A1(n1086), .A2(n1088), .ZN(n1052) );
INV_X1 U919 ( .A(n1076), .ZN(n1083) );
NAND2_X1 U920 ( .A1(n1242), .A2(n1222), .ZN(n1076) );
INV_X1 U921 ( .A(n1231), .ZN(n1059) );
XNOR2_X1 U922 ( .A(n1243), .B(n1150), .ZN(G12) );
NAND3_X1 U923 ( .A1(n1235), .A2(n1220), .A3(n1226), .ZN(n1150) );
AND3_X1 U924 ( .A1(n1069), .A2(n1231), .A3(n1048), .ZN(n1226) );
NOR2_X1 U925 ( .A1(n1221), .A2(n1222), .ZN(n1048) );
NAND3_X1 U926 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1222) );
INV_X1 U927 ( .A(n1109), .ZN(n1246) );
NOR2_X1 U928 ( .A1(n1111), .A2(G475), .ZN(n1109) );
NAND3_X1 U929 ( .A1(G475), .A2(n1111), .A3(n1247), .ZN(n1245) );
OR2_X1 U930 ( .A1(n1247), .A2(n1111), .ZN(n1244) );
NAND2_X1 U931 ( .A1(n1170), .A2(n1248), .ZN(n1111) );
XNOR2_X1 U932 ( .A(n1249), .B(n1250), .ZN(n1170) );
NOR2_X1 U933 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XOR2_X1 U934 ( .A(KEYINPUT48), .B(n1253), .Z(n1252) );
NOR2_X1 U935 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
AND2_X1 U936 ( .A1(n1255), .A2(n1254), .ZN(n1251) );
NAND2_X1 U937 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
NAND2_X1 U938 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U939 ( .A(KEYINPUT43), .B(n1260), .Z(n1258) );
NAND2_X1 U940 ( .A1(n1261), .A2(G146), .ZN(n1256) );
XNOR2_X1 U941 ( .A(n1260), .B(KEYINPUT44), .ZN(n1261) );
XNOR2_X1 U942 ( .A(n1262), .B(n1263), .ZN(n1255) );
XNOR2_X1 U943 ( .A(n1264), .B(G131), .ZN(n1263) );
NAND2_X1 U944 ( .A1(G214), .A2(n1265), .ZN(n1262) );
XNOR2_X1 U945 ( .A(G104), .B(n1266), .ZN(n1249) );
NOR2_X1 U946 ( .A1(KEYINPUT22), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U947 ( .A(G113), .B(n1268), .ZN(n1267) );
INV_X1 U948 ( .A(KEYINPUT39), .ZN(n1247) );
INV_X1 U949 ( .A(n1242), .ZN(n1221) );
XOR2_X1 U950 ( .A(n1107), .B(n1106), .Z(n1242) );
INV_X1 U951 ( .A(G478), .ZN(n1106) );
NOR2_X1 U952 ( .A1(n1163), .A2(G902), .ZN(n1107) );
INV_X1 U953 ( .A(n1166), .ZN(n1163) );
XNOR2_X1 U954 ( .A(n1269), .B(n1270), .ZN(n1166) );
AND2_X1 U955 ( .A1(n1271), .A2(G217), .ZN(n1270) );
NAND2_X1 U956 ( .A1(KEYINPUT52), .A2(n1272), .ZN(n1269) );
NAND2_X1 U957 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U958 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XNOR2_X1 U959 ( .A(n1277), .B(n1278), .ZN(n1276) );
INV_X1 U960 ( .A(n1279), .ZN(n1278) );
XOR2_X1 U961 ( .A(n1280), .B(n1281), .Z(n1275) );
XOR2_X1 U962 ( .A(n1282), .B(KEYINPUT27), .Z(n1273) );
NAND2_X1 U963 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XNOR2_X1 U964 ( .A(n1280), .B(n1281), .ZN(n1284) );
XNOR2_X1 U965 ( .A(G128), .B(n1264), .ZN(n1281) );
NAND2_X1 U966 ( .A1(KEYINPUT7), .A2(n1131), .ZN(n1280) );
XNOR2_X1 U967 ( .A(n1279), .B(n1277), .ZN(n1283) );
AND2_X1 U968 ( .A1(KEYINPUT49), .A2(n1285), .ZN(n1277) );
XNOR2_X1 U969 ( .A(n1099), .B(KEYINPUT37), .ZN(n1231) );
XOR2_X1 U970 ( .A(n1286), .B(n1287), .Z(n1099) );
NOR2_X1 U971 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
INV_X1 U972 ( .A(G217), .ZN(n1289) );
NOR2_X1 U973 ( .A1(G902), .A2(n1290), .ZN(n1288) );
NAND2_X1 U974 ( .A1(n1157), .A2(n1248), .ZN(n1286) );
XNOR2_X1 U975 ( .A(n1291), .B(n1292), .ZN(n1157) );
XOR2_X1 U976 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U977 ( .A(G110), .B(G119), .ZN(n1294) );
NAND2_X1 U978 ( .A1(n1271), .A2(G221), .ZN(n1293) );
NOR2_X1 U979 ( .A1(n1290), .A2(G953), .ZN(n1271) );
INV_X1 U980 ( .A(G234), .ZN(n1290) );
XNOR2_X1 U981 ( .A(n1127), .B(n1295), .ZN(n1291) );
XOR2_X1 U982 ( .A(G137), .B(n1260), .Z(n1127) );
XNOR2_X1 U983 ( .A(n1296), .B(G140), .ZN(n1260) );
NOR2_X1 U984 ( .A1(n1086), .A2(n1110), .ZN(n1069) );
INV_X1 U985 ( .A(n1088), .ZN(n1110) );
NAND2_X1 U986 ( .A1(G221), .A2(n1159), .ZN(n1088) );
NAND2_X1 U987 ( .A1(G234), .A2(n1248), .ZN(n1159) );
XOR2_X1 U988 ( .A(n1098), .B(KEYINPUT59), .Z(n1086) );
XNOR2_X1 U989 ( .A(n1297), .B(G469), .ZN(n1098) );
NAND2_X1 U990 ( .A1(n1298), .A2(n1248), .ZN(n1297) );
XOR2_X1 U991 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U992 ( .A(n1191), .B(n1186), .ZN(n1300) );
XOR2_X1 U993 ( .A(n1128), .B(n1301), .Z(n1186) );
XNOR2_X1 U994 ( .A(n1302), .B(n1303), .ZN(n1301) );
NAND3_X1 U995 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1302) );
NAND2_X1 U996 ( .A1(n1307), .A2(n1182), .ZN(n1306) );
NAND2_X1 U997 ( .A1(n1308), .A2(n1309), .ZN(n1305) );
INV_X1 U998 ( .A(KEYINPUT33), .ZN(n1309) );
NAND2_X1 U999 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
XNOR2_X1 U1000 ( .A(KEYINPUT58), .B(n1182), .ZN(n1311) );
INV_X1 U1001 ( .A(n1307), .ZN(n1310) );
NAND2_X1 U1002 ( .A1(KEYINPUT33), .A2(n1312), .ZN(n1304) );
NAND2_X1 U1003 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
OR3_X1 U1004 ( .A1(n1182), .A2(n1307), .A3(KEYINPUT58), .ZN(n1314) );
XOR2_X1 U1005 ( .A(G104), .B(n1315), .Z(n1307) );
XOR2_X1 U1006 ( .A(KEYINPUT50), .B(G107), .Z(n1315) );
NAND2_X1 U1007 ( .A1(KEYINPUT58), .A2(n1182), .ZN(n1313) );
XNOR2_X1 U1008 ( .A(n1316), .B(n1317), .ZN(n1128) );
NOR2_X1 U1009 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
XOR2_X1 U1010 ( .A(KEYINPUT14), .B(n1320), .Z(n1319) );
NOR2_X1 U1011 ( .A1(G143), .A2(n1259), .ZN(n1320) );
NOR2_X1 U1012 ( .A1(G146), .A2(n1264), .ZN(n1318) );
INV_X1 U1013 ( .A(G143), .ZN(n1264) );
NAND2_X1 U1014 ( .A1(KEYINPUT53), .A2(G128), .ZN(n1316) );
XOR2_X1 U1015 ( .A(G110), .B(n1321), .Z(n1191) );
NOR2_X1 U1016 ( .A1(G953), .A2(n1116), .ZN(n1321) );
INV_X1 U1017 ( .A(G227), .ZN(n1116) );
XNOR2_X1 U1018 ( .A(KEYINPUT17), .B(n1322), .ZN(n1299) );
NOR2_X1 U1019 ( .A1(G140), .A2(KEYINPUT45), .ZN(n1322) );
INV_X1 U1020 ( .A(n1234), .ZN(n1220) );
NAND2_X1 U1021 ( .A1(n1065), .A2(n1323), .ZN(n1234) );
NAND2_X1 U1022 ( .A1(n1324), .A2(n1045), .ZN(n1323) );
NAND3_X1 U1023 ( .A1(n1237), .A2(n1090), .A3(G952), .ZN(n1045) );
NAND3_X1 U1024 ( .A1(n1151), .A2(n1237), .A3(G902), .ZN(n1324) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1237) );
NOR2_X1 U1026 ( .A1(G898), .A2(n1090), .ZN(n1151) );
INV_X1 U1027 ( .A(G953), .ZN(n1090) );
NOR2_X1 U1028 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
AND2_X1 U1029 ( .A1(G214), .A2(n1198), .ZN(n1067) );
NAND2_X1 U1030 ( .A1(n1325), .A2(n1248), .ZN(n1198) );
INV_X1 U1031 ( .A(n1112), .ZN(n1066) );
NAND2_X1 U1032 ( .A1(n1326), .A2(n1327), .ZN(n1112) );
NAND2_X1 U1033 ( .A1(G210), .A2(n1328), .ZN(n1327) );
NAND2_X1 U1034 ( .A1(n1248), .A2(n1329), .ZN(n1328) );
OR2_X1 U1035 ( .A1(n1325), .A2(n1330), .ZN(n1329) );
INV_X1 U1036 ( .A(G237), .ZN(n1325) );
NAND3_X1 U1037 ( .A1(n1331), .A2(n1248), .A3(n1330), .ZN(n1326) );
XNOR2_X1 U1038 ( .A(n1196), .B(n1332), .ZN(n1330) );
NOR2_X1 U1039 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
XOR2_X1 U1040 ( .A(n1335), .B(KEYINPUT55), .Z(n1334) );
NAND2_X1 U1041 ( .A1(n1336), .A2(n1296), .ZN(n1335) );
XNOR2_X1 U1042 ( .A(n1195), .B(KEYINPUT30), .ZN(n1336) );
NOR2_X1 U1043 ( .A1(n1296), .A2(n1195), .ZN(n1333) );
INV_X1 U1044 ( .A(G125), .ZN(n1296) );
XOR2_X1 U1045 ( .A(n1152), .B(n1337), .Z(n1196) );
XOR2_X1 U1046 ( .A(n1338), .B(n1339), .Z(n1337) );
NOR2_X1 U1047 ( .A1(n1153), .A2(KEYINPUT3), .ZN(n1339) );
AND2_X1 U1048 ( .A1(n1340), .A2(n1341), .ZN(n1153) );
NAND2_X1 U1049 ( .A1(G113), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1050 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XOR2_X1 U1051 ( .A(n1345), .B(KEYINPUT18), .Z(n1340) );
NAND3_X1 U1052 ( .A1(n1344), .A2(n1346), .A3(n1343), .ZN(n1345) );
XOR2_X1 U1053 ( .A(n1347), .B(KEYINPUT63), .Z(n1343) );
NOR2_X1 U1054 ( .A1(G953), .A2(n1140), .ZN(n1338) );
INV_X1 U1055 ( .A(G224), .ZN(n1140) );
XOR2_X1 U1056 ( .A(n1348), .B(n1349), .Z(n1152) );
XNOR2_X1 U1057 ( .A(n1350), .B(G101), .ZN(n1349) );
INV_X1 U1058 ( .A(G104), .ZN(n1350) );
XNOR2_X1 U1059 ( .A(n1279), .B(n1351), .ZN(n1348) );
NOR2_X1 U1060 ( .A1(KEYINPUT28), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1061 ( .A(G107), .B(n1268), .Z(n1279) );
XOR2_X1 U1062 ( .A(G122), .B(KEYINPUT2), .Z(n1268) );
NAND2_X1 U1063 ( .A1(G210), .A2(G237), .ZN(n1331) );
INV_X1 U1064 ( .A(n1060), .ZN(n1235) );
XNOR2_X1 U1065 ( .A(n1104), .B(G472), .ZN(n1060) );
NAND2_X1 U1066 ( .A1(n1353), .A2(n1248), .ZN(n1104) );
INV_X1 U1067 ( .A(G902), .ZN(n1248) );
XOR2_X1 U1068 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1069 ( .A(n1183), .B(n1356), .ZN(n1355) );
INV_X1 U1070 ( .A(n1176), .ZN(n1356) );
XOR2_X1 U1071 ( .A(n1195), .B(n1303), .Z(n1176) );
XNOR2_X1 U1072 ( .A(n1357), .B(n1358), .ZN(n1303) );
XOR2_X1 U1073 ( .A(KEYINPUT0), .B(G131), .Z(n1358) );
NAND3_X1 U1074 ( .A1(n1359), .A2(n1360), .A3(n1361), .ZN(n1357) );
NAND2_X1 U1075 ( .A1(G137), .A2(n1362), .ZN(n1361) );
OR3_X1 U1076 ( .A1(n1362), .A2(G137), .A3(n1363), .ZN(n1360) );
INV_X1 U1077 ( .A(KEYINPUT57), .ZN(n1363) );
NAND2_X1 U1078 ( .A1(KEYINPUT32), .A2(n1364), .ZN(n1362) );
OR2_X1 U1079 ( .A1(n1364), .A2(KEYINPUT57), .ZN(n1359) );
XOR2_X1 U1080 ( .A(n1131), .B(KEYINPUT41), .Z(n1364) );
INV_X1 U1081 ( .A(G134), .ZN(n1131) );
XOR2_X1 U1082 ( .A(G143), .B(n1295), .Z(n1195) );
XNOR2_X1 U1083 ( .A(G128), .B(n1259), .ZN(n1295) );
INV_X1 U1084 ( .A(G146), .ZN(n1259) );
NAND2_X1 U1085 ( .A1(G210), .A2(n1265), .ZN(n1183) );
NOR2_X1 U1086 ( .A1(G953), .A2(G237), .ZN(n1265) );
XNOR2_X1 U1087 ( .A(n1365), .B(n1182), .ZN(n1354) );
INV_X1 U1088 ( .A(G101), .ZN(n1182) );
NAND2_X1 U1089 ( .A1(KEYINPUT34), .A2(n1184), .ZN(n1365) );
AND2_X1 U1090 ( .A1(n1366), .A2(n1367), .ZN(n1184) );
NAND2_X1 U1091 ( .A1(n1368), .A2(n1346), .ZN(n1367) );
XOR2_X1 U1092 ( .A(KEYINPUT56), .B(n1369), .Z(n1366) );
NOR2_X1 U1093 ( .A1(n1368), .A2(n1346), .ZN(n1369) );
INV_X1 U1094 ( .A(G113), .ZN(n1346) );
AND2_X1 U1095 ( .A1(n1344), .A2(n1347), .ZN(n1368) );
NAND2_X1 U1096 ( .A1(G119), .A2(n1285), .ZN(n1347) );
OR2_X1 U1097 ( .A1(n1285), .A2(G119), .ZN(n1344) );
INV_X1 U1098 ( .A(G116), .ZN(n1285) );
NAND2_X1 U1099 ( .A1(KEYINPUT31), .A2(n1352), .ZN(n1243) );
INV_X1 U1100 ( .A(G110), .ZN(n1352) );
endmodule


