//Key = 0010101100001010111010010101010101101100110100000110100100101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316;

XNOR2_X1 U734 ( .A(G107), .B(n1005), .ZN(G9) );
NOR2_X1 U735 ( .A1(n1006), .A2(n1007), .ZN(G75) );
NOR4_X1 U736 ( .A1(G953), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1007) );
INV_X1 U737 ( .A(n1011), .ZN(n1010) );
NOR2_X1 U738 ( .A1(n1012), .A2(n1013), .ZN(n1009) );
NOR2_X1 U739 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR3_X1 U740 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NOR2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U742 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR3_X1 U743 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1021) );
NOR3_X1 U744 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NOR2_X1 U745 ( .A1(n1029), .A2(n1030), .ZN(n1023) );
NOR2_X1 U746 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U747 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(n1019) );
NOR2_X1 U749 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U750 ( .A1(n1022), .A2(n1039), .A3(n1036), .ZN(n1014) );
INV_X1 U751 ( .A(n1040), .ZN(n1036) );
NOR2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
INV_X1 U753 ( .A(n1043), .ZN(n1022) );
NOR3_X1 U754 ( .A1(n1008), .A2(G953), .A3(G952), .ZN(n1006) );
AND4_X1 U755 ( .A1(n1040), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1008) );
NOR4_X1 U756 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
XOR2_X1 U757 ( .A(n1051), .B(KEYINPUT36), .Z(n1050) );
NAND2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U760 ( .A1(KEYINPUT58), .A2(n1056), .ZN(n1054) );
NAND2_X1 U761 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U762 ( .A1(n1059), .A2(n1060), .ZN(n1052) );
NAND2_X1 U763 ( .A1(n1058), .A2(n1061), .ZN(n1060) );
NAND2_X1 U764 ( .A1(KEYINPUT58), .A2(n1062), .ZN(n1061) );
INV_X1 U765 ( .A(KEYINPUT51), .ZN(n1058) );
NOR2_X1 U766 ( .A1(n1063), .A2(n1064), .ZN(n1049) );
XNOR2_X1 U767 ( .A(G478), .B(KEYINPUT9), .ZN(n1064) );
INV_X1 U768 ( .A(n1065), .ZN(n1063) );
NOR2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(n1048) );
XOR2_X1 U770 ( .A(n1068), .B(KEYINPUT53), .Z(n1045) );
NAND2_X1 U771 ( .A1(n1067), .A2(n1066), .ZN(n1068) );
XOR2_X1 U772 ( .A(n1069), .B(KEYINPUT35), .Z(n1067) );
XNOR2_X1 U773 ( .A(KEYINPUT18), .B(n1070), .ZN(n1044) );
NOR2_X1 U774 ( .A1(n1027), .A2(n1030), .ZN(n1040) );
XOR2_X1 U775 ( .A(n1071), .B(n1072), .Z(G72) );
NOR2_X1 U776 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XOR2_X1 U777 ( .A(n1075), .B(n1076), .Z(n1074) );
XNOR2_X1 U778 ( .A(n1077), .B(n1078), .ZN(n1076) );
XNOR2_X1 U779 ( .A(n1079), .B(n1080), .ZN(n1075) );
NOR2_X1 U780 ( .A1(G131), .A2(KEYINPUT56), .ZN(n1080) );
NOR2_X1 U781 ( .A1(KEYINPUT11), .A2(n1081), .ZN(n1079) );
XOR2_X1 U782 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U783 ( .A1(G140), .A2(n1084), .ZN(n1083) );
XNOR2_X1 U784 ( .A(KEYINPUT34), .B(KEYINPUT3), .ZN(n1084) );
XNOR2_X1 U785 ( .A(G125), .B(KEYINPUT8), .ZN(n1082) );
NOR2_X1 U786 ( .A1(G900), .A2(n1085), .ZN(n1073) );
NAND2_X1 U787 ( .A1(n1086), .A2(n1087), .ZN(n1071) );
NAND2_X1 U788 ( .A1(n1088), .A2(n1085), .ZN(n1087) );
NAND3_X1 U789 ( .A1(KEYINPUT55), .A2(n1089), .A3(G953), .ZN(n1086) );
NAND2_X1 U790 ( .A1(G900), .A2(G227), .ZN(n1089) );
XOR2_X1 U791 ( .A(n1090), .B(n1091), .Z(G69) );
NOR2_X1 U792 ( .A1(n1092), .A2(n1085), .ZN(n1091) );
NOR2_X1 U793 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XNOR2_X1 U794 ( .A(G224), .B(KEYINPUT5), .ZN(n1093) );
NAND2_X1 U795 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
NAND2_X1 U796 ( .A1(n1097), .A2(n1085), .ZN(n1096) );
XNOR2_X1 U797 ( .A(n1098), .B(n1099), .ZN(n1097) );
NOR2_X1 U798 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND3_X1 U799 ( .A1(G898), .A2(n1098), .A3(G953), .ZN(n1095) );
NOR2_X1 U800 ( .A1(n1102), .A2(n1103), .ZN(G66) );
XOR2_X1 U801 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U802 ( .A1(n1106), .A2(n1059), .ZN(n1104) );
INV_X1 U803 ( .A(n1057), .ZN(n1059) );
NOR2_X1 U804 ( .A1(n1102), .A2(n1107), .ZN(G63) );
XOR2_X1 U805 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U806 ( .A1(n1106), .A2(G478), .ZN(n1109) );
NOR2_X1 U807 ( .A1(n1102), .A2(n1110), .ZN(G60) );
NOR3_X1 U808 ( .A1(n1069), .A2(n1111), .A3(n1112), .ZN(n1110) );
AND3_X1 U809 ( .A1(n1113), .A2(G475), .A3(n1106), .ZN(n1112) );
NOR2_X1 U810 ( .A1(n1114), .A2(n1113), .ZN(n1111) );
NOR2_X1 U811 ( .A1(n1011), .A2(n1066), .ZN(n1114) );
XNOR2_X1 U812 ( .A(G104), .B(n1115), .ZN(G6) );
NOR2_X1 U813 ( .A1(n1102), .A2(n1116), .ZN(G57) );
XOR2_X1 U814 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U815 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U816 ( .A(n1121), .B(n1122), .Z(n1117) );
XNOR2_X1 U817 ( .A(n1123), .B(n1124), .ZN(n1122) );
NAND2_X1 U818 ( .A1(KEYINPUT6), .A2(n1125), .ZN(n1124) );
NAND2_X1 U819 ( .A1(n1126), .A2(KEYINPUT29), .ZN(n1123) );
XNOR2_X1 U820 ( .A(n1127), .B(KEYINPUT22), .ZN(n1126) );
NAND2_X1 U821 ( .A1(n1106), .A2(G472), .ZN(n1121) );
NOR2_X1 U822 ( .A1(n1102), .A2(n1128), .ZN(G54) );
XOR2_X1 U823 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U824 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U825 ( .A(G110), .B(n1133), .Z(n1132) );
NOR2_X1 U826 ( .A1(KEYINPUT42), .A2(n1134), .ZN(n1133) );
XOR2_X1 U827 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U828 ( .A(n1137), .B(n1120), .Z(n1129) );
XOR2_X1 U829 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U830 ( .A1(G140), .A2(KEYINPUT0), .ZN(n1139) );
NAND2_X1 U831 ( .A1(n1106), .A2(G469), .ZN(n1138) );
NOR2_X1 U832 ( .A1(n1102), .A2(n1140), .ZN(G51) );
XOR2_X1 U833 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U834 ( .A1(KEYINPUT30), .A2(n1143), .ZN(n1142) );
NAND2_X1 U835 ( .A1(n1106), .A2(n1144), .ZN(n1141) );
NOR2_X1 U836 ( .A1(n1145), .A2(n1011), .ZN(n1106) );
NOR3_X1 U837 ( .A1(n1088), .A2(n1101), .A3(n1146), .ZN(n1011) );
XOR2_X1 U838 ( .A(n1100), .B(KEYINPUT45), .Z(n1146) );
NAND4_X1 U839 ( .A1(n1147), .A2(n1115), .A3(n1148), .A4(n1149), .ZN(n1101) );
AND3_X1 U840 ( .A1(n1150), .A2(n1005), .A3(n1151), .ZN(n1149) );
NAND3_X1 U841 ( .A1(n1152), .A2(n1153), .A3(n1037), .ZN(n1005) );
NAND2_X1 U842 ( .A1(n1154), .A2(n1037), .ZN(n1148) );
INV_X1 U843 ( .A(n1155), .ZN(n1154) );
NAND3_X1 U844 ( .A1(n1152), .A2(n1153), .A3(n1038), .ZN(n1115) );
NAND2_X1 U845 ( .A1(n1156), .A2(n1157), .ZN(n1147) );
NAND2_X1 U846 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U847 ( .A(n1160), .B(KEYINPUT57), .Z(n1158) );
NAND4_X1 U848 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1088) );
AND4_X1 U849 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NOR2_X1 U850 ( .A1(n1169), .A2(n1170), .ZN(n1163) );
NOR2_X1 U851 ( .A1(KEYINPUT13), .A2(n1171), .ZN(n1170) );
NAND4_X1 U852 ( .A1(n1172), .A2(n1042), .A3(KEYINPUT13), .A4(n1173), .ZN(n1162) );
NAND2_X1 U853 ( .A1(n1038), .A2(n1174), .ZN(n1161) );
NAND2_X1 U854 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND4_X1 U855 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NAND2_X1 U856 ( .A1(KEYINPUT14), .A2(n1181), .ZN(n1180) );
NAND2_X1 U857 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
INV_X1 U858 ( .A(KEYINPUT14), .ZN(n1183) );
NAND2_X1 U859 ( .A1(n1032), .A2(n1184), .ZN(n1182) );
NAND2_X1 U860 ( .A1(n1041), .A2(n1172), .ZN(n1175) );
NOR2_X1 U861 ( .A1(n1085), .A2(G952), .ZN(n1102) );
XNOR2_X1 U862 ( .A(G146), .B(n1185), .ZN(G48) );
NAND4_X1 U863 ( .A1(n1177), .A2(n1038), .A3(n1152), .A4(n1186), .ZN(n1185) );
XNOR2_X1 U864 ( .A(KEYINPUT31), .B(n1178), .ZN(n1186) );
XOR2_X1 U865 ( .A(G143), .B(n1169), .Z(G45) );
AND4_X1 U866 ( .A1(n1041), .A2(n1152), .A3(n1187), .A4(n1188), .ZN(n1169) );
AND2_X1 U867 ( .A1(n1189), .A2(n1178), .ZN(n1187) );
NAND2_X1 U868 ( .A1(n1190), .A2(n1191), .ZN(G42) );
NAND2_X1 U869 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U870 ( .A(n1171), .B(KEYINPUT21), .Z(n1193) );
XNOR2_X1 U871 ( .A(KEYINPUT43), .B(G140), .ZN(n1192) );
NAND2_X1 U872 ( .A1(n1194), .A2(n1195), .ZN(n1190) );
XNOR2_X1 U873 ( .A(KEYINPUT26), .B(n1171), .ZN(n1195) );
NAND3_X1 U874 ( .A1(n1042), .A2(n1038), .A3(n1172), .ZN(n1171) );
XNOR2_X1 U875 ( .A(KEYINPUT43), .B(n1196), .ZN(n1194) );
XNOR2_X1 U876 ( .A(G137), .B(n1168), .ZN(G39) );
NAND3_X1 U877 ( .A1(n1172), .A2(n1177), .A3(n1043), .ZN(n1168) );
XNOR2_X1 U878 ( .A(G134), .B(n1167), .ZN(G36) );
NAND3_X1 U879 ( .A1(n1172), .A2(n1037), .A3(n1041), .ZN(n1167) );
INV_X1 U880 ( .A(n1197), .ZN(n1172) );
XOR2_X1 U881 ( .A(G131), .B(n1198), .Z(G33) );
NOR4_X1 U882 ( .A1(KEYINPUT61), .A2(n1173), .A3(n1197), .A4(n1199), .ZN(n1198) );
INV_X1 U883 ( .A(n1041), .ZN(n1199) );
NAND3_X1 U884 ( .A1(n1032), .A2(n1178), .A3(n1200), .ZN(n1197) );
INV_X1 U885 ( .A(n1030), .ZN(n1200) );
NAND2_X1 U886 ( .A1(n1201), .A2(n1026), .ZN(n1030) );
INV_X1 U887 ( .A(n1028), .ZN(n1201) );
XNOR2_X1 U888 ( .A(G128), .B(n1202), .ZN(G30) );
NAND2_X1 U889 ( .A1(KEYINPUT12), .A2(n1203), .ZN(n1202) );
INV_X1 U890 ( .A(n1166), .ZN(n1203) );
NAND4_X1 U891 ( .A1(n1177), .A2(n1037), .A3(n1152), .A4(n1178), .ZN(n1166) );
XNOR2_X1 U892 ( .A(G101), .B(n1150), .ZN(G3) );
NAND3_X1 U893 ( .A1(n1041), .A2(n1152), .A3(n1204), .ZN(n1150) );
INV_X1 U894 ( .A(n1181), .ZN(n1152) );
NAND2_X1 U895 ( .A1(n1156), .A2(n1032), .ZN(n1181) );
XNOR2_X1 U896 ( .A(G125), .B(n1165), .ZN(G27) );
NAND4_X1 U897 ( .A1(n1042), .A2(n1038), .A3(n1024), .A4(n1178), .ZN(n1165) );
NAND2_X1 U898 ( .A1(n1013), .A2(n1205), .ZN(n1178) );
NAND2_X1 U899 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
INV_X1 U900 ( .A(G900), .ZN(n1207) );
INV_X1 U901 ( .A(n1173), .ZN(n1038) );
NAND2_X1 U902 ( .A1(n1208), .A2(n1209), .ZN(G24) );
NAND2_X1 U903 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
INV_X1 U904 ( .A(G122), .ZN(n1211) );
NAND2_X1 U905 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
NAND2_X1 U906 ( .A1(KEYINPUT63), .A2(n1151), .ZN(n1213) );
OR2_X1 U907 ( .A1(n1214), .A2(KEYINPUT63), .ZN(n1212) );
NAND2_X1 U908 ( .A1(G122), .A2(n1214), .ZN(n1208) );
NOR2_X1 U909 ( .A1(n1215), .A2(KEYINPUT47), .ZN(n1214) );
INV_X1 U910 ( .A(n1151), .ZN(n1215) );
NAND4_X1 U911 ( .A1(n1024), .A2(n1153), .A3(n1188), .A4(n1189), .ZN(n1151) );
AND3_X1 U912 ( .A1(n1216), .A2(n1217), .A3(n1070), .ZN(n1153) );
XNOR2_X1 U913 ( .A(G119), .B(n1218), .ZN(G21) );
NAND2_X1 U914 ( .A1(n1219), .A2(n1156), .ZN(n1218) );
INV_X1 U915 ( .A(n1184), .ZN(n1156) );
XOR2_X1 U916 ( .A(n1159), .B(KEYINPUT33), .Z(n1219) );
NAND3_X1 U917 ( .A1(n1177), .A2(n1220), .A3(n1204), .ZN(n1159) );
NOR2_X1 U918 ( .A1(n1216), .A2(n1070), .ZN(n1177) );
XNOR2_X1 U919 ( .A(n1221), .B(n1222), .ZN(G18) );
NOR2_X1 U920 ( .A1(n1155), .A2(n1223), .ZN(n1222) );
XOR2_X1 U921 ( .A(KEYINPUT52), .B(n1037), .Z(n1223) );
NOR2_X1 U922 ( .A1(n1188), .A2(n1224), .ZN(n1037) );
XOR2_X1 U923 ( .A(G113), .B(n1100), .Z(G15) );
NOR2_X1 U924 ( .A1(n1155), .A2(n1173), .ZN(n1100) );
NAND2_X1 U925 ( .A1(n1224), .A2(n1188), .ZN(n1173) );
NAND3_X1 U926 ( .A1(n1024), .A2(n1217), .A3(n1041), .ZN(n1155) );
NOR2_X1 U927 ( .A1(n1018), .A2(n1070), .ZN(n1041) );
INV_X1 U928 ( .A(n1016), .ZN(n1070) );
NOR2_X1 U929 ( .A1(n1027), .A2(n1184), .ZN(n1024) );
INV_X1 U930 ( .A(n1220), .ZN(n1027) );
NOR2_X1 U931 ( .A1(n1034), .A2(n1225), .ZN(n1220) );
INV_X1 U932 ( .A(n1033), .ZN(n1225) );
XOR2_X1 U933 ( .A(G110), .B(n1226), .Z(G12) );
NOR2_X1 U934 ( .A1(n1184), .A2(n1160), .ZN(n1226) );
NAND3_X1 U935 ( .A1(n1042), .A2(n1032), .A3(n1204), .ZN(n1160) );
AND2_X1 U936 ( .A1(n1043), .A2(n1217), .ZN(n1204) );
NAND2_X1 U937 ( .A1(n1013), .A2(n1227), .ZN(n1217) );
NAND2_X1 U938 ( .A1(n1206), .A2(n1094), .ZN(n1227) );
INV_X1 U939 ( .A(G898), .ZN(n1094) );
AND3_X1 U940 ( .A1(G953), .A2(n1228), .A3(n1229), .ZN(n1206) );
XNOR2_X1 U941 ( .A(G902), .B(KEYINPUT27), .ZN(n1229) );
NAND3_X1 U942 ( .A1(n1228), .A2(n1085), .A3(G952), .ZN(n1013) );
NAND2_X1 U943 ( .A1(G237), .A2(G234), .ZN(n1228) );
NOR2_X1 U944 ( .A1(n1189), .A2(n1188), .ZN(n1043) );
XNOR2_X1 U945 ( .A(n1069), .B(n1066), .ZN(n1188) );
INV_X1 U946 ( .A(G475), .ZN(n1066) );
NOR2_X1 U947 ( .A1(n1113), .A2(G902), .ZN(n1069) );
XNOR2_X1 U948 ( .A(n1230), .B(n1231), .ZN(n1113) );
XOR2_X1 U949 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U950 ( .A(G143), .B(G131), .Z(n1233) );
XNOR2_X1 U951 ( .A(KEYINPUT60), .B(n1234), .ZN(n1232) );
INV_X1 U952 ( .A(G146), .ZN(n1234) );
XOR2_X1 U953 ( .A(n1235), .B(n1236), .Z(n1230) );
XNOR2_X1 U954 ( .A(n1237), .B(n1238), .ZN(n1236) );
NOR2_X1 U955 ( .A1(KEYINPUT19), .A2(n1239), .ZN(n1238) );
XOR2_X1 U956 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U957 ( .A(G113), .B(KEYINPUT17), .ZN(n1240) );
XOR2_X1 U958 ( .A(n1242), .B(n1243), .Z(n1235) );
AND2_X1 U959 ( .A1(n1244), .A2(G214), .ZN(n1243) );
NAND2_X1 U960 ( .A1(KEYINPUT16), .A2(n1196), .ZN(n1242) );
INV_X1 U961 ( .A(n1224), .ZN(n1189) );
NOR2_X1 U962 ( .A1(n1245), .A2(n1047), .ZN(n1224) );
NOR2_X1 U963 ( .A1(n1065), .A2(G478), .ZN(n1047) );
AND2_X1 U964 ( .A1(G478), .A2(n1065), .ZN(n1245) );
NAND2_X1 U965 ( .A1(n1108), .A2(n1145), .ZN(n1065) );
NAND2_X1 U966 ( .A1(n1246), .A2(n1247), .ZN(n1108) );
NAND4_X1 U967 ( .A1(G234), .A2(G217), .A3(n1248), .A4(n1085), .ZN(n1247) );
XOR2_X1 U968 ( .A(n1249), .B(KEYINPUT15), .Z(n1246) );
NAND2_X1 U969 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND3_X1 U970 ( .A1(G217), .A2(n1085), .A3(G234), .ZN(n1251) );
XNOR2_X1 U971 ( .A(KEYINPUT62), .B(n1248), .ZN(n1250) );
NAND3_X1 U972 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1248) );
OR2_X1 U973 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NAND3_X1 U974 ( .A1(n1257), .A2(n1255), .A3(n1258), .ZN(n1253) );
INV_X1 U975 ( .A(KEYINPUT54), .ZN(n1255) );
OR2_X1 U976 ( .A1(n1258), .A2(n1257), .ZN(n1252) );
AND2_X1 U977 ( .A1(KEYINPUT2), .A2(n1256), .ZN(n1257) );
NAND2_X1 U978 ( .A1(n1259), .A2(n1260), .ZN(n1256) );
NAND2_X1 U979 ( .A1(n1261), .A2(G107), .ZN(n1260) );
XOR2_X1 U980 ( .A(KEYINPUT40), .B(n1262), .Z(n1259) );
NOR2_X1 U981 ( .A1(G107), .A2(n1261), .ZN(n1262) );
XNOR2_X1 U982 ( .A(G116), .B(n1263), .ZN(n1261) );
NOR2_X1 U983 ( .A1(G122), .A2(KEYINPUT38), .ZN(n1263) );
XOR2_X1 U984 ( .A(n1264), .B(n1265), .Z(n1258) );
XOR2_X1 U985 ( .A(KEYINPUT41), .B(n1266), .Z(n1265) );
AND2_X1 U986 ( .A1(n1267), .A2(n1034), .ZN(n1032) );
XNOR2_X1 U987 ( .A(n1268), .B(G469), .ZN(n1034) );
NAND2_X1 U988 ( .A1(n1269), .A2(n1145), .ZN(n1268) );
XOR2_X1 U989 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U990 ( .A(n1136), .B(n1272), .ZN(n1271) );
XOR2_X1 U991 ( .A(n1273), .B(n1274), .Z(n1136) );
INV_X1 U992 ( .A(n1077), .ZN(n1274) );
XNOR2_X1 U993 ( .A(n1275), .B(KEYINPUT46), .ZN(n1077) );
NAND2_X1 U994 ( .A1(KEYINPUT49), .A2(n1276), .ZN(n1273) );
XNOR2_X1 U995 ( .A(n1120), .B(n1277), .ZN(n1270) );
XNOR2_X1 U996 ( .A(G140), .B(n1278), .ZN(n1277) );
NAND2_X1 U997 ( .A1(KEYINPUT25), .A2(n1131), .ZN(n1278) );
AND2_X1 U998 ( .A1(G227), .A2(n1085), .ZN(n1131) );
XNOR2_X1 U999 ( .A(KEYINPUT23), .B(n1033), .ZN(n1267) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1279), .ZN(n1033) );
NOR2_X1 U1001 ( .A1(n1016), .A2(n1216), .ZN(n1042) );
INV_X1 U1002 ( .A(n1018), .ZN(n1216) );
XNOR2_X1 U1003 ( .A(n1062), .B(n1057), .ZN(n1018) );
NAND2_X1 U1004 ( .A1(G217), .A2(n1279), .ZN(n1057) );
NAND2_X1 U1005 ( .A1(n1280), .A2(G234), .ZN(n1279) );
INV_X1 U1006 ( .A(n1055), .ZN(n1062) );
NAND2_X1 U1007 ( .A1(n1105), .A2(n1145), .ZN(n1055) );
XOR2_X1 U1008 ( .A(n1281), .B(n1282), .Z(n1105) );
XOR2_X1 U1009 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U1010 ( .A(n1285), .B(n1286), .ZN(n1284) );
NOR2_X1 U1011 ( .A1(KEYINPUT32), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U1012 ( .A(G110), .B(n1288), .ZN(n1287) );
NAND2_X1 U1013 ( .A1(n1289), .A2(KEYINPUT7), .ZN(n1288) );
XNOR2_X1 U1014 ( .A(G128), .B(G119), .ZN(n1289) );
NAND2_X1 U1015 ( .A1(n1290), .A2(KEYINPUT20), .ZN(n1285) );
XNOR2_X1 U1016 ( .A(G146), .B(KEYINPUT39), .ZN(n1290) );
AND3_X1 U1017 ( .A1(G221), .A2(n1085), .A3(G234), .ZN(n1283) );
XOR2_X1 U1018 ( .A(n1291), .B(n1292), .Z(n1281) );
XNOR2_X1 U1019 ( .A(KEYINPUT59), .B(n1196), .ZN(n1292) );
INV_X1 U1020 ( .A(G140), .ZN(n1196) );
XNOR2_X1 U1021 ( .A(G137), .B(G125), .ZN(n1291) );
XNOR2_X1 U1022 ( .A(n1293), .B(G472), .ZN(n1016) );
NAND2_X1 U1023 ( .A1(n1294), .A2(n1145), .ZN(n1293) );
XOR2_X1 U1024 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1025 ( .A(n1125), .B(n1120), .ZN(n1296) );
XNOR2_X1 U1026 ( .A(n1297), .B(n1078), .ZN(n1120) );
XOR2_X1 U1027 ( .A(G137), .B(n1266), .Z(n1078) );
XOR2_X1 U1028 ( .A(G134), .B(KEYINPUT10), .Z(n1266) );
XNOR2_X1 U1029 ( .A(G131), .B(KEYINPUT37), .ZN(n1297) );
XOR2_X1 U1030 ( .A(n1298), .B(n1119), .Z(n1295) );
XNOR2_X1 U1031 ( .A(n1299), .B(G101), .ZN(n1119) );
NAND2_X1 U1032 ( .A1(G210), .A2(n1244), .ZN(n1299) );
NOR2_X1 U1033 ( .A1(G953), .A2(G237), .ZN(n1244) );
NAND2_X1 U1034 ( .A1(KEYINPUT4), .A2(n1127), .ZN(n1298) );
XNOR2_X1 U1035 ( .A(n1300), .B(n1301), .ZN(n1127) );
XNOR2_X1 U1036 ( .A(n1302), .B(n1303), .ZN(n1301) );
NOR2_X1 U1037 ( .A1(G116), .A2(KEYINPUT28), .ZN(n1303) );
INV_X1 U1038 ( .A(G119), .ZN(n1302) );
NAND2_X1 U1039 ( .A1(n1028), .A2(n1026), .ZN(n1184) );
NAND2_X1 U1040 ( .A1(G214), .A2(n1304), .ZN(n1026) );
XNOR2_X1 U1041 ( .A(n1305), .B(n1144), .ZN(n1028) );
AND2_X1 U1042 ( .A1(G210), .A2(n1304), .ZN(n1144) );
NAND2_X1 U1043 ( .A1(n1280), .A2(n1306), .ZN(n1304) );
INV_X1 U1044 ( .A(G237), .ZN(n1306) );
XNOR2_X1 U1045 ( .A(G902), .B(KEYINPUT24), .ZN(n1280) );
NAND2_X1 U1046 ( .A1(n1307), .A2(n1145), .ZN(n1305) );
INV_X1 U1047 ( .A(G902), .ZN(n1145) );
XNOR2_X1 U1048 ( .A(n1143), .B(KEYINPUT1), .ZN(n1307) );
XNOR2_X1 U1049 ( .A(n1308), .B(n1309), .ZN(n1143) );
XNOR2_X1 U1050 ( .A(n1237), .B(n1310), .ZN(n1309) );
AND2_X1 U1051 ( .A1(n1085), .A2(G224), .ZN(n1310) );
INV_X1 U1052 ( .A(G953), .ZN(n1085) );
INV_X1 U1053 ( .A(G125), .ZN(n1237) );
XNOR2_X1 U1054 ( .A(n1098), .B(n1125), .ZN(n1308) );
XNOR2_X1 U1055 ( .A(n1275), .B(KEYINPUT44), .ZN(n1125) );
XNOR2_X1 U1056 ( .A(G146), .B(n1264), .ZN(n1275) );
XOR2_X1 U1057 ( .A(G128), .B(G143), .Z(n1264) );
XNOR2_X1 U1058 ( .A(n1311), .B(n1312), .ZN(n1098) );
XOR2_X1 U1059 ( .A(n1313), .B(n1300), .Z(n1312) );
XNOR2_X1 U1060 ( .A(G113), .B(KEYINPUT48), .ZN(n1300) );
NAND2_X1 U1061 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND2_X1 U1062 ( .A1(G119), .A2(n1221), .ZN(n1315) );
XOR2_X1 U1063 ( .A(KEYINPUT50), .B(n1316), .Z(n1314) );
NOR2_X1 U1064 ( .A1(G119), .A2(n1221), .ZN(n1316) );
INV_X1 U1065 ( .A(G116), .ZN(n1221) );
XNOR2_X1 U1066 ( .A(n1272), .B(n1241), .ZN(n1311) );
XNOR2_X1 U1067 ( .A(n1276), .B(G122), .ZN(n1241) );
INV_X1 U1068 ( .A(G104), .ZN(n1276) );
XOR2_X1 U1069 ( .A(G110), .B(n1135), .Z(n1272) );
XOR2_X1 U1070 ( .A(G101), .B(G107), .Z(n1135) );
endmodule


