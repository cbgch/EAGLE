//Key = 1010011001110011111100011001010001010000000100111101010101100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;

XNOR2_X1 U731 ( .A(G107), .B(n1016), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR3_X1 U733 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND3_X1 U734 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1019) );
NAND2_X1 U735 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U736 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NAND3_X1 U737 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NAND2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
OR2_X1 U740 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U741 ( .A1(n1038), .A2(n1039), .ZN(n1032) );
NAND2_X1 U742 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U744 ( .A1(n1034), .A2(n1044), .A3(n1038), .ZN(n1027) );
NAND2_X1 U745 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U746 ( .A1(n1031), .A2(n1047), .ZN(n1046) );
NAND2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U748 ( .A1(n1029), .A2(n1050), .ZN(n1045) );
NAND2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR3_X1 U751 ( .A1(n1055), .A2(G953), .A3(n1056), .ZN(n1017) );
INV_X1 U752 ( .A(n1022), .ZN(n1056) );
NAND4_X1 U753 ( .A1(n1031), .A2(n1034), .A3(n1057), .A4(n1058), .ZN(n1022) );
NOR4_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
XOR2_X1 U755 ( .A(n1063), .B(n1064), .Z(n1061) );
NOR2_X1 U756 ( .A1(G475), .A2(KEYINPUT62), .ZN(n1064) );
AND2_X1 U757 ( .A1(n1065), .A2(G478), .ZN(n1060) );
XNOR2_X1 U758 ( .A(n1066), .B(n1067), .ZN(n1057) );
XNOR2_X1 U759 ( .A(KEYINPUT26), .B(n1020), .ZN(n1055) );
XOR2_X1 U760 ( .A(n1068), .B(n1069), .Z(G72) );
NOR2_X1 U761 ( .A1(n1070), .A2(n1023), .ZN(n1069) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1068) );
NAND3_X1 U764 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
INV_X1 U765 ( .A(n1078), .ZN(n1077) );
NAND2_X1 U766 ( .A1(G953), .A2(n1072), .ZN(n1076) );
NAND2_X1 U767 ( .A1(n1079), .A2(n1023), .ZN(n1075) );
XOR2_X1 U768 ( .A(n1080), .B(KEYINPUT44), .Z(n1073) );
NAND3_X1 U769 ( .A1(n1079), .A2(n1023), .A3(n1078), .ZN(n1080) );
XOR2_X1 U770 ( .A(n1081), .B(n1082), .Z(n1078) );
XOR2_X1 U771 ( .A(n1083), .B(n1084), .Z(n1081) );
NOR2_X1 U772 ( .A1(KEYINPUT54), .A2(n1085), .ZN(n1084) );
XOR2_X1 U773 ( .A(n1086), .B(n1087), .Z(n1085) );
XNOR2_X1 U774 ( .A(KEYINPUT1), .B(n1088), .ZN(n1086) );
NOR2_X1 U775 ( .A1(KEYINPUT40), .A2(n1089), .ZN(n1088) );
NAND3_X1 U776 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1083) );
NAND2_X1 U777 ( .A1(KEYINPUT25), .A2(n1093), .ZN(n1091) );
NAND2_X1 U778 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XNOR2_X1 U779 ( .A(KEYINPUT20), .B(n1096), .ZN(n1094) );
NAND2_X1 U780 ( .A1(n1097), .A2(n1098), .ZN(n1090) );
INV_X1 U781 ( .A(KEYINPUT25), .ZN(n1098) );
NAND2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NAND2_X1 U783 ( .A1(KEYINPUT20), .A2(n1096), .ZN(n1100) );
OR3_X1 U784 ( .A1(n1101), .A2(KEYINPUT20), .A3(n1096), .ZN(n1099) );
NAND2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1079) );
XOR2_X1 U786 ( .A(n1104), .B(KEYINPUT37), .Z(n1103) );
XOR2_X1 U787 ( .A(n1105), .B(n1106), .Z(G69) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U789 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U790 ( .A1(n1111), .A2(G953), .ZN(n1110) );
XOR2_X1 U791 ( .A(n1112), .B(n1113), .Z(n1109) );
XNOR2_X1 U792 ( .A(n1114), .B(n1115), .ZN(n1113) );
NAND2_X1 U793 ( .A1(KEYINPUT53), .A2(n1116), .ZN(n1114) );
XOR2_X1 U794 ( .A(KEYINPUT21), .B(n1117), .Z(n1116) );
NAND2_X1 U795 ( .A1(G953), .A2(n1118), .ZN(n1107) );
NAND2_X1 U796 ( .A1(G224), .A2(n1119), .ZN(n1118) );
XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n1120), .ZN(n1119) );
INV_X1 U798 ( .A(G898), .ZN(n1120) );
NOR2_X1 U799 ( .A1(n1121), .A2(G953), .ZN(n1105) );
NOR2_X1 U800 ( .A1(n1122), .A2(n1123), .ZN(G66) );
XNOR2_X1 U801 ( .A(n1124), .B(n1125), .ZN(n1123) );
NOR2_X1 U802 ( .A1(n1067), .A2(n1126), .ZN(n1124) );
NOR2_X1 U803 ( .A1(n1122), .A2(n1127), .ZN(G63) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U805 ( .A1(KEYINPUT31), .A2(n1130), .ZN(n1129) );
AND2_X1 U806 ( .A1(G478), .A2(n1131), .ZN(n1128) );
NOR2_X1 U807 ( .A1(n1122), .A2(n1132), .ZN(G60) );
XOR2_X1 U808 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR3_X1 U809 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
NOR2_X1 U810 ( .A1(KEYINPUT27), .A2(n1138), .ZN(n1137) );
AND2_X1 U811 ( .A1(n1139), .A2(n1021), .ZN(n1138) );
AND2_X1 U812 ( .A1(n1126), .A2(KEYINPUT27), .ZN(n1136) );
NAND2_X1 U813 ( .A1(KEYINPUT2), .A2(n1140), .ZN(n1133) );
XNOR2_X1 U814 ( .A(G104), .B(n1141), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1122), .A2(n1142), .ZN(G57) );
XOR2_X1 U816 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U817 ( .A(KEYINPUT3), .B(n1145), .Z(n1144) );
AND2_X1 U818 ( .A1(G472), .A2(n1131), .ZN(n1145) );
NOR2_X1 U819 ( .A1(n1122), .A2(n1146), .ZN(G54) );
XOR2_X1 U820 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U821 ( .A(n1149), .B(n1150), .ZN(n1148) );
NAND3_X1 U822 ( .A1(G469), .A2(n1021), .A3(n1151), .ZN(n1149) );
XNOR2_X1 U823 ( .A(G902), .B(KEYINPUT16), .ZN(n1151) );
XOR2_X1 U824 ( .A(n1152), .B(n1153), .Z(n1147) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U826 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NAND2_X1 U827 ( .A1(n1158), .A2(n1095), .ZN(n1157) );
XOR2_X1 U828 ( .A(KEYINPUT24), .B(n1159), .Z(n1156) );
NOR2_X1 U829 ( .A1(n1095), .A2(n1158), .ZN(n1159) );
XNOR2_X1 U830 ( .A(KEYINPUT22), .B(n1160), .ZN(n1158) );
NAND2_X1 U831 ( .A1(KEYINPUT51), .A2(n1161), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1122), .A2(n1162), .ZN(G51) );
NOR3_X1 U833 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
NOR2_X1 U834 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
INV_X1 U835 ( .A(n1168), .ZN(n1167) );
NOR2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
XNOR2_X1 U837 ( .A(KEYINPUT17), .B(n1171), .ZN(n1170) );
NOR3_X1 U838 ( .A1(n1168), .A2(n1171), .A3(n1169), .ZN(n1164) );
XOR2_X1 U839 ( .A(n1172), .B(n1173), .Z(n1168) );
XOR2_X1 U840 ( .A(n1174), .B(n1175), .Z(n1172) );
AND2_X1 U841 ( .A1(n1169), .A2(n1171), .ZN(n1163) );
NAND2_X1 U842 ( .A1(n1131), .A2(n1176), .ZN(n1171) );
INV_X1 U843 ( .A(n1126), .ZN(n1131) );
NAND2_X1 U844 ( .A1(G902), .A2(n1021), .ZN(n1126) );
NAND3_X1 U845 ( .A1(n1121), .A2(n1102), .A3(n1104), .ZN(n1021) );
AND4_X1 U846 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1104) );
AND4_X1 U847 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1102) );
OR2_X1 U848 ( .A1(n1185), .A2(n1040), .ZN(n1182) );
AND4_X1 U849 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1121) );
NOR4_X1 U850 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
INV_X1 U851 ( .A(n1141), .ZN(n1192) );
NAND3_X1 U852 ( .A1(n1029), .A2(n1194), .A3(n1036), .ZN(n1141) );
AND2_X1 U853 ( .A1(n1016), .A2(n1195), .ZN(n1188) );
NAND3_X1 U854 ( .A1(n1029), .A2(n1194), .A3(n1037), .ZN(n1016) );
NAND3_X1 U855 ( .A1(n1036), .A2(n1196), .A3(n1197), .ZN(n1186) );
XNOR2_X1 U856 ( .A(KEYINPUT42), .B(n1049), .ZN(n1196) );
INV_X1 U857 ( .A(KEYINPUT15), .ZN(n1169) );
NOR2_X1 U858 ( .A1(n1023), .A2(G952), .ZN(n1122) );
XNOR2_X1 U859 ( .A(G146), .B(n1177), .ZN(G48) );
NAND3_X1 U860 ( .A1(n1198), .A2(n1199), .A3(n1036), .ZN(n1177) );
XNOR2_X1 U861 ( .A(G143), .B(n1178), .ZN(G45) );
NAND4_X1 U862 ( .A1(n1200), .A2(n1199), .A3(n1201), .A4(n1202), .ZN(n1178) );
NOR3_X1 U863 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
XNOR2_X1 U864 ( .A(G140), .B(n1179), .ZN(G42) );
NAND3_X1 U865 ( .A1(n1031), .A2(n1200), .A3(n1206), .ZN(n1179) );
XNOR2_X1 U866 ( .A(G137), .B(n1180), .ZN(G39) );
NAND3_X1 U867 ( .A1(n1198), .A2(n1031), .A3(n1038), .ZN(n1180) );
XOR2_X1 U868 ( .A(G134), .B(n1207), .Z(G36) );
NOR2_X1 U869 ( .A1(n1185), .A2(n1208), .ZN(n1207) );
XNOR2_X1 U870 ( .A(KEYINPUT48), .B(n1040), .ZN(n1208) );
NAND4_X1 U871 ( .A1(n1201), .A2(n1031), .A3(n1037), .A4(n1209), .ZN(n1185) );
XNOR2_X1 U872 ( .A(G131), .B(n1184), .ZN(G33) );
NAND4_X1 U873 ( .A1(n1201), .A2(n1036), .A3(n1210), .A4(n1031), .ZN(n1184) );
NOR2_X1 U874 ( .A1(n1211), .A2(n1053), .ZN(n1031) );
NOR2_X1 U875 ( .A1(n1203), .A2(n1040), .ZN(n1210) );
XOR2_X1 U876 ( .A(G128), .B(n1212), .Z(G30) );
NOR2_X1 U877 ( .A1(KEYINPUT7), .A2(n1183), .ZN(n1212) );
NAND3_X1 U878 ( .A1(n1037), .A2(n1199), .A3(n1198), .ZN(n1183) );
AND3_X1 U879 ( .A1(n1200), .A2(n1209), .A3(n1213), .ZN(n1198) );
XOR2_X1 U880 ( .A(G101), .B(n1191), .Z(G3) );
AND3_X1 U881 ( .A1(n1038), .A2(n1194), .A3(n1201), .ZN(n1191) );
XOR2_X1 U882 ( .A(n1214), .B(n1215), .Z(G27) );
NOR2_X1 U883 ( .A1(KEYINPUT34), .A2(n1096), .ZN(n1215) );
NAND2_X1 U884 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
OR2_X1 U885 ( .A1(n1181), .A2(KEYINPUT39), .ZN(n1217) );
NAND3_X1 U886 ( .A1(n1034), .A2(n1199), .A3(n1206), .ZN(n1181) );
AND3_X1 U887 ( .A1(n1218), .A2(n1209), .A3(n1036), .ZN(n1206) );
NAND4_X1 U888 ( .A1(n1203), .A2(n1036), .A3(n1219), .A4(KEYINPUT39), .ZN(n1216) );
NOR3_X1 U889 ( .A1(n1048), .A2(n1051), .A3(n1220), .ZN(n1219) );
INV_X1 U890 ( .A(n1199), .ZN(n1051) );
INV_X1 U891 ( .A(n1218), .ZN(n1048) );
INV_X1 U892 ( .A(n1209), .ZN(n1203) );
NAND2_X1 U893 ( .A1(n1221), .A2(n1222), .ZN(n1209) );
NAND3_X1 U894 ( .A1(n1026), .A2(n1023), .A3(G952), .ZN(n1222) );
XOR2_X1 U895 ( .A(KEYINPUT33), .B(n1223), .Z(n1221) );
AND4_X1 U896 ( .A1(n1072), .A2(n1026), .A3(G902), .A4(G953), .ZN(n1223) );
INV_X1 U897 ( .A(G900), .ZN(n1072) );
XNOR2_X1 U898 ( .A(G122), .B(n1187), .ZN(G24) );
NAND4_X1 U899 ( .A1(n1197), .A2(n1029), .A3(n1224), .A4(n1225), .ZN(n1187) );
NOR2_X1 U900 ( .A1(n1062), .A2(n1226), .ZN(n1029) );
NAND2_X1 U901 ( .A1(n1227), .A2(n1228), .ZN(G21) );
NAND2_X1 U902 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
XOR2_X1 U903 ( .A(KEYINPUT19), .B(n1231), .Z(n1227) );
NOR2_X1 U904 ( .A1(n1229), .A2(n1230), .ZN(n1231) );
XNOR2_X1 U905 ( .A(KEYINPUT35), .B(n1232), .ZN(n1230) );
NAND2_X1 U906 ( .A1(n1233), .A2(n1234), .ZN(n1229) );
NAND2_X1 U907 ( .A1(n1193), .A2(n1235), .ZN(n1234) );
INV_X1 U908 ( .A(KEYINPUT36), .ZN(n1235) );
AND3_X1 U909 ( .A1(n1038), .A2(n1213), .A3(n1197), .ZN(n1193) );
NAND4_X1 U910 ( .A1(n1213), .A2(n1236), .A3(n1197), .A4(KEYINPUT36), .ZN(n1233) );
INV_X1 U911 ( .A(n1038), .ZN(n1236) );
AND2_X1 U912 ( .A1(n1226), .A2(n1062), .ZN(n1213) );
INV_X1 U913 ( .A(n1237), .ZN(n1226) );
XOR2_X1 U914 ( .A(n1190), .B(n1238), .Z(G18) );
NOR2_X1 U915 ( .A1(KEYINPUT63), .A2(n1239), .ZN(n1238) );
AND3_X1 U916 ( .A1(n1201), .A2(n1037), .A3(n1197), .ZN(n1190) );
NOR2_X1 U917 ( .A1(n1220), .A2(n1240), .ZN(n1197) );
NOR2_X1 U918 ( .A1(n1224), .A2(n1204), .ZN(n1037) );
INV_X1 U919 ( .A(n1225), .ZN(n1204) );
XNOR2_X1 U920 ( .A(G113), .B(n1241), .ZN(G15) );
NAND4_X1 U921 ( .A1(n1242), .A2(n1201), .A3(n1243), .A4(n1036), .ZN(n1241) );
NOR2_X1 U922 ( .A1(n1225), .A2(n1205), .ZN(n1036) );
INV_X1 U923 ( .A(n1224), .ZN(n1205) );
NOR2_X1 U924 ( .A1(KEYINPUT32), .A2(n1240), .ZN(n1243) );
INV_X1 U925 ( .A(n1049), .ZN(n1201) );
NAND2_X1 U926 ( .A1(n1062), .A2(n1237), .ZN(n1049) );
XNOR2_X1 U927 ( .A(n1034), .B(KEYINPUT46), .ZN(n1242) );
INV_X1 U928 ( .A(n1220), .ZN(n1034) );
NAND2_X1 U929 ( .A1(n1043), .A2(n1244), .ZN(n1220) );
XNOR2_X1 U930 ( .A(G110), .B(n1195), .ZN(G12) );
NAND3_X1 U931 ( .A1(n1038), .A2(n1194), .A3(n1218), .ZN(n1195) );
NOR2_X1 U932 ( .A1(n1237), .A2(n1062), .ZN(n1218) );
XNOR2_X1 U933 ( .A(n1245), .B(G472), .ZN(n1062) );
OR2_X1 U934 ( .A1(n1143), .A2(G902), .ZN(n1245) );
XNOR2_X1 U935 ( .A(n1246), .B(n1247), .ZN(n1143) );
XOR2_X1 U936 ( .A(n1248), .B(n1249), .Z(n1247) );
XOR2_X1 U937 ( .A(G113), .B(G101), .Z(n1249) );
XNOR2_X1 U938 ( .A(n1232), .B(G116), .ZN(n1248) );
XOR2_X1 U939 ( .A(n1250), .B(n1161), .Z(n1246) );
XOR2_X1 U940 ( .A(n1251), .B(n1252), .Z(n1250) );
NAND2_X1 U941 ( .A1(G210), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U942 ( .A(n1066), .B(n1254), .ZN(n1237) );
NOR2_X1 U943 ( .A1(n1255), .A2(KEYINPUT13), .ZN(n1254) );
INV_X1 U944 ( .A(n1067), .ZN(n1255) );
NAND2_X1 U945 ( .A1(G217), .A2(n1256), .ZN(n1067) );
NAND2_X1 U946 ( .A1(n1257), .A2(n1125), .ZN(n1066) );
XOR2_X1 U947 ( .A(n1258), .B(n1259), .Z(n1125) );
XNOR2_X1 U948 ( .A(n1096), .B(n1260), .ZN(n1259) );
XNOR2_X1 U949 ( .A(KEYINPUT8), .B(n1261), .ZN(n1260) );
INV_X1 U950 ( .A(G146), .ZN(n1261) );
XNOR2_X1 U951 ( .A(n1262), .B(n1101), .ZN(n1258) );
NAND2_X1 U952 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NAND2_X1 U953 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
INV_X1 U954 ( .A(n1267), .ZN(n1266) );
XOR2_X1 U955 ( .A(KEYINPUT52), .B(n1268), .Z(n1265) );
NAND2_X1 U956 ( .A1(n1269), .A2(n1267), .ZN(n1263) );
XOR2_X1 U957 ( .A(n1270), .B(n1271), .Z(n1267) );
INV_X1 U958 ( .A(G137), .ZN(n1271) );
NAND2_X1 U959 ( .A1(G221), .A2(n1272), .ZN(n1270) );
XOR2_X1 U960 ( .A(KEYINPUT10), .B(n1268), .Z(n1269) );
AND2_X1 U961 ( .A1(KEYINPUT14), .A2(n1273), .ZN(n1268) );
XOR2_X1 U962 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U963 ( .A(G110), .B(G128), .ZN(n1275) );
NAND2_X1 U964 ( .A1(KEYINPUT18), .A2(n1232), .ZN(n1274) );
INV_X1 U965 ( .A(G119), .ZN(n1232) );
XNOR2_X1 U966 ( .A(KEYINPUT6), .B(n1139), .ZN(n1257) );
NOR2_X1 U967 ( .A1(n1040), .A2(n1240), .ZN(n1194) );
NAND4_X1 U968 ( .A1(n1199), .A2(n1026), .A3(n1276), .A4(n1277), .ZN(n1240) );
NAND2_X1 U969 ( .A1(n1020), .A2(n1023), .ZN(n1277) );
INV_X1 U970 ( .A(G952), .ZN(n1020) );
NAND2_X1 U971 ( .A1(G953), .A2(n1278), .ZN(n1276) );
NAND2_X1 U972 ( .A1(n1111), .A2(G902), .ZN(n1278) );
XNOR2_X1 U973 ( .A(G898), .B(KEYINPUT60), .ZN(n1111) );
NAND2_X1 U974 ( .A1(G237), .A2(G234), .ZN(n1026) );
NOR2_X1 U975 ( .A1(n1054), .A2(n1053), .ZN(n1199) );
AND2_X1 U976 ( .A1(G214), .A2(n1279), .ZN(n1053) );
INV_X1 U977 ( .A(n1211), .ZN(n1054) );
XNOR2_X1 U978 ( .A(n1280), .B(n1176), .ZN(n1211) );
AND2_X1 U979 ( .A1(G210), .A2(n1279), .ZN(n1176) );
OR2_X1 U980 ( .A1(G902), .A2(G237), .ZN(n1279) );
NAND2_X1 U981 ( .A1(n1281), .A2(n1139), .ZN(n1280) );
XOR2_X1 U982 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U983 ( .A(n1284), .B(n1175), .Z(n1283) );
AND2_X1 U984 ( .A1(G224), .A2(n1023), .ZN(n1175) );
NAND2_X1 U985 ( .A1(KEYINPUT57), .A2(n1174), .ZN(n1284) );
XNOR2_X1 U986 ( .A(G125), .B(n1252), .ZN(n1174) );
XNOR2_X1 U987 ( .A(n1285), .B(n1286), .ZN(n1252) );
NOR2_X1 U988 ( .A1(KEYINPUT28), .A2(G143), .ZN(n1286) );
XNOR2_X1 U989 ( .A(G146), .B(G128), .ZN(n1285) );
NAND2_X1 U990 ( .A1(KEYINPUT58), .A2(n1173), .ZN(n1282) );
XOR2_X1 U991 ( .A(n1287), .B(n1115), .Z(n1173) );
XOR2_X1 U992 ( .A(G122), .B(G110), .Z(n1115) );
NAND2_X1 U993 ( .A1(n1288), .A2(KEYINPUT23), .ZN(n1287) );
XOR2_X1 U994 ( .A(n1112), .B(n1117), .Z(n1288) );
XNOR2_X1 U995 ( .A(G113), .B(n1289), .ZN(n1112) );
NOR2_X1 U996 ( .A1(KEYINPUT38), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U997 ( .A(n1239), .B(n1291), .ZN(n1290) );
NOR2_X1 U998 ( .A1(G119), .A2(KEYINPUT50), .ZN(n1291) );
INV_X1 U999 ( .A(G116), .ZN(n1239) );
INV_X1 U1000 ( .A(n1200), .ZN(n1040) );
NOR2_X1 U1001 ( .A1(n1043), .A2(n1042), .ZN(n1200) );
INV_X1 U1002 ( .A(n1244), .ZN(n1042) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1256), .ZN(n1244) );
NAND2_X1 U1004 ( .A1(G234), .A2(n1139), .ZN(n1256) );
XOR2_X1 U1005 ( .A(n1292), .B(G469), .Z(n1043) );
NAND2_X1 U1006 ( .A1(n1293), .A2(n1139), .ZN(n1292) );
XOR2_X1 U1007 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U1008 ( .A(n1296), .B(n1155), .Z(n1295) );
NOR2_X1 U1009 ( .A1(n1071), .A2(G953), .ZN(n1155) );
INV_X1 U1010 ( .A(G227), .ZN(n1071) );
NAND2_X1 U1011 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
NAND2_X1 U1012 ( .A1(n1101), .A2(n1160), .ZN(n1298) );
XOR2_X1 U1013 ( .A(KEYINPUT9), .B(n1299), .Z(n1297) );
NOR2_X1 U1014 ( .A1(n1101), .A2(n1160), .ZN(n1299) );
INV_X1 U1015 ( .A(G110), .ZN(n1160) );
NAND3_X1 U1016 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1294) );
NAND2_X1 U1017 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
INV_X1 U1018 ( .A(n1150), .ZN(n1303) );
OR3_X1 U1019 ( .A1(n1304), .A2(n1305), .A3(n1161), .ZN(n1301) );
INV_X1 U1020 ( .A(KEYINPUT0), .ZN(n1304) );
NAND2_X1 U1021 ( .A1(n1161), .A2(n1305), .ZN(n1300) );
NAND2_X1 U1022 ( .A1(KEYINPUT47), .A2(n1150), .ZN(n1305) );
XNOR2_X1 U1023 ( .A(n1306), .B(n1307), .ZN(n1150) );
XOR2_X1 U1024 ( .A(KEYINPUT45), .B(KEYINPUT29), .Z(n1307) );
XOR2_X1 U1025 ( .A(n1082), .B(n1117), .Z(n1306) );
XNOR2_X1 U1026 ( .A(n1308), .B(n1309), .ZN(n1117) );
XOR2_X1 U1027 ( .A(KEYINPUT59), .B(G107), .Z(n1309) );
XNOR2_X1 U1028 ( .A(G101), .B(G104), .ZN(n1308) );
NAND3_X1 U1029 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1082) );
NAND2_X1 U1030 ( .A1(KEYINPUT56), .A2(n1313), .ZN(n1312) );
INV_X1 U1031 ( .A(n1314), .ZN(n1313) );
OR3_X1 U1032 ( .A1(n1315), .A2(KEYINPUT56), .A3(G128), .ZN(n1311) );
NAND2_X1 U1033 ( .A1(G128), .A2(n1315), .ZN(n1310) );
NAND2_X1 U1034 ( .A1(KEYINPUT5), .A2(n1314), .ZN(n1315) );
XOR2_X1 U1035 ( .A(G146), .B(G143), .Z(n1314) );
XNOR2_X1 U1036 ( .A(n1089), .B(n1087), .ZN(n1161) );
XOR2_X1 U1037 ( .A(G134), .B(G137), .Z(n1087) );
NOR2_X1 U1038 ( .A1(n1225), .A2(n1224), .ZN(n1038) );
NAND2_X1 U1039 ( .A1(n1316), .A2(n1317), .ZN(n1224) );
NAND2_X1 U1040 ( .A1(KEYINPUT30), .A2(n1135), .ZN(n1317) );
XOR2_X1 U1041 ( .A(n1063), .B(n1318), .Z(n1316) );
NOR2_X1 U1042 ( .A1(KEYINPUT30), .A2(n1135), .ZN(n1318) );
INV_X1 U1043 ( .A(G475), .ZN(n1135) );
NAND2_X1 U1044 ( .A1(n1140), .A2(n1139), .ZN(n1063) );
XOR2_X1 U1045 ( .A(n1319), .B(n1320), .Z(n1140) );
XOR2_X1 U1046 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1047 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR2_X1 U1048 ( .A1(G146), .A2(KEYINPUT41), .ZN(n1324) );
NAND2_X1 U1049 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
NAND2_X1 U1050 ( .A1(G125), .A2(n1095), .ZN(n1326) );
XNOR2_X1 U1051 ( .A(KEYINPUT43), .B(n1092), .ZN(n1325) );
NAND2_X1 U1052 ( .A1(n1101), .A2(n1096), .ZN(n1092) );
INV_X1 U1053 ( .A(G125), .ZN(n1096) );
INV_X1 U1054 ( .A(n1095), .ZN(n1101) );
XOR2_X1 U1055 ( .A(G140), .B(KEYINPUT11), .Z(n1095) );
NAND2_X1 U1056 ( .A1(KEYINPUT55), .A2(n1089), .ZN(n1321) );
INV_X1 U1057 ( .A(G131), .ZN(n1089) );
XOR2_X1 U1058 ( .A(n1327), .B(n1328), .Z(n1319) );
XNOR2_X1 U1059 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U1060 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1061 ( .A(n1333), .B(KEYINPUT49), .Z(n1332) );
NAND3_X1 U1062 ( .A1(n1253), .A2(G143), .A3(G214), .ZN(n1333) );
NOR2_X1 U1063 ( .A1(n1334), .A2(G143), .ZN(n1331) );
AND2_X1 U1064 ( .A1(n1253), .A2(G214), .ZN(n1334) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1253) );
INV_X1 U1066 ( .A(G104), .ZN(n1329) );
XNOR2_X1 U1067 ( .A(G113), .B(G122), .ZN(n1327) );
NAND2_X1 U1068 ( .A1(n1335), .A2(n1336), .ZN(n1225) );
NAND2_X1 U1069 ( .A1(G478), .A2(n1065), .ZN(n1336) );
XNOR2_X1 U1070 ( .A(n1059), .B(KEYINPUT4), .ZN(n1335) );
NOR2_X1 U1071 ( .A1(n1065), .A2(G478), .ZN(n1059) );
NAND2_X1 U1072 ( .A1(n1130), .A2(n1139), .ZN(n1065) );
INV_X1 U1073 ( .A(G902), .ZN(n1139) );
XOR2_X1 U1074 ( .A(n1337), .B(n1338), .Z(n1130) );
NOR2_X1 U1075 ( .A1(KEYINPUT12), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1076 ( .A(n1340), .B(n1341), .Z(n1339) );
XOR2_X1 U1077 ( .A(G107), .B(n1342), .Z(n1341) );
XNOR2_X1 U1078 ( .A(n1343), .B(G116), .ZN(n1342) );
INV_X1 U1079 ( .A(G122), .ZN(n1343) );
XOR2_X1 U1080 ( .A(G128), .B(n1344), .Z(n1340) );
XOR2_X1 U1081 ( .A(G143), .B(G134), .Z(n1344) );
NAND2_X1 U1082 ( .A1(G217), .A2(n1272), .ZN(n1337) );
AND2_X1 U1083 ( .A1(G234), .A2(n1023), .ZN(n1272) );
INV_X1 U1084 ( .A(G953), .ZN(n1023) );
endmodule


