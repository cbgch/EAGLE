//Key = 1010100111100000001010100011101000011100101001100110100001101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323;

XNOR2_X1 U722 ( .A(G107), .B(n1000), .ZN(G9) );
NOR2_X1 U723 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR4_X1 U724 ( .A1(G953), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1002) );
NOR2_X1 U725 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U726 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR4_X1 U727 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1009) );
NOR3_X1 U728 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n1013) );
NOR2_X1 U729 ( .A1(n1017), .A2(n1018), .ZN(n1012) );
NOR2_X1 U730 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U731 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NAND2_X1 U732 ( .A1(n1023), .A2(n1024), .ZN(n1010) );
NOR3_X1 U733 ( .A1(n1020), .A2(n1025), .A3(n1014), .ZN(n1008) );
NOR2_X1 U734 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR3_X1 U735 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NOR3_X1 U736 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NOR2_X1 U737 ( .A1(n1034), .A2(n1024), .ZN(n1029) );
NOR2_X1 U738 ( .A1(n1035), .A2(n1011), .ZN(n1026) );
NOR3_X1 U739 ( .A1(n1003), .A2(G953), .A3(G952), .ZN(n1001) );
AND4_X1 U740 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1003) );
NOR3_X1 U741 ( .A1(n1040), .A2(n1031), .A3(n1041), .ZN(n1039) );
NOR2_X1 U742 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
INV_X1 U743 ( .A(n1024), .ZN(n1031) );
NAND3_X1 U744 ( .A1(n1044), .A2(n1045), .A3(n1022), .ZN(n1040) );
NOR3_X1 U745 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1038) );
NOR2_X1 U746 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
XOR2_X1 U747 ( .A(n1051), .B(n1052), .Z(n1036) );
XOR2_X1 U748 ( .A(KEYINPUT40), .B(n1053), .Z(n1052) );
NAND2_X1 U749 ( .A1(KEYINPUT46), .A2(n1054), .ZN(n1051) );
XOR2_X1 U750 ( .A(n1055), .B(n1056), .Z(G72) );
NOR2_X1 U751 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NOR2_X1 U752 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND2_X1 U753 ( .A1(n1061), .A2(n1062), .ZN(n1055) );
NAND2_X1 U754 ( .A1(n1063), .A2(n1058), .ZN(n1062) );
XOR2_X1 U755 ( .A(n1064), .B(n1065), .Z(n1063) );
NOR3_X1 U756 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
INV_X1 U757 ( .A(n1069), .ZN(n1067) );
XNOR2_X1 U758 ( .A(n1070), .B(KEYINPUT33), .ZN(n1064) );
NAND3_X1 U759 ( .A1(n1070), .A2(G900), .A3(G953), .ZN(n1061) );
NOR2_X1 U760 ( .A1(KEYINPUT12), .A2(n1071), .ZN(n1070) );
XOR2_X1 U761 ( .A(n1072), .B(n1073), .Z(n1071) );
XNOR2_X1 U762 ( .A(n1074), .B(n1075), .ZN(n1073) );
NOR2_X1 U763 ( .A1(KEYINPUT34), .A2(n1076), .ZN(n1075) );
XOR2_X1 U764 ( .A(G134), .B(n1077), .Z(n1076) );
XOR2_X1 U765 ( .A(n1078), .B(n1079), .Z(G69) );
NOR2_X1 U766 ( .A1(n1080), .A2(n1058), .ZN(n1079) );
AND2_X1 U767 ( .A1(G224), .A2(G898), .ZN(n1080) );
NAND2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1078) );
NAND2_X1 U769 ( .A1(n1083), .A2(n1058), .ZN(n1082) );
XNOR2_X1 U770 ( .A(n1084), .B(n1085), .ZN(n1083) );
NAND3_X1 U771 ( .A1(G898), .A2(n1084), .A3(G953), .ZN(n1081) );
XNOR2_X1 U772 ( .A(n1086), .B(n1087), .ZN(n1084) );
NOR2_X1 U773 ( .A1(n1088), .A2(n1089), .ZN(G66) );
XOR2_X1 U774 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U776 ( .A1(KEYINPUT30), .A2(n1094), .ZN(n1090) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1095), .ZN(G63) );
XNOR2_X1 U778 ( .A(n1096), .B(n1097), .ZN(n1095) );
XNOR2_X1 U779 ( .A(KEYINPUT22), .B(n1098), .ZN(n1097) );
NOR3_X1 U780 ( .A1(n1093), .A2(KEYINPUT31), .A3(n1099), .ZN(n1098) );
INV_X1 U781 ( .A(G478), .ZN(n1099) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1100), .ZN(G60) );
XOR2_X1 U783 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U784 ( .A1(n1050), .A2(n1093), .ZN(n1101) );
XOR2_X1 U785 ( .A(n1103), .B(n1104), .Z(G6) );
NOR2_X1 U786 ( .A1(n1088), .A2(n1105), .ZN(G57) );
XOR2_X1 U787 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U788 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U789 ( .A(n1110), .B(n1111), .Z(n1106) );
NOR2_X1 U790 ( .A1(n1054), .A2(n1093), .ZN(n1111) );
NOR2_X1 U791 ( .A1(n1088), .A2(n1112), .ZN(G54) );
NOR2_X1 U792 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U793 ( .A(n1115), .B(n1116), .Z(n1114) );
NOR2_X1 U794 ( .A1(n1043), .A2(n1093), .ZN(n1116) );
NOR2_X1 U795 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
INV_X1 U796 ( .A(KEYINPUT60), .ZN(n1118) );
XOR2_X1 U797 ( .A(n1119), .B(n1120), .Z(n1117) );
NOR2_X1 U798 ( .A1(KEYINPUT60), .A2(n1121), .ZN(n1113) );
XOR2_X1 U799 ( .A(n1119), .B(n1122), .Z(n1121) );
NAND2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1119) );
NAND2_X1 U801 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U802 ( .A(KEYINPUT8), .B(n1127), .Z(n1123) );
NOR2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(n1127) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1125) );
NOR2_X1 U805 ( .A1(n1088), .A2(n1130), .ZN(G51) );
XNOR2_X1 U806 ( .A(n1131), .B(n1132), .ZN(n1130) );
XOR2_X1 U807 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U808 ( .A1(n1093), .A2(n1135), .ZN(n1134) );
XOR2_X1 U809 ( .A(KEYINPUT20), .B(n1136), .Z(n1135) );
NAND2_X1 U810 ( .A1(G902), .A2(n1005), .ZN(n1093) );
NAND4_X1 U811 ( .A1(n1137), .A2(n1085), .A3(n1138), .A4(n1069), .ZN(n1005) );
NAND2_X1 U812 ( .A1(n1139), .A2(n1140), .ZN(n1069) );
XOR2_X1 U813 ( .A(n1141), .B(KEYINPUT41), .Z(n1139) );
INV_X1 U814 ( .A(n1066), .ZN(n1138) );
NAND3_X1 U815 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1066) );
AND2_X1 U816 ( .A1(n1145), .A2(n1146), .ZN(n1085) );
NOR4_X1 U817 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1146) );
NOR4_X1 U818 ( .A1(n1151), .A2(n1020), .A3(n1152), .A4(n1153), .ZN(n1150) );
XOR2_X1 U819 ( .A(KEYINPUT17), .B(n1154), .Z(n1153) );
AND4_X1 U820 ( .A1(n1000), .A2(n1155), .A3(n1156), .A4(n1104), .ZN(n1145) );
NAND4_X1 U821 ( .A1(n1015), .A2(n1157), .A3(n1034), .A4(n1158), .ZN(n1104) );
NAND4_X1 U822 ( .A1(n1157), .A2(n1016), .A3(n1034), .A4(n1158), .ZN(n1000) );
XOR2_X1 U823 ( .A(n1068), .B(KEYINPUT26), .Z(n1137) );
NAND3_X1 U824 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1068) );
NAND2_X1 U825 ( .A1(n1016), .A2(n1162), .ZN(n1161) );
NAND3_X1 U826 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
NAND3_X1 U827 ( .A1(n1166), .A2(n1152), .A3(n1167), .ZN(n1164) );
INV_X1 U828 ( .A(KEYINPUT0), .ZN(n1167) );
NAND2_X1 U829 ( .A1(KEYINPUT0), .A2(n1168), .ZN(n1163) );
NOR2_X1 U830 ( .A1(KEYINPUT1), .A2(n1169), .ZN(n1133) );
XOR2_X1 U831 ( .A(KEYINPUT47), .B(n1170), .Z(n1169) );
NOR2_X1 U832 ( .A1(n1058), .A2(G952), .ZN(n1088) );
XNOR2_X1 U833 ( .A(G146), .B(n1144), .ZN(G48) );
NAND2_X1 U834 ( .A1(n1171), .A2(n1015), .ZN(n1144) );
INV_X1 U835 ( .A(n1165), .ZN(n1171) );
XOR2_X1 U836 ( .A(G143), .B(n1172), .Z(G45) );
AND2_X1 U837 ( .A1(n1141), .A2(n1140), .ZN(n1172) );
NOR4_X1 U838 ( .A1(n1152), .A2(n1151), .A3(n1173), .A4(n1174), .ZN(n1140) );
XNOR2_X1 U839 ( .A(G140), .B(n1142), .ZN(G42) );
NAND3_X1 U840 ( .A1(n1032), .A2(n1015), .A3(n1166), .ZN(n1142) );
XOR2_X1 U841 ( .A(n1175), .B(n1143), .Z(G39) );
NAND4_X1 U842 ( .A1(n1166), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1143) );
XOR2_X1 U843 ( .A(n1179), .B(n1180), .Z(G36) );
NAND2_X1 U844 ( .A1(n1168), .A2(n1016), .ZN(n1180) );
XOR2_X1 U845 ( .A(n1181), .B(n1159), .Z(G33) );
NAND2_X1 U846 ( .A1(n1168), .A2(n1015), .ZN(n1159) );
AND2_X1 U847 ( .A1(n1166), .A2(n1033), .ZN(n1168) );
AND3_X1 U848 ( .A1(n1023), .A2(n1141), .A3(n1182), .ZN(n1166) );
AND3_X1 U849 ( .A1(n1024), .A2(n1022), .A3(n1183), .ZN(n1182) );
INV_X1 U850 ( .A(n1028), .ZN(n1023) );
XOR2_X1 U851 ( .A(n1037), .B(KEYINPUT35), .Z(n1028) );
XOR2_X1 U852 ( .A(G128), .B(n1184), .Z(G30) );
NOR3_X1 U853 ( .A1(n1165), .A2(KEYINPUT16), .A3(n1185), .ZN(n1184) );
NAND4_X1 U854 ( .A1(n1178), .A2(n1157), .A3(n1177), .A4(n1141), .ZN(n1165) );
INV_X1 U855 ( .A(n1151), .ZN(n1157) );
XOR2_X1 U856 ( .A(G101), .B(n1186), .Z(G3) );
AND2_X1 U857 ( .A1(n1033), .A2(n1187), .ZN(n1186) );
INV_X1 U858 ( .A(n1152), .ZN(n1033) );
XNOR2_X1 U859 ( .A(G125), .B(n1160), .ZN(G27) );
NAND3_X1 U860 ( .A1(n1032), .A2(n1015), .A3(n1188), .ZN(n1160) );
AND3_X1 U861 ( .A1(n1017), .A2(n1141), .A3(n1189), .ZN(n1188) );
NAND2_X1 U862 ( .A1(n1007), .A2(n1190), .ZN(n1141) );
NAND4_X1 U863 ( .A1(G953), .A2(G902), .A3(n1191), .A4(n1060), .ZN(n1190) );
INV_X1 U864 ( .A(G900), .ZN(n1060) );
NAND2_X1 U865 ( .A1(n1192), .A2(n1193), .ZN(G24) );
NAND2_X1 U866 ( .A1(G122), .A2(n1156), .ZN(n1193) );
XOR2_X1 U867 ( .A(n1194), .B(KEYINPUT54), .Z(n1192) );
OR2_X1 U868 ( .A1(n1156), .A2(G122), .ZN(n1194) );
NAND4_X1 U869 ( .A1(n1048), .A2(n1034), .A3(n1017), .A4(n1195), .ZN(n1156) );
NOR3_X1 U870 ( .A1(n1035), .A2(n1154), .A3(n1174), .ZN(n1195) );
INV_X1 U871 ( .A(n1011), .ZN(n1034) );
NAND2_X1 U872 ( .A1(n1196), .A2(n1197), .ZN(n1011) );
XOR2_X1 U873 ( .A(n1198), .B(G119), .Z(G21) );
NAND2_X1 U874 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NAND2_X1 U875 ( .A1(n1149), .A2(n1201), .ZN(n1200) );
INV_X1 U876 ( .A(KEYINPUT29), .ZN(n1201) );
NOR2_X1 U877 ( .A1(n1202), .A2(n1035), .ZN(n1149) );
NAND3_X1 U878 ( .A1(n1189), .A2(n1202), .A3(KEYINPUT29), .ZN(n1199) );
NAND4_X1 U879 ( .A1(n1176), .A2(n1017), .A3(n1203), .A4(n1178), .ZN(n1202) );
NOR2_X1 U880 ( .A1(n1154), .A2(n1204), .ZN(n1203) );
INV_X1 U881 ( .A(n1014), .ZN(n1017) );
INV_X1 U882 ( .A(n1020), .ZN(n1176) );
XOR2_X1 U883 ( .A(n1148), .B(n1205), .Z(G18) );
NOR2_X1 U884 ( .A1(KEYINPUT19), .A2(n1206), .ZN(n1205) );
AND2_X1 U885 ( .A1(n1207), .A2(n1016), .ZN(n1148) );
INV_X1 U886 ( .A(n1185), .ZN(n1016) );
NAND2_X1 U887 ( .A1(n1174), .A2(n1048), .ZN(n1185) );
XOR2_X1 U888 ( .A(G113), .B(n1147), .Z(G15) );
AND2_X1 U889 ( .A1(n1015), .A2(n1207), .ZN(n1147) );
NOR4_X1 U890 ( .A1(n1152), .A2(n1014), .A3(n1035), .A4(n1154), .ZN(n1207) );
NAND2_X1 U891 ( .A1(n1021), .A2(n1022), .ZN(n1014) );
INV_X1 U892 ( .A(n1183), .ZN(n1021) );
NAND2_X1 U893 ( .A1(n1208), .A2(n1197), .ZN(n1152) );
INV_X1 U894 ( .A(n1178), .ZN(n1197) );
XOR2_X1 U895 ( .A(KEYINPUT18), .B(n1204), .Z(n1208) );
INV_X1 U896 ( .A(n1177), .ZN(n1204) );
NOR2_X1 U897 ( .A1(n1048), .A2(n1174), .ZN(n1015) );
NAND2_X1 U898 ( .A1(n1209), .A2(n1210), .ZN(G12) );
OR2_X1 U899 ( .A1(n1155), .A2(G110), .ZN(n1210) );
XOR2_X1 U900 ( .A(n1211), .B(KEYINPUT38), .Z(n1209) );
NAND2_X1 U901 ( .A1(G110), .A2(n1155), .ZN(n1211) );
NAND2_X1 U902 ( .A1(n1032), .A2(n1187), .ZN(n1155) );
NOR3_X1 U903 ( .A1(n1151), .A2(n1154), .A3(n1020), .ZN(n1187) );
NAND2_X1 U904 ( .A1(n1174), .A2(n1173), .ZN(n1020) );
INV_X1 U905 ( .A(n1048), .ZN(n1173) );
XOR2_X1 U906 ( .A(n1212), .B(n1213), .Z(n1048) );
XOR2_X1 U907 ( .A(KEYINPUT52), .B(G478), .Z(n1213) );
NAND2_X1 U908 ( .A1(n1096), .A2(n1214), .ZN(n1212) );
XNOR2_X1 U909 ( .A(n1215), .B(n1216), .ZN(n1096) );
XOR2_X1 U910 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U911 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U912 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
INV_X1 U913 ( .A(G217), .ZN(n1222) );
NAND2_X1 U914 ( .A1(n1223), .A2(n1224), .ZN(n1219) );
NAND2_X1 U915 ( .A1(G107), .A2(n1225), .ZN(n1224) );
XOR2_X1 U916 ( .A(n1226), .B(KEYINPUT3), .Z(n1223) );
OR2_X1 U917 ( .A1(n1225), .A2(G107), .ZN(n1226) );
XOR2_X1 U918 ( .A(n1206), .B(n1227), .Z(n1225) );
XOR2_X1 U919 ( .A(n1228), .B(n1229), .Z(n1215) );
XOR2_X1 U920 ( .A(KEYINPUT48), .B(G134), .Z(n1229) );
NAND2_X1 U921 ( .A1(KEYINPUT58), .A2(n1230), .ZN(n1228) );
AND3_X1 U922 ( .A1(n1231), .A2(n1232), .A3(n1045), .ZN(n1174) );
NAND2_X1 U923 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
NAND2_X1 U924 ( .A1(n1050), .A2(n1233), .ZN(n1232) );
OR3_X1 U925 ( .A1(n1050), .A2(n1049), .A3(n1233), .ZN(n1231) );
INV_X1 U926 ( .A(KEYINPUT62), .ZN(n1233) );
NOR2_X1 U927 ( .A1(n1102), .A2(n1234), .ZN(n1049) );
XNOR2_X1 U928 ( .A(n1235), .B(n1236), .ZN(n1102) );
XOR2_X1 U929 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U930 ( .A(n1239), .B(n1240), .ZN(n1238) );
NOR4_X1 U931 ( .A1(KEYINPUT59), .A2(G953), .A3(G237), .A4(n1241), .ZN(n1240) );
XNOR2_X1 U932 ( .A(G214), .B(KEYINPUT44), .ZN(n1241) );
NAND2_X1 U933 ( .A1(KEYINPUT27), .A2(n1181), .ZN(n1239) );
XOR2_X1 U934 ( .A(KEYINPUT13), .B(n1242), .Z(n1237) );
NOR2_X1 U935 ( .A1(KEYINPUT14), .A2(n1243), .ZN(n1242) );
XOR2_X1 U936 ( .A(G104), .B(n1244), .Z(n1243) );
XOR2_X1 U937 ( .A(G122), .B(G113), .Z(n1244) );
XOR2_X1 U938 ( .A(n1245), .B(n1246), .Z(n1235) );
XOR2_X1 U939 ( .A(n1247), .B(n1248), .Z(n1245) );
INV_X1 U940 ( .A(n1249), .ZN(n1248) );
NAND2_X1 U941 ( .A1(KEYINPUT45), .A2(n1074), .ZN(n1247) );
INV_X1 U942 ( .A(G475), .ZN(n1050) );
INV_X1 U943 ( .A(n1158), .ZN(n1154) );
NAND2_X1 U944 ( .A1(n1250), .A2(n1007), .ZN(n1158) );
NAND3_X1 U945 ( .A1(n1191), .A2(n1058), .A3(n1251), .ZN(n1007) );
XNOR2_X1 U946 ( .A(G952), .B(KEYINPUT2), .ZN(n1251) );
NAND4_X1 U947 ( .A1(G953), .A2(G902), .A3(n1191), .A4(n1252), .ZN(n1250) );
INV_X1 U948 ( .A(G898), .ZN(n1252) );
NAND2_X1 U949 ( .A1(G237), .A2(G234), .ZN(n1191) );
NAND3_X1 U950 ( .A1(n1183), .A2(n1022), .A3(n1189), .ZN(n1151) );
INV_X1 U951 ( .A(n1035), .ZN(n1189) );
NAND2_X1 U952 ( .A1(n1253), .A2(n1024), .ZN(n1035) );
NAND2_X1 U953 ( .A1(G214), .A2(n1254), .ZN(n1024) );
INV_X1 U954 ( .A(n1037), .ZN(n1253) );
XOR2_X1 U955 ( .A(n1255), .B(n1136), .Z(n1037) );
AND2_X1 U956 ( .A1(G210), .A2(n1254), .ZN(n1136) );
NAND2_X1 U957 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
NAND2_X1 U958 ( .A1(n1258), .A2(n1259), .ZN(n1255) );
XNOR2_X1 U959 ( .A(n1131), .B(n1170), .ZN(n1259) );
XNOR2_X1 U960 ( .A(n1260), .B(n1261), .ZN(n1170) );
INV_X1 U961 ( .A(n1072), .ZN(n1261) );
XNOR2_X1 U962 ( .A(G125), .B(n1129), .ZN(n1072) );
NAND2_X1 U963 ( .A1(G224), .A2(n1058), .ZN(n1260) );
NAND2_X1 U964 ( .A1(n1262), .A2(n1263), .ZN(n1131) );
NAND2_X1 U965 ( .A1(n1264), .A2(n1087), .ZN(n1263) );
XOR2_X1 U966 ( .A(n1265), .B(KEYINPUT6), .Z(n1262) );
OR2_X1 U967 ( .A1(n1087), .A2(n1264), .ZN(n1265) );
XOR2_X1 U968 ( .A(n1086), .B(KEYINPUT10), .Z(n1264) );
XOR2_X1 U969 ( .A(n1227), .B(n1266), .Z(n1086) );
NOR2_X1 U970 ( .A1(G110), .A2(KEYINPUT51), .ZN(n1266) );
INV_X1 U971 ( .A(G122), .ZN(n1227) );
XNOR2_X1 U972 ( .A(n1267), .B(n1268), .ZN(n1087) );
XNOR2_X1 U973 ( .A(n1269), .B(n1270), .ZN(n1268) );
NOR2_X1 U974 ( .A1(G104), .A2(KEYINPUT25), .ZN(n1270) );
NAND2_X1 U975 ( .A1(KEYINPUT50), .A2(n1271), .ZN(n1269) );
XNOR2_X1 U976 ( .A(n1272), .B(n1273), .ZN(n1267) );
XNOR2_X1 U977 ( .A(KEYINPUT11), .B(n1234), .ZN(n1258) );
INV_X1 U978 ( .A(n1214), .ZN(n1234) );
NAND2_X1 U979 ( .A1(G221), .A2(n1274), .ZN(n1022) );
NAND3_X1 U980 ( .A1(n1275), .A2(n1276), .A3(n1044), .ZN(n1183) );
NAND2_X1 U981 ( .A1(n1042), .A2(n1043), .ZN(n1044) );
NAND2_X1 U982 ( .A1(KEYINPUT24), .A2(n1043), .ZN(n1276) );
OR3_X1 U983 ( .A1(n1042), .A2(KEYINPUT24), .A3(n1043), .ZN(n1275) );
INV_X1 U984 ( .A(G469), .ZN(n1043) );
AND2_X1 U985 ( .A1(n1277), .A2(n1214), .ZN(n1042) );
XOR2_X1 U986 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U987 ( .A(n1129), .B(n1120), .Z(n1279) );
INV_X1 U988 ( .A(n1122), .ZN(n1120) );
XNOR2_X1 U989 ( .A(n1074), .B(n1280), .ZN(n1122) );
XOR2_X1 U990 ( .A(G110), .B(n1281), .Z(n1280) );
NOR2_X1 U991 ( .A1(G953), .A2(n1059), .ZN(n1281) );
INV_X1 U992 ( .A(G227), .ZN(n1059) );
XNOR2_X1 U993 ( .A(n1282), .B(n1283), .ZN(n1278) );
NAND2_X1 U994 ( .A1(KEYINPUT7), .A2(n1128), .ZN(n1283) );
XOR2_X1 U995 ( .A(n1103), .B(n1272), .Z(n1128) );
XOR2_X1 U996 ( .A(G107), .B(n1109), .Z(n1272) );
INV_X1 U997 ( .A(G104), .ZN(n1103) );
NAND2_X1 U998 ( .A1(KEYINPUT42), .A2(n1284), .ZN(n1282) );
AND2_X1 U999 ( .A1(n1178), .A2(n1196), .ZN(n1032) );
XOR2_X1 U1000 ( .A(n1177), .B(KEYINPUT49), .Z(n1196) );
XOR2_X1 U1001 ( .A(n1054), .B(n1285), .Z(n1177) );
NOR2_X1 U1002 ( .A1(n1053), .A2(KEYINPUT32), .ZN(n1285) );
AND2_X1 U1003 ( .A1(n1286), .A2(n1214), .ZN(n1053) );
XOR2_X1 U1004 ( .A(n1108), .B(n1287), .Z(n1286) );
NOR3_X1 U1005 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1287) );
NOR2_X1 U1006 ( .A1(n1291), .A2(n1109), .ZN(n1290) );
INV_X1 U1007 ( .A(n1292), .ZN(n1109) );
NOR2_X1 U1008 ( .A1(KEYINPUT15), .A2(n1293), .ZN(n1291) );
XOR2_X1 U1009 ( .A(n1110), .B(KEYINPUT56), .Z(n1293) );
NOR3_X1 U1010 ( .A1(n1292), .A2(KEYINPUT15), .A3(n1110), .ZN(n1289) );
XNOR2_X1 U1011 ( .A(G101), .B(KEYINPUT43), .ZN(n1292) );
AND2_X1 U1012 ( .A1(n1110), .A2(KEYINPUT15), .ZN(n1288) );
NAND3_X1 U1013 ( .A1(n1256), .A2(n1058), .A3(G210), .ZN(n1110) );
INV_X1 U1014 ( .A(G237), .ZN(n1256) );
XOR2_X1 U1015 ( .A(n1294), .B(n1126), .Z(n1108) );
INV_X1 U1016 ( .A(n1284), .ZN(n1126) );
XNOR2_X1 U1017 ( .A(n1077), .B(n1295), .ZN(n1284) );
NOR2_X1 U1018 ( .A1(KEYINPUT39), .A2(n1296), .ZN(n1295) );
XOR2_X1 U1019 ( .A(n1179), .B(KEYINPUT63), .Z(n1296) );
INV_X1 U1020 ( .A(G134), .ZN(n1179) );
XOR2_X1 U1021 ( .A(n1181), .B(n1175), .Z(n1077) );
INV_X1 U1022 ( .A(G137), .ZN(n1175) );
INV_X1 U1023 ( .A(G131), .ZN(n1181) );
XOR2_X1 U1024 ( .A(n1297), .B(n1129), .Z(n1294) );
XNOR2_X1 U1025 ( .A(n1298), .B(n1246), .ZN(n1129) );
INV_X1 U1026 ( .A(n1217), .ZN(n1246) );
XNOR2_X1 U1027 ( .A(G143), .B(KEYINPUT28), .ZN(n1217) );
XOR2_X1 U1028 ( .A(G146), .B(n1230), .Z(n1298) );
NAND3_X1 U1029 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1297) );
OR2_X1 U1030 ( .A1(n1273), .A2(KEYINPUT36), .ZN(n1301) );
NAND3_X1 U1031 ( .A1(KEYINPUT36), .A2(n1273), .A3(G113), .ZN(n1300) );
NAND2_X1 U1032 ( .A1(n1302), .A2(n1271), .ZN(n1299) );
INV_X1 U1033 ( .A(G113), .ZN(n1271) );
NAND2_X1 U1034 ( .A1(n1303), .A2(KEYINPUT36), .ZN(n1302) );
XNOR2_X1 U1035 ( .A(n1273), .B(KEYINPUT4), .ZN(n1303) );
XOR2_X1 U1036 ( .A(n1206), .B(n1304), .Z(n1273) );
INV_X1 U1037 ( .A(G116), .ZN(n1206) );
INV_X1 U1038 ( .A(G472), .ZN(n1054) );
XNOR2_X1 U1039 ( .A(n1046), .B(KEYINPUT37), .ZN(n1178) );
XOR2_X1 U1040 ( .A(n1305), .B(n1092), .Z(n1046) );
NAND2_X1 U1041 ( .A1(G217), .A2(n1274), .ZN(n1092) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1257), .ZN(n1274) );
INV_X1 U1043 ( .A(G902), .ZN(n1257) );
NAND2_X1 U1044 ( .A1(n1094), .A2(n1214), .ZN(n1305) );
XOR2_X1 U1045 ( .A(G902), .B(KEYINPUT9), .Z(n1214) );
XNOR2_X1 U1046 ( .A(n1306), .B(n1307), .ZN(n1094) );
XOR2_X1 U1047 ( .A(n1249), .B(n1308), .Z(n1307) );
XNOR2_X1 U1048 ( .A(n1309), .B(n1310), .ZN(n1308) );
NOR2_X1 U1049 ( .A1(KEYINPUT61), .A2(n1074), .ZN(n1310) );
XOR2_X1 U1050 ( .A(G140), .B(KEYINPUT53), .Z(n1074) );
NOR3_X1 U1051 ( .A1(n1221), .A2(KEYINPUT5), .A3(n1311), .ZN(n1309) );
INV_X1 U1052 ( .A(G221), .ZN(n1311) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1058), .ZN(n1221) );
INV_X1 U1054 ( .A(G953), .ZN(n1058) );
XNOR2_X1 U1055 ( .A(G125), .B(G146), .ZN(n1249) );
XOR2_X1 U1056 ( .A(n1312), .B(n1313), .Z(n1306) );
XOR2_X1 U1057 ( .A(KEYINPUT57), .B(G137), .Z(n1313) );
XOR2_X1 U1058 ( .A(n1314), .B(G110), .Z(n1312) );
NAND4_X1 U1059 ( .A1(n1315), .A2(n1316), .A3(n1317), .A4(n1318), .ZN(n1314) );
NAND3_X1 U1060 ( .A1(n1319), .A2(n1230), .A3(n1320), .ZN(n1318) );
INV_X1 U1061 ( .A(KEYINPUT23), .ZN(n1320) );
INV_X1 U1062 ( .A(G128), .ZN(n1230) );
OR2_X1 U1063 ( .A1(n1304), .A2(KEYINPUT21), .ZN(n1319) );
NAND3_X1 U1064 ( .A1(G128), .A2(n1321), .A3(KEYINPUT23), .ZN(n1317) );
NAND2_X1 U1065 ( .A1(KEYINPUT21), .A2(G119), .ZN(n1321) );
NAND2_X1 U1066 ( .A1(KEYINPUT55), .A2(n1304), .ZN(n1316) );
INV_X1 U1067 ( .A(G119), .ZN(n1304) );
NAND3_X1 U1068 ( .A1(n1322), .A2(n1323), .A3(G119), .ZN(n1315) );
INV_X1 U1069 ( .A(KEYINPUT55), .ZN(n1323) );
XOR2_X1 U1070 ( .A(KEYINPUT21), .B(G128), .Z(n1322) );
endmodule


