//Key = 1010100111010110011101000111110001000110111001010101101001011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328;

XNOR2_X1 U711 ( .A(G107), .B(n997), .ZN(G9) );
NAND3_X1 U712 ( .A1(n998), .A2(n999), .A3(KEYINPUT49), .ZN(n997) );
NOR2_X1 U713 ( .A1(n1000), .A2(n1001), .ZN(G75) );
NOR4_X1 U714 ( .A1(n1002), .A2(n1003), .A3(G953), .A4(n1004), .ZN(n1001) );
NOR3_X1 U715 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1003) );
INV_X1 U716 ( .A(n1008), .ZN(n1007) );
NAND3_X1 U717 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1002) );
NAND3_X1 U718 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
NAND2_X1 U719 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NAND3_X1 U720 ( .A1(n1008), .A2(n1017), .A3(n1018), .ZN(n1016) );
NAND2_X1 U721 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NAND2_X1 U722 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U723 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U724 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
INV_X1 U725 ( .A(n1027), .ZN(n1023) );
NAND2_X1 U726 ( .A1(n1028), .A2(n1029), .ZN(n1019) );
NAND2_X1 U727 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U728 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U729 ( .A1(n1034), .A2(n1035), .ZN(n1015) );
OR2_X1 U730 ( .A1(n1036), .A2(n998), .ZN(n1035) );
INV_X1 U731 ( .A(n1005), .ZN(n1034) );
NAND3_X1 U732 ( .A1(n1028), .A2(n1021), .A3(n1018), .ZN(n1005) );
INV_X1 U733 ( .A(n1037), .ZN(n1018) );
NOR3_X1 U734 ( .A1(n1004), .A2(G953), .A3(G952), .ZN(n1000) );
AND4_X1 U735 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1004) );
NOR4_X1 U736 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
XNOR2_X1 U737 ( .A(G472), .B(n1046), .ZN(n1045) );
XOR2_X1 U738 ( .A(n1047), .B(KEYINPUT45), .Z(n1044) );
XOR2_X1 U739 ( .A(KEYINPUT41), .B(n1048), .Z(n1043) );
NOR2_X1 U740 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
INV_X1 U741 ( .A(n1051), .ZN(n1050) );
NOR2_X1 U742 ( .A1(n1052), .A2(n1053), .ZN(n1049) );
NAND2_X1 U743 ( .A1(n1054), .A2(n1055), .ZN(n1042) );
XOR2_X1 U744 ( .A(n1056), .B(KEYINPUT44), .Z(n1055) );
XOR2_X1 U745 ( .A(n1057), .B(KEYINPUT31), .Z(n1054) );
NOR3_X1 U746 ( .A1(n1058), .A2(n1032), .A3(n1025), .ZN(n1040) );
XOR2_X1 U747 ( .A(n1059), .B(n1060), .Z(n1038) );
NOR2_X1 U748 ( .A1(KEYINPUT35), .A2(n1061), .ZN(n1059) );
XOR2_X1 U749 ( .A(n1062), .B(KEYINPUT26), .Z(n1061) );
XOR2_X1 U750 ( .A(n1063), .B(n1064), .Z(G72) );
NAND2_X1 U751 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND3_X1 U752 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
INV_X1 U753 ( .A(n1070), .ZN(n1069) );
XOR2_X1 U754 ( .A(KEYINPUT19), .B(n1071), .Z(n1067) );
NAND2_X1 U755 ( .A1(n1071), .A2(n1070), .ZN(n1065) );
XNOR2_X1 U756 ( .A(n1072), .B(n1073), .ZN(n1070) );
XNOR2_X1 U757 ( .A(n1074), .B(G125), .ZN(n1073) );
XNOR2_X1 U758 ( .A(n1075), .B(n1076), .ZN(n1072) );
NOR2_X1 U759 ( .A1(G953), .A2(n1011), .ZN(n1071) );
NAND2_X1 U760 ( .A1(n1077), .A2(n1068), .ZN(n1063) );
INV_X1 U761 ( .A(n1078), .ZN(n1068) );
OR2_X1 U762 ( .A1(n1079), .A2(G227), .ZN(n1077) );
NAND2_X1 U763 ( .A1(n1080), .A2(n1081), .ZN(G69) );
NAND2_X1 U764 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U765 ( .A1(G953), .A2(n1084), .ZN(n1083) );
NAND2_X1 U766 ( .A1(G898), .A2(G224), .ZN(n1084) );
NAND2_X1 U767 ( .A1(n1085), .A2(n1086), .ZN(n1080) );
NAND2_X1 U768 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U769 ( .A1(G953), .A2(n1089), .ZN(n1088) );
INV_X1 U770 ( .A(n1082), .ZN(n1085) );
XNOR2_X1 U771 ( .A(n1090), .B(n1091), .ZN(n1082) );
NOR2_X1 U772 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U773 ( .A(KEYINPUT55), .B(n1079), .ZN(n1093) );
NOR2_X1 U774 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
XOR2_X1 U775 ( .A(n1096), .B(KEYINPUT62), .Z(n1094) );
NAND2_X1 U776 ( .A1(n1097), .A2(n1087), .ZN(n1090) );
INV_X1 U777 ( .A(n1098), .ZN(n1087) );
XNOR2_X1 U778 ( .A(n1099), .B(n1100), .ZN(n1097) );
NOR2_X1 U779 ( .A1(n1101), .A2(n1102), .ZN(G66) );
XOR2_X1 U780 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND2_X1 U781 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NOR2_X1 U782 ( .A1(n1101), .A2(n1107), .ZN(G63) );
XOR2_X1 U783 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U784 ( .A1(n1105), .A2(G478), .ZN(n1108) );
NOR2_X1 U785 ( .A1(n1101), .A2(n1110), .ZN(G60) );
XOR2_X1 U786 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U787 ( .A(n1113), .B(KEYINPUT17), .Z(n1112) );
NAND2_X1 U788 ( .A1(n1105), .A2(G475), .ZN(n1113) );
XNOR2_X1 U789 ( .A(G104), .B(n1114), .ZN(G6) );
NOR2_X1 U790 ( .A1(n1101), .A2(n1115), .ZN(G57) );
XOR2_X1 U791 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U792 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U793 ( .A1(KEYINPUT57), .A2(G101), .ZN(n1118) );
XOR2_X1 U794 ( .A(n1120), .B(n1121), .Z(n1116) );
XNOR2_X1 U795 ( .A(n1122), .B(n1123), .ZN(n1121) );
NOR2_X1 U796 ( .A1(KEYINPUT39), .A2(n1124), .ZN(n1122) );
NOR3_X1 U797 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
NOR2_X1 U798 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U799 ( .A1(KEYINPUT24), .A2(n1130), .ZN(n1128) );
XNOR2_X1 U800 ( .A(KEYINPUT16), .B(n1131), .ZN(n1130) );
NOR3_X1 U801 ( .A1(n1132), .A2(KEYINPUT24), .A3(n1133), .ZN(n1126) );
AND2_X1 U802 ( .A1(n1133), .A2(KEYINPUT24), .ZN(n1125) );
NAND2_X1 U803 ( .A1(n1105), .A2(G472), .ZN(n1120) );
NOR2_X1 U804 ( .A1(n1101), .A2(n1134), .ZN(G54) );
XOR2_X1 U805 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U806 ( .A(n1137), .B(n1138), .ZN(n1136) );
XNOR2_X1 U807 ( .A(n1133), .B(n1139), .ZN(n1135) );
XOR2_X1 U808 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U809 ( .A1(KEYINPUT29), .A2(n1142), .ZN(n1141) );
NAND2_X1 U810 ( .A1(n1105), .A2(G469), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1101), .A2(n1143), .ZN(G51) );
XOR2_X1 U812 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U813 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U814 ( .A1(n1105), .A2(G210), .ZN(n1146) );
AND2_X1 U815 ( .A1(G902), .A2(n1148), .ZN(n1105) );
NAND2_X1 U816 ( .A1(n1149), .A2(n1011), .ZN(n1148) );
AND4_X1 U817 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1011) );
AND4_X1 U818 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
NAND2_X1 U819 ( .A1(n1158), .A2(n1159), .ZN(n1152) );
NAND2_X1 U820 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U821 ( .A1(n1028), .A2(n1162), .ZN(n1161) );
XOR2_X1 U822 ( .A(n1163), .B(KEYINPUT34), .Z(n1160) );
NAND2_X1 U823 ( .A1(n1164), .A2(n1021), .ZN(n1150) );
XOR2_X1 U824 ( .A(n1165), .B(KEYINPUT14), .Z(n1164) );
XNOR2_X1 U825 ( .A(n1009), .B(KEYINPUT42), .ZN(n1149) );
NOR2_X1 U826 ( .A1(n1096), .A2(n1095), .ZN(n1009) );
NAND3_X1 U827 ( .A1(n1166), .A2(n1114), .A3(n1167), .ZN(n1095) );
OR2_X1 U828 ( .A1(n1168), .A2(n1006), .ZN(n1167) );
NOR2_X1 U829 ( .A1(n1169), .A2(n1170), .ZN(n1006) );
NAND2_X1 U830 ( .A1(n1036), .A2(n999), .ZN(n1114) );
NAND2_X1 U831 ( .A1(n998), .A2(n999), .ZN(n1166) );
AND3_X1 U832 ( .A1(n1158), .A2(n1027), .A3(n1171), .ZN(n999) );
AND3_X1 U833 ( .A1(n1014), .A2(n1172), .A3(n1012), .ZN(n1171) );
NAND4_X1 U834 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1096) );
XNOR2_X1 U835 ( .A(KEYINPUT8), .B(n1177), .ZN(n1144) );
NOR2_X1 U836 ( .A1(n1079), .A2(G952), .ZN(n1101) );
XOR2_X1 U837 ( .A(n1151), .B(n1178), .Z(G48) );
XOR2_X1 U838 ( .A(KEYINPUT52), .B(G146), .Z(n1178) );
NAND3_X1 U839 ( .A1(n1179), .A2(n1158), .A3(n1036), .ZN(n1151) );
XOR2_X1 U840 ( .A(G143), .B(n1180), .Z(G45) );
NOR2_X1 U841 ( .A1(n1030), .A2(n1163), .ZN(n1180) );
NAND2_X1 U842 ( .A1(n1181), .A2(n1182), .ZN(n1163) );
NAND2_X1 U843 ( .A1(n1183), .A2(n1184), .ZN(G42) );
NAND2_X1 U844 ( .A1(n1185), .A2(n1074), .ZN(n1184) );
XOR2_X1 U845 ( .A(KEYINPUT51), .B(n1186), .Z(n1183) );
NOR2_X1 U846 ( .A1(n1185), .A2(n1074), .ZN(n1186) );
INV_X1 U847 ( .A(n1157), .ZN(n1185) );
NAND3_X1 U848 ( .A1(n1021), .A2(n1027), .A3(n1162), .ZN(n1157) );
XOR2_X1 U849 ( .A(n1156), .B(n1187), .Z(G39) );
NAND2_X1 U850 ( .A1(KEYINPUT4), .A2(G137), .ZN(n1187) );
NAND3_X1 U851 ( .A1(n1021), .A2(n1179), .A3(n1008), .ZN(n1156) );
XNOR2_X1 U852 ( .A(G134), .B(n1155), .ZN(G36) );
NAND3_X1 U853 ( .A1(n1182), .A2(n998), .A3(n1021), .ZN(n1155) );
INV_X1 U854 ( .A(n1188), .ZN(n1021) );
XNOR2_X1 U855 ( .A(n1189), .B(n1190), .ZN(G33) );
NOR2_X1 U856 ( .A1(n1188), .A2(n1165), .ZN(n1190) );
NAND2_X1 U857 ( .A1(n1036), .A2(n1182), .ZN(n1165) );
AND3_X1 U858 ( .A1(n1027), .A2(n1191), .A3(n1169), .ZN(n1182) );
NAND2_X1 U859 ( .A1(n1033), .A2(n1192), .ZN(n1188) );
XNOR2_X1 U860 ( .A(G128), .B(n1154), .ZN(G30) );
NAND3_X1 U861 ( .A1(n998), .A2(n1158), .A3(n1179), .ZN(n1154) );
AND4_X1 U862 ( .A1(n1193), .A2(n1194), .A3(n1027), .A4(n1191), .ZN(n1179) );
XOR2_X1 U863 ( .A(G101), .B(n1195), .Z(G3) );
NOR2_X1 U864 ( .A1(n1196), .A2(n1168), .ZN(n1195) );
INV_X1 U865 ( .A(n1169), .ZN(n1196) );
NAND3_X1 U866 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(G27) );
NAND2_X1 U867 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
INV_X1 U868 ( .A(KEYINPUT7), .ZN(n1201) );
NAND2_X1 U869 ( .A1(G125), .A2(n1202), .ZN(n1200) );
NAND3_X1 U870 ( .A1(KEYINPUT7), .A2(n1203), .A3(G125), .ZN(n1198) );
NAND2_X1 U871 ( .A1(KEYINPUT59), .A2(n1204), .ZN(n1203) );
NAND3_X1 U872 ( .A1(KEYINPUT59), .A2(n1204), .A3(n1177), .ZN(n1197) );
INV_X1 U873 ( .A(n1202), .ZN(n1204) );
NAND3_X1 U874 ( .A1(n1162), .A2(n1205), .A3(n1028), .ZN(n1202) );
XNOR2_X1 U875 ( .A(KEYINPUT15), .B(n1030), .ZN(n1205) );
INV_X1 U876 ( .A(n1158), .ZN(n1030) );
AND3_X1 U877 ( .A1(n1170), .A2(n1191), .A3(n1036), .ZN(n1162) );
NAND2_X1 U878 ( .A1(n1037), .A2(n1206), .ZN(n1191) );
NAND3_X1 U879 ( .A1(G902), .A2(n1207), .A3(n1078), .ZN(n1206) );
NOR2_X1 U880 ( .A1(G900), .A2(n1079), .ZN(n1078) );
XNOR2_X1 U881 ( .A(G122), .B(n1174), .ZN(G24) );
NAND4_X1 U882 ( .A1(n1208), .A2(n1181), .A3(n1014), .A4(n1012), .ZN(n1174) );
AND2_X1 U883 ( .A1(n1209), .A2(n1210), .ZN(n1181) );
XNOR2_X1 U884 ( .A(n1211), .B(KEYINPUT63), .ZN(n1209) );
XNOR2_X1 U885 ( .A(G119), .B(n1212), .ZN(G21) );
NAND2_X1 U886 ( .A1(KEYINPUT11), .A2(n1213), .ZN(n1212) );
INV_X1 U887 ( .A(n1173), .ZN(n1213) );
NAND4_X1 U888 ( .A1(n1208), .A2(n1008), .A3(n1193), .A4(n1194), .ZN(n1173) );
XNOR2_X1 U889 ( .A(G116), .B(n1175), .ZN(G18) );
NAND3_X1 U890 ( .A1(n1169), .A2(n998), .A3(n1208), .ZN(n1175) );
NOR2_X1 U891 ( .A1(n1210), .A2(n1211), .ZN(n998) );
NAND2_X1 U892 ( .A1(n1214), .A2(n1215), .ZN(G15) );
NAND2_X1 U893 ( .A1(n1216), .A2(n1176), .ZN(n1215) );
XOR2_X1 U894 ( .A(KEYINPUT46), .B(G113), .Z(n1216) );
XOR2_X1 U895 ( .A(n1217), .B(KEYINPUT56), .Z(n1214) );
NAND2_X1 U896 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U897 ( .A(n1176), .ZN(n1219) );
NAND3_X1 U898 ( .A1(n1036), .A2(n1169), .A3(n1208), .ZN(n1176) );
AND3_X1 U899 ( .A1(n1158), .A2(n1172), .A3(n1028), .ZN(n1208) );
NOR2_X1 U900 ( .A1(n1220), .A2(n1025), .ZN(n1028) );
NOR2_X1 U901 ( .A1(n1012), .A2(n1193), .ZN(n1169) );
INV_X1 U902 ( .A(n1014), .ZN(n1193) );
AND2_X1 U903 ( .A1(n1211), .A2(n1210), .ZN(n1036) );
INV_X1 U904 ( .A(n1221), .ZN(n1211) );
XNOR2_X1 U905 ( .A(G113), .B(KEYINPUT46), .ZN(n1218) );
XNOR2_X1 U906 ( .A(n1222), .B(n1223), .ZN(G12) );
NOR2_X1 U907 ( .A1(n1224), .A2(n1168), .ZN(n1223) );
NAND4_X1 U908 ( .A1(n1008), .A2(n1158), .A3(n1027), .A4(n1172), .ZN(n1168) );
NAND2_X1 U909 ( .A1(n1037), .A2(n1225), .ZN(n1172) );
NAND3_X1 U910 ( .A1(n1098), .A2(n1207), .A3(G902), .ZN(n1225) );
NOR2_X1 U911 ( .A1(n1079), .A2(G898), .ZN(n1098) );
NAND3_X1 U912 ( .A1(n1207), .A2(n1079), .A3(G952), .ZN(n1037) );
NAND2_X1 U913 ( .A1(G237), .A2(G234), .ZN(n1207) );
NOR2_X1 U914 ( .A1(n1025), .A2(n1026), .ZN(n1027) );
INV_X1 U915 ( .A(n1220), .ZN(n1026) );
NAND2_X1 U916 ( .A1(n1226), .A2(n1047), .ZN(n1220) );
NAND2_X1 U917 ( .A1(G469), .A2(n1227), .ZN(n1047) );
OR2_X1 U918 ( .A1(n1228), .A2(G902), .ZN(n1227) );
XNOR2_X1 U919 ( .A(n1058), .B(KEYINPUT10), .ZN(n1226) );
NOR3_X1 U920 ( .A1(G469), .A2(G902), .A3(n1228), .ZN(n1058) );
XOR2_X1 U921 ( .A(n1229), .B(n1230), .Z(n1228) );
NOR2_X1 U922 ( .A1(KEYINPUT48), .A2(n1231), .ZN(n1230) );
INV_X1 U923 ( .A(n1142), .ZN(n1231) );
XNOR2_X1 U924 ( .A(n1232), .B(n1233), .ZN(n1142) );
XNOR2_X1 U925 ( .A(n1074), .B(G110), .ZN(n1233) );
NAND2_X1 U926 ( .A1(G227), .A2(n1079), .ZN(n1232) );
NAND2_X1 U927 ( .A1(n1234), .A2(n1235), .ZN(n1229) );
NAND2_X1 U928 ( .A1(n1236), .A2(n1131), .ZN(n1235) );
XOR2_X1 U929 ( .A(KEYINPUT40), .B(n1237), .Z(n1234) );
NOR2_X1 U930 ( .A1(n1236), .A2(n1131), .ZN(n1237) );
AND3_X1 U931 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1236) );
NAND2_X1 U932 ( .A1(n1076), .A2(n1241), .ZN(n1240) );
NAND2_X1 U933 ( .A1(n1242), .A2(KEYINPUT25), .ZN(n1241) );
XNOR2_X1 U934 ( .A(n1137), .B(KEYINPUT2), .ZN(n1242) );
NAND3_X1 U935 ( .A1(KEYINPUT25), .A2(n1138), .A3(n1137), .ZN(n1239) );
INV_X1 U936 ( .A(n1076), .ZN(n1138) );
XOR2_X1 U937 ( .A(n1243), .B(n1244), .Z(n1076) );
OR2_X1 U938 ( .A1(n1137), .A2(KEYINPUT25), .ZN(n1238) );
AND2_X1 U939 ( .A1(G221), .A2(n1245), .ZN(n1025) );
NOR2_X1 U940 ( .A1(n1033), .A2(n1032), .ZN(n1158) );
INV_X1 U941 ( .A(n1192), .ZN(n1032) );
NAND2_X1 U942 ( .A1(G214), .A2(n1246), .ZN(n1192) );
XNOR2_X1 U943 ( .A(n1247), .B(n1060), .ZN(n1033) );
AND2_X1 U944 ( .A1(n1248), .A2(G210), .ZN(n1060) );
XOR2_X1 U945 ( .A(n1246), .B(KEYINPUT3), .Z(n1248) );
NAND2_X1 U946 ( .A1(n1249), .A2(n1250), .ZN(n1246) );
XOR2_X1 U947 ( .A(n1062), .B(KEYINPUT13), .Z(n1247) );
NAND2_X1 U948 ( .A1(n1251), .A2(n1250), .ZN(n1062) );
XOR2_X1 U949 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U950 ( .A(n1254), .B(n1147), .Z(n1253) );
XNOR2_X1 U951 ( .A(n1255), .B(n1129), .ZN(n1147) );
INV_X1 U952 ( .A(n1132), .ZN(n1129) );
XOR2_X1 U953 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U954 ( .A1(G953), .A2(n1089), .ZN(n1257) );
INV_X1 U955 ( .A(G224), .ZN(n1089) );
NAND3_X1 U956 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1256) );
OR2_X1 U957 ( .A1(n1099), .A2(KEYINPUT47), .ZN(n1260) );
NAND3_X1 U958 ( .A1(KEYINPUT47), .A2(n1099), .A3(n1261), .ZN(n1259) );
NAND2_X1 U959 ( .A1(n1100), .A2(n1262), .ZN(n1258) );
NAND2_X1 U960 ( .A1(KEYINPUT47), .A2(n1263), .ZN(n1262) );
XOR2_X1 U961 ( .A(KEYINPUT43), .B(n1099), .Z(n1263) );
XOR2_X1 U962 ( .A(n1137), .B(n1264), .Z(n1099) );
XNOR2_X1 U963 ( .A(n1265), .B(n1266), .ZN(n1264) );
NAND2_X1 U964 ( .A1(KEYINPUT18), .A2(n1267), .ZN(n1265) );
XOR2_X1 U965 ( .A(G101), .B(n1268), .Z(n1137) );
XNOR2_X1 U966 ( .A(n1269), .B(G104), .ZN(n1268) );
INV_X1 U967 ( .A(G107), .ZN(n1269) );
INV_X1 U968 ( .A(n1261), .ZN(n1100) );
XOR2_X1 U969 ( .A(G110), .B(n1270), .Z(n1261) );
NAND2_X1 U970 ( .A1(KEYINPUT27), .A2(n1177), .ZN(n1254) );
XNOR2_X1 U971 ( .A(KEYINPUT60), .B(KEYINPUT21), .ZN(n1252) );
NOR2_X1 U972 ( .A1(n1221), .A2(n1210), .ZN(n1008) );
NAND3_X1 U973 ( .A1(n1271), .A2(n1272), .A3(n1051), .ZN(n1210) );
NAND2_X1 U974 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U975 ( .A1(n1053), .A2(n1273), .ZN(n1272) );
OR3_X1 U976 ( .A1(n1053), .A2(n1052), .A3(n1273), .ZN(n1271) );
INV_X1 U977 ( .A(KEYINPUT9), .ZN(n1273) );
NOR2_X1 U978 ( .A1(n1111), .A2(G902), .ZN(n1052) );
XOR2_X1 U979 ( .A(n1274), .B(n1275), .Z(n1111) );
XOR2_X1 U980 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U981 ( .A(n1278), .B(n1279), .ZN(n1277) );
NOR2_X1 U982 ( .A1(G125), .A2(KEYINPUT20), .ZN(n1279) );
NOR2_X1 U983 ( .A1(KEYINPUT61), .A2(n1280), .ZN(n1278) );
XOR2_X1 U984 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U985 ( .A(G143), .B(n1189), .ZN(n1282) );
INV_X1 U986 ( .A(G131), .ZN(n1189) );
NAND3_X1 U987 ( .A1(n1283), .A2(n1249), .A3(G214), .ZN(n1281) );
XNOR2_X1 U988 ( .A(KEYINPUT33), .B(n1079), .ZN(n1283) );
XNOR2_X1 U989 ( .A(G104), .B(KEYINPUT1), .ZN(n1276) );
XNOR2_X1 U990 ( .A(n1270), .B(n1284), .ZN(n1274) );
XNOR2_X1 U991 ( .A(n1285), .B(n1286), .ZN(n1284) );
INV_X1 U992 ( .A(n1266), .ZN(n1285) );
INV_X1 U993 ( .A(G475), .ZN(n1053) );
NAND2_X1 U994 ( .A1(n1039), .A2(n1057), .ZN(n1221) );
NAND3_X1 U995 ( .A1(n1287), .A2(n1250), .A3(n1109), .ZN(n1057) );
INV_X1 U996 ( .A(G478), .ZN(n1287) );
NAND2_X1 U997 ( .A1(G478), .A2(n1288), .ZN(n1039) );
NAND2_X1 U998 ( .A1(n1109), .A2(n1250), .ZN(n1288) );
XOR2_X1 U999 ( .A(n1289), .B(n1290), .Z(n1109) );
XNOR2_X1 U1000 ( .A(n1291), .B(n1270), .ZN(n1290) );
XOR2_X1 U1001 ( .A(G122), .B(KEYINPUT58), .Z(n1270) );
NAND2_X1 U1002 ( .A1(G217), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1003 ( .A(n1293), .B(n1294), .Z(n1289) );
NOR2_X1 U1004 ( .A1(KEYINPUT12), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1005 ( .A(G128), .B(n1296), .Z(n1295) );
XOR2_X1 U1006 ( .A(G143), .B(G134), .Z(n1296) );
XNOR2_X1 U1007 ( .A(G107), .B(G116), .ZN(n1293) );
XNOR2_X1 U1008 ( .A(n1170), .B(KEYINPUT22), .ZN(n1224) );
NOR2_X1 U1009 ( .A1(n1014), .A2(n1194), .ZN(n1170) );
INV_X1 U1010 ( .A(n1012), .ZN(n1194) );
XNOR2_X1 U1011 ( .A(n1046), .B(n1297), .ZN(n1012) );
NOR2_X1 U1012 ( .A1(G472), .A2(KEYINPUT30), .ZN(n1297) );
NAND2_X1 U1013 ( .A1(n1298), .A2(n1250), .ZN(n1046) );
XOR2_X1 U1014 ( .A(n1119), .B(n1299), .Z(n1298) );
XOR2_X1 U1015 ( .A(n1300), .B(n1301), .Z(n1299) );
NOR2_X1 U1016 ( .A1(KEYINPUT6), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1017 ( .A(n1123), .B(G101), .Z(n1302) );
NAND3_X1 U1018 ( .A1(n1249), .A2(n1079), .A3(G210), .ZN(n1123) );
INV_X1 U1019 ( .A(G237), .ZN(n1249) );
NAND3_X1 U1020 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1300) );
OR2_X1 U1021 ( .A1(n1131), .A2(KEYINPUT37), .ZN(n1305) );
INV_X1 U1022 ( .A(n1133), .ZN(n1131) );
NAND3_X1 U1023 ( .A1(KEYINPUT37), .A2(n1306), .A3(n1132), .ZN(n1304) );
OR2_X1 U1024 ( .A1(n1132), .A2(n1306), .ZN(n1303) );
NOR2_X1 U1025 ( .A1(KEYINPUT23), .A2(n1133), .ZN(n1306) );
XNOR2_X1 U1026 ( .A(n1075), .B(KEYINPUT38), .ZN(n1133) );
XNOR2_X1 U1027 ( .A(G131), .B(n1307), .ZN(n1075) );
XNOR2_X1 U1028 ( .A(n1308), .B(G134), .ZN(n1307) );
XOR2_X1 U1029 ( .A(n1309), .B(n1310), .Z(n1132) );
INV_X1 U1030 ( .A(n1243), .ZN(n1310) );
XOR2_X1 U1031 ( .A(G146), .B(G143), .Z(n1243) );
NAND2_X1 U1032 ( .A1(KEYINPUT28), .A2(n1244), .ZN(n1309) );
XNOR2_X1 U1033 ( .A(G128), .B(KEYINPUT50), .ZN(n1244) );
XNOR2_X1 U1034 ( .A(n1266), .B(n1267), .ZN(n1119) );
XOR2_X1 U1035 ( .A(G116), .B(G119), .Z(n1267) );
XOR2_X1 U1036 ( .A(G113), .B(KEYINPUT54), .Z(n1266) );
XNOR2_X1 U1037 ( .A(n1056), .B(KEYINPUT0), .ZN(n1014) );
XOR2_X1 U1038 ( .A(n1311), .B(n1106), .Z(n1056) );
AND2_X1 U1039 ( .A1(G217), .A2(n1245), .ZN(n1106) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1250), .ZN(n1245) );
NAND2_X1 U1041 ( .A1(n1104), .A2(n1250), .ZN(n1311) );
INV_X1 U1042 ( .A(G902), .ZN(n1250) );
XNOR2_X1 U1043 ( .A(n1312), .B(n1313), .ZN(n1104) );
XNOR2_X1 U1044 ( .A(n1314), .B(n1286), .ZN(n1313) );
XNOR2_X1 U1045 ( .A(G146), .B(n1074), .ZN(n1286) );
INV_X1 U1046 ( .A(G140), .ZN(n1074) );
NAND3_X1 U1047 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1314) );
NAND2_X1 U1048 ( .A1(KEYINPUT32), .A2(n1318), .ZN(n1317) );
NAND3_X1 U1049 ( .A1(n1319), .A2(n1320), .A3(G110), .ZN(n1316) );
NAND2_X1 U1050 ( .A1(n1321), .A2(n1222), .ZN(n1315) );
NAND2_X1 U1051 ( .A1(n1322), .A2(n1320), .ZN(n1321) );
INV_X1 U1052 ( .A(KEYINPUT32), .ZN(n1320) );
XNOR2_X1 U1053 ( .A(KEYINPUT5), .B(n1318), .ZN(n1322) );
INV_X1 U1054 ( .A(n1319), .ZN(n1318) );
XOR2_X1 U1055 ( .A(G119), .B(n1323), .Z(n1319) );
XOR2_X1 U1056 ( .A(KEYINPUT36), .B(G128), .Z(n1323) );
XNOR2_X1 U1057 ( .A(n1324), .B(n1177), .ZN(n1312) );
INV_X1 U1058 ( .A(G125), .ZN(n1177) );
NAND2_X1 U1059 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1060 ( .A1(n1308), .A2(n1327), .ZN(n1326) );
NAND2_X1 U1061 ( .A1(G221), .A2(n1292), .ZN(n1327) );
INV_X1 U1062 ( .A(G137), .ZN(n1308) );
XOR2_X1 U1063 ( .A(n1328), .B(KEYINPUT53), .Z(n1325) );
NAND3_X1 U1064 ( .A1(G137), .A2(n1292), .A3(G221), .ZN(n1328) );
AND2_X1 U1065 ( .A1(G234), .A2(n1079), .ZN(n1292) );
INV_X1 U1066 ( .A(G953), .ZN(n1079) );
INV_X1 U1067 ( .A(G110), .ZN(n1222) );
endmodule


