//Key = 1001100111011010100101000100010111000001101000101110110101001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345;

XOR2_X1 U733 ( .A(n1021), .B(n1022), .Z(G9) );
NOR2_X1 U734 ( .A1(G107), .A2(KEYINPUT43), .ZN(n1022) );
NOR2_X1 U735 ( .A1(n1023), .A2(n1024), .ZN(G75) );
NOR2_X1 U736 ( .A1(G952), .A2(n1025), .ZN(n1024) );
NOR4_X1 U737 ( .A1(n1026), .A2(n1027), .A3(n1025), .A4(n1028), .ZN(n1023) );
NAND2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(n1025) );
NAND4_X1 U739 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NOR4_X1 U740 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1034) );
XOR2_X1 U741 ( .A(n1039), .B(n1040), .Z(n1036) );
NOR2_X1 U742 ( .A1(G469), .A2(n1041), .ZN(n1040) );
XOR2_X1 U743 ( .A(KEYINPUT44), .B(KEYINPUT10), .Z(n1041) );
XOR2_X1 U744 ( .A(n1042), .B(n1043), .Z(n1033) );
NAND2_X1 U745 ( .A1(KEYINPUT48), .A2(n1044), .ZN(n1042) );
XNOR2_X1 U746 ( .A(n1045), .B(KEYINPUT56), .ZN(n1031) );
NOR2_X1 U747 ( .A1(n1046), .A2(n1047), .ZN(n1027) );
INV_X1 U748 ( .A(n1032), .ZN(n1047) );
NOR3_X1 U749 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1046) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
AND2_X1 U752 ( .A1(n1055), .A2(n1035), .ZN(n1053) );
NOR3_X1 U753 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1049) );
NOR2_X1 U754 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NOR2_X1 U755 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U756 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U757 ( .A1(n1065), .A2(n1066), .ZN(n1059) );
NOR2_X1 U758 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U759 ( .A1(KEYINPUT51), .A2(n1069), .ZN(n1067) );
NOR2_X1 U760 ( .A1(n1070), .A2(n1071), .ZN(n1048) );
INV_X1 U761 ( .A(KEYINPUT51), .ZN(n1071) );
NOR4_X1 U762 ( .A1(n1066), .A2(n1069), .A3(n1058), .A4(n1056), .ZN(n1070) );
INV_X1 U763 ( .A(n1072), .ZN(n1069) );
NOR3_X1 U764 ( .A1(n1052), .A2(n1073), .A3(n1058), .ZN(n1026) );
NOR2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
OR3_X1 U767 ( .A1(n1062), .A2(n1066), .A3(n1056), .ZN(n1052) );
INV_X1 U768 ( .A(n1078), .ZN(n1062) );
NAND2_X1 U769 ( .A1(n1079), .A2(n1080), .ZN(G72) );
NAND3_X1 U770 ( .A1(n1081), .A2(n1082), .A3(G953), .ZN(n1080) );
NAND2_X1 U771 ( .A1(G900), .A2(G227), .ZN(n1081) );
XOR2_X1 U772 ( .A(n1083), .B(KEYINPUT20), .Z(n1079) );
NAND3_X1 U773 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
OR2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U775 ( .A1(n1088), .A2(n1087), .A3(n1029), .ZN(n1085) );
NAND2_X1 U776 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
XOR2_X1 U777 ( .A(KEYINPUT27), .B(n1091), .Z(n1090) );
NAND2_X1 U778 ( .A1(G953), .A2(n1092), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1088), .A2(G227), .ZN(n1092) );
INV_X1 U780 ( .A(n1082), .ZN(n1088) );
NAND2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(n1082) );
NAND2_X1 U782 ( .A1(G953), .A2(n1095), .ZN(n1094) );
XOR2_X1 U783 ( .A(n1096), .B(n1097), .Z(n1093) );
XOR2_X1 U784 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U785 ( .A(n1100), .B(KEYINPUT0), .Z(n1096) );
NAND2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U788 ( .A1(KEYINPUT33), .A2(n1105), .ZN(n1104) );
NAND2_X1 U789 ( .A1(G131), .A2(n1106), .ZN(n1105) );
INV_X1 U790 ( .A(n1107), .ZN(n1103) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1101) );
NAND2_X1 U792 ( .A1(n1106), .A2(n1110), .ZN(n1108) );
NAND2_X1 U793 ( .A1(KEYINPUT33), .A2(n1107), .ZN(n1110) );
INV_X1 U794 ( .A(KEYINPUT24), .ZN(n1106) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(G69) );
XOR2_X1 U796 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U797 ( .A1(n1115), .A2(n1029), .ZN(n1114) );
NOR2_X1 U798 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U799 ( .A1(n1118), .A2(n1119), .ZN(n1113) );
NAND2_X1 U800 ( .A1(G953), .A2(n1117), .ZN(n1119) );
XNOR2_X1 U801 ( .A(n1120), .B(n1121), .ZN(n1118) );
NAND3_X1 U802 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1120) );
NAND2_X1 U803 ( .A1(KEYINPUT28), .A2(n1125), .ZN(n1124) );
OR3_X1 U804 ( .A1(n1125), .A2(KEYINPUT28), .A3(n1126), .ZN(n1123) );
NAND2_X1 U805 ( .A1(n1126), .A2(n1127), .ZN(n1122) );
NAND2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
INV_X1 U807 ( .A(KEYINPUT28), .ZN(n1129) );
XNOR2_X1 U808 ( .A(KEYINPUT16), .B(n1130), .ZN(n1128) );
NAND2_X1 U809 ( .A1(n1029), .A2(n1131), .ZN(n1111) );
NOR2_X1 U810 ( .A1(n1132), .A2(n1133), .ZN(G66) );
NOR3_X1 U811 ( .A1(n1043), .A2(n1134), .A3(n1135), .ZN(n1133) );
AND3_X1 U812 ( .A1(n1136), .A2(n1044), .A3(n1137), .ZN(n1135) );
NOR2_X1 U813 ( .A1(n1138), .A2(n1136), .ZN(n1134) );
AND2_X1 U814 ( .A1(n1028), .A2(n1044), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1132), .A2(n1139), .ZN(G63) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U817 ( .A1(n1137), .A2(G478), .ZN(n1140) );
NOR2_X1 U818 ( .A1(n1132), .A2(n1142), .ZN(G60) );
XOR2_X1 U819 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U820 ( .A1(n1137), .A2(G475), .ZN(n1143) );
XNOR2_X1 U821 ( .A(G104), .B(n1145), .ZN(G6) );
NOR2_X1 U822 ( .A1(n1132), .A2(n1146), .ZN(G57) );
XOR2_X1 U823 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U824 ( .A(n1149), .B(n1125), .ZN(n1148) );
NAND2_X1 U825 ( .A1(n1137), .A2(G472), .ZN(n1149) );
XOR2_X1 U826 ( .A(n1150), .B(n1151), .Z(n1147) );
NOR2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XNOR2_X1 U828 ( .A(n1154), .B(KEYINPUT25), .ZN(n1153) );
NOR2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
NOR2_X1 U830 ( .A1(KEYINPUT36), .A2(n1157), .ZN(n1150) );
NOR2_X1 U831 ( .A1(n1132), .A2(n1158), .ZN(G54) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U833 ( .A(KEYINPUT34), .B(n1161), .Z(n1160) );
NOR2_X1 U834 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
AND2_X1 U835 ( .A1(n1163), .A2(n1162), .ZN(n1159) );
XNOR2_X1 U836 ( .A(n1164), .B(n1165), .ZN(n1162) );
XNOR2_X1 U837 ( .A(n1166), .B(n1167), .ZN(n1165) );
XNOR2_X1 U838 ( .A(n1168), .B(n1169), .ZN(n1164) );
XNOR2_X1 U839 ( .A(n1170), .B(n1171), .ZN(n1168) );
NOR2_X1 U840 ( .A1(KEYINPUT2), .A2(n1172), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1137), .A2(G469), .ZN(n1163) );
INV_X1 U842 ( .A(n1173), .ZN(n1137) );
NOR2_X1 U843 ( .A1(n1132), .A2(n1174), .ZN(G51) );
XOR2_X1 U844 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U845 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR2_X1 U846 ( .A1(G953), .A2(n1116), .ZN(n1178) );
NAND3_X1 U847 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1177) );
NAND2_X1 U848 ( .A1(KEYINPUT41), .A2(n1182), .ZN(n1181) );
OR3_X1 U849 ( .A1(n1183), .A2(KEYINPUT41), .A3(G125), .ZN(n1180) );
NAND2_X1 U850 ( .A1(G125), .A2(n1183), .ZN(n1179) );
NAND2_X1 U851 ( .A1(KEYINPUT63), .A2(n1184), .ZN(n1183) );
XOR2_X1 U852 ( .A(n1185), .B(n1186), .Z(n1175) );
NOR3_X1 U853 ( .A1(n1173), .A2(KEYINPUT23), .A3(n1187), .ZN(n1186) );
NAND2_X1 U854 ( .A1(G902), .A2(n1028), .ZN(n1173) );
NAND3_X1 U855 ( .A1(n1091), .A2(n1089), .A3(n1188), .ZN(n1028) );
INV_X1 U856 ( .A(n1131), .ZN(n1188) );
NAND4_X1 U857 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1131) );
AND4_X1 U858 ( .A1(n1021), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1192) );
NAND3_X1 U859 ( .A1(n1072), .A2(n1196), .A3(n1197), .ZN(n1021) );
AND2_X1 U860 ( .A1(n1198), .A2(n1145), .ZN(n1191) );
NAND3_X1 U861 ( .A1(n1197), .A2(n1196), .A3(n1068), .ZN(n1145) );
AND4_X1 U862 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1089) );
NAND3_X1 U863 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1200) );
XNOR2_X1 U864 ( .A(n1075), .B(KEYINPUT29), .ZN(n1205) );
NAND2_X1 U865 ( .A1(n1206), .A2(n1032), .ZN(n1199) );
XNOR2_X1 U866 ( .A(n1207), .B(KEYINPUT50), .ZN(n1206) );
AND3_X1 U867 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1091) );
NAND2_X1 U868 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND2_X1 U869 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND3_X1 U870 ( .A1(n1215), .A2(n1045), .A3(n1064), .ZN(n1214) );
NAND2_X1 U871 ( .A1(n1216), .A2(n1068), .ZN(n1213) );
NOR2_X1 U872 ( .A1(n1029), .A2(G952), .ZN(n1132) );
XNOR2_X1 U873 ( .A(G146), .B(n1217), .ZN(G48) );
NAND4_X1 U874 ( .A1(KEYINPUT49), .A2(n1211), .A3(n1068), .A4(n1218), .ZN(n1217) );
XOR2_X1 U875 ( .A(KEYINPUT22), .B(n1216), .Z(n1218) );
XNOR2_X1 U876 ( .A(G143), .B(n1219), .ZN(G45) );
NAND3_X1 U877 ( .A1(KEYINPUT52), .A2(n1211), .A3(n1220), .ZN(n1219) );
NOR3_X1 U878 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1220) );
XNOR2_X1 U879 ( .A(G140), .B(n1208), .ZN(G42) );
NAND3_X1 U880 ( .A1(n1068), .A2(n1063), .A3(n1224), .ZN(n1208) );
XNOR2_X1 U881 ( .A(G137), .B(n1209), .ZN(G39) );
NAND3_X1 U882 ( .A1(n1216), .A2(n1078), .A3(n1224), .ZN(n1209) );
XNOR2_X1 U883 ( .A(G134), .B(n1201), .ZN(G36) );
NAND3_X1 U884 ( .A1(n1064), .A2(n1072), .A3(n1224), .ZN(n1201) );
AND2_X1 U885 ( .A1(n1204), .A2(n1032), .ZN(n1224) );
XOR2_X1 U886 ( .A(n1225), .B(n1226), .Z(G33) );
XNOR2_X1 U887 ( .A(G131), .B(KEYINPUT35), .ZN(n1226) );
NAND2_X1 U888 ( .A1(n1207), .A2(n1032), .ZN(n1225) );
NOR2_X1 U889 ( .A1(n1076), .A2(n1227), .ZN(n1032) );
AND3_X1 U890 ( .A1(n1068), .A2(n1064), .A3(n1204), .ZN(n1207) );
XOR2_X1 U891 ( .A(n1228), .B(n1229), .Z(G30) );
NOR2_X1 U892 ( .A1(KEYINPUT54), .A2(G128), .ZN(n1229) );
NAND2_X1 U893 ( .A1(n1203), .A2(n1211), .ZN(n1228) );
AND2_X1 U894 ( .A1(n1204), .A2(n1075), .ZN(n1211) );
AND2_X1 U895 ( .A1(n1054), .A2(n1230), .ZN(n1204) );
AND2_X1 U896 ( .A1(n1216), .A2(n1072), .ZN(n1203) );
XNOR2_X1 U897 ( .A(G101), .B(n1198), .ZN(G3) );
NAND3_X1 U898 ( .A1(n1078), .A2(n1197), .A3(n1064), .ZN(n1198) );
XNOR2_X1 U899 ( .A(n1202), .B(n1231), .ZN(G27) );
NOR2_X1 U900 ( .A1(KEYINPUT37), .A2(n1232), .ZN(n1231) );
INV_X1 U901 ( .A(G125), .ZN(n1232) );
NAND4_X1 U902 ( .A1(n1068), .A2(n1233), .A3(n1234), .A4(n1063), .ZN(n1202) );
AND2_X1 U903 ( .A1(n1230), .A2(n1075), .ZN(n1234) );
NAND2_X1 U904 ( .A1(n1056), .A2(n1235), .ZN(n1230) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1095), .ZN(n1235) );
INV_X1 U906 ( .A(G900), .ZN(n1095) );
XNOR2_X1 U907 ( .A(G122), .B(n1189), .ZN(G24) );
NAND4_X1 U908 ( .A1(n1237), .A2(n1196), .A3(n1215), .A4(n1045), .ZN(n1189) );
INV_X1 U909 ( .A(n1066), .ZN(n1196) );
NAND2_X1 U910 ( .A1(n1238), .A2(n1239), .ZN(n1066) );
XNOR2_X1 U911 ( .A(n1240), .B(KEYINPUT61), .ZN(n1238) );
XNOR2_X1 U912 ( .A(G119), .B(n1190), .ZN(G21) );
NAND3_X1 U913 ( .A1(n1237), .A2(n1078), .A3(n1216), .ZN(n1190) );
NOR2_X1 U914 ( .A1(n1241), .A2(n1239), .ZN(n1216) );
INV_X1 U915 ( .A(n1240), .ZN(n1241) );
NAND2_X1 U916 ( .A1(n1242), .A2(n1243), .ZN(G18) );
NAND2_X1 U917 ( .A1(G116), .A2(n1195), .ZN(n1243) );
XOR2_X1 U918 ( .A(KEYINPUT39), .B(n1244), .Z(n1242) );
NOR2_X1 U919 ( .A1(G116), .A2(n1195), .ZN(n1244) );
NAND3_X1 U920 ( .A1(n1237), .A2(n1072), .A3(n1064), .ZN(n1195) );
NOR2_X1 U921 ( .A1(n1223), .A2(n1045), .ZN(n1072) );
XNOR2_X1 U922 ( .A(G113), .B(n1194), .ZN(G15) );
NAND3_X1 U923 ( .A1(n1064), .A2(n1237), .A3(n1068), .ZN(n1194) );
NOR2_X1 U924 ( .A1(n1222), .A2(n1215), .ZN(n1068) );
INV_X1 U925 ( .A(n1045), .ZN(n1222) );
AND2_X1 U926 ( .A1(n1233), .A2(n1245), .ZN(n1237) );
INV_X1 U927 ( .A(n1058), .ZN(n1233) );
NAND2_X1 U928 ( .A1(n1055), .A2(n1246), .ZN(n1058) );
INV_X1 U929 ( .A(n1221), .ZN(n1064) );
NAND2_X1 U930 ( .A1(n1239), .A2(n1240), .ZN(n1221) );
NAND2_X1 U931 ( .A1(n1247), .A2(n1248), .ZN(G12) );
NAND2_X1 U932 ( .A1(G110), .A2(n1193), .ZN(n1248) );
XOR2_X1 U933 ( .A(KEYINPUT46), .B(n1249), .Z(n1247) );
NOR2_X1 U934 ( .A1(G110), .A2(n1193), .ZN(n1249) );
NAND3_X1 U935 ( .A1(n1063), .A2(n1197), .A3(n1078), .ZN(n1193) );
NOR2_X1 U936 ( .A1(n1045), .A2(n1215), .ZN(n1078) );
INV_X1 U937 ( .A(n1223), .ZN(n1215) );
XOR2_X1 U938 ( .A(n1038), .B(KEYINPUT12), .Z(n1223) );
XNOR2_X1 U939 ( .A(n1250), .B(n1251), .ZN(n1038) );
XOR2_X1 U940 ( .A(KEYINPUT1), .B(G478), .Z(n1251) );
NAND2_X1 U941 ( .A1(n1141), .A2(n1252), .ZN(n1250) );
XOR2_X1 U942 ( .A(n1253), .B(n1254), .Z(n1141) );
NOR3_X1 U943 ( .A1(n1255), .A2(G953), .A3(n1256), .ZN(n1254) );
INV_X1 U944 ( .A(G234), .ZN(n1256) );
XOR2_X1 U945 ( .A(KEYINPUT4), .B(G217), .Z(n1255) );
NAND3_X1 U946 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1253) );
OR2_X1 U947 ( .A1(n1260), .A2(KEYINPUT7), .ZN(n1259) );
NAND3_X1 U948 ( .A1(KEYINPUT7), .A2(n1260), .A3(n1261), .ZN(n1258) );
NAND2_X1 U949 ( .A1(n1262), .A2(n1263), .ZN(n1257) );
NAND2_X1 U950 ( .A1(n1264), .A2(KEYINPUT7), .ZN(n1263) );
XNOR2_X1 U951 ( .A(n1260), .B(KEYINPUT3), .ZN(n1264) );
XNOR2_X1 U952 ( .A(n1265), .B(n1266), .ZN(n1260) );
XOR2_X1 U953 ( .A(G122), .B(G116), .Z(n1266) );
NAND2_X1 U954 ( .A1(KEYINPUT55), .A2(n1267), .ZN(n1265) );
INV_X1 U955 ( .A(n1261), .ZN(n1262) );
XOR2_X1 U956 ( .A(G134), .B(n1268), .Z(n1261) );
XNOR2_X1 U957 ( .A(n1269), .B(G475), .ZN(n1045) );
NAND2_X1 U958 ( .A1(n1144), .A2(n1252), .ZN(n1269) );
XOR2_X1 U959 ( .A(n1270), .B(n1271), .Z(n1144) );
XOR2_X1 U960 ( .A(G104), .B(n1272), .Z(n1271) );
XNOR2_X1 U961 ( .A(KEYINPUT60), .B(n1273), .ZN(n1272) );
XOR2_X1 U962 ( .A(n1274), .B(n1275), .Z(n1270) );
XNOR2_X1 U963 ( .A(n1276), .B(n1277), .ZN(n1275) );
NOR2_X1 U964 ( .A1(KEYINPUT13), .A2(n1278), .ZN(n1277) );
XOR2_X1 U965 ( .A(n1279), .B(n1280), .Z(n1278) );
XNOR2_X1 U966 ( .A(n1109), .B(n1281), .ZN(n1280) );
NOR3_X1 U967 ( .A1(n1282), .A2(G237), .A3(n1283), .ZN(n1281) );
XNOR2_X1 U968 ( .A(KEYINPUT5), .B(n1029), .ZN(n1282) );
XNOR2_X1 U969 ( .A(KEYINPUT53), .B(n1284), .ZN(n1279) );
NAND2_X1 U970 ( .A1(KEYINPUT57), .A2(n1285), .ZN(n1276) );
XOR2_X1 U971 ( .A(G122), .B(G113), .Z(n1285) );
AND2_X1 U972 ( .A1(n1245), .A2(n1054), .ZN(n1197) );
NOR2_X1 U973 ( .A1(n1055), .A2(n1035), .ZN(n1054) );
INV_X1 U974 ( .A(n1246), .ZN(n1035) );
NAND2_X1 U975 ( .A1(G221), .A2(n1286), .ZN(n1246) );
XOR2_X1 U976 ( .A(n1039), .B(G469), .Z(n1055) );
NAND2_X1 U977 ( .A1(n1287), .A2(n1252), .ZN(n1039) );
XOR2_X1 U978 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U979 ( .A(n1170), .B(n1166), .ZN(n1289) );
XNOR2_X1 U980 ( .A(n1290), .B(n1172), .ZN(n1288) );
NAND2_X1 U981 ( .A1(G227), .A2(n1029), .ZN(n1172) );
XNOR2_X1 U982 ( .A(n1291), .B(n1292), .ZN(n1290) );
NAND2_X1 U983 ( .A1(KEYINPUT42), .A2(n1167), .ZN(n1292) );
XNOR2_X1 U984 ( .A(n1126), .B(n1099), .ZN(n1167) );
XNOR2_X1 U985 ( .A(n1273), .B(n1268), .ZN(n1099) );
XOR2_X1 U986 ( .A(G128), .B(G143), .Z(n1268) );
NAND2_X1 U987 ( .A1(n1293), .A2(KEYINPUT19), .ZN(n1291) );
XNOR2_X1 U988 ( .A(n1294), .B(KEYINPUT59), .ZN(n1293) );
AND2_X1 U989 ( .A1(n1075), .A2(n1295), .ZN(n1245) );
NAND2_X1 U990 ( .A1(n1056), .A2(n1296), .ZN(n1295) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1117), .ZN(n1296) );
INV_X1 U992 ( .A(G898), .ZN(n1117) );
NAND3_X1 U993 ( .A1(n1236), .A2(n1029), .A3(G952), .ZN(n1056) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1236) );
AND2_X1 U995 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U996 ( .A(n1227), .ZN(n1077) );
NOR2_X1 U997 ( .A1(n1283), .A2(n1297), .ZN(n1227) );
INV_X1 U998 ( .A(G214), .ZN(n1283) );
XNOR2_X1 U999 ( .A(n1298), .B(n1299), .ZN(n1076) );
NOR2_X1 U1000 ( .A1(n1297), .A2(n1187), .ZN(n1299) );
NOR2_X1 U1001 ( .A1(G902), .A2(G237), .ZN(n1297) );
NAND2_X1 U1002 ( .A1(n1300), .A2(n1252), .ZN(n1298) );
XOR2_X1 U1003 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1004 ( .A(n1303), .B(n1304), .Z(n1302) );
NAND2_X1 U1005 ( .A1(KEYINPUT40), .A2(n1116), .ZN(n1304) );
INV_X1 U1006 ( .A(G224), .ZN(n1116) );
NAND2_X1 U1007 ( .A1(KEYINPUT11), .A2(G125), .ZN(n1303) );
XNOR2_X1 U1008 ( .A(n1185), .B(n1182), .ZN(n1301) );
NAND3_X1 U1009 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1185) );
NAND2_X1 U1010 ( .A1(KEYINPUT26), .A2(n1308), .ZN(n1307) );
OR3_X1 U1011 ( .A1(n1308), .A2(KEYINPUT26), .A3(n1121), .ZN(n1306) );
NAND2_X1 U1012 ( .A1(n1121), .A2(n1309), .ZN(n1305) );
NAND2_X1 U1013 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
INV_X1 U1014 ( .A(KEYINPUT26), .ZN(n1311) );
XOR2_X1 U1015 ( .A(KEYINPUT32), .B(n1308), .Z(n1310) );
XNOR2_X1 U1016 ( .A(n1126), .B(n1130), .ZN(n1308) );
XOR2_X1 U1017 ( .A(G101), .B(n1312), .Z(n1126) );
XNOR2_X1 U1018 ( .A(n1267), .B(G104), .ZN(n1312) );
INV_X1 U1019 ( .A(G107), .ZN(n1267) );
XOR2_X1 U1020 ( .A(G122), .B(n1169), .Z(n1121) );
NOR2_X1 U1021 ( .A1(n1240), .A2(n1239), .ZN(n1063) );
XNOR2_X1 U1022 ( .A(n1043), .B(n1044), .ZN(n1239) );
AND2_X1 U1023 ( .A1(G217), .A2(n1286), .ZN(n1044) );
NAND2_X1 U1024 ( .A1(G234), .A2(n1252), .ZN(n1286) );
NOR2_X1 U1025 ( .A1(n1136), .A2(G902), .ZN(n1043) );
XNOR2_X1 U1026 ( .A(n1313), .B(n1314), .ZN(n1136) );
XOR2_X1 U1027 ( .A(n1315), .B(n1316), .Z(n1314) );
AND3_X1 U1028 ( .A1(G221), .A2(n1029), .A3(G234), .ZN(n1315) );
INV_X1 U1029 ( .A(G953), .ZN(n1029) );
XNOR2_X1 U1030 ( .A(KEYINPUT9), .B(n1317), .ZN(n1313) );
NOR2_X1 U1031 ( .A1(KEYINPUT6), .A2(n1318), .ZN(n1317) );
XOR2_X1 U1032 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1033 ( .A(n1321), .B(n1322), .ZN(n1320) );
NOR2_X1 U1034 ( .A1(KEYINPUT62), .A2(n1274), .ZN(n1322) );
XNOR2_X1 U1035 ( .A(n1098), .B(KEYINPUT30), .ZN(n1274) );
XOR2_X1 U1036 ( .A(G125), .B(n1166), .Z(n1098) );
XOR2_X1 U1037 ( .A(G140), .B(KEYINPUT18), .Z(n1166) );
NAND2_X1 U1038 ( .A1(KEYINPUT8), .A2(n1169), .ZN(n1321) );
INV_X1 U1039 ( .A(n1294), .ZN(n1169) );
XOR2_X1 U1040 ( .A(G110), .B(KEYINPUT15), .Z(n1294) );
XOR2_X1 U1041 ( .A(G119), .B(n1323), .Z(n1319) );
XNOR2_X1 U1042 ( .A(n1273), .B(G128), .ZN(n1323) );
XOR2_X1 U1043 ( .A(n1037), .B(KEYINPUT58), .Z(n1240) );
XNOR2_X1 U1044 ( .A(n1324), .B(G472), .ZN(n1037) );
NAND2_X1 U1045 ( .A1(n1325), .A2(n1252), .ZN(n1324) );
INV_X1 U1046 ( .A(G902), .ZN(n1252) );
XNOR2_X1 U1047 ( .A(n1326), .B(n1130), .ZN(n1325) );
INV_X1 U1048 ( .A(n1125), .ZN(n1130) );
XOR2_X1 U1049 ( .A(G113), .B(n1327), .Z(n1125) );
XOR2_X1 U1050 ( .A(G119), .B(G116), .Z(n1327) );
XOR2_X1 U1051 ( .A(n1157), .B(n1328), .Z(n1326) );
NOR2_X1 U1052 ( .A1(n1154), .A2(n1329), .ZN(n1328) );
XOR2_X1 U1053 ( .A(n1330), .B(KEYINPUT21), .Z(n1329) );
NAND2_X1 U1054 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XNOR2_X1 U1055 ( .A(KEYINPUT45), .B(n1155), .ZN(n1332) );
XOR2_X1 U1056 ( .A(n1156), .B(KEYINPUT14), .Z(n1331) );
AND2_X1 U1057 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
OR3_X1 U1058 ( .A1(G237), .A2(G953), .A3(n1187), .ZN(n1156) );
INV_X1 U1059 ( .A(G210), .ZN(n1187) );
INV_X1 U1060 ( .A(G101), .ZN(n1155) );
XNOR2_X1 U1061 ( .A(n1184), .B(n1170), .ZN(n1157) );
XNOR2_X1 U1062 ( .A(n1107), .B(n1109), .ZN(n1170) );
INV_X1 U1063 ( .A(G131), .ZN(n1109) );
XOR2_X1 U1064 ( .A(G134), .B(n1316), .Z(n1107) );
XOR2_X1 U1065 ( .A(G137), .B(KEYINPUT38), .Z(n1316) );
INV_X1 U1066 ( .A(n1182), .ZN(n1184) );
NAND2_X1 U1067 ( .A1(n1333), .A2(n1334), .ZN(n1182) );
NAND3_X1 U1068 ( .A1(n1335), .A2(n1336), .A3(G128), .ZN(n1334) );
NAND2_X1 U1069 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND2_X1 U1070 ( .A1(G143), .A2(n1273), .ZN(n1337) );
NAND2_X1 U1071 ( .A1(n1339), .A2(KEYINPUT31), .ZN(n1335) );
XNOR2_X1 U1072 ( .A(n1273), .B(G143), .ZN(n1339) );
INV_X1 U1073 ( .A(G146), .ZN(n1273) );
NAND2_X1 U1074 ( .A1(n1340), .A2(n1341), .ZN(n1333) );
NAND2_X1 U1075 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1076 ( .A1(G146), .A2(n1284), .ZN(n1343) );
XNOR2_X1 U1077 ( .A(n1338), .B(n1344), .ZN(n1342) );
NOR2_X1 U1078 ( .A1(G146), .A2(n1284), .ZN(n1344) );
INV_X1 U1079 ( .A(G143), .ZN(n1284) );
INV_X1 U1080 ( .A(KEYINPUT31), .ZN(n1338) );
XOR2_X1 U1081 ( .A(n1345), .B(G128), .Z(n1340) );
XNOR2_X1 U1082 ( .A(KEYINPUT47), .B(KEYINPUT17), .ZN(n1345) );
endmodule


