//Key = 0100101001001001000111011010100110011101011110000010101100101000


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
n2287, n2288;

INV_X2 U1280 ( .A(n1885), .ZN(n1857) );
INV_X2 U1281 ( .A(U280), .ZN(n1858) );
INV_X1 U1282 ( .A(n1717), .ZN(U375) );
NAND2_X1 U1283 ( .A1(n1718), .A2(n1719), .ZN(U344) );
NAND2_X1 U1284 ( .A1(n1720), .A2(DATA_IN_7_), .ZN(n1719) );
XOR2_X1 U1285 ( .A(n1721), .B(KEYINPUT41), .Z(n1720) );
NAND2_X1 U1286 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1721), .ZN(n1718) );
NAND2_X1 U1287 ( .A1(n1722), .A2(n1723), .ZN(U343) );
NAND2_X1 U1288 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1721), .ZN(n1723) );
NAND2_X1 U1289 ( .A1(n1724), .A2(DATA_IN_6_), .ZN(n1722) );
NAND2_X1 U1290 ( .A1(n1725), .A2(n1726), .ZN(U342) );
NAND2_X1 U1291 ( .A1(n1727), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1726) );
XOR2_X1 U1292 ( .A(n1721), .B(KEYINPUT27), .Z(n1727) );
NAND2_X1 U1293 ( .A1(n1724), .A2(DATA_IN_5_), .ZN(n1725) );
NAND2_X1 U1294 ( .A1(n1728), .A2(n1729), .ZN(U341) );
NAND2_X1 U1295 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1721), .ZN(n1729) );
NAND2_X1 U1296 ( .A1(n1724), .A2(DATA_IN_4_), .ZN(n1728) );
NAND2_X1 U1297 ( .A1(n1730), .A2(n1731), .ZN(U340) );
NAND2_X1 U1298 ( .A1(n1732), .A2(n1721), .ZN(n1731) );
XOR2_X1 U1299 ( .A(RMAX_REG_3__SCAN_IN), .B(KEYINPUT8), .Z(n1732) );
NAND2_X1 U1300 ( .A1(n1724), .A2(DATA_IN_3_), .ZN(n1730) );
NAND2_X1 U1301 ( .A1(n1733), .A2(n1734), .ZN(U339) );
NAND2_X1 U1302 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1721), .ZN(n1734) );
NAND2_X1 U1303 ( .A1(n1724), .A2(DATA_IN_2_), .ZN(n1733) );
NAND2_X1 U1304 ( .A1(n1735), .A2(n1736), .ZN(U338) );
NAND2_X1 U1305 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1721), .ZN(n1736) );
NAND2_X1 U1306 ( .A1(n1724), .A2(DATA_IN_1_), .ZN(n1735) );
NAND2_X1 U1307 ( .A1(n1737), .A2(n1738), .ZN(U337) );
NAND2_X1 U1308 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1721), .ZN(n1738) );
NAND2_X1 U1309 ( .A1(n1739), .A2(n1724), .ZN(n1737) );
INV_X1 U1310 ( .A(n1721), .ZN(n1724) );
NAND2_X1 U1311 ( .A1(n1717), .A2(n1740), .ZN(n1721) );
NAND3_X1 U1312 ( .A1(n1741), .A2(n1742), .A3(n1743), .ZN(n1740) );
XOR2_X1 U1313 ( .A(n1744), .B(KEYINPUT15), .Z(n1739) );
NAND2_X1 U1314 ( .A1(n1745), .A2(n1746), .ZN(U336) );
NAND2_X1 U1315 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1747), .ZN(n1746) );
NAND2_X1 U1316 ( .A1(n1748), .A2(DATA_IN_7_), .ZN(n1745) );
NAND2_X1 U1317 ( .A1(n1749), .A2(n1750), .ZN(U335) );
NAND2_X1 U1318 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1747), .ZN(n1750) );
NAND2_X1 U1319 ( .A1(n1748), .A2(DATA_IN_6_), .ZN(n1749) );
NAND2_X1 U1320 ( .A1(n1751), .A2(n1752), .ZN(U334) );
NAND2_X1 U1321 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1747), .ZN(n1752) );
NAND2_X1 U1322 ( .A1(n1748), .A2(DATA_IN_5_), .ZN(n1751) );
NAND2_X1 U1323 ( .A1(n1753), .A2(n1754), .ZN(U333) );
NAND2_X1 U1324 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1747), .ZN(n1754) );
NAND2_X1 U1325 ( .A1(n1748), .A2(DATA_IN_4_), .ZN(n1753) );
NAND2_X1 U1326 ( .A1(n1755), .A2(n1756), .ZN(U332) );
NAND2_X1 U1327 ( .A1(n1757), .A2(RMIN_REG_3__SCAN_IN), .ZN(n1756) );
XOR2_X1 U1328 ( .A(n1747), .B(KEYINPUT11), .Z(n1757) );
NAND2_X1 U1329 ( .A1(n1748), .A2(DATA_IN_3_), .ZN(n1755) );
NAND2_X1 U1330 ( .A1(n1758), .A2(n1759), .ZN(U331) );
NAND2_X1 U1331 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1747), .ZN(n1759) );
NAND2_X1 U1332 ( .A1(n1748), .A2(DATA_IN_2_), .ZN(n1758) );
NAND2_X1 U1333 ( .A1(n1760), .A2(n1761), .ZN(U330) );
NAND2_X1 U1334 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1747), .ZN(n1761) );
NAND2_X1 U1335 ( .A1(n1748), .A2(DATA_IN_1_), .ZN(n1760) );
NAND2_X1 U1336 ( .A1(n1762), .A2(n1763), .ZN(U329) );
NAND2_X1 U1337 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1747), .ZN(n1763) );
XOR2_X1 U1338 ( .A(n1764), .B(KEYINPUT30), .Z(n1762) );
NAND2_X1 U1339 ( .A1(n1748), .A2(DATA_IN_0_), .ZN(n1764) );
INV_X1 U1340 ( .A(n1747), .ZN(n1748) );
NAND2_X1 U1341 ( .A1(n1717), .A2(n1765), .ZN(n1747) );
NAND2_X1 U1342 ( .A1(n1766), .A2(n1742), .ZN(n1765) );
NAND3_X1 U1343 ( .A1(n1743), .A2(n1741), .A3(n1767), .ZN(n1766) );
NAND2_X1 U1344 ( .A1(n1768), .A2(n1769), .ZN(n1767) );
NAND3_X1 U1345 ( .A1(n1770), .A2(n1771), .A3(n1772), .ZN(n1769) );
NAND2_X1 U1346 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1773), .ZN(n1772) );
NAND3_X1 U1347 ( .A1(n1774), .A2(n1775), .A3(n1776), .ZN(n1771) );
NAND2_X1 U1348 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1777), .ZN(n1776) );
NAND3_X1 U1349 ( .A1(n1778), .A2(n1779), .A3(n1780), .ZN(n1775) );
NAND2_X1 U1350 ( .A1(DATA_IN_4_), .A2(n1781), .ZN(n1780) );
NAND3_X1 U1351 ( .A1(n1782), .A2(n1783), .A3(n1784), .ZN(n1779) );
NAND2_X1 U1352 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1785), .ZN(n1784) );
NAND3_X1 U1353 ( .A1(n1786), .A2(n1787), .A3(n1788), .ZN(n1783) );
NAND2_X1 U1354 ( .A1(DATA_IN_3_), .A2(n1789), .ZN(n1788) );
NAND3_X1 U1355 ( .A1(n1790), .A2(n1791), .A3(n1792), .ZN(n1787) );
NAND2_X1 U1356 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1793), .ZN(n1792) );
NAND3_X1 U1357 ( .A1(n1794), .A2(n1744), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1791) );
NAND2_X1 U1358 ( .A1(DATA_IN_1_), .A2(n1795), .ZN(n1794) );
NAND2_X1 U1359 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1796), .ZN(n1790) );
NAND2_X1 U1360 ( .A1(DATA_IN_2_), .A2(n1797), .ZN(n1786) );
XOR2_X1 U1361 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT60), .Z(n1797) );
NAND2_X1 U1362 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1798), .ZN(n1782) );
NAND2_X1 U1363 ( .A1(n1799), .A2(n1800), .ZN(n1778) );
XOR2_X1 U1364 ( .A(KEYINPUT16), .B(DATA_IN_5_), .Z(n1799) );
NAND2_X1 U1365 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1801), .ZN(n1774) );
NAND2_X1 U1366 ( .A1(DATA_IN_6_), .A2(n1802), .ZN(n1770) );
NAND2_X1 U1367 ( .A1(DATA_IN_7_), .A2(n1803), .ZN(n1768) );
NAND3_X1 U1368 ( .A1(n1804), .A2(n1805), .A3(n1806), .ZN(n1741) );
NAND2_X1 U1369 ( .A1(DATA_IN_7_), .A2(n1807), .ZN(n1806) );
NAND3_X1 U1370 ( .A1(n1808), .A2(n1809), .A3(n1810), .ZN(n1805) );
NAND2_X1 U1371 ( .A1(DATA_IN_5_), .A2(n1811), .ZN(n1810) );
NAND3_X1 U1372 ( .A1(n1812), .A2(n1813), .A3(n1814), .ZN(n1809) );
NAND2_X1 U1373 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1801), .ZN(n1814) );
NAND3_X1 U1374 ( .A1(n1815), .A2(n1816), .A3(n1817), .ZN(n1813) );
NAND2_X1 U1375 ( .A1(DATA_IN_4_), .A2(n1818), .ZN(n1817) );
NAND3_X1 U1376 ( .A1(n1819), .A2(n1820), .A3(n1821), .ZN(n1816) );
NAND2_X1 U1377 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1798), .ZN(n1821) );
NAND3_X1 U1378 ( .A1(n1822), .A2(n1823), .A3(n1824), .ZN(n1820) );
NAND2_X1 U1379 ( .A1(DATA_IN_2_), .A2(n1825), .ZN(n1824) );
NAND3_X1 U1380 ( .A1(n1826), .A2(n1827), .A3(DATA_IN_0_), .ZN(n1823) );
NAND2_X1 U1381 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1796), .ZN(n1826) );
NAND2_X1 U1382 ( .A1(DATA_IN_1_), .A2(n1828), .ZN(n1822) );
XOR2_X1 U1383 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT43), .Z(n1828) );
NAND2_X1 U1384 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1793), .ZN(n1819) );
NAND2_X1 U1385 ( .A1(DATA_IN_3_), .A2(n1829), .ZN(n1815) );
NAND2_X1 U1386 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1785), .ZN(n1812) );
NAND2_X1 U1387 ( .A1(DATA_IN_6_), .A2(n1830), .ZN(n1808) );
XOR2_X1 U1388 ( .A(RMAX_REG_6__SCAN_IN), .B(KEYINPUT39), .Z(n1830) );
NAND2_X1 U1389 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1777), .ZN(n1804) );
NAND2_X1 U1390 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1773), .ZN(n1743) );
NAND2_X1 U1391 ( .A1(n1831), .A2(n1832), .ZN(U328) );
NAND2_X1 U1392 ( .A1(n1833), .A2(DATA_IN_7_), .ZN(n1832) );
NAND2_X1 U1393 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1834), .ZN(n1831) );
NAND2_X1 U1394 ( .A1(n1835), .A2(n1836), .ZN(U327) );
NAND2_X1 U1395 ( .A1(n1833), .A2(DATA_IN_6_), .ZN(n1836) );
NAND2_X1 U1396 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1834), .ZN(n1835) );
NAND2_X1 U1397 ( .A1(n1837), .A2(n1838), .ZN(U326) );
NAND2_X1 U1398 ( .A1(n1833), .A2(n1839), .ZN(n1838) );
XOR2_X1 U1399 ( .A(KEYINPUT3), .B(DATA_IN_5_), .Z(n1839) );
NAND2_X1 U1400 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1834), .ZN(n1837) );
NAND2_X1 U1401 ( .A1(n1840), .A2(n1841), .ZN(U325) );
NAND2_X1 U1402 ( .A1(n1833), .A2(DATA_IN_4_), .ZN(n1841) );
NAND2_X1 U1403 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1834), .ZN(n1840) );
NAND2_X1 U1404 ( .A1(n1842), .A2(n1843), .ZN(U324) );
NAND2_X1 U1405 ( .A1(n1833), .A2(DATA_IN_3_), .ZN(n1843) );
NAND2_X1 U1406 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1834), .ZN(n1842) );
NAND2_X1 U1407 ( .A1(n1844), .A2(n1845), .ZN(U323) );
NAND2_X1 U1408 ( .A1(n1833), .A2(DATA_IN_2_), .ZN(n1845) );
NAND2_X1 U1409 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1834), .ZN(n1844) );
NAND2_X1 U1410 ( .A1(n1846), .A2(n1847), .ZN(U322) );
NAND2_X1 U1411 ( .A1(DATA_IN_1_), .A2(n1848), .ZN(n1847) );
XOR2_X1 U1412 ( .A(KEYINPUT45), .B(n1833), .Z(n1848) );
NAND2_X1 U1413 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1834), .ZN(n1846) );
NAND2_X1 U1414 ( .A1(n1849), .A2(n1850), .ZN(U321) );
NAND2_X1 U1415 ( .A1(n1833), .A2(DATA_IN_0_), .ZN(n1850) );
AND2_X1 U1416 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1851), .ZN(n1833) );
XOR2_X1 U1417 ( .A(n1852), .B(KEYINPUT38), .Z(n1849) );
NAND2_X1 U1418 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1834), .ZN(n1852) );
NAND2_X1 U1419 ( .A1(n1717), .A2(n1851), .ZN(n1834) );
NAND2_X1 U1420 ( .A1(n1742), .A2(n1853), .ZN(n1851) );
NAND2_X1 U1421 ( .A1(n1742), .A2(n1854), .ZN(n1717) );
NAND2_X1 U1422 ( .A1(n1855), .A2(n1856), .ZN(U320) );
NAND2_X1 U1423 ( .A1(n1857), .A2(DATA_IN_7_), .ZN(n1856) );
NAND2_X1 U1424 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1858), .ZN(n1855) );
NAND2_X1 U1425 ( .A1(n1859), .A2(n1860), .ZN(U319) );
NAND2_X1 U1426 ( .A1(n1857), .A2(DATA_IN_6_), .ZN(n1860) );
NAND2_X1 U1427 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1858), .ZN(n1859) );
NAND2_X1 U1428 ( .A1(n1861), .A2(n1862), .ZN(U318) );
NAND2_X1 U1429 ( .A1(n1857), .A2(DATA_IN_5_), .ZN(n1862) );
NAND2_X1 U1430 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1858), .ZN(n1861) );
NAND2_X1 U1431 ( .A1(n1863), .A2(n1864), .ZN(U317) );
NAND2_X1 U1432 ( .A1(n1857), .A2(DATA_IN_4_), .ZN(n1864) );
XOR2_X1 U1433 ( .A(n1865), .B(KEYINPUT63), .Z(n1863) );
NAND2_X1 U1434 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1858), .ZN(n1865) );
NAND2_X1 U1435 ( .A1(n1866), .A2(n1867), .ZN(U316) );
NAND2_X1 U1436 ( .A1(n1857), .A2(DATA_IN_3_), .ZN(n1867) );
NAND2_X1 U1437 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1858), .ZN(n1866) );
NAND2_X1 U1438 ( .A1(n1868), .A2(n1869), .ZN(U315) );
NAND2_X1 U1439 ( .A1(n1857), .A2(DATA_IN_2_), .ZN(n1869) );
NAND2_X1 U1440 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1858), .ZN(n1868) );
NAND2_X1 U1441 ( .A1(n1870), .A2(n1871), .ZN(U314) );
NAND2_X1 U1442 ( .A1(n1857), .A2(DATA_IN_1_), .ZN(n1871) );
NAND2_X1 U1443 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1858), .ZN(n1870) );
NAND2_X1 U1444 ( .A1(n1872), .A2(n1873), .ZN(U313) );
NAND2_X1 U1445 ( .A1(n1857), .A2(DATA_IN_0_), .ZN(n1873) );
NAND2_X1 U1446 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1858), .ZN(n1872) );
NAND2_X1 U1447 ( .A1(n1874), .A2(n1875), .ZN(U312) );
NAND2_X1 U1448 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1857), .ZN(n1875) );
NAND2_X1 U1449 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1858), .ZN(n1874) );
NAND2_X1 U1450 ( .A1(n1876), .A2(n1877), .ZN(U311) );
NAND2_X1 U1451 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1857), .ZN(n1877) );
NAND2_X1 U1452 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1858), .ZN(n1876) );
NAND2_X1 U1453 ( .A1(n1878), .A2(n1879), .ZN(U310) );
NAND2_X1 U1454 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1857), .ZN(n1879) );
NAND2_X1 U1455 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1858), .ZN(n1878) );
NAND2_X1 U1456 ( .A1(n1880), .A2(n1881), .ZN(U309) );
NAND2_X1 U1457 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1857), .ZN(n1881) );
NAND2_X1 U1458 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1858), .ZN(n1880) );
NAND2_X1 U1459 ( .A1(n1882), .A2(n1883), .ZN(U308) );
NAND2_X1 U1460 ( .A1(n1884), .A2(REG1_REG_3__SCAN_IN), .ZN(n1883) );
XOR2_X1 U1461 ( .A(n1885), .B(KEYINPUT20), .Z(n1884) );
NAND2_X1 U1462 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1858), .ZN(n1882) );
NAND2_X1 U1463 ( .A1(n1886), .A2(n1887), .ZN(U307) );
NAND2_X1 U1464 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1857), .ZN(n1887) );
NAND2_X1 U1465 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1858), .ZN(n1886) );
NAND2_X1 U1466 ( .A1(n1888), .A2(n1889), .ZN(U306) );
NAND2_X1 U1467 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1857), .ZN(n1889) );
NAND2_X1 U1468 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1858), .ZN(n1888) );
NAND2_X1 U1469 ( .A1(n1890), .A2(n1891), .ZN(U305) );
NAND2_X1 U1470 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1858), .ZN(n1891) );
XOR2_X1 U1471 ( .A(n1892), .B(KEYINPUT7), .Z(n1890) );
NAND2_X1 U1472 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1893), .ZN(n1892) );
XOR2_X1 U1473 ( .A(KEYINPUT10), .B(n1857), .Z(n1893) );
NAND2_X1 U1474 ( .A1(n1894), .A2(n1895), .ZN(U304) );
NAND2_X1 U1475 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1857), .ZN(n1895) );
NAND2_X1 U1476 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1858), .ZN(n1894) );
NAND2_X1 U1477 ( .A1(n1896), .A2(n1897), .ZN(U303) );
NAND2_X1 U1478 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1898), .ZN(n1897) );
XOR2_X1 U1479 ( .A(KEYINPUT59), .B(n1858), .Z(n1898) );
NAND2_X1 U1480 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1857), .ZN(n1896) );
NAND2_X1 U1481 ( .A1(n1899), .A2(n1900), .ZN(U302) );
NAND2_X1 U1482 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1857), .ZN(n1900) );
NAND2_X1 U1483 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1858), .ZN(n1899) );
NAND2_X1 U1484 ( .A1(n1901), .A2(n1902), .ZN(U301) );
NAND2_X1 U1485 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1857), .ZN(n1902) );
NAND2_X1 U1486 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1858), .ZN(n1901) );
NAND2_X1 U1487 ( .A1(n1903), .A2(n1904), .ZN(U300) );
NAND2_X1 U1488 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1857), .ZN(n1904) );
NAND2_X1 U1489 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1858), .ZN(n1903) );
NAND2_X1 U1490 ( .A1(n1905), .A2(n1906), .ZN(U299) );
NAND2_X1 U1491 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1857), .ZN(n1906) );
NAND2_X1 U1492 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1858), .ZN(n1905) );
NAND2_X1 U1493 ( .A1(n1907), .A2(n1908), .ZN(U298) );
NAND2_X1 U1494 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1857), .ZN(n1908) );
NAND2_X1 U1495 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1858), .ZN(n1907) );
NAND2_X1 U1496 ( .A1(n1909), .A2(n1910), .ZN(U297) );
NAND2_X1 U1497 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1857), .ZN(n1910) );
NAND2_X1 U1498 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1858), .ZN(n1909) );
NAND2_X1 U1499 ( .A1(n1911), .A2(n1912), .ZN(U296) );
NAND2_X1 U1500 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1857), .ZN(n1912) );
NAND2_X1 U1501 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1858), .ZN(n1911) );
NAND2_X1 U1502 ( .A1(n1913), .A2(n1914), .ZN(U295) );
NAND2_X1 U1503 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1857), .ZN(n1914) );
NAND2_X1 U1504 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1858), .ZN(n1913) );
NAND2_X1 U1505 ( .A1(n1915), .A2(n1916), .ZN(U294) );
NAND2_X1 U1506 ( .A1(n1917), .A2(REG4_REG_5__SCAN_IN), .ZN(n1916) );
XOR2_X1 U1507 ( .A(U280), .B(KEYINPUT28), .Z(n1917) );
NAND2_X1 U1508 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1857), .ZN(n1915) );
NAND2_X1 U1509 ( .A1(n1918), .A2(n1919), .ZN(U293) );
NAND2_X1 U1510 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1857), .ZN(n1919) );
NAND2_X1 U1511 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1858), .ZN(n1918) );
NAND2_X1 U1512 ( .A1(n1920), .A2(n1921), .ZN(U292) );
NAND2_X1 U1513 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1857), .ZN(n1921) );
NAND2_X1 U1514 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1858), .ZN(n1920) );
NAND2_X1 U1515 ( .A1(n1922), .A2(n1923), .ZN(U291) );
NAND2_X1 U1516 ( .A1(n1924), .A2(n1858), .ZN(n1923) );
XOR2_X1 U1517 ( .A(REG4_REG_2__SCAN_IN), .B(KEYINPUT14), .Z(n1924) );
NAND2_X1 U1518 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1857), .ZN(n1922) );
NAND2_X1 U1519 ( .A1(n1925), .A2(n1926), .ZN(U290) );
NAND2_X1 U1520 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1857), .ZN(n1926) );
NAND2_X1 U1521 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1858), .ZN(n1925) );
NAND2_X1 U1522 ( .A1(n1927), .A2(n1928), .ZN(U289) );
NAND2_X1 U1523 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1857), .ZN(n1928) );
NAND2_X1 U1524 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1858), .ZN(n1927) );
NAND4_X1 U1525 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(U288));
NAND2_X1 U1526 ( .A1(n1933), .A2(n1934), .ZN(n1932) );
XOR2_X1 U1527 ( .A(REG4_REG_7__SCAN_IN), .B(KEYINPUT17), .Z(n1934) );
NAND2_X1 U1528 ( .A1(n1935), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1931) );
NAND2_X1 U1529 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1858), .ZN(n1930) );
NAND4_X1 U1530 ( .A1(n1936), .A2(n1937), .A3(n1938), .A4(n1939), .ZN(U287));
AND4_X1 U1531 ( .A1(n1929), .A2(n1940), .A3(n1941), .A4(n1942), .ZN(n1939));
OR2_X1 U1532 ( .A1(n1943), .A2(KEYINPUT1), .ZN(n1942) );
NAND4_X1 U1533 ( .A1(n1944), .A2(n1945), .A3(n1946), .A4(KEYINPUT1), .ZN(n1941) );
NAND2_X1 U1534 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1858), .ZN(n1940) );
AND2_X1 U1535 ( .A1(n1947), .A2(n1948), .ZN(n1929) );
OR3_X1 U1536 ( .A1(n1949), .A2(n1950), .A3(n1951), .ZN(n1948) );
NAND2_X1 U1537 ( .A1(n1952), .A2(n1953), .ZN(n1947) );
NAND2_X1 U1538 ( .A1(n1933), .A2(REG4_REG_6__SCAN_IN), .ZN(n1938) );
NAND3_X1 U1539 ( .A1(n1954), .A2(n1949), .A3(n1950), .ZN(n1937) );
NAND2_X1 U1540 ( .A1(n1935), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1936) );
NAND4_X1 U1541 ( .A1(n1955), .A2(n1956), .A3(n1957), .A4(n1958), .ZN(U286));
NOR3_X1 U1542 ( .A1(n1959), .A2(n1960), .A3(n1961), .ZN(n1958) );
NOR2_X1 U1543 ( .A1(n1962), .A2(n1963), .ZN(n1961) );
XOR2_X1 U1544 ( .A(n1964), .B(KEYINPUT57), .Z(n1962) );
NOR3_X1 U1545 ( .A1(n1951), .A2(n1950), .A3(n1965), .ZN(n1960) );
XOR2_X1 U1546 ( .A(n1966), .B(KEYINPUT50), .Z(n1965) );
NAND2_X1 U1547 ( .A1(n1967), .A2(n1968), .ZN(n1966) );
NOR2_X1 U1548 ( .A1(n1968), .A2(n1967), .ZN(n1950) );
AND2_X1 U1549 ( .A1(n1969), .A2(n1949), .ZN(n1967) );
NAND2_X1 U1550 ( .A1(n1970), .A2(n1971), .ZN(n1949) );
XOR2_X1 U1551 ( .A(n1972), .B(KEYINPUT51), .Z(n1969) );
NAND2_X1 U1552 ( .A1(n1973), .A2(n1974), .ZN(n1972) );
NOR2_X1 U1553 ( .A1(n1975), .A2(n1943), .ZN(n1959) );
INV_X1 U1554 ( .A(n1952), .ZN(n1943) );
NOR2_X1 U1555 ( .A1(n1976), .A2(n1946), .ZN(n1952) );
AND2_X1 U1556 ( .A1(n1977), .A2(n1978), .ZN(n1946) );
NAND2_X1 U1557 ( .A1(n1979), .A2(n1945), .ZN(n1978) );
NAND2_X1 U1558 ( .A1(n1973), .A2(n1980), .ZN(n1979) );
NOR3_X1 U1559 ( .A1(n1981), .A2(n1953), .A3(n1977), .ZN(n1975) );
INV_X1 U1560 ( .A(n1945), .ZN(n1953) );
NAND2_X1 U1561 ( .A1(n1982), .A2(n1971), .ZN(n1945) );
XOR2_X1 U1562 ( .A(n1980), .B(KEYINPUT24), .Z(n1982) );
NOR2_X1 U1563 ( .A1(n1983), .A2(n1971), .ZN(n1981) );
NAND2_X1 U1564 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1858), .ZN(n1957) );
NAND2_X1 U1565 ( .A1(n1984), .A2(n1973), .ZN(n1956) );
INV_X1 U1566 ( .A(n1971), .ZN(n1973) );
NAND2_X1 U1567 ( .A1(n1985), .A2(n1986), .ZN(n1971) );
NAND4_X1 U1568 ( .A1(n1987), .A2(n1988), .A3(n1989), .A4(n1990), .ZN(n1986));
NAND3_X1 U1569 ( .A1(n1991), .A2(KEYINPUT42), .A3(n1992), .ZN(n1990) );
INV_X1 U1570 ( .A(n1993), .ZN(n1992) );
NAND2_X1 U1571 ( .A1(n1993), .A2(n1994), .ZN(n1989) );
NAND2_X1 U1572 ( .A1(n1995), .A2(n1996), .ZN(n1994) );
NAND2_X1 U1573 ( .A1(n1997), .A2(n1998), .ZN(n1996) );
NAND2_X1 U1574 ( .A1(n1991), .A2(n1999), .ZN(n1995) );
NAND2_X1 U1575 ( .A1(KEYINPUT42), .A2(n1998), .ZN(n1999) );
INV_X1 U1576 ( .A(KEYINPUT46), .ZN(n1998) );
NAND2_X1 U1577 ( .A1(n2000), .A2(n2001), .ZN(n1988) );
NAND3_X1 U1578 ( .A1(n2001), .A2(n2002), .A3(n2003), .ZN(n1985) );
XOR2_X1 U1579 ( .A(n1993), .B(n2004), .Z(n2003) );
AND2_X1 U1580 ( .A1(KEYINPUT42), .A2(n1991), .ZN(n2004) );
INV_X1 U1581 ( .A(n1997), .ZN(n1991) );
NAND2_X1 U1582 ( .A1(n2005), .A2(n2006), .ZN(n1997) );
NAND2_X1 U1583 ( .A1(n2007), .A2(n2008), .ZN(n2006) );
NAND2_X1 U1584 ( .A1(KEYINPUT37), .A2(REG4_REG_6__SCAN_IN), .ZN(n2007) );
NAND2_X1 U1585 ( .A1(n2009), .A2(n1802), .ZN(n2005) );
INV_X1 U1586 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1802) );
NAND2_X1 U1587 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2010), .ZN(n2009) );
NAND2_X1 U1588 ( .A1(KEYINPUT37), .A2(RESTART), .ZN(n2010) );
NAND2_X1 U1589 ( .A1(n2011), .A2(n2012), .ZN(n1993) );
NAND2_X1 U1590 ( .A1(DATA_IN_6_), .A2(n2008), .ZN(n2012) );
NAND2_X1 U1591 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2011) );
NAND2_X1 U1592 ( .A1(n2013), .A2(n1987), .ZN(n2002) );
NAND2_X1 U1593 ( .A1(n2014), .A2(n2015), .ZN(n1987) );
NAND2_X1 U1594 ( .A1(n2016), .A2(n2017), .ZN(n2001) );
NAND2_X1 U1595 ( .A1(n1935), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1955) );
NAND4_X1 U1596 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(U285));
NOR3_X1 U1597 ( .A1(n2022), .A2(n2023), .A3(n2024), .ZN(n2021) );
NOR3_X1 U1598 ( .A1(n1976), .A2(n1977), .A3(n2025), .ZN(n2024) );
NOR3_X1 U1599 ( .A1(n2026), .A2(n1983), .A3(n2027), .ZN(n2025) );
AND2_X1 U1600 ( .A1(n2028), .A2(n2029), .ZN(n2027) );
INV_X1 U1601 ( .A(n1980), .ZN(n1983) );
AND2_X1 U1602 ( .A1(n2030), .A2(n2031), .ZN(n2026) );
AND3_X1 U1603 ( .A1(n2032), .A2(n2033), .A3(n2031), .ZN(n1977) );
NAND2_X1 U1604 ( .A1(n2034), .A2(n1980), .ZN(n2033) );
NAND2_X1 U1605 ( .A1(n2035), .A2(n2036), .ZN(n1980) );
XOR2_X1 U1606 ( .A(n2028), .B(KEYINPUT36), .Z(n2035) );
NAND2_X1 U1607 ( .A1(n2029), .A2(n2028), .ZN(n2034) );
XOR2_X1 U1608 ( .A(KEYINPUT34), .B(n2030), .Z(n2032) );
NOR3_X1 U1609 ( .A1(n1951), .A2(n2037), .A3(n2038), .ZN(n2023) );
NOR3_X1 U1610 ( .A1(n2029), .A2(n1970), .A3(n2039), .ZN(n2038) );
NOR2_X1 U1611 ( .A1(n2040), .A2(n2041), .ZN(n2039) );
INV_X1 U1612 ( .A(n1974), .ZN(n1970) );
INV_X1 U1613 ( .A(n1968), .ZN(n2037) );
NAND3_X1 U1614 ( .A1(n2042), .A2(n2043), .A3(n2044), .ZN(n1968) );
NAND2_X1 U1615 ( .A1(n2045), .A2(n1974), .ZN(n2042) );
NAND2_X1 U1616 ( .A1(n2046), .A2(n2036), .ZN(n1974) );
XOR2_X1 U1617 ( .A(n2047), .B(KEYINPUT35), .Z(n2046) );
NAND2_X1 U1618 ( .A1(n2029), .A2(n2047), .ZN(n2045) );
NOR2_X1 U1619 ( .A1(n2036), .A2(n2048), .ZN(n2022) );
INV_X1 U1620 ( .A(n2029), .ZN(n2036) );
NAND2_X1 U1621 ( .A1(n2049), .A2(n2050), .ZN(n2029) );
NAND2_X1 U1622 ( .A1(n2051), .A2(n2017), .ZN(n2050) );
XOR2_X1 U1623 ( .A(n2016), .B(n2013), .Z(n2051) );
NAND2_X1 U1624 ( .A1(n2052), .A2(n2015), .ZN(n2049) );
INV_X1 U1625 ( .A(n2017), .ZN(n2015) );
NAND3_X1 U1626 ( .A1(n2053), .A2(n2054), .A3(n2055), .ZN(n2017) );
NAND2_X1 U1627 ( .A1(n2056), .A2(n1800), .ZN(n2055) );
NAND2_X1 U1628 ( .A1(REG4_REG_5__SCAN_IN), .A2(n2008), .ZN(n2056) );
NAND3_X1 U1629 ( .A1(KEYINPUT6), .A2(n1964), .A3(n2008), .ZN(n2054) );
INV_X1 U1630 ( .A(REG4_REG_5__SCAN_IN), .ZN(n1964) );
OR2_X1 U1631 ( .A1(n2008), .A2(KEYINPUT6), .ZN(n2053) );
XOR2_X1 U1632 ( .A(n2057), .B(n2000), .Z(n2052) );
INV_X1 U1633 ( .A(n2013), .ZN(n2000) );
NAND2_X1 U1634 ( .A1(n2058), .A2(n2059), .ZN(n2013) );
NAND2_X1 U1635 ( .A1(RESTART), .A2(n1811), .ZN(n2059) );
NAND2_X1 U1636 ( .A1(n1801), .A2(n2008), .ZN(n2058) );
XNOR2_X1 U1637 ( .A(KEYINPUT26), .B(n2060), .ZN(n2057) );
NOR2_X1 U1638 ( .A1(KEYINPUT62), .A2(n2014), .ZN(n2060) );
INV_X1 U1639 ( .A(n2016), .ZN(n2014) );
NAND2_X1 U1640 ( .A1(n2061), .A2(n2062), .ZN(n2016) );
NAND2_X1 U1641 ( .A1(n2063), .A2(n2064), .ZN(n2062) );
OR2_X1 U1642 ( .A1(n2065), .A2(n2066), .ZN(n2061) );
NAND2_X1 U1643 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1858), .ZN(n2020) );
NAND2_X1 U1644 ( .A1(n1935), .A2(RLAST_REG_4__SCAN_IN), .ZN(n2019) );
NAND2_X1 U1645 ( .A1(n1933), .A2(REG4_REG_4__SCAN_IN), .ZN(n2018) );
NAND4_X1 U1646 ( .A1(n2067), .A2(n2068), .A3(n2069), .A4(n2070), .ZN(U284));
NOR3_X1 U1647 ( .A1(n2071), .A2(n2072), .A3(n2073), .ZN(n2070) );
AND2_X1 U1648 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1935), .ZN(n2073) );
NOR2_X1 U1649 ( .A1(n2074), .A2(n2048), .ZN(n2072) );
NOR2_X1 U1650 ( .A1(n2075), .A2(n1963), .ZN(n2071) );
NAND2_X1 U1651 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n2076), .ZN(n2069) );
XOR2_X1 U1652 ( .A(KEYINPUT53), .B(n1858), .Z(n2076) );
NAND2_X1 U1653 ( .A1(n2077), .A2(n1954), .ZN(n2068) );
XOR2_X1 U1654 ( .A(n2041), .B(n2040), .Z(n2077) );
INV_X1 U1655 ( .A(n2043), .ZN(n2040) );
NAND2_X1 U1656 ( .A1(n2047), .A2(n2078), .ZN(n2043) );
NAND2_X1 U1657 ( .A1(n2079), .A2(n2080), .ZN(n2078) );
OR2_X1 U1658 ( .A1(n2080), .A2(n2079), .ZN(n2047) );
NAND3_X1 U1659 ( .A1(n2081), .A2(n2082), .A3(n1944), .ZN(n2067) );
NAND2_X1 U1660 ( .A1(n2083), .A2(n2084), .ZN(n2082) );
NAND2_X1 U1661 ( .A1(n2031), .A2(n2030), .ZN(n2081) );
XNOR2_X1 U1662 ( .A(n2083), .B(KEYINPUT49), .ZN(n2031) );
AND2_X1 U1663 ( .A1(n2028), .A2(n2085), .ZN(n2083) );
NAND2_X1 U1664 ( .A1(n2079), .A2(n2086), .ZN(n2085) );
INV_X1 U1665 ( .A(n2074), .ZN(n2079) );
NAND2_X1 U1666 ( .A1(n2087), .A2(n2074), .ZN(n2028) );
XOR2_X1 U1667 ( .A(n2063), .B(n2088), .Z(n2074) );
NOR2_X1 U1668 ( .A1(n2089), .A2(n2090), .ZN(n2088) );
INV_X1 U1669 ( .A(n2064), .ZN(n2090) );
NAND2_X1 U1670 ( .A1(n2066), .A2(n2065), .ZN(n2064) );
NOR3_X1 U1671 ( .A1(n2065), .A2(KEYINPUT13), .A3(n2066), .ZN(n2089) );
AND2_X1 U1672 ( .A1(n2091), .A2(n2092), .ZN(n2066) );
NAND2_X1 U1673 ( .A1(n1785), .A2(n2008), .ZN(n2092) );
NAND2_X1 U1674 ( .A1(n2093), .A2(RESTART), .ZN(n2091) );
XOR2_X1 U1675 ( .A(n1818), .B(KEYINPUT22), .Z(n2093) );
NAND2_X1 U1676 ( .A1(n2094), .A2(n2095), .ZN(n2065) );
NAND2_X1 U1677 ( .A1(n2096), .A2(n2097), .ZN(n2095) );
NAND2_X1 U1678 ( .A1(n2098), .A2(n2099), .ZN(n2096) );
XOR2_X1 U1679 ( .A(n2100), .B(KEYINPUT4), .Z(n2094) );
NAND2_X1 U1680 ( .A1(n2101), .A2(n2102), .ZN(n2100) );
OR3_X1 U1681 ( .A1(n2103), .A2(n2098), .A3(KEYINPUT32), .ZN(n2102) );
NAND2_X1 U1682 ( .A1(KEYINPUT32), .A2(n2104), .ZN(n2101) );
NAND2_X1 U1683 ( .A1(n2105), .A2(n2106), .ZN(n2063) );
NAND2_X1 U1684 ( .A1(RESTART), .A2(n1781), .ZN(n2106) );
NAND2_X1 U1685 ( .A1(n2107), .A2(n2008), .ZN(n2105) );
NAND4_X1 U1686 ( .A1(n2108), .A2(n2109), .A3(n2110), .A4(n2111), .ZN(U283));
NOR3_X1 U1687 ( .A1(n2112), .A2(n2113), .A3(n2114), .ZN(n2111) );
NOR3_X1 U1688 ( .A1(n1976), .A2(n2030), .A3(n2115), .ZN(n2114) );
NOR4_X1 U1689 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2087), .ZN(n2115));
INV_X1 U1690 ( .A(n2086), .ZN(n2087) );
AND3_X1 U1691 ( .A1(KEYINPUT2), .A2(n2119), .A3(n2120), .ZN(n2117) );
INV_X1 U1692 ( .A(n2121), .ZN(n2120) );
NOR2_X1 U1693 ( .A1(KEYINPUT2), .A2(n2122), .ZN(n2116) );
INV_X1 U1694 ( .A(n2084), .ZN(n2030) );
NAND2_X1 U1695 ( .A1(n2123), .A2(n2124), .ZN(n2084) );
NAND2_X1 U1696 ( .A1(n2086), .A2(n2125), .ZN(n2124) );
NAND2_X1 U1697 ( .A1(n2126), .A2(n2127), .ZN(n2086) );
XOR2_X1 U1698 ( .A(KEYINPUT18), .B(n2128), .Z(n2127) );
INV_X1 U1699 ( .A(n1944), .ZN(n1976) );
NOR3_X1 U1700 ( .A1(n2129), .A2(n2130), .A3(n2044), .ZN(n2113) );
INV_X1 U1701 ( .A(n2041), .ZN(n2044) );
NAND2_X1 U1702 ( .A1(n2123), .A2(n2131), .ZN(n2041) );
NAND2_X1 U1703 ( .A1(n2080), .A2(n2125), .ZN(n2131) );
INV_X1 U1704 ( .A(n2118), .ZN(n2125) );
NAND2_X1 U1705 ( .A1(n2128), .A2(n2126), .ZN(n2080) );
NOR2_X1 U1706 ( .A1(n2118), .A2(n2123), .ZN(n2130) );
NOR2_X1 U1707 ( .A1(n2126), .A2(n2128), .ZN(n2118) );
XOR2_X1 U1708 ( .A(KEYINPUT21), .B(n1954), .Z(n2129) );
NOR2_X1 U1709 ( .A1(n2126), .A2(n2048), .ZN(n2112) );
AND2_X1 U1710 ( .A1(n2132), .A2(n2133), .ZN(n2126) );
NAND4_X1 U1711 ( .A1(n2134), .A2(n2097), .A3(n2135), .A4(n2136), .ZN(n2133));
OR3_X1 U1712 ( .A1(n2103), .A2(KEYINPUT40), .A3(n2098), .ZN(n2136) );
NAND2_X1 U1713 ( .A1(n2137), .A2(n2098), .ZN(n2135) );
NAND2_X1 U1714 ( .A1(n2138), .A2(n2139), .ZN(n2137) );
NAND2_X1 U1715 ( .A1(KEYINPUT40), .A2(n2099), .ZN(n2138) );
NAND2_X1 U1716 ( .A1(n2104), .A2(n2140), .ZN(n2134) );
INV_X1 U1717 ( .A(KEYINPUT54), .ZN(n2140) );
XOR2_X1 U1718 ( .A(n2141), .B(KEYINPUT33), .Z(n2132) );
NAND3_X1 U1719 ( .A1(n2142), .A2(n2143), .A3(n2144), .ZN(n2141) );
XOR2_X1 U1720 ( .A(n2097), .B(KEYINPUT44), .Z(n2144) );
NAND2_X1 U1721 ( .A1(n2145), .A2(n2146), .ZN(n2097) );
NAND2_X1 U1722 ( .A1(n2147), .A2(n2148), .ZN(n2146) );
NAND2_X1 U1723 ( .A1(n2149), .A2(n2150), .ZN(n2148) );
INV_X1 U1724 ( .A(n2151), .ZN(n2147) );
OR2_X1 U1725 ( .A1(n2150), .A2(n2149), .ZN(n2145) );
NAND2_X1 U1726 ( .A1(n2098), .A2(n2139), .ZN(n2143) );
NAND2_X1 U1727 ( .A1(n2103), .A2(KEYINPUT54), .ZN(n2139) );
INV_X1 U1728 ( .A(n2099), .ZN(n2103) );
NAND2_X1 U1729 ( .A1(KEYINPUT54), .A2(n2104), .ZN(n2142) );
NOR2_X1 U1730 ( .A1(n2099), .A2(n2098), .ZN(n2104) );
NAND2_X1 U1731 ( .A1(n2152), .A2(n2153), .ZN(n2098) );
NAND2_X1 U1732 ( .A1(RESTART), .A2(n1829), .ZN(n2153) );
NAND2_X1 U1733 ( .A1(n1798), .A2(n2008), .ZN(n2152) );
NAND2_X1 U1734 ( .A1(n2154), .A2(n2155), .ZN(n2099) );
NAND2_X1 U1735 ( .A1(RESTART), .A2(n1789), .ZN(n2155) );
NAND2_X1 U1736 ( .A1(n2075), .A2(n2008), .ZN(n2154) );
XOR2_X1 U1737 ( .A(KEYINPUT19), .B(n2156), .Z(n2110) );
NOR2_X1 U1738 ( .A1(n2157), .A2(n1963), .ZN(n2156) );
INV_X1 U1739 ( .A(n1933), .ZN(n1963) );
NAND2_X1 U1740 ( .A1(n1935), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2109) );
NAND2_X1 U1741 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1858), .ZN(n2108) );
NAND4_X1 U1742 ( .A1(n2158), .A2(n2159), .A3(n2160), .A4(n2161), .ZN(U282));
NAND2_X1 U1743 ( .A1(n1935), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2161) );
NOR2_X1 U1744 ( .A1(n2162), .A2(n2163), .ZN(n2160) );
NOR2_X1 U1745 ( .A1(n2164), .A2(n2165), .ZN(n2163) );
XOR2_X1 U1746 ( .A(KEYINPUT9), .B(n1984), .Z(n2165) );
INV_X1 U1747 ( .A(n2166), .ZN(n2164) );
NOR3_X1 U1748 ( .A1(n2167), .A2(n2123), .A3(n2168), .ZN(n2162) );
NOR2_X1 U1749 ( .A1(n2121), .A2(n2119), .ZN(n2168) );
INV_X1 U1750 ( .A(n2122), .ZN(n2123) );
NAND2_X1 U1751 ( .A1(n2121), .A2(n2119), .ZN(n2122) );
NAND2_X1 U1752 ( .A1(n2169), .A2(n2170), .ZN(n2119) );
NAND2_X1 U1753 ( .A1(n2166), .A2(n2171), .ZN(n2170) );
INV_X1 U1754 ( .A(n2128), .ZN(n2169) );
NOR2_X1 U1755 ( .A1(n2171), .A2(n2166), .ZN(n2128) );
NAND2_X1 U1756 ( .A1(n2172), .A2(n2173), .ZN(n2166) );
NAND2_X1 U1757 ( .A1(n2174), .A2(n2151), .ZN(n2173) );
XOR2_X1 U1758 ( .A(n2175), .B(KEYINPUT56), .Z(n2172) );
OR2_X1 U1759 ( .A1(n2151), .A2(n2174), .ZN(n2175) );
XOR2_X1 U1760 ( .A(n2150), .B(n2149), .Z(n2174) );
NAND2_X1 U1761 ( .A1(n2176), .A2(n2177), .ZN(n2149) );
NAND2_X1 U1762 ( .A1(RESTART), .A2(n2178), .ZN(n2177) );
NAND2_X1 U1763 ( .A1(n2157), .A2(n2008), .ZN(n2176) );
NAND3_X1 U1764 ( .A1(n2179), .A2(n2180), .A3(n2181), .ZN(n2150) );
NAND2_X1 U1765 ( .A1(n2182), .A2(n1825), .ZN(n2181) );
NAND2_X1 U1766 ( .A1(DATA_IN_2_), .A2(n2008), .ZN(n2182) );
NAND3_X1 U1767 ( .A1(KEYINPUT58), .A2(n1793), .A3(n2008), .ZN(n2180) );
OR2_X1 U1768 ( .A1(n2008), .A2(KEYINPUT58), .ZN(n2179) );
NAND2_X1 U1769 ( .A1(n2183), .A2(n2184), .ZN(n2151) );
NAND2_X1 U1770 ( .A1(n2185), .A2(n2186), .ZN(n2184) );
OR2_X1 U1771 ( .A1(n2187), .A2(n2188), .ZN(n2186) );
NAND2_X1 U1772 ( .A1(n2188), .A2(n2187), .ZN(n2183) );
NOR2_X1 U1773 ( .A1(n1954), .A2(n1944), .ZN(n2167) );
NAND2_X1 U1774 ( .A1(n1933), .A2(REG4_REG_1__SCAN_IN), .ZN(n2159) );
NAND2_X1 U1775 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1858), .ZN(n2158) );
NAND3_X1 U1776 ( .A1(n2189), .A2(n2190), .A3(n2191), .ZN(U281) );
NOR3_X1 U1777 ( .A1(n2192), .A2(n2193), .A3(n2194), .ZN(n2191) );
NOR2_X1 U1778 ( .A1(n2195), .A2(n2196), .ZN(n2194) );
INV_X1 U1779 ( .A(RLAST_REG_0__SCAN_IN), .ZN(n2196) );
XNOR2_X1 U1780 ( .A(n1935), .B(KEYINPUT47), .ZN(n2195) );
NOR2_X1 U1781 ( .A1(n2197), .A2(ENABLE), .ZN(n1935) );
NOR2_X1 U1782 ( .A1(n2198), .A2(n2199), .ZN(n2193) );
XOR2_X1 U1783 ( .A(KEYINPUT23), .B(n1933), .Z(n2199) );
NOR3_X1 U1784 ( .A1(n1853), .A2(n2197), .A3(n2200), .ZN(n1933) );
NOR2_X1 U1785 ( .A1(n2201), .A2(n2121), .ZN(n2192) );
NAND2_X1 U1786 ( .A1(n2171), .A2(n2202), .ZN(n2121) );
NAND3_X1 U1787 ( .A1(n2203), .A2(n2188), .A3(n2204), .ZN(n2202) );
OR2_X1 U1788 ( .A1(n2204), .A2(n2205), .ZN(n2171) );
AND2_X1 U1789 ( .A1(n2203), .A2(n2188), .ZN(n2205) );
NAND3_X1 U1790 ( .A1(n2206), .A2(n2207), .A3(n2208), .ZN(n2203) );
INV_X1 U1791 ( .A(n2209), .ZN(n2208) );
NAND2_X1 U1792 ( .A1(DATA_IN_0_), .A2(n2008), .ZN(n2207) );
NAND2_X1 U1793 ( .A1(RESTART), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2206) );
NOR2_X1 U1794 ( .A1(n1944), .A2(n2210), .ZN(n2201) );
XOR2_X1 U1795 ( .A(KEYINPUT48), .B(n1954), .Z(n2210) );
INV_X1 U1796 ( .A(n1951), .ZN(n1954) );
NAND4_X1 U1797 ( .A1(n2211), .A2(U280), .A3(n2212), .A4(n2213), .ZN(n1951));
NOR2_X1 U1798 ( .A1(n1854), .A2(n2008), .ZN(n2213) );
NOR4_X1 U1799 ( .A1(n1853), .A2(n2197), .A3(n2214), .A4(AVERAGE), .ZN(n1944));
NAND3_X1 U1800 ( .A1(U280), .A2(n2008), .A3(STATO_REG_1__SCAN_IN), .ZN(n2197) );
INV_X1 U1801 ( .A(ENABLE), .ZN(n1853) );
NAND2_X1 U1802 ( .A1(n1984), .A2(n2204), .ZN(n2190) );
XOR2_X1 U1803 ( .A(n2215), .B(n2187), .Z(n2204) );
NAND2_X1 U1804 ( .A1(n2216), .A2(n2217), .ZN(n2187) );
NAND2_X1 U1805 ( .A1(n2218), .A2(n2008), .ZN(n2217) );
NAND2_X1 U1806 ( .A1(DATA_IN_1_), .A2(n2219), .ZN(n2218) );
NAND2_X1 U1807 ( .A1(n2220), .A2(n2221), .ZN(n2216) );
NAND2_X1 U1808 ( .A1(DATA_IN_1_), .A2(n2222), .ZN(n2220) );
NAND2_X1 U1809 ( .A1(RESTART), .A2(n2219), .ZN(n2222) );
INV_X1 U1810 ( .A(KEYINPUT61), .ZN(n2219) );
NAND2_X1 U1811 ( .A1(KEYINPUT31), .A2(n2223), .ZN(n2215) );
XOR2_X1 U1812 ( .A(n2188), .B(n2185), .Z(n2223) );
AND2_X1 U1813 ( .A1(n2224), .A2(n2225), .ZN(n2185) );
NAND2_X1 U1814 ( .A1(REG4_REG_1__SCAN_IN), .A2(n2008), .ZN(n2225) );
NAND2_X1 U1815 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2224) );
NAND3_X1 U1816 ( .A1(n2226), .A2(n2227), .A3(n2209), .ZN(n2188) );
NAND3_X1 U1817 ( .A1(n2228), .A2(n2229), .A3(n2230), .ZN(n2209) );
NAND2_X1 U1818 ( .A1(RESTART), .A2(n2231), .ZN(n2230) );
OR2_X1 U1819 ( .A1(RMIN_REG_0__SCAN_IN), .A2(KEYINPUT0), .ZN(n2231) );
OR3_X1 U1820 ( .A1(n2198), .A2(RESTART), .A3(KEYINPUT0), .ZN(n2229) );
NAND2_X1 U1821 ( .A1(KEYINPUT0), .A2(n2198), .ZN(n2228) );
INV_X1 U1822 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2198) );
NAND2_X1 U1823 ( .A1(RESTART), .A2(n1827), .ZN(n2227) );
INV_X1 U1824 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1827) );
NAND2_X1 U1825 ( .A1(n1744), .A2(n2008), .ZN(n2226) );
INV_X1 U1826 ( .A(n2048), .ZN(n1984) );
NAND4_X1 U1827 ( .A1(STATO_REG_1__SCAN_IN), .A2(U280), .A3(n2232), .A4(n2233), .ZN(n2048) );
NAND2_X1 U1828 ( .A1(n2234), .A2(n2008), .ZN(n2233) );
INV_X1 U1829 ( .A(RESTART), .ZN(n2008) );
NAND3_X1 U1830 ( .A1(n2214), .A2(n2200), .A3(ENABLE), .ZN(n2234) );
INV_X1 U1831 ( .A(AVERAGE), .ZN(n2200) );
NAND2_X1 U1832 ( .A1(n2235), .A2(n2236), .ZN(n2214) );
NAND2_X1 U1833 ( .A1(n2237), .A2(n2238), .ZN(n2236) );
INV_X1 U1834 ( .A(REG4_REG_7__SCAN_IN), .ZN(n2238) );
OR2_X1 U1835 ( .A1(n2239), .A2(n1773), .ZN(n2237) );
NAND2_X1 U1836 ( .A1(n2239), .A2(n1773), .ZN(n2235) );
INV_X1 U1837 ( .A(DATA_IN_7_), .ZN(n1773) );
NAND2_X1 U1838 ( .A1(n2240), .A2(n2241), .ZN(n2239) );
NAND2_X1 U1839 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2242), .ZN(n2241) );
NAND2_X1 U1840 ( .A1(n1777), .A2(n2243), .ZN(n2242) );
OR2_X1 U1841 ( .A1(n2243), .A2(n1777), .ZN(n2240) );
INV_X1 U1842 ( .A(DATA_IN_6_), .ZN(n1777) );
NAND2_X1 U1843 ( .A1(n2244), .A2(n2245), .ZN(n2243) );
NAND2_X1 U1844 ( .A1(n2246), .A2(n1801), .ZN(n2245) );
INV_X1 U1845 ( .A(DATA_IN_5_), .ZN(n1801) );
NAND2_X1 U1846 ( .A1(n2247), .A2(n2248), .ZN(n2246) );
XOR2_X1 U1847 ( .A(REG4_REG_5__SCAN_IN), .B(KEYINPUT25), .Z(n2247) );
OR2_X1 U1848 ( .A1(n2248), .A2(REG4_REG_5__SCAN_IN), .ZN(n2244) );
NAND2_X1 U1849 ( .A1(n2249), .A2(n2250), .ZN(n2248) );
NAND3_X1 U1850 ( .A1(n2251), .A2(n2252), .A3(n2253), .ZN(n2250) );
NAND2_X1 U1851 ( .A1(n1785), .A2(n2107), .ZN(n2253) );
INV_X1 U1852 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2107) );
INV_X1 U1853 ( .A(DATA_IN_4_), .ZN(n1785) );
NAND3_X1 U1854 ( .A1(n2254), .A2(n2255), .A3(n2256), .ZN(n2252) );
NAND2_X1 U1855 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2256) );
NAND3_X1 U1856 ( .A1(n2257), .A2(n2258), .A3(n2259), .ZN(n2255) );
NAND2_X1 U1857 ( .A1(n1793), .A2(n2157), .ZN(n2259) );
INV_X1 U1858 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2157) );
INV_X1 U1859 ( .A(DATA_IN_2_), .ZN(n1793) );
NAND2_X1 U1860 ( .A1(n2260), .A2(n1796), .ZN(n2258) );
INV_X1 U1861 ( .A(DATA_IN_1_), .ZN(n1796) );
NAND2_X1 U1862 ( .A1(n2261), .A2(n2262), .ZN(n2260) );
XNOR2_X1 U1863 ( .A(REG4_REG_1__SCAN_IN), .B(KEYINPUT55), .ZN(n2261) );
OR2_X1 U1864 ( .A1(n2262), .A2(REG4_REG_1__SCAN_IN), .ZN(n2257) );
AND2_X1 U1865 ( .A1(n2263), .A2(REG4_REG_0__SCAN_IN), .ZN(n2262) );
XOR2_X1 U1866 ( .A(n1744), .B(KEYINPUT12), .Z(n2263) );
INV_X1 U1867 ( .A(DATA_IN_0_), .ZN(n1744) );
NAND2_X1 U1868 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2254) );
NAND2_X1 U1869 ( .A1(n1798), .A2(n2075), .ZN(n2251) );
INV_X1 U1870 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2075) );
INV_X1 U1871 ( .A(DATA_IN_3_), .ZN(n1798) );
NAND2_X1 U1872 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2249) );
NAND3_X1 U1873 ( .A1(n2212), .A2(n2211), .A3(RESTART), .ZN(n2232) );
NAND3_X1 U1874 ( .A1(n2264), .A2(n2265), .A3(n2266), .ZN(n2211) );
OR2_X1 U1875 ( .A1(RMAX_REG_6__SCAN_IN), .A2(RMIN_REG_6__SCAN_IN), .ZN(n2266) );
NAND2_X1 U1876 ( .A1(n2267), .A2(n2268), .ZN(n2265) );
NAND2_X1 U1877 ( .A1(RMIN_REG_6__SCAN_IN), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2268) );
NAND2_X1 U1878 ( .A1(n2269), .A2(n2270), .ZN(n2267) );
NAND2_X1 U1879 ( .A1(n1811), .A2(n1800), .ZN(n2270) );
INV_X1 U1880 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1800) );
INV_X1 U1881 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1811) );
NAND3_X1 U1882 ( .A1(n2271), .A2(n2272), .A3(n2273), .ZN(n2269) );
NAND2_X1 U1883 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2273) );
NAND3_X1 U1884 ( .A1(n2274), .A2(n2275), .A3(n2276), .ZN(n2272) );
NAND2_X1 U1885 ( .A1(n1818), .A2(n1781), .ZN(n2276) );
INV_X1 U1886 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1781) );
INV_X1 U1887 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1818) );
NAND3_X1 U1888 ( .A1(n2277), .A2(n2278), .A3(n2279), .ZN(n2275) );
NAND2_X1 U1889 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2279) );
NAND3_X1 U1890 ( .A1(n2280), .A2(n2281), .A3(n2282), .ZN(n2278) );
XOR2_X1 U1891 ( .A(n2283), .B(KEYINPUT5), .Z(n2282) );
NAND2_X1 U1892 ( .A1(n2178), .A2(n1825), .ZN(n2283) );
INV_X1 U1893 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1825) );
INV_X1 U1894 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n2178) );
NAND2_X1 U1895 ( .A1(n2284), .A2(n1795), .ZN(n2281) );
INV_X1 U1896 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1795) );
OR2_X1 U1897 ( .A1(n2285), .A2(n2221), .ZN(n2284) );
NAND2_X1 U1898 ( .A1(n2285), .A2(n2221), .ZN(n2280) );
INV_X1 U1899 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n2221) );
NAND2_X1 U1900 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2285) );
NAND2_X1 U1901 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n2286), .ZN(n2277) );
XOR2_X1 U1902 ( .A(RMIN_REG_3__SCAN_IN), .B(KEYINPUT29), .Z(n2286) );
NAND2_X1 U1903 ( .A1(n1829), .A2(n1789), .ZN(n2274) );
INV_X1 U1904 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1789) );
INV_X1 U1905 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1829) );
NAND2_X1 U1906 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2271) );
NAND2_X1 U1907 ( .A1(n2287), .A2(RMIN_REG_7__SCAN_IN), .ZN(n2264) );
XOR2_X1 U1908 ( .A(n1807), .B(KEYINPUT52), .Z(n2287) );
NAND2_X1 U1909 ( .A1(n1803), .A2(n1807), .ZN(n2212) );
INV_X1 U1910 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1807) );
INV_X1 U1911 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1803) );
NAND2_X1 U1912 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1858), .ZN(n2189) );
NAND2_X1 U1913 ( .A1(n1885), .A2(n2288), .ZN(U280) );
NAND2_X1 U1914 ( .A1(STATO_REG_0__SCAN_IN), .A2(n1854), .ZN(n2288) );
INV_X1 U1915 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1854) );
NAND2_X1 U1916 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1742), .ZN(n1885) );
INV_X1 U1917 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1742) );
endmodule


