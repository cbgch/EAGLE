//Key = 1000101000111011100101001101011001111111010111001110001010101011


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
n2250;

OR2_X1 U1264 ( .A1(n1749), .A2(STATO_REG_0__SCAN_IN), .ZN(n1690) );
INV_X2 U1265 ( .A(n1690), .ZN(n1691) );
INV_X2 U1266 ( .A(U280), .ZN(n1844) );
XNOR2_X1 U1267 ( .A(KEYINPUT7), .B(n1692), .ZN(U375) );
NAND2_X1 U1268 ( .A1(n1693), .A2(n1694), .ZN(U344) );
NAND2_X1 U1269 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1695), .ZN(n1694) );
NAND2_X1 U1270 ( .A1(DATA_IN_7_), .A2(n1696), .ZN(n1693) );
NAND2_X1 U1271 ( .A1(n1697), .A2(n1698), .ZN(U343) );
NAND2_X1 U1272 ( .A1(DATA_IN_6_), .A2(n1696), .ZN(n1698) );
XOR2_X1 U1273 ( .A(n1699), .B(KEYINPUT42), .Z(n1697) );
NAND2_X1 U1274 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1695), .ZN(n1699) );
NAND2_X1 U1275 ( .A1(n1700), .A2(n1701), .ZN(U342) );
NAND2_X1 U1276 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1695), .ZN(n1701) );
NAND2_X1 U1277 ( .A1(DATA_IN_5_), .A2(n1696), .ZN(n1700) );
NAND2_X1 U1278 ( .A1(n1702), .A2(n1703), .ZN(U341) );
NAND2_X1 U1279 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1695), .ZN(n1703) );
NAND2_X1 U1280 ( .A1(DATA_IN_4_), .A2(n1696), .ZN(n1702) );
NAND2_X1 U1281 ( .A1(n1704), .A2(n1705), .ZN(U340) );
NAND2_X1 U1282 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1695), .ZN(n1705) );
NAND2_X1 U1283 ( .A1(DATA_IN_3_), .A2(n1696), .ZN(n1704) );
NAND2_X1 U1284 ( .A1(n1706), .A2(n1707), .ZN(U339) );
NAND2_X1 U1285 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1695), .ZN(n1707) );
NAND2_X1 U1286 ( .A1(DATA_IN_2_), .A2(n1696), .ZN(n1706) );
NAND2_X1 U1287 ( .A1(n1708), .A2(n1709), .ZN(U338) );
NAND2_X1 U1288 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1695), .ZN(n1709) );
XOR2_X1 U1289 ( .A(KEYINPUT38), .B(n1710), .Z(n1708) );
NOR2_X1 U1290 ( .A1(n1711), .A2(n1712), .ZN(n1710) );
XOR2_X1 U1291 ( .A(n1696), .B(KEYINPUT50), .Z(n1711) );
NAND2_X1 U1292 ( .A1(n1713), .A2(n1714), .ZN(U337) );
NAND2_X1 U1293 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1695), .ZN(n1714) );
NAND2_X1 U1294 ( .A1(n1692), .A2(n1715), .ZN(n1695) );
NAND2_X1 U1295 ( .A1(n1716), .A2(n1717), .ZN(n1715) );
XNOR2_X1 U1296 ( .A(n1718), .B(KEYINPUT19), .ZN(n1716) );
NAND2_X1 U1297 ( .A1(DATA_IN_0_), .A2(n1696), .ZN(n1713) );
NAND2_X1 U1298 ( .A1(n1717), .A2(n1719), .ZN(n1696) );
NAND2_X1 U1299 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1720), .ZN(n1719) );
NAND2_X1 U1300 ( .A1(n1721), .A2(n1722), .ZN(U336) );
NAND2_X1 U1301 ( .A1(DATA_IN_7_), .A2(n1723), .ZN(n1722) );
NAND2_X1 U1302 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1724), .ZN(n1721) );
NAND2_X1 U1303 ( .A1(n1725), .A2(n1726), .ZN(U335) );
NAND2_X1 U1304 ( .A1(DATA_IN_6_), .A2(n1723), .ZN(n1726) );
NAND2_X1 U1305 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1724), .ZN(n1725) );
NAND2_X1 U1306 ( .A1(n1727), .A2(n1728), .ZN(U334) );
NAND2_X1 U1307 ( .A1(DATA_IN_5_), .A2(n1723), .ZN(n1728) );
NAND2_X1 U1308 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1724), .ZN(n1727) );
NAND2_X1 U1309 ( .A1(n1729), .A2(n1730), .ZN(U333) );
NAND2_X1 U1310 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1724), .ZN(n1730) );
XOR2_X1 U1311 ( .A(KEYINPUT11), .B(n1731), .Z(n1729) );
NOR2_X1 U1312 ( .A1(n1732), .A2(n1733), .ZN(n1731) );
NAND2_X1 U1313 ( .A1(n1734), .A2(n1735), .ZN(U332) );
NAND2_X1 U1314 ( .A1(n1736), .A2(n1724), .ZN(n1735) );
XNOR2_X1 U1315 ( .A(RMIN_REG_3__SCAN_IN), .B(KEYINPUT41), .ZN(n1736) );
NAND2_X1 U1316 ( .A1(DATA_IN_3_), .A2(n1723), .ZN(n1734) );
NAND2_X1 U1317 ( .A1(n1737), .A2(n1738), .ZN(U331) );
NAND2_X1 U1318 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1724), .ZN(n1738) );
XOR2_X1 U1319 ( .A(KEYINPUT16), .B(n1739), .Z(n1737) );
NOR2_X1 U1320 ( .A1(n1732), .A2(n1740), .ZN(n1739) );
NAND2_X1 U1321 ( .A1(n1741), .A2(n1742), .ZN(U330) );
NAND2_X1 U1322 ( .A1(n1743), .A2(DATA_IN_1_), .ZN(n1742) );
XNOR2_X1 U1323 ( .A(n1732), .B(KEYINPUT23), .ZN(n1743) );
INV_X1 U1324 ( .A(n1723), .ZN(n1732) );
NAND2_X1 U1325 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1724), .ZN(n1741) );
NAND2_X1 U1326 ( .A1(n1744), .A2(n1745), .ZN(U329) );
NAND2_X1 U1327 ( .A1(DATA_IN_0_), .A2(n1723), .ZN(n1745) );
NAND2_X1 U1328 ( .A1(n1746), .A2(n1747), .ZN(n1723) );
OR2_X1 U1329 ( .A1(n1748), .A2(n1749), .ZN(n1747) );
XNOR2_X1 U1330 ( .A(n1717), .B(KEYINPUT30), .ZN(n1746) );
NAND2_X1 U1331 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1724), .ZN(n1744) );
NAND2_X1 U1332 ( .A1(n1692), .A2(n1750), .ZN(n1724) );
NAND2_X1 U1333 ( .A1(n1748), .A2(n1717), .ZN(n1750) );
NAND2_X1 U1334 ( .A1(n1718), .A2(n1751), .ZN(n1748) );
NAND2_X1 U1335 ( .A1(n1752), .A2(n1753), .ZN(n1751) );
NAND3_X1 U1336 ( .A1(n1754), .A2(n1755), .A3(n1756), .ZN(n1753) );
NAND2_X1 U1337 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1757), .ZN(n1756) );
NAND3_X1 U1338 ( .A1(n1758), .A2(n1759), .A3(n1760), .ZN(n1755) );
NAND2_X1 U1339 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1761), .ZN(n1760) );
NAND3_X1 U1340 ( .A1(n1762), .A2(n1763), .A3(n1764), .ZN(n1759) );
NAND2_X1 U1341 ( .A1(DATA_IN_4_), .A2(n1765), .ZN(n1764) );
NAND3_X1 U1342 ( .A1(n1766), .A2(n1767), .A3(n1768), .ZN(n1763) );
NAND2_X1 U1343 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1733), .ZN(n1768) );
NAND3_X1 U1344 ( .A1(n1769), .A2(n1770), .A3(n1771), .ZN(n1767) );
NAND2_X1 U1345 ( .A1(DATA_IN_3_), .A2(n1772), .ZN(n1771) );
NAND3_X1 U1346 ( .A1(n1773), .A2(n1774), .A3(n1775), .ZN(n1770) );
NAND2_X1 U1347 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1740), .ZN(n1775) );
NAND3_X1 U1348 ( .A1(n1776), .A2(n1777), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1774) );
NAND2_X1 U1349 ( .A1(DATA_IN_1_), .A2(n1778), .ZN(n1776) );
NAND2_X1 U1350 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1712), .ZN(n1773) );
NAND2_X1 U1351 ( .A1(DATA_IN_2_), .A2(n1779), .ZN(n1769) );
NAND2_X1 U1352 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1780), .ZN(n1766) );
NAND2_X1 U1353 ( .A1(n1781), .A2(DATA_IN_5_), .ZN(n1762) );
XNOR2_X1 U1354 ( .A(RMIN_REG_5__SCAN_IN), .B(KEYINPUT13), .ZN(n1781) );
NAND2_X1 U1355 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1782), .ZN(n1758) );
NAND2_X1 U1356 ( .A1(DATA_IN_6_), .A2(n1783), .ZN(n1754) );
OR2_X1 U1357 ( .A1(n1757), .A2(RMIN_REG_7__SCAN_IN), .ZN(n1752) );
INV_X1 U1358 ( .A(n1720), .ZN(n1718) );
NAND2_X1 U1359 ( .A1(n1784), .A2(n1785), .ZN(n1720) );
NAND2_X1 U1360 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1757), .ZN(n1785) );
INV_X1 U1361 ( .A(DATA_IN_7_), .ZN(n1757) );
NAND3_X1 U1362 ( .A1(n1786), .A2(n1787), .A3(n1788), .ZN(n1784) );
NAND2_X1 U1363 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1789), .ZN(n1788) );
XNOR2_X1 U1364 ( .A(KEYINPUT0), .B(n1761), .ZN(n1789) );
NAND3_X1 U1365 ( .A1(n1790), .A2(n1791), .A3(n1792), .ZN(n1787) );
XOR2_X1 U1366 ( .A(n1793), .B(KEYINPUT53), .Z(n1792) );
NAND2_X1 U1367 ( .A1(DATA_IN_5_), .A2(n1794), .ZN(n1793) );
NAND3_X1 U1368 ( .A1(n1795), .A2(n1796), .A3(n1797), .ZN(n1791) );
NAND2_X1 U1369 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1782), .ZN(n1797) );
NAND3_X1 U1370 ( .A1(n1798), .A2(n1799), .A3(n1800), .ZN(n1796) );
NAND2_X1 U1371 ( .A1(DATA_IN_4_), .A2(n1801), .ZN(n1800) );
NAND3_X1 U1372 ( .A1(n1802), .A2(n1803), .A3(n1804), .ZN(n1799) );
NAND2_X1 U1373 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1780), .ZN(n1804) );
NAND3_X1 U1374 ( .A1(n1805), .A2(n1806), .A3(n1807), .ZN(n1803) );
NAND2_X1 U1375 ( .A1(DATA_IN_2_), .A2(n1808), .ZN(n1807) );
NAND3_X1 U1376 ( .A1(n1809), .A2(n1810), .A3(DATA_IN_0_), .ZN(n1806) );
INV_X1 U1377 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1810) );
NAND2_X1 U1378 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1712), .ZN(n1809) );
NAND2_X1 U1379 ( .A1(DATA_IN_1_), .A2(n1811), .ZN(n1805) );
NAND2_X1 U1380 ( .A1(n1812), .A2(n1740), .ZN(n1802) );
XNOR2_X1 U1381 ( .A(n1808), .B(KEYINPUT55), .ZN(n1812) );
NAND2_X1 U1382 ( .A1(DATA_IN_3_), .A2(n1813), .ZN(n1798) );
NAND2_X1 U1383 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1733), .ZN(n1795) );
NAND2_X1 U1384 ( .A1(DATA_IN_6_), .A2(n1814), .ZN(n1790) );
NAND2_X1 U1385 ( .A1(n1815), .A2(DATA_IN_7_), .ZN(n1786) );
XNOR2_X1 U1386 ( .A(RMAX_REG_7__SCAN_IN), .B(KEYINPUT32), .ZN(n1815) );
NAND2_X1 U1387 ( .A1(n1816), .A2(n1817), .ZN(U328) );
NAND2_X1 U1388 ( .A1(n1818), .A2(DATA_IN_7_), .ZN(n1817) );
NAND2_X1 U1389 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1819), .ZN(n1816) );
NAND2_X1 U1390 ( .A1(n1820), .A2(n1821), .ZN(U327) );
NAND2_X1 U1391 ( .A1(n1818), .A2(DATA_IN_6_), .ZN(n1821) );
NAND2_X1 U1392 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1819), .ZN(n1820) );
NAND2_X1 U1393 ( .A1(n1822), .A2(n1823), .ZN(U326) );
NAND2_X1 U1394 ( .A1(n1818), .A2(DATA_IN_5_), .ZN(n1823) );
NAND2_X1 U1395 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1819), .ZN(n1822) );
NAND2_X1 U1396 ( .A1(n1824), .A2(n1825), .ZN(U325) );
NAND2_X1 U1397 ( .A1(n1826), .A2(DATA_IN_4_), .ZN(n1825) );
XNOR2_X1 U1398 ( .A(n1818), .B(KEYINPUT6), .ZN(n1826) );
XOR2_X1 U1399 ( .A(KEYINPUT62), .B(n1827), .Z(n1824) );
NOR2_X1 U1400 ( .A1(n1828), .A2(n1829), .ZN(n1827) );
XNOR2_X1 U1401 ( .A(RLAST_REG_4__SCAN_IN), .B(KEYINPUT22), .ZN(n1829) );
INV_X1 U1402 ( .A(n1819), .ZN(n1828) );
NAND2_X1 U1403 ( .A1(n1830), .A2(n1831), .ZN(U324) );
NAND2_X1 U1404 ( .A1(n1818), .A2(DATA_IN_3_), .ZN(n1831) );
NAND2_X1 U1405 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1819), .ZN(n1830) );
NAND2_X1 U1406 ( .A1(n1832), .A2(n1833), .ZN(U323) );
NAND2_X1 U1407 ( .A1(n1818), .A2(DATA_IN_2_), .ZN(n1833) );
NAND2_X1 U1408 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1819), .ZN(n1832) );
NAND2_X1 U1409 ( .A1(n1834), .A2(n1835), .ZN(U322) );
NAND2_X1 U1410 ( .A1(n1818), .A2(DATA_IN_1_), .ZN(n1835) );
NAND2_X1 U1411 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1819), .ZN(n1834) );
NAND2_X1 U1412 ( .A1(n1836), .A2(n1837), .ZN(U321) );
NAND2_X1 U1413 ( .A1(n1818), .A2(DATA_IN_0_), .ZN(n1837) );
AND2_X1 U1414 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1838), .ZN(n1818) );
NAND2_X1 U1415 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1819), .ZN(n1836) );
NAND2_X1 U1416 ( .A1(n1692), .A2(n1838), .ZN(n1819) );
NAND2_X1 U1417 ( .A1(n1717), .A2(n1839), .ZN(n1838) );
NAND2_X1 U1418 ( .A1(n1840), .A2(n1749), .ZN(n1692) );
XNOR2_X1 U1419 ( .A(n1717), .B(KEYINPUT35), .ZN(n1840) );
INV_X1 U1420 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1717) );
NAND2_X1 U1421 ( .A1(n1841), .A2(n1842), .ZN(U320) );
NAND2_X1 U1422 ( .A1(DATA_IN_7_), .A2(n1843), .ZN(n1842) );
XNOR2_X1 U1423 ( .A(KEYINPUT59), .B(n1690), .ZN(n1843) );
NAND2_X1 U1424 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1844), .ZN(n1841) );
NAND2_X1 U1425 ( .A1(n1845), .A2(n1846), .ZN(U319) );
NAND2_X1 U1426 ( .A1(n1691), .A2(DATA_IN_6_), .ZN(n1846) );
NAND2_X1 U1427 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1844), .ZN(n1845) );
NAND2_X1 U1428 ( .A1(n1847), .A2(n1848), .ZN(U318) );
NAND2_X1 U1429 ( .A1(n1691), .A2(DATA_IN_5_), .ZN(n1848) );
NAND2_X1 U1430 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1844), .ZN(n1847) );
NAND2_X1 U1431 ( .A1(n1849), .A2(n1850), .ZN(U317) );
NAND2_X1 U1432 ( .A1(n1851), .A2(DATA_IN_4_), .ZN(n1850) );
XNOR2_X1 U1433 ( .A(n1691), .B(KEYINPUT34), .ZN(n1851) );
NAND2_X1 U1434 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1844), .ZN(n1849) );
NAND2_X1 U1435 ( .A1(n1852), .A2(n1853), .ZN(U316) );
NAND2_X1 U1436 ( .A1(n1691), .A2(DATA_IN_3_), .ZN(n1853) );
NAND2_X1 U1437 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1844), .ZN(n1852) );
NAND2_X1 U1438 ( .A1(n1854), .A2(n1855), .ZN(U315) );
NAND2_X1 U1439 ( .A1(n1691), .A2(DATA_IN_2_), .ZN(n1855) );
NAND2_X1 U1440 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1844), .ZN(n1854) );
NAND2_X1 U1441 ( .A1(n1856), .A2(n1857), .ZN(U314) );
NAND2_X1 U1442 ( .A1(n1691), .A2(DATA_IN_1_), .ZN(n1857) );
XOR2_X1 U1443 ( .A(n1858), .B(KEYINPUT18), .Z(n1856) );
NAND2_X1 U1444 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1844), .ZN(n1858) );
NAND2_X1 U1445 ( .A1(n1859), .A2(n1860), .ZN(U313) );
NAND2_X1 U1446 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1861), .ZN(n1860) );
XNOR2_X1 U1447 ( .A(KEYINPUT47), .B(U280), .ZN(n1861) );
NAND2_X1 U1448 ( .A1(n1691), .A2(DATA_IN_0_), .ZN(n1859) );
NAND2_X1 U1449 ( .A1(n1862), .A2(n1863), .ZN(U312) );
NAND2_X1 U1450 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1691), .ZN(n1863) );
NAND2_X1 U1451 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1844), .ZN(n1862) );
NAND2_X1 U1452 ( .A1(n1864), .A2(n1865), .ZN(U311) );
NAND2_X1 U1453 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1691), .ZN(n1865) );
NAND2_X1 U1454 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1844), .ZN(n1864) );
NAND2_X1 U1455 ( .A1(n1866), .A2(n1867), .ZN(U310) );
NAND2_X1 U1456 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1691), .ZN(n1867) );
NAND2_X1 U1457 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1844), .ZN(n1866) );
NAND2_X1 U1458 ( .A1(n1868), .A2(n1869), .ZN(U309) );
NAND2_X1 U1459 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1691), .ZN(n1869) );
NAND2_X1 U1460 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1844), .ZN(n1868) );
NAND2_X1 U1461 ( .A1(n1870), .A2(n1871), .ZN(U308) );
NAND2_X1 U1462 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1844), .ZN(n1871) );
XOR2_X1 U1463 ( .A(n1872), .B(KEYINPUT26), .Z(n1870) );
NAND2_X1 U1464 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1691), .ZN(n1872) );
NAND2_X1 U1465 ( .A1(n1873), .A2(n1874), .ZN(U307) );
NAND2_X1 U1466 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1691), .ZN(n1874) );
NAND2_X1 U1467 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1844), .ZN(n1873) );
NAND2_X1 U1468 ( .A1(n1875), .A2(n1876), .ZN(U306) );
NAND2_X1 U1469 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1691), .ZN(n1876) );
NAND2_X1 U1470 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1844), .ZN(n1875) );
NAND2_X1 U1471 ( .A1(n1877), .A2(n1878), .ZN(U305) );
NAND2_X1 U1472 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1691), .ZN(n1878) );
NAND2_X1 U1473 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1844), .ZN(n1877) );
NAND2_X1 U1474 ( .A1(n1879), .A2(n1880), .ZN(U304) );
NAND2_X1 U1475 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1691), .ZN(n1880) );
NAND2_X1 U1476 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1844), .ZN(n1879) );
NAND2_X1 U1477 ( .A1(n1881), .A2(n1882), .ZN(U303) );
NAND2_X1 U1478 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1691), .ZN(n1882) );
NAND2_X1 U1479 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1844), .ZN(n1881) );
NAND2_X1 U1480 ( .A1(n1883), .A2(n1884), .ZN(U302) );
NAND2_X1 U1481 ( .A1(n1885), .A2(n1844), .ZN(n1884) );
XNOR2_X1 U1482 ( .A(REG3_REG_5__SCAN_IN), .B(KEYINPUT39), .ZN(n1885) );
NAND2_X1 U1483 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1691), .ZN(n1883) );
NAND2_X1 U1484 ( .A1(n1886), .A2(n1887), .ZN(U301) );
NAND2_X1 U1485 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1691), .ZN(n1887) );
NAND2_X1 U1486 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1844), .ZN(n1886) );
NAND2_X1 U1487 ( .A1(n1888), .A2(n1889), .ZN(U300) );
NAND2_X1 U1488 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1691), .ZN(n1889) );
NAND2_X1 U1489 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1844), .ZN(n1888) );
NAND2_X1 U1490 ( .A1(n1890), .A2(n1891), .ZN(U299) );
NAND2_X1 U1491 ( .A1(n1892), .A2(n1691), .ZN(n1891) );
XNOR2_X1 U1492 ( .A(REG2_REG_2__SCAN_IN), .B(KEYINPUT33), .ZN(n1892) );
NAND2_X1 U1493 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1844), .ZN(n1890) );
NAND2_X1 U1494 ( .A1(n1893), .A2(n1894), .ZN(U298) );
NAND2_X1 U1495 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1691), .ZN(n1894) );
NAND2_X1 U1496 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1844), .ZN(n1893) );
NAND2_X1 U1497 ( .A1(n1895), .A2(n1896), .ZN(U297) );
NAND2_X1 U1498 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1691), .ZN(n1896) );
NAND2_X1 U1499 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1844), .ZN(n1895) );
NAND2_X1 U1500 ( .A1(n1897), .A2(n1898), .ZN(U296) );
NAND2_X1 U1501 ( .A1(n1899), .A2(n1844), .ZN(n1898) );
XNOR2_X1 U1502 ( .A(REG4_REG_7__SCAN_IN), .B(KEYINPUT48), .ZN(n1899) );
NAND2_X1 U1503 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1691), .ZN(n1897) );
NAND2_X1 U1504 ( .A1(n1900), .A2(n1901), .ZN(U295) );
NAND2_X1 U1505 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1691), .ZN(n1901) );
NAND2_X1 U1506 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1844), .ZN(n1900) );
NAND2_X1 U1507 ( .A1(n1902), .A2(n1903), .ZN(U294) );
NAND2_X1 U1508 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1691), .ZN(n1903) );
NAND2_X1 U1509 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1844), .ZN(n1902) );
NAND2_X1 U1510 ( .A1(n1904), .A2(n1905), .ZN(U293) );
NAND2_X1 U1511 ( .A1(n1906), .A2(n1691), .ZN(n1905) );
XNOR2_X1 U1512 ( .A(REG3_REG_4__SCAN_IN), .B(KEYINPUT24), .ZN(n1906) );
NAND2_X1 U1513 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1844), .ZN(n1904) );
NAND2_X1 U1514 ( .A1(n1907), .A2(n1908), .ZN(U292) );
NAND2_X1 U1515 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1691), .ZN(n1908) );
NAND2_X1 U1516 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1844), .ZN(n1907) );
NAND2_X1 U1517 ( .A1(n1909), .A2(n1910), .ZN(U291) );
NAND2_X1 U1518 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1691), .ZN(n1910) );
NAND2_X1 U1519 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1844), .ZN(n1909) );
NAND2_X1 U1520 ( .A1(n1911), .A2(n1912), .ZN(U290) );
NAND2_X1 U1521 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1691), .ZN(n1912) );
NAND2_X1 U1522 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1844), .ZN(n1911) );
NAND2_X1 U1523 ( .A1(n1913), .A2(n1914), .ZN(U289) );
NAND2_X1 U1524 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1691), .ZN(n1914) );
NAND2_X1 U1525 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1844), .ZN(n1913) );
NAND4_X1 U1526 ( .A1(n1915), .A2(n1916), .A3(n1917), .A4(n1918), .ZN(U288));
NAND2_X1 U1527 ( .A1(n1919), .A2(n1920), .ZN(n1918) );
NAND2_X1 U1528 ( .A1(n1921), .A2(REG4_REG_7__SCAN_IN), .ZN(n1917) );
NAND2_X1 U1529 ( .A1(n1922), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1916) );
NAND2_X1 U1530 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1844), .ZN(n1915) );
NAND4_X1 U1531 ( .A1(n1923), .A2(n1924), .A3(n1925), .A4(n1926), .ZN(U287));
NOR3_X1 U1532 ( .A1(n1927), .A2(n1928), .A3(n1929), .ZN(n1926) );
NOR3_X1 U1533 ( .A1(n1930), .A2(n1931), .A3(n1932), .ZN(n1929) );
AND2_X1 U1534 ( .A1(n1933), .A2(n1919), .ZN(n1931) );
XNOR2_X1 U1535 ( .A(KEYINPUT54), .B(n1934), .ZN(n1930) );
NOR3_X1 U1536 ( .A1(n1935), .A2(n1936), .A3(n1937), .ZN(n1928) );
AND2_X1 U1537 ( .A1(n1920), .A2(n1919), .ZN(n1927) );
NAND2_X1 U1538 ( .A1(n1938), .A2(n1939), .ZN(n1920) );
NAND3_X1 U1539 ( .A1(n1933), .A2(n1934), .A3(n1940), .ZN(n1939) );
XOR2_X1 U1540 ( .A(n1941), .B(KEYINPUT21), .Z(n1933) );
NAND3_X1 U1541 ( .A1(n1935), .A2(n1942), .A3(n1943), .ZN(n1938) );
NAND2_X1 U1542 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1844), .ZN(n1925) );
NAND2_X1 U1543 ( .A1(n1921), .A2(REG4_REG_6__SCAN_IN), .ZN(n1924) );
NAND2_X1 U1544 ( .A1(n1922), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1923) );
NAND4_X1 U1545 ( .A1(n1944), .A2(n1945), .A3(n1946), .A4(n1947), .ZN(U286));
NOR3_X1 U1546 ( .A1(n1948), .A2(n1949), .A3(n1950), .ZN(n1947) );
NOR2_X1 U1547 ( .A1(n1942), .A2(n1951), .ZN(n1950) );
NOR3_X1 U1548 ( .A1(n1932), .A2(n1952), .A3(n1953), .ZN(n1949) );
NOR2_X1 U1549 ( .A1(n1954), .A2(n1955), .ZN(n1953) );
INV_X1 U1550 ( .A(n1934), .ZN(n1952) );
NAND3_X1 U1551 ( .A1(n1956), .A2(n1957), .A3(n1955), .ZN(n1934) );
NAND2_X1 U1552 ( .A1(n1942), .A2(n1958), .ZN(n1957) );
NAND2_X1 U1553 ( .A1(n1941), .A2(n1919), .ZN(n1956) );
XOR2_X1 U1554 ( .A(n1954), .B(KEYINPUT2), .Z(n1941) );
AND2_X1 U1555 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1921), .ZN(n1948) );
XOR2_X1 U1556 ( .A(KEYINPUT4), .B(n1959), .Z(n1946) );
NOR3_X1 U1557 ( .A1(n1960), .A2(n1961), .A3(n1937), .ZN(n1959) );
NOR2_X1 U1558 ( .A1(n1962), .A2(n1963), .ZN(n1961) );
XNOR2_X1 U1559 ( .A(KEYINPUT8), .B(n1935), .ZN(n1960) );
NAND2_X1 U1560 ( .A1(n1962), .A2(n1963), .ZN(n1935) );
NAND2_X1 U1561 ( .A1(n1964), .A2(n1965), .ZN(n1963) );
INV_X1 U1562 ( .A(n1936), .ZN(n1965) );
NOR2_X1 U1563 ( .A1(n1958), .A2(n1954), .ZN(n1936) );
INV_X1 U1564 ( .A(n1942), .ZN(n1954) );
XOR2_X1 U1565 ( .A(KEYINPUT60), .B(n1966), .Z(n1964) );
NOR2_X1 U1566 ( .A1(n1919), .A2(n1942), .ZN(n1966) );
NAND2_X1 U1567 ( .A1(n1967), .A2(n1968), .ZN(n1942) );
NAND3_X1 U1568 ( .A1(n1969), .A2(n1970), .A3(n1971), .ZN(n1968) );
NAND2_X1 U1569 ( .A1(n1972), .A2(n1973), .ZN(n1971) );
NAND2_X1 U1570 ( .A1(n1974), .A2(n1975), .ZN(n1973) );
NAND2_X1 U1571 ( .A1(n1976), .A2(n1977), .ZN(n1975) );
XNOR2_X1 U1572 ( .A(KEYINPUT10), .B(n1978), .ZN(n1976) );
NAND3_X1 U1573 ( .A1(n1979), .A2(n1972), .A3(n1980), .ZN(n1967) );
NAND2_X1 U1574 ( .A1(n1969), .A2(n1970), .ZN(n1980) );
NAND3_X1 U1575 ( .A1(n1981), .A2(n1982), .A3(n1983), .ZN(n1970) );
NAND2_X1 U1576 ( .A1(DATA_IN_6_), .A2(n1984), .ZN(n1982) );
NAND2_X1 U1577 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1981) );
NAND3_X1 U1578 ( .A1(n1985), .A2(n1986), .A3(n1987), .ZN(n1969) );
XOR2_X1 U1579 ( .A(n1983), .B(KEYINPUT25), .Z(n1987) );
NAND2_X1 U1580 ( .A1(n1988), .A2(n1989), .ZN(n1983) );
NAND2_X1 U1581 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1984), .ZN(n1989) );
NAND2_X1 U1582 ( .A1(RESTART), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1988) );
NAND2_X1 U1583 ( .A1(RESTART), .A2(n1814), .ZN(n1986) );
NAND2_X1 U1584 ( .A1(n1761), .A2(n1984), .ZN(n1985) );
INV_X1 U1585 ( .A(DATA_IN_6_), .ZN(n1761) );
NAND2_X1 U1586 ( .A1(n1974), .A2(n1990), .ZN(n1979) );
NAND2_X1 U1587 ( .A1(n1977), .A2(n1978), .ZN(n1990) );
INV_X1 U1588 ( .A(n1958), .ZN(n1919) );
NAND2_X1 U1589 ( .A1(n1922), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1945) );
NAND2_X1 U1590 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1844), .ZN(n1944) );
NAND4_X1 U1591 ( .A1(n1991), .A2(n1992), .A3(n1993), .A4(n1994), .ZN(U285));
NOR3_X1 U1592 ( .A1(n1995), .A2(n1996), .A3(n1997), .ZN(n1994) );
NOR3_X1 U1593 ( .A1(n1937), .A2(n1962), .A3(n1998), .ZN(n1997) );
NOR2_X1 U1594 ( .A1(n1999), .A2(n2000), .ZN(n1998) );
AND2_X1 U1595 ( .A1(n2001), .A2(n1999), .ZN(n1962) );
XOR2_X1 U1596 ( .A(n2000), .B(KEYINPUT51), .Z(n2001) );
NOR3_X1 U1597 ( .A1(n2002), .A2(n2003), .A3(n1932), .ZN(n1996) );
NOR2_X1 U1598 ( .A1(n2004), .A2(n2000), .ZN(n2003) );
NOR2_X1 U1599 ( .A1(n2005), .A2(n2006), .ZN(n2004) );
XOR2_X1 U1600 ( .A(KEYINPUT46), .B(n1955), .Z(n2002) );
NOR3_X1 U1601 ( .A1(n2005), .A2(n2007), .A3(n2006), .ZN(n1955) );
INV_X1 U1602 ( .A(n2000), .ZN(n2007) );
NAND2_X1 U1603 ( .A1(n1958), .A2(n2008), .ZN(n2000) );
NAND2_X1 U1604 ( .A1(n2009), .A2(n2010), .ZN(n2008) );
NAND2_X1 U1605 ( .A1(n2011), .A2(n2012), .ZN(n2009) );
NAND3_X1 U1606 ( .A1(n2012), .A2(n2013), .A3(n2011), .ZN(n1958) );
NOR2_X1 U1607 ( .A1(n2013), .A2(n1951), .ZN(n1995) );
INV_X1 U1608 ( .A(n2010), .ZN(n2013) );
NAND3_X1 U1609 ( .A1(n2014), .A2(n2015), .A3(n2016), .ZN(n2010) );
OR2_X1 U1610 ( .A1(n1972), .A2(n1974), .ZN(n2016) );
OR2_X1 U1611 ( .A1(n1977), .A2(n1978), .ZN(n1972) );
NAND3_X1 U1612 ( .A1(n1974), .A2(n1978), .A3(n2017), .ZN(n2015) );
INV_X1 U1613 ( .A(n1977), .ZN(n2017) );
NAND2_X1 U1614 ( .A1(n2018), .A2(n1977), .ZN(n2014) );
NAND2_X1 U1615 ( .A1(n2019), .A2(n2020), .ZN(n1977) );
NAND2_X1 U1616 ( .A1(n2021), .A2(n2022), .ZN(n2020) );
NAND2_X1 U1617 ( .A1(n2023), .A2(n2024), .ZN(n2022) );
OR2_X1 U1618 ( .A1(n2024), .A2(n2023), .ZN(n2019) );
XOR2_X1 U1619 ( .A(n1978), .B(n1974), .Z(n2018) );
NAND2_X1 U1620 ( .A1(n2025), .A2(n2026), .ZN(n1974) );
NAND2_X1 U1621 ( .A1(RESTART), .A2(n1794), .ZN(n2026) );
NAND2_X1 U1622 ( .A1(n1782), .A2(n1984), .ZN(n2025) );
INV_X1 U1623 ( .A(DATA_IN_5_), .ZN(n1782) );
NAND3_X1 U1624 ( .A1(n2027), .A2(n2028), .A3(n2029), .ZN(n1978) );
OR2_X1 U1625 ( .A1(KEYINPUT63), .A2(REG4_REG_5__SCAN_IN), .ZN(n2029) );
NAND3_X1 U1626 ( .A1(KEYINPUT63), .A2(REG4_REG_5__SCAN_IN), .A3(n1984), .ZN(n2028) );
NAND2_X1 U1627 ( .A1(RESTART), .A2(n2030), .ZN(n2027) );
NAND2_X1 U1628 ( .A1(KEYINPUT63), .A2(n2031), .ZN(n2030) );
NAND2_X1 U1629 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1844), .ZN(n1993) );
NAND2_X1 U1630 ( .A1(n1921), .A2(REG4_REG_4__SCAN_IN), .ZN(n1992) );
NAND2_X1 U1631 ( .A1(n1922), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1991) );
NAND4_X1 U1632 ( .A1(n2032), .A2(n2033), .A3(n2034), .A4(n2035), .ZN(U284));
NOR3_X1 U1633 ( .A1(n2036), .A2(n2037), .A3(n2038), .ZN(n2035) );
NOR2_X1 U1634 ( .A1(n2012), .A2(n1951), .ZN(n2038) );
NOR2_X1 U1635 ( .A1(U280), .A2(n2039), .ZN(n2037) );
XNOR2_X1 U1636 ( .A(KEYINPUT5), .B(DATA_OUT_REG_3__SCAN_IN), .ZN(n2039) );
AND2_X1 U1637 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1922), .ZN(n2036) );
NAND2_X1 U1638 ( .A1(n1940), .A2(n2040), .ZN(n2034) );
XNOR2_X1 U1639 ( .A(n2041), .B(n2005), .ZN(n2040) );
NAND3_X1 U1640 ( .A1(n2042), .A2(n2043), .A3(n1943), .ZN(n2033) );
INV_X1 U1641 ( .A(n1999), .ZN(n2043) );
NOR2_X1 U1642 ( .A1(n2044), .A2(n2005), .ZN(n1999) );
NAND2_X1 U1643 ( .A1(n2005), .A2(n2044), .ZN(n2042) );
XOR2_X1 U1644 ( .A(n2011), .B(n2012), .Z(n2005) );
XNOR2_X1 U1645 ( .A(n2021), .B(n2045), .ZN(n2012) );
NOR2_X1 U1646 ( .A1(n2046), .A2(n2047), .ZN(n2045) );
NOR2_X1 U1647 ( .A1(n2048), .A2(n2049), .ZN(n2047) );
NOR2_X1 U1648 ( .A1(KEYINPUT31), .A2(n2023), .ZN(n2049) );
NOR2_X1 U1649 ( .A1(n2050), .A2(n2024), .ZN(n2048) );
NOR2_X1 U1650 ( .A1(KEYINPUT27), .A2(n2051), .ZN(n2050) );
NOR4_X1 U1651 ( .A1(KEYINPUT31), .A2(n2023), .A3(n2052), .A4(n2024), .ZN(n2046) );
NAND2_X1 U1652 ( .A1(n2053), .A2(n2054), .ZN(n2024) );
NAND2_X1 U1653 ( .A1(RESTART), .A2(n1801), .ZN(n2054) );
NAND2_X1 U1654 ( .A1(n1733), .A2(n1984), .ZN(n2053) );
INV_X1 U1655 ( .A(KEYINPUT27), .ZN(n2052) );
INV_X1 U1656 ( .A(n2051), .ZN(n2023) );
NAND3_X1 U1657 ( .A1(n2055), .A2(n2056), .A3(n2057), .ZN(n2051) );
NAND2_X1 U1658 ( .A1(KEYINPUT20), .A2(n1765), .ZN(n2057) );
NAND2_X1 U1659 ( .A1(RESTART), .A2(n2058), .ZN(n2056) );
NAND2_X1 U1660 ( .A1(n2059), .A2(n2060), .ZN(n2058) );
NAND2_X1 U1661 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n2061), .ZN(n2060) );
OR2_X1 U1662 ( .A1(n2062), .A2(KEYINPUT45), .ZN(n2059) );
NAND2_X1 U1663 ( .A1(n2063), .A2(n1984), .ZN(n2055) );
NAND2_X1 U1664 ( .A1(n2061), .A2(n2064), .ZN(n2063) );
NAND2_X1 U1665 ( .A1(KEYINPUT45), .A2(REG4_REG_4__SCAN_IN), .ZN(n2064) );
INV_X1 U1666 ( .A(KEYINPUT20), .ZN(n2061) );
AND2_X1 U1667 ( .A1(n2065), .A2(n2066), .ZN(n2021) );
NAND2_X1 U1668 ( .A1(n2067), .A2(n2068), .ZN(n2066) );
NAND2_X1 U1669 ( .A1(n2069), .A2(n2070), .ZN(n2068) );
XNOR2_X1 U1670 ( .A(KEYINPUT1), .B(n2071), .ZN(n2069) );
NAND2_X1 U1671 ( .A1(n2071), .A2(n2072), .ZN(n2065) );
NAND2_X1 U1672 ( .A1(n2073), .A2(n1921), .ZN(n2032) );
XNOR2_X1 U1673 ( .A(REG4_REG_3__SCAN_IN), .B(KEYINPUT15), .ZN(n2073) );
NAND4_X1 U1674 ( .A1(n2074), .A2(n2075), .A3(n2076), .A4(n2077), .ZN(U283));
NOR3_X1 U1675 ( .A1(n2078), .A2(n2079), .A3(n2080), .ZN(n2077) );
NOR3_X1 U1676 ( .A1(n1932), .A2(n2041), .A3(n2081), .ZN(n2080) );
NOR2_X1 U1677 ( .A1(n2082), .A2(n2083), .ZN(n2081) );
AND2_X1 U1678 ( .A1(n2084), .A2(n2085), .ZN(n2082) );
INV_X1 U1679 ( .A(n2006), .ZN(n2041) );
NAND3_X1 U1680 ( .A1(n2085), .A2(n2084), .A3(n2086), .ZN(n2006) );
OR2_X1 U1681 ( .A1(n2083), .A2(n2011), .ZN(n2086) );
XOR2_X1 U1682 ( .A(n2087), .B(KEYINPUT58), .Z(n2083) );
NOR3_X1 U1683 ( .A1(n1937), .A2(n2088), .A3(n2089), .ZN(n2079) );
NOR2_X1 U1684 ( .A1(n2090), .A2(n2091), .ZN(n2089) );
AND2_X1 U1685 ( .A1(n2092), .A2(n2093), .ZN(n2090) );
INV_X1 U1686 ( .A(n2044), .ZN(n2088) );
NAND3_X1 U1687 ( .A1(n2093), .A2(n2092), .A3(n2091), .ZN(n2044) );
NAND2_X1 U1688 ( .A1(n2094), .A2(n2087), .ZN(n2091) );
NAND2_X1 U1689 ( .A1(n2095), .A2(n2096), .ZN(n2087) );
INV_X1 U1690 ( .A(n2011), .ZN(n2094) );
NOR2_X1 U1691 ( .A1(n2096), .A2(n2095), .ZN(n2011) );
AND2_X1 U1692 ( .A1(n2095), .A2(n2097), .ZN(n2078) );
NAND2_X1 U1693 ( .A1(n2098), .A2(n2099), .ZN(n2095) );
NAND2_X1 U1694 ( .A1(n2070), .A2(n2100), .ZN(n2099) );
NAND3_X1 U1695 ( .A1(n2101), .A2(n2102), .A3(n2103), .ZN(n2100) );
NAND2_X1 U1696 ( .A1(KEYINPUT61), .A2(n2104), .ZN(n2103) );
NAND2_X1 U1697 ( .A1(n2071), .A2(n2105), .ZN(n2102) );
NAND2_X1 U1698 ( .A1(n2106), .A2(n2107), .ZN(n2105) );
OR2_X1 U1699 ( .A1(n2104), .A2(KEYINPUT61), .ZN(n2107) );
INV_X1 U1700 ( .A(n2067), .ZN(n2104) );
INV_X1 U1701 ( .A(KEYINPUT17), .ZN(n2106) );
NAND2_X1 U1702 ( .A1(n2108), .A2(n2109), .ZN(n2101) );
INV_X1 U1703 ( .A(n2071), .ZN(n2109) );
INV_X1 U1704 ( .A(n2072), .ZN(n2070) );
NAND2_X1 U1705 ( .A1(n2110), .A2(n2072), .ZN(n2098) );
NAND2_X1 U1706 ( .A1(n2111), .A2(n2112), .ZN(n2072) );
NAND2_X1 U1707 ( .A1(n2113), .A2(n2114), .ZN(n2112) );
OR2_X1 U1708 ( .A1(n2115), .A2(n2116), .ZN(n2113) );
NAND2_X1 U1709 ( .A1(n2116), .A2(n2115), .ZN(n2111) );
XNOR2_X1 U1710 ( .A(n2108), .B(n2071), .ZN(n2110) );
NAND2_X1 U1711 ( .A1(n2117), .A2(n2118), .ZN(n2071) );
NAND2_X1 U1712 ( .A1(RESTART), .A2(n1772), .ZN(n2118) );
NAND2_X1 U1713 ( .A1(n2119), .A2(n1984), .ZN(n2117) );
NOR2_X1 U1714 ( .A1(n2067), .A2(KEYINPUT17), .ZN(n2108) );
NAND2_X1 U1715 ( .A1(n2120), .A2(n2121), .ZN(n2067) );
NAND2_X1 U1716 ( .A1(RESTART), .A2(n1813), .ZN(n2121) );
NAND2_X1 U1717 ( .A1(n1780), .A2(n1984), .ZN(n2120) );
NAND2_X1 U1718 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1844), .ZN(n2076) );
NAND2_X1 U1719 ( .A1(n1921), .A2(REG4_REG_2__SCAN_IN), .ZN(n2075) );
NAND2_X1 U1720 ( .A1(n1922), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2074) );
NAND4_X1 U1721 ( .A1(n2122), .A2(n2123), .A3(n2124), .A4(n2125), .ZN(U282));
NOR3_X1 U1722 ( .A1(n2126), .A2(n2127), .A3(n2128), .ZN(n2125) );
NOR2_X1 U1723 ( .A1(n2129), .A2(n1937), .ZN(n2128) );
XNOR2_X1 U1724 ( .A(n2093), .B(n2092), .ZN(n2129) );
NAND3_X1 U1725 ( .A1(n2130), .A2(n2131), .A3(n2096), .ZN(n2093) );
OR2_X1 U1726 ( .A1(n2132), .A2(KEYINPUT29), .ZN(n2131) );
NAND3_X1 U1727 ( .A1(n2132), .A2(n2133), .A3(KEYINPUT29), .ZN(n2130) );
NOR2_X1 U1728 ( .A1(n2134), .A2(n2135), .ZN(n2127) );
XNOR2_X1 U1729 ( .A(KEYINPUT36), .B(n1932), .ZN(n2135) );
XOR2_X1 U1730 ( .A(n2085), .B(n2136), .Z(n2134) );
NOR2_X1 U1731 ( .A1(KEYINPUT52), .A2(n2084), .ZN(n2136) );
NAND2_X1 U1732 ( .A1(n2096), .A2(n2137), .ZN(n2085) );
NAND2_X1 U1733 ( .A1(n2132), .A2(n2133), .ZN(n2137) );
OR2_X1 U1734 ( .A1(n2133), .A2(n2132), .ZN(n2096) );
AND2_X1 U1735 ( .A1(n2132), .A2(n2097), .ZN(n2126) );
XOR2_X1 U1736 ( .A(n2138), .B(n2115), .Z(n2132) );
NAND2_X1 U1737 ( .A1(n2139), .A2(n2140), .ZN(n2115) );
NAND2_X1 U1738 ( .A1(RESTART), .A2(n1779), .ZN(n2140) );
NAND2_X1 U1739 ( .A1(n2141), .A2(n1984), .ZN(n2139) );
XNOR2_X1 U1740 ( .A(n2114), .B(n2116), .ZN(n2138) );
NAND2_X1 U1741 ( .A1(n2142), .A2(n2143), .ZN(n2116) );
NAND2_X1 U1742 ( .A1(n1740), .A2(n1984), .ZN(n2143) );
NAND2_X1 U1743 ( .A1(n2144), .A2(RESTART), .ZN(n2142) );
XNOR2_X1 U1744 ( .A(n1808), .B(KEYINPUT14), .ZN(n2144) );
NAND2_X1 U1745 ( .A1(n2145), .A2(n2146), .ZN(n2114) );
NAND2_X1 U1746 ( .A1(n2147), .A2(n2148), .ZN(n2146) );
NAND2_X1 U1747 ( .A1(n2149), .A2(n2150), .ZN(n2148) );
XNOR2_X1 U1748 ( .A(n2151), .B(n2152), .ZN(n2150) );
NAND2_X1 U1749 ( .A1(n2151), .A2(n2153), .ZN(n2145) );
NAND2_X1 U1750 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1844), .ZN(n2124) );
NAND2_X1 U1751 ( .A1(n1921), .A2(REG4_REG_1__SCAN_IN), .ZN(n2123) );
INV_X1 U1752 ( .A(n2154), .ZN(n1921) );
NAND2_X1 U1753 ( .A1(n1922), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2122) );
NAND4_X1 U1754 ( .A1(n2155), .A2(n2156), .A3(n2157), .A4(n2158), .ZN(U281));
NOR3_X1 U1755 ( .A1(n2159), .A2(n2160), .A3(n2161), .ZN(n2158) );
NOR2_X1 U1756 ( .A1(n2162), .A2(n2154), .ZN(n2161) );
NAND3_X1 U1757 ( .A1(ENABLE), .A2(n2163), .A3(AVERAGE), .ZN(n2154) );
XNOR2_X1 U1758 ( .A(KEYINPUT57), .B(n2164), .ZN(n2163) );
NOR2_X1 U1759 ( .A1(n1937), .A2(n2165), .ZN(n2160) );
XNOR2_X1 U1760 ( .A(KEYINPUT37), .B(n2092), .ZN(n2165) );
NAND2_X1 U1761 ( .A1(n2166), .A2(n2167), .ZN(n2092) );
NAND2_X1 U1762 ( .A1(n2168), .A2(n2169), .ZN(n2167) );
NAND2_X1 U1763 ( .A1(n2170), .A2(n2171), .ZN(n2169) );
NAND2_X1 U1764 ( .A1(n2172), .A2(n2170), .ZN(n2166) );
INV_X1 U1765 ( .A(KEYINPUT3), .ZN(n2170) );
INV_X1 U1766 ( .A(n1943), .ZN(n1937) );
NOR4_X1 U1767 ( .A1(n1839), .A2(n2164), .A3(n2173), .A4(AVERAGE), .ZN(n1943));
INV_X1 U1768 ( .A(ENABLE), .ZN(n1839) );
AND2_X1 U1769 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1922), .ZN(n2159) );
AND2_X1 U1770 ( .A1(n2174), .A2(n2175), .ZN(n1922) );
INV_X1 U1771 ( .A(n2164), .ZN(n2175) );
NAND3_X1 U1772 ( .A1(U280), .A2(n1984), .A3(STATO_REG_1__SCAN_IN), .ZN(n2164) );
XNOR2_X1 U1773 ( .A(ENABLE), .B(KEYINPUT28), .ZN(n2174) );
XOR2_X1 U1774 ( .A(n2176), .B(KEYINPUT9), .Z(n2157) );
NAND2_X1 U1775 ( .A1(n2097), .A2(n2168), .ZN(n2176) );
INV_X1 U1776 ( .A(n1951), .ZN(n2097) );
NAND4_X1 U1777 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2177), .A3(n2178), .A4(U280), .ZN(n1951) );
NAND2_X1 U1778 ( .A1(n2179), .A2(n1984), .ZN(n2177) );
NAND3_X1 U1779 ( .A1(n2173), .A2(n2180), .A3(ENABLE), .ZN(n2179) );
INV_X1 U1780 ( .A(AVERAGE), .ZN(n2180) );
NAND2_X1 U1781 ( .A1(n2181), .A2(n2182), .ZN(n2173) );
OR2_X1 U1782 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2182) );
NAND3_X1 U1783 ( .A1(n2183), .A2(n2184), .A3(n2185), .ZN(n2181) );
NAND2_X1 U1784 ( .A1(REG4_REG_7__SCAN_IN), .A2(DATA_IN_7_), .ZN(n2185) );
NAND3_X1 U1785 ( .A1(n2186), .A2(n2187), .A3(n2188), .ZN(n2184) );
NAND2_X1 U1786 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2188) );
NAND2_X1 U1787 ( .A1(n2189), .A2(n2190), .ZN(n2187) );
NAND2_X1 U1788 ( .A1(n2191), .A2(n2192), .ZN(n2190) );
NAND3_X1 U1789 ( .A1(n2193), .A2(n2194), .A3(n2195), .ZN(n2192) );
NAND2_X1 U1790 ( .A1(n1733), .A2(n2062), .ZN(n2195) );
INV_X1 U1791 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2062) );
INV_X1 U1792 ( .A(DATA_IN_4_), .ZN(n1733) );
NAND3_X1 U1793 ( .A1(n2196), .A2(n2197), .A3(n2198), .ZN(n2194) );
NAND2_X1 U1794 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2198) );
NAND3_X1 U1795 ( .A1(n2199), .A2(n2200), .A3(n2201), .ZN(n2197) );
NAND2_X1 U1796 ( .A1(n1740), .A2(n2141), .ZN(n2201) );
INV_X1 U1797 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2141) );
INV_X1 U1798 ( .A(DATA_IN_2_), .ZN(n1740) );
NAND2_X1 U1799 ( .A1(n2202), .A2(n2203), .ZN(n2200) );
NAND2_X1 U1800 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2203) );
XOR2_X1 U1801 ( .A(KEYINPUT56), .B(n2204), .Z(n2202) );
NAND2_X1 U1802 ( .A1(n1712), .A2(n2205), .ZN(n2199) );
NAND2_X1 U1803 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2196) );
NAND2_X1 U1804 ( .A1(n1780), .A2(n2119), .ZN(n2193) );
INV_X1 U1805 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2119) );
INV_X1 U1806 ( .A(DATA_IN_3_), .ZN(n1780) );
NAND2_X1 U1807 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2191) );
XOR2_X1 U1808 ( .A(KEYINPUT43), .B(n2206), .Z(n2189) );
NOR2_X1 U1809 ( .A1(DATA_IN_5_), .A2(REG4_REG_5__SCAN_IN), .ZN(n2206) );
NAND2_X1 U1810 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2186) );
OR2_X1 U1811 ( .A1(DATA_IN_6_), .A2(REG4_REG_6__SCAN_IN), .ZN(n2183) );
OR2_X1 U1812 ( .A1(n2084), .A2(n1932), .ZN(n2156) );
INV_X1 U1813 ( .A(n1940), .ZN(n1932) );
NOR3_X1 U1814 ( .A1(n1749), .A2(n1844), .A3(n2178), .ZN(n1940) );
NAND2_X1 U1815 ( .A1(n2207), .A2(RESTART), .ZN(n2178) );
XOR2_X1 U1816 ( .A(n2208), .B(KEYINPUT40), .Z(n2207) );
NAND2_X1 U1817 ( .A1(n2209), .A2(n2210), .ZN(n2208) );
NAND2_X1 U1818 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2210) );
NAND3_X1 U1819 ( .A1(n2211), .A2(n2212), .A3(n2213), .ZN(n2209) );
OR2_X1 U1820 ( .A1(RMAX_REG_7__SCAN_IN), .A2(RMIN_REG_7__SCAN_IN), .ZN(n2213) );
NAND2_X1 U1821 ( .A1(KEYINPUT44), .A2(n2214), .ZN(n2212) );
NAND2_X1 U1822 ( .A1(n2215), .A2(n2216), .ZN(n2214) );
NAND2_X1 U1823 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n2217), .ZN(n2216) );
NAND2_X1 U1824 ( .A1(n1814), .A2(n2218), .ZN(n2217) );
OR2_X1 U1825 ( .A1(n2218), .A2(n1814), .ZN(n2215) );
INV_X1 U1826 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1814) );
NAND3_X1 U1827 ( .A1(n2219), .A2(n1783), .A3(n2220), .ZN(n2211) );
INV_X1 U1828 ( .A(KEYINPUT44), .ZN(n2220) );
INV_X1 U1829 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1783) );
XNOR2_X1 U1830 ( .A(RMAX_REG_6__SCAN_IN), .B(n2218), .ZN(n2219) );
NAND2_X1 U1831 ( .A1(n2221), .A2(n2222), .ZN(n2218) );
NAND2_X1 U1832 ( .A1(n1794), .A2(n2031), .ZN(n2222) );
INV_X1 U1833 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n2031) );
INV_X1 U1834 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1794) );
NAND3_X1 U1835 ( .A1(n2223), .A2(n2224), .A3(n2225), .ZN(n2221) );
NAND2_X1 U1836 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2225) );
NAND3_X1 U1837 ( .A1(n2226), .A2(n2227), .A3(n2228), .ZN(n2224) );
NAND2_X1 U1838 ( .A1(n1801), .A2(n1765), .ZN(n2228) );
INV_X1 U1839 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1765) );
INV_X1 U1840 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1801) );
NAND3_X1 U1841 ( .A1(n2229), .A2(n2230), .A3(n2231), .ZN(n2227) );
NAND2_X1 U1842 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2231) );
NAND3_X1 U1843 ( .A1(n2232), .A2(n2233), .A3(n2234), .ZN(n2230) );
NAND2_X1 U1844 ( .A1(n1808), .A2(n1779), .ZN(n2234) );
INV_X1 U1845 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1779) );
INV_X1 U1846 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1808) );
NAND2_X1 U1847 ( .A1(n2235), .A2(n1778), .ZN(n2233) );
OR2_X1 U1848 ( .A1(n2236), .A2(n1811), .ZN(n2235) );
NAND2_X1 U1849 ( .A1(n2236), .A2(n1811), .ZN(n2232) );
NAND2_X1 U1850 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2229) );
NAND2_X1 U1851 ( .A1(n1813), .A2(n1772), .ZN(n2226) );
INV_X1 U1852 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1772) );
INV_X1 U1853 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1813) );
NAND2_X1 U1854 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2223) );
NAND3_X1 U1855 ( .A1(n2237), .A2(n2238), .A3(n2133), .ZN(n2084) );
INV_X1 U1856 ( .A(n2172), .ZN(n2133) );
NOR2_X1 U1857 ( .A1(n2168), .A2(n2239), .ZN(n2172) );
OR2_X1 U1858 ( .A1(n2239), .A2(KEYINPUT12), .ZN(n2238) );
NAND3_X1 U1859 ( .A1(n2239), .A2(n2168), .A3(KEYINPUT12), .ZN(n2237) );
XOR2_X1 U1860 ( .A(n2151), .B(n2240), .Z(n2168) );
NOR2_X1 U1861 ( .A1(n2152), .A2(n2241), .ZN(n2240) );
XNOR2_X1 U1862 ( .A(n2147), .B(n2149), .ZN(n2241) );
INV_X1 U1863 ( .A(n2153), .ZN(n2149) );
NAND2_X1 U1864 ( .A1(n2242), .A2(n2243), .ZN(n2153) );
NAND2_X1 U1865 ( .A1(RESTART), .A2(n1811), .ZN(n2243) );
INV_X1 U1866 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1811) );
NAND2_X1 U1867 ( .A1(n1712), .A2(n1984), .ZN(n2242) );
INV_X1 U1868 ( .A(DATA_IN_1_), .ZN(n1712) );
NAND2_X1 U1869 ( .A1(n2244), .A2(n2245), .ZN(n2147) );
NAND2_X1 U1870 ( .A1(RESTART), .A2(n1778), .ZN(n2245) );
INV_X1 U1871 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1778) );
NAND2_X1 U1872 ( .A1(n2205), .A2(n1984), .ZN(n2244) );
INV_X1 U1873 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2205) );
INV_X1 U1874 ( .A(KEYINPUT49), .ZN(n2152) );
INV_X1 U1875 ( .A(n2171), .ZN(n2239) );
NAND3_X1 U1876 ( .A1(n2246), .A2(n2247), .A3(n2151), .ZN(n2171) );
NAND2_X1 U1877 ( .A1(n2248), .A2(n2249), .ZN(n2151) );
NAND2_X1 U1878 ( .A1(RESTART), .A2(n2236), .ZN(n2249) );
NAND2_X1 U1879 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2236) );
OR2_X1 U1880 ( .A1(n2204), .A2(RESTART), .ZN(n2248) );
NOR2_X1 U1881 ( .A1(n2162), .A2(n1777), .ZN(n2204) );
NAND3_X1 U1882 ( .A1(n1777), .A2(n2162), .A3(n1984), .ZN(n2247) );
INV_X1 U1883 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2162) );
INV_X1 U1884 ( .A(DATA_IN_0_), .ZN(n1777) );
OR3_X1 U1885 ( .A1(RMAX_REG_0__SCAN_IN), .A2(RMIN_REG_0__SCAN_IN), .A3(n1984), .ZN(n2246) );
INV_X1 U1886 ( .A(RESTART), .ZN(n1984) );
NAND2_X1 U1887 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1844), .ZN(n2155) );
NAND2_X1 U1888 ( .A1(n1690), .A2(n2250), .ZN(U280) );
NAND2_X1 U1889 ( .A1(STATO_REG_0__SCAN_IN), .A2(n1749), .ZN(n2250) );
INV_X1 U1890 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1749) );
endmodule


