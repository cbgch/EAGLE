//Key = 0100111100111000000000110100001011011011011000011110101101100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333;

XOR2_X1 U729 ( .A(G107), .B(n1010), .Z(G9) );
NOR2_X1 U730 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
XOR2_X1 U732 ( .A(n1017), .B(KEYINPUT35), .Z(n1015) );
NAND4_X1 U733 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NAND2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND3_X1 U736 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1020) );
NAND4_X1 U737 ( .A1(n1029), .A2(n1025), .A3(n1030), .A4(n1031), .ZN(n1027) );
NAND2_X1 U738 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1024), .A2(n1036), .ZN(n1026) );
XNOR2_X1 U741 ( .A(n1037), .B(n1038), .ZN(n1019) );
NAND3_X1 U742 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1013) );
NAND2_X1 U743 ( .A1(n1018), .A2(n1042), .ZN(n1041) );
NAND2_X1 U744 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U745 ( .A1(n1045), .A2(n1025), .A3(n1024), .ZN(n1044) );
NAND2_X1 U746 ( .A1(n1046), .A2(n1047), .ZN(n1043) );
NAND3_X1 U747 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NAND2_X1 U748 ( .A1(n1024), .A2(n1051), .ZN(n1050) );
NAND4_X1 U749 ( .A1(n1029), .A2(n1052), .A3(n1025), .A4(n1034), .ZN(n1049) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1048) );
INV_X1 U751 ( .A(n1055), .ZN(n1018) );
NOR3_X1 U752 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1011) );
INV_X1 U753 ( .A(n1039), .ZN(n1056) );
NAND4_X1 U754 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1039) );
NOR4_X1 U755 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
XNOR2_X1 U756 ( .A(n1065), .B(n1066), .ZN(n1064) );
NOR2_X1 U757 ( .A1(KEYINPUT24), .A2(n1067), .ZN(n1066) );
XNOR2_X1 U758 ( .A(n1068), .B(n1069), .ZN(n1061) );
NOR2_X1 U759 ( .A1(n1022), .A2(n1032), .ZN(n1059) );
XOR2_X1 U760 ( .A(n1070), .B(n1071), .Z(n1058) );
XNOR2_X1 U761 ( .A(G472), .B(KEYINPUT47), .ZN(n1071) );
XOR2_X1 U762 ( .A(n1072), .B(n1073), .Z(n1057) );
NAND2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
XOR2_X1 U764 ( .A(KEYINPUT9), .B(KEYINPUT55), .Z(n1074) );
XOR2_X1 U765 ( .A(n1076), .B(n1077), .Z(G72) );
NOR3_X1 U766 ( .A1(n1040), .A2(KEYINPUT40), .A3(n1078), .ZN(n1077) );
AND2_X1 U767 ( .A1(G227), .A2(G900), .ZN(n1078) );
NAND2_X1 U768 ( .A1(n1079), .A2(n1080), .ZN(n1076) );
NAND3_X1 U769 ( .A1(n1081), .A2(n1082), .A3(n1016), .ZN(n1080) );
NAND2_X1 U770 ( .A1(G953), .A2(n1083), .ZN(n1082) );
NAND2_X1 U771 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U772 ( .A1(G900), .A2(n1086), .ZN(n1084) );
NAND2_X1 U773 ( .A1(n1087), .A2(n1040), .ZN(n1081) );
OR2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1087) );
INV_X1 U775 ( .A(KEYINPUT4), .ZN(n1085) );
NAND2_X1 U776 ( .A1(n1086), .A2(n1088), .ZN(n1079) );
NAND2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U778 ( .A1(G900), .A2(n1091), .ZN(n1090) );
NAND2_X1 U779 ( .A1(n1016), .A2(n1092), .ZN(n1091) );
NAND2_X1 U780 ( .A1(KEYINPUT4), .A2(G953), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1093), .A2(n1040), .ZN(n1089) );
NAND2_X1 U782 ( .A1(KEYINPUT4), .A2(n1016), .ZN(n1093) );
XOR2_X1 U783 ( .A(n1094), .B(n1095), .Z(n1086) );
XNOR2_X1 U784 ( .A(G125), .B(n1096), .ZN(n1095) );
NAND2_X1 U785 ( .A1(KEYINPUT7), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U786 ( .A(n1098), .B(n1099), .ZN(n1094) );
XOR2_X1 U787 ( .A(n1100), .B(n1101), .Z(G69) );
NOR2_X1 U788 ( .A1(n1102), .A2(n1040), .ZN(n1101) );
NOR2_X1 U789 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1100) );
XOR2_X1 U791 ( .A(KEYINPUT29), .B(KEYINPUT16), .Z(n1106) );
XOR2_X1 U792 ( .A(n1107), .B(n1108), .Z(n1105) );
AND2_X1 U793 ( .A1(n1014), .A2(n1040), .ZN(n1108) );
NAND2_X1 U794 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NAND2_X1 U795 ( .A1(G953), .A2(n1104), .ZN(n1110) );
XOR2_X1 U796 ( .A(n1111), .B(n1112), .Z(n1109) );
XOR2_X1 U797 ( .A(KEYINPUT26), .B(n1113), .Z(n1112) );
NOR2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(G66) );
XNOR2_X1 U799 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U800 ( .A1(n1118), .A2(G217), .ZN(n1116) );
NOR2_X1 U801 ( .A1(n1114), .A2(n1119), .ZN(G63) );
XOR2_X1 U802 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U803 ( .A1(n1118), .A2(G478), .ZN(n1120) );
NOR2_X1 U804 ( .A1(n1114), .A2(n1122), .ZN(G60) );
XOR2_X1 U805 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U806 ( .A1(n1118), .A2(G475), .ZN(n1123) );
XOR2_X1 U807 ( .A(G104), .B(n1125), .Z(G6) );
NOR3_X1 U808 ( .A1(n1126), .A2(KEYINPUT21), .A3(n1127), .ZN(n1125) );
NOR2_X1 U809 ( .A1(n1114), .A2(n1128), .ZN(G57) );
XOR2_X1 U810 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U811 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U812 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U813 ( .A1(n1118), .A2(G472), .ZN(n1133) );
XOR2_X1 U814 ( .A(n1135), .B(n1136), .Z(n1129) );
XNOR2_X1 U815 ( .A(n1137), .B(n1138), .ZN(n1136) );
NAND2_X1 U816 ( .A1(KEYINPUT58), .A2(n1139), .ZN(n1137) );
XNOR2_X1 U817 ( .A(n1140), .B(n1141), .ZN(n1139) );
XOR2_X1 U818 ( .A(KEYINPUT43), .B(KEYINPUT1), .Z(n1141) );
XNOR2_X1 U819 ( .A(G101), .B(n1142), .ZN(n1135) );
NOR2_X1 U820 ( .A1(n1114), .A2(n1143), .ZN(G54) );
XOR2_X1 U821 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U822 ( .A(n1146), .B(n1147), .ZN(n1145) );
XOR2_X1 U823 ( .A(n1148), .B(n1149), .Z(n1144) );
XOR2_X1 U824 ( .A(KEYINPUT12), .B(n1150), .Z(n1149) );
NOR2_X1 U825 ( .A1(KEYINPUT20), .A2(n1151), .ZN(n1150) );
NOR3_X1 U826 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
XOR2_X1 U827 ( .A(KEYINPUT61), .B(n1155), .Z(n1152) );
NOR2_X1 U828 ( .A1(n1156), .A2(n1157), .ZN(n1148) );
XOR2_X1 U829 ( .A(n1158), .B(KEYINPUT25), .Z(n1157) );
NAND2_X1 U830 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U831 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
AND3_X1 U832 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1159) );
NAND2_X1 U833 ( .A1(G140), .A2(n1164), .ZN(n1163) );
OR3_X1 U834 ( .A1(n1164), .A2(G140), .A3(KEYINPUT0), .ZN(n1162) );
NAND2_X1 U835 ( .A1(KEYINPUT33), .A2(n1165), .ZN(n1164) );
NAND2_X1 U836 ( .A1(KEYINPUT0), .A2(G110), .ZN(n1161) );
NOR2_X1 U837 ( .A1(n1040), .A2(G952), .ZN(n1114) );
NOR2_X1 U838 ( .A1(n1166), .A2(n1167), .ZN(G51) );
XOR2_X1 U839 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U841 ( .A1(n1118), .A2(n1172), .ZN(n1170) );
INV_X1 U842 ( .A(n1075), .ZN(n1172) );
NOR2_X1 U843 ( .A1(n1153), .A2(n1155), .ZN(n1118) );
NOR2_X1 U844 ( .A1(n1173), .A2(n1016), .ZN(n1155) );
NAND4_X1 U845 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1016) );
AND3_X1 U846 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
NAND2_X1 U847 ( .A1(n1024), .A2(n1181), .ZN(n1176) );
NAND3_X1 U848 ( .A1(n1036), .A2(n1052), .A3(n1182), .ZN(n1175) );
NAND2_X1 U849 ( .A1(n1183), .A2(n1184), .ZN(n1174) );
NAND3_X1 U850 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1184) );
NAND2_X1 U851 ( .A1(n1181), .A2(n1188), .ZN(n1187) );
NAND2_X1 U852 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
OR2_X1 U853 ( .A1(n1126), .A2(KEYINPUT28), .ZN(n1190) );
XNOR2_X1 U854 ( .A(KEYINPUT6), .B(n1035), .ZN(n1189) );
NAND4_X1 U855 ( .A1(n1036), .A2(n1052), .A3(n1046), .A4(n1191), .ZN(n1186) );
NAND2_X1 U856 ( .A1(KEYINPUT28), .A2(n1192), .ZN(n1185) );
NAND2_X1 U857 ( .A1(n1181), .A2(n1052), .ZN(n1192) );
XNOR2_X1 U858 ( .A(n1014), .B(KEYINPUT11), .ZN(n1173) );
NAND4_X1 U859 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1014) );
NOR4_X1 U860 ( .A1(n1197), .A2(n1198), .A3(n1010), .A4(n1199), .ZN(n1196) );
INV_X1 U861 ( .A(n1200), .ZN(n1199) );
NOR2_X1 U862 ( .A1(n1035), .A2(n1127), .ZN(n1010) );
NAND3_X1 U863 ( .A1(n1054), .A2(n1201), .A3(n1045), .ZN(n1127) );
INV_X1 U864 ( .A(n1202), .ZN(n1198) );
NOR2_X1 U865 ( .A1(n1203), .A2(n1204), .ZN(n1195) );
NOR3_X1 U866 ( .A1(n1205), .A2(n1206), .A3(n1035), .ZN(n1204) );
XNOR2_X1 U867 ( .A(n1051), .B(KEYINPUT59), .ZN(n1206) );
NAND3_X1 U868 ( .A1(n1207), .A2(n1201), .A3(n1045), .ZN(n1194) );
NAND2_X1 U869 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND4_X1 U870 ( .A1(n1036), .A2(n1053), .A3(n1210), .A4(n1211), .ZN(n1209) );
NAND2_X1 U871 ( .A1(n1052), .A2(n1054), .ZN(n1208) );
AND2_X1 U872 ( .A1(n1183), .A2(n1025), .ZN(n1054) );
OR2_X1 U873 ( .A1(n1211), .A2(n1212), .ZN(n1193) );
INV_X1 U874 ( .A(KEYINPUT52), .ZN(n1211) );
XOR2_X1 U875 ( .A(n1213), .B(n1214), .Z(n1168) );
NAND2_X1 U876 ( .A1(KEYINPUT36), .A2(n1215), .ZN(n1213) );
NOR2_X1 U877 ( .A1(G952), .A2(n1216), .ZN(n1166) );
XNOR2_X1 U878 ( .A(KEYINPUT30), .B(n1040), .ZN(n1216) );
XNOR2_X1 U879 ( .A(G146), .B(n1217), .ZN(G48) );
NAND2_X1 U880 ( .A1(n1218), .A2(n1052), .ZN(n1217) );
XOR2_X1 U881 ( .A(n1178), .B(n1219), .Z(G45) );
NOR2_X1 U882 ( .A1(G143), .A2(KEYINPUT15), .ZN(n1219) );
NAND4_X1 U883 ( .A1(n1045), .A2(n1183), .A3(n1051), .A4(n1220), .ZN(n1178) );
AND3_X1 U884 ( .A1(n1221), .A2(n1191), .A3(n1062), .ZN(n1220) );
XNOR2_X1 U885 ( .A(G140), .B(n1222), .ZN(G42) );
NAND4_X1 U886 ( .A1(KEYINPUT49), .A2(n1182), .A3(n1036), .A4(n1052), .ZN(n1222) );
XNOR2_X1 U887 ( .A(n1097), .B(n1223), .ZN(G39) );
AND2_X1 U888 ( .A1(n1181), .A2(n1024), .ZN(n1223) );
NOR3_X1 U889 ( .A1(n1033), .A2(n1032), .A3(n1224), .ZN(n1024) );
INV_X1 U890 ( .A(n1053), .ZN(n1033) );
INV_X1 U891 ( .A(n1225), .ZN(n1181) );
XOR2_X1 U892 ( .A(n1180), .B(n1226), .Z(G36) );
NAND2_X1 U893 ( .A1(KEYINPUT32), .A2(G134), .ZN(n1226) );
NAND2_X1 U894 ( .A1(n1227), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U895 ( .A(G131), .B(n1179), .ZN(G33) );
NAND3_X1 U896 ( .A1(n1052), .A2(n1051), .A3(n1182), .ZN(n1179) );
AND4_X1 U897 ( .A1(n1029), .A2(n1045), .A3(n1191), .A4(n1034), .ZN(n1182) );
XOR2_X1 U898 ( .A(n1228), .B(n1229), .Z(G30) );
AND2_X1 U899 ( .A1(n1230), .A2(n1218), .ZN(n1229) );
NOR2_X1 U900 ( .A1(n1225), .A2(n1210), .ZN(n1218) );
INV_X1 U901 ( .A(n1183), .ZN(n1210) );
NAND4_X1 U902 ( .A1(n1231), .A2(n1045), .A3(n1191), .A4(n1063), .ZN(n1225) );
NOR2_X1 U903 ( .A1(KEYINPUT19), .A2(n1232), .ZN(n1228) );
INV_X1 U904 ( .A(G128), .ZN(n1232) );
XOR2_X1 U905 ( .A(G101), .B(n1203), .Z(G3) );
AND2_X1 U906 ( .A1(n1233), .A2(n1051), .ZN(n1203) );
INV_X1 U907 ( .A(n1234), .ZN(n1051) );
XNOR2_X1 U908 ( .A(G125), .B(n1235), .ZN(G27) );
NAND3_X1 U909 ( .A1(n1236), .A2(n1052), .A3(n1237), .ZN(n1235) );
AND3_X1 U910 ( .A1(n1183), .A2(n1191), .A3(n1046), .ZN(n1237) );
NAND2_X1 U911 ( .A1(n1055), .A2(n1238), .ZN(n1191) );
NAND4_X1 U912 ( .A1(G902), .A2(G953), .A3(n1239), .A4(n1240), .ZN(n1238) );
INV_X1 U913 ( .A(G900), .ZN(n1240) );
INV_X1 U914 ( .A(n1126), .ZN(n1052) );
XNOR2_X1 U915 ( .A(n1036), .B(KEYINPUT22), .ZN(n1236) );
XNOR2_X1 U916 ( .A(G122), .B(n1202), .ZN(G24) );
NAND4_X1 U917 ( .A1(n1241), .A2(n1025), .A3(n1221), .A4(n1062), .ZN(n1202) );
NOR2_X1 U918 ( .A1(n1063), .A2(n1231), .ZN(n1025) );
XNOR2_X1 U919 ( .A(G119), .B(n1200), .ZN(G21) );
NAND4_X1 U920 ( .A1(n1053), .A2(n1241), .A3(n1231), .A4(n1063), .ZN(n1200) );
XNOR2_X1 U921 ( .A(n1242), .B(n1243), .ZN(G18) );
AND2_X1 U922 ( .A1(n1241), .A2(n1227), .ZN(n1243) );
NOR2_X1 U923 ( .A1(n1234), .A2(n1035), .ZN(n1227) );
INV_X1 U924 ( .A(n1230), .ZN(n1035) );
NOR2_X1 U925 ( .A1(n1062), .A2(n1244), .ZN(n1230) );
INV_X1 U926 ( .A(n1205), .ZN(n1241) );
XOR2_X1 U927 ( .A(n1197), .B(n1245), .Z(G15) );
NOR2_X1 U928 ( .A1(KEYINPUT56), .A2(n1246), .ZN(n1245) );
NOR3_X1 U929 ( .A1(n1205), .A2(n1234), .A3(n1126), .ZN(n1197) );
NAND2_X1 U930 ( .A1(n1244), .A2(n1062), .ZN(n1126) );
INV_X1 U931 ( .A(n1221), .ZN(n1244) );
NAND2_X1 U932 ( .A1(n1231), .A2(n1247), .ZN(n1234) );
XOR2_X1 U933 ( .A(KEYINPUT34), .B(n1248), .Z(n1247) );
NAND3_X1 U934 ( .A1(n1046), .A2(n1201), .A3(n1183), .ZN(n1205) );
NAND2_X1 U935 ( .A1(n1249), .A2(n1250), .ZN(n1046) );
NAND3_X1 U936 ( .A1(n1038), .A2(n1028), .A3(n1037), .ZN(n1250) );
INV_X1 U937 ( .A(KEYINPUT8), .ZN(n1037) );
NAND2_X1 U938 ( .A1(KEYINPUT8), .A2(n1045), .ZN(n1249) );
XOR2_X1 U939 ( .A(n1212), .B(n1251), .Z(G12) );
NAND2_X1 U940 ( .A1(KEYINPUT50), .A2(G110), .ZN(n1251) );
NAND2_X1 U941 ( .A1(n1036), .A2(n1233), .ZN(n1212) );
AND4_X1 U942 ( .A1(n1053), .A2(n1045), .A3(n1183), .A4(n1201), .ZN(n1233) );
NAND2_X1 U943 ( .A1(n1252), .A2(n1055), .ZN(n1201) );
NAND3_X1 U944 ( .A1(n1239), .A2(n1040), .A3(G952), .ZN(n1055) );
NAND4_X1 U945 ( .A1(G953), .A2(n1253), .A3(n1239), .A4(n1104), .ZN(n1252) );
INV_X1 U946 ( .A(G898), .ZN(n1104) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1239) );
XNOR2_X1 U948 ( .A(KEYINPUT51), .B(n1153), .ZN(n1253) );
NOR2_X1 U949 ( .A1(n1029), .A2(n1032), .ZN(n1183) );
INV_X1 U950 ( .A(n1034), .ZN(n1032) );
NAND2_X1 U951 ( .A1(G214), .A2(n1254), .ZN(n1034) );
INV_X1 U952 ( .A(n1224), .ZN(n1029) );
XOR2_X1 U953 ( .A(n1073), .B(n1075), .Z(n1224) );
NAND2_X1 U954 ( .A1(G210), .A2(n1254), .ZN(n1075) );
NAND2_X1 U955 ( .A1(n1255), .A2(n1153), .ZN(n1254) );
NAND2_X1 U956 ( .A1(n1256), .A2(n1153), .ZN(n1073) );
XOR2_X1 U957 ( .A(n1257), .B(n1215), .Z(n1256) );
XNOR2_X1 U958 ( .A(n1140), .B(n1258), .ZN(n1215) );
XOR2_X1 U959 ( .A(KEYINPUT38), .B(G125), .Z(n1258) );
INV_X1 U960 ( .A(n1259), .ZN(n1140) );
XNOR2_X1 U961 ( .A(n1214), .B(n1171), .ZN(n1257) );
XOR2_X1 U962 ( .A(n1111), .B(n1260), .Z(n1171) );
NOR2_X1 U963 ( .A1(n1113), .A2(KEYINPUT63), .ZN(n1260) );
AND2_X1 U964 ( .A1(n1261), .A2(n1262), .ZN(n1113) );
NAND2_X1 U965 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XNOR2_X1 U966 ( .A(KEYINPUT41), .B(n1246), .ZN(n1264) );
INV_X1 U967 ( .A(G113), .ZN(n1246) );
XNOR2_X1 U968 ( .A(G119), .B(n1265), .ZN(n1263) );
NAND2_X1 U969 ( .A1(G113), .A2(n1266), .ZN(n1261) );
XNOR2_X1 U970 ( .A(n1267), .B(n1265), .ZN(n1266) );
NOR2_X1 U971 ( .A1(KEYINPUT13), .A2(n1268), .ZN(n1265) );
XNOR2_X1 U972 ( .A(G116), .B(KEYINPUT44), .ZN(n1268) );
XOR2_X1 U973 ( .A(n1269), .B(n1270), .Z(n1111) );
XNOR2_X1 U974 ( .A(n1271), .B(n1272), .ZN(n1270) );
NOR2_X1 U975 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U976 ( .A(KEYINPUT17), .B(KEYINPUT14), .Z(n1274) );
INV_X1 U977 ( .A(G122), .ZN(n1271) );
NOR2_X1 U978 ( .A1(n1103), .A2(G953), .ZN(n1214) );
INV_X1 U979 ( .A(G224), .ZN(n1103) );
NOR2_X1 U980 ( .A1(n1038), .A2(n1022), .ZN(n1045) );
INV_X1 U981 ( .A(n1028), .ZN(n1022) );
NAND2_X1 U982 ( .A1(G221), .A2(n1275), .ZN(n1028) );
NAND2_X1 U983 ( .A1(G234), .A2(n1153), .ZN(n1275) );
XNOR2_X1 U984 ( .A(n1068), .B(n1276), .ZN(n1038) );
NOR2_X1 U985 ( .A1(KEYINPUT18), .A2(n1069), .ZN(n1276) );
XOR2_X1 U986 ( .A(n1154), .B(KEYINPUT10), .Z(n1069) );
INV_X1 U987 ( .A(G469), .ZN(n1154) );
NAND2_X1 U988 ( .A1(n1277), .A2(n1278), .ZN(n1068) );
XNOR2_X1 U989 ( .A(KEYINPUT39), .B(n1153), .ZN(n1278) );
XOR2_X1 U990 ( .A(n1279), .B(n1280), .Z(n1277) );
XNOR2_X1 U991 ( .A(n1160), .B(n1269), .ZN(n1280) );
XNOR2_X1 U992 ( .A(n1165), .B(n1146), .ZN(n1269) );
XOR2_X1 U993 ( .A(G107), .B(G101), .Z(n1146) );
INV_X1 U994 ( .A(G110), .ZN(n1165) );
NAND2_X1 U995 ( .A1(G227), .A2(n1040), .ZN(n1160) );
XOR2_X1 U996 ( .A(n1147), .B(n1099), .Z(n1279) );
XOR2_X1 U997 ( .A(KEYINPUT12), .B(G140), .Z(n1099) );
XOR2_X1 U998 ( .A(n1281), .B(n1273), .Z(n1147) );
XNOR2_X1 U999 ( .A(n1282), .B(KEYINPUT57), .ZN(n1273) );
NOR2_X1 U1000 ( .A1(n1221), .A2(n1062), .ZN(n1053) );
XNOR2_X1 U1001 ( .A(n1283), .B(G475), .ZN(n1062) );
NAND2_X1 U1002 ( .A1(n1124), .A2(n1153), .ZN(n1283) );
XOR2_X1 U1003 ( .A(n1284), .B(n1285), .Z(n1124) );
XOR2_X1 U1004 ( .A(n1282), .B(n1286), .Z(n1285) );
XNOR2_X1 U1005 ( .A(n1287), .B(n1288), .ZN(n1286) );
NOR2_X1 U1006 ( .A1(KEYINPUT37), .A2(n1289), .ZN(n1288) );
XOR2_X1 U1007 ( .A(n1290), .B(G131), .Z(n1289) );
NAND2_X1 U1008 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NAND4_X1 U1009 ( .A1(G214), .A2(G143), .A3(n1255), .A4(n1040), .ZN(n1292) );
NAND2_X1 U1010 ( .A1(n1293), .A2(n1294), .ZN(n1291) );
NAND3_X1 U1011 ( .A1(n1255), .A2(n1040), .A3(G214), .ZN(n1294) );
XNOR2_X1 U1012 ( .A(G143), .B(KEYINPUT53), .ZN(n1293) );
XNOR2_X1 U1013 ( .A(G104), .B(KEYINPUT23), .ZN(n1282) );
XOR2_X1 U1014 ( .A(n1295), .B(n1296), .Z(n1284) );
XOR2_X1 U1015 ( .A(KEYINPUT3), .B(G125), .Z(n1296) );
XNOR2_X1 U1016 ( .A(G113), .B(G122), .ZN(n1295) );
XOR2_X1 U1017 ( .A(n1065), .B(n1067), .Z(n1221) );
INV_X1 U1018 ( .A(G478), .ZN(n1067) );
NAND2_X1 U1019 ( .A1(n1121), .A2(n1153), .ZN(n1065) );
XNOR2_X1 U1020 ( .A(n1297), .B(n1298), .ZN(n1121) );
XNOR2_X1 U1021 ( .A(n1299), .B(n1300), .ZN(n1298) );
XOR2_X1 U1022 ( .A(n1301), .B(n1302), .Z(n1300) );
NOR3_X1 U1023 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1302) );
INV_X1 U1024 ( .A(G234), .ZN(n1305) );
XNOR2_X1 U1025 ( .A(KEYINPUT31), .B(n1040), .ZN(n1303) );
NAND2_X1 U1026 ( .A1(KEYINPUT54), .A2(n1242), .ZN(n1301) );
INV_X1 U1027 ( .A(G116), .ZN(n1242) );
XOR2_X1 U1028 ( .A(n1306), .B(n1307), .Z(n1297) );
XOR2_X1 U1029 ( .A(KEYINPUT42), .B(G134), .Z(n1307) );
XNOR2_X1 U1030 ( .A(G107), .B(G122), .ZN(n1306) );
NOR2_X1 U1031 ( .A1(n1231), .A2(n1248), .ZN(n1036) );
INV_X1 U1032 ( .A(n1063), .ZN(n1248) );
NAND3_X1 U1033 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1063) );
NAND2_X1 U1034 ( .A1(n1311), .A2(n1117), .ZN(n1310) );
OR3_X1 U1035 ( .A1(n1117), .A2(n1311), .A3(G902), .ZN(n1309) );
NOR2_X1 U1036 ( .A1(n1304), .A2(G234), .ZN(n1311) );
INV_X1 U1037 ( .A(G217), .ZN(n1304) );
XNOR2_X1 U1038 ( .A(n1312), .B(n1313), .ZN(n1117) );
XOR2_X1 U1039 ( .A(n1287), .B(n1314), .Z(n1313) );
XOR2_X1 U1040 ( .A(n1315), .B(n1316), .Z(n1314) );
AND3_X1 U1041 ( .A1(G221), .A2(n1040), .A3(G234), .ZN(n1316) );
NOR2_X1 U1042 ( .A1(KEYINPUT45), .A2(G125), .ZN(n1315) );
XOR2_X1 U1043 ( .A(G146), .B(G140), .Z(n1287) );
XOR2_X1 U1044 ( .A(n1317), .B(n1318), .Z(n1312) );
XNOR2_X1 U1045 ( .A(n1267), .B(G110), .ZN(n1318) );
XNOR2_X1 U1046 ( .A(G128), .B(G137), .ZN(n1317) );
NAND2_X1 U1047 ( .A1(G902), .A2(G217), .ZN(n1308) );
XNOR2_X1 U1048 ( .A(n1319), .B(n1070), .ZN(n1231) );
NAND2_X1 U1049 ( .A1(n1320), .A2(n1153), .ZN(n1070) );
INV_X1 U1050 ( .A(G902), .ZN(n1153) );
XOR2_X1 U1051 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1052 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR2_X1 U1053 ( .A1(KEYINPUT46), .A2(n1138), .ZN(n1324) );
NAND3_X1 U1054 ( .A1(n1255), .A2(n1040), .A3(G210), .ZN(n1138) );
INV_X1 U1055 ( .A(G953), .ZN(n1040) );
INV_X1 U1056 ( .A(G237), .ZN(n1255) );
NAND2_X1 U1057 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
NAND2_X1 U1058 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
XOR2_X1 U1059 ( .A(n1329), .B(KEYINPUT2), .Z(n1325) );
NAND2_X1 U1060 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XOR2_X1 U1061 ( .A(KEYINPUT5), .B(n1328), .Z(n1331) );
XNOR2_X1 U1062 ( .A(n1281), .B(KEYINPUT1), .ZN(n1328) );
XNOR2_X1 U1063 ( .A(n1142), .B(n1098), .ZN(n1281) );
XNOR2_X1 U1064 ( .A(n1259), .B(n1134), .ZN(n1098) );
XNOR2_X1 U1065 ( .A(G131), .B(G134), .ZN(n1134) );
XOR2_X1 U1066 ( .A(G146), .B(n1299), .Z(n1259) );
XOR2_X1 U1067 ( .A(G128), .B(G143), .Z(n1299) );
NOR2_X1 U1068 ( .A1(KEYINPUT27), .A2(n1097), .ZN(n1142) );
INV_X1 U1069 ( .A(G137), .ZN(n1097) );
INV_X1 U1070 ( .A(n1327), .ZN(n1330) );
XOR2_X1 U1071 ( .A(n1131), .B(KEYINPUT62), .Z(n1327) );
XOR2_X1 U1072 ( .A(G113), .B(n1332), .Z(n1131) );
XNOR2_X1 U1073 ( .A(n1267), .B(G116), .ZN(n1332) );
INV_X1 U1074 ( .A(G119), .ZN(n1267) );
XNOR2_X1 U1075 ( .A(G101), .B(KEYINPUT60), .ZN(n1321) );
NAND2_X1 U1076 ( .A1(KEYINPUT48), .A2(n1333), .ZN(n1319) );
INV_X1 U1077 ( .A(G472), .ZN(n1333) );
endmodule


