//Key = 0111111000100001111110111011010111101110010111001101110110110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271;

XNOR2_X1 U706 ( .A(G107), .B(n985), .ZN(G9) );
NOR2_X1 U707 ( .A1(n986), .A2(n987), .ZN(G75) );
NOR3_X1 U708 ( .A1(n988), .A2(n989), .A3(n990), .ZN(n987) );
NAND3_X1 U709 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n988) );
NAND2_X1 U710 ( .A1(n994), .A2(n995), .ZN(n991) );
NAND2_X1 U711 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND4_X1 U712 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(n997) );
NAND3_X1 U713 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n1000) );
NAND2_X1 U714 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U715 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND2_X1 U716 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
INV_X1 U717 ( .A(n1011), .ZN(n1007) );
NAND2_X1 U718 ( .A1(n1012), .A2(n1013), .ZN(n1003) );
NAND2_X1 U719 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U720 ( .A1(KEYINPUT2), .A2(n1016), .ZN(n1015) );
OR3_X1 U721 ( .A1(n1017), .A2(KEYINPUT2), .A3(n1012), .ZN(n1002) );
NAND3_X1 U722 ( .A1(n1012), .A2(n1018), .A3(n1005), .ZN(n996) );
NAND2_X1 U723 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND3_X1 U724 ( .A1(n1021), .A2(n1022), .A3(n998), .ZN(n1020) );
OR3_X1 U725 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NAND2_X1 U726 ( .A1(n1026), .A2(n1025), .ZN(n1021) );
XOR2_X1 U727 ( .A(n999), .B(KEYINPUT4), .Z(n1026) );
NAND2_X1 U728 ( .A1(n1027), .A2(n999), .ZN(n1019) );
INV_X1 U729 ( .A(n1028), .ZN(n994) );
AND3_X1 U730 ( .A1(n1029), .A2(n992), .A3(n993), .ZN(n986) );
NAND4_X1 U731 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n992) );
NOR4_X1 U732 ( .A1(n1034), .A2(n1025), .A3(n1035), .A4(n1036), .ZN(n1033) );
XOR2_X1 U733 ( .A(n1037), .B(KEYINPUT56), .Z(n1035) );
AND2_X1 U734 ( .A1(n1012), .A2(n998), .ZN(n1032) );
XOR2_X1 U735 ( .A(n1038), .B(n1039), .Z(n1031) );
NOR2_X1 U736 ( .A1(KEYINPUT8), .A2(n1040), .ZN(n1039) );
XOR2_X1 U737 ( .A(n1041), .B(KEYINPUT40), .Z(n1030) );
NAND2_X1 U738 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
XOR2_X1 U739 ( .A(KEYINPUT35), .B(n1044), .Z(n1042) );
XNOR2_X1 U740 ( .A(n989), .B(KEYINPUT26), .ZN(n1029) );
INV_X1 U741 ( .A(G952), .ZN(n989) );
XOR2_X1 U742 ( .A(n1045), .B(n1046), .Z(G72) );
NOR2_X1 U743 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
AND2_X1 U744 ( .A1(G227), .A2(G900), .ZN(n1047) );
XOR2_X1 U745 ( .A(n1049), .B(n1050), .Z(n1045) );
NOR2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U747 ( .A(n1053), .B(n1054), .ZN(n1052) );
XNOR2_X1 U748 ( .A(KEYINPUT5), .B(n1055), .ZN(n1053) );
NOR2_X1 U749 ( .A1(KEYINPUT9), .A2(n1056), .ZN(n1055) );
XOR2_X1 U750 ( .A(n1057), .B(n1058), .Z(n1056) );
XOR2_X1 U751 ( .A(G131), .B(n1059), .Z(n1058) );
NOR2_X1 U752 ( .A1(KEYINPUT0), .A2(n1060), .ZN(n1059) );
NAND2_X1 U753 ( .A1(n1061), .A2(KEYINPUT38), .ZN(n1057) );
XOR2_X1 U754 ( .A(n1062), .B(KEYINPUT10), .Z(n1061) );
NOR2_X1 U755 ( .A1(G900), .A2(n1063), .ZN(n1051) );
NAND2_X1 U756 ( .A1(KEYINPUT1), .A2(n1064), .ZN(n1049) );
NAND2_X1 U757 ( .A1(n1065), .A2(n1048), .ZN(n1064) );
NAND3_X1 U758 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
XOR2_X1 U759 ( .A(n1069), .B(KEYINPUT30), .Z(n1068) );
XNOR2_X1 U760 ( .A(KEYINPUT55), .B(n1070), .ZN(n1067) );
XOR2_X1 U761 ( .A(n1071), .B(n1072), .Z(G69) );
NAND2_X1 U762 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U763 ( .A1(G898), .A2(G224), .ZN(n1074) );
XNOR2_X1 U764 ( .A(G953), .B(KEYINPUT17), .ZN(n1073) );
NAND2_X1 U765 ( .A1(KEYINPUT27), .A2(n1075), .ZN(n1071) );
XOR2_X1 U766 ( .A(n1076), .B(n1077), .Z(n1075) );
NAND2_X1 U767 ( .A1(n1048), .A2(n1078), .ZN(n1077) );
NAND3_X1 U768 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1076) );
INV_X1 U769 ( .A(n1082), .ZN(n1081) );
NAND2_X1 U770 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
NAND2_X1 U771 ( .A1(n1085), .A2(n1086), .ZN(n1079) );
XOR2_X1 U772 ( .A(n1084), .B(KEYINPUT59), .Z(n1086) );
NOR2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(G66) );
XNOR2_X1 U774 ( .A(n1089), .B(n1090), .ZN(n1088) );
XOR2_X1 U775 ( .A(KEYINPUT42), .B(n1091), .Z(n1090) );
NOR2_X1 U776 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U777 ( .A(G217), .B(KEYINPUT28), .ZN(n1092) );
NOR2_X1 U778 ( .A1(n1087), .A2(n1094), .ZN(G63) );
XOR2_X1 U779 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U780 ( .A1(n1097), .A2(n1093), .ZN(n1095) );
NOR2_X1 U781 ( .A1(n1087), .A2(n1098), .ZN(G60) );
XNOR2_X1 U782 ( .A(n1099), .B(n1100), .ZN(n1098) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1093), .ZN(n1100) );
XOR2_X1 U784 ( .A(n1102), .B(n1103), .Z(G6) );
NAND2_X1 U785 ( .A1(KEYINPUT48), .A2(G104), .ZN(n1103) );
NOR2_X1 U786 ( .A1(n1087), .A2(n1104), .ZN(G57) );
XNOR2_X1 U787 ( .A(n1105), .B(n1106), .ZN(n1104) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR3_X1 U789 ( .A1(n1093), .A2(KEYINPUT39), .A3(n1040), .ZN(n1107) );
NOR2_X1 U790 ( .A1(n1087), .A2(n1109), .ZN(G54) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(n1109) );
XNOR2_X1 U792 ( .A(n1112), .B(n1113), .ZN(n1111) );
XOR2_X1 U793 ( .A(n1114), .B(n1115), .Z(n1110) );
XOR2_X1 U794 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U795 ( .A1(n1118), .A2(n1093), .ZN(n1117) );
NAND2_X1 U796 ( .A1(KEYINPUT33), .A2(n1119), .ZN(n1116) );
NOR2_X1 U797 ( .A1(n1087), .A2(n1120), .ZN(G51) );
NOR2_X1 U798 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U799 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U800 ( .A1(n1125), .A2(n1093), .ZN(n1124) );
NAND2_X1 U801 ( .A1(G902), .A2(n990), .ZN(n1093) );
NAND4_X1 U802 ( .A1(n1126), .A2(n1066), .A3(n1070), .A4(n1069), .ZN(n990) );
AND4_X1 U803 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1066) );
NOR2_X1 U804 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U805 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
XNOR2_X1 U807 ( .A(n1016), .B(KEYINPUT43), .ZN(n1136) );
INV_X1 U808 ( .A(n1078), .ZN(n1126) );
NAND4_X1 U809 ( .A1(n1137), .A2(n1102), .A3(n1138), .A4(n1139), .ZN(n1078) );
AND4_X1 U810 ( .A1(n985), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1139) );
NAND3_X1 U811 ( .A1(n1016), .A2(n999), .A3(n1143), .ZN(n985) );
NOR2_X1 U812 ( .A1(n1144), .A2(n1145), .ZN(n1138) );
NOR2_X1 U813 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND3_X1 U814 ( .A1(n1143), .A2(n999), .A3(n1135), .ZN(n1102) );
OR2_X1 U815 ( .A1(n1148), .A2(n1149), .ZN(n1137) );
NOR2_X1 U816 ( .A1(KEYINPUT63), .A2(n1150), .ZN(n1123) );
XOR2_X1 U817 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U818 ( .A1(n1153), .A2(n1154), .ZN(n1121) );
INV_X1 U819 ( .A(KEYINPUT63), .ZN(n1154) );
XNOR2_X1 U820 ( .A(n1152), .B(n1151), .ZN(n1153) );
XNOR2_X1 U821 ( .A(n1155), .B(n1156), .ZN(n1152) );
NAND2_X1 U822 ( .A1(KEYINPUT51), .A2(n1157), .ZN(n1155) );
NOR2_X1 U823 ( .A1(n1048), .A2(G952), .ZN(n1087) );
XOR2_X1 U824 ( .A(G146), .B(n1158), .Z(G48) );
NOR2_X1 U825 ( .A1(n1014), .A2(n1134), .ZN(n1158) );
XNOR2_X1 U826 ( .A(n1131), .B(n1159), .ZN(G45) );
NOR2_X1 U827 ( .A1(G143), .A2(KEYINPUT25), .ZN(n1159) );
AND3_X1 U828 ( .A1(n1160), .A2(n1023), .A3(n1161), .ZN(n1131) );
AND3_X1 U829 ( .A1(n1162), .A2(n1036), .A3(n1011), .ZN(n1161) );
XNOR2_X1 U830 ( .A(G140), .B(n1129), .ZN(G42) );
NAND3_X1 U831 ( .A1(n1135), .A2(n1024), .A3(n1163), .ZN(n1129) );
XNOR2_X1 U832 ( .A(G137), .B(n1070), .ZN(G39) );
NAND2_X1 U833 ( .A1(n1163), .A2(n1164), .ZN(n1070) );
XNOR2_X1 U834 ( .A(G134), .B(n1127), .ZN(G36) );
NAND3_X1 U835 ( .A1(n1023), .A2(n1016), .A3(n1163), .ZN(n1127) );
XNOR2_X1 U836 ( .A(G131), .B(n1069), .ZN(G33) );
NAND3_X1 U837 ( .A1(n1023), .A2(n1135), .A3(n1163), .ZN(n1069) );
AND4_X1 U838 ( .A1(n998), .A2(n1011), .A3(n1165), .A4(n1001), .ZN(n1163) );
XNOR2_X1 U839 ( .A(n1166), .B(n1167), .ZN(G30) );
NOR2_X1 U840 ( .A1(n1017), .A2(n1134), .ZN(n1167) );
NAND4_X1 U841 ( .A1(n1168), .A2(n1160), .A3(n1011), .A4(n1169), .ZN(n1134) );
XNOR2_X1 U842 ( .A(n1170), .B(n1144), .ZN(G3) );
AND3_X1 U843 ( .A1(n1005), .A2(n1143), .A3(n1023), .ZN(n1144) );
XNOR2_X1 U844 ( .A(n1171), .B(n1128), .ZN(G27) );
NAND4_X1 U845 ( .A1(n1160), .A2(n1135), .A3(n1012), .A4(n1024), .ZN(n1128) );
AND2_X1 U846 ( .A1(n1027), .A2(n1165), .ZN(n1160) );
NAND2_X1 U847 ( .A1(n1172), .A2(n1173), .ZN(n1165) );
OR4_X1 U848 ( .A1(n1174), .A2(n1063), .A3(n1175), .A4(G900), .ZN(n1173) );
INV_X1 U849 ( .A(n1176), .ZN(n1175) );
XNOR2_X1 U850 ( .A(KEYINPUT29), .B(n1028), .ZN(n1172) );
NAND2_X1 U851 ( .A1(KEYINPUT36), .A2(n1177), .ZN(n1171) );
XOR2_X1 U852 ( .A(G122), .B(n1178), .Z(G24) );
NOR3_X1 U853 ( .A1(n1149), .A2(KEYINPUT47), .A3(n1179), .ZN(n1178) );
XOR2_X1 U854 ( .A(n1148), .B(KEYINPUT11), .Z(n1179) );
NAND4_X1 U855 ( .A1(n1162), .A2(n1180), .A3(n999), .A4(n1036), .ZN(n1148) );
NAND2_X1 U856 ( .A1(n1181), .A2(n1182), .ZN(n999) );
OR3_X1 U857 ( .A1(n1169), .A2(n1168), .A3(KEYINPUT14), .ZN(n1182) );
NAND2_X1 U858 ( .A1(KEYINPUT14), .A2(n1024), .ZN(n1181) );
XNOR2_X1 U859 ( .A(n1183), .B(n1184), .ZN(G21) );
NOR2_X1 U860 ( .A1(n1185), .A2(n1147), .ZN(n1184) );
NAND3_X1 U861 ( .A1(n1027), .A2(n1186), .A3(n1164), .ZN(n1147) );
AND3_X1 U862 ( .A1(n1005), .A2(n1169), .A3(n1168), .ZN(n1164) );
INV_X1 U863 ( .A(n1187), .ZN(n1169) );
XNOR2_X1 U864 ( .A(n1012), .B(KEYINPUT54), .ZN(n1185) );
XNOR2_X1 U865 ( .A(G116), .B(n1142), .ZN(G18) );
NAND4_X1 U866 ( .A1(n1027), .A2(n1023), .A3(n1180), .A4(n1016), .ZN(n1142) );
INV_X1 U867 ( .A(n1017), .ZN(n1016) );
NAND2_X1 U868 ( .A1(n1188), .A2(n1036), .ZN(n1017) );
XOR2_X1 U869 ( .A(n1162), .B(KEYINPUT34), .Z(n1188) );
INV_X1 U870 ( .A(n1149), .ZN(n1027) );
XOR2_X1 U871 ( .A(n1189), .B(KEYINPUT41), .Z(n1149) );
XNOR2_X1 U872 ( .A(G113), .B(n1141), .ZN(G15) );
NAND4_X1 U873 ( .A1(n1023), .A2(n1135), .A3(n1180), .A4(n1189), .ZN(n1141) );
AND2_X1 U874 ( .A1(n1012), .A2(n1186), .ZN(n1180) );
INV_X1 U875 ( .A(n1146), .ZN(n1012) );
NAND2_X1 U876 ( .A1(n1010), .A2(n1190), .ZN(n1146) );
INV_X1 U877 ( .A(n1014), .ZN(n1135) );
NAND2_X1 U878 ( .A1(n1191), .A2(n1162), .ZN(n1014) );
INV_X1 U879 ( .A(n1036), .ZN(n1191) );
AND2_X1 U880 ( .A1(n1168), .A2(n1187), .ZN(n1023) );
XNOR2_X1 U881 ( .A(G110), .B(n1140), .ZN(G12) );
NAND3_X1 U882 ( .A1(n1143), .A2(n1024), .A3(n1005), .ZN(n1140) );
NOR2_X1 U883 ( .A1(n1036), .A2(n1162), .ZN(n1005) );
XOR2_X1 U884 ( .A(n1037), .B(KEYINPUT3), .Z(n1162) );
XOR2_X1 U885 ( .A(n1192), .B(n1193), .Z(n1037) );
XNOR2_X1 U886 ( .A(KEYINPUT7), .B(n1101), .ZN(n1193) );
INV_X1 U887 ( .A(G475), .ZN(n1101) );
NAND2_X1 U888 ( .A1(n1099), .A2(n1174), .ZN(n1192) );
XNOR2_X1 U889 ( .A(n1194), .B(n1195), .ZN(n1099) );
XOR2_X1 U890 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U891 ( .A(G131), .B(G104), .Z(n1197) );
XOR2_X1 U892 ( .A(KEYINPUT58), .B(G143), .Z(n1196) );
XOR2_X1 U893 ( .A(n1198), .B(n1199), .Z(n1194) );
XOR2_X1 U894 ( .A(n1200), .B(n1054), .Z(n1199) );
NAND2_X1 U895 ( .A1(n1201), .A2(G214), .ZN(n1200) );
XNOR2_X1 U896 ( .A(n1202), .B(n1203), .ZN(n1198) );
NAND2_X1 U897 ( .A1(KEYINPUT32), .A2(n1204), .ZN(n1203) );
NAND2_X1 U898 ( .A1(KEYINPUT15), .A2(n1205), .ZN(n1202) );
XOR2_X1 U899 ( .A(G122), .B(G113), .Z(n1205) );
XOR2_X1 U900 ( .A(n1206), .B(n1097), .Z(n1036) );
INV_X1 U901 ( .A(G478), .ZN(n1097) );
OR2_X1 U902 ( .A1(n1096), .A2(G902), .ZN(n1206) );
XNOR2_X1 U903 ( .A(n1207), .B(n1208), .ZN(n1096) );
XOR2_X1 U904 ( .A(n1209), .B(n1210), .Z(n1208) );
XNOR2_X1 U905 ( .A(n1166), .B(G122), .ZN(n1210) );
XOR2_X1 U906 ( .A(G143), .B(G134), .Z(n1209) );
XOR2_X1 U907 ( .A(n1211), .B(n1212), .Z(n1207) );
XNOR2_X1 U908 ( .A(G116), .B(n1213), .ZN(n1212) );
NAND3_X1 U909 ( .A1(G234), .A2(n1048), .A3(G217), .ZN(n1213) );
NAND2_X1 U910 ( .A1(KEYINPUT44), .A2(n1214), .ZN(n1211) );
NOR2_X1 U911 ( .A1(n1168), .A2(n1187), .ZN(n1024) );
NOR2_X1 U912 ( .A1(n1215), .A2(n1034), .ZN(n1187) );
NOR2_X1 U913 ( .A1(n1043), .A2(n1044), .ZN(n1034) );
AND2_X1 U914 ( .A1(n1044), .A2(n1043), .ZN(n1215) );
NAND2_X1 U915 ( .A1(n1089), .A2(n1174), .ZN(n1043) );
NAND2_X1 U916 ( .A1(n1216), .A2(n1217), .ZN(n1089) );
NAND2_X1 U917 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U918 ( .A(KEYINPUT31), .B(n1220), .Z(n1216) );
NOR2_X1 U919 ( .A1(n1218), .A2(n1219), .ZN(n1220) );
NAND2_X1 U920 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
NAND2_X1 U921 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U922 ( .A(KEYINPUT53), .B(n1225), .Z(n1221) );
NOR2_X1 U923 ( .A1(n1224), .A2(n1223), .ZN(n1225) );
NAND3_X1 U924 ( .A1(G234), .A2(n1048), .A3(G221), .ZN(n1223) );
INV_X1 U925 ( .A(G137), .ZN(n1224) );
XNOR2_X1 U926 ( .A(n1226), .B(n1227), .ZN(n1218) );
XNOR2_X1 U927 ( .A(n1228), .B(n1229), .ZN(n1227) );
XNOR2_X1 U928 ( .A(n1230), .B(n1231), .ZN(n1229) );
NOR2_X1 U929 ( .A1(KEYINPUT57), .A2(n1183), .ZN(n1231) );
NOR2_X1 U930 ( .A1(KEYINPUT12), .A2(n1054), .ZN(n1230) );
XNOR2_X1 U931 ( .A(G125), .B(G140), .ZN(n1054) );
XNOR2_X1 U932 ( .A(G110), .B(n1232), .ZN(n1226) );
XNOR2_X1 U933 ( .A(KEYINPUT60), .B(n1166), .ZN(n1232) );
AND2_X1 U934 ( .A1(G217), .A2(n1233), .ZN(n1044) );
XNOR2_X1 U935 ( .A(n1234), .B(n1038), .ZN(n1168) );
NAND2_X1 U936 ( .A1(n1235), .A2(n1174), .ZN(n1038) );
XOR2_X1 U937 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U938 ( .A(KEYINPUT62), .B(KEYINPUT16), .Z(n1237) );
XNOR2_X1 U939 ( .A(n1108), .B(n1105), .ZN(n1236) );
XOR2_X1 U940 ( .A(n1238), .B(n1170), .Z(n1105) );
INV_X1 U941 ( .A(G101), .ZN(n1170) );
NAND2_X1 U942 ( .A1(n1201), .A2(G210), .ZN(n1238) );
NOR2_X1 U943 ( .A1(G953), .A2(G237), .ZN(n1201) );
XNOR2_X1 U944 ( .A(n1239), .B(n1240), .ZN(n1108) );
XNOR2_X1 U945 ( .A(n1119), .B(n1241), .ZN(n1240) );
XOR2_X1 U946 ( .A(n1242), .B(KEYINPUT45), .Z(n1241) );
NAND2_X1 U947 ( .A1(KEYINPUT37), .A2(n1183), .ZN(n1242) );
XOR2_X1 U948 ( .A(n1243), .B(n1244), .Z(n1239) );
NAND2_X1 U949 ( .A1(KEYINPUT24), .A2(n1040), .ZN(n1234) );
INV_X1 U950 ( .A(G472), .ZN(n1040) );
AND3_X1 U951 ( .A1(n1189), .A2(n1186), .A3(n1011), .ZN(n1143) );
NOR2_X1 U952 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
INV_X1 U953 ( .A(n1190), .ZN(n1009) );
NAND2_X1 U954 ( .A1(G221), .A2(n1233), .ZN(n1190) );
NAND2_X1 U955 ( .A1(G234), .A2(n1174), .ZN(n1233) );
XNOR2_X1 U956 ( .A(n1245), .B(n1118), .ZN(n1010) );
INV_X1 U957 ( .A(G469), .ZN(n1118) );
NAND2_X1 U958 ( .A1(n1246), .A2(n1174), .ZN(n1245) );
XOR2_X1 U959 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U960 ( .A(n1249), .B(n1119), .Z(n1248) );
XNOR2_X1 U961 ( .A(n1250), .B(G131), .ZN(n1119) );
NAND2_X1 U962 ( .A1(KEYINPUT19), .A2(n1062), .ZN(n1250) );
XNOR2_X1 U963 ( .A(G134), .B(G137), .ZN(n1062) );
NOR2_X1 U964 ( .A1(KEYINPUT13), .A2(n1114), .ZN(n1249) );
XNOR2_X1 U965 ( .A(n1085), .B(KEYINPUT18), .ZN(n1114) );
XNOR2_X1 U966 ( .A(n1112), .B(n1251), .ZN(n1247) );
INV_X1 U967 ( .A(n1113), .ZN(n1251) );
XNOR2_X1 U968 ( .A(n1252), .B(n1253), .ZN(n1113) );
XNOR2_X1 U969 ( .A(G140), .B(n1254), .ZN(n1253) );
NAND2_X1 U970 ( .A1(G227), .A2(n1048), .ZN(n1252) );
XOR2_X1 U971 ( .A(n1060), .B(KEYINPUT61), .Z(n1112) );
XNOR2_X1 U972 ( .A(n1255), .B(G128), .ZN(n1060) );
NAND2_X1 U973 ( .A1(n1028), .A2(n1256), .ZN(n1186) );
NAND3_X1 U974 ( .A1(n1082), .A2(n1176), .A3(G902), .ZN(n1256) );
NOR2_X1 U975 ( .A1(n1063), .A2(G898), .ZN(n1082) );
XNOR2_X1 U976 ( .A(G953), .B(KEYINPUT21), .ZN(n1063) );
NAND3_X1 U977 ( .A1(n993), .A2(n1176), .A3(G952), .ZN(n1028) );
NAND2_X1 U978 ( .A1(n1257), .A2(G237), .ZN(n1176) );
XNOR2_X1 U979 ( .A(G234), .B(KEYINPUT20), .ZN(n1257) );
XOR2_X1 U980 ( .A(G953), .B(KEYINPUT22), .Z(n993) );
NOR2_X1 U981 ( .A1(n998), .A2(n1025), .ZN(n1189) );
INV_X1 U982 ( .A(n1001), .ZN(n1025) );
NAND2_X1 U983 ( .A1(G214), .A2(n1258), .ZN(n1001) );
XNOR2_X1 U984 ( .A(n1259), .B(n1125), .ZN(n998) );
NAND2_X1 U985 ( .A1(G210), .A2(n1258), .ZN(n1125) );
NAND2_X1 U986 ( .A1(n1260), .A2(n1174), .ZN(n1258) );
INV_X1 U987 ( .A(G237), .ZN(n1260) );
NAND3_X1 U988 ( .A1(n1261), .A2(n1174), .A3(n1262), .ZN(n1259) );
XOR2_X1 U989 ( .A(n1263), .B(KEYINPUT46), .Z(n1262) );
OR2_X1 U990 ( .A1(n1264), .A2(n1151), .ZN(n1263) );
INV_X1 U991 ( .A(G902), .ZN(n1174) );
NAND2_X1 U992 ( .A1(n1151), .A2(n1264), .ZN(n1261) );
XOR2_X1 U993 ( .A(n1156), .B(n1265), .Z(n1264) );
XOR2_X1 U994 ( .A(KEYINPUT49), .B(n1157), .Z(n1265) );
XNOR2_X1 U995 ( .A(n1177), .B(KEYINPUT23), .ZN(n1157) );
INV_X1 U996 ( .A(G125), .ZN(n1177) );
XNOR2_X1 U997 ( .A(n1243), .B(n1266), .ZN(n1156) );
AND2_X1 U998 ( .A1(n1048), .A2(G224), .ZN(n1266) );
INV_X1 U999 ( .A(G953), .ZN(n1048) );
XOR2_X1 U1000 ( .A(n1267), .B(n1255), .Z(n1243) );
XNOR2_X1 U1001 ( .A(G143), .B(n1204), .ZN(n1255) );
INV_X1 U1002 ( .A(n1228), .ZN(n1204) );
XOR2_X1 U1003 ( .A(G146), .B(KEYINPUT50), .Z(n1228) );
NAND2_X1 U1004 ( .A1(KEYINPUT52), .A2(n1166), .ZN(n1267) );
INV_X1 U1005 ( .A(G128), .ZN(n1166) );
XOR2_X1 U1006 ( .A(n1084), .B(n1083), .Z(n1151) );
INV_X1 U1007 ( .A(n1085), .ZN(n1083) );
XOR2_X1 U1008 ( .A(G101), .B(n1268), .Z(n1085) );
XNOR2_X1 U1009 ( .A(n1214), .B(G104), .ZN(n1268) );
INV_X1 U1010 ( .A(G107), .ZN(n1214) );
XOR2_X1 U1011 ( .A(n1269), .B(n1270), .Z(n1084) );
XNOR2_X1 U1012 ( .A(G122), .B(n1183), .ZN(n1270) );
INV_X1 U1013 ( .A(G119), .ZN(n1183) );
XOR2_X1 U1014 ( .A(n1271), .B(n1244), .Z(n1269) );
XOR2_X1 U1015 ( .A(G113), .B(G116), .Z(n1244) );
NAND2_X1 U1016 ( .A1(KEYINPUT6), .A2(n1254), .ZN(n1271) );
INV_X1 U1017 ( .A(G110), .ZN(n1254) );
endmodule


