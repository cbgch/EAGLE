//Key = 0011100100111101001110110100101101100010011010111110010000100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410;

XNOR2_X1 U776 ( .A(n1080), .B(n1081), .ZN(G9) );
NOR2_X1 U777 ( .A1(n1082), .A2(n1083), .ZN(G75) );
NOR4_X1 U778 ( .A1(n1084), .A2(n1085), .A3(G953), .A4(n1086), .ZN(n1083) );
NOR3_X1 U779 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
NOR2_X1 U780 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U781 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR3_X1 U782 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1090) );
NOR4_X1 U783 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
NOR2_X1 U784 ( .A1(n1093), .A2(n1101), .ZN(n1100) );
INV_X1 U785 ( .A(KEYINPUT57), .ZN(n1101) );
NOR3_X1 U786 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1099) );
NOR2_X1 U787 ( .A1(n1105), .A2(n1106), .ZN(n1098) );
NOR2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(n1095) );
NOR2_X1 U789 ( .A1(KEYINPUT57), .A2(n1093), .ZN(n1107) );
NAND2_X1 U790 ( .A1(n1109), .A2(n1110), .ZN(n1093) );
NAND2_X1 U791 ( .A1(n1111), .A2(n1112), .ZN(n1084) );
NAND3_X1 U792 ( .A1(n1113), .A2(n1108), .A3(n1114), .ZN(n1112) );
INV_X1 U793 ( .A(n1094), .ZN(n1114) );
NAND2_X1 U794 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NAND2_X1 U795 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U796 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND3_X1 U797 ( .A1(n1110), .A2(n1121), .A3(n1122), .ZN(n1120) );
NAND2_X1 U798 ( .A1(n1109), .A2(n1123), .ZN(n1119) );
NAND2_X1 U799 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND3_X1 U800 ( .A1(n1121), .A2(n1126), .A3(KEYINPUT58), .ZN(n1125) );
NAND2_X1 U801 ( .A1(n1110), .A2(n1127), .ZN(n1124) );
OR2_X1 U802 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(n1115) );
INV_X1 U804 ( .A(KEYINPUT58), .ZN(n1131) );
NAND4_X1 U805 ( .A1(n1117), .A2(n1109), .A3(n1121), .A4(n1126), .ZN(n1130) );
INV_X1 U806 ( .A(n1087), .ZN(n1117) );
NOR3_X1 U807 ( .A1(n1086), .A2(G953), .A3(G952), .ZN(n1082) );
AND4_X1 U808 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1086) );
NOR4_X1 U809 ( .A1(n1136), .A2(n1137), .A3(n1106), .A4(n1138), .ZN(n1135) );
XNOR2_X1 U810 ( .A(n1139), .B(n1140), .ZN(n1138) );
XOR2_X1 U811 ( .A(n1141), .B(KEYINPUT48), .Z(n1136) );
NAND2_X1 U812 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR3_X1 U813 ( .A1(n1144), .A2(n1145), .A3(n1097), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1143), .A2(n1142), .ZN(n1144) );
XNOR2_X1 U815 ( .A(G472), .B(KEYINPUT52), .ZN(n1142) );
NAND2_X1 U816 ( .A1(n1146), .A2(n1147), .ZN(n1133) );
XNOR2_X1 U817 ( .A(n1148), .B(n1149), .ZN(n1132) );
NAND2_X1 U818 ( .A1(KEYINPUT18), .A2(n1150), .ZN(n1149) );
XOR2_X1 U819 ( .A(n1151), .B(n1152), .Z(G72) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
INV_X1 U822 ( .A(n1157), .ZN(n1155) );
NOR3_X1 U823 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1153) );
XNOR2_X1 U824 ( .A(KEYINPUT59), .B(n1156), .ZN(n1159) );
NAND2_X1 U825 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
NAND2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U827 ( .A(n1164), .B(KEYINPUT47), .ZN(n1162) );
NOR2_X1 U828 ( .A1(G900), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U829 ( .A(n1165), .B(n1166), .ZN(n1157) );
XNOR2_X1 U830 ( .A(n1167), .B(n1168), .ZN(n1166) );
NOR2_X1 U831 ( .A1(G134), .A2(KEYINPUT61), .ZN(n1168) );
NAND2_X1 U832 ( .A1(KEYINPUT4), .A2(n1169), .ZN(n1167) );
XOR2_X1 U833 ( .A(n1170), .B(n1171), .Z(n1165) );
NAND3_X1 U834 ( .A1(G953), .A2(n1172), .A3(KEYINPUT13), .ZN(n1151) );
NAND2_X1 U835 ( .A1(G900), .A2(G227), .ZN(n1172) );
NAND2_X1 U836 ( .A1(n1173), .A2(n1174), .ZN(G69) );
NAND2_X1 U837 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND2_X1 U838 ( .A1(KEYINPUT3), .A2(n1177), .ZN(n1176) );
NAND2_X1 U839 ( .A1(G953), .A2(n1178), .ZN(n1177) );
NAND2_X1 U840 ( .A1(G898), .A2(G224), .ZN(n1178) );
INV_X1 U841 ( .A(n1179), .ZN(n1175) );
NAND3_X1 U842 ( .A1(KEYINPUT3), .A2(n1180), .A3(n1179), .ZN(n1173) );
XNOR2_X1 U843 ( .A(n1181), .B(n1182), .ZN(n1179) );
NOR2_X1 U844 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U845 ( .A(n1185), .B(n1186), .Z(n1184) );
XNOR2_X1 U846 ( .A(n1187), .B(n1188), .ZN(n1186) );
NOR2_X1 U847 ( .A1(KEYINPUT14), .A2(n1189), .ZN(n1188) );
XNOR2_X1 U848 ( .A(G122), .B(G110), .ZN(n1189) );
NOR2_X1 U849 ( .A1(KEYINPUT17), .A2(n1190), .ZN(n1187) );
XOR2_X1 U850 ( .A(n1191), .B(n1192), .Z(n1190) );
XNOR2_X1 U851 ( .A(KEYINPUT10), .B(n1193), .ZN(n1192) );
NOR2_X1 U852 ( .A1(G898), .A2(n1160), .ZN(n1183) );
NAND2_X1 U853 ( .A1(n1160), .A2(n1194), .ZN(n1181) );
NAND2_X1 U854 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
OR2_X1 U855 ( .A1(n1160), .A2(G224), .ZN(n1180) );
NOR2_X1 U856 ( .A1(n1197), .A2(n1198), .ZN(G66) );
XOR2_X1 U857 ( .A(n1199), .B(n1200), .Z(n1198) );
NAND2_X1 U858 ( .A1(n1201), .A2(n1202), .ZN(n1199) );
NOR2_X1 U859 ( .A1(n1203), .A2(n1204), .ZN(G63) );
XOR2_X1 U860 ( .A(n1205), .B(n1206), .Z(n1204) );
NAND2_X1 U861 ( .A1(n1201), .A2(G478), .ZN(n1205) );
NOR2_X1 U862 ( .A1(n1160), .A2(n1207), .ZN(n1203) );
XOR2_X1 U863 ( .A(KEYINPUT21), .B(G952), .Z(n1207) );
NOR2_X1 U864 ( .A1(n1197), .A2(n1208), .ZN(G60) );
NOR3_X1 U865 ( .A1(n1148), .A2(n1209), .A3(n1210), .ZN(n1208) );
AND3_X1 U866 ( .A1(n1211), .A2(G475), .A3(n1201), .ZN(n1210) );
NOR2_X1 U867 ( .A1(n1212), .A2(n1211), .ZN(n1209) );
NOR2_X1 U868 ( .A1(n1111), .A2(n1150), .ZN(n1212) );
INV_X1 U869 ( .A(G475), .ZN(n1150) );
XNOR2_X1 U870 ( .A(G104), .B(n1196), .ZN(G6) );
NOR2_X1 U871 ( .A1(n1197), .A2(n1213), .ZN(G57) );
XNOR2_X1 U872 ( .A(n1214), .B(n1215), .ZN(n1213) );
NAND3_X1 U873 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1214) );
OR2_X1 U874 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND3_X1 U875 ( .A1(n1220), .A2(n1219), .A3(KEYINPUT63), .ZN(n1217) );
AND2_X1 U876 ( .A1(KEYINPUT12), .A2(n1221), .ZN(n1220) );
OR2_X1 U877 ( .A1(n1221), .A2(KEYINPUT63), .ZN(n1216) );
AND2_X1 U878 ( .A1(n1201), .A2(G472), .ZN(n1221) );
NOR2_X1 U879 ( .A1(n1197), .A2(n1222), .ZN(G54) );
XOR2_X1 U880 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U881 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U882 ( .A(n1227), .B(n1228), .ZN(n1226) );
XNOR2_X1 U883 ( .A(G140), .B(n1229), .ZN(n1225) );
XNOR2_X1 U884 ( .A(n1230), .B(n1169), .ZN(n1223) );
XOR2_X1 U885 ( .A(n1231), .B(n1232), .Z(n1230) );
NAND2_X1 U886 ( .A1(n1201), .A2(G469), .ZN(n1231) );
NOR2_X1 U887 ( .A1(n1197), .A2(n1233), .ZN(G51) );
XOR2_X1 U888 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U889 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND2_X1 U890 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U891 ( .A1(n1201), .A2(n1139), .ZN(n1236) );
NOR2_X1 U892 ( .A1(n1240), .A2(n1111), .ZN(n1201) );
AND4_X1 U893 ( .A1(n1241), .A2(n1163), .A3(n1164), .A4(n1195), .ZN(n1111) );
AND4_X1 U894 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1195) );
NOR3_X1 U895 ( .A1(n1081), .A2(n1246), .A3(n1247), .ZN(n1245) );
AND3_X1 U896 ( .A1(n1248), .A2(n1249), .A3(n1121), .ZN(n1081) );
NAND2_X1 U897 ( .A1(n1250), .A2(n1251), .ZN(n1244) );
NAND3_X1 U898 ( .A1(n1252), .A2(n1253), .A3(n1254), .ZN(n1251) );
NAND2_X1 U899 ( .A1(KEYINPUT42), .A2(n1255), .ZN(n1254) );
NAND3_X1 U900 ( .A1(n1129), .A2(n1249), .A3(n1256), .ZN(n1253) );
XNOR2_X1 U901 ( .A(n1092), .B(KEYINPUT40), .ZN(n1256) );
NAND3_X1 U902 ( .A1(n1257), .A2(n1122), .A3(n1258), .ZN(n1252) );
XNOR2_X1 U903 ( .A(n1129), .B(KEYINPUT49), .ZN(n1258) );
NAND4_X1 U904 ( .A1(n1255), .A2(n1259), .A3(n1110), .A4(n1260), .ZN(n1243) );
INV_X1 U905 ( .A(KEYINPUT42), .ZN(n1260) );
INV_X1 U906 ( .A(n1106), .ZN(n1110) );
NAND3_X1 U907 ( .A1(n1128), .A2(n1248), .A3(n1109), .ZN(n1242) );
AND4_X1 U908 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1164) );
AND4_X1 U909 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1163) );
XOR2_X1 U910 ( .A(n1196), .B(KEYINPUT5), .Z(n1241) );
NAND3_X1 U911 ( .A1(n1121), .A2(n1248), .A3(n1122), .ZN(n1196) );
NOR2_X1 U912 ( .A1(n1160), .A2(G952), .ZN(n1197) );
XOR2_X1 U913 ( .A(n1269), .B(n1270), .Z(G48) );
NOR2_X1 U914 ( .A1(KEYINPUT29), .A2(n1271), .ZN(n1270) );
NAND2_X1 U915 ( .A1(n1272), .A2(n1273), .ZN(n1269) );
NAND3_X1 U916 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
NAND2_X1 U917 ( .A1(n1122), .A2(n1277), .ZN(n1275) );
OR2_X1 U918 ( .A1(n1264), .A2(n1276), .ZN(n1272) );
INV_X1 U919 ( .A(KEYINPUT46), .ZN(n1276) );
NAND3_X1 U920 ( .A1(n1274), .A2(n1277), .A3(n1122), .ZN(n1264) );
XNOR2_X1 U921 ( .A(G143), .B(n1261), .ZN(G45) );
NAND4_X1 U922 ( .A1(n1274), .A2(n1126), .A3(n1129), .A4(n1278), .ZN(n1261) );
NOR3_X1 U923 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1278) );
XNOR2_X1 U924 ( .A(G140), .B(n1262), .ZN(G42) );
NAND3_X1 U925 ( .A1(n1122), .A2(n1282), .A3(n1128), .ZN(n1262) );
XNOR2_X1 U926 ( .A(G137), .B(n1263), .ZN(G39) );
NAND4_X1 U927 ( .A1(n1109), .A2(n1282), .A3(n1137), .A4(n1283), .ZN(n1263) );
XNOR2_X1 U928 ( .A(G134), .B(n1265), .ZN(G36) );
NAND3_X1 U929 ( .A1(n1282), .A2(n1249), .A3(n1129), .ZN(n1265) );
XOR2_X1 U930 ( .A(n1267), .B(n1284), .Z(G33) );
NAND2_X1 U931 ( .A1(KEYINPUT53), .A2(G131), .ZN(n1284) );
NAND3_X1 U932 ( .A1(n1122), .A2(n1282), .A3(n1129), .ZN(n1267) );
NOR4_X1 U933 ( .A1(n1094), .A2(n1285), .A3(n1280), .A4(n1097), .ZN(n1282) );
INV_X1 U934 ( .A(n1108), .ZN(n1097) );
XOR2_X1 U935 ( .A(n1268), .B(n1286), .Z(G30) );
XOR2_X1 U936 ( .A(KEYINPUT44), .B(G128), .Z(n1286) );
NAND3_X1 U937 ( .A1(n1274), .A2(n1249), .A3(n1277), .ZN(n1268) );
AND4_X1 U938 ( .A1(n1126), .A2(n1137), .A3(n1283), .A4(n1287), .ZN(n1277) );
XOR2_X1 U939 ( .A(G101), .B(n1247), .Z(G3) );
AND3_X1 U940 ( .A1(n1129), .A2(n1248), .A3(n1109), .ZN(n1247) );
AND3_X1 U941 ( .A1(n1257), .A2(n1288), .A3(n1126), .ZN(n1248) );
INV_X1 U942 ( .A(n1285), .ZN(n1126) );
NAND2_X1 U943 ( .A1(n1289), .A2(n1290), .ZN(G27) );
OR2_X1 U944 ( .A1(n1266), .A2(G125), .ZN(n1290) );
XOR2_X1 U945 ( .A(n1291), .B(KEYINPUT56), .Z(n1289) );
NAND2_X1 U946 ( .A1(G125), .A2(n1266), .ZN(n1291) );
NAND4_X1 U947 ( .A1(n1128), .A2(n1122), .A3(n1292), .A4(n1274), .ZN(n1266) );
NOR2_X1 U948 ( .A1(n1280), .A2(n1106), .ZN(n1292) );
INV_X1 U949 ( .A(n1287), .ZN(n1280) );
NAND2_X1 U950 ( .A1(n1087), .A2(n1293), .ZN(n1287) );
NAND4_X1 U951 ( .A1(G953), .A2(G902), .A3(n1294), .A4(n1295), .ZN(n1293) );
INV_X1 U952 ( .A(G900), .ZN(n1295) );
INV_X1 U953 ( .A(n1296), .ZN(n1128) );
XOR2_X1 U954 ( .A(G122), .B(n1246), .Z(G24) );
AND3_X1 U955 ( .A1(n1274), .A2(n1250), .A3(n1297), .ZN(n1246) );
NOR3_X1 U956 ( .A1(n1089), .A2(n1281), .A3(n1279), .ZN(n1297) );
INV_X1 U957 ( .A(n1121), .ZN(n1089) );
NOR2_X1 U958 ( .A1(n1283), .A2(n1137), .ZN(n1121) );
XOR2_X1 U959 ( .A(n1298), .B(G119), .Z(G21) );
NAND2_X1 U960 ( .A1(KEYINPUT15), .A2(n1299), .ZN(n1298) );
NAND2_X1 U961 ( .A1(n1255), .A2(n1250), .ZN(n1299) );
AND4_X1 U962 ( .A1(n1274), .A2(n1109), .A3(n1137), .A4(n1283), .ZN(n1255) );
INV_X1 U963 ( .A(n1300), .ZN(n1283) );
INV_X1 U964 ( .A(n1092), .ZN(n1274) );
XNOR2_X1 U965 ( .A(G116), .B(n1301), .ZN(G18) );
NOR2_X1 U966 ( .A1(KEYINPUT0), .A2(n1302), .ZN(n1301) );
NOR3_X1 U967 ( .A1(n1303), .A2(n1105), .A3(n1092), .ZN(n1302) );
XNOR2_X1 U968 ( .A(n1304), .B(KEYINPUT28), .ZN(n1092) );
INV_X1 U969 ( .A(n1249), .ZN(n1105) );
NOR2_X1 U970 ( .A1(n1305), .A2(n1281), .ZN(n1249) );
XOR2_X1 U971 ( .A(n1306), .B(KEYINPUT30), .Z(n1281) );
XOR2_X1 U972 ( .A(KEYINPUT38), .B(n1279), .Z(n1305) );
XNOR2_X1 U973 ( .A(G113), .B(n1307), .ZN(G15) );
NAND4_X1 U974 ( .A1(KEYINPUT41), .A2(n1308), .A3(n1257), .A4(n1122), .ZN(n1307) );
NOR2_X1 U975 ( .A1(n1306), .A2(n1279), .ZN(n1122) );
INV_X1 U976 ( .A(n1303), .ZN(n1308) );
NAND2_X1 U977 ( .A1(n1250), .A2(n1129), .ZN(n1303) );
NOR2_X1 U978 ( .A1(n1137), .A2(n1300), .ZN(n1129) );
NOR2_X1 U979 ( .A1(n1106), .A2(n1259), .ZN(n1250) );
NAND2_X1 U980 ( .A1(n1309), .A2(n1102), .ZN(n1106) );
INV_X1 U981 ( .A(n1104), .ZN(n1309) );
XNOR2_X1 U982 ( .A(G110), .B(n1310), .ZN(G12) );
NAND3_X1 U983 ( .A1(n1311), .A2(n1109), .A3(n1312), .ZN(n1310) );
NOR3_X1 U984 ( .A1(n1296), .A2(n1259), .A3(n1285), .ZN(n1312) );
NAND2_X1 U985 ( .A1(n1104), .A2(n1102), .ZN(n1285) );
NAND2_X1 U986 ( .A1(G221), .A2(n1313), .ZN(n1102) );
XNOR2_X1 U987 ( .A(n1314), .B(G469), .ZN(n1104) );
NAND2_X1 U988 ( .A1(n1315), .A2(n1240), .ZN(n1314) );
XOR2_X1 U989 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U990 ( .A(n1232), .B(n1169), .ZN(n1317) );
XNOR2_X1 U991 ( .A(G128), .B(n1318), .ZN(n1169) );
NOR2_X1 U992 ( .A1(KEYINPUT43), .A2(n1319), .ZN(n1318) );
XNOR2_X1 U993 ( .A(G146), .B(G143), .ZN(n1319) );
XOR2_X1 U994 ( .A(n1320), .B(n1321), .Z(n1316) );
XOR2_X1 U995 ( .A(n1228), .B(n1322), .Z(n1321) );
NOR2_X1 U996 ( .A1(KEYINPUT45), .A2(n1323), .ZN(n1322) );
XOR2_X1 U997 ( .A(n1324), .B(G140), .Z(n1323) );
NAND2_X1 U998 ( .A1(KEYINPUT34), .A2(G110), .ZN(n1324) );
NAND2_X1 U999 ( .A1(G227), .A2(n1160), .ZN(n1228) );
NAND2_X1 U1000 ( .A1(KEYINPUT11), .A2(n1227), .ZN(n1320) );
AND3_X1 U1001 ( .A1(n1325), .A2(n1326), .A3(n1327), .ZN(n1227) );
NAND2_X1 U1002 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
OR4_X1 U1003 ( .A1(n1328), .A2(KEYINPUT32), .A3(n1329), .A4(G101), .ZN(n1326) );
INV_X1 U1004 ( .A(KEYINPUT50), .ZN(n1329) );
NAND2_X1 U1005 ( .A1(G101), .A2(n1330), .ZN(n1325) );
OR2_X1 U1006 ( .A1(n1328), .A2(KEYINPUT32), .ZN(n1330) );
NAND3_X1 U1007 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1328) );
OR2_X1 U1008 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND3_X1 U1009 ( .A1(n1335), .A2(n1334), .A3(KEYINPUT19), .ZN(n1332) );
XOR2_X1 U1010 ( .A(n1080), .B(KEYINPUT24), .Z(n1334) );
NOR2_X1 U1011 ( .A1(G104), .A2(KEYINPUT51), .ZN(n1335) );
OR2_X1 U1012 ( .A1(n1336), .A2(KEYINPUT19), .ZN(n1331) );
INV_X1 U1013 ( .A(n1288), .ZN(n1259) );
NAND2_X1 U1014 ( .A1(n1087), .A2(n1337), .ZN(n1288) );
NAND4_X1 U1015 ( .A1(G953), .A2(G902), .A3(n1294), .A4(n1338), .ZN(n1337) );
INV_X1 U1016 ( .A(G898), .ZN(n1338) );
NAND3_X1 U1017 ( .A1(n1294), .A2(n1160), .A3(G952), .ZN(n1087) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1294) );
NAND2_X1 U1019 ( .A1(n1300), .A2(n1137), .ZN(n1296) );
XNOR2_X1 U1020 ( .A(n1339), .B(n1202), .ZN(n1137) );
AND2_X1 U1021 ( .A1(G217), .A2(n1313), .ZN(n1202) );
NAND2_X1 U1022 ( .A1(n1340), .A2(n1240), .ZN(n1313) );
XNOR2_X1 U1023 ( .A(G234), .B(KEYINPUT23), .ZN(n1340) );
NAND2_X1 U1024 ( .A1(n1200), .A2(n1240), .ZN(n1339) );
XOR2_X1 U1025 ( .A(n1341), .B(n1342), .Z(n1200) );
XOR2_X1 U1026 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1027 ( .A(G137), .B(G128), .Z(n1344) );
XOR2_X1 U1028 ( .A(KEYINPUT33), .B(KEYINPUT22), .Z(n1343) );
XOR2_X1 U1029 ( .A(n1345), .B(n1346), .Z(n1341) );
XNOR2_X1 U1030 ( .A(n1229), .B(n1347), .ZN(n1346) );
NOR2_X1 U1031 ( .A1(G119), .A2(KEYINPUT27), .ZN(n1347) );
XOR2_X1 U1032 ( .A(n1348), .B(n1349), .Z(n1345) );
AND3_X1 U1033 ( .A1(G221), .A2(n1160), .A3(G234), .ZN(n1349) );
XNOR2_X1 U1034 ( .A(n1143), .B(G472), .ZN(n1300) );
AND2_X1 U1035 ( .A1(n1350), .A2(n1240), .ZN(n1143) );
XNOR2_X1 U1036 ( .A(n1219), .B(n1215), .ZN(n1350) );
XNOR2_X1 U1037 ( .A(n1351), .B(G101), .ZN(n1215) );
NAND2_X1 U1038 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1039 ( .A(KEYINPUT54), .B(G210), .Z(n1353) );
XNOR2_X1 U1040 ( .A(n1354), .B(n1232), .ZN(n1219) );
XNOR2_X1 U1041 ( .A(n1170), .B(n1355), .ZN(n1232) );
NOR2_X1 U1042 ( .A1(G134), .A2(KEYINPUT62), .ZN(n1355) );
XNOR2_X1 U1043 ( .A(G131), .B(n1356), .ZN(n1170) );
XOR2_X1 U1044 ( .A(KEYINPUT55), .B(G137), .Z(n1356) );
XOR2_X1 U1045 ( .A(n1357), .B(n1358), .Z(n1354) );
NOR2_X1 U1046 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
XOR2_X1 U1047 ( .A(KEYINPUT8), .B(n1361), .Z(n1360) );
NOR2_X1 U1048 ( .A1(n1362), .A2(n1193), .ZN(n1361) );
AND2_X1 U1049 ( .A1(n1193), .A2(n1362), .ZN(n1359) );
INV_X1 U1050 ( .A(G113), .ZN(n1193) );
INV_X1 U1051 ( .A(n1103), .ZN(n1109) );
NAND2_X1 U1052 ( .A1(n1279), .A2(n1363), .ZN(n1103) );
XNOR2_X1 U1053 ( .A(KEYINPUT26), .B(n1306), .ZN(n1363) );
NAND3_X1 U1054 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1306) );
INV_X1 U1055 ( .A(n1145), .ZN(n1366) );
NOR2_X1 U1056 ( .A1(n1147), .A2(n1146), .ZN(n1145) );
NAND3_X1 U1057 ( .A1(n1146), .A2(n1147), .A3(n1367), .ZN(n1365) );
XNOR2_X1 U1058 ( .A(G478), .B(KEYINPUT7), .ZN(n1146) );
OR2_X1 U1059 ( .A1(n1367), .A2(n1147), .ZN(n1364) );
NAND2_X1 U1060 ( .A1(n1206), .A2(n1240), .ZN(n1147) );
XNOR2_X1 U1061 ( .A(n1368), .B(n1369), .ZN(n1206) );
XOR2_X1 U1062 ( .A(n1370), .B(n1371), .Z(n1369) );
XOR2_X1 U1063 ( .A(G128), .B(G122), .Z(n1371) );
XNOR2_X1 U1064 ( .A(n1372), .B(G134), .ZN(n1370) );
XOR2_X1 U1065 ( .A(n1373), .B(n1374), .Z(n1368) );
AND3_X1 U1066 ( .A1(G217), .A2(n1160), .A3(G234), .ZN(n1374) );
XNOR2_X1 U1067 ( .A(G116), .B(G107), .ZN(n1373) );
INV_X1 U1068 ( .A(KEYINPUT35), .ZN(n1367) );
XNOR2_X1 U1069 ( .A(n1148), .B(G475), .ZN(n1279) );
NOR2_X1 U1070 ( .A1(n1211), .A2(G902), .ZN(n1148) );
XNOR2_X1 U1071 ( .A(n1375), .B(n1376), .ZN(n1211) );
NOR2_X1 U1072 ( .A1(n1377), .A2(n1378), .ZN(n1376) );
XOR2_X1 U1073 ( .A(KEYINPUT37), .B(n1379), .Z(n1378) );
NOR2_X1 U1074 ( .A1(n1380), .A2(n1336), .ZN(n1379) );
INV_X1 U1075 ( .A(G104), .ZN(n1336) );
NOR2_X1 U1076 ( .A1(G104), .A2(n1381), .ZN(n1377) );
XNOR2_X1 U1077 ( .A(n1382), .B(KEYINPUT20), .ZN(n1381) );
NAND2_X1 U1078 ( .A1(KEYINPUT31), .A2(n1383), .ZN(n1375) );
XOR2_X1 U1079 ( .A(n1384), .B(n1385), .Z(n1383) );
XOR2_X1 U1080 ( .A(n1348), .B(n1386), .Z(n1385) );
NOR2_X1 U1081 ( .A1(G131), .A2(KEYINPUT6), .ZN(n1386) );
XNOR2_X1 U1082 ( .A(G146), .B(n1171), .ZN(n1348) );
XOR2_X1 U1083 ( .A(G125), .B(G140), .Z(n1171) );
XNOR2_X1 U1084 ( .A(n1387), .B(n1372), .ZN(n1384) );
NAND2_X1 U1085 ( .A1(G214), .A2(n1352), .ZN(n1387) );
NOR2_X1 U1086 ( .A1(G953), .A2(G237), .ZN(n1352) );
XOR2_X1 U1087 ( .A(n1257), .B(KEYINPUT39), .Z(n1311) );
XOR2_X1 U1088 ( .A(n1304), .B(KEYINPUT25), .Z(n1257) );
NAND2_X1 U1089 ( .A1(n1094), .A2(n1108), .ZN(n1304) );
NAND2_X1 U1090 ( .A1(G214), .A2(n1388), .ZN(n1108) );
NAND2_X1 U1091 ( .A1(n1389), .A2(n1390), .ZN(n1094) );
OR2_X1 U1092 ( .A1(n1140), .A2(n1139), .ZN(n1390) );
INV_X1 U1093 ( .A(n1391), .ZN(n1139) );
XOR2_X1 U1094 ( .A(n1392), .B(KEYINPUT9), .Z(n1389) );
NAND2_X1 U1095 ( .A1(n1393), .A2(n1140), .ZN(n1392) );
NAND2_X1 U1096 ( .A1(n1394), .A2(n1240), .ZN(n1140) );
XOR2_X1 U1097 ( .A(n1395), .B(n1234), .Z(n1394) );
XNOR2_X1 U1098 ( .A(n1396), .B(n1397), .ZN(n1234) );
XNOR2_X1 U1099 ( .A(n1229), .B(n1191), .ZN(n1397) );
NOR2_X1 U1100 ( .A1(KEYINPUT36), .A2(n1362), .ZN(n1191) );
XNOR2_X1 U1101 ( .A(G116), .B(G119), .ZN(n1362) );
INV_X1 U1102 ( .A(G110), .ZN(n1229) );
XNOR2_X1 U1103 ( .A(n1185), .B(n1380), .ZN(n1396) );
INV_X1 U1104 ( .A(n1382), .ZN(n1380) );
XOR2_X1 U1105 ( .A(G113), .B(G122), .Z(n1382) );
XNOR2_X1 U1106 ( .A(G101), .B(n1398), .ZN(n1185) );
XNOR2_X1 U1107 ( .A(n1080), .B(G104), .ZN(n1398) );
INV_X1 U1108 ( .A(G107), .ZN(n1080) );
NAND2_X1 U1109 ( .A1(n1399), .A2(n1239), .ZN(n1395) );
NAND3_X1 U1110 ( .A1(G224), .A2(n1160), .A3(n1400), .ZN(n1239) );
XOR2_X1 U1111 ( .A(n1357), .B(G125), .Z(n1400) );
XOR2_X1 U1112 ( .A(n1238), .B(KEYINPUT60), .Z(n1399) );
NAND2_X1 U1113 ( .A1(n1401), .A2(n1402), .ZN(n1238) );
NAND2_X1 U1114 ( .A1(G224), .A2(n1160), .ZN(n1402) );
INV_X1 U1115 ( .A(G953), .ZN(n1160) );
XNOR2_X1 U1116 ( .A(G125), .B(n1357), .ZN(n1401) );
NAND2_X1 U1117 ( .A1(n1403), .A2(n1404), .ZN(n1357) );
NAND2_X1 U1118 ( .A1(G128), .A2(n1405), .ZN(n1404) );
XOR2_X1 U1119 ( .A(KEYINPUT2), .B(n1406), .Z(n1403) );
NOR2_X1 U1120 ( .A1(G128), .A2(n1405), .ZN(n1406) );
NAND2_X1 U1121 ( .A1(n1407), .A2(n1408), .ZN(n1405) );
NAND2_X1 U1122 ( .A1(G143), .A2(n1271), .ZN(n1408) );
INV_X1 U1123 ( .A(G146), .ZN(n1271) );
XOR2_X1 U1124 ( .A(n1409), .B(KEYINPUT1), .Z(n1407) );
NAND2_X1 U1125 ( .A1(G146), .A2(n1372), .ZN(n1409) );
INV_X1 U1126 ( .A(G143), .ZN(n1372) );
XNOR2_X1 U1127 ( .A(KEYINPUT16), .B(n1391), .ZN(n1393) );
NAND2_X1 U1128 ( .A1(G210), .A2(n1388), .ZN(n1391) );
NAND2_X1 U1129 ( .A1(n1410), .A2(n1240), .ZN(n1388) );
INV_X1 U1130 ( .A(G902), .ZN(n1240) );
INV_X1 U1131 ( .A(G237), .ZN(n1410) );
endmodule


