//Key = 1111011110001110100110100110111001011100100110001010101001111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410;

XOR2_X1 U771 ( .A(G107), .B(n1059), .Z(G9) );
NOR2_X1 U772 ( .A1(n1060), .A2(n1061), .ZN(G75) );
XOR2_X1 U773 ( .A(KEYINPUT51), .B(n1062), .Z(n1061) );
AND3_X1 U774 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NOR4_X1 U775 ( .A1(n1066), .A2(n1067), .A3(n1065), .A4(n1068), .ZN(n1060) );
INV_X1 U776 ( .A(G952), .ZN(n1065) );
NAND4_X1 U777 ( .A1(n1069), .A2(n1070), .A3(n1063), .A4(n1064), .ZN(n1066) );
NAND4_X1 U778 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1063) );
NOR4_X1 U779 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
XOR2_X1 U780 ( .A(n1079), .B(n1080), .Z(n1078) );
XOR2_X1 U781 ( .A(n1081), .B(n1082), .Z(n1077) );
XNOR2_X1 U782 ( .A(G475), .B(KEYINPUT34), .ZN(n1082) );
XOR2_X1 U783 ( .A(n1083), .B(n1084), .Z(n1076) );
XNOR2_X1 U784 ( .A(n1085), .B(KEYINPUT50), .ZN(n1084) );
NAND2_X1 U785 ( .A1(KEYINPUT2), .A2(n1086), .ZN(n1083) );
NOR2_X1 U786 ( .A1(n1087), .A2(n1088), .ZN(n1073) );
XOR2_X1 U787 ( .A(n1089), .B(KEYINPUT11), .Z(n1088) );
NAND3_X1 U788 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
OR2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND3_X1 U790 ( .A1(n1094), .A2(n1093), .A3(G472), .ZN(n1091) );
NAND2_X1 U791 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
NAND2_X1 U792 ( .A1(n1097), .A2(n1093), .ZN(n1095) );
INV_X1 U793 ( .A(KEYINPUT32), .ZN(n1093) );
XOR2_X1 U794 ( .A(n1094), .B(KEYINPUT49), .Z(n1097) );
XNOR2_X1 U795 ( .A(n1098), .B(n1099), .ZN(n1087) );
NAND2_X1 U796 ( .A1(KEYINPUT52), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U797 ( .A(KEYINPUT1), .B(n1101), .ZN(n1100) );
NAND2_X1 U798 ( .A1(n1102), .A2(n1103), .ZN(n1070) );
NAND2_X1 U799 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND3_X1 U800 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
NAND2_X1 U801 ( .A1(n1109), .A2(n1110), .ZN(n1104) );
NAND2_X1 U802 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U804 ( .A(KEYINPUT8), .B(n1115), .Z(n1114) );
NAND2_X1 U805 ( .A1(n1107), .A2(n1116), .ZN(n1069) );
NAND3_X1 U806 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
NAND2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND4_X1 U808 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1102), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1125), .A2(n1106), .ZN(n1124) );
NAND4_X1 U810 ( .A1(n1126), .A2(n1122), .A3(n1102), .A4(n1071), .ZN(n1118) );
INV_X1 U811 ( .A(n1127), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NOR3_X1 U813 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1125), .A2(n1133), .ZN(n1128) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1121), .ZN(n1133) );
INV_X1 U816 ( .A(KEYINPUT33), .ZN(n1121) );
NAND2_X1 U817 ( .A1(n1109), .A2(n1135), .ZN(n1117) );
NAND2_X1 U818 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U819 ( .A1(n1138), .A2(n1075), .ZN(n1137) );
AND2_X1 U820 ( .A1(n1108), .A2(n1071), .ZN(n1109) );
NOR3_X1 U821 ( .A1(n1130), .A2(n1134), .A3(n1127), .ZN(n1108) );
XOR2_X1 U822 ( .A(n1139), .B(n1140), .Z(G72) );
XOR2_X1 U823 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U824 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
AND2_X1 U825 ( .A1(G227), .A2(G900), .ZN(n1143) );
NAND2_X1 U826 ( .A1(n1145), .A2(n1146), .ZN(n1141) );
INV_X1 U827 ( .A(n1147), .ZN(n1146) );
XOR2_X1 U828 ( .A(n1148), .B(n1149), .Z(n1145) );
XOR2_X1 U829 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U830 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U831 ( .A(n1154), .B(KEYINPUT61), .Z(n1152) );
NAND2_X1 U832 ( .A1(n1155), .A2(n1156), .ZN(n1150) );
NAND2_X1 U833 ( .A1(G131), .A2(n1157), .ZN(n1156) );
XOR2_X1 U834 ( .A(KEYINPUT44), .B(n1158), .Z(n1155) );
NOR2_X1 U835 ( .A1(G131), .A2(n1157), .ZN(n1158) );
XOR2_X1 U836 ( .A(G137), .B(G134), .Z(n1157) );
NAND4_X1 U837 ( .A1(KEYINPUT37), .A2(n1064), .A3(n1159), .A4(n1160), .ZN(n1139) );
NAND3_X1 U838 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
INV_X1 U839 ( .A(KEYINPUT60), .ZN(n1163) );
NAND2_X1 U840 ( .A1(KEYINPUT60), .A2(n1164), .ZN(n1159) );
XOR2_X1 U841 ( .A(n1165), .B(n1166), .Z(G69) );
XOR2_X1 U842 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1144), .ZN(n1168) );
XOR2_X1 U844 ( .A(G953), .B(KEYINPUT19), .Z(n1144) );
AND2_X1 U845 ( .A1(G224), .A2(G898), .ZN(n1169) );
NAND2_X1 U846 ( .A1(n1170), .A2(n1171), .ZN(n1167) );
INV_X1 U847 ( .A(n1172), .ZN(n1171) );
NAND2_X1 U848 ( .A1(n1064), .A2(n1067), .ZN(n1165) );
NOR2_X1 U849 ( .A1(n1173), .A2(n1174), .ZN(G66) );
XOR2_X1 U850 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U851 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U852 ( .A1(n1173), .A2(n1179), .ZN(G63) );
XOR2_X1 U853 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U854 ( .A1(n1079), .A2(n1178), .ZN(n1181) );
INV_X1 U855 ( .A(G478), .ZN(n1079) );
NOR2_X1 U856 ( .A1(n1173), .A2(n1182), .ZN(G60) );
XOR2_X1 U857 ( .A(n1183), .B(n1184), .Z(n1182) );
XNOR2_X1 U858 ( .A(n1185), .B(KEYINPUT20), .ZN(n1184) );
NAND3_X1 U859 ( .A1(n1186), .A2(G475), .A3(KEYINPUT25), .ZN(n1185) );
INV_X1 U860 ( .A(n1178), .ZN(n1186) );
XOR2_X1 U861 ( .A(G104), .B(n1187), .Z(G6) );
NOR2_X1 U862 ( .A1(n1173), .A2(n1188), .ZN(G57) );
NOR2_X1 U863 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U864 ( .A(KEYINPUT55), .B(n1191), .Z(n1190) );
NOR2_X1 U865 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
AND2_X1 U866 ( .A1(n1193), .A2(n1192), .ZN(n1189) );
AND2_X1 U867 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
NAND2_X1 U868 ( .A1(KEYINPUT15), .A2(G101), .ZN(n1195) );
NAND2_X1 U869 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
INV_X1 U870 ( .A(KEYINPUT15), .ZN(n1197) );
NAND2_X1 U871 ( .A1(n1198), .A2(n1199), .ZN(n1193) );
NAND2_X1 U872 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U873 ( .A(KEYINPUT16), .B(n1202), .Z(n1200) );
NOR2_X1 U874 ( .A1(n1096), .A2(n1178), .ZN(n1202) );
OR3_X1 U875 ( .A1(n1178), .A2(n1096), .A3(n1201), .ZN(n1198) );
XOR2_X1 U876 ( .A(n1203), .B(n1204), .Z(n1201) );
NOR2_X1 U877 ( .A1(KEYINPUT18), .A2(n1205), .ZN(n1204) );
INV_X1 U878 ( .A(G472), .ZN(n1096) );
NOR2_X1 U879 ( .A1(n1173), .A2(n1206), .ZN(G54) );
XOR2_X1 U880 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U881 ( .A(n1148), .B(n1209), .Z(n1208) );
XOR2_X1 U882 ( .A(n1210), .B(n1211), .Z(n1209) );
NOR2_X1 U883 ( .A1(n1086), .A2(n1178), .ZN(n1210) );
XOR2_X1 U884 ( .A(G146), .B(n1212), .Z(n1148) );
XOR2_X1 U885 ( .A(n1213), .B(n1214), .Z(n1207) );
XOR2_X1 U886 ( .A(KEYINPUT17), .B(n1215), .Z(n1214) );
NOR4_X1 U887 ( .A1(n1216), .A2(n1217), .A3(KEYINPUT4), .A4(n1218), .ZN(n1215) );
INV_X1 U888 ( .A(n1219), .ZN(n1218) );
NOR3_X1 U889 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1217) );
NOR2_X1 U890 ( .A1(G110), .A2(n1223), .ZN(n1216) );
XOR2_X1 U891 ( .A(n1224), .B(n1221), .Z(n1223) );
NOR2_X1 U892 ( .A1(KEYINPUT24), .A2(n1225), .ZN(n1213) );
XOR2_X1 U893 ( .A(G101), .B(n1226), .Z(n1225) );
XOR2_X1 U894 ( .A(G107), .B(G104), .Z(n1226) );
NOR2_X1 U895 ( .A1(n1173), .A2(n1227), .ZN(G51) );
XOR2_X1 U896 ( .A(n1228), .B(n1170), .Z(n1227) );
XOR2_X1 U897 ( .A(n1229), .B(n1230), .Z(n1228) );
NOR3_X1 U898 ( .A1(n1178), .A2(KEYINPUT62), .A3(n1099), .ZN(n1230) );
NAND2_X1 U899 ( .A1(G902), .A2(n1231), .ZN(n1178) );
NAND2_X1 U900 ( .A1(n1232), .A2(n1164), .ZN(n1231) );
INV_X1 U901 ( .A(n1068), .ZN(n1164) );
NAND4_X1 U902 ( .A1(n1162), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1068) );
NOR4_X1 U903 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NOR2_X1 U904 ( .A1(n1240), .A2(n1161), .ZN(n1234) );
NAND2_X1 U905 ( .A1(n1241), .A2(n1242), .ZN(n1162) );
XOR2_X1 U906 ( .A(n1243), .B(KEYINPUT12), .Z(n1241) );
XOR2_X1 U907 ( .A(n1067), .B(KEYINPUT22), .Z(n1232) );
NAND4_X1 U908 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1067) );
NOR4_X1 U909 ( .A1(n1059), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1247) );
AND3_X1 U910 ( .A1(n1132), .A2(n1102), .A3(n1251), .ZN(n1059) );
NOR2_X1 U911 ( .A1(n1187), .A2(n1252), .ZN(n1246) );
AND3_X1 U912 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1252) );
AND3_X1 U913 ( .A1(n1251), .A2(n1102), .A3(n1131), .ZN(n1187) );
NAND2_X1 U914 ( .A1(n1256), .A2(n1257), .ZN(n1229) );
INV_X1 U915 ( .A(n1258), .ZN(n1256) );
NOR2_X1 U916 ( .A1(n1064), .A2(G952), .ZN(n1173) );
XOR2_X1 U917 ( .A(G146), .B(n1259), .Z(G48) );
NOR3_X1 U918 ( .A1(n1243), .A2(KEYINPUT46), .A3(n1111), .ZN(n1259) );
NAND4_X1 U919 ( .A1(n1260), .A2(n1131), .A3(n1254), .A4(n1075), .ZN(n1243) );
XOR2_X1 U920 ( .A(n1240), .B(n1261), .Z(G45) );
NOR2_X1 U921 ( .A1(KEYINPUT39), .A2(n1262), .ZN(n1261) );
INV_X1 U922 ( .A(G143), .ZN(n1262) );
AND4_X1 U923 ( .A1(n1260), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(n1240) );
NOR2_X1 U924 ( .A1(n1266), .A2(n1111), .ZN(n1264) );
NAND3_X1 U925 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(G42) );
NAND2_X1 U926 ( .A1(n1239), .A2(n1270), .ZN(n1269) );
NAND2_X1 U927 ( .A1(KEYINPUT45), .A2(n1271), .ZN(n1268) );
NAND2_X1 U928 ( .A1(n1272), .A2(G140), .ZN(n1271) );
XNOR2_X1 U929 ( .A(n1239), .B(KEYINPUT9), .ZN(n1272) );
NAND2_X1 U930 ( .A1(n1273), .A2(n1274), .ZN(n1267) );
INV_X1 U931 ( .A(KEYINPUT45), .ZN(n1274) );
NAND2_X1 U932 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
OR3_X1 U933 ( .A1(n1270), .A2(n1239), .A3(KEYINPUT9), .ZN(n1276) );
NAND2_X1 U934 ( .A1(KEYINPUT9), .A2(n1239), .ZN(n1275) );
AND3_X1 U935 ( .A1(n1138), .A2(n1075), .A3(n1277), .ZN(n1239) );
XOR2_X1 U936 ( .A(n1278), .B(n1233), .Z(G39) );
NAND4_X1 U937 ( .A1(n1107), .A2(n1260), .A3(n1255), .A4(n1254), .ZN(n1233) );
XOR2_X1 U938 ( .A(n1279), .B(n1280), .Z(G36) );
XOR2_X1 U939 ( .A(n1281), .B(KEYINPUT21), .Z(n1280) );
NAND2_X1 U940 ( .A1(KEYINPUT29), .A2(n1238), .ZN(n1279) );
AND4_X1 U941 ( .A1(n1107), .A2(n1260), .A3(n1263), .A4(n1132), .ZN(n1238) );
XNOR2_X1 U942 ( .A(G131), .B(n1282), .ZN(G33) );
NOR2_X1 U943 ( .A1(n1237), .A2(KEYINPUT10), .ZN(n1282) );
AND2_X1 U944 ( .A1(n1277), .A2(n1263), .ZN(n1237) );
AND3_X1 U945 ( .A1(n1260), .A2(n1131), .A3(n1107), .ZN(n1277) );
NOR2_X1 U946 ( .A1(n1115), .A2(n1113), .ZN(n1107) );
INV_X1 U947 ( .A(n1072), .ZN(n1113) );
NAND2_X1 U948 ( .A1(n1283), .A2(n1284), .ZN(G30) );
NAND2_X1 U949 ( .A1(n1236), .A2(n1285), .ZN(n1284) );
XOR2_X1 U950 ( .A(KEYINPUT59), .B(n1286), .Z(n1283) );
NOR2_X1 U951 ( .A1(n1236), .A2(n1285), .ZN(n1286) );
AND4_X1 U952 ( .A1(n1254), .A2(n1075), .A3(n1242), .A4(n1287), .ZN(n1236) );
AND2_X1 U953 ( .A1(n1132), .A2(n1260), .ZN(n1287) );
NOR3_X1 U954 ( .A1(n1106), .A2(n1125), .A3(n1288), .ZN(n1260) );
XOR2_X1 U955 ( .A(n1289), .B(n1244), .Z(G3) );
NAND3_X1 U956 ( .A1(n1123), .A2(n1251), .A3(n1263), .ZN(n1244) );
INV_X1 U957 ( .A(n1134), .ZN(n1123) );
XOR2_X1 U958 ( .A(G125), .B(n1161), .Z(G27) );
AND4_X1 U959 ( .A1(n1138), .A2(n1125), .A3(n1131), .A4(n1290), .ZN(n1161) );
NOR4_X1 U960 ( .A1(n1106), .A2(n1291), .A3(n1288), .A4(n1111), .ZN(n1290) );
AND2_X1 U961 ( .A1(n1292), .A2(n1293), .ZN(n1288) );
NAND3_X1 U962 ( .A1(G902), .A2(n1294), .A3(n1147), .ZN(n1293) );
NOR2_X1 U963 ( .A1(n1064), .A2(G900), .ZN(n1147) );
XOR2_X1 U964 ( .A(n1127), .B(KEYINPUT47), .Z(n1292) );
INV_X1 U965 ( .A(n1071), .ZN(n1106) );
XNOR2_X1 U966 ( .A(G122), .B(n1245), .ZN(G24) );
NAND4_X1 U967 ( .A1(n1265), .A2(n1253), .A3(n1102), .A4(n1295), .ZN(n1245) );
NOR2_X1 U968 ( .A1(n1075), .A2(n1254), .ZN(n1102) );
XNOR2_X1 U969 ( .A(G119), .B(n1296), .ZN(G21) );
NAND4_X1 U970 ( .A1(KEYINPUT48), .A2(n1253), .A3(n1255), .A4(n1254), .ZN(n1296) );
XOR2_X1 U971 ( .A(G116), .B(n1250), .Z(G18) );
AND3_X1 U972 ( .A1(n1263), .A2(n1132), .A3(n1253), .ZN(n1250) );
NOR2_X1 U973 ( .A1(n1265), .A2(n1266), .ZN(n1132) );
XOR2_X1 U974 ( .A(G113), .B(n1249), .Z(G15) );
AND3_X1 U975 ( .A1(n1131), .A2(n1263), .A3(n1253), .ZN(n1249) );
AND3_X1 U976 ( .A1(n1297), .A2(n1071), .A3(n1125), .ZN(n1253) );
INV_X1 U977 ( .A(n1130), .ZN(n1125) );
INV_X1 U978 ( .A(n1136), .ZN(n1263) );
NAND2_X1 U979 ( .A1(n1291), .A2(n1254), .ZN(n1136) );
INV_X1 U980 ( .A(n1138), .ZN(n1254) );
NOR2_X1 U981 ( .A1(n1298), .A2(n1295), .ZN(n1131) );
INV_X1 U982 ( .A(n1266), .ZN(n1295) );
XOR2_X1 U983 ( .A(G110), .B(n1248), .Z(G12) );
AND3_X1 U984 ( .A1(n1138), .A2(n1251), .A3(n1255), .ZN(n1248) );
NOR2_X1 U985 ( .A1(n1134), .A2(n1291), .ZN(n1255) );
INV_X1 U986 ( .A(n1075), .ZN(n1291) );
NAND3_X1 U987 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1075) );
NAND2_X1 U988 ( .A1(G217), .A2(G902), .ZN(n1301) );
OR3_X1 U989 ( .A1(n1175), .A2(G902), .A3(n1302), .ZN(n1300) );
NAND2_X1 U990 ( .A1(n1302), .A2(n1175), .ZN(n1299) );
XOR2_X1 U991 ( .A(n1303), .B(n1304), .Z(n1175) );
XOR2_X1 U992 ( .A(KEYINPUT31), .B(G137), .Z(n1304) );
XOR2_X1 U993 ( .A(n1305), .B(n1306), .Z(n1303) );
AND2_X1 U994 ( .A1(G221), .A2(n1307), .ZN(n1306) );
NAND2_X1 U995 ( .A1(n1308), .A2(KEYINPUT26), .ZN(n1305) );
XOR2_X1 U996 ( .A(n1309), .B(n1310), .Z(n1308) );
XOR2_X1 U997 ( .A(G110), .B(n1311), .Z(n1310) );
NOR2_X1 U998 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
XOR2_X1 U999 ( .A(n1314), .B(KEYINPUT5), .Z(n1313) );
NAND2_X1 U1000 ( .A1(G125), .A2(n1315), .ZN(n1314) );
NOR2_X1 U1001 ( .A1(n1316), .A2(n1315), .ZN(n1312) );
XOR2_X1 U1002 ( .A(KEYINPUT57), .B(G140), .Z(n1315) );
XOR2_X1 U1003 ( .A(KEYINPUT38), .B(G125), .Z(n1316) );
XNOR2_X1 U1004 ( .A(G119), .B(n1317), .ZN(n1309) );
XOR2_X1 U1005 ( .A(G146), .B(G128), .Z(n1317) );
NOR2_X1 U1006 ( .A1(n1177), .A2(G234), .ZN(n1302) );
INV_X1 U1007 ( .A(G217), .ZN(n1177) );
NAND2_X1 U1008 ( .A1(n1266), .A2(n1298), .ZN(n1134) );
INV_X1 U1009 ( .A(n1265), .ZN(n1298) );
XOR2_X1 U1010 ( .A(n1318), .B(G475), .Z(n1265) );
NAND2_X1 U1011 ( .A1(KEYINPUT6), .A2(n1081), .ZN(n1318) );
NAND2_X1 U1012 ( .A1(n1183), .A2(n1319), .ZN(n1081) );
XOR2_X1 U1013 ( .A(n1320), .B(n1321), .Z(n1183) );
XNOR2_X1 U1014 ( .A(n1322), .B(n1323), .ZN(n1321) );
NAND2_X1 U1015 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1016 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
INV_X1 U1017 ( .A(KEYINPUT27), .ZN(n1327) );
NAND2_X1 U1018 ( .A1(n1153), .A2(n1154), .ZN(n1326) );
NAND2_X1 U1019 ( .A1(G140), .A2(n1328), .ZN(n1154) );
NAND2_X1 U1020 ( .A1(G125), .A2(n1270), .ZN(n1153) );
NAND2_X1 U1021 ( .A1(KEYINPUT27), .A2(n1329), .ZN(n1324) );
XOR2_X1 U1022 ( .A(n1328), .B(G140), .Z(n1329) );
XNOR2_X1 U1023 ( .A(n1330), .B(n1331), .ZN(n1320) );
NAND2_X1 U1024 ( .A1(n1332), .A2(KEYINPUT43), .ZN(n1331) );
XOR2_X1 U1025 ( .A(n1333), .B(G122), .Z(n1332) );
NAND2_X1 U1026 ( .A1(KEYINPUT3), .A2(n1334), .ZN(n1333) );
INV_X1 U1027 ( .A(G113), .ZN(n1334) );
NAND2_X1 U1028 ( .A1(KEYINPUT0), .A2(n1335), .ZN(n1330) );
XOR2_X1 U1029 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1030 ( .A(G143), .B(G131), .Z(n1337) );
AND2_X1 U1031 ( .A1(G214), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1032 ( .A(n1339), .B(G478), .Z(n1266) );
NAND2_X1 U1033 ( .A1(KEYINPUT40), .A2(n1340), .ZN(n1339) );
INV_X1 U1034 ( .A(n1080), .ZN(n1340) );
NAND2_X1 U1035 ( .A1(n1341), .A2(n1319), .ZN(n1080) );
XOR2_X1 U1036 ( .A(n1180), .B(KEYINPUT30), .Z(n1341) );
XOR2_X1 U1037 ( .A(n1342), .B(n1343), .Z(n1180) );
XOR2_X1 U1038 ( .A(n1281), .B(n1344), .Z(n1343) );
NAND2_X1 U1039 ( .A1(G217), .A2(n1307), .ZN(n1344) );
AND2_X1 U1040 ( .A1(G234), .A2(n1064), .ZN(n1307) );
INV_X1 U1041 ( .A(G134), .ZN(n1281) );
XNOR2_X1 U1042 ( .A(n1345), .B(n1346), .ZN(n1342) );
AND3_X1 U1043 ( .A1(n1071), .A2(n1130), .A3(n1297), .ZN(n1251) );
AND2_X1 U1044 ( .A1(n1242), .A2(n1347), .ZN(n1297) );
NAND2_X1 U1045 ( .A1(n1127), .A2(n1348), .ZN(n1347) );
NAND3_X1 U1046 ( .A1(n1172), .A2(n1294), .A3(G902), .ZN(n1348) );
NOR2_X1 U1047 ( .A1(n1064), .A2(G898), .ZN(n1172) );
NAND3_X1 U1048 ( .A1(n1294), .A2(n1064), .A3(G952), .ZN(n1127) );
NAND2_X1 U1049 ( .A1(G234), .A2(G237), .ZN(n1294) );
INV_X1 U1050 ( .A(n1111), .ZN(n1242) );
NAND2_X1 U1051 ( .A1(n1115), .A2(n1072), .ZN(n1111) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1349), .ZN(n1072) );
XOR2_X1 U1053 ( .A(n1101), .B(n1099), .Z(n1115) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1349), .ZN(n1099) );
NAND2_X1 U1055 ( .A1(n1350), .A2(n1319), .ZN(n1349) );
XNOR2_X1 U1056 ( .A(G237), .B(KEYINPUT53), .ZN(n1350) );
NAND2_X1 U1057 ( .A1(n1351), .A2(n1319), .ZN(n1101) );
XNOR2_X1 U1058 ( .A(n1352), .B(n1170), .ZN(n1351) );
XNOR2_X1 U1059 ( .A(n1353), .B(n1354), .ZN(n1170) );
XOR2_X1 U1060 ( .A(n1355), .B(n1346), .Z(n1354) );
XOR2_X1 U1061 ( .A(G116), .B(G122), .Z(n1346) );
XOR2_X1 U1062 ( .A(n1356), .B(n1357), .Z(n1353) );
XOR2_X1 U1063 ( .A(G110), .B(G101), .Z(n1357) );
NAND3_X1 U1064 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1356) );
NAND2_X1 U1065 ( .A1(KEYINPUT56), .A2(G104), .ZN(n1360) );
NAND3_X1 U1066 ( .A1(n1361), .A2(n1362), .A3(G107), .ZN(n1359) );
INV_X1 U1067 ( .A(G104), .ZN(n1361) );
NAND2_X1 U1068 ( .A1(n1363), .A2(n1364), .ZN(n1358) );
NAND2_X1 U1069 ( .A1(n1365), .A2(n1362), .ZN(n1363) );
INV_X1 U1070 ( .A(KEYINPUT56), .ZN(n1362) );
XOR2_X1 U1071 ( .A(KEYINPUT63), .B(G104), .Z(n1365) );
NAND3_X1 U1072 ( .A1(n1366), .A2(n1367), .A3(n1257), .ZN(n1352) );
NAND3_X1 U1073 ( .A1(n1368), .A2(n1369), .A3(G125), .ZN(n1257) );
NAND2_X1 U1074 ( .A1(n1370), .A2(n1371), .ZN(n1367) );
INV_X1 U1075 ( .A(KEYINPUT28), .ZN(n1371) );
XOR2_X1 U1076 ( .A(n1372), .B(n1373), .Z(n1370) );
NAND2_X1 U1077 ( .A1(n1374), .A2(n1328), .ZN(n1372) );
NAND2_X1 U1078 ( .A1(KEYINPUT28), .A2(n1258), .ZN(n1366) );
NAND2_X1 U1079 ( .A1(n1375), .A2(n1376), .ZN(n1258) );
NAND2_X1 U1080 ( .A1(n1377), .A2(n1328), .ZN(n1376) );
INV_X1 U1081 ( .A(G125), .ZN(n1328) );
XOR2_X1 U1082 ( .A(n1369), .B(n1368), .Z(n1377) );
INV_X1 U1083 ( .A(n1374), .ZN(n1368) );
NAND3_X1 U1084 ( .A1(n1373), .A2(n1374), .A3(G125), .ZN(n1375) );
INV_X1 U1085 ( .A(n1369), .ZN(n1373) );
NAND2_X1 U1086 ( .A1(G224), .A2(n1064), .ZN(n1369) );
NAND2_X1 U1087 ( .A1(n1378), .A2(n1379), .ZN(n1130) );
NAND2_X1 U1088 ( .A1(n1085), .A2(n1086), .ZN(n1379) );
XOR2_X1 U1089 ( .A(KEYINPUT35), .B(n1380), .Z(n1378) );
NOR2_X1 U1090 ( .A1(n1085), .A2(n1086), .ZN(n1380) );
INV_X1 U1091 ( .A(G469), .ZN(n1086) );
AND2_X1 U1092 ( .A1(n1381), .A2(n1319), .ZN(n1085) );
XOR2_X1 U1093 ( .A(n1382), .B(n1383), .Z(n1381) );
XOR2_X1 U1094 ( .A(n1384), .B(n1322), .Z(n1383) );
XOR2_X1 U1095 ( .A(G146), .B(G104), .Z(n1322) );
XNOR2_X1 U1096 ( .A(n1211), .B(n1345), .ZN(n1384) );
XNOR2_X1 U1097 ( .A(n1364), .B(n1212), .ZN(n1345) );
XOR2_X1 U1098 ( .A(G128), .B(G143), .Z(n1212) );
INV_X1 U1099 ( .A(G107), .ZN(n1364) );
XOR2_X1 U1100 ( .A(n1385), .B(n1386), .Z(n1382) );
XOR2_X1 U1101 ( .A(KEYINPUT42), .B(G101), .Z(n1386) );
NAND3_X1 U1102 ( .A1(n1387), .A2(n1388), .A3(n1219), .ZN(n1385) );
NAND3_X1 U1103 ( .A1(G110), .A2(n1222), .A3(n1221), .ZN(n1219) );
NAND2_X1 U1104 ( .A1(n1389), .A2(n1220), .ZN(n1388) );
INV_X1 U1105 ( .A(G110), .ZN(n1220) );
XOR2_X1 U1106 ( .A(n1224), .B(n1390), .Z(n1389) );
NAND2_X1 U1107 ( .A1(n1391), .A2(G110), .ZN(n1387) );
NAND2_X1 U1108 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NAND2_X1 U1109 ( .A1(n1222), .A2(n1394), .ZN(n1393) );
NAND2_X1 U1110 ( .A1(n1390), .A2(n1224), .ZN(n1392) );
INV_X1 U1111 ( .A(n1222), .ZN(n1224) );
NAND2_X1 U1112 ( .A1(G227), .A2(n1064), .ZN(n1222) );
NOR2_X1 U1113 ( .A1(n1394), .A2(n1221), .ZN(n1390) );
XOR2_X1 U1114 ( .A(n1270), .B(KEYINPUT41), .Z(n1221) );
INV_X1 U1115 ( .A(G140), .ZN(n1270) );
INV_X1 U1116 ( .A(KEYINPUT58), .ZN(n1394) );
NAND2_X1 U1117 ( .A1(G221), .A2(n1395), .ZN(n1071) );
NAND2_X1 U1118 ( .A1(G234), .A2(n1319), .ZN(n1395) );
XOR2_X1 U1119 ( .A(n1094), .B(G472), .Z(n1138) );
NAND2_X1 U1120 ( .A1(n1396), .A2(n1319), .ZN(n1094) );
INV_X1 U1121 ( .A(G902), .ZN(n1319) );
XOR2_X1 U1122 ( .A(n1397), .B(n1398), .Z(n1396) );
XNOR2_X1 U1123 ( .A(KEYINPUT7), .B(n1196), .ZN(n1398) );
NAND2_X1 U1124 ( .A1(n1399), .A2(n1400), .ZN(n1196) );
NAND3_X1 U1125 ( .A1(G210), .A2(G101), .A3(n1338), .ZN(n1400) );
NAND2_X1 U1126 ( .A1(n1289), .A2(n1401), .ZN(n1399) );
NAND2_X1 U1127 ( .A1(n1338), .A2(G210), .ZN(n1401) );
AND2_X1 U1128 ( .A1(n1402), .A2(n1064), .ZN(n1338) );
INV_X1 U1129 ( .A(G953), .ZN(n1064) );
XOR2_X1 U1130 ( .A(KEYINPUT13), .B(G237), .Z(n1402) );
INV_X1 U1131 ( .A(G101), .ZN(n1289) );
XOR2_X1 U1132 ( .A(n1205), .B(n1403), .Z(n1397) );
INV_X1 U1133 ( .A(n1203), .ZN(n1403) );
XOR2_X1 U1134 ( .A(n1404), .B(n1355), .Z(n1203) );
XOR2_X1 U1135 ( .A(G113), .B(G119), .Z(n1355) );
INV_X1 U1136 ( .A(G116), .ZN(n1404) );
XOR2_X1 U1137 ( .A(n1211), .B(n1374), .Z(n1205) );
XOR2_X1 U1138 ( .A(n1405), .B(n1406), .Z(n1374) );
NOR2_X1 U1139 ( .A1(KEYINPUT23), .A2(n1285), .ZN(n1406) );
INV_X1 U1140 ( .A(G128), .ZN(n1285) );
XOR2_X1 U1141 ( .A(n1407), .B(G146), .Z(n1405) );
NAND2_X1 U1142 ( .A1(KEYINPUT54), .A2(n1408), .ZN(n1407) );
XOR2_X1 U1143 ( .A(KEYINPUT14), .B(G143), .Z(n1408) );
XNOR2_X1 U1144 ( .A(n1409), .B(n1410), .ZN(n1211) );
XOR2_X1 U1145 ( .A(G134), .B(G131), .Z(n1410) );
NAND2_X1 U1146 ( .A1(KEYINPUT36), .A2(n1278), .ZN(n1409) );
INV_X1 U1147 ( .A(G137), .ZN(n1278) );
endmodule


