//Key = 1100001101010010110101000100111110001000011011000101101100001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340;

XOR2_X1 U740 ( .A(n1026), .B(n1027), .Z(G9) );
NAND4_X1 U741 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
OR2_X1 U742 ( .A1(n1032), .A2(KEYINPUT35), .ZN(n1031) );
NAND2_X1 U743 ( .A1(KEYINPUT35), .A2(n1033), .ZN(n1030) );
OR3_X1 U744 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NOR2_X1 U745 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U747 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U748 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
XOR2_X1 U749 ( .A(KEYINPUT8), .B(n1046), .Z(n1045) );
NOR4_X1 U750 ( .A1(n1034), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1046) );
NOR4_X1 U751 ( .A1(n1050), .A2(n1051), .A3(n1048), .A4(n1049), .ZN(n1044) );
OR3_X1 U752 ( .A1(n1047), .A2(KEYINPUT40), .A3(n1052), .ZN(n1050) );
NAND3_X1 U753 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1039) );
NAND3_X1 U754 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
INV_X1 U755 ( .A(n1049), .ZN(n1058) );
NAND2_X1 U756 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND3_X1 U757 ( .A1(n1029), .A2(n1061), .A3(n1062), .ZN(n1060) );
OR2_X1 U758 ( .A1(n1063), .A2(n1028), .ZN(n1061) );
NAND2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(n1059) );
NAND2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U761 ( .A1(n1062), .A2(n1068), .ZN(n1067) );
NAND2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U763 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U764 ( .A1(n1029), .A2(n1073), .ZN(n1066) );
NAND3_X1 U765 ( .A1(n1074), .A2(n1036), .A3(n1075), .ZN(n1073) );
NAND2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
INV_X1 U767 ( .A(n1078), .ZN(n1036) );
NAND2_X1 U768 ( .A1(KEYINPUT40), .A2(n1062), .ZN(n1074) );
NOR3_X1 U769 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1037) );
INV_X1 U770 ( .A(n1053), .ZN(n1079) );
NAND4_X1 U771 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1053) );
NOR4_X1 U772 ( .A1(n1076), .A2(n1084), .A3(n1085), .A4(n1072), .ZN(n1083) );
XOR2_X1 U773 ( .A(n1086), .B(G478), .Z(n1082) );
XNOR2_X1 U774 ( .A(n1087), .B(n1088), .ZN(n1081) );
XOR2_X1 U775 ( .A(n1089), .B(G472), .Z(n1080) );
XOR2_X1 U776 ( .A(n1090), .B(n1091), .Z(G72) );
XOR2_X1 U777 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR2_X1 U778 ( .A1(G953), .A2(n1094), .ZN(n1093) );
NOR2_X1 U779 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR4_X1 U780 ( .A1(KEYINPUT37), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1092) );
XOR2_X1 U781 ( .A(KEYINPUT58), .B(n1100), .Z(n1099) );
NOR2_X1 U782 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
AND2_X1 U783 ( .A1(n1102), .A2(n1101), .ZN(n1097) );
XNOR2_X1 U784 ( .A(n1103), .B(n1104), .ZN(n1101) );
XOR2_X1 U785 ( .A(n1105), .B(G137), .Z(n1103) );
NAND2_X1 U786 ( .A1(n1106), .A2(n1107), .ZN(n1102) );
NAND2_X1 U787 ( .A1(G140), .A2(n1108), .ZN(n1107) );
XOR2_X1 U788 ( .A(KEYINPUT28), .B(n1109), .Z(n1106) );
NOR2_X1 U789 ( .A1(G140), .A2(n1108), .ZN(n1109) );
NOR2_X1 U790 ( .A1(n1110), .A2(n1111), .ZN(n1090) );
AND2_X1 U791 ( .A1(G227), .A2(G900), .ZN(n1110) );
XOR2_X1 U792 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U793 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U794 ( .A1(n1116), .A2(n1111), .ZN(n1115) );
XOR2_X1 U795 ( .A(G953), .B(KEYINPUT11), .Z(n1111) );
NOR2_X1 U796 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U797 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
NAND2_X1 U798 ( .A1(n1121), .A2(n1118), .ZN(n1120) );
XOR2_X1 U799 ( .A(KEYINPUT34), .B(G953), .Z(n1121) );
XNOR2_X1 U800 ( .A(n1122), .B(n1123), .ZN(n1119) );
NAND3_X1 U801 ( .A1(n1124), .A2(n1054), .A3(KEYINPUT36), .ZN(n1112) );
NOR2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XOR2_X1 U803 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U804 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
NOR2_X1 U805 ( .A1(n1125), .A2(n1131), .ZN(G63) );
NOR3_X1 U806 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR3_X1 U807 ( .A1(n1135), .A2(n1136), .A3(n1130), .ZN(n1134) );
NOR2_X1 U808 ( .A1(n1137), .A2(n1138), .ZN(n1133) );
NOR2_X1 U809 ( .A1(n1139), .A2(n1136), .ZN(n1137) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1140), .ZN(G60) );
XOR2_X1 U811 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND3_X1 U812 ( .A1(n1143), .A2(n1041), .A3(G475), .ZN(n1141) );
XOR2_X1 U813 ( .A(KEYINPUT20), .B(G902), .Z(n1143) );
XNOR2_X1 U814 ( .A(G104), .B(n1144), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1125), .A2(n1145), .ZN(G57) );
XOR2_X1 U816 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U817 ( .A(n1148), .B(n1149), .ZN(n1147) );
XOR2_X1 U818 ( .A(n1150), .B(n1151), .Z(n1148) );
XOR2_X1 U819 ( .A(n1152), .B(n1153), .Z(n1146) );
NOR2_X1 U820 ( .A1(G101), .A2(KEYINPUT33), .ZN(n1153) );
XOR2_X1 U821 ( .A(n1154), .B(n1155), .Z(n1152) );
NOR2_X1 U822 ( .A1(n1156), .A2(n1130), .ZN(n1155) );
NOR2_X1 U823 ( .A1(n1125), .A2(n1157), .ZN(G54) );
XOR2_X1 U824 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U825 ( .A1(n1160), .A2(n1130), .ZN(n1159) );
INV_X1 U826 ( .A(G469), .ZN(n1160) );
NAND2_X1 U827 ( .A1(n1161), .A2(KEYINPUT29), .ZN(n1158) );
XNOR2_X1 U828 ( .A(n1149), .B(n1162), .ZN(n1161) );
XOR2_X1 U829 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U830 ( .A1(KEYINPUT59), .A2(n1165), .ZN(n1164) );
NOR2_X1 U831 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
NOR2_X1 U832 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NOR2_X1 U833 ( .A1(n1125), .A2(n1170), .ZN(G51) );
XOR2_X1 U834 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U835 ( .A1(n1088), .A2(n1130), .ZN(n1172) );
NAND2_X1 U836 ( .A1(G902), .A2(n1041), .ZN(n1130) );
INV_X1 U837 ( .A(n1139), .ZN(n1041) );
NOR3_X1 U838 ( .A1(n1096), .A2(n1173), .A3(n1124), .ZN(n1139) );
NAND4_X1 U839 ( .A1(n1144), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1124) );
AND4_X1 U840 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NAND2_X1 U841 ( .A1(n1028), .A2(n1181), .ZN(n1175) );
NAND2_X1 U842 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U843 ( .A1(n1032), .A2(n1029), .ZN(n1183) );
NAND2_X1 U844 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
NAND3_X1 U845 ( .A1(n1032), .A2(n1029), .A3(n1063), .ZN(n1144) );
XOR2_X1 U846 ( .A(KEYINPUT2), .B(n1095), .Z(n1173) );
NAND4_X1 U847 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1095) );
NAND4_X1 U848 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1096) );
NAND2_X1 U849 ( .A1(n1194), .A2(KEYINPUT52), .ZN(n1171) );
XOR2_X1 U850 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U851 ( .A(n1197), .B(n1198), .Z(n1196) );
NAND2_X1 U852 ( .A1(KEYINPUT9), .A2(n1199), .ZN(n1198) );
XOR2_X1 U853 ( .A(n1150), .B(n1200), .Z(n1195) );
NOR2_X1 U854 ( .A1(G125), .A2(KEYINPUT38), .ZN(n1200) );
NOR2_X1 U855 ( .A1(n1054), .A2(G952), .ZN(n1125) );
XNOR2_X1 U856 ( .A(G146), .B(n1190), .ZN(G48) );
NAND3_X1 U857 ( .A1(n1063), .A2(n1078), .A3(n1201), .ZN(n1190) );
XOR2_X1 U858 ( .A(n1191), .B(n1202), .Z(G45) );
NAND2_X1 U859 ( .A1(KEYINPUT25), .A2(G143), .ZN(n1202) );
NAND4_X1 U860 ( .A1(n1203), .A2(n1078), .A3(n1204), .A4(n1084), .ZN(n1191) );
XNOR2_X1 U861 ( .A(n1192), .B(n1205), .ZN(G42) );
XOR2_X1 U862 ( .A(KEYINPUT57), .B(G140), .Z(n1205) );
NAND3_X1 U863 ( .A1(n1062), .A2(n1206), .A3(n1207), .ZN(n1192) );
XOR2_X1 U864 ( .A(n1193), .B(n1208), .Z(G39) );
NAND2_X1 U865 ( .A1(KEYINPUT14), .A2(G137), .ZN(n1208) );
NAND3_X1 U866 ( .A1(n1062), .A2(n1064), .A3(n1201), .ZN(n1193) );
XOR2_X1 U867 ( .A(n1186), .B(n1209), .Z(G36) );
NAND2_X1 U868 ( .A1(KEYINPUT21), .A2(G134), .ZN(n1209) );
NAND3_X1 U869 ( .A1(n1062), .A2(n1028), .A3(n1203), .ZN(n1186) );
XNOR2_X1 U870 ( .A(G131), .B(n1187), .ZN(G33) );
NAND3_X1 U871 ( .A1(n1062), .A2(n1063), .A3(n1203), .ZN(n1187) );
AND3_X1 U872 ( .A1(n1206), .A2(n1210), .A3(n1184), .ZN(n1203) );
INV_X1 U873 ( .A(n1043), .ZN(n1062) );
NAND2_X1 U874 ( .A1(n1077), .A2(n1211), .ZN(n1043) );
XNOR2_X1 U875 ( .A(n1212), .B(n1188), .ZN(G30) );
NAND3_X1 U876 ( .A1(n1028), .A2(n1078), .A3(n1201), .ZN(n1188) );
AND4_X1 U877 ( .A1(n1206), .A2(n1072), .A3(n1210), .A4(n1213), .ZN(n1201) );
INV_X1 U878 ( .A(n1214), .ZN(n1028) );
XOR2_X1 U879 ( .A(n1215), .B(KEYINPUT54), .Z(n1212) );
XNOR2_X1 U880 ( .A(G101), .B(n1174), .ZN(G3) );
NAND3_X1 U881 ( .A1(n1032), .A2(n1064), .A3(n1184), .ZN(n1174) );
XOR2_X1 U882 ( .A(n1108), .B(n1189), .Z(G27) );
NAND3_X1 U883 ( .A1(n1056), .A2(n1078), .A3(n1207), .ZN(n1189) );
AND4_X1 U884 ( .A1(n1063), .A2(n1071), .A3(n1072), .A4(n1210), .ZN(n1207) );
NAND2_X1 U885 ( .A1(n1049), .A2(n1216), .ZN(n1210) );
NAND3_X1 U886 ( .A1(G902), .A2(n1217), .A3(n1098), .ZN(n1216) );
NOR2_X1 U887 ( .A1(n1054), .A2(G900), .ZN(n1098) );
XOR2_X1 U888 ( .A(n1218), .B(n1219), .Z(G24) );
NOR2_X1 U889 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NOR2_X1 U890 ( .A1(n1222), .A2(n1177), .ZN(n1221) );
NAND4_X1 U891 ( .A1(n1185), .A2(n1029), .A3(n1204), .A4(n1084), .ZN(n1177) );
INV_X1 U892 ( .A(n1223), .ZN(n1084) );
INV_X1 U893 ( .A(KEYINPUT62), .ZN(n1222) );
NOR4_X1 U894 ( .A1(KEYINPUT62), .A2(n1224), .A3(n1225), .A4(n1047), .ZN(n1220) );
INV_X1 U895 ( .A(n1029), .ZN(n1047) );
NOR2_X1 U896 ( .A1(n1213), .A2(n1072), .ZN(n1029) );
NOR2_X1 U897 ( .A1(n1223), .A2(n1226), .ZN(n1225) );
NAND2_X1 U898 ( .A1(KEYINPUT19), .A2(G122), .ZN(n1218) );
XNOR2_X1 U899 ( .A(G119), .B(n1180), .ZN(G21) );
NAND4_X1 U900 ( .A1(n1064), .A2(n1185), .A3(n1072), .A4(n1213), .ZN(n1180) );
XOR2_X1 U901 ( .A(G116), .B(n1227), .Z(G18) );
NOR4_X1 U902 ( .A1(KEYINPUT56), .A2(n1214), .A3(n1224), .A4(n1069), .ZN(n1227) );
NAND2_X1 U903 ( .A1(n1223), .A2(n1204), .ZN(n1214) );
XNOR2_X1 U904 ( .A(G113), .B(n1179), .ZN(G15) );
NAND3_X1 U905 ( .A1(n1184), .A2(n1185), .A3(n1063), .ZN(n1179) );
NOR2_X1 U906 ( .A1(n1204), .A2(n1223), .ZN(n1063) );
INV_X1 U907 ( .A(n1224), .ZN(n1185) );
NAND3_X1 U908 ( .A1(n1078), .A2(n1035), .A3(n1056), .ZN(n1224) );
INV_X1 U909 ( .A(n1085), .ZN(n1056) );
NAND2_X1 U910 ( .A1(n1228), .A2(n1051), .ZN(n1085) );
INV_X1 U911 ( .A(n1052), .ZN(n1228) );
INV_X1 U912 ( .A(n1069), .ZN(n1184) );
NAND2_X1 U913 ( .A1(n1229), .A2(n1213), .ZN(n1069) );
XNOR2_X1 U914 ( .A(n1072), .B(KEYINPUT47), .ZN(n1229) );
XNOR2_X1 U915 ( .A(G110), .B(n1178), .ZN(G12) );
NAND4_X1 U916 ( .A1(n1032), .A2(n1064), .A3(n1071), .A4(n1072), .ZN(n1178) );
XNOR2_X1 U917 ( .A(n1230), .B(n1231), .ZN(n1072) );
NOR2_X1 U918 ( .A1(n1129), .A2(n1232), .ZN(n1231) );
XNOR2_X1 U919 ( .A(KEYINPUT24), .B(n1233), .ZN(n1232) );
INV_X1 U920 ( .A(G217), .ZN(n1129) );
OR2_X1 U921 ( .A1(n1128), .A2(G902), .ZN(n1230) );
XNOR2_X1 U922 ( .A(n1234), .B(n1235), .ZN(n1128) );
XOR2_X1 U923 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND3_X1 U924 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1236) );
NAND2_X1 U925 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND2_X1 U926 ( .A1(KEYINPUT61), .A2(n1243), .ZN(n1239) );
NAND2_X1 U927 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
INV_X1 U928 ( .A(n1241), .ZN(n1245) );
XNOR2_X1 U929 ( .A(KEYINPUT18), .B(n1242), .ZN(n1244) );
NAND2_X1 U930 ( .A1(n1246), .A2(n1247), .ZN(n1238) );
INV_X1 U931 ( .A(KEYINPUT61), .ZN(n1247) );
NAND2_X1 U932 ( .A1(n1248), .A2(n1249), .ZN(n1246) );
OR3_X1 U933 ( .A1(n1242), .A2(n1241), .A3(KEYINPUT18), .ZN(n1249) );
XOR2_X1 U934 ( .A(n1250), .B(KEYINPUT12), .Z(n1241) );
NAND2_X1 U935 ( .A1(KEYINPUT18), .A2(n1242), .ZN(n1248) );
NAND3_X1 U936 ( .A1(G221), .A2(G234), .A3(n1251), .ZN(n1242) );
XOR2_X1 U937 ( .A(n1252), .B(KEYINPUT48), .Z(n1251) );
XOR2_X1 U938 ( .A(n1253), .B(n1254), .Z(n1234) );
NOR2_X1 U939 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U940 ( .A(n1257), .B(KEYINPUT30), .Z(n1256) );
NAND2_X1 U941 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NOR2_X1 U942 ( .A1(n1258), .A2(n1259), .ZN(n1255) );
XOR2_X1 U943 ( .A(KEYINPUT46), .B(G110), .Z(n1259) );
XNOR2_X1 U944 ( .A(G119), .B(n1260), .ZN(n1258) );
NOR2_X1 U945 ( .A1(G128), .A2(KEYINPUT43), .ZN(n1260) );
NAND2_X1 U946 ( .A1(KEYINPUT6), .A2(n1108), .ZN(n1253) );
INV_X1 U947 ( .A(n1213), .ZN(n1071) );
NAND3_X1 U948 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1213) );
NAND2_X1 U949 ( .A1(n1264), .A2(n1089), .ZN(n1263) );
NAND2_X1 U950 ( .A1(n1265), .A2(KEYINPUT44), .ZN(n1264) );
XOR2_X1 U951 ( .A(n1156), .B(KEYINPUT5), .Z(n1265) );
NAND3_X1 U952 ( .A1(KEYINPUT44), .A2(n1266), .A3(n1156), .ZN(n1262) );
INV_X1 U953 ( .A(n1089), .ZN(n1266) );
NAND2_X1 U954 ( .A1(n1267), .A2(n1268), .ZN(n1089) );
XOR2_X1 U955 ( .A(n1269), .B(n1270), .Z(n1267) );
XNOR2_X1 U956 ( .A(n1271), .B(n1154), .ZN(n1270) );
NAND2_X1 U957 ( .A1(G210), .A2(n1272), .ZN(n1154) );
NAND2_X1 U958 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
OR2_X1 U959 ( .A1(n1151), .A2(n1275), .ZN(n1274) );
XOR2_X1 U960 ( .A(n1276), .B(KEYINPUT23), .Z(n1273) );
NAND2_X1 U961 ( .A1(n1277), .A2(n1275), .ZN(n1276) );
XNOR2_X1 U962 ( .A(n1149), .B(n1278), .ZN(n1275) );
NOR2_X1 U963 ( .A1(KEYINPUT26), .A2(n1150), .ZN(n1278) );
XNOR2_X1 U964 ( .A(n1151), .B(KEYINPUT32), .ZN(n1277) );
XOR2_X1 U965 ( .A(n1279), .B(n1280), .Z(n1151) );
NOR2_X1 U966 ( .A1(G116), .A2(KEYINPUT50), .ZN(n1280) );
XNOR2_X1 U967 ( .A(G101), .B(KEYINPUT27), .ZN(n1269) );
OR2_X1 U968 ( .A1(n1156), .A2(KEYINPUT44), .ZN(n1261) );
INV_X1 U969 ( .A(G472), .ZN(n1156) );
INV_X1 U970 ( .A(n1048), .ZN(n1064) );
NAND2_X1 U971 ( .A1(n1223), .A2(n1226), .ZN(n1048) );
INV_X1 U972 ( .A(n1204), .ZN(n1226) );
XOR2_X1 U973 ( .A(n1281), .B(n1132), .Z(n1204) );
INV_X1 U974 ( .A(n1086), .ZN(n1132) );
NAND2_X1 U975 ( .A1(n1135), .A2(n1268), .ZN(n1086) );
INV_X1 U976 ( .A(n1138), .ZN(n1135) );
XOR2_X1 U977 ( .A(n1282), .B(n1283), .Z(n1138) );
XOR2_X1 U978 ( .A(G116), .B(n1284), .Z(n1283) );
XOR2_X1 U979 ( .A(G134), .B(G122), .Z(n1284) );
XOR2_X1 U980 ( .A(n1285), .B(n1286), .Z(n1282) );
AND3_X1 U981 ( .A1(G234), .A2(G217), .A3(n1252), .ZN(n1286) );
XOR2_X1 U982 ( .A(n1026), .B(n1287), .Z(n1285) );
NOR2_X1 U983 ( .A1(KEYINPUT13), .A2(n1288), .ZN(n1287) );
XOR2_X1 U984 ( .A(n1215), .B(G143), .Z(n1288) );
INV_X1 U985 ( .A(G128), .ZN(n1215) );
NAND2_X1 U986 ( .A1(KEYINPUT45), .A2(n1136), .ZN(n1281) );
INV_X1 U987 ( .A(G478), .ZN(n1136) );
XOR2_X1 U988 ( .A(n1289), .B(G475), .Z(n1223) );
NAND2_X1 U989 ( .A1(n1142), .A2(n1268), .ZN(n1289) );
XNOR2_X1 U990 ( .A(n1290), .B(n1291), .ZN(n1142) );
XOR2_X1 U991 ( .A(KEYINPUT0), .B(G131), .Z(n1291) );
XOR2_X1 U992 ( .A(n1292), .B(n1293), .Z(n1290) );
XOR2_X1 U993 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U994 ( .A(G125), .B(G122), .Z(n1295) );
XOR2_X1 U995 ( .A(KEYINPUT63), .B(G143), .Z(n1294) );
XOR2_X1 U996 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U997 ( .A(G113), .B(G104), .Z(n1297) );
XOR2_X1 U998 ( .A(n1298), .B(n1299), .Z(n1296) );
INV_X1 U999 ( .A(n1237), .ZN(n1299) );
XNOR2_X1 U1000 ( .A(G140), .B(G146), .ZN(n1237) );
NAND2_X1 U1001 ( .A1(G214), .A2(n1272), .ZN(n1298) );
NOR2_X1 U1002 ( .A1(n1300), .A2(G237), .ZN(n1272) );
AND3_X1 U1003 ( .A1(n1206), .A2(n1035), .A3(n1078), .ZN(n1032) );
NOR2_X1 U1004 ( .A1(n1077), .A2(n1076), .ZN(n1078) );
INV_X1 U1005 ( .A(n1211), .ZN(n1076) );
NAND2_X1 U1006 ( .A1(G214), .A2(n1301), .ZN(n1211) );
XOR2_X1 U1007 ( .A(n1302), .B(n1088), .Z(n1077) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1301), .ZN(n1088) );
NAND2_X1 U1009 ( .A1(n1303), .A2(n1268), .ZN(n1301) );
INV_X1 U1010 ( .A(G237), .ZN(n1303) );
NAND2_X1 U1011 ( .A1(KEYINPUT16), .A2(n1304), .ZN(n1302) );
XNOR2_X1 U1012 ( .A(KEYINPUT60), .B(n1087), .ZN(n1304) );
NAND2_X1 U1013 ( .A1(n1305), .A2(n1268), .ZN(n1087) );
XOR2_X1 U1014 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1015 ( .A(n1150), .B(n1308), .Z(n1307) );
XOR2_X1 U1016 ( .A(n1309), .B(n1199), .Z(n1308) );
NOR2_X1 U1017 ( .A1(n1117), .A2(n1300), .ZN(n1199) );
INV_X1 U1018 ( .A(n1252), .ZN(n1300) );
INV_X1 U1019 ( .A(G224), .ZN(n1117) );
NAND2_X1 U1020 ( .A1(KEYINPUT31), .A2(n1108), .ZN(n1309) );
INV_X1 U1021 ( .A(G125), .ZN(n1108) );
XNOR2_X1 U1022 ( .A(n1310), .B(G146), .ZN(n1150) );
XOR2_X1 U1023 ( .A(n1197), .B(n1311), .Z(n1306) );
XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(KEYINPUT4), .ZN(n1311) );
NAND2_X1 U1025 ( .A1(n1312), .A2(n1313), .ZN(n1197) );
NAND2_X1 U1026 ( .A1(n1123), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1027 ( .A(KEYINPUT41), .B(n1315), .Z(n1312) );
NOR2_X1 U1028 ( .A1(n1123), .A2(n1314), .ZN(n1315) );
NAND2_X1 U1029 ( .A1(n1316), .A2(n1317), .ZN(n1314) );
OR2_X1 U1030 ( .A1(n1122), .A2(KEYINPUT53), .ZN(n1317) );
XNOR2_X1 U1031 ( .A(n1318), .B(n1319), .ZN(n1122) );
NAND3_X1 U1032 ( .A1(n1319), .A2(n1318), .A3(KEYINPUT53), .ZN(n1316) );
XOR2_X1 U1033 ( .A(n1320), .B(n1321), .Z(n1318) );
NOR2_X1 U1034 ( .A1(KEYINPUT39), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1035 ( .A(G104), .B(n1026), .Z(n1322) );
INV_X1 U1036 ( .A(G107), .ZN(n1026) );
XNOR2_X1 U1037 ( .A(G101), .B(KEYINPUT7), .ZN(n1320) );
XOR2_X1 U1038 ( .A(G116), .B(n1279), .Z(n1319) );
XOR2_X1 U1039 ( .A(G113), .B(G119), .Z(n1279) );
XNOR2_X1 U1040 ( .A(G110), .B(G122), .ZN(n1123) );
NAND2_X1 U1041 ( .A1(n1049), .A2(n1323), .ZN(n1035) );
NAND4_X1 U1042 ( .A1(G902), .A2(G953), .A3(n1217), .A4(n1118), .ZN(n1323) );
INV_X1 U1043 ( .A(G898), .ZN(n1118) );
NAND3_X1 U1044 ( .A1(n1217), .A2(n1054), .A3(G952), .ZN(n1049) );
NAND2_X1 U1045 ( .A1(G237), .A2(G234), .ZN(n1217) );
INV_X1 U1046 ( .A(n1034), .ZN(n1206) );
NAND2_X1 U1047 ( .A1(n1052), .A2(n1051), .ZN(n1034) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1233), .ZN(n1051) );
NAND2_X1 U1049 ( .A1(G234), .A2(n1268), .ZN(n1233) );
XNOR2_X1 U1050 ( .A(n1324), .B(G469), .ZN(n1052) );
NAND2_X1 U1051 ( .A1(n1325), .A2(n1268), .ZN(n1324) );
INV_X1 U1052 ( .A(G902), .ZN(n1268) );
XOR2_X1 U1053 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1054 ( .A(KEYINPUT1), .B(n1328), .Z(n1327) );
NOR3_X1 U1055 ( .A1(n1167), .A2(n1329), .A3(n1330), .ZN(n1328) );
AND2_X1 U1056 ( .A1(n1169), .A2(KEYINPUT10), .ZN(n1330) );
NOR3_X1 U1057 ( .A1(KEYINPUT10), .A2(n1168), .A3(n1169), .ZN(n1329) );
AND2_X1 U1058 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U1059 ( .A(G110), .B(n1331), .Z(n1169) );
XOR2_X1 U1060 ( .A(KEYINPUT55), .B(G140), .Z(n1331) );
AND2_X1 U1061 ( .A1(G227), .A2(n1252), .ZN(n1168) );
XOR2_X1 U1062 ( .A(n1054), .B(KEYINPUT22), .Z(n1252) );
INV_X1 U1063 ( .A(G953), .ZN(n1054) );
XNOR2_X1 U1064 ( .A(n1165), .B(n1149), .ZN(n1326) );
NAND2_X1 U1065 ( .A1(n1332), .A2(n1333), .ZN(n1149) );
NAND2_X1 U1066 ( .A1(n1104), .A2(G137), .ZN(n1333) );
NAND2_X1 U1067 ( .A1(n1334), .A2(n1250), .ZN(n1332) );
INV_X1 U1068 ( .A(G137), .ZN(n1250) );
XNOR2_X1 U1069 ( .A(n1104), .B(KEYINPUT15), .ZN(n1334) );
XOR2_X1 U1070 ( .A(G131), .B(G134), .Z(n1104) );
XOR2_X1 U1071 ( .A(n1105), .B(n1335), .Z(n1165) );
XNOR2_X1 U1072 ( .A(G101), .B(n1336), .ZN(n1335) );
NAND2_X1 U1073 ( .A1(KEYINPUT49), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1074 ( .A(G107), .B(G104), .Z(n1337) );
XOR2_X1 U1075 ( .A(n1338), .B(n1310), .Z(n1105) );
XNOR2_X1 U1076 ( .A(n1339), .B(n1340), .ZN(n1310) );
XOR2_X1 U1077 ( .A(G143), .B(G128), .Z(n1340) );
XNOR2_X1 U1078 ( .A(KEYINPUT3), .B(KEYINPUT17), .ZN(n1339) );
NAND2_X1 U1079 ( .A1(KEYINPUT42), .A2(G146), .ZN(n1338) );
endmodule


