//Key = 0011010000101111100110100101111110011001000101101010001000101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
n1422, n1423, n1424, n1425, n1426;

XNOR2_X1 U776 ( .A(G107), .B(n1082), .ZN(G9) );
NAND3_X1 U777 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(G75) );
NOR4_X1 U779 ( .A1(n1088), .A2(n1089), .A3(G953), .A4(n1090), .ZN(n1087) );
NOR3_X1 U780 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1089) );
XOR2_X1 U781 ( .A(n1094), .B(KEYINPUT61), .Z(n1092) );
NAND3_X1 U782 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1088) );
NAND3_X1 U783 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1096) );
NAND2_X1 U784 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND3_X1 U785 ( .A1(n1084), .A2(n1103), .A3(n1104), .ZN(n1102) );
NAND2_X1 U786 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
NAND2_X1 U787 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
INV_X1 U788 ( .A(n1109), .ZN(n1105) );
NAND2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1101) );
NAND2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U791 ( .A1(n1104), .A2(n1114), .ZN(n1113) );
OR2_X1 U792 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U793 ( .A1(n1084), .A2(n1117), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XNOR2_X1 U795 ( .A(n1120), .B(KEYINPUT18), .ZN(n1118) );
NAND2_X1 U796 ( .A1(n1121), .A2(n1122), .ZN(n1095) );
XOR2_X1 U797 ( .A(n1094), .B(KEYINPUT20), .Z(n1121) );
NAND4_X1 U798 ( .A1(n1104), .A2(n1110), .A3(n1084), .A4(n1099), .ZN(n1094) );
NOR3_X1 U799 ( .A1(n1090), .A2(G953), .A3(G952), .ZN(n1086) );
AND4_X1 U800 ( .A1(n1123), .A2(n1100), .A3(n1124), .A4(n1125), .ZN(n1090) );
NOR4_X1 U801 ( .A1(n1107), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1125) );
NOR2_X1 U802 ( .A1(n1129), .A2(n1130), .ZN(n1126) );
NOR2_X1 U803 ( .A1(G902), .A2(n1131), .ZN(n1129) );
NOR2_X1 U804 ( .A1(n1132), .A2(n1133), .ZN(n1124) );
XNOR2_X1 U805 ( .A(n1134), .B(n1135), .ZN(n1133) );
XOR2_X1 U806 ( .A(KEYINPUT63), .B(n1136), .Z(n1132) );
XOR2_X1 U807 ( .A(n1137), .B(n1138), .Z(G72) );
NOR2_X1 U808 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U809 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NAND2_X1 U810 ( .A1(n1143), .A2(n1144), .ZN(n1137) );
NAND2_X1 U811 ( .A1(n1145), .A2(n1140), .ZN(n1144) );
XOR2_X1 U812 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U813 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NAND3_X1 U814 ( .A1(G900), .A2(n1147), .A3(G953), .ZN(n1143) );
XNOR2_X1 U815 ( .A(n1150), .B(n1151), .ZN(n1147) );
XOR2_X1 U816 ( .A(n1152), .B(KEYINPUT16), .Z(n1150) );
NAND2_X1 U817 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U818 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U819 ( .A(n1157), .B(KEYINPUT55), .Z(n1153) );
OR2_X1 U820 ( .A1(n1156), .A2(n1155), .ZN(n1157) );
XNOR2_X1 U821 ( .A(n1158), .B(n1159), .ZN(n1156) );
NOR2_X1 U822 ( .A1(G131), .A2(KEYINPUT52), .ZN(n1159) );
XOR2_X1 U823 ( .A(n1160), .B(G134), .Z(n1158) );
NAND2_X1 U824 ( .A1(KEYINPUT12), .A2(n1161), .ZN(n1160) );
XOR2_X1 U825 ( .A(n1162), .B(n1163), .Z(G69) );
NOR2_X1 U826 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U827 ( .A(n1166), .B(n1167), .ZN(n1165) );
NOR2_X1 U828 ( .A1(n1140), .A2(n1168), .ZN(n1164) );
XNOR2_X1 U829 ( .A(KEYINPUT6), .B(n1169), .ZN(n1168) );
NAND2_X1 U830 ( .A1(n1170), .A2(n1171), .ZN(n1162) );
NAND2_X1 U831 ( .A1(n1172), .A2(n1140), .ZN(n1171) );
NAND3_X1 U832 ( .A1(KEYINPUT25), .A2(n1173), .A3(G953), .ZN(n1170) );
NAND2_X1 U833 ( .A1(G898), .A2(G224), .ZN(n1173) );
NOR2_X1 U834 ( .A1(n1174), .A2(n1175), .ZN(G66) );
NOR3_X1 U835 ( .A1(n1134), .A2(n1176), .A3(n1177), .ZN(n1175) );
AND3_X1 U836 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
NOR2_X1 U837 ( .A1(n1181), .A2(n1178), .ZN(n1176) );
NOR2_X1 U838 ( .A1(n1097), .A2(n1135), .ZN(n1181) );
NOR2_X1 U839 ( .A1(n1174), .A2(n1182), .ZN(G63) );
NOR2_X1 U840 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
XOR2_X1 U841 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U842 ( .A1(KEYINPUT4), .A2(n1187), .ZN(n1186) );
AND2_X1 U843 ( .A1(G478), .A2(n1180), .ZN(n1185) );
AND2_X1 U844 ( .A1(n1187), .A2(KEYINPUT4), .ZN(n1183) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1188), .ZN(G60) );
XNOR2_X1 U846 ( .A(n1189), .B(n1131), .ZN(n1188) );
NAND3_X1 U847 ( .A1(n1180), .A2(n1190), .A3(KEYINPUT46), .ZN(n1189) );
XNOR2_X1 U848 ( .A(KEYINPUT26), .B(n1130), .ZN(n1190) );
INV_X1 U849 ( .A(G475), .ZN(n1130) );
XNOR2_X1 U850 ( .A(G104), .B(n1191), .ZN(G6) );
NOR2_X1 U851 ( .A1(n1174), .A2(n1192), .ZN(G57) );
XOR2_X1 U852 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U853 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(n1196) );
AND2_X1 U855 ( .A1(G472), .A2(n1180), .ZN(n1197) );
XOR2_X1 U856 ( .A(n1199), .B(n1200), .Z(n1193) );
XNOR2_X1 U857 ( .A(G101), .B(KEYINPUT28), .ZN(n1200) );
NOR2_X1 U858 ( .A1(n1174), .A2(n1201), .ZN(G54) );
NOR2_X1 U859 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XOR2_X1 U860 ( .A(n1204), .B(KEYINPUT31), .Z(n1203) );
NAND2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NOR2_X1 U862 ( .A1(n1205), .A2(n1206), .ZN(n1202) );
XNOR2_X1 U863 ( .A(n1207), .B(n1208), .ZN(n1206) );
XOR2_X1 U864 ( .A(n1209), .B(n1210), .Z(n1207) );
NAND2_X1 U865 ( .A1(KEYINPUT13), .A2(n1155), .ZN(n1209) );
AND2_X1 U866 ( .A1(n1180), .A2(G469), .ZN(n1205) );
NOR3_X1 U867 ( .A1(n1174), .A2(n1211), .A3(n1212), .ZN(G51) );
NOR2_X1 U868 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
INV_X1 U869 ( .A(n1215), .ZN(n1214) );
NOR2_X1 U870 ( .A1(n1216), .A2(n1217), .ZN(n1213) );
NOR3_X1 U871 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
AND2_X1 U872 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
INV_X1 U873 ( .A(KEYINPUT48), .ZN(n1218) );
NOR2_X1 U874 ( .A1(n1221), .A2(n1215), .ZN(n1211) );
XNOR2_X1 U875 ( .A(n1222), .B(n1223), .ZN(n1215) );
NOR2_X1 U876 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NOR2_X1 U877 ( .A1(n1219), .A2(n1220), .ZN(n1221) );
INV_X1 U878 ( .A(KEYINPUT54), .ZN(n1220) );
NAND2_X1 U879 ( .A1(n1180), .A2(G210), .ZN(n1219) );
NOR2_X1 U880 ( .A1(n1226), .A2(n1097), .ZN(n1180) );
AND3_X1 U881 ( .A1(n1227), .A2(n1228), .A3(n1148), .ZN(n1097) );
NOR3_X1 U882 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1148) );
OR4_X1 U883 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1231) );
NOR3_X1 U884 ( .A1(n1236), .A2(n1120), .A3(n1237), .ZN(n1235) );
AND2_X1 U885 ( .A1(n1236), .A2(n1238), .ZN(n1234) );
INV_X1 U886 ( .A(KEYINPUT59), .ZN(n1236) );
NOR4_X1 U887 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1233) );
NAND3_X1 U888 ( .A1(n1115), .A2(n1109), .A3(n1083), .ZN(n1240) );
INV_X1 U889 ( .A(KEYINPUT56), .ZN(n1239) );
NOR2_X1 U890 ( .A1(KEYINPUT56), .A2(n1243), .ZN(n1232) );
XOR2_X1 U891 ( .A(KEYINPUT21), .B(n1149), .Z(n1228) );
AND4_X1 U892 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1149) );
OR3_X1 U893 ( .A1(n1248), .A2(n1241), .A3(n1249), .ZN(n1245) );
INV_X1 U894 ( .A(n1172), .ZN(n1227) );
NAND4_X1 U895 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1172) );
AND4_X1 U896 ( .A1(n1191), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1253) );
NAND3_X1 U897 ( .A1(n1085), .A2(n1084), .A3(n1120), .ZN(n1191) );
NOR3_X1 U898 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1252) );
NOR2_X1 U899 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U900 ( .A(KEYINPUT5), .ZN(n1260) );
NOR4_X1 U901 ( .A1(KEYINPUT5), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1258) );
NAND3_X1 U902 ( .A1(n1265), .A2(n1266), .A3(n1115), .ZN(n1262) );
NOR3_X1 U903 ( .A1(n1267), .A2(n1119), .A3(n1268), .ZN(n1257) );
XOR2_X1 U904 ( .A(n1084), .B(KEYINPUT36), .Z(n1267) );
NOR2_X1 U905 ( .A1(n1140), .A2(G952), .ZN(n1174) );
XNOR2_X1 U906 ( .A(n1246), .B(n1269), .ZN(G48) );
NOR2_X1 U907 ( .A1(KEYINPUT17), .A2(n1270), .ZN(n1269) );
OR3_X1 U908 ( .A1(n1248), .A2(n1266), .A3(n1263), .ZN(n1246) );
XNOR2_X1 U909 ( .A(G143), .B(n1271), .ZN(G45) );
NAND2_X1 U910 ( .A1(KEYINPUT27), .A2(n1272), .ZN(n1271) );
INV_X1 U911 ( .A(n1244), .ZN(n1272) );
NAND4_X1 U912 ( .A1(n1273), .A2(n1122), .A3(n1115), .A4(n1274), .ZN(n1244) );
AND3_X1 U913 ( .A1(n1109), .A2(n1275), .A3(n1242), .ZN(n1274) );
XNOR2_X1 U914 ( .A(G140), .B(n1247), .ZN(G42) );
NAND3_X1 U915 ( .A1(n1120), .A2(n1276), .A3(n1116), .ZN(n1247) );
XNOR2_X1 U916 ( .A(n1161), .B(n1277), .ZN(G39) );
NOR4_X1 U917 ( .A1(KEYINPUT9), .A2(n1241), .A3(n1248), .A4(n1249), .ZN(n1277) );
INV_X1 U918 ( .A(n1104), .ZN(n1249) );
INV_X1 U919 ( .A(n1100), .ZN(n1241) );
XOR2_X1 U920 ( .A(n1243), .B(n1278), .Z(G36) );
XOR2_X1 U921 ( .A(KEYINPUT32), .B(G134), .Z(n1278) );
NAND3_X1 U922 ( .A1(n1083), .A2(n1115), .A3(n1276), .ZN(n1243) );
XOR2_X1 U923 ( .A(n1279), .B(n1229), .Z(G33) );
AND3_X1 U924 ( .A1(n1276), .A2(n1115), .A3(n1120), .ZN(n1229) );
AND3_X1 U925 ( .A1(n1109), .A2(n1242), .A3(n1100), .ZN(n1276) );
NOR2_X1 U926 ( .A1(n1093), .A2(n1280), .ZN(n1100) );
INV_X1 U927 ( .A(n1091), .ZN(n1280) );
NAND2_X1 U928 ( .A1(KEYINPUT30), .A2(n1281), .ZN(n1279) );
XOR2_X1 U929 ( .A(G128), .B(n1230), .Z(G30) );
NOR3_X1 U930 ( .A1(n1119), .A2(n1266), .A3(n1248), .ZN(n1230) );
NAND4_X1 U931 ( .A1(n1282), .A2(n1109), .A3(n1283), .A4(n1242), .ZN(n1248) );
XNOR2_X1 U932 ( .A(G101), .B(n1250), .ZN(G3) );
NAND3_X1 U933 ( .A1(n1085), .A2(n1115), .A3(n1104), .ZN(n1250) );
XOR2_X1 U934 ( .A(G125), .B(n1238), .Z(G27) );
NOR2_X1 U935 ( .A1(n1237), .A2(n1263), .ZN(n1238) );
INV_X1 U936 ( .A(n1120), .ZN(n1263) );
NAND4_X1 U937 ( .A1(n1110), .A2(n1116), .A3(n1122), .A4(n1242), .ZN(n1237) );
NAND2_X1 U938 ( .A1(n1284), .A2(n1285), .ZN(n1242) );
NAND2_X1 U939 ( .A1(n1286), .A2(n1142), .ZN(n1285) );
INV_X1 U940 ( .A(G900), .ZN(n1142) );
XNOR2_X1 U941 ( .A(G122), .B(n1251), .ZN(G24) );
NAND4_X1 U942 ( .A1(n1273), .A2(n1287), .A3(n1084), .A4(n1275), .ZN(n1251) );
NAND2_X1 U943 ( .A1(n1288), .A2(n1289), .ZN(n1084) );
OR3_X1 U944 ( .A1(n1282), .A2(n1283), .A3(KEYINPUT7), .ZN(n1289) );
NAND2_X1 U945 ( .A1(KEYINPUT7), .A2(n1115), .ZN(n1288) );
XNOR2_X1 U946 ( .A(G119), .B(n1256), .ZN(G21) );
NAND4_X1 U947 ( .A1(n1287), .A2(n1104), .A3(n1282), .A4(n1283), .ZN(n1256) );
NAND2_X1 U948 ( .A1(n1290), .A2(n1291), .ZN(G18) );
NAND2_X1 U949 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U950 ( .A(n1255), .B(KEYINPUT50), .Z(n1292) );
NAND2_X1 U951 ( .A1(G116), .A2(n1294), .ZN(n1290) );
XOR2_X1 U952 ( .A(n1255), .B(KEYINPUT23), .Z(n1294) );
NAND3_X1 U953 ( .A1(n1083), .A2(n1115), .A3(n1287), .ZN(n1255) );
INV_X1 U954 ( .A(n1119), .ZN(n1083) );
NAND2_X1 U955 ( .A1(n1295), .A2(n1273), .ZN(n1119) );
XNOR2_X1 U956 ( .A(G113), .B(n1261), .ZN(G15) );
NAND3_X1 U957 ( .A1(n1120), .A2(n1115), .A3(n1287), .ZN(n1261) );
AND3_X1 U958 ( .A1(n1122), .A2(n1265), .A3(n1110), .ZN(n1287) );
INV_X1 U959 ( .A(n1264), .ZN(n1110) );
NAND2_X1 U960 ( .A1(n1108), .A2(n1296), .ZN(n1264) );
NOR2_X1 U961 ( .A1(n1282), .A2(n1297), .ZN(n1115) );
INV_X1 U962 ( .A(n1283), .ZN(n1297) );
NOR2_X1 U963 ( .A1(n1273), .A2(n1295), .ZN(n1120) );
XNOR2_X1 U964 ( .A(G110), .B(n1254), .ZN(G12) );
NAND3_X1 U965 ( .A1(n1116), .A2(n1085), .A3(n1104), .ZN(n1254) );
NOR2_X1 U966 ( .A1(n1275), .A2(n1273), .ZN(n1104) );
XNOR2_X1 U967 ( .A(n1127), .B(KEYINPUT2), .ZN(n1273) );
XNOR2_X1 U968 ( .A(n1298), .B(G478), .ZN(n1127) );
OR2_X1 U969 ( .A1(n1187), .A2(G902), .ZN(n1298) );
XNOR2_X1 U970 ( .A(n1299), .B(n1300), .ZN(n1187) );
XOR2_X1 U971 ( .A(n1301), .B(n1302), .Z(n1300) );
AND2_X1 U972 ( .A1(n1303), .A2(G217), .ZN(n1302) );
NOR2_X1 U973 ( .A1(KEYINPUT57), .A2(n1304), .ZN(n1301) );
XNOR2_X1 U974 ( .A(G134), .B(n1305), .ZN(n1304) );
NOR2_X1 U975 ( .A1(KEYINPUT1), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U976 ( .A(n1307), .B(G128), .ZN(n1306) );
XNOR2_X1 U977 ( .A(G107), .B(n1308), .ZN(n1299) );
XNOR2_X1 U978 ( .A(n1309), .B(G116), .ZN(n1308) );
INV_X1 U979 ( .A(n1295), .ZN(n1275) );
NOR2_X1 U980 ( .A1(n1310), .A2(n1136), .ZN(n1295) );
NOR3_X1 U981 ( .A1(G475), .A2(G902), .A3(n1131), .ZN(n1136) );
AND2_X1 U982 ( .A1(G475), .A2(n1311), .ZN(n1310) );
NAND2_X1 U983 ( .A1(n1312), .A2(n1226), .ZN(n1311) );
INV_X1 U984 ( .A(n1131), .ZN(n1312) );
XNOR2_X1 U985 ( .A(n1313), .B(n1314), .ZN(n1131) );
XOR2_X1 U986 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U987 ( .A(G113), .B(n1317), .ZN(n1316) );
XNOR2_X1 U988 ( .A(n1307), .B(G131), .ZN(n1315) );
XOR2_X1 U989 ( .A(n1318), .B(n1319), .Z(n1313) );
NOR2_X1 U990 ( .A1(KEYINPUT37), .A2(n1309), .ZN(n1319) );
XOR2_X1 U991 ( .A(n1320), .B(n1321), .Z(n1318) );
NOR2_X1 U992 ( .A1(n1322), .A2(KEYINPUT49), .ZN(n1321) );
NOR2_X1 U993 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U994 ( .A(n1325), .B(KEYINPUT58), .Z(n1324) );
NAND2_X1 U995 ( .A1(n1326), .A2(n1270), .ZN(n1325) );
NOR2_X1 U996 ( .A1(n1326), .A2(n1270), .ZN(n1323) );
NAND2_X1 U997 ( .A1(n1327), .A2(G214), .ZN(n1320) );
INV_X1 U998 ( .A(n1268), .ZN(n1085) );
NAND3_X1 U999 ( .A1(n1109), .A2(n1265), .A3(n1122), .ZN(n1268) );
INV_X1 U1000 ( .A(n1266), .ZN(n1122) );
NAND2_X1 U1001 ( .A1(n1093), .A2(n1091), .ZN(n1266) );
NAND2_X1 U1002 ( .A1(G214), .A2(n1328), .ZN(n1091) );
NAND2_X1 U1003 ( .A1(n1226), .A2(n1329), .ZN(n1328) );
NAND2_X1 U1004 ( .A1(n1330), .A2(n1331), .ZN(n1093) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1332), .ZN(n1331) );
NAND2_X1 U1006 ( .A1(n1226), .A2(n1333), .ZN(n1332) );
OR2_X1 U1007 ( .A1(n1329), .A2(n1334), .ZN(n1333) );
INV_X1 U1008 ( .A(G237), .ZN(n1329) );
NAND3_X1 U1009 ( .A1(n1335), .A2(n1226), .A3(n1334), .ZN(n1330) );
XNOR2_X1 U1010 ( .A(n1222), .B(n1336), .ZN(n1334) );
NOR2_X1 U1011 ( .A1(n1225), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1012 ( .A(n1224), .B(KEYINPUT3), .ZN(n1337) );
NOR3_X1 U1013 ( .A1(n1338), .A2(G953), .A3(n1339), .ZN(n1224) );
INV_X1 U1014 ( .A(G224), .ZN(n1338) );
AND2_X1 U1015 ( .A1(n1339), .A2(n1340), .ZN(n1225) );
NAND2_X1 U1016 ( .A1(G224), .A2(n1140), .ZN(n1340) );
XNOR2_X1 U1017 ( .A(n1341), .B(G125), .ZN(n1339) );
NAND3_X1 U1018 ( .A1(n1342), .A2(n1343), .A3(n1344), .ZN(n1222) );
NAND2_X1 U1019 ( .A1(n1167), .A2(n1166), .ZN(n1344) );
NAND2_X1 U1020 ( .A1(n1345), .A2(n1346), .ZN(n1343) );
INV_X1 U1021 ( .A(KEYINPUT29), .ZN(n1346) );
NAND2_X1 U1022 ( .A1(n1347), .A2(n1348), .ZN(n1345) );
INV_X1 U1023 ( .A(n1166), .ZN(n1348) );
XNOR2_X1 U1024 ( .A(n1167), .B(KEYINPUT41), .ZN(n1347) );
NAND2_X1 U1025 ( .A1(KEYINPUT29), .A2(n1349), .ZN(n1342) );
NAND2_X1 U1026 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
OR3_X1 U1027 ( .A1(n1166), .A2(n1167), .A3(KEYINPUT41), .ZN(n1351) );
XNOR2_X1 U1028 ( .A(n1352), .B(n1353), .ZN(n1166) );
XOR2_X1 U1029 ( .A(n1354), .B(n1355), .Z(n1353) );
NOR2_X1 U1030 ( .A1(G104), .A2(KEYINPUT24), .ZN(n1354) );
XOR2_X1 U1031 ( .A(n1356), .B(n1357), .Z(n1352) );
XOR2_X1 U1032 ( .A(KEYINPUT33), .B(G113), .Z(n1357) );
NAND3_X1 U1033 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1356) );
NAND2_X1 U1034 ( .A1(KEYINPUT11), .A2(G119), .ZN(n1360) );
NAND3_X1 U1035 ( .A1(n1361), .A2(n1362), .A3(G116), .ZN(n1359) );
NAND2_X1 U1036 ( .A1(n1363), .A2(n1293), .ZN(n1358) );
INV_X1 U1037 ( .A(G116), .ZN(n1293) );
NAND2_X1 U1038 ( .A1(n1364), .A2(n1362), .ZN(n1363) );
INV_X1 U1039 ( .A(KEYINPUT11), .ZN(n1362) );
XNOR2_X1 U1040 ( .A(G119), .B(KEYINPUT51), .ZN(n1364) );
NAND2_X1 U1041 ( .A1(KEYINPUT41), .A2(n1167), .ZN(n1350) );
AND3_X1 U1042 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1167) );
NAND2_X1 U1043 ( .A1(n1368), .A2(n1309), .ZN(n1367) );
NAND2_X1 U1044 ( .A1(KEYINPUT53), .A2(n1369), .ZN(n1366) );
NAND2_X1 U1045 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
XNOR2_X1 U1046 ( .A(KEYINPUT44), .B(n1309), .ZN(n1371) );
INV_X1 U1047 ( .A(n1368), .ZN(n1370) );
NAND2_X1 U1048 ( .A1(n1372), .A2(n1373), .ZN(n1365) );
INV_X1 U1049 ( .A(KEYINPUT53), .ZN(n1373) );
NAND2_X1 U1050 ( .A1(n1374), .A2(n1375), .ZN(n1372) );
OR3_X1 U1051 ( .A1(n1309), .A2(n1368), .A3(KEYINPUT44), .ZN(n1375) );
NAND2_X1 U1052 ( .A1(KEYINPUT44), .A2(n1309), .ZN(n1374) );
INV_X1 U1053 ( .A(G122), .ZN(n1309) );
NAND2_X1 U1054 ( .A1(G210), .A2(G237), .ZN(n1335) );
NAND2_X1 U1055 ( .A1(n1284), .A2(n1376), .ZN(n1265) );
NAND2_X1 U1056 ( .A1(n1286), .A2(n1169), .ZN(n1376) );
INV_X1 U1057 ( .A(G898), .ZN(n1169) );
AND3_X1 U1058 ( .A1(G902), .A2(n1099), .A3(G953), .ZN(n1286) );
NAND3_X1 U1059 ( .A1(G952), .A2(n1099), .A3(n1377), .ZN(n1284) );
XNOR2_X1 U1060 ( .A(G953), .B(KEYINPUT47), .ZN(n1377) );
NAND2_X1 U1061 ( .A1(G234), .A2(G237), .ZN(n1099) );
NOR2_X1 U1062 ( .A1(n1108), .A2(n1107), .ZN(n1109) );
INV_X1 U1063 ( .A(n1296), .ZN(n1107) );
NAND2_X1 U1064 ( .A1(G221), .A2(n1378), .ZN(n1296) );
XOR2_X1 U1065 ( .A(n1128), .B(KEYINPUT19), .Z(n1108) );
XNOR2_X1 U1066 ( .A(n1379), .B(G469), .ZN(n1128) );
NAND2_X1 U1067 ( .A1(n1380), .A2(n1226), .ZN(n1379) );
XNOR2_X1 U1068 ( .A(n1210), .B(n1381), .ZN(n1380) );
XNOR2_X1 U1069 ( .A(n1155), .B(n1382), .ZN(n1381) );
NAND2_X1 U1070 ( .A1(KEYINPUT45), .A2(n1208), .ZN(n1382) );
XNOR2_X1 U1071 ( .A(n1383), .B(n1355), .ZN(n1208) );
XNOR2_X1 U1072 ( .A(n1384), .B(G101), .ZN(n1355) );
INV_X1 U1073 ( .A(G107), .ZN(n1384) );
NAND2_X1 U1074 ( .A1(n1385), .A2(n1317), .ZN(n1383) );
INV_X1 U1075 ( .A(G104), .ZN(n1317) );
XOR2_X1 U1076 ( .A(KEYINPUT62), .B(KEYINPUT43), .Z(n1385) );
AND3_X1 U1077 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n1155) );
XNOR2_X1 U1078 ( .A(n1389), .B(n1390), .ZN(n1210) );
XOR2_X1 U1079 ( .A(G140), .B(n1391), .Z(n1390) );
NOR2_X1 U1080 ( .A1(G953), .A2(n1141), .ZN(n1391) );
INV_X1 U1081 ( .A(G227), .ZN(n1141) );
XNOR2_X1 U1082 ( .A(n1198), .B(n1368), .ZN(n1389) );
AND2_X1 U1083 ( .A1(n1392), .A2(n1282), .ZN(n1116) );
XNOR2_X1 U1084 ( .A(n1134), .B(n1393), .ZN(n1282) );
NOR2_X1 U1085 ( .A1(n1179), .A2(KEYINPUT8), .ZN(n1393) );
INV_X1 U1086 ( .A(n1135), .ZN(n1179) );
NAND2_X1 U1087 ( .A1(G217), .A2(n1378), .ZN(n1135) );
NAND2_X1 U1088 ( .A1(G234), .A2(n1226), .ZN(n1378) );
NOR2_X1 U1089 ( .A1(n1178), .A2(G902), .ZN(n1134) );
XNOR2_X1 U1090 ( .A(n1394), .B(n1395), .ZN(n1178) );
NOR2_X1 U1091 ( .A1(KEYINPUT34), .A2(n1396), .ZN(n1395) );
XNOR2_X1 U1092 ( .A(n1397), .B(n1161), .ZN(n1396) );
NAND2_X1 U1093 ( .A1(n1303), .A2(G221), .ZN(n1397) );
AND2_X1 U1094 ( .A1(G234), .A2(n1140), .ZN(n1303) );
INV_X1 U1095 ( .A(G953), .ZN(n1140) );
NAND2_X1 U1096 ( .A1(n1398), .A2(n1399), .ZN(n1394) );
NAND2_X1 U1097 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
XOR2_X1 U1098 ( .A(KEYINPUT14), .B(n1402), .Z(n1398) );
NOR2_X1 U1099 ( .A1(n1400), .A2(n1401), .ZN(n1402) );
XNOR2_X1 U1100 ( .A(n1403), .B(n1368), .ZN(n1401) );
XOR2_X1 U1101 ( .A(G110), .B(KEYINPUT38), .Z(n1368) );
XNOR2_X1 U1102 ( .A(G128), .B(G119), .ZN(n1403) );
XNOR2_X1 U1103 ( .A(G146), .B(n1151), .ZN(n1400) );
INV_X1 U1104 ( .A(n1326), .ZN(n1151) );
XNOR2_X1 U1105 ( .A(G125), .B(G140), .ZN(n1326) );
XNOR2_X1 U1106 ( .A(KEYINPUT7), .B(n1283), .ZN(n1392) );
XNOR2_X1 U1107 ( .A(n1123), .B(KEYINPUT42), .ZN(n1283) );
XOR2_X1 U1108 ( .A(n1404), .B(n1405), .Z(n1123) );
XOR2_X1 U1109 ( .A(KEYINPUT0), .B(G472), .Z(n1405) );
NAND2_X1 U1110 ( .A1(n1406), .A2(n1226), .ZN(n1404) );
INV_X1 U1111 ( .A(G902), .ZN(n1226) );
XOR2_X1 U1112 ( .A(n1407), .B(n1408), .Z(n1406) );
XOR2_X1 U1113 ( .A(n1409), .B(n1410), .Z(n1408) );
XOR2_X1 U1114 ( .A(n1199), .B(KEYINPUT40), .Z(n1410) );
NAND2_X1 U1115 ( .A1(n1327), .A2(G210), .ZN(n1199) );
NOR2_X1 U1116 ( .A1(G953), .A2(G237), .ZN(n1327) );
NAND2_X1 U1117 ( .A1(KEYINPUT22), .A2(n1198), .ZN(n1409) );
XNOR2_X1 U1118 ( .A(n1411), .B(n1412), .ZN(n1198) );
XOR2_X1 U1119 ( .A(KEYINPUT10), .B(G134), .Z(n1412) );
XNOR2_X1 U1120 ( .A(n1413), .B(n1281), .ZN(n1411) );
INV_X1 U1121 ( .A(G131), .ZN(n1281) );
NAND2_X1 U1122 ( .A1(KEYINPUT39), .A2(n1161), .ZN(n1413) );
INV_X1 U1123 ( .A(G137), .ZN(n1161) );
XOR2_X1 U1124 ( .A(n1414), .B(n1195), .Z(n1407) );
XNOR2_X1 U1125 ( .A(n1415), .B(n1416), .ZN(n1195) );
XNOR2_X1 U1126 ( .A(n1361), .B(G116), .ZN(n1416) );
INV_X1 U1127 ( .A(G119), .ZN(n1361) );
XOR2_X1 U1128 ( .A(n1341), .B(G113), .Z(n1415) );
NAND3_X1 U1129 ( .A1(n1417), .A2(n1418), .A3(n1387), .ZN(n1341) );
NAND3_X1 U1130 ( .A1(n1419), .A2(n1270), .A3(G143), .ZN(n1387) );
NAND2_X1 U1131 ( .A1(KEYINPUT15), .A2(n1420), .ZN(n1418) );
NAND2_X1 U1132 ( .A1(n1386), .A2(n1388), .ZN(n1420) );
NAND3_X1 U1133 ( .A1(n1307), .A2(n1270), .A3(n1421), .ZN(n1388) );
INV_X1 U1134 ( .A(G146), .ZN(n1270) );
NAND2_X1 U1135 ( .A1(n1422), .A2(G146), .ZN(n1386) );
XNOR2_X1 U1136 ( .A(G143), .B(n1421), .ZN(n1422) );
NAND2_X1 U1137 ( .A1(n1423), .A2(n1424), .ZN(n1417) );
INV_X1 U1138 ( .A(KEYINPUT15), .ZN(n1424) );
XNOR2_X1 U1139 ( .A(n1425), .B(n1419), .ZN(n1423) );
INV_X1 U1140 ( .A(n1421), .ZN(n1419) );
XOR2_X1 U1141 ( .A(G128), .B(KEYINPUT60), .Z(n1421) );
NAND2_X1 U1142 ( .A1(G146), .A2(n1307), .ZN(n1425) );
INV_X1 U1143 ( .A(G143), .ZN(n1307) );
NAND2_X1 U1144 ( .A1(KEYINPUT35), .A2(n1426), .ZN(n1414) );
INV_X1 U1145 ( .A(G101), .ZN(n1426) );
endmodule


