//Key = 0011100011101100010100110001110111001011111000010011110001000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413;

XNOR2_X1 U771 ( .A(G107), .B(n1072), .ZN(G9) );
NAND3_X1 U772 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
XNOR2_X1 U773 ( .A(n1076), .B(KEYINPUT33), .ZN(n1075) );
NOR2_X1 U774 ( .A1(n1077), .A2(n1078), .ZN(G75) );
NOR4_X1 U775 ( .A1(G953), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1078) );
NOR2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR3_X1 U778 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U780 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NOR2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NOR2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR2_X1 U785 ( .A1(n1101), .A2(n1102), .ZN(n1093) );
NOR2_X1 U786 ( .A1(n1076), .A2(n1103), .ZN(n1101) );
NOR3_X1 U787 ( .A1(n1102), .A2(n1104), .A3(n1096), .ZN(n1089) );
NOR4_X1 U788 ( .A1(n1105), .A2(n1096), .A3(n1092), .A4(n1102), .ZN(n1084) );
INV_X1 U789 ( .A(n1106), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1086), .ZN(n1107) );
NOR3_X1 U792 ( .A1(n1087), .A2(n1109), .A3(n1110), .ZN(n1104) );
NOR3_X1 U793 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1077) );
AND4_X1 U794 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1079) );
NOR4_X1 U795 ( .A1(n1115), .A2(n1087), .A3(n1116), .A4(n1117), .ZN(n1114) );
INV_X1 U796 ( .A(n1118), .ZN(n1117) );
NOR2_X1 U797 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
XOR2_X1 U798 ( .A(n1121), .B(KEYINPUT48), .Z(n1120) );
INV_X1 U799 ( .A(n1122), .ZN(n1087) );
NOR2_X1 U800 ( .A1(n1102), .A2(n1123), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U802 ( .A(n1126), .B(KEYINPUT58), .Z(n1125) );
NAND2_X1 U803 ( .A1(KEYINPUT52), .A2(n1127), .ZN(n1124) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1112) );
XNOR2_X1 U805 ( .A(n1130), .B(G475), .ZN(n1111) );
XOR2_X1 U806 ( .A(n1131), .B(n1132), .Z(G72) );
NOR2_X1 U807 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
AND2_X1 U808 ( .A1(G227), .A2(G900), .ZN(n1133) );
NAND2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(n1131) );
NAND2_X1 U810 ( .A1(n1137), .A2(n1134), .ZN(n1136) );
XNOR2_X1 U811 ( .A(n1138), .B(n1139), .ZN(n1137) );
NAND3_X1 U812 ( .A1(n1138), .A2(G900), .A3(G953), .ZN(n1135) );
NOR2_X1 U813 ( .A1(KEYINPUT14), .A2(n1140), .ZN(n1138) );
XOR2_X1 U814 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U815 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U816 ( .A(G140), .B(G131), .Z(n1144) );
NOR2_X1 U817 ( .A1(G137), .A2(KEYINPUT45), .ZN(n1143) );
XOR2_X1 U818 ( .A(n1145), .B(n1146), .Z(n1141) );
XOR2_X1 U819 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U820 ( .A1(KEYINPUT56), .A2(n1149), .ZN(n1147) );
XOR2_X1 U821 ( .A(n1150), .B(n1151), .Z(G69) );
XOR2_X1 U822 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U823 ( .A1(KEYINPUT27), .A2(n1154), .ZN(n1153) );
NAND2_X1 U824 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U825 ( .A(KEYINPUT62), .B(n1157), .Z(n1156) );
NOR2_X1 U826 ( .A1(G898), .A2(n1134), .ZN(n1157) );
XOR2_X1 U827 ( .A(n1158), .B(n1159), .Z(n1155) );
NAND2_X1 U828 ( .A1(KEYINPUT9), .A2(n1160), .ZN(n1158) );
NAND2_X1 U829 ( .A1(n1134), .A2(n1161), .ZN(n1152) );
NAND2_X1 U830 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U831 ( .A1(G953), .A2(n1164), .ZN(n1150) );
NAND2_X1 U832 ( .A1(G898), .A2(G224), .ZN(n1164) );
NOR2_X1 U833 ( .A1(n1165), .A2(n1166), .ZN(G66) );
XNOR2_X1 U834 ( .A(n1167), .B(n1168), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1171), .ZN(G63) );
XOR2_X1 U837 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U838 ( .A(KEYINPUT15), .B(n1174), .Z(n1173) );
NOR2_X1 U839 ( .A1(n1129), .A2(n1170), .ZN(n1174) );
NOR2_X1 U840 ( .A1(n1165), .A2(n1175), .ZN(G60) );
NOR3_X1 U841 ( .A1(n1130), .A2(n1176), .A3(n1177), .ZN(n1175) );
AND3_X1 U842 ( .A1(n1178), .A2(G475), .A3(n1179), .ZN(n1177) );
NOR2_X1 U843 ( .A1(n1180), .A2(n1178), .ZN(n1176) );
AND2_X1 U844 ( .A1(n1081), .A2(G475), .ZN(n1180) );
XOR2_X1 U845 ( .A(G104), .B(n1181), .Z(G6) );
NOR2_X1 U846 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U847 ( .A1(n1165), .A2(n1184), .ZN(G57) );
XOR2_X1 U848 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U849 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR3_X1 U850 ( .A1(n1170), .A2(KEYINPUT54), .A3(n1121), .ZN(n1188) );
NOR2_X1 U851 ( .A1(n1165), .A2(n1189), .ZN(G54) );
XOR2_X1 U852 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U853 ( .A1(KEYINPUT59), .A2(n1192), .ZN(n1191) );
XOR2_X1 U854 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U855 ( .A(n1195), .B(G110), .Z(n1194) );
NAND2_X1 U856 ( .A1(KEYINPUT2), .A2(n1196), .ZN(n1195) );
NAND2_X1 U857 ( .A1(n1179), .A2(G469), .ZN(n1190) );
NOR3_X1 U858 ( .A1(n1165), .A2(n1197), .A3(n1198), .ZN(G51) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NOR2_X1 U860 ( .A1(n1201), .A2(n1202), .ZN(n1199) );
NOR2_X1 U861 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NOR2_X1 U862 ( .A1(n1205), .A2(n1206), .ZN(n1201) );
NOR2_X1 U863 ( .A1(n1207), .A2(n1208), .ZN(n1197) );
NOR2_X1 U864 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NOR2_X1 U865 ( .A1(n1204), .A2(n1206), .ZN(n1210) );
XNOR2_X1 U866 ( .A(KEYINPUT13), .B(n1211), .ZN(n1206) );
NOR2_X1 U867 ( .A1(n1205), .A2(n1203), .ZN(n1209) );
XOR2_X1 U868 ( .A(KEYINPUT39), .B(n1211), .Z(n1203) );
AND2_X1 U869 ( .A1(n1179), .A2(n1127), .ZN(n1211) );
INV_X1 U870 ( .A(n1170), .ZN(n1179) );
NAND2_X1 U871 ( .A1(G902), .A2(n1081), .ZN(n1170) );
NAND3_X1 U872 ( .A1(n1162), .A2(n1212), .A3(n1139), .ZN(n1081) );
AND4_X1 U873 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1139) );
NOR4_X1 U874 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
INV_X1 U875 ( .A(n1221), .ZN(n1220) );
NOR2_X1 U876 ( .A1(n1222), .A2(n1223), .ZN(n1215) );
NAND2_X1 U877 ( .A1(n1108), .A2(n1224), .ZN(n1214) );
NAND2_X1 U878 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND4_X1 U879 ( .A1(n1227), .A2(n1076), .A3(n1228), .A4(n1229), .ZN(n1226) );
NOR2_X1 U880 ( .A1(KEYINPUT41), .A2(n1098), .ZN(n1228) );
XOR2_X1 U881 ( .A(n1230), .B(KEYINPUT37), .Z(n1225) );
NAND2_X1 U882 ( .A1(KEYINPUT41), .A2(n1231), .ZN(n1213) );
XNOR2_X1 U883 ( .A(KEYINPUT12), .B(n1163), .ZN(n1212) );
NAND2_X1 U884 ( .A1(n1232), .A2(n1108), .ZN(n1163) );
XOR2_X1 U885 ( .A(n1183), .B(KEYINPUT29), .Z(n1232) );
NAND3_X1 U886 ( .A1(n1074), .A2(n1233), .A3(n1103), .ZN(n1183) );
AND4_X1 U887 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1162) );
NOR4_X1 U888 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1237) );
INV_X1 U889 ( .A(n1242), .ZN(n1241) );
NAND3_X1 U890 ( .A1(n1074), .A2(n1076), .A3(n1073), .ZN(n1236) );
NAND4_X1 U891 ( .A1(n1243), .A2(n1244), .A3(n1103), .A4(n1110), .ZN(n1234) );
XOR2_X1 U892 ( .A(n1182), .B(KEYINPUT31), .Z(n1243) );
INV_X1 U893 ( .A(n1204), .ZN(n1205) );
XNOR2_X1 U894 ( .A(n1245), .B(n1246), .ZN(n1204) );
NOR2_X1 U895 ( .A1(KEYINPUT0), .A2(n1247), .ZN(n1246) );
NOR2_X1 U896 ( .A1(n1134), .A2(G952), .ZN(n1165) );
XOR2_X1 U897 ( .A(G146), .B(n1223), .Z(G48) );
AND2_X1 U898 ( .A1(n1248), .A2(n1103), .ZN(n1223) );
XOR2_X1 U899 ( .A(G143), .B(n1249), .Z(G45) );
NOR2_X1 U900 ( .A1(n1182), .A2(n1230), .ZN(n1249) );
NAND4_X1 U901 ( .A1(n1110), .A2(n1229), .A3(n1098), .A4(n1250), .ZN(n1230) );
AND2_X1 U902 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U903 ( .A1(n1253), .A2(n1254), .ZN(G42) );
NAND2_X1 U904 ( .A1(G140), .A2(n1255), .ZN(n1254) );
XOR2_X1 U905 ( .A(n1256), .B(KEYINPUT7), .Z(n1253) );
NAND2_X1 U906 ( .A1(n1222), .A2(n1196), .ZN(n1256) );
INV_X1 U907 ( .A(n1255), .ZN(n1222) );
NAND3_X1 U908 ( .A1(n1103), .A2(n1257), .A3(n1109), .ZN(n1255) );
XOR2_X1 U909 ( .A(G137), .B(n1219), .Z(G39) );
AND3_X1 U910 ( .A1(n1257), .A2(n1106), .A3(n1227), .ZN(n1219) );
XOR2_X1 U911 ( .A(G134), .B(n1218), .Z(G36) );
AND3_X1 U912 ( .A1(n1076), .A2(n1110), .A3(n1257), .ZN(n1218) );
XOR2_X1 U913 ( .A(G131), .B(n1217), .Z(G33) );
AND3_X1 U914 ( .A1(n1257), .A2(n1110), .A3(n1103), .ZN(n1217) );
AND4_X1 U915 ( .A1(n1098), .A2(n1258), .A3(n1229), .A4(n1122), .ZN(n1257) );
INV_X1 U916 ( .A(n1086), .ZN(n1258) );
XOR2_X1 U917 ( .A(G128), .B(n1231), .Z(G30) );
AND2_X1 U918 ( .A1(n1248), .A2(n1076), .ZN(n1231) );
AND4_X1 U919 ( .A1(n1227), .A2(n1108), .A3(n1098), .A4(n1229), .ZN(n1248) );
XOR2_X1 U920 ( .A(n1259), .B(n1235), .Z(G3) );
NAND3_X1 U921 ( .A1(n1106), .A2(n1110), .A3(n1073), .ZN(n1235) );
XOR2_X1 U922 ( .A(n1149), .B(n1221), .Z(G27) );
NAND4_X1 U923 ( .A1(n1109), .A2(n1103), .A3(n1260), .A4(n1261), .ZN(n1221) );
AND2_X1 U924 ( .A1(n1229), .A2(n1108), .ZN(n1260) );
NAND2_X1 U925 ( .A1(n1083), .A2(n1262), .ZN(n1229) );
NAND2_X1 U926 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
INV_X1 U927 ( .A(G900), .ZN(n1264) );
NAND2_X1 U928 ( .A1(n1265), .A2(n1266), .ZN(G24) );
NAND2_X1 U929 ( .A1(G122), .A2(n1242), .ZN(n1266) );
XOR2_X1 U930 ( .A(KEYINPUT38), .B(n1267), .Z(n1265) );
NOR2_X1 U931 ( .A1(G122), .A2(n1242), .ZN(n1267) );
NAND4_X1 U932 ( .A1(n1268), .A2(n1074), .A3(n1252), .A4(n1251), .ZN(n1242) );
INV_X1 U933 ( .A(n1092), .ZN(n1074) );
NAND3_X1 U934 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(G21) );
NAND2_X1 U935 ( .A1(n1240), .A2(n1272), .ZN(n1271) );
NAND2_X1 U936 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U937 ( .A(KEYINPUT44), .B(G119), .Z(n1273) );
INV_X1 U938 ( .A(n1275), .ZN(n1240) );
NAND3_X1 U939 ( .A1(G119), .A2(n1275), .A3(n1274), .ZN(n1270) );
INV_X1 U940 ( .A(KEYINPUT11), .ZN(n1274) );
NAND3_X1 U941 ( .A1(n1227), .A2(n1106), .A3(n1268), .ZN(n1275) );
NOR2_X1 U942 ( .A1(n1118), .A2(n1276), .ZN(n1227) );
NAND2_X1 U943 ( .A1(KEYINPUT11), .A2(n1277), .ZN(n1269) );
XOR2_X1 U944 ( .A(G116), .B(n1239), .Z(G18) );
AND3_X1 U945 ( .A1(n1076), .A2(n1110), .A3(n1268), .ZN(n1239) );
AND2_X1 U946 ( .A1(n1252), .A2(n1278), .ZN(n1076) );
XOR2_X1 U947 ( .A(KEYINPUT20), .B(n1279), .Z(n1278) );
XOR2_X1 U948 ( .A(n1280), .B(n1281), .Z(G15) );
NOR2_X1 U949 ( .A1(KEYINPUT21), .A2(n1282), .ZN(n1281) );
AND3_X1 U950 ( .A1(n1268), .A2(n1110), .A3(n1103), .ZN(n1280) );
NAND2_X1 U951 ( .A1(n1283), .A2(n1284), .ZN(n1110) );
OR2_X1 U952 ( .A1(n1092), .A2(KEYINPUT10), .ZN(n1284) );
NAND2_X1 U953 ( .A1(n1276), .A2(n1118), .ZN(n1092) );
NAND3_X1 U954 ( .A1(n1118), .A2(n1285), .A3(KEYINPUT10), .ZN(n1283) );
AND2_X1 U955 ( .A1(n1244), .A2(n1108), .ZN(n1268) );
AND2_X1 U956 ( .A1(n1261), .A2(n1286), .ZN(n1244) );
INV_X1 U957 ( .A(n1102), .ZN(n1261) );
NAND2_X1 U958 ( .A1(n1287), .A2(n1100), .ZN(n1102) );
XOR2_X1 U959 ( .A(n1288), .B(n1289), .Z(G12) );
NAND2_X1 U960 ( .A1(KEYINPUT40), .A2(n1238), .ZN(n1289) );
AND3_X1 U961 ( .A1(n1073), .A2(n1106), .A3(n1109), .ZN(n1238) );
NOR2_X1 U962 ( .A1(n1285), .A2(n1118), .ZN(n1109) );
XNOR2_X1 U963 ( .A(n1290), .B(n1169), .ZN(n1118) );
NAND2_X1 U964 ( .A1(G217), .A2(n1291), .ZN(n1169) );
NAND2_X1 U965 ( .A1(n1167), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U966 ( .A(n1293), .B(n1294), .ZN(n1167) );
XNOR2_X1 U967 ( .A(n1295), .B(n1296), .ZN(n1294) );
NAND4_X1 U968 ( .A1(KEYINPUT47), .A2(n1297), .A3(n1298), .A4(n1299), .ZN(n1295) );
NAND2_X1 U969 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
INV_X1 U970 ( .A(KEYINPUT28), .ZN(n1301) );
NAND2_X1 U971 ( .A1(n1302), .A2(n1303), .ZN(n1300) );
XOR2_X1 U972 ( .A(KEYINPUT51), .B(G110), .Z(n1303) );
NAND2_X1 U973 ( .A1(KEYINPUT28), .A2(n1304), .ZN(n1298) );
NAND2_X1 U974 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NAND3_X1 U975 ( .A1(KEYINPUT51), .A2(n1302), .A3(n1288), .ZN(n1306) );
INV_X1 U976 ( .A(n1307), .ZN(n1302) );
OR2_X1 U977 ( .A1(n1288), .A2(KEYINPUT51), .ZN(n1305) );
NAND2_X1 U978 ( .A1(G110), .A2(n1307), .ZN(n1297) );
XNOR2_X1 U979 ( .A(n1277), .B(G128), .ZN(n1307) );
XNOR2_X1 U980 ( .A(G146), .B(n1308), .ZN(n1293) );
NOR2_X1 U981 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U982 ( .A(KEYINPUT6), .B(n1311), .Z(n1310) );
NOR3_X1 U983 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1311) );
NOR2_X1 U984 ( .A1(n1315), .A2(G137), .ZN(n1309) );
NOR2_X1 U985 ( .A1(n1313), .A2(n1312), .ZN(n1315) );
INV_X1 U986 ( .A(G221), .ZN(n1313) );
INV_X1 U987 ( .A(n1276), .ZN(n1285) );
NOR2_X1 U988 ( .A1(n1316), .A2(n1115), .ZN(n1276) );
NOR2_X1 U989 ( .A1(n1317), .A2(G472), .ZN(n1115) );
NOR2_X1 U990 ( .A1(n1121), .A2(n1119), .ZN(n1316) );
INV_X1 U991 ( .A(n1317), .ZN(n1119) );
NAND2_X1 U992 ( .A1(n1318), .A2(n1292), .ZN(n1317) );
XOR2_X1 U993 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U994 ( .A(n1187), .B(n1185), .Z(n1320) );
XOR2_X1 U995 ( .A(n1321), .B(G101), .Z(n1185) );
NAND2_X1 U996 ( .A1(n1322), .A2(G210), .ZN(n1321) );
XOR2_X1 U997 ( .A(n1323), .B(n1324), .Z(n1187) );
XOR2_X1 U998 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U999 ( .A(G119), .B(G116), .Z(n1326) );
NOR2_X1 U1000 ( .A1(KEYINPUT35), .A2(n1327), .ZN(n1325) );
XOR2_X1 U1001 ( .A(n1282), .B(KEYINPUT34), .Z(n1327) );
XNOR2_X1 U1002 ( .A(n1328), .B(n1329), .ZN(n1323) );
XOR2_X1 U1003 ( .A(KEYINPUT57), .B(KEYINPUT46), .Z(n1319) );
INV_X1 U1004 ( .A(G472), .ZN(n1121) );
NAND2_X1 U1005 ( .A1(n1330), .A2(n1331), .ZN(n1106) );
OR3_X1 U1006 ( .A1(n1251), .A2(n1252), .A3(KEYINPUT20), .ZN(n1331) );
NAND2_X1 U1007 ( .A1(KEYINPUT20), .A2(n1103), .ZN(n1330) );
NOR2_X1 U1008 ( .A1(n1279), .A2(n1252), .ZN(n1103) );
XOR2_X1 U1009 ( .A(n1332), .B(n1128), .Z(n1252) );
NOR2_X1 U1010 ( .A1(n1172), .A2(G902), .ZN(n1128) );
XNOR2_X1 U1011 ( .A(n1333), .B(n1334), .ZN(n1172) );
XOR2_X1 U1012 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U1013 ( .A(n1337), .B(n1338), .Z(n1336) );
NOR2_X1 U1014 ( .A1(n1339), .A2(n1312), .ZN(n1338) );
NAND2_X1 U1015 ( .A1(n1340), .A2(n1134), .ZN(n1312) );
XOR2_X1 U1016 ( .A(KEYINPUT26), .B(G234), .Z(n1340) );
INV_X1 U1017 ( .A(G217), .ZN(n1339) );
NAND2_X1 U1018 ( .A1(n1341), .A2(n1342), .ZN(n1337) );
NAND2_X1 U1019 ( .A1(G143), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1020 ( .A(n1344), .B(KEYINPUT5), .Z(n1341) );
NAND2_X1 U1021 ( .A1(G128), .A2(n1345), .ZN(n1344) );
INV_X1 U1022 ( .A(G143), .ZN(n1345) );
XNOR2_X1 U1023 ( .A(G107), .B(n1346), .ZN(n1333) );
XOR2_X1 U1024 ( .A(G122), .B(G116), .Z(n1346) );
NAND2_X1 U1025 ( .A1(KEYINPUT36), .A2(n1129), .ZN(n1332) );
INV_X1 U1026 ( .A(G478), .ZN(n1129) );
INV_X1 U1027 ( .A(n1251), .ZN(n1279) );
XNOR2_X1 U1028 ( .A(n1130), .B(n1347), .ZN(n1251) );
NOR2_X1 U1029 ( .A1(G475), .A2(KEYINPUT1), .ZN(n1347) );
NOR2_X1 U1030 ( .A1(n1178), .A2(G902), .ZN(n1130) );
XOR2_X1 U1031 ( .A(n1348), .B(n1349), .Z(n1178) );
XOR2_X1 U1032 ( .A(n1350), .B(n1296), .Z(n1349) );
XOR2_X1 U1033 ( .A(n1149), .B(n1196), .Z(n1296) );
INV_X1 U1034 ( .A(G140), .ZN(n1196) );
INV_X1 U1035 ( .A(G125), .ZN(n1149) );
XOR2_X1 U1036 ( .A(n1351), .B(n1352), .Z(n1348) );
AND2_X1 U1037 ( .A1(G214), .A2(n1322), .ZN(n1352) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1322) );
XOR2_X1 U1039 ( .A(n1353), .B(n1354), .Z(n1351) );
NOR2_X1 U1040 ( .A1(KEYINPUT18), .A2(n1355), .ZN(n1354) );
XOR2_X1 U1041 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1042 ( .A(n1282), .B(n1358), .Z(n1357) );
NOR2_X1 U1043 ( .A1(G122), .A2(KEYINPUT49), .ZN(n1358) );
NAND2_X1 U1044 ( .A1(KEYINPUT42), .A2(G104), .ZN(n1356) );
AND2_X1 U1045 ( .A1(n1108), .A2(n1233), .ZN(n1073) );
AND2_X1 U1046 ( .A1(n1098), .A2(n1286), .ZN(n1233) );
NAND2_X1 U1047 ( .A1(n1083), .A2(n1359), .ZN(n1286) );
NAND2_X1 U1048 ( .A1(n1263), .A2(n1360), .ZN(n1359) );
INV_X1 U1049 ( .A(G898), .ZN(n1360) );
AND3_X1 U1050 ( .A1(G953), .A2(n1361), .A3(n1362), .ZN(n1263) );
XOR2_X1 U1051 ( .A(n1292), .B(KEYINPUT17), .Z(n1362) );
NAND3_X1 U1052 ( .A1(n1361), .A2(n1134), .A3(G952), .ZN(n1083) );
NAND2_X1 U1053 ( .A1(G237), .A2(G234), .ZN(n1361) );
AND2_X1 U1054 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U1055 ( .A1(G221), .A2(n1291), .ZN(n1100) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1292), .ZN(n1291) );
INV_X1 U1057 ( .A(n1287), .ZN(n1099) );
XOR2_X1 U1058 ( .A(n1363), .B(G469), .Z(n1287) );
NAND2_X1 U1059 ( .A1(n1364), .A2(n1292), .ZN(n1363) );
XOR2_X1 U1060 ( .A(n1365), .B(n1366), .Z(n1364) );
INV_X1 U1061 ( .A(n1193), .ZN(n1366) );
XOR2_X1 U1062 ( .A(n1367), .B(n1368), .Z(n1193) );
XOR2_X1 U1063 ( .A(n1369), .B(n1370), .Z(n1368) );
XOR2_X1 U1064 ( .A(n1371), .B(G101), .Z(n1370) );
NAND2_X1 U1065 ( .A1(G227), .A2(n1372), .ZN(n1371) );
XOR2_X1 U1066 ( .A(KEYINPUT3), .B(G953), .Z(n1372) );
XNOR2_X1 U1067 ( .A(G104), .B(KEYINPUT23), .ZN(n1369) );
XOR2_X1 U1068 ( .A(n1373), .B(n1374), .Z(n1367) );
INV_X1 U1069 ( .A(n1145), .ZN(n1374) );
XOR2_X1 U1070 ( .A(n1343), .B(n1350), .Z(n1145) );
XOR2_X1 U1071 ( .A(n1328), .B(n1375), .Z(n1373) );
NOR2_X1 U1072 ( .A1(G107), .A2(KEYINPUT55), .ZN(n1375) );
NAND3_X1 U1073 ( .A1(n1376), .A2(n1377), .A3(n1378), .ZN(n1328) );
NAND2_X1 U1074 ( .A1(G131), .A2(n1379), .ZN(n1378) );
NAND2_X1 U1075 ( .A1(KEYINPUT16), .A2(n1380), .ZN(n1377) );
NAND2_X1 U1076 ( .A1(n1381), .A2(n1353), .ZN(n1380) );
XOR2_X1 U1077 ( .A(KEYINPUT32), .B(n1379), .Z(n1381) );
NAND2_X1 U1078 ( .A1(n1382), .A2(n1383), .ZN(n1376) );
INV_X1 U1079 ( .A(KEYINPUT16), .ZN(n1383) );
NAND2_X1 U1080 ( .A1(n1384), .A2(n1385), .ZN(n1382) );
NAND3_X1 U1081 ( .A1(KEYINPUT32), .A2(n1353), .A3(n1386), .ZN(n1385) );
INV_X1 U1082 ( .A(G131), .ZN(n1353) );
OR2_X1 U1083 ( .A1(n1386), .A2(KEYINPUT32), .ZN(n1384) );
INV_X1 U1084 ( .A(n1379), .ZN(n1386) );
XNOR2_X1 U1085 ( .A(n1314), .B(n1148), .ZN(n1379) );
INV_X1 U1086 ( .A(n1335), .ZN(n1148) );
XNOR2_X1 U1087 ( .A(G134), .B(KEYINPUT43), .ZN(n1335) );
INV_X1 U1088 ( .A(G137), .ZN(n1314) );
NAND2_X1 U1089 ( .A1(n1387), .A2(KEYINPUT19), .ZN(n1365) );
XOR2_X1 U1090 ( .A(n1288), .B(n1388), .Z(n1387) );
XOR2_X1 U1091 ( .A(KEYINPUT60), .B(G140), .Z(n1388) );
INV_X1 U1092 ( .A(n1182), .ZN(n1108) );
NAND2_X1 U1093 ( .A1(n1389), .A2(n1086), .ZN(n1182) );
XOR2_X1 U1094 ( .A(n1126), .B(n1390), .Z(n1086) );
XOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1127), .Z(n1390) );
AND2_X1 U1096 ( .A1(G210), .A2(n1391), .ZN(n1127) );
NAND2_X1 U1097 ( .A1(n1392), .A2(n1292), .ZN(n1126) );
XOR2_X1 U1098 ( .A(n1393), .B(n1207), .Z(n1392) );
INV_X1 U1099 ( .A(n1200), .ZN(n1207) );
XNOR2_X1 U1100 ( .A(n1159), .B(n1160), .ZN(n1200) );
XOR2_X1 U1101 ( .A(n1394), .B(n1282), .Z(n1160) );
INV_X1 U1102 ( .A(G113), .ZN(n1282) );
NAND2_X1 U1103 ( .A1(n1395), .A2(n1396), .ZN(n1394) );
NAND2_X1 U1104 ( .A1(G116), .A2(n1277), .ZN(n1396) );
XOR2_X1 U1105 ( .A(KEYINPUT22), .B(n1397), .Z(n1395) );
NOR2_X1 U1106 ( .A1(G116), .A2(n1277), .ZN(n1397) );
INV_X1 U1107 ( .A(G119), .ZN(n1277) );
XNOR2_X1 U1108 ( .A(n1398), .B(n1399), .ZN(n1159) );
XOR2_X1 U1109 ( .A(n1400), .B(n1401), .Z(n1399) );
NAND3_X1 U1110 ( .A1(n1402), .A2(n1403), .A3(n1404), .ZN(n1401) );
OR2_X1 U1111 ( .A1(n1405), .A2(n1406), .ZN(n1404) );
NAND3_X1 U1112 ( .A1(n1406), .A2(n1405), .A3(KEYINPUT63), .ZN(n1403) );
INV_X1 U1113 ( .A(G122), .ZN(n1405) );
NOR2_X1 U1114 ( .A1(G110), .A2(KEYINPUT30), .ZN(n1406) );
OR2_X1 U1115 ( .A1(n1288), .A2(KEYINPUT63), .ZN(n1402) );
NAND2_X1 U1116 ( .A1(KEYINPUT4), .A2(n1407), .ZN(n1400) );
XOR2_X1 U1117 ( .A(G107), .B(G104), .Z(n1407) );
XOR2_X1 U1118 ( .A(n1259), .B(KEYINPUT53), .Z(n1398) );
INV_X1 U1119 ( .A(G101), .ZN(n1259) );
XOR2_X1 U1120 ( .A(n1247), .B(n1245), .Z(n1393) );
XNOR2_X1 U1121 ( .A(n1329), .B(G125), .ZN(n1245) );
NAND3_X1 U1122 ( .A1(n1408), .A2(n1409), .A3(n1410), .ZN(n1329) );
OR2_X1 U1123 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
NAND3_X1 U1124 ( .A1(n1412), .A2(n1411), .A3(KEYINPUT8), .ZN(n1409) );
XOR2_X1 U1125 ( .A(n1350), .B(KEYINPUT25), .Z(n1411) );
XOR2_X1 U1126 ( .A(G146), .B(G143), .Z(n1350) );
NOR2_X1 U1127 ( .A1(G128), .A2(KEYINPUT24), .ZN(n1412) );
OR2_X1 U1128 ( .A1(n1343), .A2(KEYINPUT8), .ZN(n1408) );
INV_X1 U1129 ( .A(G128), .ZN(n1343) );
NAND2_X1 U1130 ( .A1(G224), .A2(n1134), .ZN(n1247) );
INV_X1 U1131 ( .A(G953), .ZN(n1134) );
XOR2_X1 U1132 ( .A(n1122), .B(KEYINPUT61), .Z(n1389) );
NAND2_X1 U1133 ( .A1(G214), .A2(n1391), .ZN(n1122) );
NAND2_X1 U1134 ( .A1(n1292), .A2(n1413), .ZN(n1391) );
INV_X1 U1135 ( .A(G237), .ZN(n1413) );
INV_X1 U1136 ( .A(G902), .ZN(n1292) );
INV_X1 U1137 ( .A(G110), .ZN(n1288) );
endmodule


