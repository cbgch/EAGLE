//Key = 0001100010011010011101111001111110100110100000000010111010010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313;

XOR2_X1 U710 ( .A(n989), .B(n990), .Z(G9) );
XOR2_X1 U711 ( .A(KEYINPUT37), .B(G107), .Z(n990) );
NOR2_X1 U712 ( .A1(n991), .A2(n992), .ZN(G75) );
NOR4_X1 U713 ( .A1(n993), .A2(n994), .A3(G953), .A4(n995), .ZN(n992) );
NOR3_X1 U714 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n994) );
NAND3_X1 U715 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n996) );
NAND2_X1 U716 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
XNOR2_X1 U717 ( .A(n1004), .B(KEYINPUT61), .ZN(n1002) );
NAND3_X1 U718 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n993) );
NAND4_X1 U719 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1006) );
NAND2_X1 U720 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND3_X1 U721 ( .A1(n999), .A2(n1014), .A3(n1015), .ZN(n1013) );
NAND2_X1 U722 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND2_X1 U723 ( .A1(n1001), .A2(n1018), .ZN(n1012) );
NAND2_X1 U724 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U725 ( .A1(n1015), .A2(n1021), .ZN(n1020) );
NAND2_X1 U726 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U727 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U728 ( .A1(n999), .A2(n1026), .ZN(n1019) );
NAND2_X1 U729 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U730 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
INV_X1 U731 ( .A(n998), .ZN(n1009) );
NOR3_X1 U732 ( .A1(n995), .A2(G953), .A3(G952), .ZN(n991) );
AND4_X1 U733 ( .A1(n1031), .A2(n999), .A3(n1032), .A4(n1033), .ZN(n995) );
NOR4_X1 U734 ( .A1(n1029), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1033) );
XOR2_X1 U735 ( .A(n1037), .B(n1038), .Z(n1034) );
NOR2_X1 U736 ( .A1(G472), .A2(KEYINPUT36), .ZN(n1038) );
XOR2_X1 U737 ( .A(n1039), .B(n1040), .Z(n1032) );
XNOR2_X1 U738 ( .A(n1041), .B(KEYINPUT45), .ZN(n1039) );
XNOR2_X1 U739 ( .A(n1042), .B(n1030), .ZN(n1031) );
XNOR2_X1 U740 ( .A(KEYINPUT4), .B(KEYINPUT12), .ZN(n1042) );
XOR2_X1 U741 ( .A(n1043), .B(n1044), .Z(G72) );
XOR2_X1 U742 ( .A(n1045), .B(n1046), .Z(n1044) );
NOR2_X1 U743 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
AND2_X1 U744 ( .A1(G227), .A2(G900), .ZN(n1047) );
NAND2_X1 U745 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
NAND2_X1 U746 ( .A1(G953), .A2(n1051), .ZN(n1050) );
XOR2_X1 U747 ( .A(KEYINPUT14), .B(G900), .Z(n1051) );
XOR2_X1 U748 ( .A(n1052), .B(n1053), .Z(n1049) );
XOR2_X1 U749 ( .A(n1054), .B(n1055), .Z(n1053) );
NAND2_X1 U750 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U751 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
XNOR2_X1 U752 ( .A(KEYINPUT25), .B(n1060), .ZN(n1058) );
NAND2_X1 U753 ( .A1(G125), .A2(n1061), .ZN(n1056) );
XNOR2_X1 U754 ( .A(n1062), .B(KEYINPUT0), .ZN(n1061) );
XNOR2_X1 U755 ( .A(KEYINPUT8), .B(n1063), .ZN(n1052) );
NAND2_X1 U756 ( .A1(n1064), .A2(n1065), .ZN(n1043) );
XOR2_X1 U757 ( .A(n1066), .B(n1067), .Z(G69) );
XOR2_X1 U758 ( .A(n1068), .B(n1069), .Z(n1067) );
OR2_X1 U759 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U760 ( .A1(n1072), .A2(n1073), .ZN(n1068) );
NAND2_X1 U761 ( .A1(G898), .A2(G224), .ZN(n1073) );
INV_X1 U762 ( .A(n1048), .ZN(n1072) );
XOR2_X1 U763 ( .A(G953), .B(KEYINPUT18), .Z(n1048) );
NOR2_X1 U764 ( .A1(n1007), .A2(G953), .ZN(n1066) );
NOR2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(G66) );
XNOR2_X1 U766 ( .A(n1076), .B(n1077), .ZN(n1075) );
NOR2_X1 U767 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NOR2_X1 U768 ( .A1(n1074), .A2(n1080), .ZN(G63) );
XOR2_X1 U769 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U770 ( .A1(n1083), .A2(n1079), .ZN(n1081) );
NOR2_X1 U771 ( .A1(n1074), .A2(n1084), .ZN(G60) );
NOR3_X1 U772 ( .A1(n1041), .A2(n1085), .A3(n1086), .ZN(n1084) );
NOR2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U774 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U775 ( .A1(n1065), .A2(n1091), .ZN(n1089) );
NOR3_X1 U776 ( .A1(n1092), .A2(n1090), .A3(n1079), .ZN(n1085) );
XNOR2_X1 U777 ( .A(G104), .B(n1093), .ZN(G6) );
NOR2_X1 U778 ( .A1(n1074), .A2(n1094), .ZN(G57) );
XOR2_X1 U779 ( .A(n1095), .B(n1096), .Z(n1094) );
XOR2_X1 U780 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U781 ( .A1(G101), .A2(KEYINPUT7), .ZN(n1098) );
AND2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
XNOR2_X1 U783 ( .A(n1101), .B(n1102), .ZN(n1095) );
NOR2_X1 U784 ( .A1(n1079), .A2(n1103), .ZN(n1102) );
INV_X1 U785 ( .A(G472), .ZN(n1103) );
NOR2_X1 U786 ( .A1(n1074), .A2(n1104), .ZN(G54) );
XOR2_X1 U787 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U788 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U789 ( .A(n1109), .B(n1110), .Z(n1105) );
NOR2_X1 U790 ( .A1(KEYINPUT46), .A2(n1063), .ZN(n1110) );
XOR2_X1 U791 ( .A(n1111), .B(n1112), .Z(n1109) );
NOR2_X1 U792 ( .A1(n1113), .A2(n1079), .ZN(n1112) );
NOR2_X1 U793 ( .A1(n1074), .A2(n1114), .ZN(G51) );
XOR2_X1 U794 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U795 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U796 ( .A1(n1119), .A2(n1079), .ZN(n1118) );
NAND2_X1 U797 ( .A1(G902), .A2(n1120), .ZN(n1079) );
NAND2_X1 U798 ( .A1(n1007), .A2(n1005), .ZN(n1120) );
INV_X1 U799 ( .A(n1065), .ZN(n1005) );
NAND4_X1 U800 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1065) );
NOR4_X1 U801 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1124) );
NOR3_X1 U802 ( .A1(n1129), .A2(n1130), .A3(n1017), .ZN(n1128) );
XNOR2_X1 U803 ( .A(n1131), .B(KEYINPUT5), .ZN(n1130) );
INV_X1 U804 ( .A(n1132), .ZN(n1126) );
INV_X1 U805 ( .A(n1133), .ZN(n1125) );
NOR2_X1 U806 ( .A1(n1134), .A2(n1135), .ZN(n1123) );
INV_X1 U807 ( .A(n1091), .ZN(n1007) );
NAND4_X1 U808 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1091) );
AND4_X1 U809 ( .A1(n989), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1139) );
NAND3_X1 U810 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n989) );
AND2_X1 U811 ( .A1(n1146), .A2(n1093), .ZN(n1138) );
NAND3_X1 U812 ( .A1(n1143), .A2(n1144), .A3(n1147), .ZN(n1093) );
XNOR2_X1 U813 ( .A(G125), .B(n1148), .ZN(n1115) );
NOR2_X1 U814 ( .A1(KEYINPUT26), .A2(n1149), .ZN(n1148) );
NOR2_X1 U815 ( .A1(n1064), .A2(G952), .ZN(n1074) );
NAND2_X1 U816 ( .A1(n1150), .A2(n1151), .ZN(G48) );
NAND2_X1 U817 ( .A1(n1152), .A2(n1122), .ZN(n1151) );
INV_X1 U818 ( .A(n1153), .ZN(n1122) );
NAND2_X1 U819 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
OR2_X1 U820 ( .A1(KEYINPUT13), .A2(KEYINPUT32), .ZN(n1155) );
NAND3_X1 U821 ( .A1(n1156), .A2(n1157), .A3(KEYINPUT32), .ZN(n1150) );
NAND2_X1 U822 ( .A1(G146), .A2(n1158), .ZN(n1157) );
NAND2_X1 U823 ( .A1(n1159), .A2(n1154), .ZN(n1156) );
INV_X1 U824 ( .A(G146), .ZN(n1154) );
NAND2_X1 U825 ( .A1(n1153), .A2(n1158), .ZN(n1159) );
INV_X1 U826 ( .A(KEYINPUT13), .ZN(n1158) );
NOR3_X1 U827 ( .A1(n1016), .A2(n1027), .A3(n1129), .ZN(n1153) );
INV_X1 U828 ( .A(n1147), .ZN(n1016) );
XOR2_X1 U829 ( .A(G143), .B(n1160), .Z(G45) );
NOR2_X1 U830 ( .A1(KEYINPUT51), .A2(n1121), .ZN(n1160) );
NAND4_X1 U831 ( .A1(n1161), .A2(n1131), .A3(n1036), .A4(n1162), .ZN(n1121) );
XOR2_X1 U832 ( .A(G140), .B(n1135), .Z(G42) );
AND4_X1 U833 ( .A1(n1015), .A2(n1147), .A3(n1163), .A4(n1004), .ZN(n1135) );
NOR2_X1 U834 ( .A1(n1164), .A2(n1022), .ZN(n1163) );
XNOR2_X1 U835 ( .A(n1165), .B(n1127), .ZN(G39) );
NOR3_X1 U836 ( .A1(n997), .A2(n1166), .A3(n1129), .ZN(n1127) );
INV_X1 U837 ( .A(n1001), .ZN(n1166) );
INV_X1 U838 ( .A(n1015), .ZN(n997) );
XOR2_X1 U839 ( .A(G134), .B(n1134), .Z(G36) );
AND3_X1 U840 ( .A1(n1015), .A2(n1145), .A3(n1161), .ZN(n1134) );
NAND2_X1 U841 ( .A1(n1167), .A2(n1168), .ZN(G33) );
OR2_X1 U842 ( .A1(n1132), .A2(G131), .ZN(n1168) );
XOR2_X1 U843 ( .A(n1169), .B(KEYINPUT9), .Z(n1167) );
NAND2_X1 U844 ( .A1(G131), .A2(n1132), .ZN(n1169) );
NAND3_X1 U845 ( .A1(n1015), .A2(n1147), .A3(n1161), .ZN(n1132) );
NOR3_X1 U846 ( .A1(n1022), .A2(n1164), .A3(n1003), .ZN(n1161) );
INV_X1 U847 ( .A(n1143), .ZN(n1022) );
NOR2_X1 U848 ( .A1(n1170), .A2(n1029), .ZN(n1015) );
XNOR2_X1 U849 ( .A(n1171), .B(n1172), .ZN(G30) );
NOR3_X1 U850 ( .A1(n1129), .A2(n1027), .A3(n1017), .ZN(n1172) );
INV_X1 U851 ( .A(n1145), .ZN(n1017) );
NAND4_X1 U852 ( .A1(n1143), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1129) );
XOR2_X1 U853 ( .A(n1146), .B(n1176), .Z(G3) );
NAND2_X1 U854 ( .A1(KEYINPUT50), .A2(G101), .ZN(n1176) );
NAND2_X1 U855 ( .A1(n1177), .A2(n1178), .ZN(n1146) );
XNOR2_X1 U856 ( .A(G125), .B(n1133), .ZN(G27) );
NAND4_X1 U857 ( .A1(n1147), .A2(n1004), .A3(n1179), .A4(n999), .ZN(n1133) );
NOR2_X1 U858 ( .A1(n1164), .A2(n1027), .ZN(n1179) );
INV_X1 U859 ( .A(n1131), .ZN(n1027) );
INV_X1 U860 ( .A(n1175), .ZN(n1164) );
NAND2_X1 U861 ( .A1(n1180), .A2(n998), .ZN(n1175) );
XOR2_X1 U862 ( .A(KEYINPUT3), .B(n1181), .Z(n1180) );
NOR4_X1 U863 ( .A1(G900), .A2(n1182), .A3(n1064), .A4(n1183), .ZN(n1181) );
INV_X1 U864 ( .A(n1184), .ZN(n1182) );
XNOR2_X1 U865 ( .A(G122), .B(n1136), .ZN(G24) );
NAND4_X1 U866 ( .A1(n999), .A2(n1144), .A3(n1036), .A4(n1162), .ZN(n1136) );
AND3_X1 U867 ( .A1(n1008), .A2(n1010), .A3(n1185), .ZN(n1144) );
XNOR2_X1 U868 ( .A(G119), .B(n1137), .ZN(G21) );
NAND4_X1 U869 ( .A1(n1186), .A2(n1001), .A3(n1173), .A4(n1174), .ZN(n1137) );
XNOR2_X1 U870 ( .A(G116), .B(n1142), .ZN(G18) );
NAND3_X1 U871 ( .A1(n1186), .A2(n1145), .A3(n1177), .ZN(n1142) );
NOR2_X1 U872 ( .A1(n1162), .A2(n1187), .ZN(n1145) );
INV_X1 U873 ( .A(n1036), .ZN(n1187) );
XNOR2_X1 U874 ( .A(G113), .B(n1141), .ZN(G15) );
NAND3_X1 U875 ( .A1(n1177), .A2(n1186), .A3(n1147), .ZN(n1141) );
NOR2_X1 U876 ( .A1(n1036), .A2(n1188), .ZN(n1147) );
INV_X1 U877 ( .A(n1162), .ZN(n1188) );
AND2_X1 U878 ( .A1(n999), .A2(n1185), .ZN(n1186) );
NOR2_X1 U879 ( .A1(n1189), .A2(n1024), .ZN(n999) );
INV_X1 U880 ( .A(n1003), .ZN(n1177) );
NAND2_X1 U881 ( .A1(n1008), .A2(n1173), .ZN(n1003) );
XOR2_X1 U882 ( .A(n1010), .B(KEYINPUT29), .Z(n1173) );
INV_X1 U883 ( .A(n1174), .ZN(n1008) );
XNOR2_X1 U884 ( .A(G110), .B(n1140), .ZN(G12) );
NAND2_X1 U885 ( .A1(n1004), .A2(n1178), .ZN(n1140) );
AND3_X1 U886 ( .A1(n1143), .A2(n1185), .A3(n1001), .ZN(n1178) );
NOR2_X1 U887 ( .A1(n1036), .A2(n1162), .ZN(n1001) );
NAND2_X1 U888 ( .A1(n1190), .A2(n1191), .ZN(n1162) );
NAND2_X1 U889 ( .A1(n1192), .A2(n1040), .ZN(n1191) );
XOR2_X1 U890 ( .A(KEYINPUT62), .B(n1193), .Z(n1190) );
NOR2_X1 U891 ( .A1(n1040), .A2(n1192), .ZN(n1193) );
XNOR2_X1 U892 ( .A(KEYINPUT40), .B(n1194), .ZN(n1192) );
INV_X1 U893 ( .A(n1041), .ZN(n1194) );
NOR2_X1 U894 ( .A1(n1088), .A2(G902), .ZN(n1041) );
INV_X1 U895 ( .A(n1092), .ZN(n1088) );
XNOR2_X1 U896 ( .A(n1195), .B(n1196), .ZN(n1092) );
NOR2_X1 U897 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U898 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U899 ( .A(n1201), .B(KEYINPUT2), .Z(n1200) );
AND2_X1 U900 ( .A1(n1201), .A2(n1199), .ZN(n1197) );
XOR2_X1 U901 ( .A(n1202), .B(n1060), .Z(n1199) );
XNOR2_X1 U902 ( .A(G125), .B(n1203), .ZN(n1202) );
NOR2_X1 U903 ( .A1(KEYINPUT41), .A2(n1204), .ZN(n1203) );
NAND3_X1 U904 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1201) );
NAND2_X1 U905 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U906 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XNOR2_X1 U907 ( .A(n1212), .B(n1213), .ZN(n1208) );
NAND4_X1 U908 ( .A1(n1210), .A2(n1211), .A3(n1214), .A4(n1215), .ZN(n1206) );
XNOR2_X1 U909 ( .A(n1212), .B(n1216), .ZN(n1214) );
NAND3_X1 U910 ( .A1(n1217), .A2(n1064), .A3(G214), .ZN(n1212) );
INV_X1 U911 ( .A(KEYINPUT1), .ZN(n1211) );
OR2_X1 U912 ( .A1(n1210), .A2(n1215), .ZN(n1205) );
INV_X1 U913 ( .A(KEYINPUT48), .ZN(n1215) );
XNOR2_X1 U914 ( .A(G131), .B(KEYINPUT16), .ZN(n1210) );
NAND3_X1 U915 ( .A1(n1218), .A2(n1219), .A3(KEYINPUT38), .ZN(n1195) );
NAND2_X1 U916 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
INV_X1 U917 ( .A(KEYINPUT47), .ZN(n1221) );
XNOR2_X1 U918 ( .A(n1222), .B(n1223), .ZN(n1220) );
NAND3_X1 U919 ( .A1(G104), .A2(n1223), .A3(KEYINPUT47), .ZN(n1218) );
XOR2_X1 U920 ( .A(G113), .B(G122), .Z(n1223) );
XNOR2_X1 U921 ( .A(n1090), .B(KEYINPUT42), .ZN(n1040) );
INV_X1 U922 ( .A(G475), .ZN(n1090) );
XOR2_X1 U923 ( .A(n1224), .B(n1083), .Z(n1036) );
INV_X1 U924 ( .A(G478), .ZN(n1083) );
OR2_X1 U925 ( .A1(n1082), .A2(G902), .ZN(n1224) );
XNOR2_X1 U926 ( .A(n1225), .B(n1226), .ZN(n1082) );
AND2_X1 U927 ( .A1(n1227), .A2(G217), .ZN(n1226) );
NAND2_X1 U928 ( .A1(KEYINPUT23), .A2(n1228), .ZN(n1225) );
XOR2_X1 U929 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U930 ( .A(n1231), .B(G107), .Z(n1230) );
NAND3_X1 U931 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
NAND2_X1 U932 ( .A1(KEYINPUT63), .A2(n1213), .ZN(n1234) );
NAND3_X1 U933 ( .A1(n1216), .A2(n1235), .A3(G128), .ZN(n1233) );
NAND2_X1 U934 ( .A1(n1236), .A2(n1171), .ZN(n1232) );
NAND2_X1 U935 ( .A1(n1237), .A2(n1235), .ZN(n1236) );
INV_X1 U936 ( .A(KEYINPUT63), .ZN(n1235) );
XNOR2_X1 U937 ( .A(KEYINPUT53), .B(n1216), .ZN(n1237) );
INV_X1 U938 ( .A(n1213), .ZN(n1216) );
XNOR2_X1 U939 ( .A(G116), .B(n1238), .ZN(n1229) );
XOR2_X1 U940 ( .A(G134), .B(G122), .Z(n1238) );
AND2_X1 U941 ( .A1(n1131), .A2(n1239), .ZN(n1185) );
NAND2_X1 U942 ( .A1(n1240), .A2(n998), .ZN(n1239) );
NAND3_X1 U943 ( .A1(n1184), .A2(n1064), .A3(G952), .ZN(n998) );
NAND3_X1 U944 ( .A1(n1071), .A2(n1184), .A3(G902), .ZN(n1240) );
NAND2_X1 U945 ( .A1(G234), .A2(G237), .ZN(n1184) );
NOR2_X1 U946 ( .A1(n1064), .A2(G898), .ZN(n1071) );
NOR2_X1 U947 ( .A1(n1030), .A2(n1029), .ZN(n1131) );
AND2_X1 U948 ( .A1(G214), .A2(n1241), .ZN(n1029) );
INV_X1 U949 ( .A(n1170), .ZN(n1030) );
XOR2_X1 U950 ( .A(n1242), .B(n1119), .Z(n1170) );
NAND2_X1 U951 ( .A1(G210), .A2(n1241), .ZN(n1119) );
NAND2_X1 U952 ( .A1(n1243), .A2(n1183), .ZN(n1241) );
NAND2_X1 U953 ( .A1(n1244), .A2(n1183), .ZN(n1242) );
XOR2_X1 U954 ( .A(n1245), .B(n1246), .Z(n1244) );
XNOR2_X1 U955 ( .A(n1247), .B(KEYINPUT30), .ZN(n1246) );
NAND2_X1 U956 ( .A1(KEYINPUT22), .A2(n1059), .ZN(n1247) );
INV_X1 U957 ( .A(G125), .ZN(n1059) );
XNOR2_X1 U958 ( .A(n1117), .B(n1149), .ZN(n1245) );
XOR2_X1 U959 ( .A(n1248), .B(n1070), .Z(n1117) );
XNOR2_X1 U960 ( .A(n1249), .B(n1250), .ZN(n1070) );
XOR2_X1 U961 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U962 ( .A(n1253), .B(n1254), .ZN(n1249) );
XNOR2_X1 U963 ( .A(G122), .B(n1222), .ZN(n1254) );
NAND2_X1 U964 ( .A1(n1255), .A2(n1064), .ZN(n1248) );
XOR2_X1 U965 ( .A(KEYINPUT58), .B(G224), .Z(n1255) );
NOR2_X1 U966 ( .A1(n1025), .A2(n1024), .ZN(n1143) );
AND2_X1 U967 ( .A1(G221), .A2(n1256), .ZN(n1024) );
INV_X1 U968 ( .A(n1189), .ZN(n1025) );
XOR2_X1 U969 ( .A(n1257), .B(n1113), .Z(n1189) );
INV_X1 U970 ( .A(G469), .ZN(n1113) );
NAND2_X1 U971 ( .A1(n1258), .A2(n1183), .ZN(n1257) );
XOR2_X1 U972 ( .A(n1259), .B(n1260), .Z(n1258) );
NOR2_X1 U973 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U974 ( .A(n1263), .B(KEYINPUT17), .Z(n1262) );
NAND2_X1 U975 ( .A1(n1107), .A2(n1264), .ZN(n1263) );
NOR2_X1 U976 ( .A1(n1107), .A2(n1264), .ZN(n1261) );
XOR2_X1 U977 ( .A(n1265), .B(n1266), .Z(n1107) );
XOR2_X1 U978 ( .A(KEYINPUT28), .B(n1267), .Z(n1266) );
NOR2_X1 U979 ( .A1(KEYINPUT10), .A2(n1222), .ZN(n1267) );
INV_X1 U980 ( .A(G104), .ZN(n1222) );
XOR2_X1 U981 ( .A(n1054), .B(n1252), .Z(n1265) );
XOR2_X1 U982 ( .A(G101), .B(n1268), .Z(n1252) );
XOR2_X1 U983 ( .A(KEYINPUT54), .B(G107), .Z(n1268) );
XNOR2_X1 U984 ( .A(n1269), .B(n1171), .ZN(n1054) );
NAND2_X1 U985 ( .A1(KEYINPUT21), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U986 ( .A(n1271), .B(n1213), .ZN(n1270) );
NAND3_X1 U987 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1259) );
OR2_X1 U988 ( .A1(n1111), .A2(KEYINPUT11), .ZN(n1274) );
NAND3_X1 U989 ( .A1(KEYINPUT11), .A2(n1111), .A3(n1275), .ZN(n1273) );
INV_X1 U990 ( .A(n1108), .ZN(n1275) );
NAND2_X1 U991 ( .A1(n1108), .A2(n1276), .ZN(n1272) );
NAND2_X1 U992 ( .A1(n1277), .A2(KEYINPUT11), .ZN(n1276) );
XOR2_X1 U993 ( .A(n1111), .B(KEYINPUT35), .Z(n1277) );
NAND2_X1 U994 ( .A1(G227), .A2(n1278), .ZN(n1111) );
XNOR2_X1 U995 ( .A(KEYINPUT24), .B(n1064), .ZN(n1278) );
AND2_X1 U996 ( .A1(n1010), .A2(n1174), .ZN(n1004) );
XOR2_X1 U997 ( .A(n1035), .B(KEYINPUT15), .Z(n1174) );
XOR2_X1 U998 ( .A(n1279), .B(n1078), .Z(n1035) );
NAND2_X1 U999 ( .A1(G217), .A2(n1256), .ZN(n1078) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1183), .ZN(n1256) );
NAND2_X1 U1001 ( .A1(n1076), .A2(n1183), .ZN(n1279) );
XNOR2_X1 U1002 ( .A(n1280), .B(n1281), .ZN(n1076) );
XNOR2_X1 U1003 ( .A(G137), .B(n1282), .ZN(n1281) );
XNOR2_X1 U1004 ( .A(KEYINPUT34), .B(KEYINPUT31), .ZN(n1282) );
XOR2_X1 U1005 ( .A(n1283), .B(n1284), .Z(n1280) );
NOR2_X1 U1006 ( .A1(G125), .A2(KEYINPUT60), .ZN(n1284) );
XOR2_X1 U1007 ( .A(n1285), .B(n1286), .Z(n1283) );
XOR2_X1 U1008 ( .A(n1204), .B(n1287), .Z(n1286) );
NAND2_X1 U1009 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U1010 ( .A1(KEYINPUT56), .A2(n1290), .ZN(n1289) );
INV_X1 U1011 ( .A(n1291), .ZN(n1290) );
NAND2_X1 U1012 ( .A1(KEYINPUT6), .A2(n1291), .ZN(n1288) );
XNOR2_X1 U1013 ( .A(n1292), .B(KEYINPUT52), .ZN(n1204) );
XNOR2_X1 U1014 ( .A(n1293), .B(n1108), .ZN(n1285) );
XOR2_X1 U1015 ( .A(n1251), .B(n1060), .Z(n1108) );
INV_X1 U1016 ( .A(n1062), .ZN(n1060) );
XOR2_X1 U1017 ( .A(G140), .B(KEYINPUT20), .Z(n1062) );
XOR2_X1 U1018 ( .A(G110), .B(KEYINPUT43), .Z(n1251) );
XNOR2_X1 U1019 ( .A(n1294), .B(n1171), .ZN(n1293) );
INV_X1 U1020 ( .A(G128), .ZN(n1171) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1227), .ZN(n1294) );
AND2_X1 U1022 ( .A1(G234), .A2(n1064), .ZN(n1227) );
XNOR2_X1 U1023 ( .A(n1037), .B(n1295), .ZN(n1010) );
NOR2_X1 U1024 ( .A1(G472), .A2(KEYINPUT44), .ZN(n1295) );
NAND2_X1 U1025 ( .A1(n1296), .A2(n1183), .ZN(n1037) );
INV_X1 U1026 ( .A(G902), .ZN(n1183) );
XOR2_X1 U1027 ( .A(n1101), .B(n1297), .Z(n1296) );
XOR2_X1 U1028 ( .A(n1298), .B(G101), .Z(n1297) );
NAND2_X1 U1029 ( .A1(n1299), .A2(n1099), .ZN(n1298) );
NAND3_X1 U1030 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1099) );
XNOR2_X1 U1031 ( .A(n1149), .B(n1264), .ZN(n1302) );
NAND2_X1 U1032 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
INV_X1 U1033 ( .A(n1253), .ZN(n1303) );
NAND3_X1 U1034 ( .A1(G113), .A2(n1305), .A3(KEYINPUT55), .ZN(n1300) );
XOR2_X1 U1035 ( .A(n1100), .B(KEYINPUT49), .Z(n1299) );
NAND3_X1 U1036 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1100) );
XNOR2_X1 U1037 ( .A(n1063), .B(n1149), .ZN(n1308) );
XNOR2_X1 U1038 ( .A(n1309), .B(n1271), .ZN(n1149) );
INV_X1 U1039 ( .A(n1292), .ZN(n1271) );
XOR2_X1 U1040 ( .A(G146), .B(KEYINPUT59), .Z(n1292) );
XNOR2_X1 U1041 ( .A(n1310), .B(n1311), .ZN(n1309) );
NOR2_X1 U1042 ( .A1(G128), .A2(KEYINPUT39), .ZN(n1311) );
NOR2_X1 U1043 ( .A1(KEYINPUT33), .A2(n1213), .ZN(n1310) );
XOR2_X1 U1044 ( .A(G143), .B(KEYINPUT57), .Z(n1213) );
INV_X1 U1045 ( .A(n1264), .ZN(n1063) );
XOR2_X1 U1046 ( .A(G131), .B(n1312), .Z(n1264) );
XNOR2_X1 U1047 ( .A(n1165), .B(G134), .ZN(n1312) );
INV_X1 U1048 ( .A(G137), .ZN(n1165) );
NAND2_X1 U1049 ( .A1(KEYINPUT55), .A2(n1313), .ZN(n1307) );
NAND2_X1 U1050 ( .A1(n1305), .A2(G113), .ZN(n1313) );
NAND2_X1 U1051 ( .A1(n1253), .A2(n1304), .ZN(n1306) );
INV_X1 U1052 ( .A(KEYINPUT55), .ZN(n1304) );
XNOR2_X1 U1053 ( .A(n1305), .B(G113), .ZN(n1253) );
XNOR2_X1 U1054 ( .A(G116), .B(n1291), .ZN(n1305) );
XOR2_X1 U1055 ( .A(G119), .B(KEYINPUT19), .Z(n1291) );
NAND3_X1 U1056 ( .A1(n1217), .A2(n1064), .A3(G210), .ZN(n1101) );
INV_X1 U1057 ( .A(G953), .ZN(n1064) );
XNOR2_X1 U1058 ( .A(n1243), .B(KEYINPUT27), .ZN(n1217) );
INV_X1 U1059 ( .A(G237), .ZN(n1243) );
endmodule


