//Key = 0101000001011010111110011011011100100101101000110000000001010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346;

NAND2_X1 U745 ( .A1(n1035), .A2(n1036), .ZN(G9) );
NAND2_X1 U746 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
XOR2_X1 U747 ( .A(KEYINPUT3), .B(n1039), .Z(n1035) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1039) );
NOR2_X1 U749 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR4_X1 U750 ( .A1(G953), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1041) );
NOR2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U752 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
INV_X1 U754 ( .A(n1051), .ZN(n1050) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1049) );
NOR2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR3_X1 U757 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1054) );
NOR2_X1 U758 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U759 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR3_X1 U761 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1057) );
NOR2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1056) );
XNOR2_X1 U763 ( .A(n1070), .B(KEYINPUT28), .ZN(n1068) );
NOR3_X1 U764 ( .A1(n1065), .A2(n1071), .A3(n1060), .ZN(n1052) );
NOR2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U766 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR4_X1 U767 ( .A1(n1076), .A2(n1055), .A3(n1060), .A4(n1065), .ZN(n1047) );
INV_X1 U768 ( .A(n1077), .ZN(n1055) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR3_X1 U770 ( .A1(n1042), .A2(G953), .A3(G952), .ZN(n1040) );
AND4_X1 U771 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1042) );
NOR3_X1 U772 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
XNOR2_X1 U773 ( .A(KEYINPUT7), .B(n1087), .ZN(n1086) );
XNOR2_X1 U774 ( .A(KEYINPUT6), .B(n1088), .ZN(n1085) );
NAND3_X1 U775 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1084) );
XNOR2_X1 U776 ( .A(n1092), .B(G472), .ZN(n1091) );
NOR3_X1 U777 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1082) );
XOR2_X1 U778 ( .A(KEYINPUT47), .B(n1096), .Z(n1080) );
XOR2_X1 U779 ( .A(n1097), .B(n1098), .Z(G72) );
NOR2_X1 U780 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR3_X1 U781 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1100) );
NOR2_X1 U782 ( .A1(G953), .A2(n1104), .ZN(n1099) );
XOR2_X1 U783 ( .A(n1105), .B(n1102), .Z(n1104) );
XOR2_X1 U784 ( .A(n1106), .B(n1107), .Z(n1102) );
XNOR2_X1 U785 ( .A(n1108), .B(n1109), .ZN(n1107) );
XNOR2_X1 U786 ( .A(n1110), .B(G137), .ZN(n1109) );
XOR2_X1 U787 ( .A(n1111), .B(n1112), .Z(n1106) );
XNOR2_X1 U788 ( .A(n1113), .B(n1114), .ZN(n1112) );
NOR2_X1 U789 ( .A1(G125), .A2(KEYINPUT54), .ZN(n1114) );
NAND2_X1 U790 ( .A1(KEYINPUT9), .A2(n1115), .ZN(n1113) );
NAND3_X1 U791 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1105) );
XNOR2_X1 U792 ( .A(KEYINPUT57), .B(n1119), .ZN(n1117) );
NAND3_X1 U793 ( .A1(n1120), .A2(n1121), .A3(KEYINPUT46), .ZN(n1097) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1121) );
XOR2_X1 U795 ( .A(n1122), .B(n1123), .Z(G69) );
XOR2_X1 U796 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND2_X1 U797 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U798 ( .A1(G953), .A2(n1128), .ZN(n1127) );
XOR2_X1 U799 ( .A(n1129), .B(n1130), .Z(n1126) );
XNOR2_X1 U800 ( .A(n1131), .B(n1132), .ZN(n1130) );
XOR2_X1 U801 ( .A(n1133), .B(KEYINPUT41), .Z(n1129) );
NAND2_X1 U802 ( .A1(n1120), .A2(n1134), .ZN(n1124) );
NAND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1134) );
XNOR2_X1 U804 ( .A(n1101), .B(KEYINPUT53), .ZN(n1120) );
NOR2_X1 U805 ( .A1(n1135), .A2(G953), .ZN(n1122) );
NOR2_X1 U806 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XNOR2_X1 U807 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U808 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U809 ( .A1(n1136), .A2(n1142), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1143), .B(n1144), .ZN(n1142) );
XOR2_X1 U811 ( .A(n1145), .B(KEYINPUT50), .Z(n1144) );
NAND3_X1 U812 ( .A1(n1146), .A2(n1044), .A3(G478), .ZN(n1145) );
XNOR2_X1 U813 ( .A(KEYINPUT35), .B(n1147), .ZN(n1146) );
NOR2_X1 U814 ( .A1(n1136), .A2(n1148), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U816 ( .A1(n1151), .A2(n1141), .ZN(n1150) );
NAND3_X1 U817 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(G6) );
OR2_X1 U818 ( .A1(G104), .A2(KEYINPUT31), .ZN(n1154) );
NAND3_X1 U819 ( .A1(KEYINPUT31), .A2(G104), .A3(n1155), .ZN(n1153) );
NAND2_X1 U820 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
NAND2_X1 U821 ( .A1(KEYINPUT31), .A2(n1158), .ZN(n1157) );
XOR2_X1 U822 ( .A(KEYINPUT8), .B(G104), .Z(n1158) );
INV_X1 U823 ( .A(n1155), .ZN(n1156) );
NOR2_X1 U824 ( .A1(n1136), .A2(n1159), .ZN(G57) );
XOR2_X1 U825 ( .A(n1160), .B(n1161), .Z(n1159) );
XNOR2_X1 U826 ( .A(G101), .B(n1162), .ZN(n1161) );
NAND2_X1 U827 ( .A1(KEYINPUT61), .A2(n1163), .ZN(n1162) );
XOR2_X1 U828 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U829 ( .A(n1166), .B(n1167), .Z(n1160) );
NOR2_X1 U830 ( .A1(n1168), .A2(n1141), .ZN(n1167) );
NAND2_X1 U831 ( .A1(KEYINPUT29), .A2(n1169), .ZN(n1166) );
NOR2_X1 U832 ( .A1(n1136), .A2(n1170), .ZN(G54) );
XOR2_X1 U833 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U834 ( .A1(n1173), .A2(n1141), .ZN(n1172) );
XNOR2_X1 U835 ( .A(G469), .B(KEYINPUT22), .ZN(n1173) );
NAND2_X1 U836 ( .A1(KEYINPUT17), .A2(n1174), .ZN(n1171) );
XOR2_X1 U837 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U838 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR2_X1 U839 ( .A1(KEYINPUT48), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U840 ( .A(G110), .B(G140), .ZN(n1179) );
NAND2_X1 U841 ( .A1(n1180), .A2(n1181), .ZN(n1175) );
NAND2_X1 U842 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XOR2_X1 U843 ( .A(KEYINPUT16), .B(n1184), .Z(n1180) );
NOR2_X1 U844 ( .A1(n1182), .A2(n1183), .ZN(n1184) );
XOR2_X1 U845 ( .A(n1111), .B(n1185), .Z(n1182) );
AND2_X1 U846 ( .A1(KEYINPUT30), .A2(n1131), .ZN(n1185) );
NOR2_X1 U847 ( .A1(n1136), .A2(n1186), .ZN(G51) );
XNOR2_X1 U848 ( .A(n1187), .B(n1188), .ZN(n1186) );
XOR2_X1 U849 ( .A(KEYINPUT2), .B(n1189), .Z(n1188) );
NOR2_X1 U850 ( .A1(n1190), .A2(n1141), .ZN(n1189) );
NAND2_X1 U851 ( .A1(G902), .A2(n1044), .ZN(n1141) );
NAND3_X1 U852 ( .A1(n1118), .A2(n1191), .A3(n1135), .ZN(n1044) );
AND2_X1 U853 ( .A1(n1192), .A2(n1193), .ZN(n1135) );
NOR4_X1 U854 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1037), .ZN(n1193) );
AND3_X1 U855 ( .A1(n1078), .A2(n1197), .A3(n1198), .ZN(n1037) );
INV_X1 U856 ( .A(n1199), .ZN(n1194) );
AND4_X1 U857 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1155), .ZN(n1192) );
NAND3_X1 U858 ( .A1(n1198), .A2(n1197), .A3(n1079), .ZN(n1155) );
XOR2_X1 U859 ( .A(KEYINPUT49), .B(n1203), .Z(n1191) );
AND2_X1 U860 ( .A1(n1119), .A2(n1116), .ZN(n1203) );
AND3_X1 U861 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1116) );
AND4_X1 U862 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1118) );
NAND4_X1 U863 ( .A1(n1211), .A2(n1070), .A3(n1073), .A4(n1212), .ZN(n1208) );
XNOR2_X1 U864 ( .A(KEYINPUT37), .B(n1213), .ZN(n1212) );
NAND4_X1 U865 ( .A1(n1214), .A2(n1062), .A3(n1215), .A4(n1216), .ZN(n1207) );
AND2_X1 U866 ( .A1(G953), .A2(n1217), .ZN(n1136) );
XOR2_X1 U867 ( .A(KEYINPUT27), .B(G952), .Z(n1217) );
XNOR2_X1 U868 ( .A(n1218), .B(n1209), .ZN(G48) );
NAND3_X1 U869 ( .A1(n1079), .A2(n1062), .A3(n1219), .ZN(n1209) );
XNOR2_X1 U870 ( .A(G146), .B(KEYINPUT24), .ZN(n1218) );
XOR2_X1 U871 ( .A(n1220), .B(n1221), .Z(G45) );
NAND4_X1 U872 ( .A1(n1214), .A2(n1222), .A3(n1215), .A4(n1216), .ZN(n1221) );
XOR2_X1 U873 ( .A(KEYINPUT60), .B(n1062), .Z(n1222) );
NAND2_X1 U874 ( .A1(KEYINPUT39), .A2(n1223), .ZN(n1220) );
XNOR2_X1 U875 ( .A(KEYINPUT62), .B(n1224), .ZN(n1223) );
XOR2_X1 U876 ( .A(n1225), .B(n1226), .Z(G42) );
NOR2_X1 U877 ( .A1(KEYINPUT15), .A2(n1110), .ZN(n1226) );
NOR3_X1 U878 ( .A1(n1227), .A2(n1228), .A3(n1065), .ZN(n1225) );
INV_X1 U879 ( .A(n1070), .ZN(n1065) );
XNOR2_X1 U880 ( .A(G137), .B(n1210), .ZN(G39) );
NAND3_X1 U881 ( .A1(n1070), .A2(n1051), .A3(n1219), .ZN(n1210) );
XNOR2_X1 U882 ( .A(G134), .B(n1119), .ZN(G36) );
NAND3_X1 U883 ( .A1(n1070), .A2(n1078), .A3(n1214), .ZN(n1119) );
XNOR2_X1 U884 ( .A(G131), .B(n1206), .ZN(G33) );
NAND3_X1 U885 ( .A1(n1070), .A2(n1079), .A3(n1214), .ZN(n1206) );
NOR2_X1 U886 ( .A1(n1228), .A2(n1069), .ZN(n1214) );
NOR2_X1 U887 ( .A1(n1063), .A2(n1093), .ZN(n1070) );
INV_X1 U888 ( .A(n1064), .ZN(n1093) );
XNOR2_X1 U889 ( .A(n1229), .B(n1230), .ZN(G30) );
NOR2_X1 U890 ( .A1(KEYINPUT36), .A2(n1204), .ZN(n1230) );
NAND3_X1 U891 ( .A1(n1078), .A2(n1062), .A3(n1219), .ZN(n1204) );
NOR3_X1 U892 ( .A1(n1231), .A2(n1066), .A3(n1228), .ZN(n1219) );
NAND2_X1 U893 ( .A1(n1073), .A2(n1213), .ZN(n1228) );
INV_X1 U894 ( .A(n1232), .ZN(n1066) );
NAND2_X1 U895 ( .A1(n1233), .A2(n1234), .ZN(G3) );
NAND2_X1 U896 ( .A1(n1196), .A2(n1235), .ZN(n1234) );
XOR2_X1 U897 ( .A(KEYINPUT1), .B(n1236), .Z(n1233) );
NOR2_X1 U898 ( .A1(n1196), .A2(n1235), .ZN(n1236) );
AND3_X1 U899 ( .A1(n1051), .A2(n1198), .A3(n1237), .ZN(n1196) );
XNOR2_X1 U900 ( .A(G125), .B(n1205), .ZN(G27) );
NAND4_X1 U901 ( .A1(n1211), .A2(n1062), .A3(n1077), .A4(n1213), .ZN(n1205) );
NAND2_X1 U902 ( .A1(n1046), .A2(n1238), .ZN(n1213) );
NAND4_X1 U903 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1103), .ZN(n1238) );
INV_X1 U904 ( .A(G900), .ZN(n1103) );
INV_X1 U905 ( .A(n1227), .ZN(n1211) );
NAND3_X1 U906 ( .A1(n1231), .A2(n1232), .A3(n1079), .ZN(n1227) );
XNOR2_X1 U907 ( .A(G122), .B(n1202), .ZN(G24) );
NAND4_X1 U908 ( .A1(n1240), .A2(n1197), .A3(n1215), .A4(n1216), .ZN(n1202) );
INV_X1 U909 ( .A(n1060), .ZN(n1197) );
NAND2_X1 U910 ( .A1(n1241), .A2(n1231), .ZN(n1060) );
XNOR2_X1 U911 ( .A(G119), .B(n1201), .ZN(G21) );
NAND4_X1 U912 ( .A1(n1240), .A2(n1051), .A3(n1067), .A4(n1232), .ZN(n1201) );
XNOR2_X1 U913 ( .A(n1200), .B(n1242), .ZN(G18) );
NOR2_X1 U914 ( .A1(KEYINPUT51), .A2(n1243), .ZN(n1242) );
NAND3_X1 U915 ( .A1(n1237), .A2(n1078), .A3(n1240), .ZN(n1200) );
AND3_X1 U916 ( .A1(n1077), .A2(n1244), .A3(n1062), .ZN(n1240) );
XOR2_X1 U917 ( .A(n1245), .B(KEYINPUT10), .Z(n1062) );
NOR2_X1 U918 ( .A1(n1215), .A2(n1246), .ZN(n1078) );
XNOR2_X1 U919 ( .A(n1195), .B(n1247), .ZN(G15) );
XOR2_X1 U920 ( .A(KEYINPUT18), .B(G113), .Z(n1247) );
AND3_X1 U921 ( .A1(n1079), .A2(n1237), .A3(n1248), .ZN(n1195) );
AND3_X1 U922 ( .A1(n1245), .A2(n1244), .A3(n1077), .ZN(n1248) );
NAND2_X1 U923 ( .A1(n1249), .A2(n1250), .ZN(n1077) );
OR3_X1 U924 ( .A1(n1074), .A2(n1095), .A3(KEYINPUT21), .ZN(n1250) );
NAND2_X1 U925 ( .A1(KEYINPUT21), .A2(n1073), .ZN(n1249) );
INV_X1 U926 ( .A(n1069), .ZN(n1237) );
NAND2_X1 U927 ( .A1(n1241), .A2(n1067), .ZN(n1069) );
XNOR2_X1 U928 ( .A(n1232), .B(KEYINPUT55), .ZN(n1241) );
NOR2_X1 U929 ( .A1(n1216), .A2(n1087), .ZN(n1079) );
INV_X1 U930 ( .A(n1215), .ZN(n1087) );
XNOR2_X1 U931 ( .A(G110), .B(n1199), .ZN(G12) );
NAND4_X1 U932 ( .A1(n1051), .A2(n1198), .A3(n1231), .A4(n1232), .ZN(n1199) );
XNOR2_X1 U933 ( .A(n1090), .B(KEYINPUT56), .ZN(n1232) );
XNOR2_X1 U934 ( .A(n1251), .B(n1140), .ZN(n1090) );
NAND2_X1 U935 ( .A1(G217), .A2(n1252), .ZN(n1140) );
NAND2_X1 U936 ( .A1(n1138), .A2(n1147), .ZN(n1251) );
XNOR2_X1 U937 ( .A(n1253), .B(n1254), .ZN(n1138) );
XOR2_X1 U938 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U939 ( .A(G137), .B(n1257), .ZN(n1256) );
XOR2_X1 U940 ( .A(KEYINPUT44), .B(G146), .Z(n1255) );
XOR2_X1 U941 ( .A(n1258), .B(n1259), .Z(n1253) );
NOR2_X1 U942 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U943 ( .A(n1262), .B(KEYINPUT11), .Z(n1261) );
NAND2_X1 U944 ( .A1(G125), .A2(n1110), .ZN(n1262) );
NOR2_X1 U945 ( .A1(G125), .A2(n1110), .ZN(n1260) );
XOR2_X1 U946 ( .A(n1263), .B(n1264), .Z(n1258) );
AND2_X1 U947 ( .A1(G221), .A2(n1265), .ZN(n1264) );
NAND2_X1 U948 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
NAND2_X1 U949 ( .A1(n1268), .A2(n1229), .ZN(n1267) );
XNOR2_X1 U950 ( .A(G119), .B(KEYINPUT59), .ZN(n1268) );
XOR2_X1 U951 ( .A(KEYINPUT19), .B(n1269), .Z(n1266) );
NOR2_X1 U952 ( .A1(G119), .A2(n1229), .ZN(n1269) );
INV_X1 U953 ( .A(G128), .ZN(n1229) );
INV_X1 U954 ( .A(n1067), .ZN(n1231) );
XOR2_X1 U955 ( .A(n1270), .B(n1168), .Z(n1067) );
INV_X1 U956 ( .A(G472), .ZN(n1168) );
NAND2_X1 U957 ( .A1(KEYINPUT42), .A2(n1092), .ZN(n1270) );
AND2_X1 U958 ( .A1(n1271), .A2(n1147), .ZN(n1092) );
XOR2_X1 U959 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U960 ( .A(n1274), .B(n1164), .ZN(n1273) );
XNOR2_X1 U961 ( .A(n1133), .B(n1183), .ZN(n1164) );
NAND2_X1 U962 ( .A1(KEYINPUT12), .A2(n1165), .ZN(n1274) );
XNOR2_X1 U963 ( .A(n1169), .B(n1275), .ZN(n1272) );
XNOR2_X1 U964 ( .A(KEYINPUT14), .B(n1235), .ZN(n1275) );
INV_X1 U965 ( .A(G101), .ZN(n1235) );
AND3_X1 U966 ( .A1(n1276), .A2(n1101), .A3(G210), .ZN(n1169) );
AND3_X1 U967 ( .A1(n1245), .A2(n1244), .A3(n1073), .ZN(n1198) );
NOR2_X1 U968 ( .A1(n1089), .A2(n1095), .ZN(n1073) );
INV_X1 U969 ( .A(n1075), .ZN(n1095) );
NAND2_X1 U970 ( .A1(n1277), .A2(n1252), .ZN(n1075) );
NAND2_X1 U971 ( .A1(G234), .A2(n1147), .ZN(n1252) );
XNOR2_X1 U972 ( .A(G221), .B(KEYINPUT26), .ZN(n1277) );
INV_X1 U973 ( .A(n1074), .ZN(n1089) );
XNOR2_X1 U974 ( .A(n1278), .B(G469), .ZN(n1074) );
NAND2_X1 U975 ( .A1(n1279), .A2(n1147), .ZN(n1278) );
XOR2_X1 U976 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U977 ( .A(n1111), .B(n1282), .Z(n1281) );
XNOR2_X1 U978 ( .A(n1183), .B(n1131), .ZN(n1282) );
XNOR2_X1 U979 ( .A(n1283), .B(n1284), .ZN(n1183) );
XNOR2_X1 U980 ( .A(n1115), .B(n1285), .ZN(n1284) );
NOR2_X1 U981 ( .A1(G137), .A2(KEYINPUT0), .ZN(n1285) );
INV_X1 U982 ( .A(G131), .ZN(n1115) );
XNOR2_X1 U983 ( .A(G134), .B(KEYINPUT4), .ZN(n1283) );
XOR2_X1 U984 ( .A(n1286), .B(n1287), .Z(n1111) );
XOR2_X1 U985 ( .A(KEYINPUT45), .B(KEYINPUT40), .Z(n1287) );
XNOR2_X1 U986 ( .A(G128), .B(n1288), .ZN(n1286) );
XOR2_X1 U987 ( .A(n1289), .B(n1290), .Z(n1280) );
NOR2_X1 U988 ( .A1(KEYINPUT38), .A2(n1110), .ZN(n1290) );
XNOR2_X1 U989 ( .A(n1257), .B(n1177), .ZN(n1289) );
NAND2_X1 U990 ( .A1(G227), .A2(n1101), .ZN(n1177) );
INV_X1 U991 ( .A(G110), .ZN(n1257) );
NAND2_X1 U992 ( .A1(n1046), .A2(n1291), .ZN(n1244) );
NAND4_X1 U993 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1128), .ZN(n1291) );
INV_X1 U994 ( .A(G898), .ZN(n1128) );
NAND3_X1 U995 ( .A1(n1239), .A2(n1101), .A3(G952), .ZN(n1046) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1239) );
AND2_X1 U997 ( .A1(n1064), .A2(n1063), .ZN(n1245) );
NAND2_X1 U998 ( .A1(n1081), .A2(n1088), .ZN(n1063) );
NAND3_X1 U999 ( .A1(n1190), .A2(n1147), .A3(n1187), .ZN(n1088) );
NAND2_X1 U1000 ( .A1(n1292), .A2(n1293), .ZN(n1081) );
NAND2_X1 U1001 ( .A1(n1187), .A2(n1147), .ZN(n1293) );
XOR2_X1 U1002 ( .A(n1294), .B(n1295), .Z(n1187) );
XOR2_X1 U1003 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1004 ( .A(n1133), .B(n1298), .Z(n1297) );
AND2_X1 U1005 ( .A1(n1101), .A2(G224), .ZN(n1298) );
XNOR2_X1 U1006 ( .A(G113), .B(n1299), .ZN(n1133) );
XNOR2_X1 U1007 ( .A(n1300), .B(G116), .ZN(n1299) );
INV_X1 U1008 ( .A(G119), .ZN(n1300) );
XNOR2_X1 U1009 ( .A(G125), .B(KEYINPUT25), .ZN(n1296) );
XOR2_X1 U1010 ( .A(n1301), .B(n1302), .Z(n1294) );
NOR2_X1 U1011 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NOR2_X1 U1012 ( .A1(KEYINPUT33), .A2(n1305), .ZN(n1304) );
NOR2_X1 U1013 ( .A1(KEYINPUT23), .A2(n1131), .ZN(n1303) );
INV_X1 U1014 ( .A(n1305), .ZN(n1131) );
XOR2_X1 U1015 ( .A(G101), .B(n1306), .Z(n1305) );
XNOR2_X1 U1016 ( .A(n1038), .B(G104), .ZN(n1306) );
XNOR2_X1 U1017 ( .A(n1132), .B(n1165), .ZN(n1301) );
XNOR2_X1 U1018 ( .A(n1307), .B(G128), .ZN(n1165) );
NAND2_X1 U1019 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U1020 ( .A1(G146), .A2(n1224), .ZN(n1309) );
XOR2_X1 U1021 ( .A(n1310), .B(KEYINPUT32), .Z(n1308) );
OR2_X1 U1022 ( .A1(n1224), .A2(G146), .ZN(n1310) );
XNOR2_X1 U1023 ( .A(G110), .B(n1311), .ZN(n1132) );
INV_X1 U1024 ( .A(n1190), .ZN(n1292) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1312), .ZN(n1190) );
NAND2_X1 U1026 ( .A1(G214), .A2(n1312), .ZN(n1064) );
NAND2_X1 U1027 ( .A1(n1276), .A2(n1147), .ZN(n1312) );
NOR2_X1 U1028 ( .A1(n1216), .A2(n1215), .ZN(n1051) );
XOR2_X1 U1029 ( .A(n1313), .B(n1151), .Z(n1215) );
INV_X1 U1030 ( .A(G475), .ZN(n1151) );
NAND2_X1 U1031 ( .A1(n1149), .A2(n1147), .ZN(n1313) );
INV_X1 U1032 ( .A(G902), .ZN(n1147) );
XNOR2_X1 U1033 ( .A(n1314), .B(n1315), .ZN(n1149) );
XOR2_X1 U1034 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1035 ( .A(n1311), .B(G113), .ZN(n1317) );
XNOR2_X1 U1036 ( .A(n1110), .B(G131), .ZN(n1316) );
INV_X1 U1037 ( .A(G140), .ZN(n1110) );
XOR2_X1 U1038 ( .A(n1318), .B(n1319), .Z(n1314) );
XNOR2_X1 U1039 ( .A(G104), .B(n1320), .ZN(n1319) );
NAND2_X1 U1040 ( .A1(KEYINPUT63), .A2(G125), .ZN(n1320) );
XOR2_X1 U1041 ( .A(n1321), .B(n1288), .Z(n1318) );
XNOR2_X1 U1042 ( .A(G146), .B(n1224), .ZN(n1288) );
NAND3_X1 U1043 ( .A1(n1276), .A2(n1101), .A3(G214), .ZN(n1321) );
INV_X1 U1044 ( .A(G237), .ZN(n1276) );
INV_X1 U1045 ( .A(n1246), .ZN(n1216) );
NOR2_X1 U1046 ( .A1(n1094), .A2(n1096), .ZN(n1246) );
NOR3_X1 U1047 ( .A1(G478), .A2(G902), .A3(n1143), .ZN(n1096) );
AND2_X1 U1048 ( .A1(G478), .A2(n1322), .ZN(n1094) );
OR2_X1 U1049 ( .A1(n1143), .A2(G902), .ZN(n1322) );
XNOR2_X1 U1050 ( .A(n1323), .B(n1324), .ZN(n1143) );
NOR3_X1 U1051 ( .A1(n1325), .A2(KEYINPUT58), .A3(n1326), .ZN(n1324) );
NOR2_X1 U1052 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
XNOR2_X1 U1053 ( .A(n1329), .B(n1038), .ZN(n1327) );
INV_X1 U1054 ( .A(G107), .ZN(n1038) );
XOR2_X1 U1055 ( .A(KEYINPUT13), .B(n1330), .Z(n1325) );
NOR2_X1 U1056 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XNOR2_X1 U1057 ( .A(G107), .B(n1329), .ZN(n1332) );
NAND3_X1 U1058 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1329) );
NAND2_X1 U1059 ( .A1(KEYINPUT43), .A2(n1311), .ZN(n1335) );
INV_X1 U1060 ( .A(G122), .ZN(n1311) );
NAND3_X1 U1061 ( .A1(G122), .A2(n1336), .A3(n1243), .ZN(n1334) );
INV_X1 U1062 ( .A(G116), .ZN(n1243) );
NAND2_X1 U1063 ( .A1(G116), .A2(n1337), .ZN(n1333) );
NAND2_X1 U1064 ( .A1(n1338), .A2(n1336), .ZN(n1337) );
INV_X1 U1065 ( .A(KEYINPUT43), .ZN(n1336) );
XNOR2_X1 U1066 ( .A(G122), .B(KEYINPUT20), .ZN(n1338) );
INV_X1 U1067 ( .A(n1328), .ZN(n1331) );
NAND2_X1 U1068 ( .A1(n1339), .A2(n1340), .ZN(n1328) );
NAND3_X1 U1069 ( .A1(KEYINPUT34), .A2(G128), .A3(n1341), .ZN(n1340) );
XNOR2_X1 U1070 ( .A(G134), .B(n1342), .ZN(n1341) );
NOR2_X1 U1071 ( .A1(G143), .A2(KEYINPUT5), .ZN(n1342) );
NAND2_X1 U1072 ( .A1(n1343), .A2(n1344), .ZN(n1339) );
NAND2_X1 U1073 ( .A1(KEYINPUT34), .A2(G128), .ZN(n1344) );
XNOR2_X1 U1074 ( .A(n1345), .B(n1108), .ZN(n1343) );
INV_X1 U1075 ( .A(G134), .ZN(n1108) );
OR2_X1 U1076 ( .A1(n1224), .A2(KEYINPUT5), .ZN(n1345) );
INV_X1 U1077 ( .A(G143), .ZN(n1224) );
NAND2_X1 U1078 ( .A1(G217), .A2(n1265), .ZN(n1323) );
AND2_X1 U1079 ( .A1(n1346), .A2(n1101), .ZN(n1265) );
INV_X1 U1080 ( .A(G953), .ZN(n1101) );
XOR2_X1 U1081 ( .A(KEYINPUT52), .B(G234), .Z(n1346) );
endmodule


