//Key = 1000011001011101000111000111000011111100110110010100111011001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385;

XOR2_X1 U756 ( .A(G107), .B(n1057), .Z(G9) );
NOR2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(G75) );
NOR4_X1 U758 ( .A1(G953), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1059) );
NOR2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U760 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U761 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
INV_X1 U762 ( .A(n1069), .ZN(n1068) );
NOR2_X1 U763 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR3_X1 U765 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1072) );
NOR3_X1 U766 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
NOR2_X1 U767 ( .A1(n1080), .A2(n1081), .ZN(n1074) );
NOR2_X1 U768 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR2_X1 U769 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR3_X1 U770 ( .A1(n1081), .A2(n1086), .A3(n1078), .ZN(n1070) );
NOR2_X1 U771 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U772 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR4_X1 U773 ( .A1(n1091), .A2(n1073), .A3(n1078), .A4(n1081), .ZN(n1065) );
NOR2_X1 U774 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR3_X1 U775 ( .A1(n1060), .A2(G953), .A3(G952), .ZN(n1058) );
AND4_X1 U776 ( .A1(n1094), .A2(n1069), .A3(n1095), .A4(n1096), .ZN(n1060) );
NOR4_X1 U777 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XOR2_X1 U778 ( .A(n1101), .B(n1102), .Z(n1099) );
NOR2_X1 U779 ( .A1(n1103), .A2(KEYINPUT39), .ZN(n1102) );
XOR2_X1 U780 ( .A(n1104), .B(n1105), .Z(n1095) );
NOR2_X1 U781 ( .A1(KEYINPUT63), .A2(n1106), .ZN(n1105) );
XNOR2_X1 U782 ( .A(n1107), .B(G472), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1108), .A2(n1109), .ZN(G72) );
NAND2_X1 U784 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
OR2_X1 U785 ( .A1(n1112), .A2(G227), .ZN(n1111) );
NAND3_X1 U786 ( .A1(G953), .A2(n1113), .A3(n1114), .ZN(n1108) );
INV_X1 U787 ( .A(n1110), .ZN(n1114) );
XNOR2_X1 U788 ( .A(n1115), .B(n1116), .ZN(n1110) );
NOR2_X1 U789 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U790 ( .A(n1119), .B(n1120), .Z(n1118) );
XNOR2_X1 U791 ( .A(n1121), .B(n1122), .ZN(n1120) );
NOR2_X1 U792 ( .A1(KEYINPUT55), .A2(n1123), .ZN(n1122) );
XOR2_X1 U793 ( .A(n1124), .B(n1125), .Z(n1123) );
XNOR2_X1 U794 ( .A(n1126), .B(n1127), .ZN(n1125) );
NAND2_X1 U795 ( .A1(KEYINPUT54), .A2(n1128), .ZN(n1127) );
NAND2_X1 U796 ( .A1(n1112), .A2(n1129), .ZN(n1115) );
NAND2_X1 U797 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U798 ( .A1(G900), .A2(G227), .ZN(n1113) );
NAND2_X1 U799 ( .A1(n1132), .A2(n1133), .ZN(G69) );
NAND3_X1 U800 ( .A1(G953), .A2(n1134), .A3(n1135), .ZN(n1133) );
XOR2_X1 U801 ( .A(KEYINPUT40), .B(n1136), .Z(n1132) );
NOR2_X1 U802 ( .A1(n1135), .A2(n1137), .ZN(n1136) );
AND2_X1 U803 ( .A1(n1134), .A2(G953), .ZN(n1137) );
NAND2_X1 U804 ( .A1(G224), .A2(G898), .ZN(n1134) );
AND2_X1 U805 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
NAND3_X1 U806 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
NAND2_X1 U807 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
NAND3_X1 U808 ( .A1(n1145), .A2(n1144), .A3(n1143), .ZN(n1138) );
XNOR2_X1 U809 ( .A(KEYINPUT22), .B(G953), .ZN(n1143) );
NAND2_X1 U810 ( .A1(n1142), .A2(n1141), .ZN(n1145) );
XOR2_X1 U811 ( .A(n1146), .B(n1147), .Z(n1142) );
NOR2_X1 U812 ( .A1(KEYINPUT50), .A2(n1148), .ZN(n1146) );
NOR2_X1 U813 ( .A1(n1149), .A2(n1150), .ZN(G66) );
XOR2_X1 U814 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U815 ( .A1(n1104), .A2(n1153), .ZN(n1151) );
NOR2_X1 U816 ( .A1(n1149), .A2(n1154), .ZN(G63) );
XNOR2_X1 U817 ( .A(n1155), .B(n1156), .ZN(n1154) );
AND2_X1 U818 ( .A1(G478), .A2(n1157), .ZN(n1156) );
NOR3_X1 U819 ( .A1(n1158), .A2(n1149), .A3(n1159), .ZN(G60) );
NOR4_X1 U820 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1153), .ZN(n1159) );
NOR2_X1 U821 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
NOR2_X1 U822 ( .A1(KEYINPUT3), .A2(n1165), .ZN(n1163) );
NOR2_X1 U823 ( .A1(KEYINPUT3), .A2(n1166), .ZN(n1160) );
NOR2_X1 U824 ( .A1(n1167), .A2(n1168), .ZN(n1158) );
NOR2_X1 U825 ( .A1(n1164), .A2(n1165), .ZN(n1168) );
INV_X1 U826 ( .A(KEYINPUT52), .ZN(n1165) );
NOR2_X1 U827 ( .A1(n1162), .A2(n1153), .ZN(n1167) );
XNOR2_X1 U828 ( .A(n1169), .B(n1170), .ZN(G6) );
XNOR2_X1 U829 ( .A(G104), .B(KEYINPUT18), .ZN(n1170) );
NOR3_X1 U830 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(G57) );
NOR2_X1 U831 ( .A1(G101), .A2(n1174), .ZN(n1173) );
XOR2_X1 U832 ( .A(KEYINPUT51), .B(n1175), .Z(n1174) );
AND2_X1 U833 ( .A1(G101), .A2(n1175), .ZN(n1172) );
XOR2_X1 U834 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U835 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
NAND4_X1 U836 ( .A1(n1180), .A2(n1181), .A3(G472), .A4(n1062), .ZN(n1179) );
XOR2_X1 U837 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U838 ( .A(KEYINPUT36), .B(G902), .ZN(n1180) );
NAND2_X1 U839 ( .A1(n1184), .A2(n1185), .ZN(n1178) );
NAND3_X1 U840 ( .A1(n1186), .A2(n1187), .A3(G472), .ZN(n1185) );
NAND2_X1 U841 ( .A1(KEYINPUT36), .A2(n1153), .ZN(n1187) );
NAND2_X1 U842 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
INV_X1 U843 ( .A(KEYINPUT36), .ZN(n1189) );
NAND2_X1 U844 ( .A1(n1062), .A2(n1190), .ZN(n1188) );
XNOR2_X1 U845 ( .A(n1182), .B(n1183), .ZN(n1184) );
NAND2_X1 U846 ( .A1(KEYINPUT0), .A2(n1191), .ZN(n1182) );
NOR2_X1 U847 ( .A1(n1192), .A2(n1112), .ZN(n1171) );
XNOR2_X1 U848 ( .A(G952), .B(KEYINPUT47), .ZN(n1192) );
NOR2_X1 U849 ( .A1(n1149), .A2(n1193), .ZN(G54) );
XOR2_X1 U850 ( .A(n1194), .B(n1195), .Z(n1193) );
XOR2_X1 U851 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U852 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND2_X1 U853 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U854 ( .A(n1202), .B(KEYINPUT2), .Z(n1198) );
OR2_X1 U855 ( .A1(n1201), .A2(n1200), .ZN(n1202) );
XOR2_X1 U856 ( .A(n1203), .B(G134), .Z(n1200) );
XNOR2_X1 U857 ( .A(n1204), .B(n1205), .ZN(n1201) );
XNOR2_X1 U858 ( .A(n1206), .B(KEYINPUT23), .ZN(n1204) );
NAND2_X1 U859 ( .A1(n1207), .A2(n1208), .ZN(n1196) );
OR2_X1 U860 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U861 ( .A(n1211), .B(KEYINPUT16), .Z(n1207) );
NAND2_X1 U862 ( .A1(n1212), .A2(n1210), .ZN(n1211) );
XNOR2_X1 U863 ( .A(n1209), .B(KEYINPUT9), .ZN(n1212) );
AND2_X1 U864 ( .A1(G469), .A2(n1157), .ZN(n1194) );
NOR2_X1 U865 ( .A1(n1149), .A2(n1213), .ZN(G51) );
XOR2_X1 U866 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U867 ( .A1(KEYINPUT1), .A2(n1216), .ZN(n1215) );
XOR2_X1 U868 ( .A(n1217), .B(n1218), .Z(n1216) );
NOR2_X1 U869 ( .A1(G125), .A2(KEYINPUT46), .ZN(n1218) );
NAND2_X1 U870 ( .A1(n1157), .A2(n1103), .ZN(n1214) );
INV_X1 U871 ( .A(n1153), .ZN(n1157) );
NAND2_X1 U872 ( .A1(G902), .A2(n1062), .ZN(n1153) );
NAND3_X1 U873 ( .A1(n1130), .A2(n1219), .A3(n1220), .ZN(n1062) );
INV_X1 U874 ( .A(n1144), .ZN(n1220) );
NAND4_X1 U875 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1144) );
NOR4_X1 U876 ( .A1(n1225), .A2(n1226), .A3(n1169), .A4(n1057), .ZN(n1224) );
AND3_X1 U877 ( .A1(n1092), .A2(n1227), .A3(n1228), .ZN(n1057) );
AND3_X1 U878 ( .A1(n1228), .A2(n1227), .A3(n1093), .ZN(n1169) );
NOR3_X1 U879 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1223) );
NOR3_X1 U880 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
NOR4_X1 U881 ( .A1(n1235), .A2(n1078), .A3(n1236), .A4(n1237), .ZN(n1233) );
XNOR2_X1 U882 ( .A(n1238), .B(KEYINPUT13), .ZN(n1235) );
INV_X1 U883 ( .A(KEYINPUT17), .ZN(n1232) );
NOR2_X1 U884 ( .A1(KEYINPUT17), .A2(n1239), .ZN(n1230) );
NOR2_X1 U885 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR2_X1 U886 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
INV_X1 U887 ( .A(KEYINPUT13), .ZN(n1242) );
NOR2_X1 U888 ( .A1(KEYINPUT13), .A2(n1244), .ZN(n1240) );
NAND4_X1 U889 ( .A1(n1238), .A2(n1093), .A3(n1088), .A4(n1075), .ZN(n1244) );
NOR2_X1 U890 ( .A1(n1245), .A2(n1246), .ZN(n1229) );
XOR2_X1 U891 ( .A(KEYINPUT30), .B(n1131), .Z(n1219) );
AND4_X1 U892 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1131) );
NAND3_X1 U893 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1247) );
XNOR2_X1 U894 ( .A(n1254), .B(KEYINPUT49), .ZN(n1253) );
INV_X1 U895 ( .A(n1255), .ZN(n1251) );
NOR4_X1 U896 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1130) );
NOR2_X1 U897 ( .A1(n1112), .A2(G952), .ZN(n1149) );
XNOR2_X1 U898 ( .A(n1260), .B(n1257), .ZN(G48) );
AND3_X1 U899 ( .A1(n1093), .A2(n1254), .A3(n1261), .ZN(n1257) );
XOR2_X1 U900 ( .A(n1262), .B(n1263), .Z(G45) );
XNOR2_X1 U901 ( .A(KEYINPUT28), .B(n1264), .ZN(n1263) );
NAND3_X1 U902 ( .A1(n1265), .A2(n1266), .A3(KEYINPUT12), .ZN(n1262) );
NAND2_X1 U903 ( .A1(n1256), .A2(n1267), .ZN(n1266) );
INV_X1 U904 ( .A(KEYINPUT59), .ZN(n1267) );
NOR2_X1 U905 ( .A1(n1268), .A2(n1234), .ZN(n1256) );
NAND3_X1 U906 ( .A1(n1254), .A2(n1268), .A3(KEYINPUT59), .ZN(n1265) );
NAND4_X1 U907 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1268) );
NOR2_X1 U908 ( .A1(n1273), .A2(n1236), .ZN(n1272) );
XOR2_X1 U909 ( .A(G140), .B(n1258), .Z(G42) );
NOR3_X1 U910 ( .A1(n1081), .A2(n1273), .A3(n1255), .ZN(n1258) );
INV_X1 U911 ( .A(n1274), .ZN(n1081) );
XOR2_X1 U912 ( .A(G137), .B(n1259), .Z(G39) );
AND3_X1 U913 ( .A1(n1274), .A2(n1069), .A3(n1261), .ZN(n1259) );
XNOR2_X1 U914 ( .A(G134), .B(n1248), .ZN(G36) );
NAND2_X1 U915 ( .A1(n1275), .A2(n1092), .ZN(n1248) );
XNOR2_X1 U916 ( .A(G131), .B(n1249), .ZN(G33) );
NAND2_X1 U917 ( .A1(n1275), .A2(n1093), .ZN(n1249) );
AND4_X1 U918 ( .A1(n1274), .A2(n1088), .A3(n1083), .A4(n1270), .ZN(n1275) );
NOR2_X1 U919 ( .A1(n1079), .A2(n1098), .ZN(n1274) );
XNOR2_X1 U920 ( .A(G128), .B(n1250), .ZN(G30) );
NAND3_X1 U921 ( .A1(n1092), .A2(n1254), .A3(n1261), .ZN(n1250) );
AND4_X1 U922 ( .A1(n1089), .A2(n1083), .A3(n1276), .A4(n1270), .ZN(n1261) );
INV_X1 U923 ( .A(n1273), .ZN(n1083) );
XOR2_X1 U924 ( .A(n1277), .B(n1226), .Z(G3) );
AND3_X1 U925 ( .A1(n1069), .A2(n1228), .A3(n1088), .ZN(n1226) );
NAND2_X1 U926 ( .A1(KEYINPUT57), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U927 ( .A(n1121), .B(n1279), .ZN(G27) );
NOR2_X1 U928 ( .A1(n1245), .A2(n1255), .ZN(n1279) );
NAND4_X1 U929 ( .A1(n1093), .A2(n1276), .A3(n1280), .A4(n1270), .ZN(n1255) );
NAND2_X1 U930 ( .A1(n1064), .A2(n1281), .ZN(n1270) );
NAND3_X1 U931 ( .A1(G902), .A2(n1282), .A3(n1117), .ZN(n1281) );
NOR2_X1 U932 ( .A1(n1112), .A2(G900), .ZN(n1117) );
XNOR2_X1 U933 ( .A(n1283), .B(n1284), .ZN(G24) );
NOR3_X1 U934 ( .A1(n1285), .A2(n1234), .A3(n1246), .ZN(n1284) );
NAND4_X1 U935 ( .A1(n1227), .A2(n1271), .A3(n1269), .A4(n1286), .ZN(n1246) );
INV_X1 U936 ( .A(n1073), .ZN(n1227) );
NAND2_X1 U937 ( .A1(n1287), .A2(n1280), .ZN(n1073) );
XNOR2_X1 U938 ( .A(KEYINPUT33), .B(n1090), .ZN(n1287) );
XNOR2_X1 U939 ( .A(KEYINPUT56), .B(n1078), .ZN(n1285) );
XNOR2_X1 U940 ( .A(G119), .B(n1221), .ZN(G21) );
NAND4_X1 U941 ( .A1(n1089), .A2(n1075), .A3(n1288), .A4(n1069), .ZN(n1221) );
NOR2_X1 U942 ( .A1(n1238), .A2(n1090), .ZN(n1288) );
INV_X1 U943 ( .A(n1276), .ZN(n1090) );
INV_X1 U944 ( .A(n1280), .ZN(n1089) );
XOR2_X1 U945 ( .A(n1225), .B(n1289), .Z(G18) );
NOR2_X1 U946 ( .A1(KEYINPUT7), .A2(n1290), .ZN(n1289) );
AND2_X1 U947 ( .A1(n1291), .A2(n1092), .ZN(n1225) );
NOR2_X1 U948 ( .A1(n1269), .A2(n1292), .ZN(n1092) );
XNOR2_X1 U949 ( .A(G113), .B(n1243), .ZN(G15) );
NAND2_X1 U950 ( .A1(n1093), .A2(n1291), .ZN(n1243) );
NOR3_X1 U951 ( .A1(n1245), .A2(n1238), .A3(n1236), .ZN(n1291) );
INV_X1 U952 ( .A(n1088), .ZN(n1236) );
NOR2_X1 U953 ( .A1(n1280), .A2(n1276), .ZN(n1088) );
INV_X1 U954 ( .A(n1075), .ZN(n1245) );
NOR2_X1 U955 ( .A1(n1078), .A2(n1234), .ZN(n1075) );
INV_X1 U956 ( .A(n1252), .ZN(n1078) );
NOR2_X1 U957 ( .A1(n1084), .A2(n1097), .ZN(n1252) );
INV_X1 U958 ( .A(n1085), .ZN(n1097) );
XNOR2_X1 U959 ( .A(n1100), .B(KEYINPUT21), .ZN(n1084) );
INV_X1 U960 ( .A(n1237), .ZN(n1093) );
NAND2_X1 U961 ( .A1(n1292), .A2(n1269), .ZN(n1237) );
INV_X1 U962 ( .A(n1271), .ZN(n1292) );
XNOR2_X1 U963 ( .A(G110), .B(n1222), .ZN(G12) );
NAND4_X1 U964 ( .A1(n1069), .A2(n1228), .A3(n1276), .A4(n1280), .ZN(n1222) );
XOR2_X1 U965 ( .A(G472), .B(n1293), .Z(n1280) );
NOR2_X1 U966 ( .A1(n1107), .A2(KEYINPUT4), .ZN(n1293) );
AND2_X1 U967 ( .A1(n1294), .A2(n1190), .ZN(n1107) );
XOR2_X1 U968 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U969 ( .A(G101), .B(n1177), .ZN(n1296) );
NAND2_X1 U970 ( .A1(n1297), .A2(G210), .ZN(n1177) );
XNOR2_X1 U971 ( .A(n1191), .B(n1183), .ZN(n1295) );
XOR2_X1 U972 ( .A(G113), .B(n1298), .Z(n1183) );
XNOR2_X1 U973 ( .A(n1299), .B(n1300), .ZN(n1191) );
XOR2_X1 U974 ( .A(n1106), .B(n1104), .Z(n1276) );
NAND2_X1 U975 ( .A1(G217), .A2(n1301), .ZN(n1104) );
OR2_X1 U976 ( .A1(n1152), .A2(G902), .ZN(n1106) );
XNOR2_X1 U977 ( .A(n1302), .B(n1303), .ZN(n1152) );
XNOR2_X1 U978 ( .A(n1304), .B(n1305), .ZN(n1303) );
NOR2_X1 U979 ( .A1(G119), .A2(KEYINPUT58), .ZN(n1305) );
NAND2_X1 U980 ( .A1(KEYINPUT34), .A2(n1260), .ZN(n1304) );
XOR2_X1 U981 ( .A(n1306), .B(n1307), .Z(n1302) );
NOR3_X1 U982 ( .A1(n1308), .A2(KEYINPUT38), .A3(n1309), .ZN(n1307) );
INV_X1 U983 ( .A(G221), .ZN(n1309) );
XOR2_X1 U984 ( .A(n1310), .B(n1311), .Z(n1306) );
XNOR2_X1 U985 ( .A(G128), .B(n1312), .ZN(n1311) );
XNOR2_X1 U986 ( .A(KEYINPUT60), .B(KEYINPUT45), .ZN(n1312) );
XNOR2_X1 U987 ( .A(n1209), .B(n1313), .ZN(n1310) );
XNOR2_X1 U988 ( .A(n1121), .B(n1314), .ZN(n1313) );
NOR3_X1 U989 ( .A1(n1234), .A2(n1238), .A3(n1273), .ZN(n1228) );
NAND2_X1 U990 ( .A1(n1100), .A2(n1085), .ZN(n1273) );
NAND2_X1 U991 ( .A1(G221), .A2(n1301), .ZN(n1085) );
NAND2_X1 U992 ( .A1(G234), .A2(n1190), .ZN(n1301) );
XNOR2_X1 U993 ( .A(n1315), .B(G469), .ZN(n1100) );
NAND2_X1 U994 ( .A1(n1316), .A2(n1190), .ZN(n1315) );
XOR2_X1 U995 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U996 ( .A(n1205), .B(n1209), .ZN(n1318) );
XOR2_X1 U997 ( .A(G110), .B(n1119), .Z(n1209) );
XNOR2_X1 U998 ( .A(n1319), .B(n1126), .ZN(n1205) );
NOR2_X1 U999 ( .A1(KEYINPUT31), .A2(n1320), .ZN(n1126) );
NAND2_X1 U1000 ( .A1(n1321), .A2(n1322), .ZN(n1319) );
NAND2_X1 U1001 ( .A1(n1323), .A2(n1278), .ZN(n1322) );
XOR2_X1 U1002 ( .A(KEYINPUT61), .B(n1324), .Z(n1321) );
NOR2_X1 U1003 ( .A1(n1323), .A2(n1278), .ZN(n1324) );
XOR2_X1 U1004 ( .A(n1325), .B(n1326), .Z(n1323) );
NOR2_X1 U1005 ( .A1(G104), .A2(n1327), .ZN(n1326) );
XNOR2_X1 U1006 ( .A(KEYINPUT29), .B(KEYINPUT20), .ZN(n1327) );
XNOR2_X1 U1007 ( .A(G107), .B(KEYINPUT6), .ZN(n1325) );
XOR2_X1 U1008 ( .A(n1299), .B(n1210), .Z(n1317) );
AND2_X1 U1009 ( .A1(G227), .A2(n1112), .ZN(n1210) );
XNOR2_X1 U1010 ( .A(n1124), .B(G134), .ZN(n1299) );
XOR2_X1 U1011 ( .A(n1203), .B(n1328), .Z(n1124) );
INV_X1 U1012 ( .A(n1206), .ZN(n1328) );
XNOR2_X1 U1013 ( .A(G131), .B(n1314), .ZN(n1203) );
XOR2_X1 U1014 ( .A(G137), .B(KEYINPUT35), .Z(n1314) );
INV_X1 U1015 ( .A(n1286), .ZN(n1238) );
NAND2_X1 U1016 ( .A1(n1329), .A2(n1330), .ZN(n1286) );
NAND3_X1 U1017 ( .A1(n1331), .A2(n1282), .A3(G902), .ZN(n1330) );
INV_X1 U1018 ( .A(n1141), .ZN(n1331) );
NAND2_X1 U1019 ( .A1(G953), .A2(n1332), .ZN(n1141) );
XOR2_X1 U1020 ( .A(KEYINPUT11), .B(G898), .Z(n1332) );
XNOR2_X1 U1021 ( .A(KEYINPUT27), .B(n1064), .ZN(n1329) );
NAND3_X1 U1022 ( .A1(n1282), .A2(n1112), .A3(G952), .ZN(n1064) );
NAND2_X1 U1023 ( .A1(G237), .A2(G234), .ZN(n1282) );
INV_X1 U1024 ( .A(n1254), .ZN(n1234) );
NOR2_X1 U1025 ( .A1(n1333), .A2(n1098), .ZN(n1254) );
INV_X1 U1026 ( .A(n1077), .ZN(n1098) );
NAND2_X1 U1027 ( .A1(n1334), .A2(G214), .ZN(n1077) );
XOR2_X1 U1028 ( .A(n1335), .B(KEYINPUT10), .Z(n1334) );
INV_X1 U1029 ( .A(n1079), .ZN(n1333) );
XNOR2_X1 U1030 ( .A(n1101), .B(n1103), .ZN(n1079) );
AND2_X1 U1031 ( .A1(G210), .A2(n1335), .ZN(n1103) );
NAND2_X1 U1032 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
INV_X1 U1033 ( .A(G237), .ZN(n1337) );
XNOR2_X1 U1034 ( .A(KEYINPUT44), .B(n1190), .ZN(n1336) );
NAND2_X1 U1035 ( .A1(n1338), .A2(n1190), .ZN(n1101) );
XNOR2_X1 U1036 ( .A(n1217), .B(n1121), .ZN(n1338) );
XOR2_X1 U1037 ( .A(n1339), .B(n1340), .Z(n1217) );
XNOR2_X1 U1038 ( .A(n1206), .B(n1341), .ZN(n1340) );
XOR2_X1 U1039 ( .A(n1342), .B(n1300), .Z(n1341) );
NOR2_X1 U1040 ( .A1(KEYINPUT42), .A2(n1343), .ZN(n1300) );
XNOR2_X1 U1041 ( .A(n1320), .B(KEYINPUT32), .ZN(n1343) );
XOR2_X1 U1042 ( .A(G128), .B(KEYINPUT26), .Z(n1320) );
NAND2_X1 U1043 ( .A1(G224), .A2(n1112), .ZN(n1342) );
XOR2_X1 U1044 ( .A(G143), .B(n1344), .Z(n1206) );
XNOR2_X1 U1045 ( .A(KEYINPUT14), .B(n1260), .ZN(n1344) );
XOR2_X1 U1046 ( .A(n1345), .B(n1147), .Z(n1339) );
XNOR2_X1 U1047 ( .A(n1346), .B(G122), .ZN(n1147) );
INV_X1 U1048 ( .A(G110), .ZN(n1346) );
NAND2_X1 U1049 ( .A1(n1347), .A2(n1348), .ZN(n1345) );
NAND2_X1 U1050 ( .A1(KEYINPUT15), .A2(n1148), .ZN(n1348) );
XNOR2_X1 U1051 ( .A(n1349), .B(n1350), .ZN(n1148) );
XOR2_X1 U1052 ( .A(n1351), .B(n1352), .Z(n1350) );
NAND3_X1 U1053 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1347) );
INV_X1 U1054 ( .A(KEYINPUT15), .ZN(n1355) );
XOR2_X1 U1055 ( .A(G104), .B(n1352), .Z(n1354) );
XNOR2_X1 U1056 ( .A(G107), .B(n1278), .ZN(n1352) );
INV_X1 U1057 ( .A(G101), .ZN(n1278) );
XNOR2_X1 U1058 ( .A(G113), .B(n1349), .ZN(n1353) );
NAND2_X1 U1059 ( .A1(n1356), .A2(n1357), .ZN(n1349) );
OR2_X1 U1060 ( .A1(n1298), .A2(KEYINPUT8), .ZN(n1357) );
XOR2_X1 U1061 ( .A(G116), .B(G119), .Z(n1298) );
NAND3_X1 U1062 ( .A1(G116), .A2(n1358), .A3(KEYINPUT8), .ZN(n1356) );
INV_X1 U1063 ( .A(G119), .ZN(n1358) );
NOR2_X1 U1064 ( .A1(n1271), .A2(n1269), .ZN(n1069) );
XOR2_X1 U1065 ( .A(n1359), .B(n1162), .Z(n1269) );
INV_X1 U1066 ( .A(G475), .ZN(n1162) );
NAND2_X1 U1067 ( .A1(n1360), .A2(n1190), .ZN(n1359) );
XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n1166), .ZN(n1360) );
INV_X1 U1069 ( .A(n1164), .ZN(n1166) );
XNOR2_X1 U1070 ( .A(n1361), .B(n1362), .ZN(n1164) );
XOR2_X1 U1071 ( .A(n1363), .B(n1351), .Z(n1362) );
XOR2_X1 U1072 ( .A(G104), .B(G113), .Z(n1351) );
NOR2_X1 U1073 ( .A1(KEYINPUT62), .A2(n1283), .ZN(n1363) );
INV_X1 U1074 ( .A(G122), .ZN(n1283) );
XOR2_X1 U1075 ( .A(n1364), .B(n1365), .Z(n1361) );
XOR2_X1 U1076 ( .A(G131), .B(n1366), .Z(n1365) );
NOR2_X1 U1077 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
XOR2_X1 U1078 ( .A(n1369), .B(KEYINPUT5), .Z(n1368) );
NAND2_X1 U1079 ( .A1(G146), .A2(n1370), .ZN(n1369) );
XOR2_X1 U1080 ( .A(KEYINPUT37), .B(n1371), .Z(n1370) );
AND2_X1 U1081 ( .A1(n1260), .A2(n1371), .ZN(n1367) );
XOR2_X1 U1082 ( .A(n1119), .B(n1372), .Z(n1371) );
NOR2_X1 U1083 ( .A1(KEYINPUT24), .A2(n1121), .ZN(n1372) );
INV_X1 U1084 ( .A(G125), .ZN(n1121) );
XOR2_X1 U1085 ( .A(G140), .B(KEYINPUT41), .Z(n1119) );
INV_X1 U1086 ( .A(G146), .ZN(n1260) );
NAND2_X1 U1087 ( .A1(n1373), .A2(KEYINPUT43), .ZN(n1364) );
XNOR2_X1 U1088 ( .A(n1374), .B(n1264), .ZN(n1373) );
INV_X1 U1089 ( .A(G143), .ZN(n1264) );
NAND2_X1 U1090 ( .A1(n1297), .A2(G214), .ZN(n1374) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1297) );
XNOR2_X1 U1092 ( .A(n1375), .B(G478), .ZN(n1271) );
NAND2_X1 U1093 ( .A1(n1155), .A2(n1190), .ZN(n1375) );
INV_X1 U1094 ( .A(G902), .ZN(n1190) );
XNOR2_X1 U1095 ( .A(n1376), .B(n1377), .ZN(n1155) );
NOR2_X1 U1096 ( .A1(KEYINPUT48), .A2(n1378), .ZN(n1377) );
XOR2_X1 U1097 ( .A(n1379), .B(n1380), .Z(n1378) );
XOR2_X1 U1098 ( .A(n1381), .B(n1382), .Z(n1380) );
XNOR2_X1 U1099 ( .A(n1290), .B(G107), .ZN(n1382) );
INV_X1 U1100 ( .A(G116), .ZN(n1290) );
NAND2_X1 U1101 ( .A1(KEYINPUT19), .A2(G143), .ZN(n1381) );
XOR2_X1 U1102 ( .A(n1383), .B(n1384), .Z(n1379) );
XNOR2_X1 U1103 ( .A(KEYINPUT25), .B(n1128), .ZN(n1384) );
INV_X1 U1104 ( .A(G134), .ZN(n1128) );
XNOR2_X1 U1105 ( .A(G122), .B(G128), .ZN(n1383) );
NAND2_X1 U1106 ( .A1(G217), .A2(n1385), .ZN(n1376) );
INV_X1 U1107 ( .A(n1308), .ZN(n1385) );
NAND2_X1 U1108 ( .A1(G234), .A2(n1112), .ZN(n1308) );
INV_X1 U1109 ( .A(G953), .ZN(n1112) );
endmodule


