//Key = 1111100101001100101000100111110100000101110010000101111100001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;

XNOR2_X1 U704 ( .A(G107), .B(n959), .ZN(G9) );
NAND3_X1 U705 ( .A1(n960), .A2(n961), .A3(n962), .ZN(G75) );
NOR3_X1 U706 ( .A1(n963), .A2(G953), .A3(n964), .ZN(n962) );
NOR4_X1 U707 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(n964) );
NOR2_X1 U708 ( .A1(n969), .A2(n970), .ZN(n967) );
NAND3_X1 U709 ( .A1(n971), .A2(n972), .A3(n973), .ZN(n965) );
NAND2_X1 U710 ( .A1(KEYINPUT9), .A2(n974), .ZN(n972) );
OR3_X1 U711 ( .A1(n975), .A2(KEYINPUT9), .A3(n974), .ZN(n971) );
NOR4_X1 U712 ( .A1(n976), .A2(n977), .A3(n978), .A4(n979), .ZN(n963) );
XNOR2_X1 U713 ( .A(G469), .B(n980), .ZN(n979) );
NOR2_X1 U714 ( .A1(n981), .A2(KEYINPUT17), .ZN(n980) );
NOR2_X1 U715 ( .A1(n982), .A2(n983), .ZN(n978) );
XNOR2_X1 U716 ( .A(KEYINPUT3), .B(n984), .ZN(n983) );
XNOR2_X1 U717 ( .A(n985), .B(KEYINPUT13), .ZN(n982) );
NAND3_X1 U718 ( .A1(n986), .A2(n987), .A3(n988), .ZN(n977) );
NAND4_X1 U719 ( .A1(n989), .A2(n990), .A3(n991), .A4(n992), .ZN(n976) );
XNOR2_X1 U720 ( .A(n993), .B(n994), .ZN(n990) );
NAND2_X1 U721 ( .A1(KEYINPUT31), .A2(n995), .ZN(n993) );
XNOR2_X1 U722 ( .A(n996), .B(n997), .ZN(n989) );
NAND3_X1 U723 ( .A1(n998), .A2(n999), .A3(n973), .ZN(n961) );
INV_X1 U724 ( .A(n1000), .ZN(n973) );
NAND2_X1 U725 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NAND3_X1 U726 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
NAND3_X1 U727 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1004) );
NAND2_X1 U728 ( .A1(KEYINPUT23), .A2(n988), .ZN(n1007) );
OR3_X1 U729 ( .A1(n1009), .A2(KEYINPUT23), .A3(n988), .ZN(n1006) );
NAND2_X1 U730 ( .A1(n1010), .A2(n1011), .ZN(n1001) );
NAND2_X1 U731 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U732 ( .A1(n1005), .A2(n1014), .ZN(n1013) );
OR2_X1 U733 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U734 ( .A1(n1003), .A2(n1017), .ZN(n1012) );
NAND2_X1 U735 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
OR2_X1 U736 ( .A1(n986), .A2(n1020), .ZN(n1019) );
XOR2_X1 U737 ( .A(n1021), .B(n1022), .Z(G72) );
XOR2_X1 U738 ( .A(n1023), .B(n1024), .Z(n1022) );
NOR3_X1 U739 ( .A1(n1025), .A2(KEYINPUT48), .A3(n1026), .ZN(n1024) );
NOR2_X1 U740 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XOR2_X1 U741 ( .A(n1029), .B(KEYINPUT53), .Z(n1027) );
XNOR2_X1 U742 ( .A(KEYINPUT38), .B(n1030), .ZN(n1025) );
NAND3_X1 U743 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1023) );
XOR2_X1 U744 ( .A(n1034), .B(KEYINPUT15), .Z(n1033) );
NAND2_X1 U745 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
XNOR2_X1 U746 ( .A(n1037), .B(KEYINPUT24), .ZN(n1035) );
OR2_X1 U747 ( .A1(n1036), .A2(n1038), .ZN(n1032) );
XOR2_X1 U748 ( .A(n1039), .B(n1040), .Z(n1036) );
NAND2_X1 U749 ( .A1(G953), .A2(n1041), .ZN(n1031) );
NAND2_X1 U750 ( .A1(G953), .A2(n1042), .ZN(n1021) );
NAND2_X1 U751 ( .A1(G900), .A2(G227), .ZN(n1042) );
XOR2_X1 U752 ( .A(n1043), .B(n1044), .Z(G69) );
XOR2_X1 U753 ( .A(n1045), .B(n1046), .Z(n1044) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
XNOR2_X1 U755 ( .A(KEYINPUT60), .B(n1030), .ZN(n1048) );
AND2_X1 U756 ( .A1(G224), .A2(G898), .ZN(n1047) );
NAND2_X1 U757 ( .A1(n1030), .A2(n1049), .ZN(n1045) );
NAND3_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
XOR2_X1 U759 ( .A(n1053), .B(KEYINPUT46), .Z(n1052) );
XNOR2_X1 U760 ( .A(KEYINPUT6), .B(n1054), .ZN(n1051) );
OR3_X1 U761 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1043) );
XNOR2_X1 U762 ( .A(n1058), .B(KEYINPUT32), .ZN(n1057) );
NAND2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U764 ( .A1(n1061), .A2(n1062), .ZN(G66) );
XOR2_X1 U765 ( .A(n1063), .B(n1064), .Z(n1062) );
NOR2_X1 U766 ( .A1(n997), .A2(n1065), .ZN(n1064) );
NAND2_X1 U767 ( .A1(KEYINPUT0), .A2(n1066), .ZN(n1063) );
NOR2_X1 U768 ( .A1(n1061), .A2(n1067), .ZN(G63) );
XOR2_X1 U769 ( .A(n1068), .B(n1069), .Z(n1067) );
AND2_X1 U770 ( .A1(G478), .A2(n1070), .ZN(n1069) );
NOR2_X1 U771 ( .A1(n1061), .A2(n1071), .ZN(G60) );
XOR2_X1 U772 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U773 ( .A1(n984), .A2(n1065), .ZN(n1072) );
XOR2_X1 U774 ( .A(n1074), .B(n1075), .Z(G6) );
XOR2_X1 U775 ( .A(KEYINPUT62), .B(G104), .Z(n1075) );
NAND3_X1 U776 ( .A1(n1076), .A2(n1077), .A3(KEYINPUT55), .ZN(n1074) );
NOR2_X1 U777 ( .A1(n1061), .A2(n1078), .ZN(G57) );
XNOR2_X1 U778 ( .A(n1079), .B(n1080), .ZN(n1078) );
NAND2_X1 U779 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U780 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
INV_X1 U781 ( .A(n1085), .ZN(n1083) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
XOR2_X1 U783 ( .A(n1084), .B(KEYINPUT54), .Z(n1086) );
NAND2_X1 U784 ( .A1(n1070), .A2(G472), .ZN(n1084) );
XNOR2_X1 U785 ( .A(n1087), .B(n1088), .ZN(n1085) );
NOR2_X1 U786 ( .A1(KEYINPUT30), .A2(n1089), .ZN(n1088) );
NOR2_X1 U787 ( .A1(n1061), .A2(n1090), .ZN(G54) );
XOR2_X1 U788 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U789 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U790 ( .A1(n1095), .A2(n1065), .ZN(n1094) );
NOR2_X1 U791 ( .A1(KEYINPUT61), .A2(n1096), .ZN(n1093) );
XOR2_X1 U792 ( .A(n1039), .B(n1097), .Z(n1096) );
NAND2_X1 U793 ( .A1(n1098), .A2(n1099), .ZN(n1091) );
OR2_X1 U794 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XOR2_X1 U795 ( .A(n1102), .B(KEYINPUT21), .Z(n1098) );
NAND2_X1 U796 ( .A1(n1100), .A2(n1101), .ZN(n1102) );
XNOR2_X1 U797 ( .A(n1103), .B(KEYINPUT14), .ZN(n1100) );
NOR3_X1 U798 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(G51) );
NOR3_X1 U799 ( .A1(n1107), .A2(G953), .A3(G952), .ZN(n1106) );
AND2_X1 U800 ( .A1(n1107), .A2(n1061), .ZN(n1105) );
NOR2_X1 U801 ( .A1(n1030), .A2(G952), .ZN(n1061) );
INV_X1 U802 ( .A(KEYINPUT11), .ZN(n1107) );
NOR2_X1 U803 ( .A1(n1108), .A2(n1109), .ZN(n1104) );
XOR2_X1 U804 ( .A(n1110), .B(KEYINPUT26), .Z(n1109) );
NAND2_X1 U805 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
OR2_X1 U806 ( .A1(n1065), .A2(n994), .ZN(n1112) );
NOR3_X1 U807 ( .A1(n1065), .A2(n1111), .A3(n994), .ZN(n1108) );
XOR2_X1 U808 ( .A(n1113), .B(n1114), .Z(n1111) );
NAND2_X1 U809 ( .A1(n1115), .A2(KEYINPUT39), .ZN(n1113) );
XOR2_X1 U810 ( .A(n1116), .B(KEYINPUT35), .Z(n1115) );
INV_X1 U811 ( .A(n1070), .ZN(n1065) );
NOR2_X1 U812 ( .A1(n1117), .A2(n960), .ZN(n1070) );
AND4_X1 U813 ( .A1(n1029), .A2(n1053), .A3(n1050), .A4(n1118), .ZN(n960) );
NOR2_X1 U814 ( .A1(n1028), .A2(n1054), .ZN(n1118) );
NAND3_X1 U815 ( .A1(n1119), .A2(n959), .A3(n1120), .ZN(n1054) );
NAND2_X1 U816 ( .A1(n1077), .A2(n1121), .ZN(n1120) );
OR2_X1 U817 ( .A1(n1122), .A2(n1076), .ZN(n1121) );
NOR2_X1 U818 ( .A1(n1123), .A2(n968), .ZN(n1076) );
NAND3_X1 U819 ( .A1(n969), .A2(n1003), .A3(n1077), .ZN(n959) );
NAND4_X1 U820 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1028) );
NOR4_X1 U821 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1127) );
INV_X1 U822 ( .A(n1132), .ZN(n1131) );
NAND4_X1 U823 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n975), .ZN(n1126) );
XNOR2_X1 U824 ( .A(n1005), .B(KEYINPUT44), .ZN(n1133) );
AND3_X1 U825 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1050) );
NAND3_X1 U826 ( .A1(n1016), .A2(n969), .A3(n1139), .ZN(n1138) );
XNOR2_X1 U827 ( .A(G146), .B(n1124), .ZN(G48) );
NAND4_X1 U828 ( .A1(n1134), .A2(n975), .A3(n1140), .A4(n1141), .ZN(n1124) );
XNOR2_X1 U829 ( .A(G143), .B(n1029), .ZN(G45) );
NAND4_X1 U830 ( .A1(n1142), .A2(n1140), .A3(n1143), .A4(n1144), .ZN(n1029) );
XNOR2_X1 U831 ( .A(G140), .B(n1145), .ZN(G42) );
NAND3_X1 U832 ( .A1(n1135), .A2(n1134), .A3(n970), .ZN(n1145) );
XNOR2_X1 U833 ( .A(G137), .B(n1125), .ZN(G39) );
NAND4_X1 U834 ( .A1(n1005), .A2(n1134), .A3(n998), .A4(n1141), .ZN(n1125) );
XOR2_X1 U835 ( .A(G134), .B(n1130), .Z(G36) );
AND3_X1 U836 ( .A1(n1142), .A2(n969), .A3(n1005), .ZN(n1130) );
INV_X1 U837 ( .A(n974), .ZN(n1005) );
XNOR2_X1 U838 ( .A(G131), .B(n1146), .ZN(G33) );
NAND2_X1 U839 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U840 ( .A1(KEYINPUT59), .A2(n1129), .ZN(n1148) );
OR2_X1 U841 ( .A1(KEYINPUT42), .A2(n1129), .ZN(n1147) );
AND2_X1 U842 ( .A1(n970), .A2(n1142), .ZN(n1129) );
NOR3_X1 U843 ( .A1(n1008), .A2(n1149), .A3(n1150), .ZN(n1142) );
NOR2_X1 U844 ( .A1(n974), .A2(n1123), .ZN(n970) );
NAND2_X1 U845 ( .A1(n1151), .A2(n986), .ZN(n974) );
XOR2_X1 U846 ( .A(n1128), .B(n1152), .Z(G30) );
NOR2_X1 U847 ( .A1(KEYINPUT43), .A2(n1153), .ZN(n1152) );
AND4_X1 U848 ( .A1(n1134), .A2(n969), .A3(n1140), .A4(n1141), .ZN(n1128) );
NOR3_X1 U849 ( .A1(n1008), .A2(n1149), .A3(n1154), .ZN(n1134) );
XNOR2_X1 U850 ( .A(G101), .B(n1119), .ZN(G3) );
NAND3_X1 U851 ( .A1(n998), .A2(n1077), .A3(n1016), .ZN(n1119) );
XNOR2_X1 U852 ( .A(G125), .B(n1132), .ZN(G27) );
NAND4_X1 U853 ( .A1(n1010), .A2(n1015), .A3(n1155), .A4(n975), .ZN(n1132) );
NOR2_X1 U854 ( .A1(n1149), .A2(n1018), .ZN(n1155) );
AND2_X1 U855 ( .A1(n1000), .A2(n1156), .ZN(n1149) );
NAND4_X1 U856 ( .A1(G902), .A2(G953), .A3(n1157), .A4(n1041), .ZN(n1156) );
INV_X1 U857 ( .A(G900), .ZN(n1041) );
INV_X1 U858 ( .A(n966), .ZN(n1010) );
XNOR2_X1 U859 ( .A(G122), .B(n1136), .ZN(G24) );
NAND4_X1 U860 ( .A1(n1139), .A2(n1003), .A3(n1143), .A4(n1144), .ZN(n1136) );
INV_X1 U861 ( .A(n968), .ZN(n1003) );
NAND2_X1 U862 ( .A1(n1158), .A2(n1135), .ZN(n968) );
INV_X1 U863 ( .A(n1141), .ZN(n1135) );
XNOR2_X1 U864 ( .A(G119), .B(n1137), .ZN(G21) );
NAND4_X1 U865 ( .A1(n1139), .A2(n998), .A3(n1159), .A4(n1141), .ZN(n1137) );
INV_X1 U866 ( .A(n1154), .ZN(n1159) );
XNOR2_X1 U867 ( .A(G116), .B(n1160), .ZN(G18) );
NAND4_X1 U868 ( .A1(KEYINPUT2), .A2(n1139), .A3(n1016), .A4(n969), .ZN(n1160) );
AND2_X1 U869 ( .A1(n1161), .A2(n1143), .ZN(n969) );
XNOR2_X1 U870 ( .A(G113), .B(n1053), .ZN(G15) );
NAND3_X1 U871 ( .A1(n975), .A2(n1016), .A3(n1139), .ZN(n1053) );
NOR2_X1 U872 ( .A1(n966), .A2(n1162), .ZN(n1139) );
NAND2_X1 U873 ( .A1(n1163), .A2(n988), .ZN(n966) );
INV_X1 U874 ( .A(n1009), .ZN(n1163) );
INV_X1 U875 ( .A(n1150), .ZN(n1016) );
NAND2_X1 U876 ( .A1(n1158), .A2(n1141), .ZN(n1150) );
XNOR2_X1 U877 ( .A(KEYINPUT51), .B(n1154), .ZN(n1158) );
INV_X1 U878 ( .A(n1123), .ZN(n975) );
NAND2_X1 U879 ( .A1(n991), .A2(n1144), .ZN(n1123) );
XNOR2_X1 U880 ( .A(G110), .B(n1164), .ZN(G12) );
NAND3_X1 U881 ( .A1(n1122), .A2(n1077), .A3(KEYINPUT22), .ZN(n1164) );
NOR2_X1 U882 ( .A1(n1162), .A2(n1008), .ZN(n1077) );
NAND2_X1 U883 ( .A1(n1009), .A2(n988), .ZN(n1008) );
NAND2_X1 U884 ( .A1(G221), .A2(n1165), .ZN(n988) );
XNOR2_X1 U885 ( .A(n981), .B(n1095), .ZN(n1009) );
INV_X1 U886 ( .A(G469), .ZN(n1095) );
AND2_X1 U887 ( .A1(n1166), .A2(n1117), .ZN(n981) );
XOR2_X1 U888 ( .A(n1103), .B(n1167), .Z(n1166) );
XNOR2_X1 U889 ( .A(n1168), .B(n1101), .ZN(n1167) );
NAND2_X1 U890 ( .A1(G227), .A2(n1030), .ZN(n1101) );
NAND2_X1 U891 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
OR2_X1 U892 ( .A1(n1039), .A2(n1097), .ZN(n1170) );
XOR2_X1 U893 ( .A(n1171), .B(KEYINPUT10), .Z(n1169) );
NAND2_X1 U894 ( .A1(n1097), .A2(n1039), .ZN(n1171) );
XOR2_X1 U895 ( .A(n1040), .B(n1172), .Z(n1097) );
XOR2_X1 U896 ( .A(G104), .B(n1173), .Z(n1172) );
XNOR2_X1 U897 ( .A(G146), .B(n1174), .ZN(n1040) );
XNOR2_X1 U898 ( .A(G140), .B(G110), .ZN(n1103) );
NAND2_X1 U899 ( .A1(n1140), .A2(n1175), .ZN(n1162) );
NAND2_X1 U900 ( .A1(n1000), .A2(n1176), .ZN(n1175) );
NAND3_X1 U901 ( .A1(n1056), .A2(n1157), .A3(G902), .ZN(n1176) );
NOR2_X1 U902 ( .A1(n1030), .A2(G898), .ZN(n1056) );
NAND3_X1 U903 ( .A1(n1157), .A2(n1030), .A3(G952), .ZN(n1000) );
NAND2_X1 U904 ( .A1(G237), .A2(G234), .ZN(n1157) );
INV_X1 U905 ( .A(n1018), .ZN(n1140) );
NAND2_X1 U906 ( .A1(n1020), .A2(n986), .ZN(n1018) );
NAND2_X1 U907 ( .A1(G214), .A2(n1177), .ZN(n986) );
INV_X1 U908 ( .A(n1151), .ZN(n1020) );
XNOR2_X1 U909 ( .A(n1178), .B(n994), .ZN(n1151) );
NAND2_X1 U910 ( .A1(G210), .A2(n1177), .ZN(n994) );
NAND2_X1 U911 ( .A1(n1179), .A2(n1117), .ZN(n1177) );
XNOR2_X1 U912 ( .A(n995), .B(KEYINPUT45), .ZN(n1178) );
AND2_X1 U913 ( .A1(n1180), .A2(n1117), .ZN(n995) );
XNOR2_X1 U914 ( .A(n1114), .B(n1181), .ZN(n1180) );
XNOR2_X1 U915 ( .A(KEYINPUT49), .B(n1116), .ZN(n1181) );
NAND2_X1 U916 ( .A1(n1182), .A2(n1183), .ZN(n1116) );
NAND2_X1 U917 ( .A1(n1059), .A2(n1184), .ZN(n1183) );
NAND2_X1 U918 ( .A1(KEYINPUT52), .A2(n1185), .ZN(n1184) );
INV_X1 U919 ( .A(n1060), .ZN(n1185) );
NAND2_X1 U920 ( .A1(n1055), .A2(KEYINPUT52), .ZN(n1182) );
NOR2_X1 U921 ( .A1(n1060), .A2(n1059), .ZN(n1055) );
XNOR2_X1 U922 ( .A(G122), .B(n1186), .ZN(n1059) );
NOR2_X1 U923 ( .A1(KEYINPUT20), .A2(n1187), .ZN(n1186) );
INV_X1 U924 ( .A(G110), .ZN(n1187) );
XNOR2_X1 U925 ( .A(n1188), .B(n1189), .ZN(n1060) );
XNOR2_X1 U926 ( .A(G116), .B(n1190), .ZN(n1189) );
XNOR2_X1 U927 ( .A(KEYINPUT50), .B(KEYINPUT37), .ZN(n1190) );
XOR2_X1 U928 ( .A(n1191), .B(n1173), .Z(n1188) );
XNOR2_X1 U929 ( .A(n1192), .B(G107), .ZN(n1173) );
INV_X1 U930 ( .A(G101), .ZN(n1192) );
XOR2_X1 U931 ( .A(n1193), .B(n1194), .Z(n1191) );
NAND2_X1 U932 ( .A1(KEYINPUT7), .A2(n1195), .ZN(n1193) );
XNOR2_X1 U933 ( .A(n1196), .B(n1197), .ZN(n1114) );
AND2_X1 U934 ( .A1(n1030), .A2(G224), .ZN(n1197) );
XNOR2_X1 U935 ( .A(n1089), .B(n1198), .ZN(n1196) );
INV_X1 U936 ( .A(G125), .ZN(n1198) );
AND2_X1 U937 ( .A1(n1015), .A2(n998), .ZN(n1122) );
AND2_X1 U938 ( .A1(n1161), .A2(n991), .ZN(n998) );
INV_X1 U939 ( .A(n1143), .ZN(n991) );
XNOR2_X1 U940 ( .A(n1199), .B(G478), .ZN(n1143) );
NAND2_X1 U941 ( .A1(n1200), .A2(n1117), .ZN(n1199) );
XOR2_X1 U942 ( .A(n1068), .B(KEYINPUT25), .Z(n1200) );
XOR2_X1 U943 ( .A(n1201), .B(n1202), .Z(n1068) );
XNOR2_X1 U944 ( .A(n1203), .B(n1204), .ZN(n1202) );
XNOR2_X1 U945 ( .A(n1205), .B(n1206), .ZN(n1204) );
NOR2_X1 U946 ( .A1(KEYINPUT47), .A2(n1207), .ZN(n1206) );
INV_X1 U947 ( .A(G107), .ZN(n1207) );
NOR2_X1 U948 ( .A1(KEYINPUT34), .A2(n1174), .ZN(n1205) );
XNOR2_X1 U949 ( .A(n1153), .B(n1208), .ZN(n1174) );
XOR2_X1 U950 ( .A(n1209), .B(n1210), .Z(n1201) );
XOR2_X1 U951 ( .A(G122), .B(G116), .Z(n1210) );
NAND3_X1 U952 ( .A1(G234), .A2(n1030), .A3(G217), .ZN(n1209) );
XOR2_X1 U953 ( .A(n1144), .B(KEYINPUT12), .Z(n1161) );
NAND2_X1 U954 ( .A1(n987), .A2(n1211), .ZN(n1144) );
OR2_X1 U955 ( .A1(n984), .A2(n985), .ZN(n1211) );
NAND2_X1 U956 ( .A1(n985), .A2(n984), .ZN(n987) );
INV_X1 U957 ( .A(G475), .ZN(n984) );
NOR2_X1 U958 ( .A1(n1073), .A2(G902), .ZN(n985) );
XNOR2_X1 U959 ( .A(n1212), .B(n1194), .ZN(n1073) );
XOR2_X1 U960 ( .A(G104), .B(G113), .Z(n1194) );
XOR2_X1 U961 ( .A(n1213), .B(G122), .Z(n1212) );
NAND2_X1 U962 ( .A1(n1214), .A2(KEYINPUT28), .ZN(n1213) );
XOR2_X1 U963 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U964 ( .A(n1038), .B(n1217), .ZN(n1216) );
XOR2_X1 U965 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR2_X1 U966 ( .A1(G146), .A2(KEYINPUT8), .ZN(n1219) );
AND3_X1 U967 ( .A1(G214), .A2(n1030), .A3(n1179), .ZN(n1218) );
XOR2_X1 U968 ( .A(n1220), .B(n1221), .Z(n1215) );
XNOR2_X1 U969 ( .A(n1208), .B(G131), .ZN(n1221) );
XNOR2_X1 U970 ( .A(KEYINPUT33), .B(KEYINPUT1), .ZN(n1220) );
NOR2_X1 U971 ( .A1(n1141), .A2(n1154), .ZN(n1015) );
XOR2_X1 U972 ( .A(n1222), .B(n996), .Z(n1154) );
NAND2_X1 U973 ( .A1(n1066), .A2(n1117), .ZN(n996) );
XOR2_X1 U974 ( .A(n1223), .B(n1224), .Z(n1066) );
XOR2_X1 U975 ( .A(n1225), .B(n1226), .Z(n1224) );
NAND2_X1 U976 ( .A1(n1227), .A2(KEYINPUT27), .ZN(n1226) );
XOR2_X1 U977 ( .A(n1228), .B(n1229), .Z(n1227) );
NAND3_X1 U978 ( .A1(G234), .A2(n1030), .A3(G221), .ZN(n1228) );
NAND3_X1 U979 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1225) );
NAND2_X1 U980 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND3_X1 U981 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1233) );
NAND2_X1 U982 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U983 ( .A1(KEYINPUT40), .A2(n1240), .ZN(n1236) );
NAND2_X1 U984 ( .A1(n1037), .A2(n1241), .ZN(n1240) );
NAND2_X1 U985 ( .A1(KEYINPUT29), .A2(KEYINPUT19), .ZN(n1241) );
OR2_X1 U986 ( .A1(n1038), .A2(KEYINPUT40), .ZN(n1235) );
INV_X1 U987 ( .A(n1037), .ZN(n1038) );
NAND4_X1 U988 ( .A1(n1037), .A2(n1238), .A3(G146), .A4(KEYINPUT29), .ZN(n1231) );
INV_X1 U989 ( .A(KEYINPUT19), .ZN(n1238) );
NAND2_X1 U990 ( .A1(n1242), .A2(n1239), .ZN(n1230) );
INV_X1 U991 ( .A(KEYINPUT29), .ZN(n1239) );
NAND2_X1 U992 ( .A1(n1037), .A2(n1243), .ZN(n1242) );
NAND2_X1 U993 ( .A1(KEYINPUT19), .A2(G146), .ZN(n1243) );
XOR2_X1 U994 ( .A(G125), .B(G140), .Z(n1037) );
XNOR2_X1 U995 ( .A(G110), .B(n1244), .ZN(n1223) );
XNOR2_X1 U996 ( .A(n1153), .B(G119), .ZN(n1244) );
NAND2_X1 U997 ( .A1(KEYINPUT16), .A2(n997), .ZN(n1222) );
NAND2_X1 U998 ( .A1(G217), .A2(n1165), .ZN(n997) );
NAND2_X1 U999 ( .A1(G234), .A2(n1117), .ZN(n1165) );
XNOR2_X1 U1000 ( .A(n992), .B(KEYINPUT5), .ZN(n1141) );
XOR2_X1 U1001 ( .A(n1245), .B(G472), .Z(n992) );
NAND2_X1 U1002 ( .A1(n1246), .A2(n1117), .ZN(n1245) );
INV_X1 U1003 ( .A(G902), .ZN(n1117) );
XOR2_X1 U1004 ( .A(n1247), .B(n1248), .Z(n1246) );
XNOR2_X1 U1005 ( .A(KEYINPUT18), .B(n1089), .ZN(n1248) );
NAND3_X1 U1006 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1089) );
NAND2_X1 U1007 ( .A1(KEYINPUT36), .A2(n1252), .ZN(n1251) );
NAND3_X1 U1008 ( .A1(n1253), .A2(n1254), .A3(n1153), .ZN(n1250) );
INV_X1 U1009 ( .A(KEYINPUT36), .ZN(n1254) );
OR2_X1 U1010 ( .A1(n1153), .A2(n1253), .ZN(n1249) );
NOR2_X1 U1011 ( .A1(n1255), .A2(n1252), .ZN(n1253) );
XOR2_X1 U1012 ( .A(n1256), .B(n1208), .Z(n1252) );
INV_X1 U1013 ( .A(G143), .ZN(n1208) );
NAND2_X1 U1014 ( .A1(KEYINPUT63), .A2(n1234), .ZN(n1256) );
INV_X1 U1015 ( .A(G146), .ZN(n1234) );
INV_X1 U1016 ( .A(KEYINPUT4), .ZN(n1255) );
INV_X1 U1017 ( .A(G128), .ZN(n1153) );
XOR2_X1 U1018 ( .A(n1087), .B(n1257), .Z(n1247) );
NOR2_X1 U1019 ( .A1(KEYINPUT56), .A2(n1080), .ZN(n1257) );
XOR2_X1 U1020 ( .A(n1258), .B(G101), .Z(n1080) );
NAND3_X1 U1021 ( .A1(n1179), .A2(n1030), .A3(G210), .ZN(n1258) );
INV_X1 U1022 ( .A(G953), .ZN(n1030) );
INV_X1 U1023 ( .A(G237), .ZN(n1179) );
XOR2_X1 U1024 ( .A(n1259), .B(n1260), .Z(n1087) );
XOR2_X1 U1025 ( .A(G116), .B(n1261), .Z(n1260) );
XNOR2_X1 U1026 ( .A(KEYINPUT41), .B(n1195), .ZN(n1261) );
INV_X1 U1027 ( .A(G119), .ZN(n1195) );
XNOR2_X1 U1028 ( .A(n1039), .B(G113), .ZN(n1259) );
XNOR2_X1 U1029 ( .A(n1262), .B(n1203), .ZN(n1039) );
XOR2_X1 U1030 ( .A(G134), .B(KEYINPUT57), .Z(n1203) );
XNOR2_X1 U1031 ( .A(G131), .B(n1229), .ZN(n1262) );
XOR2_X1 U1032 ( .A(G137), .B(KEYINPUT58), .Z(n1229) );
endmodule


