//Key = 1111001111110111100011110110011101100100010010010011001111101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
n1431, n1432, n1433, n1434, n1435, n1436, n1437;

XOR2_X1 U766 ( .A(G107), .B(n1081), .Z(G9) );
NOR2_X1 U767 ( .A1(n1082), .A2(n1083), .ZN(G75) );
NOR4_X1 U768 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1083) );
NOR4_X1 U769 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1086) );
INV_X1 U770 ( .A(n1092), .ZN(n1089) );
NOR2_X1 U771 ( .A1(n1093), .A2(n1094), .ZN(n1088) );
NOR2_X1 U772 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U773 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NOR3_X1 U774 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1097) );
NOR2_X1 U775 ( .A1(n1102), .A2(n1103), .ZN(n1093) );
NOR2_X1 U776 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR2_X1 U777 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
XOR2_X1 U778 ( .A(n1108), .B(KEYINPUT0), .Z(n1106) );
NAND3_X1 U779 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1084) );
NAND4_X1 U780 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1111) );
NAND2_X1 U781 ( .A1(n1116), .A2(n1091), .ZN(n1115) );
NAND2_X1 U782 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
INV_X1 U783 ( .A(KEYINPUT7), .ZN(n1118) );
NAND4_X1 U784 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1114) );
INV_X1 U785 ( .A(n1091), .ZN(n1122) );
NAND2_X1 U786 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1125), .ZN(n1120) );
OR2_X1 U788 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U789 ( .A1(KEYINPUT7), .A2(n1117), .ZN(n1119) );
NOR3_X1 U790 ( .A1(n1128), .A2(G953), .A3(n1129), .ZN(n1082) );
INV_X1 U791 ( .A(n1109), .ZN(n1129) );
NAND4_X1 U792 ( .A1(n1130), .A2(n1113), .A3(n1131), .A4(n1132), .ZN(n1109) );
NOR3_X1 U793 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
XOR2_X1 U794 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U795 ( .A(n1138), .B(KEYINPUT1), .Z(n1136) );
NOR2_X1 U796 ( .A1(n1139), .A2(n1140), .ZN(n1134) );
NAND3_X1 U797 ( .A1(n1141), .A2(n1142), .A3(n1099), .ZN(n1133) );
NOR3_X1 U798 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1131) );
NOR2_X1 U799 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
INV_X1 U800 ( .A(KEYINPUT52), .ZN(n1147) );
XNOR2_X1 U801 ( .A(KEYINPUT22), .B(n1148), .ZN(n1146) );
NOR2_X1 U802 ( .A1(KEYINPUT52), .A2(n1149), .ZN(n1144) );
XOR2_X1 U803 ( .A(KEYINPUT22), .B(n1101), .Z(n1149) );
INV_X1 U804 ( .A(n1150), .ZN(n1101) );
XOR2_X1 U805 ( .A(n1151), .B(n1152), .Z(n1143) );
XOR2_X1 U806 ( .A(n1153), .B(G478), .Z(n1130) );
XOR2_X1 U807 ( .A(n1087), .B(KEYINPUT26), .Z(n1128) );
INV_X1 U808 ( .A(G952), .ZN(n1087) );
XOR2_X1 U809 ( .A(n1154), .B(n1155), .Z(G72) );
XOR2_X1 U810 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U811 ( .A1(n1158), .A2(n1110), .ZN(n1157) );
NOR2_X1 U812 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NAND2_X1 U813 ( .A1(n1161), .A2(n1162), .ZN(n1156) );
XOR2_X1 U814 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U815 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND3_X1 U816 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1166) );
NAND2_X1 U817 ( .A1(KEYINPUT61), .A2(n1170), .ZN(n1169) );
NAND3_X1 U818 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1168) );
INV_X1 U819 ( .A(KEYINPUT61), .ZN(n1172) );
OR2_X1 U820 ( .A1(n1173), .A2(n1171), .ZN(n1167) );
NOR2_X1 U821 ( .A1(KEYINPUT4), .A2(n1170), .ZN(n1171) );
XNOR2_X1 U822 ( .A(n1174), .B(n1175), .ZN(n1170) );
NAND2_X1 U823 ( .A1(KEYINPUT20), .A2(G131), .ZN(n1174) );
NOR2_X1 U824 ( .A1(KEYINPUT43), .A2(n1176), .ZN(n1163) );
XOR2_X1 U825 ( .A(n1177), .B(KEYINPUT62), .Z(n1161) );
NAND2_X1 U826 ( .A1(G953), .A2(n1160), .ZN(n1177) );
NAND2_X1 U827 ( .A1(n1110), .A2(n1178), .ZN(n1154) );
NAND2_X1 U828 ( .A1(n1179), .A2(n1180), .ZN(G69) );
NAND2_X1 U829 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U830 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
NAND3_X1 U831 ( .A1(KEYINPUT41), .A2(n1185), .A3(n1110), .ZN(n1184) );
NAND3_X1 U832 ( .A1(n1186), .A2(n1187), .A3(G953), .ZN(n1183) );
OR3_X1 U833 ( .A1(n1185), .A2(n1188), .A3(n1182), .ZN(n1179) );
NAND2_X1 U834 ( .A1(n1189), .A2(n1190), .ZN(n1182) );
NAND2_X1 U835 ( .A1(G953), .A2(n1191), .ZN(n1190) );
XOR2_X1 U836 ( .A(n1192), .B(n1193), .Z(n1189) );
NAND2_X1 U837 ( .A1(KEYINPUT50), .A2(n1194), .ZN(n1192) );
AND2_X1 U838 ( .A1(n1195), .A2(n1196), .ZN(n1188) );
NAND3_X1 U839 ( .A1(n1197), .A2(n1186), .A3(G953), .ZN(n1196) );
NAND2_X1 U840 ( .A1(KEYINPUT41), .A2(n1187), .ZN(n1197) );
INV_X1 U841 ( .A(KEYINPUT49), .ZN(n1187) );
NAND2_X1 U842 ( .A1(KEYINPUT41), .A2(n1198), .ZN(n1195) );
NAND2_X1 U843 ( .A1(G953), .A2(n1186), .ZN(n1198) );
NAND2_X1 U844 ( .A1(G898), .A2(G224), .ZN(n1186) );
NOR2_X1 U845 ( .A1(n1199), .A2(n1200), .ZN(G66) );
NOR3_X1 U846 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
AND3_X1 U847 ( .A1(n1204), .A2(n1137), .A3(n1205), .ZN(n1203) );
NOR2_X1 U848 ( .A1(n1206), .A2(n1204), .ZN(n1202) );
NOR2_X1 U849 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR3_X1 U850 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(G63) );
AND2_X1 U851 ( .A1(KEYINPUT8), .A2(n1199), .ZN(n1211) );
NOR3_X1 U852 ( .A1(KEYINPUT8), .A2(G953), .A3(G952), .ZN(n1210) );
NOR3_X1 U853 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1209) );
NOR3_X1 U854 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
NOR2_X1 U855 ( .A1(n1218), .A2(n1219), .ZN(n1213) );
NOR2_X1 U856 ( .A1(n1207), .A2(n1216), .ZN(n1218) );
INV_X1 U857 ( .A(G478), .ZN(n1216) );
INV_X1 U858 ( .A(n1153), .ZN(n1212) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1220), .ZN(G60) );
XOR2_X1 U860 ( .A(n1221), .B(n1222), .Z(n1220) );
NOR2_X1 U861 ( .A1(n1140), .A2(n1217), .ZN(n1221) );
XOR2_X1 U862 ( .A(G104), .B(n1223), .Z(G6) );
NOR2_X1 U863 ( .A1(n1199), .A2(n1224), .ZN(G57) );
XOR2_X1 U864 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U865 ( .A(n1227), .B(n1228), .Z(n1225) );
NOR2_X1 U866 ( .A1(n1151), .A2(n1217), .ZN(n1228) );
NAND3_X1 U867 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1227) );
NAND2_X1 U868 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND3_X1 U869 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1232) );
NAND2_X1 U870 ( .A1(KEYINPUT2), .A2(n1237), .ZN(n1236) );
OR2_X1 U871 ( .A1(n1238), .A2(KEYINPUT37), .ZN(n1235) );
NAND2_X1 U872 ( .A1(KEYINPUT37), .A2(n1239), .ZN(n1234) );
NAND2_X1 U873 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NAND2_X1 U874 ( .A1(KEYINPUT25), .A2(n1242), .ZN(n1241) );
NAND4_X1 U875 ( .A1(n1240), .A2(G101), .A3(KEYINPUT2), .A4(KEYINPUT25), .ZN(n1230) );
NAND2_X1 U876 ( .A1(n1243), .A2(n1237), .ZN(n1229) );
INV_X1 U877 ( .A(KEYINPUT25), .ZN(n1237) );
NAND2_X1 U878 ( .A1(n1240), .A2(n1244), .ZN(n1243) );
NAND2_X1 U879 ( .A1(G101), .A2(n1242), .ZN(n1244) );
INV_X1 U880 ( .A(KEYINPUT2), .ZN(n1242) );
INV_X1 U881 ( .A(n1238), .ZN(n1240) );
NOR2_X1 U882 ( .A1(n1199), .A2(n1245), .ZN(G54) );
NOR3_X1 U883 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1245) );
NOR2_X1 U884 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NOR2_X1 U885 ( .A1(KEYINPUT28), .A2(n1251), .ZN(n1249) );
XNOR2_X1 U886 ( .A(KEYINPUT47), .B(n1252), .ZN(n1251) );
NOR3_X1 U887 ( .A1(n1253), .A2(KEYINPUT28), .A3(n1252), .ZN(n1247) );
INV_X1 U888 ( .A(n1250), .ZN(n1253) );
XOR2_X1 U889 ( .A(n1254), .B(n1255), .Z(n1250) );
XNOR2_X1 U890 ( .A(n1256), .B(n1257), .ZN(n1254) );
NOR2_X1 U891 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U892 ( .A(n1260), .B(KEYINPUT21), .Z(n1259) );
NAND2_X1 U893 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NOR2_X1 U894 ( .A1(n1262), .A2(n1261), .ZN(n1258) );
XOR2_X1 U895 ( .A(n1173), .B(n1263), .Z(n1261) );
NOR2_X1 U896 ( .A1(KEYINPUT19), .A2(n1264), .ZN(n1263) );
AND2_X1 U897 ( .A1(n1252), .A2(KEYINPUT28), .ZN(n1246) );
NAND2_X1 U898 ( .A1(n1205), .A2(G469), .ZN(n1252) );
NOR2_X1 U899 ( .A1(n1199), .A2(n1265), .ZN(G51) );
XOR2_X1 U900 ( .A(n1266), .B(n1267), .Z(n1265) );
NOR2_X1 U901 ( .A1(KEYINPUT38), .A2(n1268), .ZN(n1267) );
XOR2_X1 U902 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U903 ( .A(n1271), .B(KEYINPUT40), .Z(n1270) );
NAND2_X1 U904 ( .A1(n1272), .A2(n1273), .ZN(n1269) );
NAND2_X1 U905 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U906 ( .A(n1176), .B(KEYINPUT30), .Z(n1274) );
NAND2_X1 U907 ( .A1(n1276), .A2(n1277), .ZN(n1272) );
XOR2_X1 U908 ( .A(n1176), .B(KEYINPUT24), .Z(n1277) );
INV_X1 U909 ( .A(n1275), .ZN(n1276) );
NAND2_X1 U910 ( .A1(n1205), .A2(n1278), .ZN(n1266) );
INV_X1 U911 ( .A(n1217), .ZN(n1205) );
NAND2_X1 U912 ( .A1(G902), .A2(n1085), .ZN(n1217) );
INV_X1 U913 ( .A(n1207), .ZN(n1085) );
NOR2_X1 U914 ( .A1(n1185), .A2(n1178), .ZN(n1207) );
NAND4_X1 U915 ( .A1(n1279), .A2(n1280), .A3(n1281), .A4(n1282), .ZN(n1178) );
NOR4_X1 U916 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1282) );
AND2_X1 U917 ( .A1(n1287), .A2(n1288), .ZN(n1281) );
NAND2_X1 U918 ( .A1(n1289), .A2(n1105), .ZN(n1279) );
INV_X1 U919 ( .A(n1290), .ZN(n1289) );
NAND4_X1 U920 ( .A1(n1291), .A2(n1292), .A3(n1293), .A4(n1294), .ZN(n1185) );
NOR4_X1 U921 ( .A1(n1295), .A2(n1081), .A3(n1223), .A4(n1296), .ZN(n1294) );
NOR3_X1 U922 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1296) );
AND3_X1 U923 ( .A1(n1300), .A2(n1092), .A3(n1126), .ZN(n1223) );
AND3_X1 U924 ( .A1(n1127), .A2(n1092), .A3(n1300), .ZN(n1081) );
INV_X1 U925 ( .A(n1301), .ZN(n1295) );
NOR2_X1 U926 ( .A1(n1302), .A2(n1303), .ZN(n1293) );
NOR2_X1 U927 ( .A1(n1110), .A2(G952), .ZN(n1199) );
XNOR2_X1 U928 ( .A(G146), .B(n1280), .ZN(G48) );
NAND3_X1 U929 ( .A1(n1126), .A2(n1098), .A3(n1304), .ZN(n1280) );
XOR2_X1 U930 ( .A(G143), .B(n1305), .Z(G45) );
NOR2_X1 U931 ( .A1(n1290), .A2(n1306), .ZN(n1305) );
XOR2_X1 U932 ( .A(KEYINPUT57), .B(n1105), .Z(n1306) );
NAND3_X1 U933 ( .A1(n1123), .A2(n1098), .A3(n1307), .ZN(n1290) );
AND3_X1 U934 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1307) );
XOR2_X1 U935 ( .A(n1287), .B(n1311), .Z(G42) );
XOR2_X1 U936 ( .A(n1165), .B(KEYINPUT39), .Z(n1311) );
NAND3_X1 U937 ( .A1(n1126), .A2(n1312), .A3(n1313), .ZN(n1287) );
XOR2_X1 U938 ( .A(G137), .B(n1286), .Z(G39) );
AND3_X1 U939 ( .A1(n1304), .A2(n1124), .A3(n1112), .ZN(n1286) );
XNOR2_X1 U940 ( .A(n1285), .B(n1314), .ZN(G36) );
XOR2_X1 U941 ( .A(KEYINPUT16), .B(G134), .Z(n1314) );
AND3_X1 U942 ( .A1(n1123), .A2(n1127), .A3(n1313), .ZN(n1285) );
XOR2_X1 U943 ( .A(G131), .B(n1284), .Z(G33) );
AND3_X1 U944 ( .A1(n1126), .A2(n1123), .A3(n1313), .ZN(n1284) );
AND3_X1 U945 ( .A1(n1105), .A2(n1310), .A3(n1112), .ZN(n1313) );
INV_X1 U946 ( .A(n1103), .ZN(n1112) );
NAND3_X1 U947 ( .A1(n1099), .A2(n1142), .A3(n1150), .ZN(n1103) );
XOR2_X1 U948 ( .A(G128), .B(n1283), .Z(G30) );
AND3_X1 U949 ( .A1(n1127), .A2(n1098), .A3(n1304), .ZN(n1283) );
AND4_X1 U950 ( .A1(n1105), .A2(n1315), .A3(n1310), .A4(n1316), .ZN(n1304) );
XOR2_X1 U951 ( .A(n1233), .B(n1301), .Z(G3) );
NAND3_X1 U952 ( .A1(n1124), .A2(n1300), .A3(n1123), .ZN(n1301) );
XOR2_X1 U953 ( .A(n1176), .B(n1288), .Z(G27) );
NAND4_X1 U954 ( .A1(n1098), .A2(n1310), .A3(n1113), .A4(n1317), .ZN(n1288) );
NOR2_X1 U955 ( .A1(n1318), .A2(n1297), .ZN(n1317) );
NAND2_X1 U956 ( .A1(n1091), .A2(n1319), .ZN(n1310) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1320), .A4(n1160), .ZN(n1319) );
INV_X1 U958 ( .A(G900), .ZN(n1160) );
XNOR2_X1 U959 ( .A(G122), .B(n1321), .ZN(G24) );
NOR2_X1 U960 ( .A1(n1322), .A2(KEYINPUT35), .ZN(n1321) );
INV_X1 U961 ( .A(n1291), .ZN(n1322) );
NAND4_X1 U962 ( .A1(n1323), .A2(n1092), .A3(n1308), .A4(n1309), .ZN(n1291) );
NOR2_X1 U963 ( .A1(n1316), .A2(n1324), .ZN(n1092) );
XNOR2_X1 U964 ( .A(G119), .B(n1292), .ZN(G21) );
NAND4_X1 U965 ( .A1(n1323), .A2(n1124), .A3(n1315), .A4(n1316), .ZN(n1292) );
XOR2_X1 U966 ( .A(n1325), .B(n1303), .Z(G18) );
AND3_X1 U967 ( .A1(n1123), .A2(n1127), .A3(n1323), .ZN(n1303) );
INV_X1 U968 ( .A(n1299), .ZN(n1323) );
NAND3_X1 U969 ( .A1(n1098), .A2(n1326), .A3(n1113), .ZN(n1299) );
NOR2_X1 U970 ( .A1(n1309), .A2(n1327), .ZN(n1127) );
XOR2_X1 U971 ( .A(n1328), .B(KEYINPUT34), .Z(n1325) );
XNOR2_X1 U972 ( .A(G113), .B(n1329), .ZN(G15) );
NAND4_X1 U973 ( .A1(n1330), .A2(n1126), .A3(n1331), .A4(n1123), .ZN(n1329) );
INV_X1 U974 ( .A(n1298), .ZN(n1123) );
NAND2_X1 U975 ( .A1(n1332), .A2(n1315), .ZN(n1298) );
XNOR2_X1 U976 ( .A(n1324), .B(KEYINPUT6), .ZN(n1315) );
AND2_X1 U977 ( .A1(n1326), .A2(n1113), .ZN(n1331) );
INV_X1 U978 ( .A(n1096), .ZN(n1113) );
NAND2_X1 U979 ( .A1(n1108), .A2(n1107), .ZN(n1096) );
INV_X1 U980 ( .A(n1297), .ZN(n1126) );
NAND2_X1 U981 ( .A1(n1327), .A2(n1309), .ZN(n1297) );
XNOR2_X1 U982 ( .A(n1098), .B(KEYINPUT23), .ZN(n1330) );
XOR2_X1 U983 ( .A(G110), .B(n1302), .Z(G12) );
AND2_X1 U984 ( .A1(n1117), .A2(n1300), .ZN(n1302) );
AND3_X1 U985 ( .A1(n1098), .A2(n1326), .A3(n1105), .ZN(n1300) );
AND2_X1 U986 ( .A1(n1333), .A2(n1107), .ZN(n1105) );
NAND2_X1 U987 ( .A1(G221), .A2(n1334), .ZN(n1107) );
INV_X1 U988 ( .A(n1108), .ZN(n1333) );
XOR2_X1 U989 ( .A(n1335), .B(G469), .Z(n1108) );
NAND3_X1 U990 ( .A1(n1336), .A2(n1337), .A3(n1338), .ZN(n1335) );
XOR2_X1 U991 ( .A(KEYINPUT14), .B(G902), .Z(n1338) );
NAND2_X1 U992 ( .A1(n1339), .A2(n1340), .ZN(n1337) );
NAND2_X1 U993 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U994 ( .A(n1343), .B(n1344), .Z(n1339) );
NAND2_X1 U995 ( .A1(KEYINPUT54), .A2(n1345), .ZN(n1343) );
NAND3_X1 U996 ( .A1(n1346), .A2(n1342), .A3(n1341), .ZN(n1336) );
INV_X1 U997 ( .A(n1262), .ZN(n1341) );
INV_X1 U998 ( .A(KEYINPUT45), .ZN(n1342) );
XOR2_X1 U999 ( .A(n1347), .B(n1344), .Z(n1346) );
XNOR2_X1 U1000 ( .A(n1255), .B(n1348), .ZN(n1344) );
XNOR2_X1 U1001 ( .A(n1349), .B(KEYINPUT42), .ZN(n1348) );
NAND2_X1 U1002 ( .A1(KEYINPUT55), .A2(n1256), .ZN(n1349) );
NOR2_X1 U1003 ( .A1(n1159), .A2(G953), .ZN(n1256) );
INV_X1 U1004 ( .A(G227), .ZN(n1159) );
XOR2_X1 U1005 ( .A(n1350), .B(n1165), .Z(n1255) );
INV_X1 U1006 ( .A(G110), .ZN(n1350) );
NAND2_X1 U1007 ( .A1(KEYINPUT54), .A2(n1351), .ZN(n1347) );
INV_X1 U1008 ( .A(n1345), .ZN(n1351) );
XNOR2_X1 U1009 ( .A(n1173), .B(n1264), .ZN(n1345) );
XNOR2_X1 U1010 ( .A(n1352), .B(n1353), .ZN(n1264) );
XOR2_X1 U1011 ( .A(KEYINPUT46), .B(G107), .Z(n1353) );
XOR2_X1 U1012 ( .A(G104), .B(n1233), .Z(n1352) );
XNOR2_X1 U1013 ( .A(n1354), .B(n1355), .ZN(n1173) );
INV_X1 U1014 ( .A(G128), .ZN(n1354) );
NAND2_X1 U1015 ( .A1(n1356), .A2(n1091), .ZN(n1326) );
NAND3_X1 U1016 ( .A1(n1320), .A2(n1110), .A3(G952), .ZN(n1091) );
NAND4_X1 U1017 ( .A1(G953), .A2(G902), .A3(n1320), .A4(n1191), .ZN(n1356) );
INV_X1 U1018 ( .A(G898), .ZN(n1191) );
NAND2_X1 U1019 ( .A1(G237), .A2(G234), .ZN(n1320) );
AND2_X1 U1020 ( .A1(n1357), .A2(n1099), .ZN(n1098) );
NAND2_X1 U1021 ( .A1(n1358), .A2(G214), .ZN(n1099) );
XOR2_X1 U1022 ( .A(n1359), .B(KEYINPUT48), .Z(n1358) );
NAND2_X1 U1023 ( .A1(n1150), .A2(n1142), .ZN(n1357) );
INV_X1 U1024 ( .A(n1100), .ZN(n1142) );
NOR2_X1 U1025 ( .A1(n1148), .A2(n1278), .ZN(n1100) );
NAND2_X1 U1026 ( .A1(n1278), .A2(n1148), .ZN(n1150) );
NAND2_X1 U1027 ( .A1(n1360), .A2(n1361), .ZN(n1148) );
XOR2_X1 U1028 ( .A(n1271), .B(n1362), .Z(n1360) );
XOR2_X1 U1029 ( .A(n1275), .B(G125), .Z(n1362) );
XOR2_X1 U1030 ( .A(n1363), .B(n1364), .Z(n1271) );
XOR2_X1 U1031 ( .A(KEYINPUT17), .B(n1365), .Z(n1364) );
AND2_X1 U1032 ( .A1(n1110), .A2(G224), .ZN(n1365) );
XOR2_X1 U1033 ( .A(n1366), .B(n1193), .Z(n1363) );
XNOR2_X1 U1034 ( .A(n1367), .B(n1368), .ZN(n1193) );
XOR2_X1 U1035 ( .A(n1369), .B(n1370), .Z(n1368) );
NAND2_X1 U1036 ( .A1(KEYINPUT51), .A2(n1371), .ZN(n1369) );
XOR2_X1 U1037 ( .A(n1372), .B(n1373), .Z(n1367) );
XNOR2_X1 U1038 ( .A(G104), .B(n1374), .ZN(n1373) );
NAND2_X1 U1039 ( .A1(n1375), .A2(KEYINPUT3), .ZN(n1374) );
XOR2_X1 U1040 ( .A(n1233), .B(KEYINPUT12), .Z(n1375) );
INV_X1 U1041 ( .A(G101), .ZN(n1233) );
NAND2_X1 U1042 ( .A1(KEYINPUT13), .A2(n1328), .ZN(n1372) );
INV_X1 U1043 ( .A(G116), .ZN(n1328) );
NAND2_X1 U1044 ( .A1(n1376), .A2(n1377), .ZN(n1366) );
NAND2_X1 U1045 ( .A1(KEYINPUT27), .A2(n1194), .ZN(n1377) );
OR2_X1 U1046 ( .A1(KEYINPUT53), .A2(n1194), .ZN(n1376) );
XOR2_X1 U1047 ( .A(G110), .B(n1378), .Z(n1194) );
AND2_X1 U1048 ( .A1(G210), .A2(n1359), .ZN(n1278) );
NAND2_X1 U1049 ( .A1(n1361), .A2(n1379), .ZN(n1359) );
INV_X1 U1050 ( .A(G237), .ZN(n1379) );
NOR2_X1 U1051 ( .A1(n1318), .A2(n1090), .ZN(n1117) );
INV_X1 U1052 ( .A(n1124), .ZN(n1090) );
NOR2_X1 U1053 ( .A1(n1308), .A2(n1309), .ZN(n1124) );
NAND2_X1 U1054 ( .A1(n1380), .A2(n1141), .ZN(n1309) );
NAND2_X1 U1055 ( .A1(n1139), .A2(n1140), .ZN(n1141) );
INV_X1 U1056 ( .A(G475), .ZN(n1140) );
NAND2_X1 U1057 ( .A1(G475), .A2(n1381), .ZN(n1380) );
XOR2_X1 U1058 ( .A(KEYINPUT9), .B(n1139), .Z(n1381) );
NOR2_X1 U1059 ( .A1(n1222), .A2(G902), .ZN(n1139) );
XNOR2_X1 U1060 ( .A(n1382), .B(n1383), .ZN(n1222) );
XOR2_X1 U1061 ( .A(G113), .B(G104), .Z(n1383) );
XOR2_X1 U1062 ( .A(n1384), .B(n1378), .Z(n1382) );
INV_X1 U1063 ( .A(n1385), .ZN(n1378) );
NAND2_X1 U1064 ( .A1(n1386), .A2(n1387), .ZN(n1384) );
NAND2_X1 U1065 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
XOR2_X1 U1066 ( .A(KEYINPUT29), .B(n1390), .Z(n1386) );
NOR2_X1 U1067 ( .A1(n1388), .A2(n1389), .ZN(n1390) );
XNOR2_X1 U1068 ( .A(n1391), .B(n1392), .ZN(n1389) );
XOR2_X1 U1069 ( .A(G143), .B(G131), .Z(n1392) );
NAND2_X1 U1070 ( .A1(n1393), .A2(G214), .ZN(n1391) );
XOR2_X1 U1071 ( .A(n1394), .B(n1395), .Z(n1388) );
XOR2_X1 U1072 ( .A(n1165), .B(G125), .Z(n1394) );
INV_X1 U1073 ( .A(G140), .ZN(n1165) );
INV_X1 U1074 ( .A(n1327), .ZN(n1308) );
XOR2_X1 U1075 ( .A(n1396), .B(n1397), .Z(n1327) );
XOR2_X1 U1076 ( .A(KEYINPUT33), .B(G478), .Z(n1397) );
NAND2_X1 U1077 ( .A1(KEYINPUT15), .A2(n1153), .ZN(n1396) );
NAND2_X1 U1078 ( .A1(n1215), .A2(n1361), .ZN(n1153) );
INV_X1 U1079 ( .A(n1219), .ZN(n1215) );
XOR2_X1 U1080 ( .A(n1398), .B(n1399), .Z(n1219) );
AND2_X1 U1081 ( .A1(n1400), .A2(G217), .ZN(n1399) );
NAND2_X1 U1082 ( .A1(KEYINPUT58), .A2(n1401), .ZN(n1398) );
XOR2_X1 U1083 ( .A(n1402), .B(n1403), .Z(n1401) );
XOR2_X1 U1084 ( .A(n1385), .B(n1404), .Z(n1403) );
NOR2_X1 U1085 ( .A1(KEYINPUT63), .A2(n1405), .ZN(n1404) );
XOR2_X1 U1086 ( .A(n1406), .B(n1407), .Z(n1405) );
XOR2_X1 U1087 ( .A(G128), .B(n1408), .Z(n1407) );
NOR2_X1 U1088 ( .A1(KEYINPUT36), .A2(n1409), .ZN(n1408) );
INV_X1 U1089 ( .A(G143), .ZN(n1409) );
XNOR2_X1 U1090 ( .A(G122), .B(KEYINPUT31), .ZN(n1385) );
XOR2_X1 U1091 ( .A(n1371), .B(G116), .Z(n1402) );
INV_X1 U1092 ( .A(G107), .ZN(n1371) );
INV_X1 U1093 ( .A(n1312), .ZN(n1318) );
NOR2_X1 U1094 ( .A1(n1324), .A2(n1332), .ZN(n1312) );
INV_X1 U1095 ( .A(n1316), .ZN(n1332) );
NAND2_X1 U1096 ( .A1(n1410), .A2(n1411), .ZN(n1316) );
NAND2_X1 U1097 ( .A1(n1412), .A2(n1208), .ZN(n1411) );
NAND2_X1 U1098 ( .A1(n1138), .A2(n1413), .ZN(n1412) );
NAND2_X1 U1099 ( .A1(KEYINPUT59), .A2(KEYINPUT56), .ZN(n1413) );
NAND3_X1 U1100 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(n1410) );
INV_X1 U1101 ( .A(KEYINPUT59), .ZN(n1416) );
OR2_X1 U1102 ( .A1(n1201), .A2(KEYINPUT56), .ZN(n1415) );
NAND2_X1 U1103 ( .A1(KEYINPUT56), .A2(n1417), .ZN(n1414) );
NAND2_X1 U1104 ( .A1(n1137), .A2(n1138), .ZN(n1417) );
INV_X1 U1105 ( .A(n1201), .ZN(n1138) );
NOR2_X1 U1106 ( .A1(n1204), .A2(G902), .ZN(n1201) );
XNOR2_X1 U1107 ( .A(n1418), .B(n1419), .ZN(n1204) );
XOR2_X1 U1108 ( .A(n1420), .B(n1421), .Z(n1419) );
XOR2_X1 U1109 ( .A(G128), .B(G119), .Z(n1421) );
XOR2_X1 U1110 ( .A(G140), .B(G137), .Z(n1420) );
XOR2_X1 U1111 ( .A(n1422), .B(n1423), .Z(n1418) );
XOR2_X1 U1112 ( .A(n1424), .B(n1395), .Z(n1423) );
XOR2_X1 U1113 ( .A(G146), .B(KEYINPUT60), .Z(n1395) );
NOR2_X1 U1114 ( .A1(KEYINPUT32), .A2(n1176), .ZN(n1424) );
INV_X1 U1115 ( .A(G125), .ZN(n1176) );
XOR2_X1 U1116 ( .A(n1425), .B(G110), .Z(n1422) );
NAND2_X1 U1117 ( .A1(n1400), .A2(G221), .ZN(n1425) );
AND2_X1 U1118 ( .A1(G234), .A2(n1110), .ZN(n1400) );
INV_X1 U1119 ( .A(G953), .ZN(n1110) );
INV_X1 U1120 ( .A(n1208), .ZN(n1137) );
NAND2_X1 U1121 ( .A1(G217), .A2(n1334), .ZN(n1208) );
NAND2_X1 U1122 ( .A1(G234), .A2(n1361), .ZN(n1334) );
XNOR2_X1 U1123 ( .A(n1426), .B(n1152), .ZN(n1324) );
NAND2_X1 U1124 ( .A1(n1427), .A2(n1361), .ZN(n1152) );
INV_X1 U1125 ( .A(G902), .ZN(n1361) );
XOR2_X1 U1126 ( .A(n1428), .B(n1429), .Z(n1427) );
XOR2_X1 U1127 ( .A(n1238), .B(G101), .Z(n1429) );
NAND2_X1 U1128 ( .A1(n1393), .A2(G210), .ZN(n1238) );
NOR2_X1 U1129 ( .A1(G953), .A2(G237), .ZN(n1393) );
NAND2_X1 U1130 ( .A1(KEYINPUT11), .A2(n1226), .ZN(n1428) );
XNOR2_X1 U1131 ( .A(n1430), .B(n1431), .ZN(n1226) );
XOR2_X1 U1132 ( .A(n1275), .B(n1370), .Z(n1431) );
XNOR2_X1 U1133 ( .A(G113), .B(G119), .ZN(n1370) );
NAND2_X1 U1134 ( .A1(n1432), .A2(n1433), .ZN(n1275) );
NAND2_X1 U1135 ( .A1(G128), .A2(n1355), .ZN(n1433) );
XOR2_X1 U1136 ( .A(KEYINPUT10), .B(n1434), .Z(n1432) );
NOR2_X1 U1137 ( .A1(G128), .A2(n1355), .ZN(n1434) );
XOR2_X1 U1138 ( .A(G146), .B(G143), .Z(n1355) );
XOR2_X1 U1139 ( .A(n1262), .B(G116), .Z(n1430) );
NAND2_X1 U1140 ( .A1(n1435), .A2(n1436), .ZN(n1262) );
NAND2_X1 U1141 ( .A1(G131), .A2(n1175), .ZN(n1436) );
XOR2_X1 U1142 ( .A(n1437), .B(KEYINPUT5), .Z(n1435) );
OR2_X1 U1143 ( .A1(n1175), .A2(G131), .ZN(n1437) );
XOR2_X1 U1144 ( .A(G137), .B(n1406), .Z(n1175) );
XOR2_X1 U1145 ( .A(G134), .B(KEYINPUT18), .Z(n1406) );
NAND2_X1 U1146 ( .A1(KEYINPUT44), .A2(n1151), .ZN(n1426) );
INV_X1 U1147 ( .A(G472), .ZN(n1151) );
endmodule


