//Key = 0011000101110110011110001010100110101101100001101101011010100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;

XNOR2_X1 U713 ( .A(G107), .B(n979), .ZN(G9) );
NOR2_X1 U714 ( .A1(n980), .A2(n981), .ZN(G75) );
NOR3_X1 U715 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n981) );
NOR4_X1 U716 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n983) );
NOR2_X1 U717 ( .A1(n989), .A2(n990), .ZN(n985) );
NOR2_X1 U718 ( .A1(n991), .A2(n992), .ZN(n990) );
NOR3_X1 U719 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n989) );
NOR3_X1 U720 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n995) );
NOR2_X1 U721 ( .A1(n999), .A2(n1000), .ZN(n994) );
NAND3_X1 U722 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n982) );
NAND4_X1 U723 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1003) );
NOR2_X1 U724 ( .A1(n996), .A2(n992), .ZN(n1007) );
INV_X1 U725 ( .A(n999), .ZN(n992) );
NAND3_X1 U726 ( .A1(n1008), .A2(n1009), .A3(n988), .ZN(n1005) );
NAND2_X1 U727 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
INV_X1 U728 ( .A(KEYINPUT2), .ZN(n1011) );
NAND2_X1 U729 ( .A1(KEYINPUT15), .A2(n1012), .ZN(n1008) );
NAND4_X1 U730 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1004) );
INV_X1 U731 ( .A(n988), .ZN(n1016) );
NOR2_X1 U732 ( .A1(n1017), .A2(n1018), .ZN(n1015) );
NOR2_X1 U733 ( .A1(n1019), .A2(n986), .ZN(n1018) );
AND2_X1 U734 ( .A1(n1020), .A2(n1021), .ZN(n1017) );
NAND2_X1 U735 ( .A1(KEYINPUT2), .A2(n1010), .ZN(n1014) );
NAND2_X1 U736 ( .A1(n1012), .A2(n1022), .ZN(n1013) );
INV_X1 U737 ( .A(KEYINPUT15), .ZN(n1022) );
NOR3_X1 U738 ( .A1(n986), .A2(n1023), .A3(n1024), .ZN(n1012) );
INV_X1 U739 ( .A(n1025), .ZN(n986) );
NOR3_X1 U740 ( .A1(n1026), .A2(G953), .A3(G952), .ZN(n980) );
INV_X1 U741 ( .A(n1001), .ZN(n1026) );
NAND4_X1 U742 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1001) );
NOR4_X1 U743 ( .A1(n996), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1030) );
XOR2_X1 U744 ( .A(n1034), .B(KEYINPUT40), .Z(n1033) );
XOR2_X1 U745 ( .A(n1035), .B(n1036), .Z(n1032) );
NOR2_X1 U746 ( .A1(KEYINPUT5), .A2(n1037), .ZN(n1036) );
XOR2_X1 U747 ( .A(n1038), .B(KEYINPUT39), .Z(n1035) );
INV_X1 U748 ( .A(n1000), .ZN(n996) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1029) );
XNOR2_X1 U750 ( .A(G469), .B(n1041), .ZN(n1040) );
XOR2_X1 U751 ( .A(n1042), .B(n1043), .Z(n1028) );
XOR2_X1 U752 ( .A(n1044), .B(KEYINPUT1), .Z(n1027) );
XOR2_X1 U753 ( .A(n1045), .B(n1046), .Z(G72) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U755 ( .A1(G953), .A2(n1049), .ZN(n1048) );
XOR2_X1 U756 ( .A(n1050), .B(KEYINPUT53), .Z(n1049) );
NAND2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1002), .ZN(n1047) );
NOR2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XNOR2_X1 U760 ( .A(G227), .B(KEYINPUT8), .ZN(n1054) );
NAND2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(n1045) );
XOR2_X1 U762 ( .A(n1058), .B(n1059), .Z(n1056) );
XOR2_X1 U763 ( .A(n1060), .B(G125), .Z(n1059) );
INV_X1 U764 ( .A(G140), .ZN(n1060) );
NAND3_X1 U765 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1058) );
OR2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND3_X1 U767 ( .A1(n1065), .A2(n1064), .A3(KEYINPUT49), .ZN(n1062) );
NOR2_X1 U768 ( .A1(KEYINPUT21), .A2(n1066), .ZN(n1065) );
NAND2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(n1061) );
INV_X1 U770 ( .A(KEYINPUT49), .ZN(n1067) );
XOR2_X1 U771 ( .A(n1068), .B(n1069), .Z(n1066) );
XOR2_X1 U772 ( .A(n1070), .B(n1071), .Z(G69) );
NOR2_X1 U773 ( .A1(n1072), .A2(n1002), .ZN(n1071) );
NOR2_X1 U774 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U775 ( .A1(n1075), .A2(n1076), .ZN(n1070) );
NAND2_X1 U776 ( .A1(n1077), .A2(n1002), .ZN(n1076) );
XNOR2_X1 U777 ( .A(n1078), .B(n1079), .ZN(n1077) );
NAND3_X1 U778 ( .A1(G898), .A2(n1079), .A3(G953), .ZN(n1075) );
XOR2_X1 U779 ( .A(n1080), .B(KEYINPUT6), .Z(n1079) );
NOR2_X1 U780 ( .A1(n1081), .A2(n1082), .ZN(G66) );
XOR2_X1 U781 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND2_X1 U782 ( .A1(KEYINPUT56), .A2(n1085), .ZN(n1084) );
NAND2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U784 ( .A(G217), .B(n1088), .ZN(n1087) );
XNOR2_X1 U785 ( .A(KEYINPUT36), .B(KEYINPUT31), .ZN(n1088) );
NOR2_X1 U786 ( .A1(G952), .A2(n1089), .ZN(n1081) );
XOR2_X1 U787 ( .A(KEYINPUT51), .B(G953), .Z(n1089) );
NOR2_X1 U788 ( .A1(n1090), .A2(n1091), .ZN(G63) );
XOR2_X1 U789 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR2_X1 U790 ( .A1(n1094), .A2(KEYINPUT35), .ZN(n1093) );
AND2_X1 U791 ( .A1(G478), .A2(n1086), .ZN(n1094) );
NOR2_X1 U792 ( .A1(n1090), .A2(n1095), .ZN(G60) );
XNOR2_X1 U793 ( .A(n1096), .B(n1097), .ZN(n1095) );
NOR2_X1 U794 ( .A1(n1038), .A2(n1098), .ZN(n1096) );
INV_X1 U795 ( .A(G475), .ZN(n1038) );
XOR2_X1 U796 ( .A(n1099), .B(n1100), .Z(G6) );
NOR2_X1 U797 ( .A1(G104), .A2(KEYINPUT60), .ZN(n1100) );
NAND2_X1 U798 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U799 ( .A1(n1090), .A2(n1103), .ZN(G57) );
XOR2_X1 U800 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U801 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U802 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U803 ( .A(n1110), .B(KEYINPUT50), .Z(n1109) );
INV_X1 U804 ( .A(n1111), .ZN(n1108) );
NOR2_X1 U805 ( .A1(n1111), .A2(n1112), .ZN(n1106) );
XOR2_X1 U806 ( .A(n1110), .B(KEYINPUT18), .Z(n1112) );
XNOR2_X1 U807 ( .A(n1113), .B(n1114), .ZN(n1111) );
XOR2_X1 U808 ( .A(n1115), .B(n1116), .Z(n1104) );
NOR2_X1 U809 ( .A1(KEYINPUT62), .A2(n1117), .ZN(n1116) );
NAND3_X1 U810 ( .A1(n1118), .A2(n1119), .A3(G472), .ZN(n1115) );
OR2_X1 U811 ( .A1(n1086), .A2(KEYINPUT55), .ZN(n1119) );
NAND2_X1 U812 ( .A1(KEYINPUT55), .A2(n1120), .ZN(n1118) );
OR2_X1 U813 ( .A1(n984), .A2(n1121), .ZN(n1120) );
NOR2_X1 U814 ( .A1(n1090), .A2(n1122), .ZN(G54) );
XOR2_X1 U815 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U816 ( .A1(n1086), .A2(G469), .ZN(n1123) );
NOR2_X1 U817 ( .A1(n1090), .A2(n1125), .ZN(G51) );
XOR2_X1 U818 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U819 ( .A1(KEYINPUT0), .A2(n1128), .ZN(n1127) );
XOR2_X1 U820 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U821 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U822 ( .A1(G125), .A2(KEYINPUT43), .ZN(n1132) );
XOR2_X1 U823 ( .A(n1080), .B(n1114), .Z(n1129) );
NAND2_X1 U824 ( .A1(n1086), .A2(n1043), .ZN(n1126) );
INV_X1 U825 ( .A(n1133), .ZN(n1043) );
INV_X1 U826 ( .A(n1098), .ZN(n1086) );
NAND2_X1 U827 ( .A1(G902), .A2(n984), .ZN(n1098) );
NAND3_X1 U828 ( .A1(n1051), .A2(n1134), .A3(n1078), .ZN(n984) );
AND4_X1 U829 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1078) );
AND4_X1 U830 ( .A1(n1139), .A2(n1140), .A3(n979), .A4(n1141), .ZN(n1138) );
INV_X1 U831 ( .A(n1142), .ZN(n1141) );
NAND4_X1 U832 ( .A1(n999), .A2(n1143), .A3(n1020), .A4(n1144), .ZN(n979) );
NAND2_X1 U833 ( .A1(n1102), .A2(n1145), .ZN(n1137) );
NAND2_X1 U834 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
OR2_X1 U835 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U836 ( .A(KEYINPUT32), .B(n1101), .Z(n1146) );
AND4_X1 U837 ( .A1(n1150), .A2(n999), .A3(n1151), .A4(n1144), .ZN(n1101) );
XOR2_X1 U838 ( .A(KEYINPUT11), .B(n1152), .Z(n1134) );
NOR4_X1 U839 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1051) );
OR4_X1 U840 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
NOR3_X1 U841 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
XOR2_X1 U842 ( .A(KEYINPUT26), .B(n1150), .Z(n1161) );
AND3_X1 U843 ( .A1(n1164), .A2(n1165), .A3(KEYINPUT29), .ZN(n1158) );
NOR2_X1 U844 ( .A1(n1164), .A2(n1166), .ZN(n1157) );
NOR2_X1 U845 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U846 ( .A1(KEYINPUT29), .A2(n1169), .ZN(n1168) );
INV_X1 U847 ( .A(n1170), .ZN(n1164) );
NOR2_X1 U848 ( .A1(n1002), .A2(G952), .ZN(n1090) );
XOR2_X1 U849 ( .A(n1068), .B(n1171), .Z(G48) );
NAND2_X1 U850 ( .A1(KEYINPUT34), .A2(n1152), .ZN(n1171) );
INV_X1 U851 ( .A(n1052), .ZN(n1152) );
NAND2_X1 U852 ( .A1(n1172), .A2(n1150), .ZN(n1052) );
XOR2_X1 U853 ( .A(n1173), .B(n1174), .Z(G45) );
NAND3_X1 U854 ( .A1(n1167), .A2(n1170), .A3(KEYINPUT14), .ZN(n1174) );
AND4_X1 U855 ( .A1(n998), .A2(n1143), .A3(n1175), .A4(n1176), .ZN(n1167) );
XOR2_X1 U856 ( .A(G140), .B(n1177), .Z(G42) );
NOR3_X1 U857 ( .A1(n1163), .A2(n1178), .A3(n1179), .ZN(n1177) );
XOR2_X1 U858 ( .A(n1162), .B(KEYINPUT41), .Z(n1178) );
XOR2_X1 U859 ( .A(G137), .B(n1159), .Z(G39) );
AND4_X1 U860 ( .A1(n1180), .A2(n1025), .A3(n1181), .A4(n1039), .ZN(n1159) );
XOR2_X1 U861 ( .A(G134), .B(n1155), .Z(G36) );
AND3_X1 U862 ( .A1(n998), .A2(n1020), .A3(n1180), .ZN(n1155) );
INV_X1 U863 ( .A(n1163), .ZN(n1180) );
XNOR2_X1 U864 ( .A(G131), .B(n1182), .ZN(G33) );
NAND2_X1 U865 ( .A1(KEYINPUT10), .A2(n1153), .ZN(n1182) );
NOR3_X1 U866 ( .A1(n1149), .A2(n1179), .A3(n1163), .ZN(n1153) );
NAND4_X1 U867 ( .A1(n1006), .A2(n1151), .A3(n1170), .A4(n1000), .ZN(n1163) );
XOR2_X1 U868 ( .A(G128), .B(n1154), .Z(G30) );
AND2_X1 U869 ( .A1(n1172), .A2(n1020), .ZN(n1154) );
AND4_X1 U870 ( .A1(n1143), .A2(n1181), .A3(n1039), .A4(n1170), .ZN(n1172) );
NOR2_X1 U871 ( .A1(n991), .A2(n1019), .ZN(n1143) );
XOR2_X1 U872 ( .A(G101), .B(n1183), .Z(G3) );
NOR3_X1 U873 ( .A1(n1184), .A2(n1149), .A3(n1148), .ZN(n1183) );
XOR2_X1 U874 ( .A(KEYINPUT17), .B(n1102), .Z(n1184) );
XOR2_X1 U875 ( .A(n1185), .B(G125), .Z(G27) );
NAND2_X1 U876 ( .A1(KEYINPUT13), .A2(n1186), .ZN(n1185) );
NAND2_X1 U877 ( .A1(n1165), .A2(n1170), .ZN(n1186) );
NAND2_X1 U878 ( .A1(n988), .A2(n1187), .ZN(n1170) );
NAND3_X1 U879 ( .A1(G902), .A2(n1188), .A3(n1189), .ZN(n1187) );
INV_X1 U880 ( .A(n1057), .ZN(n1189) );
NAND2_X1 U881 ( .A1(G953), .A2(n1055), .ZN(n1057) );
INV_X1 U882 ( .A(G900), .ZN(n1055) );
INV_X1 U883 ( .A(n1169), .ZN(n1165) );
NAND3_X1 U884 ( .A1(n997), .A2(n1102), .A3(n1010), .ZN(n1169) );
NOR2_X1 U885 ( .A1(n1179), .A2(n987), .ZN(n1010) );
INV_X1 U886 ( .A(n1021), .ZN(n987) );
XOR2_X1 U887 ( .A(n1190), .B(n1135), .Z(G24) );
NAND4_X1 U888 ( .A1(n1191), .A2(n999), .A3(n1175), .A4(n1176), .ZN(n1135) );
NOR2_X1 U889 ( .A1(n1039), .A2(n1181), .ZN(n999) );
XNOR2_X1 U890 ( .A(G119), .B(n1136), .ZN(G21) );
NAND4_X1 U891 ( .A1(n1191), .A2(n1025), .A3(n1181), .A4(n1039), .ZN(n1136) );
INV_X1 U892 ( .A(n1044), .ZN(n1181) );
XNOR2_X1 U893 ( .A(G116), .B(n1140), .ZN(G18) );
NAND3_X1 U894 ( .A1(n1191), .A2(n1020), .A3(n998), .ZN(n1140) );
NAND2_X1 U895 ( .A1(n1192), .A2(n1193), .ZN(n1020) );
OR3_X1 U896 ( .A1(n1034), .A2(n1176), .A3(KEYINPUT4), .ZN(n1193) );
NAND2_X1 U897 ( .A1(KEYINPUT4), .A2(n1025), .ZN(n1192) );
XNOR2_X1 U898 ( .A(G113), .B(n1139), .ZN(G15) );
NAND3_X1 U899 ( .A1(n1150), .A2(n1191), .A3(n998), .ZN(n1139) );
INV_X1 U900 ( .A(n1149), .ZN(n998) );
NAND2_X1 U901 ( .A1(n1044), .A2(n1039), .ZN(n1149) );
AND3_X1 U902 ( .A1(n1102), .A2(n1144), .A3(n1021), .ZN(n1191) );
NOR2_X1 U903 ( .A1(n1024), .A2(n1031), .ZN(n1021) );
INV_X1 U904 ( .A(n991), .ZN(n1102) );
INV_X1 U905 ( .A(n1179), .ZN(n1150) );
NAND2_X1 U906 ( .A1(n1034), .A2(n1176), .ZN(n1179) );
XOR2_X1 U907 ( .A(G110), .B(n1142), .Z(G12) );
NOR3_X1 U908 ( .A1(n1148), .A2(n991), .A3(n1162), .ZN(n1142) );
INV_X1 U909 ( .A(n997), .ZN(n1162) );
NOR2_X1 U910 ( .A1(n1039), .A2(n1044), .ZN(n997) );
XOR2_X1 U911 ( .A(n1194), .B(n1195), .Z(n1044) );
NOR2_X1 U912 ( .A1(G902), .A2(n1083), .ZN(n1195) );
NAND2_X1 U913 ( .A1(n1196), .A2(n1197), .ZN(n1083) );
NAND2_X1 U914 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NAND2_X1 U915 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U916 ( .A1(KEYINPUT37), .A2(n1202), .ZN(n1201) );
INV_X1 U917 ( .A(KEYINPUT27), .ZN(n1200) );
NAND2_X1 U918 ( .A1(n1203), .A2(n1204), .ZN(n1196) );
NAND2_X1 U919 ( .A1(KEYINPUT37), .A2(n1205), .ZN(n1204) );
OR2_X1 U920 ( .A1(n1198), .A2(KEYINPUT27), .ZN(n1205) );
XOR2_X1 U921 ( .A(n1206), .B(G137), .Z(n1198) );
NAND2_X1 U922 ( .A1(G221), .A2(n1207), .ZN(n1206) );
INV_X1 U923 ( .A(n1202), .ZN(n1203) );
XNOR2_X1 U924 ( .A(n1208), .B(n1209), .ZN(n1202) );
XOR2_X1 U925 ( .A(G110), .B(n1210), .Z(n1209) );
NOR2_X1 U926 ( .A1(KEYINPUT16), .A2(n1211), .ZN(n1210) );
XNOR2_X1 U927 ( .A(G128), .B(n1212), .ZN(n1211) );
NAND2_X1 U928 ( .A1(G217), .A2(n1213), .ZN(n1194) );
XNOR2_X1 U929 ( .A(n1214), .B(G472), .ZN(n1039) );
NAND2_X1 U930 ( .A1(n1215), .A2(n1121), .ZN(n1214) );
XOR2_X1 U931 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U932 ( .A(n1110), .B(n1117), .Z(n1217) );
AND2_X1 U933 ( .A1(n1218), .A2(n1219), .ZN(n1117) );
NAND2_X1 U934 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
INV_X1 U935 ( .A(G101), .ZN(n1221) );
NAND2_X1 U936 ( .A1(G210), .A2(n1222), .ZN(n1220) );
NAND3_X1 U937 ( .A1(G210), .A2(n1222), .A3(G101), .ZN(n1218) );
XOR2_X1 U938 ( .A(n1223), .B(n1224), .Z(n1110) );
NOR2_X1 U939 ( .A1(KEYINPUT52), .A2(n1212), .ZN(n1224) );
XOR2_X1 U940 ( .A(n1225), .B(KEYINPUT20), .Z(n1216) );
NAND3_X1 U941 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1225) );
NAND2_X1 U942 ( .A1(n1114), .A2(n1229), .ZN(n1228) );
NAND2_X1 U943 ( .A1(KEYINPUT59), .A2(n1230), .ZN(n1227) );
NAND2_X1 U944 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U945 ( .A(KEYINPUT28), .B(n1229), .Z(n1232) );
INV_X1 U946 ( .A(n1113), .ZN(n1229) );
NAND2_X1 U947 ( .A1(n1233), .A2(n1234), .ZN(n1226) );
INV_X1 U948 ( .A(KEYINPUT59), .ZN(n1234) );
NAND2_X1 U949 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
NAND3_X1 U950 ( .A1(KEYINPUT28), .A2(n1231), .A3(n1113), .ZN(n1236) );
OR2_X1 U951 ( .A1(n1113), .A2(KEYINPUT28), .ZN(n1235) );
NAND2_X1 U952 ( .A1(n993), .A2(n1000), .ZN(n991) );
NAND2_X1 U953 ( .A1(G214), .A2(n1237), .ZN(n1000) );
INV_X1 U954 ( .A(n1006), .ZN(n993) );
XOR2_X1 U955 ( .A(n1133), .B(n1238), .Z(n1006) );
NOR2_X1 U956 ( .A1(KEYINPUT57), .A2(n1042), .ZN(n1238) );
NAND2_X1 U957 ( .A1(n1239), .A2(n1121), .ZN(n1042) );
XOR2_X1 U958 ( .A(n1240), .B(n1241), .Z(n1239) );
INV_X1 U959 ( .A(n1080), .ZN(n1241) );
XOR2_X1 U960 ( .A(n1242), .B(n1243), .Z(n1080) );
XOR2_X1 U961 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U962 ( .A(G104), .B(n1246), .Z(n1245) );
XOR2_X1 U963 ( .A(KEYINPUT47), .B(KEYINPUT24), .Z(n1244) );
XOR2_X1 U964 ( .A(n1223), .B(n1247), .Z(n1242) );
XNOR2_X1 U965 ( .A(n1248), .B(n1212), .ZN(n1247) );
XNOR2_X1 U966 ( .A(G119), .B(KEYINPUT7), .ZN(n1212) );
XNOR2_X1 U967 ( .A(G116), .B(G113), .ZN(n1223) );
NAND3_X1 U968 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1240) );
NAND2_X1 U969 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
NAND2_X1 U970 ( .A1(KEYINPUT58), .A2(n1254), .ZN(n1253) );
XOR2_X1 U971 ( .A(KEYINPUT22), .B(n1131), .Z(n1254) );
INV_X1 U972 ( .A(n1255), .ZN(n1252) );
NAND3_X1 U973 ( .A1(KEYINPUT58), .A2(n1255), .A3(n1131), .ZN(n1250) );
XOR2_X1 U974 ( .A(G125), .B(n1114), .Z(n1255) );
INV_X1 U975 ( .A(n1231), .ZN(n1114) );
XOR2_X1 U976 ( .A(n1256), .B(n1257), .Z(n1231) );
XOR2_X1 U977 ( .A(n1173), .B(n1258), .Z(n1257) );
NAND2_X1 U978 ( .A1(KEYINPUT61), .A2(G128), .ZN(n1258) );
INV_X1 U979 ( .A(G143), .ZN(n1173) );
NAND2_X1 U980 ( .A1(KEYINPUT48), .A2(n1068), .ZN(n1256) );
INV_X1 U981 ( .A(G146), .ZN(n1068) );
OR2_X1 U982 ( .A1(n1131), .A2(KEYINPUT58), .ZN(n1249) );
NOR2_X1 U983 ( .A1(n1073), .A2(G953), .ZN(n1131) );
INV_X1 U984 ( .A(G224), .ZN(n1073) );
NAND2_X1 U985 ( .A1(G210), .A2(n1237), .ZN(n1133) );
NAND2_X1 U986 ( .A1(n1259), .A2(n1121), .ZN(n1237) );
INV_X1 U987 ( .A(G237), .ZN(n1259) );
NAND3_X1 U988 ( .A1(n1151), .A2(n1144), .A3(n1025), .ZN(n1148) );
NOR2_X1 U989 ( .A1(n1176), .A2(n1175), .ZN(n1025) );
INV_X1 U990 ( .A(n1034), .ZN(n1175) );
XOR2_X1 U991 ( .A(n1260), .B(G478), .Z(n1034) );
NAND2_X1 U992 ( .A1(n1092), .A2(n1121), .ZN(n1260) );
XOR2_X1 U993 ( .A(n1261), .B(n1262), .Z(n1092) );
XOR2_X1 U994 ( .A(n1069), .B(n1246), .Z(n1262) );
XOR2_X1 U995 ( .A(G107), .B(G122), .Z(n1246) );
XOR2_X1 U996 ( .A(n1263), .B(n1264), .Z(n1261) );
XNOR2_X1 U997 ( .A(G116), .B(n1265), .ZN(n1263) );
NOR2_X1 U998 ( .A1(n1266), .A2(KEYINPUT33), .ZN(n1265) );
AND2_X1 U999 ( .A1(n1207), .A2(G217), .ZN(n1266) );
AND2_X1 U1000 ( .A1(G234), .A2(n1002), .ZN(n1207) );
XNOR2_X1 U1001 ( .A(n1037), .B(G475), .ZN(n1176) );
NAND2_X1 U1002 ( .A1(n1267), .A2(n1097), .ZN(n1037) );
XOR2_X1 U1003 ( .A(n1268), .B(n1269), .Z(n1097) );
XOR2_X1 U1004 ( .A(n1270), .B(n1208), .Z(n1269) );
XOR2_X1 U1005 ( .A(G125), .B(n1271), .Z(n1208) );
NOR2_X1 U1006 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
XOR2_X1 U1007 ( .A(n1274), .B(KEYINPUT46), .Z(n1273) );
NAND2_X1 U1008 ( .A1(G113), .A2(n1190), .ZN(n1274) );
NOR2_X1 U1009 ( .A1(G113), .A2(n1190), .ZN(n1272) );
INV_X1 U1010 ( .A(G122), .ZN(n1190) );
XOR2_X1 U1011 ( .A(n1275), .B(n1276), .Z(n1268) );
NOR2_X1 U1012 ( .A1(KEYINPUT42), .A2(G104), .ZN(n1276) );
NAND2_X1 U1013 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
NAND2_X1 U1014 ( .A1(n1279), .A2(G131), .ZN(n1278) );
XOR2_X1 U1015 ( .A(KEYINPUT54), .B(n1280), .Z(n1277) );
NOR2_X1 U1016 ( .A1(G131), .A2(n1279), .ZN(n1280) );
XOR2_X1 U1017 ( .A(n1281), .B(n1282), .Z(n1279) );
XOR2_X1 U1018 ( .A(KEYINPUT38), .B(G143), .Z(n1282) );
NAND2_X1 U1019 ( .A1(G214), .A2(n1222), .ZN(n1281) );
NOR2_X1 U1020 ( .A1(G953), .A2(G237), .ZN(n1222) );
XOR2_X1 U1021 ( .A(n1121), .B(KEYINPUT30), .Z(n1267) );
NAND2_X1 U1022 ( .A1(n988), .A2(n1283), .ZN(n1144) );
NAND4_X1 U1023 ( .A1(G953), .A2(G902), .A3(n1188), .A4(n1074), .ZN(n1283) );
INV_X1 U1024 ( .A(G898), .ZN(n1074) );
NAND3_X1 U1025 ( .A1(n1188), .A2(n1002), .A3(G952), .ZN(n988) );
NAND2_X1 U1026 ( .A1(G237), .A2(G234), .ZN(n1188) );
INV_X1 U1027 ( .A(n1019), .ZN(n1151) );
NAND2_X1 U1028 ( .A1(n1284), .A2(n1024), .ZN(n1019) );
XOR2_X1 U1029 ( .A(G469), .B(n1285), .Z(n1024) );
NOR2_X1 U1030 ( .A1(KEYINPUT12), .A2(n1041), .ZN(n1285) );
NAND2_X1 U1031 ( .A1(n1286), .A2(n1121), .ZN(n1041) );
XNOR2_X1 U1032 ( .A(n1124), .B(KEYINPUT19), .ZN(n1286) );
XNOR2_X1 U1033 ( .A(n1287), .B(n1288), .ZN(n1124) );
XOR2_X1 U1034 ( .A(n1113), .B(n1289), .Z(n1288) );
XNOR2_X1 U1035 ( .A(n1248), .B(n1271), .ZN(n1289) );
XOR2_X1 U1036 ( .A(G140), .B(G146), .Z(n1271) );
XNOR2_X1 U1037 ( .A(n1290), .B(G101), .ZN(n1248) );
INV_X1 U1038 ( .A(G110), .ZN(n1290) );
XNOR2_X1 U1039 ( .A(n1291), .B(n1064), .ZN(n1113) );
XOR2_X1 U1040 ( .A(n1292), .B(n1264), .Z(n1064) );
XOR2_X1 U1041 ( .A(G134), .B(KEYINPUT44), .Z(n1264) );
XNOR2_X1 U1042 ( .A(G137), .B(G131), .ZN(n1292) );
XNOR2_X1 U1043 ( .A(KEYINPUT45), .B(KEYINPUT25), .ZN(n1291) );
XOR2_X1 U1044 ( .A(n1293), .B(n1294), .Z(n1287) );
XOR2_X1 U1045 ( .A(n1295), .B(n1069), .Z(n1294) );
XOR2_X1 U1046 ( .A(G128), .B(G143), .Z(n1069) );
AND2_X1 U1047 ( .A1(n1002), .A2(G227), .ZN(n1295) );
INV_X1 U1048 ( .A(G953), .ZN(n1002) );
XOR2_X1 U1049 ( .A(n1296), .B(KEYINPUT63), .Z(n1293) );
NAND2_X1 U1050 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
OR2_X1 U1051 ( .A1(n1299), .A2(G107), .ZN(n1298) );
XOR2_X1 U1052 ( .A(n1300), .B(KEYINPUT23), .Z(n1297) );
NAND2_X1 U1053 ( .A1(G107), .A2(n1299), .ZN(n1300) );
XOR2_X1 U1054 ( .A(G104), .B(KEYINPUT3), .Z(n1299) );
XOR2_X1 U1055 ( .A(KEYINPUT9), .B(n1031), .Z(n1284) );
INV_X1 U1056 ( .A(n1023), .ZN(n1031) );
NAND2_X1 U1057 ( .A1(G221), .A2(n1213), .ZN(n1023) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1121), .ZN(n1213) );
INV_X1 U1059 ( .A(G902), .ZN(n1121) );
endmodule


