//Key = 1100100100010110101011010111001101010110011001100101011010111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374;

XNOR2_X1 U750 ( .A(G107), .B(n1042), .ZN(G9) );
NAND3_X1 U751 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(G75) );
NAND2_X1 U752 ( .A1(G952), .A2(n1046), .ZN(n1045) );
NAND3_X1 U753 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND3_X1 U756 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND2_X1 U757 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
OR2_X1 U759 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1057) );
NAND2_X1 U761 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
OR3_X1 U762 ( .A1(n1067), .A2(KEYINPUT61), .A3(n1068), .ZN(n1066) );
NAND2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
INV_X1 U764 ( .A(KEYINPUT63), .ZN(n1070) );
NAND3_X1 U765 ( .A1(n1063), .A2(n1071), .A3(n1059), .ZN(n1052) );
NAND2_X1 U766 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U767 ( .A1(n1056), .A2(n1074), .ZN(n1073) );
OR2_X1 U768 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U769 ( .A1(n1054), .A2(n1077), .ZN(n1072) );
NAND3_X1 U770 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
NAND2_X1 U771 ( .A1(KEYINPUT61), .A2(n1056), .ZN(n1080) );
INV_X1 U772 ( .A(n1081), .ZN(n1079) );
NAND2_X1 U773 ( .A1(n1082), .A2(n1083), .ZN(n1078) );
NAND2_X1 U774 ( .A1(KEYINPUT63), .A2(n1084), .ZN(n1047) );
NAND4_X1 U775 ( .A1(n1054), .A2(n1050), .A3(n1069), .A4(n1085), .ZN(n1084) );
NOR2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XNOR2_X1 U777 ( .A(KEYINPUT14), .B(n1088), .ZN(n1050) );
NAND4_X1 U778 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1043) );
NOR4_X1 U779 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1092) );
XNOR2_X1 U780 ( .A(n1097), .B(n1098), .ZN(n1096) );
XNOR2_X1 U781 ( .A(KEYINPUT6), .B(n1099), .ZN(n1095) );
NOR2_X1 U782 ( .A1(n1082), .A2(n1100), .ZN(n1091) );
XOR2_X1 U783 ( .A(n1101), .B(n1102), .Z(n1090) );
NOR2_X1 U784 ( .A1(n1103), .A2(KEYINPUT47), .ZN(n1102) );
XOR2_X1 U785 ( .A(KEYINPUT29), .B(n1104), .Z(n1089) );
NOR2_X1 U786 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U787 ( .A(n1107), .B(KEYINPUT59), .Z(n1106) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U789 ( .A(n1110), .B(KEYINPUT13), .ZN(n1108) );
NOR2_X1 U790 ( .A1(n1110), .A2(n1109), .ZN(n1105) );
XOR2_X1 U791 ( .A(n1111), .B(n1112), .Z(G72) );
NAND2_X1 U792 ( .A1(G953), .A2(n1113), .ZN(n1112) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1113) );
NAND3_X1 U794 ( .A1(n1114), .A2(n1115), .A3(KEYINPUT42), .ZN(n1111) );
NAND2_X1 U795 ( .A1(KEYINPUT18), .A2(n1116), .ZN(n1115) );
NAND3_X1 U796 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1116) );
OR2_X1 U797 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND3_X1 U798 ( .A1(n1120), .A2(n1121), .A3(n1044), .ZN(n1118) );
NAND2_X1 U799 ( .A1(G953), .A2(n1122), .ZN(n1117) );
NAND2_X1 U800 ( .A1(G900), .A2(n1120), .ZN(n1122) );
OR4_X1 U801 ( .A1(n1123), .A2(G953), .A3(n1120), .A4(KEYINPUT18), .ZN(n1114) );
NAND2_X1 U802 ( .A1(n1124), .A2(n1125), .ZN(n1120) );
NAND2_X1 U803 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
OR2_X1 U804 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U805 ( .A1(n1130), .A2(n1131), .ZN(n1124) );
INV_X1 U806 ( .A(n1126), .ZN(n1131) );
XNOR2_X1 U807 ( .A(n1132), .B(n1133), .ZN(n1126) );
NOR2_X1 U808 ( .A1(KEYINPUT32), .A2(n1134), .ZN(n1133) );
NAND2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
OR2_X1 U810 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U811 ( .A(n1139), .B(KEYINPUT50), .Z(n1135) );
NAND2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1139) );
XOR2_X1 U813 ( .A(G137), .B(n1140), .Z(n1137) );
NOR2_X1 U814 ( .A1(G134), .A2(KEYINPUT3), .ZN(n1140) );
XNOR2_X1 U815 ( .A(G140), .B(G125), .ZN(n1130) );
INV_X1 U816 ( .A(n1121), .ZN(n1123) );
NAND2_X1 U817 ( .A1(n1141), .A2(n1142), .ZN(G69) );
NAND2_X1 U818 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U819 ( .A1(G953), .A2(n1145), .ZN(n1144) );
NAND3_X1 U820 ( .A1(G953), .A2(n1146), .A3(n1147), .ZN(n1141) );
INV_X1 U821 ( .A(n1143), .ZN(n1147) );
XNOR2_X1 U822 ( .A(n1148), .B(n1149), .ZN(n1143) );
NOR3_X1 U823 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1149) );
NOR2_X1 U824 ( .A1(G898), .A2(n1044), .ZN(n1152) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
XOR2_X1 U826 ( .A(n1155), .B(KEYINPUT23), .Z(n1150) );
NAND2_X1 U827 ( .A1(n1153), .A2(n1156), .ZN(n1155) );
XNOR2_X1 U828 ( .A(KEYINPUT51), .B(n1154), .ZN(n1156) );
XOR2_X1 U829 ( .A(n1157), .B(n1158), .Z(n1154) );
XNOR2_X1 U830 ( .A(n1159), .B(KEYINPUT7), .ZN(n1158) );
NAND2_X1 U831 ( .A1(KEYINPUT35), .A2(n1160), .ZN(n1159) );
XNOR2_X1 U832 ( .A(G110), .B(n1161), .ZN(n1153) );
NAND3_X1 U833 ( .A1(n1162), .A2(n1044), .A3(KEYINPUT58), .ZN(n1148) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1146) );
NOR2_X1 U835 ( .A1(n1163), .A2(n1164), .ZN(G66) );
XNOR2_X1 U836 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U837 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U838 ( .A1(n1163), .A2(n1169), .ZN(G63) );
XNOR2_X1 U839 ( .A(n1170), .B(n1171), .ZN(n1169) );
AND2_X1 U840 ( .A1(G478), .A2(n1172), .ZN(n1170) );
NOR2_X1 U841 ( .A1(n1163), .A2(n1173), .ZN(G60) );
NOR3_X1 U842 ( .A1(n1098), .A2(n1174), .A3(n1175), .ZN(n1173) );
AND3_X1 U843 ( .A1(n1176), .A2(G475), .A3(n1172), .ZN(n1175) );
NOR2_X1 U844 ( .A1(n1177), .A2(n1176), .ZN(n1174) );
NOR2_X1 U845 ( .A1(n1049), .A2(n1097), .ZN(n1177) );
XNOR2_X1 U846 ( .A(G104), .B(n1178), .ZN(G6) );
NAND2_X1 U847 ( .A1(KEYINPUT53), .A2(n1179), .ZN(n1178) );
INV_X1 U848 ( .A(n1180), .ZN(n1179) );
NOR2_X1 U849 ( .A1(n1163), .A2(n1181), .ZN(G57) );
XOR2_X1 U850 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U851 ( .A(n1184), .B(n1185), .ZN(n1183) );
XOR2_X1 U852 ( .A(n1186), .B(n1187), .Z(n1182) );
AND2_X1 U853 ( .A1(G472), .A2(n1172), .ZN(n1187) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
NOR2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U856 ( .A1(KEYINPUT28), .A2(n1192), .ZN(n1191) );
NOR2_X1 U857 ( .A1(n1193), .A2(n1194), .ZN(n1190) );
AND2_X1 U858 ( .A1(n1192), .A2(KEYINPUT19), .ZN(n1193) );
NOR4_X1 U859 ( .A1(KEYINPUT28), .A2(KEYINPUT19), .A3(n1192), .A4(n1194), .ZN(n1188) );
NOR2_X1 U860 ( .A1(n1163), .A2(n1195), .ZN(G54) );
XOR2_X1 U861 ( .A(n1196), .B(n1197), .Z(n1195) );
XOR2_X1 U862 ( .A(n1198), .B(n1199), .Z(n1197) );
NOR2_X1 U863 ( .A1(n1109), .A2(n1168), .ZN(n1198) );
INV_X1 U864 ( .A(n1172), .ZN(n1168) );
XOR2_X1 U865 ( .A(n1200), .B(n1201), .Z(n1196) );
NAND2_X1 U866 ( .A1(n1202), .A2(KEYINPUT60), .ZN(n1201) );
XNOR2_X1 U867 ( .A(G140), .B(n1203), .ZN(n1202) );
NAND2_X1 U868 ( .A1(KEYINPUT25), .A2(n1204), .ZN(n1200) );
XOR2_X1 U869 ( .A(KEYINPUT36), .B(n1205), .Z(n1204) );
NOR2_X1 U870 ( .A1(n1163), .A2(n1206), .ZN(G51) );
XOR2_X1 U871 ( .A(n1207), .B(n1208), .Z(n1206) );
NAND2_X1 U872 ( .A1(n1172), .A2(n1101), .ZN(n1208) );
NOR2_X1 U873 ( .A1(n1209), .A2(n1049), .ZN(n1172) );
NOR2_X1 U874 ( .A1(n1162), .A2(n1121), .ZN(n1049) );
NAND4_X1 U875 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1121) );
NOR4_X1 U876 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
INV_X1 U877 ( .A(n1218), .ZN(n1215) );
NOR2_X1 U878 ( .A1(n1219), .A2(n1220), .ZN(n1212) );
NOR3_X1 U879 ( .A1(n1087), .A2(n1086), .A3(n1221), .ZN(n1220) );
INV_X1 U880 ( .A(n1063), .ZN(n1086) );
INV_X1 U881 ( .A(n1222), .ZN(n1219) );
NAND4_X1 U882 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1162) );
AND4_X1 U883 ( .A1(n1180), .A2(n1042), .A3(n1227), .A4(n1228), .ZN(n1226) );
NAND4_X1 U884 ( .A1(n1069), .A2(n1062), .A3(n1054), .A4(n1229), .ZN(n1042) );
NAND4_X1 U885 ( .A1(n1061), .A2(n1069), .A3(n1054), .A4(n1229), .ZN(n1180) );
AND2_X1 U886 ( .A1(n1230), .A2(n1231), .ZN(n1225) );
NAND2_X1 U887 ( .A1(n1232), .A2(KEYINPUT27), .ZN(n1207) );
XOR2_X1 U888 ( .A(n1233), .B(n1234), .Z(n1232) );
NOR2_X1 U889 ( .A1(KEYINPUT17), .A2(n1235), .ZN(n1234) );
NOR2_X1 U890 ( .A1(n1044), .A2(G952), .ZN(n1163) );
XNOR2_X1 U891 ( .A(G146), .B(n1210), .ZN(G48) );
NAND3_X1 U892 ( .A1(n1061), .A2(n1081), .A3(n1236), .ZN(n1210) );
XNOR2_X1 U893 ( .A(G143), .B(n1211), .ZN(G45) );
NAND4_X1 U894 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1081), .ZN(n1211) );
XNOR2_X1 U895 ( .A(G140), .B(n1222), .ZN(G42) );
NAND4_X1 U896 ( .A1(n1056), .A2(n1240), .A3(n1099), .A4(n1061), .ZN(n1222) );
XNOR2_X1 U897 ( .A(G137), .B(n1241), .ZN(G39) );
NAND4_X1 U898 ( .A1(KEYINPUT31), .A2(n1056), .A3(n1236), .A4(n1063), .ZN(n1241) );
XNOR2_X1 U899 ( .A(n1217), .B(n1242), .ZN(G36) );
XOR2_X1 U900 ( .A(KEYINPUT0), .B(G134), .Z(n1242) );
AND3_X1 U901 ( .A1(n1238), .A2(n1062), .A3(n1056), .ZN(n1217) );
XOR2_X1 U902 ( .A(n1216), .B(n1243), .Z(G33) );
NOR2_X1 U903 ( .A1(KEYINPUT40), .A2(n1138), .ZN(n1243) );
AND3_X1 U904 ( .A1(n1238), .A2(n1061), .A3(n1056), .ZN(n1216) );
INV_X1 U905 ( .A(n1087), .ZN(n1056) );
NAND2_X1 U906 ( .A1(n1083), .A2(n1244), .ZN(n1087) );
AND3_X1 U907 ( .A1(n1069), .A2(n1245), .A3(n1075), .ZN(n1238) );
XNOR2_X1 U908 ( .A(G128), .B(n1218), .ZN(G30) );
NAND3_X1 U909 ( .A1(n1062), .A2(n1081), .A3(n1236), .ZN(n1218) );
INV_X1 U910 ( .A(n1221), .ZN(n1236) );
NAND2_X1 U911 ( .A1(n1240), .A2(n1246), .ZN(n1221) );
AND3_X1 U912 ( .A1(n1093), .A2(n1245), .A3(n1069), .ZN(n1240) );
XNOR2_X1 U913 ( .A(G101), .B(n1223), .ZN(G3) );
NAND3_X1 U914 ( .A1(n1247), .A2(n1069), .A3(n1075), .ZN(n1223) );
NAND2_X1 U915 ( .A1(n1248), .A2(n1249), .ZN(G27) );
NAND2_X1 U916 ( .A1(n1214), .A2(n1235), .ZN(n1249) );
XOR2_X1 U917 ( .A(KEYINPUT33), .B(n1250), .Z(n1248) );
NOR2_X1 U918 ( .A1(n1214), .A2(n1235), .ZN(n1250) );
AND4_X1 U919 ( .A1(n1061), .A2(n1059), .A3(n1251), .A4(n1076), .ZN(n1214) );
AND2_X1 U920 ( .A1(n1245), .A2(n1081), .ZN(n1251) );
NAND2_X1 U921 ( .A1(n1252), .A2(n1253), .ZN(n1245) );
XOR2_X1 U922 ( .A(n1254), .B(KEYINPUT39), .Z(n1252) );
NAND3_X1 U923 ( .A1(n1088), .A2(n1255), .A3(n1256), .ZN(n1254) );
INV_X1 U924 ( .A(G900), .ZN(n1255) );
NAND3_X1 U925 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(G24) );
NAND2_X1 U926 ( .A1(KEYINPUT15), .A2(n1228), .ZN(n1259) );
OR3_X1 U927 ( .A1(n1228), .A2(KEYINPUT15), .A3(G122), .ZN(n1258) );
NAND2_X1 U928 ( .A1(G122), .A2(n1260), .ZN(n1257) );
NAND2_X1 U929 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
INV_X1 U930 ( .A(KEYINPUT15), .ZN(n1262) );
XOR2_X1 U931 ( .A(n1228), .B(KEYINPUT45), .Z(n1261) );
NAND4_X1 U932 ( .A1(n1239), .A2(n1229), .A3(n1054), .A4(n1263), .ZN(n1228) );
AND2_X1 U933 ( .A1(n1059), .A2(n1237), .ZN(n1263) );
NOR2_X1 U934 ( .A1(n1264), .A2(n1093), .ZN(n1054) );
XNOR2_X1 U935 ( .A(G119), .B(n1265), .ZN(G21) );
NAND2_X1 U936 ( .A1(KEYINPUT21), .A2(n1266), .ZN(n1265) );
INV_X1 U937 ( .A(n1224), .ZN(n1266) );
NAND4_X1 U938 ( .A1(n1246), .A2(n1059), .A3(n1247), .A4(n1093), .ZN(n1224) );
XNOR2_X1 U939 ( .A(n1264), .B(KEYINPUT41), .ZN(n1246) );
XNOR2_X1 U940 ( .A(G116), .B(n1231), .ZN(G18) );
NAND4_X1 U941 ( .A1(n1075), .A2(n1059), .A3(n1062), .A4(n1229), .ZN(n1231) );
AND2_X1 U942 ( .A1(n1239), .A2(n1267), .ZN(n1062) );
XNOR2_X1 U943 ( .A(G113), .B(n1227), .ZN(G15) );
NAND4_X1 U944 ( .A1(n1061), .A2(n1075), .A3(n1059), .A4(n1229), .ZN(n1227) );
NOR2_X1 U945 ( .A1(n1067), .A2(n1100), .ZN(n1059) );
INV_X1 U946 ( .A(n1068), .ZN(n1100) );
NOR2_X1 U947 ( .A1(n1093), .A2(n1099), .ZN(n1075) );
NOR2_X1 U948 ( .A1(n1267), .A2(n1239), .ZN(n1061) );
XNOR2_X1 U949 ( .A(G110), .B(n1230), .ZN(G12) );
NAND3_X1 U950 ( .A1(n1076), .A2(n1069), .A3(n1247), .ZN(n1230) );
AND2_X1 U951 ( .A1(n1063), .A2(n1229), .ZN(n1247) );
AND2_X1 U952 ( .A1(n1081), .A2(n1268), .ZN(n1229) );
NAND2_X1 U953 ( .A1(n1253), .A2(n1269), .ZN(n1268) );
NAND3_X1 U954 ( .A1(n1256), .A2(n1270), .A3(n1271), .ZN(n1269) );
XOR2_X1 U955 ( .A(n1088), .B(KEYINPUT2), .Z(n1271) );
INV_X1 U956 ( .A(G898), .ZN(n1270) );
AND2_X1 U957 ( .A1(n1272), .A2(G953), .ZN(n1256) );
XNOR2_X1 U958 ( .A(G902), .B(KEYINPUT4), .ZN(n1272) );
NAND3_X1 U959 ( .A1(n1088), .A2(n1044), .A3(G952), .ZN(n1253) );
NAND2_X1 U960 ( .A1(G237), .A2(G234), .ZN(n1088) );
NOR2_X1 U961 ( .A1(n1083), .A2(n1082), .ZN(n1081) );
INV_X1 U962 ( .A(n1244), .ZN(n1082) );
NAND2_X1 U963 ( .A1(G214), .A2(n1273), .ZN(n1244) );
XNOR2_X1 U964 ( .A(n1103), .B(n1101), .ZN(n1083) );
AND2_X1 U965 ( .A1(G210), .A2(n1273), .ZN(n1101) );
NAND2_X1 U966 ( .A1(n1274), .A2(n1209), .ZN(n1273) );
XNOR2_X1 U967 ( .A(KEYINPUT20), .B(n1275), .ZN(n1274) );
AND2_X1 U968 ( .A1(n1276), .A2(n1209), .ZN(n1103) );
XNOR2_X1 U969 ( .A(G125), .B(n1233), .ZN(n1276) );
XOR2_X1 U970 ( .A(n1277), .B(n1278), .Z(n1233) );
XNOR2_X1 U971 ( .A(n1194), .B(n1279), .ZN(n1278) );
XOR2_X1 U972 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U973 ( .A(n1282), .B(n1283), .Z(n1277) );
XOR2_X1 U974 ( .A(G110), .B(n1284), .Z(n1283) );
NOR2_X1 U975 ( .A1(G953), .A2(n1145), .ZN(n1284) );
INV_X1 U976 ( .A(G224), .ZN(n1145) );
NAND2_X1 U977 ( .A1(KEYINPUT49), .A2(n1157), .ZN(n1282) );
XNOR2_X1 U978 ( .A(n1285), .B(n1286), .ZN(n1157) );
NAND2_X1 U979 ( .A1(n1287), .A2(KEYINPUT11), .ZN(n1285) );
XNOR2_X1 U980 ( .A(G107), .B(n1288), .ZN(n1287) );
NOR2_X1 U981 ( .A1(G104), .A2(KEYINPUT43), .ZN(n1288) );
NOR2_X1 U982 ( .A1(n1239), .A2(n1237), .ZN(n1063) );
INV_X1 U983 ( .A(n1267), .ZN(n1237) );
XNOR2_X1 U984 ( .A(n1289), .B(n1098), .ZN(n1267) );
NOR2_X1 U985 ( .A1(n1176), .A2(G902), .ZN(n1098) );
XOR2_X1 U986 ( .A(n1290), .B(n1291), .Z(n1176) );
XNOR2_X1 U987 ( .A(n1292), .B(n1293), .ZN(n1291) );
NAND2_X1 U988 ( .A1(n1294), .A2(n1295), .ZN(n1292) );
INV_X1 U989 ( .A(n1128), .ZN(n1295) );
XNOR2_X1 U990 ( .A(n1129), .B(KEYINPUT22), .ZN(n1294) );
XOR2_X1 U991 ( .A(n1296), .B(n1297), .Z(n1290) );
NOR2_X1 U992 ( .A1(KEYINPUT8), .A2(n1298), .ZN(n1297) );
NOR2_X1 U993 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NOR2_X1 U994 ( .A1(G104), .A2(n1301), .ZN(n1300) );
NOR2_X1 U995 ( .A1(n1302), .A2(KEYINPUT62), .ZN(n1301) );
NOR2_X1 U996 ( .A1(KEYINPUT52), .A2(n1303), .ZN(n1302) );
INV_X1 U997 ( .A(n1304), .ZN(n1303) );
NOR2_X1 U998 ( .A1(n1305), .A2(n1304), .ZN(n1299) );
XOR2_X1 U999 ( .A(G113), .B(n1161), .Z(n1304) );
NOR2_X1 U1000 ( .A1(n1306), .A2(KEYINPUT52), .ZN(n1305) );
NOR2_X1 U1001 ( .A1(KEYINPUT62), .A2(n1307), .ZN(n1306) );
INV_X1 U1002 ( .A(G104), .ZN(n1307) );
XNOR2_X1 U1003 ( .A(n1308), .B(n1138), .ZN(n1296) );
INV_X1 U1004 ( .A(G131), .ZN(n1138) );
NAND3_X1 U1005 ( .A1(G214), .A2(n1044), .A3(n1309), .ZN(n1308) );
XNOR2_X1 U1006 ( .A(G237), .B(KEYINPUT9), .ZN(n1309) );
NAND2_X1 U1007 ( .A1(KEYINPUT37), .A2(n1097), .ZN(n1289) );
INV_X1 U1008 ( .A(G475), .ZN(n1097) );
XNOR2_X1 U1009 ( .A(n1094), .B(KEYINPUT16), .ZN(n1239) );
XNOR2_X1 U1010 ( .A(n1310), .B(G478), .ZN(n1094) );
NAND2_X1 U1011 ( .A1(n1311), .A2(n1171), .ZN(n1310) );
XOR2_X1 U1012 ( .A(n1312), .B(n1313), .Z(n1171) );
XOR2_X1 U1013 ( .A(n1314), .B(n1315), .Z(n1313) );
XNOR2_X1 U1014 ( .A(G107), .B(G134), .ZN(n1315) );
NAND3_X1 U1015 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1314) );
NAND2_X1 U1016 ( .A1(G143), .A2(n1319), .ZN(n1318) );
NAND2_X1 U1017 ( .A1(KEYINPUT5), .A2(n1320), .ZN(n1317) );
NAND2_X1 U1018 ( .A1(n1321), .A2(G128), .ZN(n1320) );
XNOR2_X1 U1019 ( .A(KEYINPUT44), .B(G143), .ZN(n1321) );
NAND2_X1 U1020 ( .A1(n1322), .A2(n1323), .ZN(n1316) );
INV_X1 U1021 ( .A(KEYINPUT5), .ZN(n1323) );
NAND2_X1 U1022 ( .A1(n1324), .A2(n1325), .ZN(n1322) );
OR3_X1 U1023 ( .A1(n1319), .A2(G143), .A3(KEYINPUT44), .ZN(n1325) );
NAND2_X1 U1024 ( .A1(KEYINPUT44), .A2(G143), .ZN(n1324) );
XNOR2_X1 U1025 ( .A(n1280), .B(n1326), .ZN(n1312) );
AND2_X1 U1026 ( .A1(n1327), .A2(G217), .ZN(n1326) );
XOR2_X1 U1027 ( .A(G116), .B(n1161), .Z(n1280) );
XOR2_X1 U1028 ( .A(G122), .B(KEYINPUT10), .Z(n1161) );
XNOR2_X1 U1029 ( .A(G902), .B(KEYINPUT12), .ZN(n1311) );
AND2_X1 U1030 ( .A1(n1067), .A2(n1068), .ZN(n1069) );
NAND2_X1 U1031 ( .A1(G221), .A2(n1328), .ZN(n1068) );
XNOR2_X1 U1032 ( .A(n1110), .B(n1109), .ZN(n1067) );
INV_X1 U1033 ( .A(G469), .ZN(n1109) );
AND2_X1 U1034 ( .A1(n1329), .A2(n1209), .ZN(n1110) );
XOR2_X1 U1035 ( .A(n1330), .B(n1199), .Z(n1329) );
XNOR2_X1 U1036 ( .A(n1192), .B(KEYINPUT54), .ZN(n1199) );
INV_X1 U1037 ( .A(n1331), .ZN(n1192) );
XOR2_X1 U1038 ( .A(n1332), .B(n1205), .Z(n1330) );
XNOR2_X1 U1039 ( .A(n1333), .B(n1134), .ZN(n1205) );
NAND2_X1 U1040 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1041 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XNOR2_X1 U1042 ( .A(KEYINPUT55), .B(n1286), .ZN(n1337) );
XNOR2_X1 U1043 ( .A(n1338), .B(G104), .ZN(n1336) );
INV_X1 U1044 ( .A(G107), .ZN(n1338) );
XOR2_X1 U1045 ( .A(n1339), .B(KEYINPUT24), .Z(n1334) );
NAND2_X1 U1046 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XNOR2_X1 U1047 ( .A(KEYINPUT55), .B(G101), .ZN(n1341) );
XNOR2_X1 U1048 ( .A(G107), .B(G104), .ZN(n1340) );
NAND3_X1 U1049 ( .A1(n1342), .A2(n1343), .A3(KEYINPUT38), .ZN(n1332) );
NAND2_X1 U1050 ( .A1(n1203), .A2(n1344), .ZN(n1343) );
NAND2_X1 U1051 ( .A1(n1345), .A2(G140), .ZN(n1342) );
XOR2_X1 U1052 ( .A(KEYINPUT56), .B(n1203), .Z(n1345) );
XOR2_X1 U1053 ( .A(G110), .B(n1346), .Z(n1203) );
AND2_X1 U1054 ( .A1(n1044), .A2(G227), .ZN(n1346) );
AND2_X1 U1055 ( .A1(n1099), .A2(n1093), .ZN(n1076) );
XOR2_X1 U1056 ( .A(n1347), .B(n1167), .Z(n1093) );
NAND2_X1 U1057 ( .A1(G217), .A2(n1328), .ZN(n1167) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1209), .ZN(n1328) );
NAND2_X1 U1059 ( .A1(n1165), .A2(n1209), .ZN(n1347) );
XNOR2_X1 U1060 ( .A(n1348), .B(n1349), .ZN(n1165) );
XNOR2_X1 U1061 ( .A(n1350), .B(n1351), .ZN(n1349) );
NAND2_X1 U1062 ( .A1(n1327), .A2(G221), .ZN(n1350) );
AND2_X1 U1063 ( .A1(G234), .A2(n1044), .ZN(n1327) );
XOR2_X1 U1064 ( .A(n1352), .B(n1353), .Z(n1348) );
NOR2_X1 U1065 ( .A1(KEYINPUT57), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1066 ( .A(n1355), .B(G110), .Z(n1354) );
NAND3_X1 U1067 ( .A1(n1356), .A2(n1357), .A3(KEYINPUT30), .ZN(n1355) );
NAND2_X1 U1068 ( .A1(KEYINPUT46), .A2(n1358), .ZN(n1357) );
XNOR2_X1 U1069 ( .A(G119), .B(G128), .ZN(n1358) );
NAND3_X1 U1070 ( .A1(G119), .A2(n1319), .A3(n1359), .ZN(n1356) );
INV_X1 U1071 ( .A(KEYINPUT46), .ZN(n1359) );
INV_X1 U1072 ( .A(G128), .ZN(n1319) );
XNOR2_X1 U1073 ( .A(G137), .B(n1360), .ZN(n1352) );
NOR2_X1 U1074 ( .A1(n1128), .A2(n1361), .ZN(n1360) );
XOR2_X1 U1075 ( .A(n1362), .B(KEYINPUT34), .Z(n1361) );
NAND2_X1 U1076 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
OR2_X1 U1077 ( .A1(G125), .A2(KEYINPUT1), .ZN(n1364) );
NAND2_X1 U1078 ( .A1(n1129), .A2(KEYINPUT1), .ZN(n1363) );
NOR2_X1 U1079 ( .A1(n1235), .A2(G140), .ZN(n1129) );
INV_X1 U1080 ( .A(G125), .ZN(n1235) );
NOR2_X1 U1081 ( .A1(n1344), .A2(G125), .ZN(n1128) );
INV_X1 U1082 ( .A(G140), .ZN(n1344) );
INV_X1 U1083 ( .A(n1264), .ZN(n1099) );
XNOR2_X1 U1084 ( .A(n1365), .B(G472), .ZN(n1264) );
NAND2_X1 U1085 ( .A1(n1366), .A2(n1209), .ZN(n1365) );
INV_X1 U1086 ( .A(G902), .ZN(n1209) );
XNOR2_X1 U1087 ( .A(n1367), .B(n1184), .ZN(n1366) );
XOR2_X1 U1088 ( .A(n1368), .B(n1286), .Z(n1184) );
INV_X1 U1089 ( .A(G101), .ZN(n1286) );
NAND3_X1 U1090 ( .A1(n1275), .A2(n1044), .A3(G210), .ZN(n1368) );
INV_X1 U1091 ( .A(G953), .ZN(n1044) );
INV_X1 U1092 ( .A(G237), .ZN(n1275) );
NAND2_X1 U1093 ( .A1(n1369), .A2(n1370), .ZN(n1367) );
NAND2_X1 U1094 ( .A1(n1185), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1095 ( .A(n1372), .B(KEYINPUT48), .Z(n1369) );
OR2_X1 U1096 ( .A1(n1371), .A2(n1185), .ZN(n1372) );
INV_X1 U1097 ( .A(n1160), .ZN(n1185) );
XOR2_X1 U1098 ( .A(G116), .B(n1281), .Z(n1160) );
XNOR2_X1 U1099 ( .A(n1373), .B(G119), .ZN(n1281) );
INV_X1 U1100 ( .A(G113), .ZN(n1373) );
XNOR2_X1 U1101 ( .A(n1331), .B(n1194), .ZN(n1371) );
INV_X1 U1102 ( .A(n1134), .ZN(n1194) );
XOR2_X1 U1103 ( .A(G128), .B(n1293), .Z(n1134) );
XOR2_X1 U1104 ( .A(G143), .B(n1351), .Z(n1293) );
XOR2_X1 U1105 ( .A(G146), .B(KEYINPUT26), .Z(n1351) );
XOR2_X1 U1106 ( .A(G131), .B(n1374), .Z(n1331) );
XOR2_X1 U1107 ( .A(G137), .B(G134), .Z(n1374) );
endmodule


