//Key = 0010101100001011010011101000010101011000110010100110100000011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360;

XOR2_X1 U750 ( .A(n1039), .B(n1040), .Z(G9) );
NAND3_X1 U751 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR4_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
INV_X1 U754 ( .A(G952), .ZN(n1049) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
XOR2_X1 U756 ( .A(KEYINPUT21), .B(n1052), .Z(n1051) );
AND4_X1 U757 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NAND4_X1 U758 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1046) );
NAND4_X1 U759 ( .A1(n1061), .A2(n1053), .A3(n1062), .A4(n1063), .ZN(n1058) );
AND3_X1 U760 ( .A1(n1054), .A2(n1064), .A3(n1041), .ZN(n1063) );
XOR2_X1 U761 ( .A(n1050), .B(KEYINPUT29), .Z(n1062) );
XNOR2_X1 U762 ( .A(n1042), .B(KEYINPUT33), .ZN(n1061) );
NAND4_X1 U763 ( .A1(n1053), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1057) );
NAND2_X1 U764 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U765 ( .A1(n1055), .A2(n1069), .ZN(n1068) );
NAND3_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1054), .ZN(n1065) );
NAND2_X1 U767 ( .A1(n1055), .A2(n1072), .ZN(n1071) );
NAND2_X1 U768 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
OR2_X1 U769 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
INV_X1 U770 ( .A(n1077), .ZN(n1073) );
AND2_X1 U771 ( .A1(n1042), .A2(n1078), .ZN(n1055) );
NAND2_X1 U772 ( .A1(n1069), .A2(n1079), .ZN(n1070) );
NAND2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1082), .ZN(n1081) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1042), .ZN(n1080) );
NOR2_X1 U776 ( .A1(KEYINPUT57), .A2(n1084), .ZN(n1053) );
INV_X1 U777 ( .A(n1085), .ZN(n1084) );
NOR3_X1 U778 ( .A1(n1086), .A2(G953), .A3(n1087), .ZN(n1044) );
INV_X1 U779 ( .A(n1059), .ZN(n1087) );
NAND4_X1 U780 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1059) );
NOR3_X1 U781 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
XOR2_X1 U782 ( .A(n1095), .B(KEYINPUT52), .Z(n1094) );
NAND2_X1 U783 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U784 ( .A1(n1096), .A2(n1097), .ZN(n1093) );
NAND3_X1 U785 ( .A1(n1098), .A2(n1075), .A3(n1064), .ZN(n1092) );
NOR3_X1 U786 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1090) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1089) );
XOR2_X1 U788 ( .A(n1104), .B(KEYINPUT53), .Z(n1088) );
XOR2_X1 U789 ( .A(KEYINPUT10), .B(G952), .Z(n1086) );
NAND2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(G72) );
NAND3_X1 U791 ( .A1(G953), .A2(n1107), .A3(n1108), .ZN(n1106) );
XOR2_X1 U792 ( .A(KEYINPUT20), .B(n1109), .Z(n1105) );
NOR2_X1 U793 ( .A1(n1110), .A2(n1108), .ZN(n1109) );
XOR2_X1 U794 ( .A(n1111), .B(n1112), .Z(n1108) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U796 ( .A(n1060), .B(KEYINPUT22), .Z(n1114) );
INV_X1 U797 ( .A(n1115), .ZN(n1113) );
NAND3_X1 U798 ( .A1(n1116), .A2(n1117), .A3(KEYINPUT6), .ZN(n1111) );
NAND2_X1 U799 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1116) );
NOR2_X1 U801 ( .A1(KEYINPUT0), .A2(n1121), .ZN(n1119) );
XOR2_X1 U802 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND2_X1 U803 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
XNOR2_X1 U804 ( .A(n1126), .B(n1127), .ZN(n1125) );
NAND2_X1 U805 ( .A1(KEYINPUT4), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U806 ( .A(KEYINPUT54), .B(KEYINPUT27), .ZN(n1124) );
AND2_X1 U807 ( .A1(n1107), .A2(G953), .ZN(n1110) );
NAND2_X1 U808 ( .A1(G900), .A2(G227), .ZN(n1107) );
NAND2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(G69) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U811 ( .A(n1133), .B(KEYINPUT38), .Z(n1131) );
NAND2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(n1129) );
XOR2_X1 U813 ( .A(KEYINPUT7), .B(n1132), .Z(n1135) );
AND2_X1 U814 ( .A1(G953), .A2(n1136), .ZN(n1132) );
NAND2_X1 U815 ( .A1(G898), .A2(G224), .ZN(n1136) );
XNOR2_X1 U816 ( .A(n1137), .B(n1133), .ZN(n1134) );
NAND2_X1 U817 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
NAND2_X1 U818 ( .A1(G953), .A2(n1140), .ZN(n1139) );
XOR2_X1 U819 ( .A(n1141), .B(KEYINPUT19), .Z(n1138) );
NAND2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
NAND2_X1 U821 ( .A1(n1144), .A2(n1060), .ZN(n1143) );
INV_X1 U822 ( .A(KEYINPUT38), .ZN(n1142) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1146), .ZN(G66) );
XOR2_X1 U824 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U825 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
NOR2_X1 U826 ( .A1(n1145), .A2(n1151), .ZN(G63) );
NOR2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U828 ( .A(KEYINPUT56), .B(n1154), .Z(n1153) );
AND2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U830 ( .A1(n1156), .A2(n1155), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1150), .A2(n1097), .ZN(n1156) );
INV_X1 U832 ( .A(G478), .ZN(n1097) );
NOR2_X1 U833 ( .A1(n1145), .A2(n1157), .ZN(G60) );
NOR3_X1 U834 ( .A1(n1102), .A2(n1158), .A3(n1159), .ZN(n1157) );
NOR3_X1 U835 ( .A1(n1160), .A2(n1103), .A3(n1150), .ZN(n1159) );
INV_X1 U836 ( .A(G475), .ZN(n1103) );
INV_X1 U837 ( .A(n1161), .ZN(n1160) );
NOR2_X1 U838 ( .A1(n1162), .A2(n1161), .ZN(n1158) );
AND2_X1 U839 ( .A1(n1047), .A2(G475), .ZN(n1162) );
XOR2_X1 U840 ( .A(G104), .B(n1163), .Z(G6) );
NOR2_X1 U841 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR3_X1 U842 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(G57) );
NOR3_X1 U843 ( .A1(n1169), .A2(G953), .A3(G952), .ZN(n1168) );
AND2_X1 U844 ( .A1(n1169), .A2(n1145), .ZN(n1167) );
INV_X1 U845 ( .A(KEYINPUT34), .ZN(n1169) );
XOR2_X1 U846 ( .A(n1170), .B(n1171), .Z(n1166) );
NOR2_X1 U847 ( .A1(KEYINPUT42), .A2(n1172), .ZN(n1171) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U849 ( .A(n1175), .B(n1176), .ZN(n1173) );
NOR2_X1 U850 ( .A1(n1177), .A2(n1150), .ZN(n1176) );
INV_X1 U851 ( .A(G472), .ZN(n1177) );
XNOR2_X1 U852 ( .A(G101), .B(n1178), .ZN(n1170) );
NOR3_X1 U853 ( .A1(n1145), .A2(n1179), .A3(n1180), .ZN(G54) );
NOR2_X1 U854 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U855 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U856 ( .A1(KEYINPUT35), .A2(n1185), .ZN(n1183) );
INV_X1 U857 ( .A(KEYINPUT55), .ZN(n1181) );
NOR2_X1 U858 ( .A1(KEYINPUT55), .A2(n1186), .ZN(n1179) );
XOR2_X1 U859 ( .A(n1187), .B(n1184), .Z(n1186) );
XNOR2_X1 U860 ( .A(n1188), .B(n1189), .ZN(n1184) );
XOR2_X1 U861 ( .A(n1190), .B(n1191), .Z(n1189) );
NAND2_X1 U862 ( .A1(KEYINPUT60), .A2(n1123), .ZN(n1190) );
XOR2_X1 U863 ( .A(n1192), .B(n1193), .Z(n1188) );
NOR2_X1 U864 ( .A1(n1194), .A2(n1150), .ZN(n1193) );
INV_X1 U865 ( .A(G469), .ZN(n1194) );
NAND2_X1 U866 ( .A1(KEYINPUT63), .A2(n1175), .ZN(n1192) );
NAND2_X1 U867 ( .A1(KEYINPUT35), .A2(n1195), .ZN(n1187) );
INV_X1 U868 ( .A(n1185), .ZN(n1195) );
NOR2_X1 U869 ( .A1(n1145), .A2(n1196), .ZN(G51) );
XNOR2_X1 U870 ( .A(n1197), .B(n1198), .ZN(n1196) );
NOR2_X1 U871 ( .A1(n1199), .A2(n1150), .ZN(n1198) );
NAND2_X1 U872 ( .A1(G902), .A2(n1047), .ZN(n1150) );
NAND3_X1 U873 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1047) );
INV_X1 U874 ( .A(n1144), .ZN(n1202) );
NAND4_X1 U875 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1144) );
NOR4_X1 U876 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
NOR2_X1 U877 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
NOR2_X1 U878 ( .A1(n1213), .A2(n1164), .ZN(n1212) );
XOR2_X1 U879 ( .A(n1165), .B(KEYINPUT25), .Z(n1213) );
NAND4_X1 U880 ( .A1(n1083), .A2(n1042), .A3(n1214), .A4(n1215), .ZN(n1165) );
NAND4_X1 U881 ( .A1(n1041), .A2(n1042), .A3(n1216), .A4(n1217), .ZN(n1204) );
NAND2_X1 U882 ( .A1(KEYINPUT41), .A2(n1218), .ZN(n1217) );
NAND2_X1 U883 ( .A1(n1219), .A2(n1220), .ZN(n1216) );
INV_X1 U884 ( .A(KEYINPUT41), .ZN(n1220) );
NAND3_X1 U885 ( .A1(n1164), .A2(n1215), .A3(n1214), .ZN(n1219) );
NAND2_X1 U886 ( .A1(n1221), .A2(n1222), .ZN(n1201) );
INV_X1 U887 ( .A(KEYINPUT12), .ZN(n1222) );
NAND2_X1 U888 ( .A1(KEYINPUT12), .A2(n1115), .ZN(n1200) );
NAND4_X1 U889 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1115) );
AND3_X1 U890 ( .A1(n1227), .A2(n1221), .A3(n1228), .ZN(n1226) );
NAND3_X1 U891 ( .A1(n1229), .A2(n1230), .A3(n1069), .ZN(n1225) );
NAND2_X1 U892 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U893 ( .A1(n1083), .A2(n1082), .ZN(n1232) );
OR2_X1 U894 ( .A1(n1233), .A2(n1234), .ZN(n1082) );
NOR2_X1 U895 ( .A1(n1060), .A2(G952), .ZN(n1145) );
XNOR2_X1 U896 ( .A(G146), .B(n1223), .ZN(G48) );
NAND2_X1 U897 ( .A1(n1235), .A2(n1083), .ZN(n1223) );
XOR2_X1 U898 ( .A(n1236), .B(n1224), .Z(G45) );
NAND4_X1 U899 ( .A1(n1077), .A2(n1229), .A3(n1237), .A4(n1233), .ZN(n1224) );
AND2_X1 U900 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XNOR2_X1 U901 ( .A(G140), .B(n1240), .ZN(G42) );
NAND4_X1 U902 ( .A1(n1241), .A2(n1229), .A3(n1234), .A4(n1083), .ZN(n1240) );
XOR2_X1 U903 ( .A(n1050), .B(KEYINPUT2), .Z(n1241) );
XNOR2_X1 U904 ( .A(G137), .B(n1242), .ZN(G39) );
NAND4_X1 U905 ( .A1(n1069), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1242) );
OR2_X1 U906 ( .A1(n1229), .A2(KEYINPUT61), .ZN(n1245) );
NAND2_X1 U907 ( .A1(KEYINPUT61), .A2(n1246), .ZN(n1244) );
NAND2_X1 U908 ( .A1(n1247), .A2(n1214), .ZN(n1246) );
XOR2_X1 U909 ( .A(n1128), .B(n1227), .Z(G36) );
NAND4_X1 U910 ( .A1(n1069), .A2(n1229), .A3(n1233), .A4(n1041), .ZN(n1227) );
XNOR2_X1 U911 ( .A(G131), .B(n1248), .ZN(G33) );
NAND4_X1 U912 ( .A1(n1069), .A2(n1083), .A3(n1249), .A4(n1233), .ZN(n1248) );
NOR2_X1 U913 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
XNOR2_X1 U914 ( .A(n1247), .B(KEYINPUT24), .ZN(n1250) );
INV_X1 U915 ( .A(n1050), .ZN(n1069) );
NAND2_X1 U916 ( .A1(n1252), .A2(n1075), .ZN(n1050) );
INV_X1 U917 ( .A(n1076), .ZN(n1252) );
XNOR2_X1 U918 ( .A(G128), .B(n1228), .ZN(G30) );
NAND2_X1 U919 ( .A1(n1235), .A2(n1041), .ZN(n1228) );
AND4_X1 U920 ( .A1(n1253), .A2(n1229), .A3(n1077), .A4(n1099), .ZN(n1235) );
NOR2_X1 U921 ( .A1(n1251), .A2(n1247), .ZN(n1229) );
XOR2_X1 U922 ( .A(G101), .B(n1210), .Z(G3) );
AND3_X1 U923 ( .A1(n1043), .A2(n1078), .A3(n1233), .ZN(n1210) );
XNOR2_X1 U924 ( .A(G125), .B(n1221), .ZN(G27) );
NAND4_X1 U925 ( .A1(n1077), .A2(n1083), .A3(n1234), .A4(n1254), .ZN(n1221) );
NOR3_X1 U926 ( .A1(n1067), .A2(n1056), .A3(n1247), .ZN(n1254) );
AND2_X1 U927 ( .A1(n1255), .A2(n1256), .ZN(n1247) );
NAND4_X1 U928 ( .A1(G953), .A2(G902), .A3(n1085), .A4(n1118), .ZN(n1256) );
INV_X1 U929 ( .A(G900), .ZN(n1118) );
INV_X1 U930 ( .A(n1064), .ZN(n1056) );
XOR2_X1 U931 ( .A(G122), .B(n1211), .Z(G24) );
AND4_X1 U932 ( .A1(n1239), .A2(n1257), .A3(n1042), .A4(n1238), .ZN(n1211) );
NOR2_X1 U933 ( .A1(n1099), .A2(n1253), .ZN(n1042) );
XOR2_X1 U934 ( .A(G119), .B(n1209), .Z(G21) );
AND2_X1 U935 ( .A1(n1243), .A2(n1257), .ZN(n1209) );
INV_X1 U936 ( .A(n1231), .ZN(n1243) );
NAND3_X1 U937 ( .A1(n1078), .A2(n1099), .A3(n1253), .ZN(n1231) );
XOR2_X1 U938 ( .A(n1208), .B(n1258), .Z(G18) );
NOR2_X1 U939 ( .A1(KEYINPUT9), .A2(n1259), .ZN(n1258) );
INV_X1 U940 ( .A(G116), .ZN(n1259) );
AND3_X1 U941 ( .A1(n1233), .A2(n1041), .A3(n1257), .ZN(n1208) );
AND2_X1 U942 ( .A1(n1077), .A2(n1260), .ZN(n1257) );
XOR2_X1 U943 ( .A(n1164), .B(KEYINPUT44), .Z(n1077) );
XOR2_X1 U944 ( .A(n1261), .B(n1262), .Z(G15) );
XNOR2_X1 U945 ( .A(G113), .B(KEYINPUT28), .ZN(n1262) );
NAND2_X1 U946 ( .A1(KEYINPUT40), .A2(n1207), .ZN(n1261) );
AND4_X1 U947 ( .A1(n1260), .A2(n1083), .A3(n1233), .A4(n1263), .ZN(n1207) );
AND2_X1 U948 ( .A1(n1264), .A2(n1099), .ZN(n1233) );
AND2_X1 U949 ( .A1(n1265), .A2(n1239), .ZN(n1083) );
XOR2_X1 U950 ( .A(KEYINPUT58), .B(n1266), .Z(n1265) );
AND3_X1 U951 ( .A1(n1064), .A2(n1215), .A3(n1054), .ZN(n1260) );
XOR2_X1 U952 ( .A(G110), .B(n1267), .Z(G12) );
NOR2_X1 U953 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NOR2_X1 U954 ( .A1(KEYINPUT37), .A2(n1270), .ZN(n1269) );
INV_X1 U955 ( .A(n1203), .ZN(n1270) );
NOR2_X1 U956 ( .A1(KEYINPUT50), .A2(n1203), .ZN(n1268) );
NAND3_X1 U957 ( .A1(n1043), .A2(n1078), .A3(n1234), .ZN(n1203) );
NOR2_X1 U958 ( .A1(n1264), .A2(n1099), .ZN(n1234) );
XNOR2_X1 U959 ( .A(n1271), .B(G472), .ZN(n1099) );
NAND2_X1 U960 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XOR2_X1 U961 ( .A(n1274), .B(n1275), .Z(n1272) );
XOR2_X1 U962 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U963 ( .A(G101), .B(KEYINPUT36), .ZN(n1277) );
NAND2_X1 U964 ( .A1(KEYINPUT59), .A2(n1175), .ZN(n1276) );
XOR2_X1 U965 ( .A(n1278), .B(n1174), .Z(n1274) );
XNOR2_X1 U966 ( .A(n1279), .B(n1280), .ZN(n1174) );
XNOR2_X1 U967 ( .A(G113), .B(n1281), .ZN(n1279) );
NAND2_X1 U968 ( .A1(KEYINPUT15), .A2(n1178), .ZN(n1278) );
NOR3_X1 U969 ( .A1(G237), .A2(G953), .A3(n1199), .ZN(n1178) );
INV_X1 U970 ( .A(G210), .ZN(n1199) );
INV_X1 U971 ( .A(n1253), .ZN(n1264) );
XNOR2_X1 U972 ( .A(n1100), .B(KEYINPUT17), .ZN(n1253) );
XOR2_X1 U973 ( .A(n1282), .B(n1149), .Z(n1100) );
NAND2_X1 U974 ( .A1(G217), .A2(n1283), .ZN(n1149) );
OR2_X1 U975 ( .A1(n1148), .A2(G902), .ZN(n1282) );
XNOR2_X1 U976 ( .A(n1284), .B(n1285), .ZN(n1148) );
XOR2_X1 U977 ( .A(G137), .B(n1286), .Z(n1285) );
NOR2_X1 U978 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XOR2_X1 U979 ( .A(KEYINPUT13), .B(n1289), .Z(n1288) );
NOR2_X1 U980 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
AND2_X1 U981 ( .A1(n1291), .A2(n1290), .ZN(n1287) );
XOR2_X1 U982 ( .A(n1292), .B(n1293), .Z(n1290) );
NOR2_X1 U983 ( .A1(KEYINPUT43), .A2(G119), .ZN(n1293) );
XOR2_X1 U984 ( .A(G128), .B(n1294), .Z(n1292) );
NAND2_X1 U985 ( .A1(n1295), .A2(n1296), .ZN(n1291) );
NAND2_X1 U986 ( .A1(KEYINPUT16), .A2(n1297), .ZN(n1296) );
NAND2_X1 U987 ( .A1(G146), .A2(n1120), .ZN(n1297) );
NAND2_X1 U988 ( .A1(n1298), .A2(n1299), .ZN(n1295) );
INV_X1 U989 ( .A(KEYINPUT16), .ZN(n1299) );
NAND3_X1 U990 ( .A1(G234), .A2(n1060), .A3(G221), .ZN(n1284) );
NAND2_X1 U991 ( .A1(n1300), .A2(n1301), .ZN(n1078) );
OR3_X1 U992 ( .A1(n1239), .A2(n1238), .A3(KEYINPUT58), .ZN(n1301) );
NAND2_X1 U993 ( .A1(KEYINPUT58), .A2(n1041), .ZN(n1300) );
NOR2_X1 U994 ( .A1(n1239), .A2(n1266), .ZN(n1041) );
INV_X1 U995 ( .A(n1238), .ZN(n1266) );
XOR2_X1 U996 ( .A(n1096), .B(G478), .Z(n1238) );
NOR2_X1 U997 ( .A1(n1302), .A2(n1155), .ZN(n1096) );
XNOR2_X1 U998 ( .A(n1303), .B(n1304), .ZN(n1155) );
NOR3_X1 U999 ( .A1(n1305), .A2(G953), .A3(n1306), .ZN(n1304) );
XNOR2_X1 U1000 ( .A(G234), .B(KEYINPUT32), .ZN(n1306) );
INV_X1 U1001 ( .A(G217), .ZN(n1305) );
NAND2_X1 U1002 ( .A1(n1307), .A2(n1308), .ZN(n1303) );
NAND2_X1 U1003 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U1004 ( .A(KEYINPUT49), .B(n1311), .Z(n1307) );
NOR2_X1 U1005 ( .A1(n1309), .A2(n1310), .ZN(n1311) );
XOR2_X1 U1006 ( .A(G134), .B(n1312), .Z(n1310) );
NOR2_X1 U1007 ( .A1(KEYINPUT11), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1008 ( .A(n1039), .B(n1314), .Z(n1309) );
XOR2_X1 U1009 ( .A(G122), .B(G116), .Z(n1314) );
INV_X1 U1010 ( .A(G107), .ZN(n1039) );
XOR2_X1 U1011 ( .A(G902), .B(KEYINPUT30), .Z(n1302) );
XNOR2_X1 U1012 ( .A(n1102), .B(n1315), .ZN(n1239) );
NOR2_X1 U1013 ( .A1(G475), .A2(KEYINPUT5), .ZN(n1315) );
NOR2_X1 U1014 ( .A1(n1161), .A2(G902), .ZN(n1102) );
XNOR2_X1 U1015 ( .A(n1316), .B(n1317), .ZN(n1161) );
XOR2_X1 U1016 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1017 ( .A(G104), .B(n1320), .Z(n1319) );
NOR2_X1 U1018 ( .A1(KEYINPUT47), .A2(n1236), .ZN(n1320) );
XOR2_X1 U1019 ( .A(G122), .B(G113), .Z(n1318) );
XOR2_X1 U1020 ( .A(n1298), .B(n1321), .Z(n1316) );
XOR2_X1 U1021 ( .A(n1322), .B(n1323), .Z(n1321) );
NOR2_X1 U1022 ( .A1(G131), .A2(KEYINPUT8), .ZN(n1323) );
AND3_X1 U1023 ( .A1(G214), .A2(n1060), .A3(n1324), .ZN(n1322) );
XNOR2_X1 U1024 ( .A(G146), .B(n1120), .ZN(n1298) );
XOR2_X1 U1025 ( .A(G125), .B(G140), .Z(n1120) );
INV_X1 U1026 ( .A(n1218), .ZN(n1043) );
NAND3_X1 U1027 ( .A1(n1214), .A2(n1215), .A3(n1263), .ZN(n1218) );
INV_X1 U1028 ( .A(n1164), .ZN(n1263) );
NAND2_X1 U1029 ( .A1(n1075), .A2(n1076), .ZN(n1164) );
NAND2_X1 U1030 ( .A1(n1104), .A2(n1098), .ZN(n1076) );
NAND3_X1 U1031 ( .A1(n1325), .A2(n1273), .A3(n1197), .ZN(n1098) );
NAND2_X1 U1032 ( .A1(G210), .A2(n1326), .ZN(n1325) );
NAND3_X1 U1033 ( .A1(n1326), .A2(n1327), .A3(G210), .ZN(n1104) );
NAND2_X1 U1034 ( .A1(n1197), .A2(n1273), .ZN(n1327) );
XNOR2_X1 U1035 ( .A(n1328), .B(n1329), .ZN(n1197) );
XOR2_X1 U1036 ( .A(G125), .B(n1330), .Z(n1329) );
AND2_X1 U1037 ( .A1(n1060), .A2(G224), .ZN(n1330) );
XOR2_X1 U1038 ( .A(n1141), .B(n1280), .Z(n1328) );
XOR2_X1 U1039 ( .A(n1123), .B(KEYINPUT62), .Z(n1280) );
XOR2_X1 U1040 ( .A(n1331), .B(n1332), .Z(n1141) );
XOR2_X1 U1041 ( .A(n1333), .B(n1191), .Z(n1332) );
NAND3_X1 U1042 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1333) );
OR2_X1 U1043 ( .A1(n1337), .A2(G113), .ZN(n1336) );
NAND2_X1 U1044 ( .A1(KEYINPUT18), .A2(n1338), .ZN(n1335) );
NAND2_X1 U1045 ( .A1(n1339), .A2(n1337), .ZN(n1338) );
XNOR2_X1 U1046 ( .A(KEYINPUT31), .B(G113), .ZN(n1339) );
NAND2_X1 U1047 ( .A1(n1340), .A2(n1341), .ZN(n1334) );
INV_X1 U1048 ( .A(KEYINPUT18), .ZN(n1341) );
NAND2_X1 U1049 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
OR2_X1 U1050 ( .A1(G113), .A2(KEYINPUT31), .ZN(n1343) );
NAND3_X1 U1051 ( .A1(G113), .A2(n1337), .A3(KEYINPUT31), .ZN(n1342) );
XNOR2_X1 U1052 ( .A(n1344), .B(n1281), .ZN(n1337) );
XOR2_X1 U1053 ( .A(G116), .B(G119), .Z(n1281) );
XNOR2_X1 U1054 ( .A(KEYINPUT39), .B(KEYINPUT3), .ZN(n1344) );
XOR2_X1 U1055 ( .A(n1294), .B(n1345), .Z(n1331) );
XOR2_X1 U1056 ( .A(KEYINPUT45), .B(G122), .Z(n1345) );
INV_X1 U1057 ( .A(G110), .ZN(n1294) );
XNOR2_X1 U1058 ( .A(n1346), .B(KEYINPUT46), .ZN(n1326) );
NAND2_X1 U1059 ( .A1(G214), .A2(n1346), .ZN(n1075) );
NAND2_X1 U1060 ( .A1(n1273), .A2(n1324), .ZN(n1346) );
INV_X1 U1061 ( .A(G237), .ZN(n1324) );
NAND2_X1 U1062 ( .A1(n1347), .A2(n1255), .ZN(n1215) );
NAND3_X1 U1063 ( .A1(n1085), .A2(n1060), .A3(n1348), .ZN(n1255) );
XOR2_X1 U1064 ( .A(KEYINPUT48), .B(G952), .Z(n1348) );
NAND4_X1 U1065 ( .A1(G953), .A2(G902), .A3(n1085), .A4(n1140), .ZN(n1347) );
INV_X1 U1066 ( .A(G898), .ZN(n1140) );
NAND2_X1 U1067 ( .A1(G237), .A2(G234), .ZN(n1085) );
INV_X1 U1068 ( .A(n1251), .ZN(n1214) );
NAND2_X1 U1069 ( .A1(n1067), .A2(n1064), .ZN(n1251) );
NAND2_X1 U1070 ( .A1(G221), .A2(n1283), .ZN(n1064) );
NAND2_X1 U1071 ( .A1(G234), .A2(n1273), .ZN(n1283) );
INV_X1 U1072 ( .A(n1054), .ZN(n1067) );
XNOR2_X1 U1073 ( .A(n1101), .B(KEYINPUT26), .ZN(n1054) );
XNOR2_X1 U1074 ( .A(n1349), .B(G469), .ZN(n1101) );
NAND2_X1 U1075 ( .A1(n1350), .A2(n1273), .ZN(n1349) );
INV_X1 U1076 ( .A(G902), .ZN(n1273) );
XOR2_X1 U1077 ( .A(n1351), .B(n1352), .Z(n1350) );
XOR2_X1 U1078 ( .A(n1185), .B(n1175), .Z(n1352) );
XNOR2_X1 U1079 ( .A(n1353), .B(n1127), .ZN(n1175) );
XOR2_X1 U1080 ( .A(G131), .B(G137), .Z(n1127) );
XOR2_X1 U1081 ( .A(n1128), .B(KEYINPUT51), .Z(n1353) );
INV_X1 U1082 ( .A(G134), .ZN(n1128) );
XOR2_X1 U1083 ( .A(n1354), .B(n1355), .Z(n1185) );
XOR2_X1 U1084 ( .A(G110), .B(n1356), .Z(n1355) );
AND2_X1 U1085 ( .A1(n1060), .A2(G227), .ZN(n1356) );
INV_X1 U1086 ( .A(G953), .ZN(n1060) );
XNOR2_X1 U1087 ( .A(G140), .B(KEYINPUT14), .ZN(n1354) );
XNOR2_X1 U1088 ( .A(KEYINPUT23), .B(n1357), .ZN(n1351) );
NOR2_X1 U1089 ( .A1(KEYINPUT1), .A2(n1358), .ZN(n1357) );
XOR2_X1 U1090 ( .A(n1123), .B(n1359), .Z(n1358) );
INV_X1 U1091 ( .A(n1191), .ZN(n1359) );
XNOR2_X1 U1092 ( .A(G101), .B(n1360), .ZN(n1191) );
XOR2_X1 U1093 ( .A(G107), .B(G104), .Z(n1360) );
XNOR2_X1 U1094 ( .A(G146), .B(n1313), .ZN(n1123) );
XOR2_X1 U1095 ( .A(G128), .B(n1236), .Z(n1313) );
INV_X1 U1096 ( .A(G143), .ZN(n1236) );
endmodule


