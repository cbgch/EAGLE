//Key = 1111000000000011001110101110010101101110000110100001111101001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287;

XOR2_X1 U726 ( .A(G107), .B(n984), .Z(G9) );
NOR2_X1 U727 ( .A1(n985), .A2(n986), .ZN(G75) );
AND3_X1 U728 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
INV_X1 U729 ( .A(G952), .ZN(n989) );
NOR3_X1 U730 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n985) );
NOR2_X1 U731 ( .A1(n993), .A2(n994), .ZN(n991) );
NOR3_X1 U732 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n993) );
INV_X1 U733 ( .A(n998), .ZN(n996) );
NAND3_X1 U734 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n995) );
NAND3_X1 U735 ( .A1(n1002), .A2(n988), .A3(n987), .ZN(n990) );
NAND4_X1 U736 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n987) );
NOR4_X1 U737 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
XOR2_X1 U738 ( .A(n1011), .B(G472), .Z(n1008) );
NAND2_X1 U739 ( .A1(KEYINPUT19), .A2(n1012), .ZN(n1011) );
NOR2_X1 U740 ( .A1(n1013), .A2(n1014), .ZN(n1005) );
XOR2_X1 U741 ( .A(n1015), .B(n1016), .Z(n1014) );
NAND2_X1 U742 ( .A1(n1017), .A2(n1018), .ZN(n1004) );
NAND2_X1 U743 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NAND2_X1 U744 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
OR2_X1 U745 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
INV_X1 U746 ( .A(KEYINPUT29), .ZN(n1022) );
NAND2_X1 U747 ( .A1(n1023), .A2(G475), .ZN(n1003) );
NOR2_X1 U748 ( .A1(n1024), .A2(KEYINPUT17), .ZN(n1023) );
NAND3_X1 U749 ( .A1(n1025), .A2(n1000), .A3(n1026), .ZN(n1002) );
INV_X1 U750 ( .A(n997), .ZN(n1026) );
XNOR2_X1 U751 ( .A(n1027), .B(KEYINPUT46), .ZN(n997) );
NAND2_X1 U752 ( .A1(n1028), .A2(n1029), .ZN(n1025) );
NAND4_X1 U753 ( .A1(n998), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
NAND2_X1 U754 ( .A1(n1009), .A2(n1033), .ZN(n1032) );
NAND2_X1 U755 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
XNOR2_X1 U756 ( .A(n1036), .B(KEYINPUT55), .ZN(n1034) );
NAND4_X1 U757 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1031) );
NAND2_X1 U758 ( .A1(n1001), .A2(n994), .ZN(n1039) );
INV_X1 U759 ( .A(KEYINPUT11), .ZN(n994) );
NAND3_X1 U760 ( .A1(n1041), .A2(n1042), .A3(n1035), .ZN(n1038) );
NAND2_X1 U761 ( .A1(n1036), .A2(n1043), .ZN(n1037) );
NAND2_X1 U762 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U763 ( .A1(n1007), .A2(n1046), .ZN(n1045) );
INV_X1 U764 ( .A(n1047), .ZN(n1044) );
NAND3_X1 U765 ( .A1(n1035), .A2(n1048), .A3(n1036), .ZN(n1028) );
NAND2_X1 U766 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U767 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XNOR2_X1 U768 ( .A(n998), .B(KEYINPUT62), .ZN(n1051) );
NAND2_X1 U769 ( .A1(n999), .A2(n1053), .ZN(n1049) );
NAND2_X1 U770 ( .A1(n1054), .A2(n1055), .ZN(G72) );
NAND2_X1 U771 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U772 ( .A1(n1058), .A2(n1059), .ZN(n1054) );
INV_X1 U773 ( .A(n1056), .ZN(n1059) );
NOR2_X1 U774 ( .A1(KEYINPUT4), .A2(n1060), .ZN(n1056) );
XOR2_X1 U775 ( .A(n1061), .B(n1062), .Z(n1060) );
NOR2_X1 U776 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
XOR2_X1 U777 ( .A(KEYINPUT18), .B(n1065), .Z(n1064) );
NOR2_X1 U778 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR3_X1 U779 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NOR2_X1 U780 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U781 ( .A1(n1073), .A2(n1074), .ZN(n1069) );
NOR2_X1 U782 ( .A1(n1075), .A2(n1076), .ZN(n1068) );
NOR4_X1 U783 ( .A1(n1077), .A2(n1078), .A3(n1076), .A4(n1075), .ZN(n1066) );
INV_X1 U784 ( .A(KEYINPUT52), .ZN(n1076) );
NOR2_X1 U785 ( .A1(n1072), .A2(n1074), .ZN(n1078) );
INV_X1 U786 ( .A(n1071), .ZN(n1074) );
XOR2_X1 U787 ( .A(n1079), .B(n1073), .Z(n1072) );
XNOR2_X1 U788 ( .A(KEYINPUT9), .B(KEYINPUT21), .ZN(n1079) );
NOR2_X1 U789 ( .A1(n1071), .A2(n1073), .ZN(n1077) );
NAND2_X1 U790 ( .A1(n988), .A2(n1080), .ZN(n1061) );
NAND3_X1 U791 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
NAND2_X1 U792 ( .A1(n1084), .A2(n1057), .ZN(n1058) );
NAND2_X1 U793 ( .A1(G953), .A2(n1085), .ZN(n1057) );
INV_X1 U794 ( .A(n1063), .ZN(n1084) );
XOR2_X1 U795 ( .A(n1086), .B(n1087), .Z(G69) );
XOR2_X1 U796 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND3_X1 U797 ( .A1(n1090), .A2(n988), .A3(KEYINPUT36), .ZN(n1089) );
NAND2_X1 U798 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
NAND2_X1 U799 ( .A1(G953), .A2(n1093), .ZN(n1092) );
XOR2_X1 U800 ( .A(n1094), .B(KEYINPUT38), .Z(n1091) );
NOR3_X1 U801 ( .A1(n988), .A2(KEYINPUT12), .A3(n1095), .ZN(n1086) );
AND2_X1 U802 ( .A1(G224), .A2(G898), .ZN(n1095) );
NOR3_X1 U803 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(G66) );
NOR3_X1 U804 ( .A1(n1099), .A2(G953), .A3(G952), .ZN(n1098) );
AND2_X1 U805 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
INV_X1 U806 ( .A(KEYINPUT5), .ZN(n1099) );
XNOR2_X1 U807 ( .A(n1101), .B(n1102), .ZN(n1096) );
NOR2_X1 U808 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U809 ( .A1(n1100), .A2(n1105), .ZN(G63) );
XOR2_X1 U810 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U811 ( .A1(n1108), .A2(n1104), .ZN(n1107) );
NAND2_X1 U812 ( .A1(KEYINPUT25), .A2(n1109), .ZN(n1106) );
NOR2_X1 U813 ( .A1(n1110), .A2(n1111), .ZN(G60) );
XOR2_X1 U814 ( .A(KEYINPUT45), .B(n1100), .Z(n1111) );
XOR2_X1 U815 ( .A(n1112), .B(n1113), .Z(n1110) );
NOR2_X1 U816 ( .A1(n1018), .A2(n1104), .ZN(n1113) );
INV_X1 U817 ( .A(G475), .ZN(n1018) );
XNOR2_X1 U818 ( .A(G104), .B(n1114), .ZN(G6) );
NOR2_X1 U819 ( .A1(n1115), .A2(n1116), .ZN(G57) );
XOR2_X1 U820 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND3_X1 U821 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1117) );
NAND2_X1 U822 ( .A1(KEYINPUT30), .A2(n1122), .ZN(n1121) );
NAND3_X1 U823 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1120) );
INV_X1 U824 ( .A(KEYINPUT30), .ZN(n1124) );
OR2_X1 U825 ( .A1(n1125), .A2(n1123), .ZN(n1119) );
AND3_X1 U826 ( .A1(G472), .A2(n992), .A3(n1126), .ZN(n1123) );
XNOR2_X1 U827 ( .A(G902), .B(KEYINPUT61), .ZN(n1126) );
NOR2_X1 U828 ( .A1(KEYINPUT63), .A2(n1122), .ZN(n1125) );
XNOR2_X1 U829 ( .A(n1127), .B(n1128), .ZN(n1122) );
NOR2_X1 U830 ( .A1(n1129), .A2(n988), .ZN(n1115) );
XNOR2_X1 U831 ( .A(G952), .B(KEYINPUT20), .ZN(n1129) );
NOR2_X1 U832 ( .A1(n1100), .A2(n1130), .ZN(G54) );
XOR2_X1 U833 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U834 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U835 ( .A1(n1135), .A2(n1104), .ZN(n1134) );
NOR2_X1 U836 ( .A1(KEYINPUT59), .A2(n1136), .ZN(n1133) );
XOR2_X1 U837 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U838 ( .A(G110), .B(n1139), .Z(n1138) );
XNOR2_X1 U839 ( .A(G140), .B(KEYINPUT37), .ZN(n1137) );
NOR2_X1 U840 ( .A1(n1140), .A2(n1141), .ZN(n1131) );
XOR2_X1 U841 ( .A(KEYINPUT35), .B(n1142), .Z(n1141) );
AND2_X1 U842 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U843 ( .A1(n1100), .A2(n1145), .ZN(G51) );
XOR2_X1 U844 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U845 ( .A(n1148), .B(n1149), .ZN(n1147) );
XNOR2_X1 U846 ( .A(n1150), .B(n1151), .ZN(n1146) );
NOR2_X1 U847 ( .A1(n1016), .A2(n1104), .ZN(n1151) );
NAND2_X1 U848 ( .A1(G902), .A2(n992), .ZN(n1104) );
NAND4_X1 U849 ( .A1(n1152), .A2(n1153), .A3(n1083), .A4(n1154), .ZN(n992) );
XNOR2_X1 U850 ( .A(KEYINPUT31), .B(n1082), .ZN(n1154) );
AND4_X1 U851 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1083) );
NOR2_X1 U852 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND3_X1 U853 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1155) );
OR2_X1 U854 ( .A1(n1053), .A2(KEYINPUT32), .ZN(n1162) );
OR2_X1 U855 ( .A1(n1164), .A2(n1165), .ZN(n1053) );
NAND2_X1 U856 ( .A1(KEYINPUT32), .A2(n1165), .ZN(n1161) );
INV_X1 U857 ( .A(n1090), .ZN(n1153) );
NAND4_X1 U858 ( .A1(n1166), .A2(n1114), .A3(n1167), .A4(n1168), .ZN(n1090) );
NOR4_X1 U859 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n984), .ZN(n1168) );
AND3_X1 U860 ( .A1(n1165), .A2(n1172), .A3(n1173), .ZN(n984) );
NAND2_X1 U861 ( .A1(n1174), .A2(n1175), .ZN(n1167) );
NAND2_X1 U862 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND2_X1 U863 ( .A1(n1009), .A2(n1030), .ZN(n1177) );
XOR2_X1 U864 ( .A(KEYINPUT54), .B(n1052), .Z(n1176) );
NAND3_X1 U865 ( .A1(n1173), .A2(n1172), .A3(n1164), .ZN(n1114) );
NAND4_X1 U866 ( .A1(n1036), .A2(n1172), .A3(n1178), .A4(n1010), .ZN(n1166) );
XOR2_X1 U867 ( .A(n1081), .B(KEYINPUT28), .Z(n1152) );
NOR2_X1 U868 ( .A1(n988), .A2(G952), .ZN(n1100) );
XNOR2_X1 U869 ( .A(G146), .B(n1156), .ZN(G48) );
NAND3_X1 U870 ( .A1(n1164), .A2(n1047), .A3(n1179), .ZN(n1156) );
XNOR2_X1 U871 ( .A(G143), .B(n1158), .ZN(G45) );
NAND4_X1 U872 ( .A1(n1180), .A2(n1047), .A3(n1178), .A4(n1010), .ZN(n1158) );
XOR2_X1 U873 ( .A(G140), .B(n1160), .Z(G42) );
AND2_X1 U874 ( .A1(n1181), .A2(n1001), .ZN(n1160) );
AND2_X1 U875 ( .A1(n1035), .A2(n1173), .ZN(n1001) );
XNOR2_X1 U876 ( .A(G137), .B(n1081), .ZN(G39) );
NAND3_X1 U877 ( .A1(n998), .A2(n1035), .A3(n1179), .ZN(n1081) );
XOR2_X1 U878 ( .A(G134), .B(n1182), .Z(G36) );
AND2_X1 U879 ( .A1(n1165), .A2(n1163), .ZN(n1182) );
AND2_X1 U880 ( .A1(n1180), .A2(n1035), .ZN(n1163) );
XNOR2_X1 U881 ( .A(G131), .B(n1183), .ZN(G33) );
NAND3_X1 U882 ( .A1(n1164), .A2(n1184), .A3(n1180), .ZN(n1183) );
AND3_X1 U883 ( .A1(n1052), .A2(n1173), .A3(n1185), .ZN(n1180) );
XOR2_X1 U884 ( .A(KEYINPUT58), .B(n1035), .Z(n1184) );
AND2_X1 U885 ( .A1(n1046), .A2(n1186), .ZN(n1035) );
XOR2_X1 U886 ( .A(G128), .B(n1187), .Z(G30) );
NOR2_X1 U887 ( .A1(KEYINPUT42), .A2(n1082), .ZN(n1187) );
NAND3_X1 U888 ( .A1(n1165), .A2(n1047), .A3(n1179), .ZN(n1082) );
AND4_X1 U889 ( .A1(n1185), .A2(n1173), .A3(n1009), .A4(n1188), .ZN(n1179) );
NAND2_X1 U890 ( .A1(n1189), .A2(n1190), .ZN(G3) );
NAND4_X1 U891 ( .A1(n1174), .A2(n1052), .A3(n1191), .A4(n1192), .ZN(n1190) );
NAND2_X1 U892 ( .A1(KEYINPUT53), .A2(G101), .ZN(n1192) );
OR2_X1 U893 ( .A1(G101), .A2(KEYINPUT1), .ZN(n1191) );
NAND3_X1 U894 ( .A1(G101), .A2(n1193), .A3(KEYINPUT53), .ZN(n1189) );
NAND3_X1 U895 ( .A1(n1174), .A2(n1052), .A3(KEYINPUT1), .ZN(n1193) );
INV_X1 U896 ( .A(n1194), .ZN(n1174) );
XOR2_X1 U897 ( .A(G125), .B(n1159), .Z(G27) );
AND3_X1 U898 ( .A1(n1036), .A2(n1047), .A3(n1181), .ZN(n1159) );
AND4_X1 U899 ( .A1(n1185), .A2(n1164), .A3(n1009), .A4(n1030), .ZN(n1181) );
AND2_X1 U900 ( .A1(n1195), .A2(n1000), .ZN(n1185) );
NAND2_X1 U901 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U902 ( .A1(n1063), .A2(G902), .ZN(n1197) );
NOR2_X1 U903 ( .A1(G900), .A2(n988), .ZN(n1063) );
OR2_X1 U904 ( .A1(n1027), .A2(G953), .ZN(n1196) );
XNOR2_X1 U905 ( .A(G122), .B(n1198), .ZN(G24) );
NAND4_X1 U906 ( .A1(n1172), .A2(n1199), .A3(n1178), .A4(n1010), .ZN(n1198) );
XNOR2_X1 U907 ( .A(KEYINPUT23), .B(n1013), .ZN(n1199) );
AND2_X1 U908 ( .A1(n1200), .A2(n999), .ZN(n1172) );
NOR2_X1 U909 ( .A1(n1009), .A2(n1201), .ZN(n999) );
XOR2_X1 U910 ( .A(n1202), .B(n1171), .Z(G21) );
AND4_X1 U911 ( .A1(n1203), .A2(n998), .A3(n1009), .A4(n1188), .ZN(n1171) );
NAND2_X1 U912 ( .A1(KEYINPUT33), .A2(n1204), .ZN(n1202) );
XNOR2_X1 U913 ( .A(n1170), .B(n1205), .ZN(G18) );
XOR2_X1 U914 ( .A(KEYINPUT2), .B(G116), .Z(n1205) );
AND3_X1 U915 ( .A1(n1052), .A2(n1165), .A3(n1203), .ZN(n1170) );
NOR2_X1 U916 ( .A1(n1178), .A2(n1206), .ZN(n1165) );
XOR2_X1 U917 ( .A(G113), .B(n1169), .Z(G15) );
AND3_X1 U918 ( .A1(n1164), .A2(n1052), .A3(n1203), .ZN(n1169) );
AND2_X1 U919 ( .A1(n1036), .A2(n1200), .ZN(n1203) );
INV_X1 U920 ( .A(n1013), .ZN(n1036) );
NAND2_X1 U921 ( .A1(n1041), .A2(n1207), .ZN(n1013) );
AND2_X1 U922 ( .A1(n1040), .A2(n1188), .ZN(n1052) );
AND2_X1 U923 ( .A1(n1206), .A2(n1178), .ZN(n1164) );
INV_X1 U924 ( .A(n1010), .ZN(n1206) );
XOR2_X1 U925 ( .A(G110), .B(n1208), .Z(G12) );
NOR3_X1 U926 ( .A1(n1194), .A2(n1201), .A3(n1040), .ZN(n1208) );
INV_X1 U927 ( .A(n1009), .ZN(n1040) );
XOR2_X1 U928 ( .A(n1209), .B(n1103), .Z(n1009) );
NAND2_X1 U929 ( .A1(G217), .A2(n1210), .ZN(n1103) );
NAND2_X1 U930 ( .A1(n1101), .A2(n1211), .ZN(n1209) );
XNOR2_X1 U931 ( .A(n1212), .B(n1213), .ZN(n1101) );
XNOR2_X1 U932 ( .A(n1073), .B(n1214), .ZN(n1213) );
XOR2_X1 U933 ( .A(n1215), .B(n1216), .Z(n1212) );
NAND2_X1 U934 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
NAND4_X1 U935 ( .A1(G137), .A2(G221), .A3(G234), .A4(n988), .ZN(n1218) );
NAND2_X1 U936 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
NAND3_X1 U937 ( .A1(G234), .A2(n988), .A3(G221), .ZN(n1220) );
XOR2_X1 U938 ( .A(KEYINPUT57), .B(G137), .Z(n1219) );
INV_X1 U939 ( .A(n1030), .ZN(n1201) );
XOR2_X1 U940 ( .A(n1188), .B(KEYINPUT15), .Z(n1030) );
XNOR2_X1 U941 ( .A(n1012), .B(G472), .ZN(n1188) );
NAND2_X1 U942 ( .A1(n1221), .A2(n1211), .ZN(n1012) );
XOR2_X1 U943 ( .A(n1222), .B(n1118), .Z(n1221) );
XOR2_X1 U944 ( .A(n1223), .B(G101), .Z(n1118) );
NAND2_X1 U945 ( .A1(G210), .A2(n1224), .ZN(n1223) );
NAND2_X1 U946 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
OR2_X1 U947 ( .A1(n1128), .A2(n1144), .ZN(n1226) );
NAND2_X1 U948 ( .A1(n1227), .A2(n1144), .ZN(n1225) );
XNOR2_X1 U949 ( .A(n1128), .B(KEYINPUT22), .ZN(n1227) );
XNOR2_X1 U950 ( .A(n1228), .B(n1229), .ZN(n1128) );
XNOR2_X1 U951 ( .A(n1204), .B(G116), .ZN(n1229) );
XNOR2_X1 U952 ( .A(n1148), .B(G113), .ZN(n1228) );
NAND3_X1 U953 ( .A1(n1173), .A2(n1200), .A3(n998), .ZN(n1194) );
NOR2_X1 U954 ( .A1(n1010), .A2(n1178), .ZN(n998) );
XOR2_X1 U955 ( .A(n1024), .B(G475), .Z(n1178) );
INV_X1 U956 ( .A(n1021), .ZN(n1024) );
NAND2_X1 U957 ( .A1(n1230), .A2(n1211), .ZN(n1021) );
XOR2_X1 U958 ( .A(n1112), .B(KEYINPUT43), .Z(n1230) );
XOR2_X1 U959 ( .A(n1231), .B(n1232), .Z(n1112) );
XOR2_X1 U960 ( .A(G131), .B(n1233), .Z(n1232) );
XOR2_X1 U961 ( .A(G146), .B(G143), .Z(n1233) );
XOR2_X1 U962 ( .A(n1234), .B(n1235), .Z(n1231) );
XNOR2_X1 U963 ( .A(n1236), .B(n1073), .ZN(n1234) );
XNOR2_X1 U964 ( .A(G125), .B(G140), .ZN(n1073) );
NAND2_X1 U965 ( .A1(G214), .A2(n1224), .ZN(n1236) );
NOR2_X1 U966 ( .A1(G953), .A2(G237), .ZN(n1224) );
XNOR2_X1 U967 ( .A(n1237), .B(n1238), .ZN(n1010) );
XNOR2_X1 U968 ( .A(KEYINPUT13), .B(n1108), .ZN(n1238) );
INV_X1 U969 ( .A(G478), .ZN(n1108) );
NAND2_X1 U970 ( .A1(n1109), .A2(n1211), .ZN(n1237) );
XOR2_X1 U971 ( .A(n1239), .B(n1240), .Z(n1109) );
NOR2_X1 U972 ( .A1(KEYINPUT49), .A2(n1241), .ZN(n1240) );
XOR2_X1 U973 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U974 ( .A(n1244), .B(n1245), .ZN(n1243) );
INV_X1 U975 ( .A(n1246), .ZN(n1245) );
NOR2_X1 U976 ( .A1(KEYINPUT50), .A2(n1247), .ZN(n1244) );
NOR2_X1 U977 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XOR2_X1 U978 ( .A(n1250), .B(KEYINPUT34), .Z(n1249) );
NAND2_X1 U979 ( .A1(G134), .A2(n1251), .ZN(n1250) );
NOR2_X1 U980 ( .A1(G134), .A2(n1251), .ZN(n1248) );
XOR2_X1 U981 ( .A(G128), .B(G143), .Z(n1251) );
XNOR2_X1 U982 ( .A(G122), .B(KEYINPUT16), .ZN(n1242) );
NAND3_X1 U983 ( .A1(G234), .A2(n988), .A3(G217), .ZN(n1239) );
AND4_X1 U984 ( .A1(n1047), .A2(n1000), .A3(n1252), .A4(n1253), .ZN(n1200) );
NAND2_X1 U985 ( .A1(G953), .A2(n1254), .ZN(n1253) );
NAND2_X1 U986 ( .A1(G902), .A2(n1093), .ZN(n1254) );
INV_X1 U987 ( .A(G898), .ZN(n1093) );
NAND2_X1 U988 ( .A1(n1027), .A2(n988), .ZN(n1252) );
XNOR2_X1 U989 ( .A(G952), .B(KEYINPUT56), .ZN(n1027) );
NAND2_X1 U990 ( .A1(G237), .A2(G234), .ZN(n1000) );
NOR2_X1 U991 ( .A1(n1046), .A2(n1255), .ZN(n1047) );
XNOR2_X1 U992 ( .A(KEYINPUT0), .B(n1007), .ZN(n1255) );
INV_X1 U993 ( .A(n1186), .ZN(n1007) );
NAND2_X1 U994 ( .A1(G214), .A2(n1256), .ZN(n1186) );
XOR2_X1 U995 ( .A(n1257), .B(n1016), .Z(n1046) );
NAND2_X1 U996 ( .A1(G210), .A2(n1256), .ZN(n1016) );
NAND2_X1 U997 ( .A1(n1258), .A2(n1211), .ZN(n1256) );
XNOR2_X1 U998 ( .A(G237), .B(KEYINPUT8), .ZN(n1258) );
NAND2_X1 U999 ( .A1(KEYINPUT60), .A2(n1015), .ZN(n1257) );
NAND2_X1 U1000 ( .A1(n1259), .A2(n1211), .ZN(n1015) );
XOR2_X1 U1001 ( .A(n1149), .B(n1260), .Z(n1259) );
XNOR2_X1 U1002 ( .A(n1261), .B(n1262), .ZN(n1260) );
NOR2_X1 U1003 ( .A1(KEYINPUT47), .A2(n1148), .ZN(n1262) );
NOR2_X1 U1004 ( .A1(KEYINPUT40), .A2(n1150), .ZN(n1261) );
NAND2_X1 U1005 ( .A1(G224), .A2(n988), .ZN(n1150) );
INV_X1 U1006 ( .A(G953), .ZN(n988) );
XOR2_X1 U1007 ( .A(n1094), .B(G125), .Z(n1149) );
XOR2_X1 U1008 ( .A(n1263), .B(n1264), .Z(n1094) );
XOR2_X1 U1009 ( .A(n1235), .B(n1265), .Z(n1264) );
XOR2_X1 U1010 ( .A(G104), .B(n1266), .Z(n1235) );
XOR2_X1 U1011 ( .A(G122), .B(G113), .Z(n1266) );
XNOR2_X1 U1012 ( .A(n1246), .B(n1267), .ZN(n1263) );
XOR2_X1 U1013 ( .A(KEYINPUT44), .B(n1214), .Z(n1267) );
XNOR2_X1 U1014 ( .A(n1204), .B(G110), .ZN(n1214) );
INV_X1 U1015 ( .A(G119), .ZN(n1204) );
XOR2_X1 U1016 ( .A(G107), .B(G116), .Z(n1246) );
NOR2_X1 U1017 ( .A1(n1041), .A2(n1042), .ZN(n1173) );
INV_X1 U1018 ( .A(n1207), .ZN(n1042) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1210), .ZN(n1207) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1211), .ZN(n1210) );
XNOR2_X1 U1021 ( .A(n1268), .B(n1135), .ZN(n1041) );
INV_X1 U1022 ( .A(G469), .ZN(n1135) );
NAND2_X1 U1023 ( .A1(n1269), .A2(n1211), .ZN(n1268) );
INV_X1 U1024 ( .A(G902), .ZN(n1211) );
XOR2_X1 U1025 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U1026 ( .A(n1139), .B(n1272), .ZN(n1271) );
NAND3_X1 U1027 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1272) );
NAND2_X1 U1028 ( .A1(KEYINPUT48), .A2(n1140), .ZN(n1275) );
NOR2_X1 U1029 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
OR3_X1 U1030 ( .A1(n1127), .A2(KEYINPUT48), .A3(n1143), .ZN(n1274) );
NAND2_X1 U1031 ( .A1(n1276), .A2(n1143), .ZN(n1273) );
XNOR2_X1 U1032 ( .A(n1277), .B(n1278), .ZN(n1143) );
XOR2_X1 U1033 ( .A(G104), .B(n1279), .Z(n1278) );
XOR2_X1 U1034 ( .A(KEYINPUT26), .B(G107), .Z(n1279) );
XNOR2_X1 U1035 ( .A(n1071), .B(n1265), .ZN(n1277) );
XOR2_X1 U1036 ( .A(G101), .B(KEYINPUT39), .Z(n1265) );
XNOR2_X1 U1037 ( .A(n1280), .B(n1281), .ZN(n1071) );
XNOR2_X1 U1038 ( .A(KEYINPUT10), .B(n1282), .ZN(n1281) );
INV_X1 U1039 ( .A(n1148), .ZN(n1282) );
XOR2_X1 U1040 ( .A(G143), .B(n1216), .Z(n1148) );
XOR2_X1 U1041 ( .A(G128), .B(G146), .Z(n1216) );
XNOR2_X1 U1042 ( .A(KEYINPUT3), .B(KEYINPUT27), .ZN(n1280) );
XNOR2_X1 U1043 ( .A(KEYINPUT7), .B(n1144), .ZN(n1276) );
INV_X1 U1044 ( .A(n1127), .ZN(n1144) );
XOR2_X1 U1045 ( .A(n1075), .B(KEYINPUT24), .Z(n1127) );
XOR2_X1 U1046 ( .A(G131), .B(n1283), .Z(n1075) );
XOR2_X1 U1047 ( .A(G137), .B(G134), .Z(n1283) );
NOR2_X1 U1048 ( .A1(n1085), .A2(G953), .ZN(n1139) );
INV_X1 U1049 ( .A(G227), .ZN(n1085) );
XNOR2_X1 U1050 ( .A(KEYINPUT41), .B(n1284), .ZN(n1270) );
NOR2_X1 U1051 ( .A1(KEYINPUT6), .A2(n1285), .ZN(n1284) );
XOR2_X1 U1052 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U1053 ( .A(G140), .B(KEYINPUT14), .ZN(n1287) );
NAND2_X1 U1054 ( .A1(KEYINPUT51), .A2(G110), .ZN(n1286) );
endmodule


