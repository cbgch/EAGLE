//Key = 1010010011000000110001111110010111010011111011000010100101010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342;

XNOR2_X1 U738 ( .A(G107), .B(n1027), .ZN(G9) );
NAND4_X1 U739 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
NOR2_X1 U740 ( .A1(KEYINPUT30), .A2(n1032), .ZN(n1030) );
NOR2_X1 U741 ( .A1(n1033), .A2(n1034), .ZN(G75) );
NOR4_X1 U742 ( .A1(G953), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1034) );
NOR2_X1 U743 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U744 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NOR2_X1 U745 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NOR2_X1 U746 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U747 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR3_X1 U748 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1046) );
NOR2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U750 ( .A1(n1028), .A2(n1053), .ZN(n1051) );
NOR3_X1 U751 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1049) );
NOR2_X1 U752 ( .A1(n1057), .A2(n1058), .ZN(n1048) );
XNOR2_X1 U753 ( .A(n1059), .B(KEYINPUT14), .ZN(n1057) );
NOR3_X1 U754 ( .A1(n1052), .A2(n1060), .A3(n1055), .ZN(n1044) );
NOR2_X1 U755 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR2_X1 U756 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR4_X1 U757 ( .A1(n1065), .A2(n1055), .A3(n1052), .A4(n1047), .ZN(n1040) );
INV_X1 U758 ( .A(n1066), .ZN(n1047) );
NOR2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR3_X1 U761 ( .A1(n1035), .A2(G953), .A3(G952), .ZN(n1033) );
AND4_X1 U762 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1035) );
NOR4_X1 U763 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
XNOR2_X1 U764 ( .A(n1079), .B(n1080), .ZN(n1078) );
XNOR2_X1 U765 ( .A(G472), .B(KEYINPUT3), .ZN(n1080) );
XOR2_X1 U766 ( .A(G475), .B(n1081), .Z(n1077) );
AND2_X1 U767 ( .A1(n1063), .A2(n1054), .ZN(n1073) );
XNOR2_X1 U768 ( .A(KEYINPUT0), .B(n1082), .ZN(n1072) );
XOR2_X1 U769 ( .A(n1083), .B(n1084), .Z(n1071) );
NAND2_X1 U770 ( .A1(KEYINPUT50), .A2(n1085), .ZN(n1084) );
XOR2_X1 U771 ( .A(n1086), .B(n1087), .Z(G72) );
XOR2_X1 U772 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U773 ( .A1(n1090), .A2(G953), .ZN(n1089) );
NOR2_X1 U774 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NOR2_X1 U775 ( .A1(KEYINPUT1), .A2(n1093), .ZN(n1088) );
NOR2_X1 U776 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
AND2_X1 U777 ( .A1(G227), .A2(G900), .ZN(n1094) );
NAND2_X1 U778 ( .A1(n1096), .A2(n1097), .ZN(n1086) );
INV_X1 U779 ( .A(n1098), .ZN(n1097) );
XOR2_X1 U780 ( .A(n1099), .B(n1100), .Z(n1096) );
XNOR2_X1 U781 ( .A(n1101), .B(n1102), .ZN(n1100) );
NOR2_X1 U782 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U783 ( .A(KEYINPUT27), .B(n1105), .Z(n1104) );
NOR2_X1 U784 ( .A1(G125), .A2(n1106), .ZN(n1105) );
NOR2_X1 U785 ( .A1(G140), .A2(n1107), .ZN(n1103) );
XOR2_X1 U786 ( .A(n1108), .B(KEYINPUT40), .Z(n1099) );
NAND2_X1 U787 ( .A1(n1109), .A2(KEYINPUT5), .ZN(n1108) );
XNOR2_X1 U788 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U789 ( .A1(KEYINPUT15), .A2(n1112), .ZN(n1111) );
XOR2_X1 U790 ( .A(n1113), .B(n1114), .Z(G69) );
NOR2_X1 U791 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U792 ( .A(n1117), .B(KEYINPUT23), .Z(n1116) );
NAND3_X1 U793 ( .A1(n1118), .A2(n1095), .A3(n1119), .ZN(n1117) );
NAND2_X1 U794 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
INV_X1 U795 ( .A(n1122), .ZN(n1121) );
XNOR2_X1 U796 ( .A(n1123), .B(n1124), .ZN(n1120) );
NOR3_X1 U797 ( .A1(n1125), .A2(n1122), .A3(n1118), .ZN(n1115) );
XNOR2_X1 U798 ( .A(n1126), .B(n1123), .ZN(n1125) );
INV_X1 U799 ( .A(n1124), .ZN(n1126) );
NAND3_X1 U800 ( .A1(G953), .A2(n1127), .A3(KEYINPUT55), .ZN(n1113) );
NAND2_X1 U801 ( .A1(G898), .A2(G224), .ZN(n1127) );
NOR3_X1 U802 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(G66) );
AND2_X1 U803 ( .A1(KEYINPUT29), .A2(n1131), .ZN(n1130) );
NOR3_X1 U804 ( .A1(KEYINPUT29), .A2(n1095), .A3(n1132), .ZN(n1129) );
INV_X1 U805 ( .A(G952), .ZN(n1132) );
XOR2_X1 U806 ( .A(n1133), .B(n1134), .Z(n1128) );
NAND2_X1 U807 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR2_X1 U808 ( .A1(n1131), .A2(n1137), .ZN(G63) );
XOR2_X1 U809 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U810 ( .A1(n1135), .A2(G478), .ZN(n1138) );
NOR2_X1 U811 ( .A1(n1131), .A2(n1140), .ZN(G60) );
NOR3_X1 U812 ( .A1(n1081), .A2(n1141), .A3(n1142), .ZN(n1140) );
AND3_X1 U813 ( .A1(n1143), .A2(G475), .A3(n1135), .ZN(n1142) );
NOR2_X1 U814 ( .A1(n1144), .A2(n1143), .ZN(n1141) );
AND2_X1 U815 ( .A1(n1037), .A2(G475), .ZN(n1144) );
XOR2_X1 U816 ( .A(G104), .B(n1145), .Z(G6) );
NOR2_X1 U817 ( .A1(n1131), .A2(n1146), .ZN(G57) );
XOR2_X1 U818 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U819 ( .A(n1149), .B(n1150), .ZN(n1148) );
XNOR2_X1 U820 ( .A(n1151), .B(n1152), .ZN(n1147) );
NOR2_X1 U821 ( .A1(KEYINPUT12), .A2(n1153), .ZN(n1152) );
NOR3_X1 U822 ( .A1(n1154), .A2(KEYINPUT36), .A3(n1155), .ZN(n1151) );
NOR2_X1 U823 ( .A1(n1131), .A2(n1156), .ZN(G54) );
XOR2_X1 U824 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U825 ( .A1(n1135), .A2(G469), .ZN(n1158) );
NAND2_X1 U826 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U827 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U828 ( .A(KEYINPUT19), .B(n1163), .Z(n1161) );
XOR2_X1 U829 ( .A(n1164), .B(KEYINPUT48), .Z(n1159) );
OR2_X1 U830 ( .A1(n1162), .A2(n1163), .ZN(n1164) );
XNOR2_X1 U831 ( .A(n1165), .B(n1166), .ZN(n1162) );
NOR2_X1 U832 ( .A1(n1167), .A2(n1168), .ZN(G51) );
XOR2_X1 U833 ( .A(KEYINPUT20), .B(n1131), .Z(n1168) );
NOR2_X1 U834 ( .A1(n1095), .A2(G952), .ZN(n1131) );
XOR2_X1 U835 ( .A(n1169), .B(n1170), .Z(n1167) );
XNOR2_X1 U836 ( .A(n1171), .B(n1172), .ZN(n1170) );
XNOR2_X1 U837 ( .A(n1173), .B(n1174), .ZN(n1172) );
NOR2_X1 U838 ( .A1(G125), .A2(KEYINPUT7), .ZN(n1174) );
XOR2_X1 U839 ( .A(n1175), .B(n1176), .Z(n1169) );
XOR2_X1 U840 ( .A(n1177), .B(KEYINPUT33), .Z(n1176) );
NAND2_X1 U841 ( .A1(n1135), .A2(n1178), .ZN(n1175) );
INV_X1 U842 ( .A(n1154), .ZN(n1135) );
NAND2_X1 U843 ( .A1(G902), .A2(n1037), .ZN(n1154) );
OR3_X1 U844 ( .A1(n1092), .A2(n1179), .A3(n1118), .ZN(n1037) );
NAND4_X1 U845 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1118) );
AND4_X1 U846 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
NAND2_X1 U847 ( .A1(KEYINPUT25), .A2(n1145), .ZN(n1182) );
AND4_X1 U848 ( .A1(n1053), .A2(n1029), .A3(n1031), .A4(n1188), .ZN(n1145) );
NAND3_X1 U849 ( .A1(n1189), .A2(n1190), .A3(KEYINPUT24), .ZN(n1181) );
NAND2_X1 U850 ( .A1(n1191), .A2(n1188), .ZN(n1180) );
NAND2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
OR4_X1 U852 ( .A1(n1194), .A2(n1052), .A3(n1062), .A4(KEYINPUT24), .ZN(n1193) );
NAND3_X1 U853 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1192) );
NAND2_X1 U854 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
OR3_X1 U855 ( .A1(n1043), .A2(KEYINPUT25), .A3(n1200), .ZN(n1198) );
INV_X1 U856 ( .A(n1029), .ZN(n1043) );
NAND3_X1 U857 ( .A1(n1201), .A2(n1202), .A3(n1062), .ZN(n1195) );
NAND2_X1 U858 ( .A1(n1028), .A2(n1029), .ZN(n1202) );
NAND2_X1 U859 ( .A1(n1068), .A2(n1059), .ZN(n1201) );
XOR2_X1 U860 ( .A(KEYINPUT10), .B(n1091), .Z(n1179) );
NAND4_X1 U861 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1091) );
NAND4_X1 U862 ( .A1(n1207), .A2(n1066), .A3(n1189), .A4(n1197), .ZN(n1203) );
XOR2_X1 U863 ( .A(n1208), .B(KEYINPUT28), .Z(n1207) );
NAND4_X1 U864 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1092) );
NAND2_X1 U865 ( .A1(n1213), .A2(n1214), .ZN(n1209) );
XNOR2_X1 U866 ( .A(n1053), .B(KEYINPUT41), .ZN(n1213) );
XNOR2_X1 U867 ( .A(n1215), .B(n1216), .ZN(G48) );
NOR2_X1 U868 ( .A1(n1200), .A2(n1217), .ZN(n1216) );
XNOR2_X1 U869 ( .A(G143), .B(n1210), .ZN(G45) );
NAND3_X1 U870 ( .A1(n1068), .A2(n1031), .A3(n1218), .ZN(n1210) );
AND3_X1 U871 ( .A1(n1076), .A2(n1219), .A3(n1208), .ZN(n1218) );
XNOR2_X1 U872 ( .A(n1220), .B(n1211), .ZN(G42) );
NAND2_X1 U873 ( .A1(n1221), .A2(n1222), .ZN(n1211) );
NAND2_X1 U874 ( .A1(KEYINPUT52), .A2(n1106), .ZN(n1220) );
XNOR2_X1 U875 ( .A(G137), .B(n1212), .ZN(G39) );
NAND3_X1 U876 ( .A1(n1223), .A2(n1070), .A3(n1222), .ZN(n1212) );
NAND2_X1 U877 ( .A1(n1224), .A2(n1225), .ZN(G36) );
NAND2_X1 U878 ( .A1(KEYINPUT63), .A2(G134), .ZN(n1225) );
XOR2_X1 U879 ( .A(n1226), .B(n1227), .Z(n1224) );
NOR2_X1 U880 ( .A1(n1194), .A2(n1228), .ZN(n1227) );
NOR2_X1 U881 ( .A1(G134), .A2(KEYINPUT63), .ZN(n1226) );
XNOR2_X1 U882 ( .A(G131), .B(n1204), .ZN(G33) );
NAND3_X1 U883 ( .A1(n1068), .A2(n1053), .A3(n1222), .ZN(n1204) );
INV_X1 U884 ( .A(n1228), .ZN(n1222) );
NAND3_X1 U885 ( .A1(n1197), .A2(n1208), .A3(n1066), .ZN(n1228) );
NOR2_X1 U886 ( .A1(n1064), .A2(n1229), .ZN(n1066) );
XOR2_X1 U887 ( .A(n1230), .B(KEYINPUT4), .Z(n1064) );
XNOR2_X1 U888 ( .A(n1231), .B(n1206), .ZN(G30) );
NAND2_X1 U889 ( .A1(n1214), .A2(n1028), .ZN(n1206) );
INV_X1 U890 ( .A(n1217), .ZN(n1214) );
NAND4_X1 U891 ( .A1(n1031), .A2(n1070), .A3(n1075), .A4(n1208), .ZN(n1217) );
XNOR2_X1 U892 ( .A(G128), .B(KEYINPUT59), .ZN(n1231) );
XNOR2_X1 U893 ( .A(G101), .B(n1232), .ZN(G3) );
NAND4_X1 U894 ( .A1(n1233), .A2(n1068), .A3(n1234), .A4(n1059), .ZN(n1232) );
NOR2_X1 U895 ( .A1(n1032), .A2(n1199), .ZN(n1234) );
XNOR2_X1 U896 ( .A(n1197), .B(KEYINPUT44), .ZN(n1233) );
INV_X1 U897 ( .A(n1058), .ZN(n1197) );
XNOR2_X1 U898 ( .A(G125), .B(n1205), .ZN(G27) );
NAND4_X1 U899 ( .A1(n1221), .A2(n1235), .A3(n1062), .A4(n1208), .ZN(n1205) );
NAND2_X1 U900 ( .A1(n1039), .A2(n1236), .ZN(n1208) );
NAND3_X1 U901 ( .A1(G902), .A2(n1237), .A3(n1098), .ZN(n1236) );
NOR2_X1 U902 ( .A1(n1238), .A2(G900), .ZN(n1098) );
NOR3_X1 U903 ( .A1(n1070), .A2(n1069), .A3(n1200), .ZN(n1221) );
XNOR2_X1 U904 ( .A(G122), .B(n1187), .ZN(G24) );
NAND4_X1 U905 ( .A1(n1190), .A2(n1029), .A3(n1076), .A4(n1219), .ZN(n1187) );
NOR2_X1 U906 ( .A1(n1075), .A2(n1070), .ZN(n1029) );
XNOR2_X1 U907 ( .A(G119), .B(n1239), .ZN(G21) );
NOR2_X1 U908 ( .A1(n1240), .A2(KEYINPUT13), .ZN(n1239) );
INV_X1 U909 ( .A(n1186), .ZN(n1240) );
NAND3_X1 U910 ( .A1(n1223), .A2(n1070), .A3(n1190), .ZN(n1186) );
XNOR2_X1 U911 ( .A(n1241), .B(n1242), .ZN(G18) );
AND2_X1 U912 ( .A1(n1190), .A2(n1189), .ZN(n1242) );
INV_X1 U913 ( .A(n1194), .ZN(n1189) );
NAND2_X1 U914 ( .A1(n1068), .A2(n1028), .ZN(n1194) );
NOR2_X1 U915 ( .A1(n1219), .A2(n1243), .ZN(n1028) );
XNOR2_X1 U916 ( .A(G113), .B(n1185), .ZN(G15) );
NAND3_X1 U917 ( .A1(n1190), .A2(n1053), .A3(n1068), .ZN(n1185) );
NOR2_X1 U918 ( .A1(n1075), .A2(n1244), .ZN(n1068) );
INV_X1 U919 ( .A(n1200), .ZN(n1053) );
NAND2_X1 U920 ( .A1(n1243), .A2(n1219), .ZN(n1200) );
INV_X1 U921 ( .A(n1076), .ZN(n1243) );
NOR3_X1 U922 ( .A1(n1199), .A2(n1032), .A3(n1052), .ZN(n1190) );
INV_X1 U923 ( .A(n1235), .ZN(n1052) );
NOR2_X1 U924 ( .A1(n1056), .A2(n1245), .ZN(n1235) );
INV_X1 U925 ( .A(n1054), .ZN(n1245) );
INV_X1 U926 ( .A(n1188), .ZN(n1032) );
XOR2_X1 U927 ( .A(n1184), .B(n1246), .Z(G12) );
XNOR2_X1 U928 ( .A(G110), .B(KEYINPUT51), .ZN(n1246) );
NAND4_X1 U929 ( .A1(n1223), .A2(n1031), .A3(n1244), .A4(n1188), .ZN(n1184) );
NAND2_X1 U930 ( .A1(n1039), .A2(n1247), .ZN(n1188) );
NAND3_X1 U931 ( .A1(n1122), .A2(n1237), .A3(G902), .ZN(n1247) );
NOR2_X1 U932 ( .A1(n1238), .A2(G898), .ZN(n1122) );
XNOR2_X1 U933 ( .A(n1095), .B(KEYINPUT22), .ZN(n1238) );
NAND3_X1 U934 ( .A1(n1237), .A2(n1095), .A3(G952), .ZN(n1039) );
NAND2_X1 U935 ( .A1(G237), .A2(G234), .ZN(n1237) );
INV_X1 U936 ( .A(n1070), .ZN(n1244) );
XOR2_X1 U937 ( .A(n1248), .B(n1155), .Z(n1070) );
INV_X1 U938 ( .A(G472), .ZN(n1155) );
NAND2_X1 U939 ( .A1(KEYINPUT38), .A2(n1079), .ZN(n1248) );
AND2_X1 U940 ( .A1(n1249), .A2(n1250), .ZN(n1079) );
XOR2_X1 U941 ( .A(n1251), .B(n1153), .Z(n1249) );
AND2_X1 U942 ( .A1(n1252), .A2(n1253), .ZN(n1153) );
NAND2_X1 U943 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U944 ( .A(G101), .ZN(n1255) );
NAND2_X1 U945 ( .A1(G210), .A2(n1256), .ZN(n1254) );
NAND3_X1 U946 ( .A1(G210), .A2(n1256), .A3(G101), .ZN(n1252) );
XNOR2_X1 U947 ( .A(n1150), .B(n1257), .ZN(n1251) );
NOR2_X1 U948 ( .A1(KEYINPUT37), .A2(n1149), .ZN(n1257) );
XOR2_X1 U949 ( .A(n1258), .B(n1259), .Z(n1149) );
INV_X1 U950 ( .A(n1260), .ZN(n1259) );
NAND2_X1 U951 ( .A1(KEYINPUT31), .A2(n1241), .ZN(n1258) );
XNOR2_X1 U952 ( .A(n1166), .B(n1261), .ZN(n1150) );
NOR2_X1 U953 ( .A1(n1199), .A2(n1058), .ZN(n1031) );
NAND2_X1 U954 ( .A1(n1056), .A2(n1054), .ZN(n1058) );
NAND2_X1 U955 ( .A1(n1262), .A2(n1263), .ZN(n1054) );
XOR2_X1 U956 ( .A(KEYINPUT62), .B(G221), .Z(n1262) );
XOR2_X1 U957 ( .A(n1083), .B(n1085), .Z(n1056) );
INV_X1 U958 ( .A(G469), .ZN(n1085) );
NAND2_X1 U959 ( .A1(n1264), .A2(n1250), .ZN(n1083) );
XOR2_X1 U960 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U961 ( .A(n1267), .B(KEYINPUT8), .ZN(n1266) );
NAND2_X1 U962 ( .A1(KEYINPUT2), .A2(n1165), .ZN(n1267) );
XNOR2_X1 U963 ( .A(n1268), .B(n1269), .ZN(n1165) );
INV_X1 U964 ( .A(n1101), .ZN(n1269) );
XNOR2_X1 U965 ( .A(n1270), .B(n1271), .ZN(n1101) );
XNOR2_X1 U966 ( .A(KEYINPUT21), .B(n1272), .ZN(n1271) );
NAND2_X1 U967 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
XOR2_X1 U968 ( .A(KEYINPUT17), .B(n1275), .Z(n1273) );
XNOR2_X1 U969 ( .A(n1276), .B(G107), .ZN(n1268) );
XNOR2_X1 U970 ( .A(n1166), .B(n1163), .ZN(n1265) );
XNOR2_X1 U971 ( .A(n1277), .B(n1278), .ZN(n1163) );
XNOR2_X1 U972 ( .A(n1106), .B(G110), .ZN(n1278) );
NAND2_X1 U973 ( .A1(G227), .A2(n1095), .ZN(n1277) );
XOR2_X1 U974 ( .A(n1279), .B(n1280), .Z(n1166) );
INV_X1 U975 ( .A(n1110), .ZN(n1280) );
XOR2_X1 U976 ( .A(G137), .B(G134), .Z(n1110) );
NAND2_X1 U977 ( .A1(KEYINPUT45), .A2(n1112), .ZN(n1279) );
INV_X1 U978 ( .A(G131), .ZN(n1112) );
INV_X1 U979 ( .A(n1062), .ZN(n1199) );
NOR2_X1 U980 ( .A1(n1229), .A2(n1082), .ZN(n1062) );
INV_X1 U981 ( .A(n1230), .ZN(n1082) );
XNOR2_X1 U982 ( .A(n1281), .B(n1178), .ZN(n1230) );
AND2_X1 U983 ( .A1(G210), .A2(n1282), .ZN(n1178) );
NAND2_X1 U984 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
XNOR2_X1 U985 ( .A(n1285), .B(n1286), .ZN(n1284) );
INV_X1 U986 ( .A(n1173), .ZN(n1286) );
XOR2_X1 U987 ( .A(n1287), .B(n1124), .Z(n1173) );
XOR2_X1 U988 ( .A(G110), .B(n1288), .Z(n1124) );
NAND2_X1 U989 ( .A1(KEYINPUT57), .A2(n1123), .ZN(n1287) );
XOR2_X1 U990 ( .A(n1289), .B(n1290), .Z(n1123) );
XNOR2_X1 U991 ( .A(n1241), .B(n1291), .ZN(n1290) );
NOR2_X1 U992 ( .A1(KEYINPUT53), .A2(n1292), .ZN(n1291) );
INV_X1 U993 ( .A(G107), .ZN(n1292) );
INV_X1 U994 ( .A(G116), .ZN(n1241) );
XNOR2_X1 U995 ( .A(n1260), .B(n1276), .ZN(n1289) );
XOR2_X1 U996 ( .A(G101), .B(n1293), .Z(n1276) );
XOR2_X1 U997 ( .A(G119), .B(n1294), .Z(n1260) );
NAND2_X1 U998 ( .A1(KEYINPUT35), .A2(n1295), .ZN(n1285) );
XNOR2_X1 U999 ( .A(n1261), .B(n1296), .ZN(n1295) );
XNOR2_X1 U1000 ( .A(G125), .B(n1177), .ZN(n1296) );
NAND2_X1 U1001 ( .A1(G224), .A2(n1095), .ZN(n1177) );
INV_X1 U1002 ( .A(n1171), .ZN(n1261) );
XOR2_X1 U1003 ( .A(n1297), .B(n1272), .Z(n1171) );
NAND2_X1 U1004 ( .A1(KEYINPUT39), .A2(n1298), .ZN(n1297) );
NAND2_X1 U1005 ( .A1(n1299), .A2(n1274), .ZN(n1298) );
NAND2_X1 U1006 ( .A1(G146), .A2(n1300), .ZN(n1274) );
XOR2_X1 U1007 ( .A(KEYINPUT32), .B(n1275), .Z(n1299) );
NOR2_X1 U1008 ( .A1(n1300), .A2(G146), .ZN(n1275) );
XNOR2_X1 U1009 ( .A(G902), .B(KEYINPUT18), .ZN(n1283) );
XOR2_X1 U1010 ( .A(n1063), .B(KEYINPUT26), .Z(n1229) );
NAND2_X1 U1011 ( .A1(G214), .A2(n1282), .ZN(n1063) );
NAND2_X1 U1012 ( .A1(n1301), .A2(n1250), .ZN(n1282) );
INV_X1 U1013 ( .A(G237), .ZN(n1301) );
NOR2_X1 U1014 ( .A1(n1055), .A2(n1069), .ZN(n1223) );
INV_X1 U1015 ( .A(n1075), .ZN(n1069) );
XNOR2_X1 U1016 ( .A(n1302), .B(n1136), .ZN(n1075) );
AND2_X1 U1017 ( .A1(G217), .A2(n1263), .ZN(n1136) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1250), .ZN(n1263) );
NAND2_X1 U1019 ( .A1(n1134), .A2(n1250), .ZN(n1302) );
XOR2_X1 U1020 ( .A(n1303), .B(n1304), .Z(n1134) );
XNOR2_X1 U1021 ( .A(n1305), .B(n1306), .ZN(n1304) );
NOR2_X1 U1022 ( .A1(KEYINPUT54), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U1023 ( .A(G110), .B(n1308), .ZN(n1307) );
XNOR2_X1 U1024 ( .A(n1272), .B(G119), .ZN(n1308) );
INV_X1 U1025 ( .A(G128), .ZN(n1272) );
NAND2_X1 U1026 ( .A1(KEYINPUT9), .A2(n1309), .ZN(n1305) );
XNOR2_X1 U1027 ( .A(G137), .B(n1310), .ZN(n1309) );
NAND3_X1 U1028 ( .A1(n1311), .A2(n1095), .A3(G221), .ZN(n1310) );
NAND2_X1 U1029 ( .A1(n1312), .A2(n1313), .ZN(n1303) );
NAND2_X1 U1030 ( .A1(n1314), .A2(n1215), .ZN(n1313) );
XOR2_X1 U1031 ( .A(KEYINPUT46), .B(n1315), .Z(n1314) );
NAND2_X1 U1032 ( .A1(n1316), .A2(G146), .ZN(n1312) );
XOR2_X1 U1033 ( .A(KEYINPUT16), .B(n1315), .Z(n1316) );
XNOR2_X1 U1034 ( .A(n1317), .B(KEYINPUT60), .ZN(n1315) );
INV_X1 U1035 ( .A(n1059), .ZN(n1055) );
NOR2_X1 U1036 ( .A1(n1076), .A2(n1219), .ZN(n1059) );
NAND2_X1 U1037 ( .A1(n1318), .A2(n1319), .ZN(n1219) );
OR2_X1 U1038 ( .A1(n1320), .A2(G475), .ZN(n1319) );
XOR2_X1 U1039 ( .A(n1321), .B(KEYINPUT58), .Z(n1318) );
NAND2_X1 U1040 ( .A1(G475), .A2(n1320), .ZN(n1321) );
XOR2_X1 U1041 ( .A(n1081), .B(KEYINPUT42), .Z(n1320) );
NOR2_X1 U1042 ( .A1(n1143), .A2(G902), .ZN(n1081) );
XOR2_X1 U1043 ( .A(n1322), .B(n1323), .Z(n1143) );
XOR2_X1 U1044 ( .A(n1324), .B(n1325), .Z(n1323) );
XNOR2_X1 U1045 ( .A(n1326), .B(n1327), .ZN(n1325) );
NOR2_X1 U1046 ( .A1(KEYINPUT6), .A2(n1328), .ZN(n1327) );
XNOR2_X1 U1047 ( .A(G122), .B(n1294), .ZN(n1328) );
XOR2_X1 U1048 ( .A(G113), .B(KEYINPUT47), .Z(n1294) );
NAND2_X1 U1049 ( .A1(KEYINPUT61), .A2(G143), .ZN(n1326) );
XNOR2_X1 U1050 ( .A(n1215), .B(G131), .ZN(n1324) );
INV_X1 U1051 ( .A(G146), .ZN(n1215) );
XNOR2_X1 U1052 ( .A(n1329), .B(n1317), .ZN(n1322) );
XNOR2_X1 U1053 ( .A(n1106), .B(n1107), .ZN(n1317) );
INV_X1 U1054 ( .A(G125), .ZN(n1107) );
INV_X1 U1055 ( .A(G140), .ZN(n1106) );
XOR2_X1 U1056 ( .A(n1330), .B(n1293), .Z(n1329) );
XOR2_X1 U1057 ( .A(G104), .B(KEYINPUT49), .Z(n1293) );
NAND2_X1 U1058 ( .A1(G214), .A2(n1256), .ZN(n1330) );
NOR2_X1 U1059 ( .A1(G953), .A2(G237), .ZN(n1256) );
XNOR2_X1 U1060 ( .A(n1331), .B(G478), .ZN(n1076) );
NAND2_X1 U1061 ( .A1(n1139), .A2(n1250), .ZN(n1331) );
INV_X1 U1062 ( .A(G902), .ZN(n1250) );
XNOR2_X1 U1063 ( .A(n1332), .B(n1333), .ZN(n1139) );
NOR2_X1 U1064 ( .A1(KEYINPUT34), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1065 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1066 ( .A(n1288), .B(G116), .ZN(n1336) );
INV_X1 U1067 ( .A(G122), .ZN(n1288) );
XNOR2_X1 U1068 ( .A(G107), .B(n1337), .ZN(n1335) );
NOR2_X1 U1069 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
XOR2_X1 U1070 ( .A(KEYINPUT43), .B(n1340), .Z(n1339) );
NOR2_X1 U1071 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
AND2_X1 U1072 ( .A1(n1342), .A2(n1341), .ZN(n1338) );
XOR2_X1 U1073 ( .A(G134), .B(KEYINPUT56), .Z(n1341) );
XNOR2_X1 U1074 ( .A(G128), .B(n1300), .ZN(n1342) );
INV_X1 U1075 ( .A(G143), .ZN(n1300) );
NAND3_X1 U1076 ( .A1(n1311), .A2(n1095), .A3(G217), .ZN(n1332) );
INV_X1 U1077 ( .A(G953), .ZN(n1095) );
XOR2_X1 U1078 ( .A(G234), .B(KEYINPUT11), .Z(n1311) );
endmodule


