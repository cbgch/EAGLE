//Key = 0000100111010010110111100110111000100010110011111101000010100100


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
n2251, n2252;

OR2_X1 U1263 ( .A1(n2252), .A2(n1692), .ZN(U280) );
OR2_X1 U1264 ( .A1(n1843), .A2(STATO_REG_0__SCAN_IN), .ZN(n1691) );
INV_X2 U1265 ( .A(n1691), .ZN(n1692) );
INV_X2 U1266 ( .A(U280), .ZN(n1693) );
NOR4_X2 U1267 ( .A1(n1842), .A2(n2163), .A3(n2168), .A4(AVERAGE), .ZN(n1947));
XOR2_X1 U1268 ( .A(n1694), .B(KEYINPUT19), .Z(U375) );
NAND2_X1 U1269 ( .A1(n1695), .A2(n1696), .ZN(U344) );
NAND2_X1 U1270 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1697), .ZN(n1696) );
NAND2_X1 U1271 ( .A1(n1698), .A2(DATA_IN_7_), .ZN(n1695) );
NAND2_X1 U1272 ( .A1(n1699), .A2(n1700), .ZN(U343) );
NAND2_X1 U1273 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1697), .ZN(n1700) );
NAND2_X1 U1274 ( .A1(n1698), .A2(DATA_IN_6_), .ZN(n1699) );
NAND2_X1 U1275 ( .A1(n1701), .A2(n1702), .ZN(U342) );
NAND2_X1 U1276 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1697), .ZN(n1702) );
NAND2_X1 U1277 ( .A1(n1698), .A2(DATA_IN_5_), .ZN(n1701) );
NAND2_X1 U1278 ( .A1(n1703), .A2(n1704), .ZN(U341) );
NAND2_X1 U1279 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1697), .ZN(n1704) );
NAND2_X1 U1280 ( .A1(n1698), .A2(n1705), .ZN(n1703) );
XOR2_X1 U1281 ( .A(n1706), .B(KEYINPUT4), .Z(n1705) );
NAND2_X1 U1282 ( .A1(n1707), .A2(n1708), .ZN(U340) );
NAND2_X1 U1283 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1697), .ZN(n1708) );
NAND2_X1 U1284 ( .A1(n1698), .A2(DATA_IN_3_), .ZN(n1707) );
NAND2_X1 U1285 ( .A1(n1709), .A2(n1710), .ZN(U339) );
NAND2_X1 U1286 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1697), .ZN(n1710) );
NAND2_X1 U1287 ( .A1(n1698), .A2(DATA_IN_2_), .ZN(n1709) );
NAND2_X1 U1288 ( .A1(n1711), .A2(n1712), .ZN(U338) );
NAND2_X1 U1289 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1697), .ZN(n1712) );
NAND2_X1 U1290 ( .A1(n1698), .A2(DATA_IN_1_), .ZN(n1711) );
NAND2_X1 U1291 ( .A1(n1713), .A2(n1714), .ZN(U337) );
NAND2_X1 U1292 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1697), .ZN(n1714) );
NAND2_X1 U1293 ( .A1(n1698), .A2(DATA_IN_0_), .ZN(n1713) );
INV_X1 U1294 ( .A(n1697), .ZN(n1698) );
NAND2_X1 U1295 ( .A1(n1694), .A2(n1715), .ZN(n1697) );
NAND3_X1 U1296 ( .A1(n1716), .A2(n1717), .A3(n1718), .ZN(n1715) );
NAND2_X1 U1297 ( .A1(n1719), .A2(n1720), .ZN(U336) );
NAND2_X1 U1298 ( .A1(n1721), .A2(DATA_IN_7_), .ZN(n1720) );
NAND2_X1 U1299 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1722), .ZN(n1719) );
NAND2_X1 U1300 ( .A1(n1723), .A2(n1724), .ZN(U335) );
NAND2_X1 U1301 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1725), .ZN(n1724) );
XNOR2_X1 U1302 ( .A(KEYINPUT47), .B(n1722), .ZN(n1725) );
NAND2_X1 U1303 ( .A1(n1721), .A2(DATA_IN_6_), .ZN(n1723) );
NAND2_X1 U1304 ( .A1(n1726), .A2(n1727), .ZN(U334) );
NAND2_X1 U1305 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1722), .ZN(n1727) );
XOR2_X1 U1306 ( .A(n1728), .B(KEYINPUT52), .Z(n1726) );
NAND2_X1 U1307 ( .A1(n1721), .A2(DATA_IN_5_), .ZN(n1728) );
NAND2_X1 U1308 ( .A1(n1729), .A2(n1730), .ZN(U333) );
NAND2_X1 U1309 ( .A1(n1731), .A2(DATA_IN_4_), .ZN(n1730) );
XOR2_X1 U1310 ( .A(n1732), .B(KEYINPUT26), .Z(n1731) );
NAND2_X1 U1311 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1722), .ZN(n1729) );
NAND2_X1 U1312 ( .A1(n1733), .A2(n1734), .ZN(U332) );
NAND2_X1 U1313 ( .A1(n1721), .A2(DATA_IN_3_), .ZN(n1734) );
NAND2_X1 U1314 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1722), .ZN(n1733) );
NAND2_X1 U1315 ( .A1(n1735), .A2(n1736), .ZN(U331) );
NAND2_X1 U1316 ( .A1(n1721), .A2(DATA_IN_2_), .ZN(n1736) );
NAND2_X1 U1317 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1722), .ZN(n1735) );
NAND2_X1 U1318 ( .A1(n1737), .A2(n1738), .ZN(U330) );
NAND2_X1 U1319 ( .A1(n1721), .A2(n1739), .ZN(n1738) );
XOR2_X1 U1320 ( .A(KEYINPUT13), .B(DATA_IN_1_), .Z(n1739) );
NAND2_X1 U1321 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1722), .ZN(n1737) );
NAND2_X1 U1322 ( .A1(n1740), .A2(n1741), .ZN(U329) );
NAND2_X1 U1323 ( .A1(DATA_IN_0_), .A2(n1742), .ZN(n1741) );
XOR2_X1 U1324 ( .A(KEYINPUT37), .B(n1721), .Z(n1742) );
INV_X1 U1325 ( .A(n1732), .ZN(n1721) );
NAND2_X1 U1326 ( .A1(n1743), .A2(n1744), .ZN(n1732) );
NAND2_X1 U1327 ( .A1(n1745), .A2(n1717), .ZN(n1744) );
NAND2_X1 U1328 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1722), .ZN(n1740) );
NAND2_X1 U1329 ( .A1(n1743), .A2(n1746), .ZN(n1722) );
NAND2_X1 U1330 ( .A1(n1747), .A2(n1717), .ZN(n1746) );
XNOR2_X1 U1331 ( .A(n1745), .B(KEYINPUT7), .ZN(n1747) );
AND2_X1 U1332 ( .A1(n1748), .A2(n1749), .ZN(n1745) );
NAND3_X1 U1333 ( .A1(n1750), .A2(n1751), .A3(n1752), .ZN(n1749) );
NAND2_X1 U1334 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1753), .ZN(n1752) );
NAND3_X1 U1335 ( .A1(n1754), .A2(n1755), .A3(n1756), .ZN(n1751) );
NAND2_X1 U1336 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1757), .ZN(n1756) );
NAND3_X1 U1337 ( .A1(n1758), .A2(n1759), .A3(n1760), .ZN(n1755) );
NAND2_X1 U1338 ( .A1(DATA_IN_5_), .A2(n1761), .ZN(n1760) );
NAND3_X1 U1339 ( .A1(n1762), .A2(n1763), .A3(n1764), .ZN(n1759) );
NAND2_X1 U1340 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1706), .ZN(n1764) );
NAND3_X1 U1341 ( .A1(n1765), .A2(n1766), .A3(n1767), .ZN(n1763) );
NAND2_X1 U1342 ( .A1(DATA_IN_3_), .A2(n1768), .ZN(n1767) );
NAND3_X1 U1343 ( .A1(n1769), .A2(n1770), .A3(n1771), .ZN(n1766) );
NAND2_X1 U1344 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1772), .ZN(n1771) );
XOR2_X1 U1345 ( .A(KEYINPUT38), .B(DATA_IN_2_), .Z(n1772) );
NAND3_X1 U1346 ( .A1(n1773), .A2(n1774), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1770) );
NAND2_X1 U1347 ( .A1(DATA_IN_1_), .A2(n1775), .ZN(n1773) );
NAND2_X1 U1348 ( .A1(n1776), .A2(n1777), .ZN(n1769) );
INV_X1 U1349 ( .A(DATA_IN_1_), .ZN(n1777) );
XOR2_X1 U1350 ( .A(RMIN_REG_1__SCAN_IN), .B(KEYINPUT39), .Z(n1776) );
NAND2_X1 U1351 ( .A1(DATA_IN_2_), .A2(n1778), .ZN(n1765) );
NAND2_X1 U1352 ( .A1(n1779), .A2(RMIN_REG_3__SCAN_IN), .ZN(n1762) );
XNOR2_X1 U1353 ( .A(DATA_IN_3_), .B(KEYINPUT15), .ZN(n1779) );
NAND2_X1 U1354 ( .A1(DATA_IN_4_), .A2(n1780), .ZN(n1758) );
NAND2_X1 U1355 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1781), .ZN(n1754) );
XOR2_X1 U1356 ( .A(KEYINPUT48), .B(DATA_IN_5_), .Z(n1781) );
NAND2_X1 U1357 ( .A1(DATA_IN_6_), .A2(n1782), .ZN(n1750) );
NAND2_X1 U1358 ( .A1(DATA_IN_7_), .A2(n1783), .ZN(n1748) );
AND2_X1 U1359 ( .A1(n1694), .A2(n1784), .ZN(n1743) );
NAND2_X1 U1360 ( .A1(n1785), .A2(n1717), .ZN(n1784) );
NAND2_X1 U1361 ( .A1(n1716), .A2(n1718), .ZN(n1785) );
NAND2_X1 U1362 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1753), .ZN(n1718) );
NAND3_X1 U1363 ( .A1(n1786), .A2(n1787), .A3(n1788), .ZN(n1716) );
XOR2_X1 U1364 ( .A(n1789), .B(KEYINPUT63), .Z(n1788) );
NAND2_X1 U1365 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1757), .ZN(n1789) );
NAND3_X1 U1366 ( .A1(n1790), .A2(n1791), .A3(n1792), .ZN(n1787) );
OR2_X1 U1367 ( .A1(n1757), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1792) );
NAND3_X1 U1368 ( .A1(n1793), .A2(n1794), .A3(n1795), .ZN(n1791) );
NAND2_X1 U1369 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1706), .ZN(n1795) );
NAND3_X1 U1370 ( .A1(n1796), .A2(n1797), .A3(n1798), .ZN(n1794) );
NAND2_X1 U1371 ( .A1(DATA_IN_3_), .A2(n1799), .ZN(n1798) );
NAND3_X1 U1372 ( .A1(n1800), .A2(n1801), .A3(n1802), .ZN(n1797) );
OR2_X1 U1373 ( .A1(n1803), .A2(DATA_IN_2_), .ZN(n1802) );
NAND3_X1 U1374 ( .A1(n1804), .A2(n1805), .A3(n1806), .ZN(n1801) );
XOR2_X1 U1375 ( .A(KEYINPUT46), .B(n1807), .Z(n1806) );
NOR3_X1 U1376 ( .A1(n1774), .A2(RMAX_REG_0__SCAN_IN), .A3(n1808), .ZN(n1807));
NOR2_X1 U1377 ( .A1(DATA_IN_1_), .A2(n1809), .ZN(n1808) );
NAND2_X1 U1378 ( .A1(DATA_IN_1_), .A2(n1809), .ZN(n1805) );
NAND2_X1 U1379 ( .A1(DATA_IN_2_), .A2(n1803), .ZN(n1804) );
NAND2_X1 U1380 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1810), .ZN(n1800) );
XOR2_X1 U1381 ( .A(KEYINPUT20), .B(DATA_IN_3_), .Z(n1810) );
NAND2_X1 U1382 ( .A1(n1811), .A2(n1812), .ZN(n1796) );
XOR2_X1 U1383 ( .A(KEYINPUT27), .B(DATA_IN_4_), .Z(n1811) );
NAND2_X1 U1384 ( .A1(n1813), .A2(RMAX_REG_5__SCAN_IN), .ZN(n1793) );
XOR2_X1 U1385 ( .A(n1814), .B(KEYINPUT3), .Z(n1813) );
NAND2_X1 U1386 ( .A1(DATA_IN_5_), .A2(n1815), .ZN(n1790) );
NAND2_X1 U1387 ( .A1(DATA_IN_7_), .A2(n1816), .ZN(n1786) );
NAND2_X1 U1388 ( .A1(n1817), .A2(n1818), .ZN(U328) );
NAND2_X1 U1389 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1819), .ZN(n1818) );
XOR2_X1 U1390 ( .A(KEYINPUT56), .B(n1820), .Z(n1817) );
NOR2_X1 U1391 ( .A1(n1753), .A2(n1821), .ZN(n1820) );
NAND2_X1 U1392 ( .A1(n1822), .A2(n1823), .ZN(U327) );
NAND2_X1 U1393 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1819), .ZN(n1823) );
XOR2_X1 U1394 ( .A(n1824), .B(KEYINPUT33), .Z(n1822) );
NAND2_X1 U1395 ( .A1(n1825), .A2(DATA_IN_6_), .ZN(n1824) );
NAND2_X1 U1396 ( .A1(n1826), .A2(n1827), .ZN(U326) );
NAND2_X1 U1397 ( .A1(n1825), .A2(DATA_IN_5_), .ZN(n1827) );
NAND2_X1 U1398 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1819), .ZN(n1826) );
NAND2_X1 U1399 ( .A1(n1828), .A2(n1829), .ZN(U325) );
NAND2_X1 U1400 ( .A1(n1825), .A2(DATA_IN_4_), .ZN(n1829) );
NAND2_X1 U1401 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1819), .ZN(n1828) );
NAND2_X1 U1402 ( .A1(n1830), .A2(n1831), .ZN(U324) );
NAND2_X1 U1403 ( .A1(DATA_IN_3_), .A2(n1832), .ZN(n1831) );
XOR2_X1 U1404 ( .A(KEYINPUT6), .B(n1825), .Z(n1832) );
NAND2_X1 U1405 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1819), .ZN(n1830) );
NAND2_X1 U1406 ( .A1(n1833), .A2(n1834), .ZN(U323) );
NAND2_X1 U1407 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1835), .ZN(n1834) );
XNOR2_X1 U1408 ( .A(KEYINPUT44), .B(n1819), .ZN(n1835) );
NAND2_X1 U1409 ( .A1(n1825), .A2(DATA_IN_2_), .ZN(n1833) );
NAND2_X1 U1410 ( .A1(n1836), .A2(n1837), .ZN(U322) );
NAND2_X1 U1411 ( .A1(n1825), .A2(DATA_IN_1_), .ZN(n1837) );
NAND2_X1 U1412 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1819), .ZN(n1836) );
NAND2_X1 U1413 ( .A1(n1838), .A2(n1839), .ZN(U321) );
NAND2_X1 U1414 ( .A1(n1825), .A2(DATA_IN_0_), .ZN(n1839) );
INV_X1 U1415 ( .A(n1821), .ZN(n1825) );
NAND2_X1 U1416 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1840), .ZN(n1821) );
NAND2_X1 U1417 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1819), .ZN(n1838) );
NAND2_X1 U1418 ( .A1(n1694), .A2(n1840), .ZN(n1819) );
NAND2_X1 U1419 ( .A1(n1841), .A2(n1842), .ZN(n1840) );
XOR2_X1 U1420 ( .A(STATO_REG_0__SCAN_IN), .B(KEYINPUT30), .Z(n1841) );
NAND2_X1 U1421 ( .A1(n1843), .A2(n1717), .ZN(n1694) );
NAND2_X1 U1422 ( .A1(n1844), .A2(n1845), .ZN(U320) );
NAND2_X1 U1423 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1693), .ZN(n1845) );
NAND2_X1 U1424 ( .A1(n1692), .A2(DATA_IN_7_), .ZN(n1844) );
NAND2_X1 U1425 ( .A1(n1846), .A2(n1847), .ZN(U319) );
NAND2_X1 U1426 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1693), .ZN(n1847) );
NAND2_X1 U1427 ( .A1(n1692), .A2(DATA_IN_6_), .ZN(n1846) );
NAND2_X1 U1428 ( .A1(n1848), .A2(n1849), .ZN(U318) );
NAND2_X1 U1429 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1693), .ZN(n1849) );
NAND2_X1 U1430 ( .A1(n1692), .A2(DATA_IN_5_), .ZN(n1848) );
NAND2_X1 U1431 ( .A1(n1850), .A2(n1851), .ZN(U317) );
NAND2_X1 U1432 ( .A1(n1692), .A2(n1852), .ZN(n1851) );
XOR2_X1 U1433 ( .A(KEYINPUT32), .B(DATA_IN_4_), .Z(n1852) );
NAND2_X1 U1434 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1693), .ZN(n1850) );
NAND2_X1 U1435 ( .A1(n1853), .A2(n1854), .ZN(U316) );
NAND2_X1 U1436 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1693), .ZN(n1854) );
NAND2_X1 U1437 ( .A1(n1692), .A2(DATA_IN_3_), .ZN(n1853) );
NAND2_X1 U1438 ( .A1(n1855), .A2(n1856), .ZN(U315) );
NAND2_X1 U1439 ( .A1(n1692), .A2(n1857), .ZN(n1856) );
XOR2_X1 U1440 ( .A(KEYINPUT31), .B(DATA_IN_2_), .Z(n1857) );
NAND2_X1 U1441 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1693), .ZN(n1855) );
NAND2_X1 U1442 ( .A1(n1858), .A2(n1859), .ZN(U314) );
NAND2_X1 U1443 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1693), .ZN(n1859) );
NAND2_X1 U1444 ( .A1(n1692), .A2(DATA_IN_1_), .ZN(n1858) );
NAND2_X1 U1445 ( .A1(n1860), .A2(n1861), .ZN(U313) );
NAND2_X1 U1446 ( .A1(n1692), .A2(n1862), .ZN(n1861) );
XOR2_X1 U1447 ( .A(KEYINPUT43), .B(DATA_IN_0_), .Z(n1862) );
NAND2_X1 U1448 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1693), .ZN(n1860) );
NAND2_X1 U1449 ( .A1(n1863), .A2(n1864), .ZN(U312) );
NAND2_X1 U1450 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1693), .ZN(n1864) );
NAND2_X1 U1451 ( .A1(n1692), .A2(REG1_REG_7__SCAN_IN), .ZN(n1863) );
NAND2_X1 U1452 ( .A1(n1865), .A2(n1866), .ZN(U311) );
NAND2_X1 U1453 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1693), .ZN(n1866) );
NAND2_X1 U1454 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1692), .ZN(n1865) );
NAND2_X1 U1455 ( .A1(n1867), .A2(n1868), .ZN(U310) );
NAND2_X1 U1456 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1693), .ZN(n1868) );
NAND2_X1 U1457 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1692), .ZN(n1867) );
NAND2_X1 U1458 ( .A1(n1869), .A2(n1870), .ZN(U309) );
NAND2_X1 U1459 ( .A1(n1871), .A2(n1693), .ZN(n1870) );
XOR2_X1 U1460 ( .A(REG2_REG_4__SCAN_IN), .B(KEYINPUT1), .Z(n1871) );
NAND2_X1 U1461 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1692), .ZN(n1869) );
NAND2_X1 U1462 ( .A1(n1872), .A2(n1873), .ZN(U308) );
NAND2_X1 U1463 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1693), .ZN(n1873) );
XOR2_X1 U1464 ( .A(KEYINPUT25), .B(n1874), .Z(n1872) );
AND2_X1 U1465 ( .A1(n1692), .A2(REG1_REG_3__SCAN_IN), .ZN(n1874) );
NAND2_X1 U1466 ( .A1(n1875), .A2(n1876), .ZN(U307) );
NAND2_X1 U1467 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1693), .ZN(n1876) );
NAND2_X1 U1468 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1692), .ZN(n1875) );
NAND2_X1 U1469 ( .A1(n1877), .A2(n1878), .ZN(U306) );
NAND2_X1 U1470 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1693), .ZN(n1878) );
NAND2_X1 U1471 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1692), .ZN(n1877) );
NAND2_X1 U1472 ( .A1(n1879), .A2(n1880), .ZN(U305) );
NAND2_X1 U1473 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1693), .ZN(n1880) );
NAND2_X1 U1474 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1692), .ZN(n1879) );
NAND2_X1 U1475 ( .A1(n1881), .A2(n1882), .ZN(U304) );
NAND2_X1 U1476 ( .A1(n1692), .A2(n1883), .ZN(n1882) );
XOR2_X1 U1477 ( .A(REG2_REG_7__SCAN_IN), .B(KEYINPUT18), .Z(n1883) );
NAND2_X1 U1478 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1693), .ZN(n1881) );
NAND2_X1 U1479 ( .A1(n1884), .A2(n1885), .ZN(U303) );
NAND2_X1 U1480 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1693), .ZN(n1885) );
NAND2_X1 U1481 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1692), .ZN(n1884) );
NAND2_X1 U1482 ( .A1(n1886), .A2(n1887), .ZN(U302) );
NAND2_X1 U1483 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1693), .ZN(n1887) );
NAND2_X1 U1484 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1692), .ZN(n1886) );
NAND2_X1 U1485 ( .A1(n1888), .A2(n1889), .ZN(U301) );
NAND2_X1 U1486 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1693), .ZN(n1889) );
NAND2_X1 U1487 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1692), .ZN(n1888) );
NAND2_X1 U1488 ( .A1(n1890), .A2(n1891), .ZN(U300) );
NAND2_X1 U1489 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1693), .ZN(n1891) );
NAND2_X1 U1490 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1692), .ZN(n1890) );
NAND2_X1 U1491 ( .A1(n1892), .A2(n1893), .ZN(U299) );
NAND2_X1 U1492 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1693), .ZN(n1893) );
NAND2_X1 U1493 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1692), .ZN(n1892) );
NAND2_X1 U1494 ( .A1(n1894), .A2(n1895), .ZN(U298) );
NAND2_X1 U1495 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1693), .ZN(n1895) );
NAND2_X1 U1496 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1692), .ZN(n1894) );
NAND2_X1 U1497 ( .A1(n1896), .A2(n1897), .ZN(U297) );
NAND2_X1 U1498 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1693), .ZN(n1897) );
NAND2_X1 U1499 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1692), .ZN(n1896) );
NAND2_X1 U1500 ( .A1(n1898), .A2(n1899), .ZN(U296) );
NAND2_X1 U1501 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1693), .ZN(n1899) );
NAND2_X1 U1502 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1692), .ZN(n1898) );
NAND2_X1 U1503 ( .A1(n1900), .A2(n1901), .ZN(U295) );
NAND2_X1 U1504 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1693), .ZN(n1901) );
NAND2_X1 U1505 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1692), .ZN(n1900) );
NAND2_X1 U1506 ( .A1(n1902), .A2(n1903), .ZN(U294) );
NAND2_X1 U1507 ( .A1(n1904), .A2(n1692), .ZN(n1903) );
XNOR2_X1 U1508 ( .A(REG3_REG_5__SCAN_IN), .B(KEYINPUT45), .ZN(n1904) );
NAND2_X1 U1509 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1693), .ZN(n1902) );
NAND2_X1 U1510 ( .A1(n1905), .A2(n1906), .ZN(U293) );
NAND2_X1 U1511 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1907), .ZN(n1906) );
XOR2_X1 U1512 ( .A(KEYINPUT57), .B(n1693), .Z(n1907) );
NAND2_X1 U1513 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1692), .ZN(n1905) );
NAND2_X1 U1514 ( .A1(n1908), .A2(n1909), .ZN(U292) );
NAND2_X1 U1515 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1693), .ZN(n1909) );
NAND2_X1 U1516 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1692), .ZN(n1908) );
NAND2_X1 U1517 ( .A1(n1910), .A2(n1911), .ZN(U291) );
NAND2_X1 U1518 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1693), .ZN(n1911) );
NAND2_X1 U1519 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1692), .ZN(n1910) );
NAND2_X1 U1520 ( .A1(n1912), .A2(n1913), .ZN(U290) );
NAND2_X1 U1521 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1693), .ZN(n1913) );
NAND2_X1 U1522 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1692), .ZN(n1912) );
NAND2_X1 U1523 ( .A1(n1914), .A2(n1915), .ZN(U289) );
NAND2_X1 U1524 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1693), .ZN(n1915) );
NAND2_X1 U1525 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1692), .ZN(n1914) );
NAND4_X1 U1526 ( .A1(n1916), .A2(n1917), .A3(n1918), .A4(n1919), .ZN(U288));
NOR2_X1 U1527 ( .A1(n1920), .A2(n1921), .ZN(n1919) );
NOR2_X1 U1528 ( .A1(n1922), .A2(n1923), .ZN(n1921) );
AND2_X1 U1529 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1924), .ZN(n1920) );
NAND2_X1 U1530 ( .A1(n1925), .A2(n1926), .ZN(n1918) );
INV_X1 U1531 ( .A(n1927), .ZN(n1925) );
NAND3_X1 U1532 ( .A1(n1928), .A2(n1929), .A3(n1930), .ZN(n1917) );
XOR2_X1 U1533 ( .A(n1931), .B(KEYINPUT8), .Z(n1930) );
NAND2_X1 U1534 ( .A1(n1932), .A2(DATA_OUT_REG_7__SCAN_IN), .ZN(n1916) );
XOR2_X1 U1535 ( .A(U280), .B(KEYINPUT41), .Z(n1932) );
NAND4_X1 U1536 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(U287));
NOR3_X1 U1537 ( .A1(n1937), .A2(n1938), .A3(n1939), .ZN(n1936) );
AND2_X1 U1538 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1924), .ZN(n1939) );
NOR2_X1 U1539 ( .A1(n1940), .A2(n1931), .ZN(n1938) );
XOR2_X1 U1540 ( .A(n1941), .B(n1942), .Z(n1940) );
NOR2_X1 U1541 ( .A1(n1943), .A2(n1923), .ZN(n1937) );
NAND2_X1 U1542 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1693), .ZN(n1935) );
OR2_X1 U1543 ( .A1(n1927), .A2(n1944), .ZN(n1934) );
NAND4_X1 U1544 ( .A1(n1945), .A2(n1946), .A3(n1947), .A4(n1944), .ZN(n1933));
NOR2_X1 U1545 ( .A1(n1948), .A2(n1926), .ZN(n1944) );
INV_X1 U1546 ( .A(KEYINPUT40), .ZN(n1948) );
NAND4_X1 U1547 ( .A1(n1949), .A2(n1950), .A3(n1951), .A4(n1952), .ZN(U286));
NOR3_X1 U1548 ( .A1(n1953), .A2(n1954), .A3(n1955), .ZN(n1952) );
NOR2_X1 U1549 ( .A1(n1956), .A2(n1927), .ZN(n1955) );
NAND2_X1 U1550 ( .A1(n1947), .A2(n1957), .ZN(n1927) );
NAND2_X1 U1551 ( .A1(n1945), .A2(n1946), .ZN(n1957) );
NOR2_X1 U1552 ( .A1(n1945), .A2(n1946), .ZN(n1956) );
NAND2_X1 U1553 ( .A1(n1958), .A2(n1959), .ZN(n1946) );
NAND2_X1 U1554 ( .A1(n1960), .A2(n1961), .ZN(n1959) );
XNOR2_X1 U1555 ( .A(n1926), .B(KEYINPUT24), .ZN(n1958) );
NOR2_X1 U1556 ( .A1(n1961), .A2(n1960), .ZN(n1926) );
NOR3_X1 U1557 ( .A1(n1931), .A2(n1942), .A3(n1962), .ZN(n1954) );
NOR3_X1 U1558 ( .A1(n1963), .A2(n1964), .A3(n1928), .ZN(n1962) );
INV_X1 U1559 ( .A(n1941), .ZN(n1928) );
NOR2_X1 U1560 ( .A1(n1965), .A2(n1966), .ZN(n1963) );
INV_X1 U1561 ( .A(n1929), .ZN(n1942) );
NAND2_X1 U1562 ( .A1(n1964), .A2(n1967), .ZN(n1929) );
NAND2_X1 U1563 ( .A1(n1968), .A2(n1941), .ZN(n1967) );
NAND2_X1 U1564 ( .A1(n1965), .A2(n1966), .ZN(n1941) );
NAND2_X1 U1565 ( .A1(n1960), .A2(n1969), .ZN(n1968) );
INV_X1 U1566 ( .A(n1966), .ZN(n1960) );
NOR2_X1 U1567 ( .A1(n1966), .A2(n1970), .ZN(n1953) );
NAND2_X1 U1568 ( .A1(n1971), .A2(n1972), .ZN(n1966) );
NAND3_X1 U1569 ( .A1(n1973), .A2(n1974), .A3(n1975), .ZN(n1972) );
NAND2_X1 U1570 ( .A1(n1976), .A2(n1977), .ZN(n1974) );
NAND2_X1 U1571 ( .A1(n1978), .A2(n1979), .ZN(n1977) );
NAND2_X1 U1572 ( .A1(n1980), .A2(n1981), .ZN(n1973) );
NAND4_X1 U1573 ( .A1(n1982), .A2(n1983), .A3(n1984), .A4(n1985), .ZN(n1971));
NAND3_X1 U1574 ( .A1(n1986), .A2(n1987), .A3(n1988), .ZN(n1985) );
INV_X1 U1575 ( .A(KEYINPUT21), .ZN(n1988) );
NAND2_X1 U1576 ( .A1(n1975), .A2(KEYINPUT21), .ZN(n1984) );
XNOR2_X1 U1577 ( .A(n1987), .B(n1989), .ZN(n1975) );
NOR2_X1 U1578 ( .A1(n1986), .A2(KEYINPUT60), .ZN(n1989) );
AND2_X1 U1579 ( .A1(n1990), .A2(n1991), .ZN(n1986) );
NAND2_X1 U1580 ( .A1(n1992), .A2(n1993), .ZN(n1991) );
XOR2_X1 U1581 ( .A(KEYINPUT23), .B(DATA_IN_6_), .Z(n1992) );
NAND2_X1 U1582 ( .A1(RESTART), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1990) );
NAND2_X1 U1583 ( .A1(n1994), .A2(n1995), .ZN(n1987) );
NAND2_X1 U1584 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1993), .ZN(n1995) );
NAND2_X1 U1585 ( .A1(RESTART), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1994) );
NAND2_X1 U1586 ( .A1(n1979), .A2(n1996), .ZN(n1983) );
NAND2_X1 U1587 ( .A1(n1976), .A2(n1997), .ZN(n1996) );
XOR2_X1 U1588 ( .A(KEYINPUT17), .B(n1978), .Z(n1997) );
INV_X1 U1589 ( .A(n1998), .ZN(n1976) );
NAND2_X1 U1590 ( .A1(n1978), .A2(n1998), .ZN(n1982) );
NAND2_X1 U1591 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1693), .ZN(n1951) );
NAND2_X1 U1592 ( .A1(n1924), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1950) );
NAND2_X1 U1593 ( .A1(n1999), .A2(REG4_REG_5__SCAN_IN), .ZN(n1949) );
NAND4_X1 U1594 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(U285));
NOR3_X1 U1595 ( .A1(n2004), .A2(n2005), .A3(n2006), .ZN(n2003) );
NOR3_X1 U1596 ( .A1(n1931), .A2(n1964), .A3(n2007), .ZN(n2006) );
NOR2_X1 U1597 ( .A1(n2008), .A2(n2009), .ZN(n2007) );
AND2_X1 U1598 ( .A1(n2008), .A2(n2009), .ZN(n1964) );
NAND3_X1 U1599 ( .A1(n2010), .A2(n2011), .A3(n1969), .ZN(n2009) );
INV_X1 U1600 ( .A(n1965), .ZN(n1969) );
NOR2_X1 U1601 ( .A1(n2012), .A2(n2013), .ZN(n1965) );
NAND3_X1 U1602 ( .A1(KEYINPUT9), .A2(n2013), .A3(n2012), .ZN(n2011) );
OR2_X1 U1603 ( .A1(n2012), .A2(KEYINPUT9), .ZN(n2010) );
NOR3_X1 U1604 ( .A1(n2014), .A2(n1945), .A3(n2015), .ZN(n2005) );
NOR2_X1 U1605 ( .A1(n2016), .A2(n2017), .ZN(n2015) );
AND2_X1 U1606 ( .A1(n2016), .A2(n2017), .ZN(n1945) );
NAND2_X1 U1607 ( .A1(n1961), .A2(n2018), .ZN(n2017) );
NAND2_X1 U1608 ( .A1(n2013), .A2(n2019), .ZN(n2018) );
OR2_X1 U1609 ( .A1(n2019), .A2(n2013), .ZN(n1961) );
INV_X1 U1610 ( .A(n2020), .ZN(n2013) );
NOR2_X1 U1611 ( .A1(n2020), .A2(n1970), .ZN(n2004) );
XOR2_X1 U1612 ( .A(n2021), .B(n1979), .Z(n2020) );
INV_X1 U1613 ( .A(n1980), .ZN(n1979) );
NAND2_X1 U1614 ( .A1(n2022), .A2(n2023), .ZN(n1980) );
NAND2_X1 U1615 ( .A1(n2024), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2023) );
XOR2_X1 U1616 ( .A(n2025), .B(KEYINPUT28), .Z(n2024) );
XOR2_X1 U1617 ( .A(KEYINPUT11), .B(n2026), .Z(n2022) );
NOR2_X1 U1618 ( .A1(n2027), .A2(n2028), .ZN(n2026) );
XOR2_X1 U1619 ( .A(n1998), .B(n1978), .Z(n2021) );
INV_X1 U1620 ( .A(n1981), .ZN(n1978) );
NAND2_X1 U1621 ( .A1(n2029), .A2(n2030), .ZN(n1981) );
NAND2_X1 U1622 ( .A1(DATA_IN_5_), .A2(n1993), .ZN(n2030) );
NAND2_X1 U1623 ( .A1(RESTART), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2029) );
NAND2_X1 U1624 ( .A1(n2031), .A2(n2032), .ZN(n1998) );
NAND2_X1 U1625 ( .A1(n2033), .A2(n2034), .ZN(n2032) );
NAND2_X1 U1626 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
OR2_X1 U1627 ( .A1(n2036), .A2(n2035), .ZN(n2031) );
NAND2_X1 U1628 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1693), .ZN(n2002) );
NAND2_X1 U1629 ( .A1(n1924), .A2(RLAST_REG_4__SCAN_IN), .ZN(n2001) );
NAND2_X1 U1630 ( .A1(n1999), .A2(REG4_REG_4__SCAN_IN), .ZN(n2000) );
NAND4_X1 U1631 ( .A1(n2037), .A2(n2038), .A3(n2039), .A4(n2040), .ZN(U284));
NOR3_X1 U1632 ( .A1(n2041), .A2(n2042), .A3(n2043), .ZN(n2040) );
NOR3_X1 U1633 ( .A1(n2014), .A2(n2016), .A3(n2044), .ZN(n2043) );
NOR2_X1 U1634 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
AND2_X1 U1635 ( .A1(n2045), .A2(n2046), .ZN(n2016) );
NAND2_X1 U1636 ( .A1(n2019), .A2(n2047), .ZN(n2046) );
NAND2_X1 U1637 ( .A1(n2048), .A2(n2049), .ZN(n2047) );
OR2_X1 U1638 ( .A1(n2049), .A2(n2048), .ZN(n2019) );
NOR3_X1 U1639 ( .A1(n1931), .A2(n2008), .A3(n2050), .ZN(n2042) );
NOR2_X1 U1640 ( .A1(n2051), .A2(n2052), .ZN(n2050) );
AND2_X1 U1641 ( .A1(n2051), .A2(n2052), .ZN(n2008) );
NAND2_X1 U1642 ( .A1(n2012), .A2(n2053), .ZN(n2052) );
NAND2_X1 U1643 ( .A1(n2048), .A2(n2054), .ZN(n2053) );
OR2_X1 U1644 ( .A1(n2054), .A2(n2048), .ZN(n2012) );
NOR2_X1 U1645 ( .A1(n2055), .A2(n1970), .ZN(n2041) );
INV_X1 U1646 ( .A(n2048), .ZN(n2055) );
XNOR2_X1 U1647 ( .A(n2056), .B(n2035), .ZN(n2048) );
NAND2_X1 U1648 ( .A1(n2057), .A2(n2058), .ZN(n2035) );
NAND2_X1 U1649 ( .A1(n2059), .A2(n2060), .ZN(n2058) );
NAND2_X1 U1650 ( .A1(n2061), .A2(n2062), .ZN(n2060) );
XOR2_X1 U1651 ( .A(KEYINPUT49), .B(n2063), .Z(n2057) );
NOR2_X1 U1652 ( .A1(n2062), .A2(n2061), .ZN(n2063) );
XOR2_X1 U1653 ( .A(n2033), .B(n2036), .Z(n2056) );
NAND2_X1 U1654 ( .A1(n2064), .A2(n2065), .ZN(n2036) );
NAND2_X1 U1655 ( .A1(RESTART), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2065) );
XOR2_X1 U1656 ( .A(KEYINPUT34), .B(n2066), .Z(n2064) );
NOR2_X1 U1657 ( .A1(n2027), .A2(n2067), .ZN(n2066) );
AND2_X1 U1658 ( .A1(n2068), .A2(n2069), .ZN(n2033) );
NAND2_X1 U1659 ( .A1(DATA_IN_4_), .A2(n1993), .ZN(n2069) );
NAND2_X1 U1660 ( .A1(RESTART), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2068) );
NAND2_X1 U1661 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1693), .ZN(n2039) );
NAND2_X1 U1662 ( .A1(n1924), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2038) );
NAND2_X1 U1663 ( .A1(n1999), .A2(REG4_REG_3__SCAN_IN), .ZN(n2037) );
NAND4_X1 U1664 ( .A1(n2070), .A2(n2071), .A3(n2072), .A4(n2073), .ZN(U283));
NOR3_X1 U1665 ( .A1(n2074), .A2(n2075), .A3(n2076), .ZN(n2073) );
NOR2_X1 U1666 ( .A1(n1931), .A2(n2077), .ZN(n2076) );
XOR2_X1 U1667 ( .A(KEYINPUT29), .B(n2078), .Z(n2077) );
NOR2_X1 U1668 ( .A1(n2051), .A2(n2079), .ZN(n2078) );
NOR2_X1 U1669 ( .A1(n2080), .A2(n2081), .ZN(n2079) );
NOR2_X1 U1670 ( .A1(n2082), .A2(n2083), .ZN(n2080) );
XOR2_X1 U1671 ( .A(KEYINPUT14), .B(n2084), .Z(n2083) );
AND3_X1 U1672 ( .A1(n2081), .A2(n2085), .A3(n2084), .ZN(n2051) );
NAND2_X1 U1673 ( .A1(n2086), .A2(n2054), .ZN(n2081) );
NAND2_X1 U1674 ( .A1(n2087), .A2(n2088), .ZN(n2054) );
XOR2_X1 U1675 ( .A(KEYINPUT0), .B(n2089), .Z(n2088) );
XOR2_X1 U1676 ( .A(n2090), .B(KEYINPUT50), .Z(n2086) );
INV_X1 U1677 ( .A(n2091), .ZN(n1931) );
NOR3_X1 U1678 ( .A1(n2014), .A2(n2045), .A3(n2092), .ZN(n2075) );
NOR2_X1 U1679 ( .A1(n2093), .A2(n2094), .ZN(n2092) );
NOR2_X1 U1680 ( .A1(n2095), .A2(n2096), .ZN(n2093) );
AND3_X1 U1681 ( .A1(n2094), .A2(n2097), .A3(n2084), .ZN(n2045) );
NAND2_X1 U1682 ( .A1(n2049), .A2(n2090), .ZN(n2094) );
NAND2_X1 U1683 ( .A1(n2098), .A2(n2099), .ZN(n2090) );
NAND2_X1 U1684 ( .A1(n2100), .A2(n2087), .ZN(n2049) );
XOR2_X1 U1685 ( .A(n2099), .B(KEYINPUT22), .Z(n2100) );
INV_X1 U1686 ( .A(n1947), .ZN(n2014) );
NOR2_X1 U1687 ( .A1(n2087), .A2(n1970), .ZN(n2074) );
INV_X1 U1688 ( .A(n2098), .ZN(n2087) );
XNOR2_X1 U1689 ( .A(n2061), .B(n2101), .ZN(n2098) );
NOR2_X1 U1690 ( .A1(n2102), .A2(n2103), .ZN(n2101) );
NOR3_X1 U1691 ( .A1(n2104), .A2(KEYINPUT54), .A3(n2062), .ZN(n2103) );
INV_X1 U1692 ( .A(n2105), .ZN(n2062) );
NOR2_X1 U1693 ( .A1(n2059), .A2(n2105), .ZN(n2102) );
NAND2_X1 U1694 ( .A1(n2106), .A2(n2107), .ZN(n2105) );
NAND2_X1 U1695 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1993), .ZN(n2107) );
NAND2_X1 U1696 ( .A1(RESTART), .A2(RMIN_REG_3__SCAN_IN), .ZN(n2106) );
INV_X1 U1697 ( .A(n2104), .ZN(n2059) );
NAND2_X1 U1698 ( .A1(n2108), .A2(n2109), .ZN(n2104) );
NAND2_X1 U1699 ( .A1(n2110), .A2(n2111), .ZN(n2109) );
NAND2_X1 U1700 ( .A1(n2112), .A2(n2113), .ZN(n2111) );
OR2_X1 U1701 ( .A1(n2113), .A2(n2112), .ZN(n2108) );
AND2_X1 U1702 ( .A1(n2114), .A2(n2115), .ZN(n2061) );
NAND2_X1 U1703 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n2116), .ZN(n2115) );
XOR2_X1 U1704 ( .A(RESTART), .B(KEYINPUT55), .Z(n2116) );
NAND2_X1 U1705 ( .A1(DATA_IN_3_), .A2(n1993), .ZN(n2114) );
XOR2_X1 U1706 ( .A(n2117), .B(KEYINPUT5), .Z(n2072) );
NAND2_X1 U1707 ( .A1(REG4_REG_2__SCAN_IN), .A2(n2118), .ZN(n2117) );
XOR2_X1 U1708 ( .A(KEYINPUT59), .B(n1999), .Z(n2118) );
NAND2_X1 U1709 ( .A1(n1924), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2071) );
NAND2_X1 U1710 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1693), .ZN(n2070) );
NAND4_X1 U1711 ( .A1(n2119), .A2(n2120), .A3(n2121), .A4(n2122), .ZN(U282));
NOR3_X1 U1712 ( .A1(n2123), .A2(n2124), .A3(n2125), .ZN(n2122) );
AND2_X1 U1713 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1924), .ZN(n2125) );
NOR2_X1 U1714 ( .A1(n2126), .A2(n1970), .ZN(n2124) );
NOR2_X1 U1715 ( .A1(n2127), .A2(n1923), .ZN(n2123) );
NAND2_X1 U1716 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1693), .ZN(n2121) );
NAND2_X1 U1717 ( .A1(n2084), .A2(n2128), .ZN(n2120) );
NAND2_X1 U1718 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
NAND2_X1 U1719 ( .A1(n2095), .A2(n1947), .ZN(n2130) );
INV_X1 U1720 ( .A(n2097), .ZN(n2095) );
NAND2_X1 U1721 ( .A1(n2082), .A2(n2091), .ZN(n2129) );
INV_X1 U1722 ( .A(n2085), .ZN(n2082) );
INV_X1 U1723 ( .A(n2096), .ZN(n2084) );
NAND2_X1 U1724 ( .A1(n2096), .A2(n2131), .ZN(n2119) );
NAND2_X1 U1725 ( .A1(n2132), .A2(n2133), .ZN(n2131) );
NAND2_X1 U1726 ( .A1(n1947), .A2(n2097), .ZN(n2133) );
NAND2_X1 U1727 ( .A1(n2134), .A2(n2135), .ZN(n2097) );
NAND2_X1 U1728 ( .A1(n2136), .A2(n2137), .ZN(n2135) );
XOR2_X1 U1729 ( .A(n2138), .B(KEYINPUT61), .Z(n2136) );
NAND2_X1 U1730 ( .A1(n2091), .A2(n2085), .ZN(n2132) );
NAND2_X1 U1731 ( .A1(n2134), .A2(n2139), .ZN(n2085) );
NAND2_X1 U1732 ( .A1(n2140), .A2(n2137), .ZN(n2139) );
AND2_X1 U1733 ( .A1(n2099), .A2(n2141), .ZN(n2134) );
NAND2_X1 U1734 ( .A1(n2142), .A2(n2137), .ZN(n2141) );
INV_X1 U1735 ( .A(n2089), .ZN(n2099) );
NOR3_X1 U1736 ( .A1(n2142), .A2(n2140), .A3(n2137), .ZN(n2089) );
INV_X1 U1737 ( .A(n2126), .ZN(n2137) );
XNOR2_X1 U1738 ( .A(n2110), .B(n2143), .ZN(n2126) );
XNOR2_X1 U1739 ( .A(n2113), .B(n2112), .ZN(n2143) );
AND2_X1 U1740 ( .A1(n2144), .A2(n2145), .ZN(n2112) );
NAND2_X1 U1741 ( .A1(n2146), .A2(n2147), .ZN(n2145) );
NAND2_X1 U1742 ( .A1(n2148), .A2(n2149), .ZN(n2147) );
NAND2_X1 U1743 ( .A1(n2150), .A2(n2151), .ZN(n2144) );
NAND2_X1 U1744 ( .A1(n2152), .A2(n2153), .ZN(n2113) );
NAND2_X1 U1745 ( .A1(DATA_IN_2_), .A2(n1993), .ZN(n2153) );
NAND2_X1 U1746 ( .A1(RESTART), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2152) );
AND2_X1 U1747 ( .A1(n2154), .A2(n2155), .ZN(n2110) );
NAND2_X1 U1748 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1993), .ZN(n2155) );
NAND2_X1 U1749 ( .A1(RESTART), .A2(RMIN_REG_2__SCAN_IN), .ZN(n2154) );
NAND4_X1 U1750 ( .A1(n2156), .A2(n2157), .A3(n2158), .A4(n2159), .ZN(U281));
NOR3_X1 U1751 ( .A1(n2160), .A2(n2161), .A3(n2162), .ZN(n2159) );
AND2_X1 U1752 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1924), .ZN(n2162) );
NOR2_X1 U1753 ( .A1(n2163), .A2(ENABLE), .ZN(n1924) );
NOR2_X1 U1754 ( .A1(n1970), .A2(n2164), .ZN(n2161) );
XOR2_X1 U1755 ( .A(n2142), .B(KEYINPUT58), .Z(n2164) );
NAND4_X1 U1756 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2165), .A3(n2166), .A4(U280), .ZN(n1970) );
NAND2_X1 U1757 ( .A1(n1993), .A2(n2167), .ZN(n2165) );
NAND3_X1 U1758 ( .A1(n2168), .A2(n2169), .A3(ENABLE), .ZN(n2167) );
NOR2_X1 U1759 ( .A1(n2170), .A2(n1923), .ZN(n2160) );
INV_X1 U1760 ( .A(n1999), .ZN(n1923) );
NOR3_X1 U1761 ( .A1(n1842), .A2(n2163), .A3(n2169), .ZN(n1999) );
INV_X1 U1762 ( .A(AVERAGE), .ZN(n2169) );
XOR2_X1 U1763 ( .A(n2171), .B(KEYINPUT62), .Z(n2158) );
NAND2_X1 U1764 ( .A1(n2091), .A2(n2096), .ZN(n2171) );
NOR3_X1 U1765 ( .A1(n1843), .A2(n1693), .A3(n2166), .ZN(n2091) );
NAND3_X1 U1766 ( .A1(n2172), .A2(n2173), .A3(RESTART), .ZN(n2166) );
NAND2_X1 U1767 ( .A1(n2174), .A2(n2175), .ZN(n2173) );
NAND2_X1 U1768 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2175) );
NAND2_X1 U1769 ( .A1(n2176), .A2(n2177), .ZN(n2174) );
NAND2_X1 U1770 ( .A1(RMIN_REG_6__SCAN_IN), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2177) );
NAND3_X1 U1771 ( .A1(n2178), .A2(n2179), .A3(n2180), .ZN(n2176) );
NAND2_X1 U1772 ( .A1(n1815), .A2(n1761), .ZN(n2180) );
INV_X1 U1773 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1761) );
INV_X1 U1774 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1815) );
NAND3_X1 U1775 ( .A1(n2181), .A2(n2182), .A3(n2183), .ZN(n2179) );
NAND2_X1 U1776 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2183) );
NAND3_X1 U1777 ( .A1(n2184), .A2(n2185), .A3(n2186), .ZN(n2182) );
XOR2_X1 U1778 ( .A(n2187), .B(KEYINPUT12), .Z(n2186) );
NAND2_X1 U1779 ( .A1(n1780), .A2(n1812), .ZN(n2187) );
INV_X1 U1780 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1812) );
INV_X1 U1781 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1780) );
NAND3_X1 U1782 ( .A1(n2188), .A2(n2189), .A3(n2190), .ZN(n2185) );
NAND2_X1 U1783 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2190) );
NAND3_X1 U1784 ( .A1(n2191), .A2(n2192), .A3(n2193), .ZN(n2189) );
NAND2_X1 U1785 ( .A1(n1803), .A2(n1778), .ZN(n2193) );
INV_X1 U1786 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1778) );
INV_X1 U1787 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1803) );
NAND2_X1 U1788 ( .A1(n2194), .A2(n1775), .ZN(n2192) );
INV_X1 U1789 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1775) );
OR2_X1 U1790 ( .A1(n2195), .A2(n1809), .ZN(n2194) );
NAND2_X1 U1791 ( .A1(n2195), .A2(n1809), .ZN(n2191) );
INV_X1 U1792 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1809) );
NAND2_X1 U1793 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2195) );
NAND2_X1 U1794 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2188) );
NAND2_X1 U1795 ( .A1(n1799), .A2(n1768), .ZN(n2184) );
INV_X1 U1796 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1768) );
INV_X1 U1797 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1799) );
NAND2_X1 U1798 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2181) );
NAND2_X1 U1799 ( .A1(n2196), .A2(n1782), .ZN(n2178) );
INV_X1 U1800 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1782) );
XNOR2_X1 U1801 ( .A(RMAX_REG_6__SCAN_IN), .B(KEYINPUT42), .ZN(n2196) );
NAND2_X1 U1802 ( .A1(n1816), .A2(n1783), .ZN(n2172) );
INV_X1 U1803 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1783) );
INV_X1 U1804 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1816) );
NAND2_X1 U1805 ( .A1(n1947), .A2(n2096), .ZN(n2157) );
XOR2_X1 U1806 ( .A(n2142), .B(n2140), .Z(n2096) );
INV_X1 U1807 ( .A(n2138), .ZN(n2140) );
NAND2_X1 U1808 ( .A1(n2197), .A2(n2198), .ZN(n2138) );
NAND2_X1 U1809 ( .A1(n2199), .A2(n2200), .ZN(n2198) );
NAND2_X1 U1810 ( .A1(n2201), .A2(n2202), .ZN(n2200) );
INV_X1 U1811 ( .A(KEYINPUT35), .ZN(n2201) );
INV_X1 U1812 ( .A(n2203), .ZN(n2199) );
OR2_X1 U1813 ( .A1(n2151), .A2(KEYINPUT35), .ZN(n2197) );
NAND2_X1 U1814 ( .A1(n2204), .A2(n2205), .ZN(n2142) );
NAND2_X1 U1815 ( .A1(n2206), .A2(n2149), .ZN(n2205) );
NAND2_X1 U1816 ( .A1(n2207), .A2(n2208), .ZN(n2206) );
NAND2_X1 U1817 ( .A1(n2209), .A2(n2151), .ZN(n2208) );
NAND2_X1 U1818 ( .A1(n2210), .A2(n2211), .ZN(n2209) );
NAND2_X1 U1819 ( .A1(n2212), .A2(n2210), .ZN(n2207) );
NAND2_X1 U1820 ( .A1(n2213), .A2(n2150), .ZN(n2204) );
INV_X1 U1821 ( .A(n2149), .ZN(n2150) );
NAND2_X1 U1822 ( .A1(n2214), .A2(n2215), .ZN(n2149) );
NAND2_X1 U1823 ( .A1(DATA_IN_1_), .A2(n1993), .ZN(n2215) );
NAND2_X1 U1824 ( .A1(RESTART), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2214) );
XOR2_X1 U1825 ( .A(KEYINPUT10), .B(n2216), .Z(n2213) );
NOR2_X1 U1826 ( .A1(n2212), .A2(n2217), .ZN(n2216) );
NOR2_X1 U1827 ( .A1(n2211), .A2(n2148), .ZN(n2217) );
XOR2_X1 U1828 ( .A(n2151), .B(n2210), .Z(n2148) );
INV_X1 U1829 ( .A(KEYINPUT2), .ZN(n2210) );
NOR2_X1 U1830 ( .A1(n2151), .A2(n2146), .ZN(n2212) );
INV_X1 U1831 ( .A(n2211), .ZN(n2146) );
NAND2_X1 U1832 ( .A1(n2218), .A2(n2219), .ZN(n2211) );
NAND2_X1 U1833 ( .A1(n2220), .A2(n1993), .ZN(n2219) );
XOR2_X1 U1834 ( .A(REG4_REG_1__SCAN_IN), .B(KEYINPUT36), .Z(n2220) );
NAND2_X1 U1835 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2218) );
NAND2_X1 U1836 ( .A1(n2203), .A2(n2202), .ZN(n2151) );
NAND2_X1 U1837 ( .A1(n2221), .A2(n2222), .ZN(n2202) );
NAND2_X1 U1838 ( .A1(DATA_IN_0_), .A2(n1993), .ZN(n2222) );
NAND2_X1 U1839 ( .A1(RESTART), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2221) );
NAND2_X1 U1840 ( .A1(n2223), .A2(n2224), .ZN(n2203) );
NAND2_X1 U1841 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n2225), .ZN(n2224) );
XOR2_X1 U1842 ( .A(RESTART), .B(KEYINPUT53), .Z(n2225) );
NAND2_X1 U1843 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1993), .ZN(n2223) );
NAND2_X1 U1844 ( .A1(n2226), .A2(n2227), .ZN(n2168) );
NAND2_X1 U1845 ( .A1(n2228), .A2(n1922), .ZN(n2227) );
INV_X1 U1846 ( .A(REG4_REG_7__SCAN_IN), .ZN(n1922) );
OR2_X1 U1847 ( .A1(n2229), .A2(n1753), .ZN(n2228) );
NAND2_X1 U1848 ( .A1(n2229), .A2(n1753), .ZN(n2226) );
INV_X1 U1849 ( .A(DATA_IN_7_), .ZN(n1753) );
NAND2_X1 U1850 ( .A1(n2230), .A2(n2231), .ZN(n2229) );
NAND2_X1 U1851 ( .A1(n2232), .A2(n2233), .ZN(n2231) );
NAND2_X1 U1852 ( .A1(n1943), .A2(n1757), .ZN(n2233) );
INV_X1 U1853 ( .A(DATA_IN_6_), .ZN(n1757) );
INV_X1 U1854 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1943) );
NAND2_X1 U1855 ( .A1(n2234), .A2(n2235), .ZN(n2232) );
NAND2_X1 U1856 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2235) );
NAND2_X1 U1857 ( .A1(n2236), .A2(n2237), .ZN(n2234) );
NAND2_X1 U1858 ( .A1(n2238), .A2(n2239), .ZN(n2237) );
NAND3_X1 U1859 ( .A1(n2240), .A2(n2241), .A3(n2242), .ZN(n2239) );
NAND2_X1 U1860 ( .A1(n1706), .A2(n2067), .ZN(n2242) );
INV_X1 U1861 ( .A(REG4_REG_4__SCAN_IN), .ZN(n2067) );
NAND3_X1 U1862 ( .A1(n2243), .A2(n2244), .A3(n2245), .ZN(n2241) );
NAND2_X1 U1863 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2245) );
NAND3_X1 U1864 ( .A1(n2246), .A2(n2247), .A3(n2248), .ZN(n2244) );
OR2_X1 U1865 ( .A1(DATA_IN_2_), .A2(REG4_REG_2__SCAN_IN), .ZN(n2248) );
NAND2_X1 U1866 ( .A1(n2249), .A2(n2127), .ZN(n2247) );
INV_X1 U1867 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2127) );
NAND2_X1 U1868 ( .A1(n2250), .A2(DATA_IN_1_), .ZN(n2249) );
OR2_X1 U1869 ( .A1(n2250), .A2(DATA_IN_1_), .ZN(n2246) );
NOR2_X1 U1870 ( .A1(n2170), .A2(n1774), .ZN(n2250) );
INV_X1 U1871 ( .A(DATA_IN_0_), .ZN(n1774) );
INV_X1 U1872 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2170) );
NAND2_X1 U1873 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2243) );
OR2_X1 U1874 ( .A1(DATA_IN_3_), .A2(REG4_REG_3__SCAN_IN), .ZN(n2240) );
NAND2_X1 U1875 ( .A1(n2251), .A2(REG4_REG_4__SCAN_IN), .ZN(n2238) );
XOR2_X1 U1876 ( .A(n1706), .B(KEYINPUT16), .Z(n2251) );
INV_X1 U1877 ( .A(DATA_IN_4_), .ZN(n1706) );
NAND2_X1 U1878 ( .A1(n1814), .A2(n2028), .ZN(n2236) );
INV_X1 U1879 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2028) );
INV_X1 U1880 ( .A(DATA_IN_5_), .ZN(n1814) );
NAND2_X1 U1881 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2230) );
NAND3_X1 U1882 ( .A1(n1993), .A2(U280), .A3(STATO_REG_1__SCAN_IN), .ZN(n2163) );
INV_X1 U1883 ( .A(n2027), .ZN(n1993) );
XOR2_X1 U1884 ( .A(n2025), .B(KEYINPUT51), .Z(n2027) );
INV_X1 U1885 ( .A(RESTART), .ZN(n2025) );
INV_X1 U1886 ( .A(ENABLE), .ZN(n1842) );
NAND2_X1 U1887 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1693), .ZN(n2156) );
INV_X1 U1888 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1843) );
NOR2_X1 U1889 ( .A1(n1717), .A2(STATO_REG_1__SCAN_IN), .ZN(n2252) );
INV_X1 U1890 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1717) );
endmodule


