//Key = 1010110010011010000111101101001110100110101011011010101010111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356;

XNOR2_X1 U740 ( .A(G107), .B(n1021), .ZN(G9) );
NOR2_X1 U741 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U742 ( .A1(G953), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1023) );
NOR2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR2_X1 U744 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U746 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U751 ( .A1(KEYINPUT10), .A2(n1043), .ZN(n1042) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1041) );
XNOR2_X1 U753 ( .A(n1046), .B(KEYINPUT48), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1037) );
NOR2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
AND2_X1 U756 ( .A1(n1051), .A2(KEYINPUT25), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1052), .A2(n1048), .ZN(n1033) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1040), .ZN(n1054) );
NOR2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR3_X1 U762 ( .A1(n1060), .A2(KEYINPUT25), .A3(n1061), .ZN(n1053) );
NOR3_X1 U763 ( .A1(n1036), .A2(n1062), .A3(n1040), .ZN(n1029) );
NOR2_X1 U764 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U765 ( .A1(n1065), .A2(n1048), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
AND3_X1 U767 ( .A1(KEYINPUT10), .A2(n1032), .A3(n1068), .ZN(n1063) );
NOR3_X1 U768 ( .A1(n1024), .A2(G953), .A3(G952), .ZN(n1022) );
AND2_X1 U769 ( .A1(n1069), .A2(n1070), .ZN(n1024) );
NOR4_X1 U770 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NOR2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1073) );
NOR2_X1 U773 ( .A1(G472), .A2(n1079), .ZN(n1078) );
NOR2_X1 U774 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U775 ( .A1(KEYINPUT49), .A2(n1082), .ZN(n1080) );
NOR2_X1 U776 ( .A1(n1083), .A2(n1084), .ZN(n1077) );
NOR2_X1 U777 ( .A1(n1085), .A2(KEYINPUT49), .ZN(n1083) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1081), .ZN(n1085) );
INV_X1 U779 ( .A(KEYINPUT47), .ZN(n1081) );
INV_X1 U780 ( .A(n1087), .ZN(n1071) );
NOR4_X1 U781 ( .A1(n1088), .A2(n1058), .A3(n1048), .A4(n1089), .ZN(n1069) );
XNOR2_X1 U782 ( .A(G475), .B(n1090), .ZN(n1089) );
XOR2_X1 U783 ( .A(n1091), .B(n1092), .Z(G72) );
XOR2_X1 U784 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U785 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U786 ( .A(n1097), .B(n1098), .Z(n1096) );
XOR2_X1 U787 ( .A(n1099), .B(n1100), .Z(n1098) );
XNOR2_X1 U788 ( .A(KEYINPUT9), .B(n1101), .ZN(n1100) );
XNOR2_X1 U789 ( .A(n1102), .B(n1103), .ZN(n1097) );
NOR2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1095) );
XNOR2_X1 U791 ( .A(KEYINPUT28), .B(n1106), .ZN(n1105) );
NAND2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(n1093) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U794 ( .A(G953), .B(KEYINPUT33), .ZN(n1107) );
NAND2_X1 U795 ( .A1(G953), .A2(n1111), .ZN(n1091) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1111) );
XOR2_X1 U797 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U798 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U799 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NAND2_X1 U800 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NAND2_X1 U801 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U802 ( .A(G953), .B(KEYINPUT12), .ZN(n1119) );
XOR2_X1 U803 ( .A(n1121), .B(n1122), .Z(n1117) );
NAND2_X1 U804 ( .A1(G953), .A2(n1123), .ZN(n1112) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1123) );
NOR2_X1 U806 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XNOR2_X1 U807 ( .A(n1126), .B(n1127), .ZN(n1125) );
NOR2_X1 U808 ( .A1(n1076), .A2(n1128), .ZN(n1127) );
NOR2_X1 U809 ( .A1(n1124), .A2(n1129), .ZN(G63) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U811 ( .A1(KEYINPUT46), .A2(n1132), .ZN(n1131) );
XNOR2_X1 U812 ( .A(n1133), .B(KEYINPUT23), .ZN(n1132) );
NAND2_X1 U813 ( .A1(n1134), .A2(G478), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1124), .A2(n1135), .ZN(G60) );
XNOR2_X1 U815 ( .A(n1136), .B(n1137), .ZN(n1135) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1128), .ZN(n1137) );
NAND2_X1 U817 ( .A1(n1139), .A2(n1140), .ZN(G6) );
NAND2_X1 U818 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XNOR2_X1 U819 ( .A(KEYINPUT55), .B(n1143), .ZN(n1141) );
NAND2_X1 U820 ( .A1(n1144), .A2(G104), .ZN(n1139) );
XNOR2_X1 U821 ( .A(KEYINPUT44), .B(n1143), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1124), .A2(n1145), .ZN(G57) );
XOR2_X1 U823 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U824 ( .A(n1148), .B(n1149), .ZN(n1147) );
XOR2_X1 U825 ( .A(n1150), .B(n1151), .Z(n1146) );
NOR2_X1 U826 ( .A1(n1086), .A2(n1128), .ZN(n1151) );
NAND2_X1 U827 ( .A1(KEYINPUT59), .A2(n1152), .ZN(n1150) );
NOR2_X1 U828 ( .A1(n1153), .A2(n1154), .ZN(G54) );
XOR2_X1 U829 ( .A(KEYINPUT35), .B(n1124), .Z(n1154) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1153) );
AND2_X1 U831 ( .A1(G469), .A2(n1134), .ZN(n1156) );
INV_X1 U832 ( .A(n1128), .ZN(n1134) );
NAND2_X1 U833 ( .A1(n1157), .A2(KEYINPUT38), .ZN(n1155) );
XOR2_X1 U834 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U836 ( .A1(KEYINPUT58), .A2(n1162), .ZN(n1161) );
OR3_X1 U837 ( .A1(n1163), .A2(n1164), .A3(KEYINPUT58), .ZN(n1160) );
NOR2_X1 U838 ( .A1(n1124), .A2(n1165), .ZN(G51) );
XOR2_X1 U839 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U840 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1166) );
NOR3_X1 U842 ( .A1(n1128), .A2(KEYINPUT13), .A3(n1172), .ZN(n1171) );
NAND2_X1 U843 ( .A1(n1173), .A2(n1026), .ZN(n1128) );
NAND3_X1 U844 ( .A1(n1116), .A2(n1109), .A3(n1174), .ZN(n1026) );
XNOR2_X1 U845 ( .A(n1110), .B(KEYINPUT27), .ZN(n1174) );
AND4_X1 U846 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1110) );
NAND2_X1 U847 ( .A1(n1179), .A2(n1180), .ZN(n1175) );
INV_X1 U848 ( .A(n1181), .ZN(n1180) );
XNOR2_X1 U849 ( .A(n1182), .B(KEYINPUT0), .ZN(n1179) );
AND4_X1 U850 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1109) );
AND4_X1 U851 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1116) );
AND4_X1 U852 ( .A1(n1143), .A2(n1021), .A3(n1191), .A4(n1192), .ZN(n1190) );
NAND3_X1 U853 ( .A1(n1193), .A2(n1067), .A3(n1194), .ZN(n1021) );
NAND3_X1 U854 ( .A1(n1194), .A2(n1193), .A3(n1066), .ZN(n1143) );
AND2_X1 U855 ( .A1(n1195), .A2(n1196), .ZN(n1189) );
NAND4_X1 U856 ( .A1(n1050), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1188) );
NAND2_X1 U857 ( .A1(KEYINPUT22), .A2(n1200), .ZN(n1199) );
NAND2_X1 U858 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
INV_X1 U859 ( .A(KEYINPUT22), .ZN(n1202) );
NAND3_X1 U860 ( .A1(n1043), .A2(n1203), .A3(n1057), .ZN(n1201) );
NAND3_X1 U861 ( .A1(n1193), .A2(n1182), .A3(n1204), .ZN(n1187) );
XNOR2_X1 U862 ( .A(G902), .B(KEYINPUT37), .ZN(n1173) );
NOR2_X1 U863 ( .A1(n1104), .A2(G952), .ZN(n1124) );
XNOR2_X1 U864 ( .A(G146), .B(n1176), .ZN(G48) );
NAND3_X1 U865 ( .A1(n1066), .A2(n1068), .A3(n1205), .ZN(n1176) );
XNOR2_X1 U866 ( .A(n1206), .B(n1207), .ZN(G45) );
NOR2_X1 U867 ( .A1(n1208), .A2(n1181), .ZN(n1207) );
NAND2_X1 U868 ( .A1(n1209), .A2(n1068), .ZN(n1181) );
XNOR2_X1 U869 ( .A(G140), .B(n1177), .ZN(G42) );
NAND4_X1 U870 ( .A1(n1051), .A2(n1066), .A3(n1210), .A4(n1211), .ZN(n1177) );
NOR2_X1 U871 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
INV_X1 U872 ( .A(n1060), .ZN(n1051) );
XNOR2_X1 U873 ( .A(G137), .B(n1178), .ZN(G39) );
NAND3_X1 U874 ( .A1(n1197), .A2(n1211), .A3(n1205), .ZN(n1178) );
XOR2_X1 U875 ( .A(n1183), .B(n1214), .Z(G36) );
NOR2_X1 U876 ( .A1(G134), .A2(KEYINPUT3), .ZN(n1214) );
NAND3_X1 U877 ( .A1(n1211), .A2(n1067), .A3(n1209), .ZN(n1183) );
XNOR2_X1 U878 ( .A(G131), .B(n1184), .ZN(G33) );
NAND3_X1 U879 ( .A1(n1066), .A2(n1211), .A3(n1209), .ZN(n1184) );
NOR3_X1 U880 ( .A1(n1213), .A2(n1212), .A3(n1215), .ZN(n1209) );
INV_X1 U881 ( .A(n1048), .ZN(n1211) );
NAND2_X1 U882 ( .A1(n1216), .A2(n1045), .ZN(n1048) );
INV_X1 U883 ( .A(n1046), .ZN(n1216) );
XNOR2_X1 U884 ( .A(n1217), .B(n1185), .ZN(G30) );
NAND3_X1 U885 ( .A1(n1068), .A2(n1067), .A3(n1205), .ZN(n1185) );
NOR4_X1 U886 ( .A1(n1218), .A2(n1213), .A3(n1212), .A4(n1219), .ZN(n1205) );
INV_X1 U887 ( .A(n1220), .ZN(n1212) );
XNOR2_X1 U888 ( .A(G128), .B(KEYINPUT54), .ZN(n1217) );
XNOR2_X1 U889 ( .A(n1221), .B(n1222), .ZN(G3) );
NOR2_X1 U890 ( .A1(n1223), .A2(n1215), .ZN(n1222) );
INV_X1 U891 ( .A(n1050), .ZN(n1215) );
XNOR2_X1 U892 ( .A(G125), .B(n1186), .ZN(G27) );
NAND4_X1 U893 ( .A1(n1068), .A2(n1220), .A3(n1066), .A4(n1224), .ZN(n1186) );
NOR2_X1 U894 ( .A1(n1060), .A2(n1036), .ZN(n1224) );
INV_X1 U895 ( .A(n1061), .ZN(n1036) );
NAND2_X1 U896 ( .A1(n1028), .A2(n1225), .ZN(n1220) );
NAND4_X1 U897 ( .A1(G953), .A2(G902), .A3(n1226), .A4(n1106), .ZN(n1225) );
INV_X1 U898 ( .A(G900), .ZN(n1106) );
XOR2_X1 U899 ( .A(G122), .B(n1227), .Z(G24) );
NOR3_X1 U900 ( .A1(n1228), .A2(n1229), .A3(n1208), .ZN(n1227) );
XNOR2_X1 U901 ( .A(n1193), .B(KEYINPUT63), .ZN(n1229) );
INV_X1 U902 ( .A(n1040), .ZN(n1193) );
NAND2_X1 U903 ( .A1(n1219), .A2(n1218), .ZN(n1040) );
XNOR2_X1 U904 ( .A(G119), .B(n1196), .ZN(G21) );
OR4_X1 U905 ( .A1(n1228), .A2(n1218), .A3(n1032), .A4(n1219), .ZN(n1196) );
INV_X1 U906 ( .A(n1230), .ZN(n1219) );
XNOR2_X1 U907 ( .A(G116), .B(n1195), .ZN(G18) );
NAND3_X1 U908 ( .A1(n1204), .A2(n1067), .A3(n1050), .ZN(n1195) );
NAND2_X1 U909 ( .A1(n1231), .A2(n1232), .ZN(n1067) );
OR2_X1 U910 ( .A1(n1208), .A2(KEYINPUT24), .ZN(n1232) );
INV_X1 U911 ( .A(n1182), .ZN(n1208) );
NOR2_X1 U912 ( .A1(n1233), .A2(n1234), .ZN(n1182) );
NAND3_X1 U913 ( .A1(n1233), .A2(n1088), .A3(KEYINPUT24), .ZN(n1231) );
XNOR2_X1 U914 ( .A(G113), .B(n1192), .ZN(G15) );
NAND3_X1 U915 ( .A1(n1204), .A2(n1066), .A3(n1050), .ZN(n1192) );
NOR2_X1 U916 ( .A1(n1218), .A2(n1230), .ZN(n1050) );
NOR2_X1 U917 ( .A1(n1233), .A2(n1088), .ZN(n1066) );
INV_X1 U918 ( .A(n1234), .ZN(n1088) );
INV_X1 U919 ( .A(n1228), .ZN(n1204) );
NAND3_X1 U920 ( .A1(n1068), .A2(n1203), .A3(n1061), .ZN(n1228) );
NOR2_X1 U921 ( .A1(n1058), .A2(n1235), .ZN(n1061) );
XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n1072), .ZN(n1235) );
INV_X1 U923 ( .A(n1059), .ZN(n1072) );
XNOR2_X1 U924 ( .A(G110), .B(n1191), .ZN(G12) );
OR2_X1 U925 ( .A1(n1060), .A2(n1223), .ZN(n1191) );
NAND2_X1 U926 ( .A1(n1197), .A2(n1194), .ZN(n1223) );
INV_X1 U927 ( .A(n1200), .ZN(n1194) );
NAND3_X1 U928 ( .A1(n1057), .A2(n1203), .A3(n1068), .ZN(n1200) );
INV_X1 U929 ( .A(n1043), .ZN(n1068) );
NAND2_X1 U930 ( .A1(n1046), .A2(n1045), .ZN(n1043) );
NAND2_X1 U931 ( .A1(G214), .A2(n1236), .ZN(n1045) );
XOR2_X1 U932 ( .A(n1237), .B(n1172), .Z(n1046) );
NAND2_X1 U933 ( .A1(G210), .A2(n1236), .ZN(n1172) );
NAND2_X1 U934 ( .A1(n1238), .A2(n1239), .ZN(n1236) );
INV_X1 U935 ( .A(G237), .ZN(n1238) );
NAND2_X1 U936 ( .A1(n1240), .A2(n1239), .ZN(n1237) );
XOR2_X1 U937 ( .A(n1241), .B(n1168), .Z(n1240) );
XOR2_X1 U938 ( .A(n1121), .B(n1242), .Z(n1168) );
NOR2_X1 U939 ( .A1(KEYINPUT53), .A2(n1122), .ZN(n1242) );
XNOR2_X1 U940 ( .A(n1243), .B(n1244), .ZN(n1122) );
XOR2_X1 U941 ( .A(G119), .B(n1245), .Z(n1244) );
NOR2_X1 U942 ( .A1(G116), .A2(KEYINPUT41), .ZN(n1245) );
XOR2_X1 U943 ( .A(n1246), .B(n1247), .Z(n1121) );
XNOR2_X1 U944 ( .A(n1248), .B(n1249), .ZN(n1247) );
XOR2_X1 U945 ( .A(KEYINPUT29), .B(G122), .Z(n1249) );
XNOR2_X1 U946 ( .A(G101), .B(n1250), .ZN(n1246) );
NOR2_X1 U947 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NOR3_X1 U948 ( .A1(KEYINPUT31), .A2(G107), .A3(n1142), .ZN(n1252) );
INV_X1 U949 ( .A(G104), .ZN(n1142) );
NOR2_X1 U950 ( .A1(n1253), .A2(n1254), .ZN(n1251) );
INV_X1 U951 ( .A(KEYINPUT31), .ZN(n1254) );
NAND3_X1 U952 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1241) );
NAND2_X1 U953 ( .A1(n1170), .A2(n1258), .ZN(n1257) );
OR3_X1 U954 ( .A1(n1258), .A2(n1170), .A3(n1169), .ZN(n1256) );
INV_X1 U955 ( .A(KEYINPUT11), .ZN(n1258) );
NAND2_X1 U956 ( .A1(n1169), .A2(n1259), .ZN(n1255) );
NAND2_X1 U957 ( .A1(KEYINPUT11), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U958 ( .A(KEYINPUT43), .B(n1170), .ZN(n1260) );
NAND2_X1 U959 ( .A1(G224), .A2(n1104), .ZN(n1170) );
XNOR2_X1 U960 ( .A(n1261), .B(G125), .ZN(n1169) );
NAND2_X1 U961 ( .A1(n1262), .A2(n1028), .ZN(n1203) );
NAND3_X1 U962 ( .A1(n1226), .A2(n1104), .A3(G952), .ZN(n1028) );
NAND4_X1 U963 ( .A1(G953), .A2(G902), .A3(n1226), .A4(n1120), .ZN(n1262) );
INV_X1 U964 ( .A(G898), .ZN(n1120) );
NAND2_X1 U965 ( .A1(G237), .A2(G234), .ZN(n1226) );
INV_X1 U966 ( .A(n1213), .ZN(n1057) );
NAND2_X1 U967 ( .A1(n1263), .A2(n1059), .ZN(n1213) );
NAND2_X1 U968 ( .A1(G221), .A2(n1264), .ZN(n1059) );
XNOR2_X1 U969 ( .A(n1058), .B(KEYINPUT21), .ZN(n1263) );
XNOR2_X1 U970 ( .A(n1265), .B(G469), .ZN(n1058) );
NAND2_X1 U971 ( .A1(n1266), .A2(n1239), .ZN(n1265) );
XNOR2_X1 U972 ( .A(n1267), .B(n1158), .ZN(n1266) );
NAND2_X1 U973 ( .A1(n1268), .A2(n1269), .ZN(n1158) );
NAND3_X1 U974 ( .A1(n1270), .A2(n1104), .A3(n1271), .ZN(n1269) );
XNOR2_X1 U975 ( .A(G110), .B(G140), .ZN(n1271) );
NAND2_X1 U976 ( .A1(n1272), .A2(n1273), .ZN(n1268) );
NAND2_X1 U977 ( .A1(n1270), .A2(n1104), .ZN(n1273) );
XOR2_X1 U978 ( .A(KEYINPUT18), .B(G227), .Z(n1270) );
XNOR2_X1 U979 ( .A(n1274), .B(G110), .ZN(n1272) );
INV_X1 U980 ( .A(G140), .ZN(n1274) );
NOR2_X1 U981 ( .A1(KEYINPUT26), .A2(n1162), .ZN(n1267) );
XOR2_X1 U982 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U983 ( .A(n1275), .B(n1253), .Z(n1163) );
XNOR2_X1 U984 ( .A(n1276), .B(G104), .ZN(n1253) );
INV_X1 U985 ( .A(G107), .ZN(n1276) );
XNOR2_X1 U986 ( .A(n1277), .B(n1278), .ZN(n1275) );
INV_X1 U987 ( .A(n1102), .ZN(n1278) );
XNOR2_X1 U988 ( .A(n1279), .B(n1280), .ZN(n1102) );
XOR2_X1 U989 ( .A(G146), .B(n1281), .Z(n1280) );
NOR2_X1 U990 ( .A1(KEYINPUT15), .A2(n1282), .ZN(n1281) );
NAND2_X1 U991 ( .A1(KEYINPUT42), .A2(n1206), .ZN(n1279) );
NAND2_X1 U992 ( .A1(KEYINPUT14), .A2(n1221), .ZN(n1277) );
INV_X1 U993 ( .A(n1032), .ZN(n1197) );
NAND2_X1 U994 ( .A1(n1283), .A2(n1234), .ZN(n1032) );
XNOR2_X1 U995 ( .A(n1284), .B(n1285), .ZN(n1234) );
XOR2_X1 U996 ( .A(KEYINPUT60), .B(G478), .Z(n1285) );
NAND2_X1 U997 ( .A1(n1133), .A2(n1239), .ZN(n1284) );
XNOR2_X1 U998 ( .A(n1286), .B(n1287), .ZN(n1133) );
XOR2_X1 U999 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U1000 ( .A(G107), .B(n1290), .ZN(n1289) );
AND3_X1 U1001 ( .A1(G217), .A2(n1104), .A3(G234), .ZN(n1290) );
NAND2_X1 U1002 ( .A1(n1291), .A2(KEYINPUT34), .ZN(n1288) );
XNOR2_X1 U1003 ( .A(G122), .B(n1292), .ZN(n1291) );
NOR2_X1 U1004 ( .A1(G116), .A2(KEYINPUT7), .ZN(n1292) );
XNOR2_X1 U1005 ( .A(G128), .B(n1293), .ZN(n1286) );
XNOR2_X1 U1006 ( .A(n1206), .B(G134), .ZN(n1293) );
XNOR2_X1 U1007 ( .A(n1233), .B(KEYINPUT24), .ZN(n1283) );
XOR2_X1 U1008 ( .A(n1294), .B(n1090), .Z(n1233) );
NAND2_X1 U1009 ( .A1(n1239), .A2(n1136), .ZN(n1090) );
NAND2_X1 U1010 ( .A1(n1295), .A2(n1296), .ZN(n1136) );
NAND2_X1 U1011 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U1012 ( .A(KEYINPUT62), .B(n1299), .Z(n1295) );
NOR2_X1 U1013 ( .A1(n1298), .A2(n1297), .ZN(n1299) );
XOR2_X1 U1014 ( .A(n1300), .B(n1301), .Z(n1297) );
XOR2_X1 U1015 ( .A(G131), .B(n1302), .Z(n1301) );
XNOR2_X1 U1016 ( .A(G146), .B(n1206), .ZN(n1302) );
XOR2_X1 U1017 ( .A(n1303), .B(n1099), .Z(n1300) );
XOR2_X1 U1018 ( .A(G125), .B(G140), .Z(n1099) );
NAND2_X1 U1019 ( .A1(n1304), .A2(G214), .ZN(n1303) );
AND2_X1 U1020 ( .A1(n1305), .A2(n1306), .ZN(n1298) );
NAND2_X1 U1021 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XNOR2_X1 U1022 ( .A(n1309), .B(n1310), .ZN(n1308) );
INV_X1 U1023 ( .A(G113), .ZN(n1309) );
XNOR2_X1 U1024 ( .A(G104), .B(KEYINPUT1), .ZN(n1307) );
NAND2_X1 U1025 ( .A1(n1311), .A2(G104), .ZN(n1305) );
XNOR2_X1 U1026 ( .A(G113), .B(n1310), .ZN(n1311) );
NOR2_X1 U1027 ( .A1(KEYINPUT57), .A2(G122), .ZN(n1310) );
NAND2_X1 U1028 ( .A1(KEYINPUT45), .A2(n1138), .ZN(n1294) );
INV_X1 U1029 ( .A(G475), .ZN(n1138) );
NAND2_X1 U1030 ( .A1(n1218), .A2(n1230), .ZN(n1060) );
NAND2_X1 U1031 ( .A1(n1312), .A2(n1087), .ZN(n1230) );
NAND2_X1 U1032 ( .A1(n1075), .A2(n1076), .ZN(n1087) );
NAND2_X1 U1033 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
INV_X1 U1034 ( .A(n1075), .ZN(n1314) );
NOR2_X1 U1035 ( .A1(n1315), .A2(G902), .ZN(n1075) );
INV_X1 U1036 ( .A(n1126), .ZN(n1315) );
XNOR2_X1 U1037 ( .A(n1316), .B(n1317), .ZN(n1126) );
XOR2_X1 U1038 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1039 ( .A(n1282), .B(G119), .ZN(n1319) );
XOR2_X1 U1040 ( .A(KEYINPUT32), .B(G137), .Z(n1318) );
XOR2_X1 U1041 ( .A(n1320), .B(n1321), .Z(n1316) );
AND3_X1 U1042 ( .A1(G221), .A2(n1104), .A3(G234), .ZN(n1321) );
INV_X1 U1043 ( .A(G953), .ZN(n1104) );
XNOR2_X1 U1044 ( .A(n1322), .B(n1248), .ZN(n1320) );
INV_X1 U1045 ( .A(G110), .ZN(n1248) );
NAND2_X1 U1046 ( .A1(n1323), .A2(KEYINPUT30), .ZN(n1322) );
XOR2_X1 U1047 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U1048 ( .A(KEYINPUT19), .B(G146), .Z(n1325) );
XNOR2_X1 U1049 ( .A(G140), .B(n1326), .ZN(n1324) );
NOR2_X1 U1050 ( .A1(KEYINPUT6), .A2(n1327), .ZN(n1326) );
XNOR2_X1 U1051 ( .A(G125), .B(KEYINPUT8), .ZN(n1327) );
XOR2_X1 U1052 ( .A(n1076), .B(KEYINPUT52), .Z(n1313) );
NAND2_X1 U1053 ( .A1(G217), .A2(n1264), .ZN(n1076) );
NAND2_X1 U1054 ( .A1(G234), .A2(n1239), .ZN(n1264) );
NAND3_X1 U1055 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1218) );
OR2_X1 U1056 ( .A1(n1084), .A2(KEYINPUT61), .ZN(n1330) );
NAND3_X1 U1057 ( .A1(KEYINPUT61), .A2(n1331), .A3(n1086), .ZN(n1329) );
OR2_X1 U1058 ( .A1(n1086), .A2(n1331), .ZN(n1328) );
NOR2_X1 U1059 ( .A1(n1082), .A2(KEYINPUT39), .ZN(n1331) );
INV_X1 U1060 ( .A(n1084), .ZN(n1082) );
NAND2_X1 U1061 ( .A1(n1332), .A2(n1239), .ZN(n1084) );
INV_X1 U1062 ( .A(G902), .ZN(n1239) );
XOR2_X1 U1063 ( .A(n1333), .B(n1152), .Z(n1332) );
XNOR2_X1 U1064 ( .A(n1334), .B(n1221), .ZN(n1152) );
INV_X1 U1065 ( .A(G101), .ZN(n1221) );
NAND2_X1 U1066 ( .A1(n1304), .A2(G210), .ZN(n1334) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1304) );
NAND2_X1 U1068 ( .A1(n1335), .A2(KEYINPUT2), .ZN(n1333) );
XNOR2_X1 U1069 ( .A(n1148), .B(n1336), .ZN(n1335) );
XOR2_X1 U1070 ( .A(KEYINPUT16), .B(n1337), .Z(n1336) );
NOR2_X1 U1071 ( .A1(KEYINPUT36), .A2(n1149), .ZN(n1337) );
XOR2_X1 U1072 ( .A(n1243), .B(n1338), .Z(n1149) );
XOR2_X1 U1073 ( .A(G116), .B(n1339), .Z(n1338) );
NOR2_X1 U1074 ( .A1(G119), .A2(KEYINPUT51), .ZN(n1339) );
XNOR2_X1 U1075 ( .A(G113), .B(KEYINPUT56), .ZN(n1243) );
XNOR2_X1 U1076 ( .A(n1261), .B(n1164), .ZN(n1148) );
XNOR2_X1 U1077 ( .A(n1340), .B(n1103), .ZN(n1164) );
XOR2_X1 U1078 ( .A(G131), .B(G137), .Z(n1103) );
NAND2_X1 U1079 ( .A1(KEYINPUT50), .A2(n1101), .ZN(n1340) );
INV_X1 U1080 ( .A(G134), .ZN(n1101) );
NAND3_X1 U1081 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1261) );
NAND2_X1 U1082 ( .A1(n1344), .A2(n1282), .ZN(n1343) );
INV_X1 U1083 ( .A(G128), .ZN(n1282) );
NAND3_X1 U1084 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1344) );
NAND2_X1 U1085 ( .A1(KEYINPUT20), .A2(KEYINPUT17), .ZN(n1347) );
NAND2_X1 U1086 ( .A1(KEYINPUT4), .A2(n1348), .ZN(n1346) );
NAND2_X1 U1087 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1088 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NAND2_X1 U1089 ( .A1(n1349), .A2(n1353), .ZN(n1345) );
INV_X1 U1090 ( .A(KEYINPUT4), .ZN(n1353) );
NAND4_X1 U1091 ( .A1(n1349), .A2(G128), .A3(KEYINPUT20), .A4(n1351), .ZN(n1342) );
INV_X1 U1092 ( .A(KEYINPUT17), .ZN(n1351) );
NAND2_X1 U1093 ( .A1(KEYINPUT17), .A2(n1354), .ZN(n1341) );
NAND2_X1 U1094 ( .A1(n1349), .A2(n1355), .ZN(n1354) );
NAND2_X1 U1095 ( .A1(G128), .A2(n1352), .ZN(n1355) );
INV_X1 U1096 ( .A(KEYINPUT20), .ZN(n1352) );
XOR2_X1 U1097 ( .A(n1356), .B(G146), .Z(n1349) );
NAND2_X1 U1098 ( .A1(KEYINPUT5), .A2(n1206), .ZN(n1356) );
INV_X1 U1099 ( .A(G143), .ZN(n1206) );
INV_X1 U1100 ( .A(G472), .ZN(n1086) );
endmodule


