//Key = 1101001110111110101100010000001100110011111110100110101111101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373;

XOR2_X1 U743 ( .A(n1038), .B(n1039), .Z(G9) );
NOR2_X1 U744 ( .A1(G107), .A2(KEYINPUT5), .ZN(n1039) );
NOR2_X1 U745 ( .A1(n1040), .A2(n1041), .ZN(G75) );
NOR3_X1 U746 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
INV_X1 U747 ( .A(n1045), .ZN(n1043) );
NAND3_X1 U748 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1042) );
NAND3_X1 U749 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND3_X1 U750 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1049) );
XOR2_X1 U751 ( .A(KEYINPUT41), .B(n1055), .Z(n1054) );
AND2_X1 U752 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND3_X1 U753 ( .A1(n1058), .A2(n1059), .A3(n1057), .ZN(n1053) );
NAND3_X1 U754 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1052) );
NAND3_X1 U755 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NAND2_X1 U756 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U757 ( .A1(n1068), .A2(n1069), .ZN(n1063) );
OR2_X1 U758 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND3_X1 U759 ( .A1(n1060), .A2(n1072), .A3(n1057), .ZN(n1046) );
AND3_X1 U760 ( .A1(n1068), .A2(n1067), .A3(n1062), .ZN(n1057) );
INV_X1 U761 ( .A(n1073), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND2_X1 U763 ( .A1(n1076), .A2(n1051), .ZN(n1075) );
NOR3_X1 U764 ( .A1(n1044), .A2(G952), .A3(n1077), .ZN(n1040) );
INV_X1 U765 ( .A(n1047), .ZN(n1077) );
NAND4_X1 U766 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1047) );
NOR3_X1 U767 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
XOR2_X1 U768 ( .A(n1085), .B(KEYINPUT60), .Z(n1084) );
NOR2_X1 U769 ( .A1(n1086), .A2(n1087), .ZN(n1083) );
XOR2_X1 U770 ( .A(n1088), .B(KEYINPUT31), .Z(n1080) );
NAND3_X1 U771 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
NOR3_X1 U772 ( .A1(n1076), .A2(n1059), .A3(n1092), .ZN(n1091) );
XNOR2_X1 U773 ( .A(KEYINPUT19), .B(n1058), .ZN(n1089) );
XNOR2_X1 U774 ( .A(n1093), .B(G472), .ZN(n1079) );
XOR2_X1 U775 ( .A(n1094), .B(n1095), .Z(n1078) );
XOR2_X1 U776 ( .A(KEYINPUT3), .B(n1096), .Z(n1095) );
NAND2_X1 U777 ( .A1(KEYINPUT8), .A2(n1097), .ZN(n1094) );
XOR2_X1 U778 ( .A(n1098), .B(n1099), .Z(G72) );
NAND2_X1 U779 ( .A1(G953), .A2(n1100), .ZN(n1099) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1100) );
NAND4_X1 U781 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1098) );
NAND3_X1 U782 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
INV_X1 U783 ( .A(KEYINPUT53), .ZN(n1106) );
OR2_X1 U784 ( .A1(n1107), .A2(n1105), .ZN(n1103) );
NOR2_X1 U785 ( .A1(KEYINPUT25), .A2(n1108), .ZN(n1105) );
AND2_X1 U786 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NAND2_X1 U787 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U788 ( .A(KEYINPUT28), .B(n1113), .Z(n1111) );
XOR2_X1 U789 ( .A(KEYINPUT11), .B(n1114), .Z(n1109) );
NOR2_X1 U790 ( .A1(n1113), .A2(n1112), .ZN(n1114) );
XNOR2_X1 U791 ( .A(n1115), .B(n1116), .ZN(n1112) );
XNOR2_X1 U792 ( .A(n1117), .B(n1118), .ZN(n1116) );
XNOR2_X1 U793 ( .A(KEYINPUT54), .B(n1119), .ZN(n1118) );
INV_X1 U794 ( .A(G137), .ZN(n1119) );
XNOR2_X1 U795 ( .A(n1120), .B(n1121), .ZN(n1115) );
INV_X1 U796 ( .A(G131), .ZN(n1121) );
NAND2_X1 U797 ( .A1(KEYINPUT52), .A2(n1122), .ZN(n1120) );
NAND2_X1 U798 ( .A1(G953), .A2(n1123), .ZN(n1102) );
NAND2_X1 U799 ( .A1(KEYINPUT53), .A2(n1108), .ZN(n1101) );
NAND2_X1 U800 ( .A1(n1124), .A2(n1125), .ZN(n1108) );
XOR2_X1 U801 ( .A(n1126), .B(n1127), .Z(G69) );
XOR2_X1 U802 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U804 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR2_X1 U805 ( .A1(G898), .A2(n1124), .ZN(n1130) );
NAND2_X1 U806 ( .A1(n1124), .A2(n1134), .ZN(n1128) );
NAND2_X1 U807 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U808 ( .A(KEYINPUT40), .B(n1137), .Z(n1136) );
INV_X1 U809 ( .A(n1138), .ZN(n1135) );
NAND2_X1 U810 ( .A1(G953), .A2(n1139), .ZN(n1126) );
NAND2_X1 U811 ( .A1(G898), .A2(G224), .ZN(n1139) );
NOR2_X1 U812 ( .A1(n1140), .A2(n1141), .ZN(G66) );
XOR2_X1 U813 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND3_X1 U814 ( .A1(n1144), .A2(n1145), .A3(KEYINPUT16), .ZN(n1142) );
NOR2_X1 U815 ( .A1(n1140), .A2(n1146), .ZN(G63) );
XOR2_X1 U816 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U817 ( .A1(n1087), .A2(n1149), .ZN(n1148) );
NOR2_X1 U818 ( .A1(n1140), .A2(n1150), .ZN(G60) );
NOR3_X1 U819 ( .A1(n1096), .A2(n1151), .A3(n1152), .ZN(n1150) );
NOR3_X1 U820 ( .A1(n1153), .A2(n1097), .A3(n1149), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1151) );
NOR2_X1 U822 ( .A1(n1045), .A2(n1097), .ZN(n1155) );
XNOR2_X1 U823 ( .A(G104), .B(n1156), .ZN(G6) );
NOR2_X1 U824 ( .A1(n1140), .A2(n1157), .ZN(G57) );
XOR2_X1 U825 ( .A(n1158), .B(n1159), .Z(n1157) );
XNOR2_X1 U826 ( .A(n1160), .B(n1161), .ZN(n1159) );
XOR2_X1 U827 ( .A(n1162), .B(n1163), .Z(n1158) );
NOR2_X1 U828 ( .A1(n1164), .A2(n1149), .ZN(n1163) );
NAND2_X1 U829 ( .A1(KEYINPUT55), .A2(n1165), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1140), .A2(n1166), .ZN(G54) );
XOR2_X1 U831 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U832 ( .A(n1169), .B(n1122), .ZN(n1168) );
INV_X1 U833 ( .A(n1170), .ZN(n1122) );
XOR2_X1 U834 ( .A(KEYINPUT17), .B(n1171), .Z(n1167) );
AND2_X1 U835 ( .A1(G469), .A2(n1144), .ZN(n1171) );
NOR2_X1 U836 ( .A1(n1140), .A2(n1172), .ZN(G51) );
XOR2_X1 U837 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U838 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U839 ( .A1(n1177), .A2(n1149), .ZN(n1176) );
INV_X1 U840 ( .A(n1144), .ZN(n1149) );
NOR2_X1 U841 ( .A1(n1178), .A2(n1045), .ZN(n1144) );
NOR3_X1 U842 ( .A1(n1138), .A2(n1137), .A3(n1125), .ZN(n1045) );
NAND4_X1 U843 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1125) );
AND4_X1 U844 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
NOR2_X1 U845 ( .A1(n1187), .A2(n1188), .ZN(n1181) );
NOR2_X1 U846 ( .A1(n1074), .A2(n1189), .ZN(n1188) );
AND3_X1 U847 ( .A1(n1066), .A2(n1071), .A3(n1190), .ZN(n1187) );
NAND4_X1 U848 ( .A1(n1191), .A2(n1156), .A3(n1192), .A4(n1193), .ZN(n1138) );
AND4_X1 U849 ( .A1(n1038), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1193) );
NAND3_X1 U850 ( .A1(n1197), .A2(n1068), .A3(n1070), .ZN(n1038) );
NAND4_X1 U851 ( .A1(n1066), .A2(n1071), .A3(n1198), .A4(n1199), .ZN(n1192) );
NAND2_X1 U852 ( .A1(KEYINPUT46), .A2(n1200), .ZN(n1199) );
NAND2_X1 U853 ( .A1(n1201), .A2(n1202), .ZN(n1198) );
INV_X1 U854 ( .A(KEYINPUT46), .ZN(n1202) );
NAND3_X1 U855 ( .A1(n1074), .A2(n1203), .A3(n1060), .ZN(n1201) );
NAND3_X1 U856 ( .A1(n1197), .A2(n1068), .A3(n1071), .ZN(n1156) );
NAND3_X1 U857 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1191) );
XOR2_X1 U858 ( .A(n1067), .B(KEYINPUT33), .Z(n1204) );
NOR2_X1 U859 ( .A1(KEYINPUT26), .A2(n1207), .ZN(n1175) );
XNOR2_X1 U860 ( .A(n1208), .B(n1209), .ZN(n1207) );
NAND2_X1 U861 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U862 ( .A(n1212), .B(KEYINPUT20), .Z(n1210) );
NOR2_X1 U863 ( .A1(n1124), .A2(G952), .ZN(n1140) );
XNOR2_X1 U864 ( .A(G146), .B(n1186), .ZN(G48) );
NAND4_X1 U865 ( .A1(n1205), .A2(n1213), .A3(n1071), .A4(n1214), .ZN(n1186) );
XOR2_X1 U866 ( .A(n1185), .B(n1215), .Z(G45) );
NOR2_X1 U867 ( .A1(G143), .A2(KEYINPUT29), .ZN(n1215) );
NAND3_X1 U868 ( .A1(n1066), .A2(n1213), .A3(n1216), .ZN(n1185) );
NOR3_X1 U869 ( .A1(n1074), .A2(n1217), .A3(n1218), .ZN(n1216) );
INV_X1 U870 ( .A(n1214), .ZN(n1074) );
XNOR2_X1 U871 ( .A(G140), .B(n1179), .ZN(G42) );
NAND4_X1 U872 ( .A1(n1190), .A2(n1071), .A3(n1219), .A4(n1220), .ZN(n1179) );
XNOR2_X1 U873 ( .A(n1221), .B(n1180), .ZN(G39) );
OR2_X1 U874 ( .A1(n1222), .A2(n1223), .ZN(n1180) );
XNOR2_X1 U875 ( .A(G137), .B(KEYINPUT13), .ZN(n1221) );
XNOR2_X1 U876 ( .A(G134), .B(n1184), .ZN(G36) );
NAND3_X1 U877 ( .A1(n1190), .A2(n1070), .A3(n1066), .ZN(n1184) );
XNOR2_X1 U878 ( .A(G131), .B(n1224), .ZN(G33) );
NAND3_X1 U879 ( .A1(n1190), .A2(n1071), .A3(n1225), .ZN(n1224) );
XNOR2_X1 U880 ( .A(n1066), .B(KEYINPUT62), .ZN(n1225) );
INV_X1 U881 ( .A(n1223), .ZN(n1190) );
NAND3_X1 U882 ( .A1(n1213), .A2(n1050), .A3(n1051), .ZN(n1223) );
XNOR2_X1 U883 ( .A(G128), .B(n1226), .ZN(G30) );
NAND2_X1 U884 ( .A1(n1227), .A2(n1214), .ZN(n1226) );
XOR2_X1 U885 ( .A(n1189), .B(KEYINPUT34), .Z(n1227) );
NAND3_X1 U886 ( .A1(n1213), .A2(n1070), .A3(n1205), .ZN(n1189) );
AND2_X1 U887 ( .A1(n1056), .A2(n1228), .ZN(n1213) );
XOR2_X1 U888 ( .A(n1196), .B(n1229), .Z(G3) );
NAND2_X1 U889 ( .A1(KEYINPUT42), .A2(G101), .ZN(n1229) );
NAND3_X1 U890 ( .A1(n1197), .A2(n1067), .A3(n1066), .ZN(n1196) );
INV_X1 U891 ( .A(n1230), .ZN(n1197) );
XNOR2_X1 U892 ( .A(G125), .B(n1183), .ZN(G27) );
NAND4_X1 U893 ( .A1(n1219), .A2(n1071), .A3(n1060), .A4(n1231), .ZN(n1183) );
AND3_X1 U894 ( .A1(n1220), .A2(n1228), .A3(n1214), .ZN(n1231) );
NAND2_X1 U895 ( .A1(n1073), .A2(n1232), .ZN(n1228) );
NAND4_X1 U896 ( .A1(G902), .A2(G953), .A3(n1233), .A4(n1123), .ZN(n1232) );
INV_X1 U897 ( .A(G900), .ZN(n1123) );
XOR2_X1 U898 ( .A(n1195), .B(n1234), .Z(G24) );
XOR2_X1 U899 ( .A(KEYINPUT10), .B(G122), .Z(n1234) );
NAND4_X1 U900 ( .A1(n1206), .A2(n1068), .A3(n1235), .A4(n1236), .ZN(n1195) );
NOR2_X1 U901 ( .A1(n1237), .A2(n1219), .ZN(n1068) );
XOR2_X1 U902 ( .A(G119), .B(n1238), .Z(G21) );
NOR2_X1 U903 ( .A1(n1222), .A2(n1200), .ZN(n1238) );
NAND2_X1 U904 ( .A1(n1205), .A2(n1067), .ZN(n1222) );
AND2_X1 U905 ( .A1(n1219), .A2(n1237), .ZN(n1205) );
XNOR2_X1 U906 ( .A(G116), .B(n1194), .ZN(G18) );
NAND3_X1 U907 ( .A1(n1066), .A2(n1070), .A3(n1206), .ZN(n1194) );
NAND2_X1 U908 ( .A1(n1239), .A2(n1240), .ZN(G15) );
NAND2_X1 U909 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND2_X1 U910 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
OR2_X1 U911 ( .A1(n1245), .A2(KEYINPUT63), .ZN(n1244) );
NAND3_X1 U912 ( .A1(n1246), .A2(n1247), .A3(KEYINPUT63), .ZN(n1239) );
NAND2_X1 U913 ( .A1(n1243), .A2(n1245), .ZN(n1247) );
INV_X1 U914 ( .A(KEYINPUT6), .ZN(n1245) );
NAND2_X1 U915 ( .A1(KEYINPUT6), .A2(n1248), .ZN(n1246) );
NAND2_X1 U916 ( .A1(G113), .A2(n1243), .ZN(n1248) );
NAND3_X1 U917 ( .A1(n1066), .A2(n1071), .A3(n1206), .ZN(n1243) );
INV_X1 U918 ( .A(n1200), .ZN(n1206) );
NAND3_X1 U919 ( .A1(n1214), .A2(n1203), .A3(n1060), .ZN(n1200) );
AND2_X1 U920 ( .A1(n1249), .A2(n1058), .ZN(n1060) );
XNOR2_X1 U921 ( .A(n1059), .B(KEYINPUT4), .ZN(n1249) );
NOR2_X1 U922 ( .A1(n1236), .A2(n1218), .ZN(n1071) );
NOR2_X1 U923 ( .A1(n1219), .A2(n1220), .ZN(n1066) );
XOR2_X1 U924 ( .A(G110), .B(n1137), .Z(G12) );
NOR2_X1 U925 ( .A1(n1064), .A2(n1230), .ZN(n1137) );
NAND3_X1 U926 ( .A1(n1056), .A2(n1203), .A3(n1214), .ZN(n1230) );
NOR2_X1 U927 ( .A1(n1076), .A2(n1051), .ZN(n1214) );
AND2_X1 U928 ( .A1(n1250), .A2(n1090), .ZN(n1051) );
NAND2_X1 U929 ( .A1(n1251), .A2(n1177), .ZN(n1090) );
XOR2_X1 U930 ( .A(KEYINPUT43), .B(n1092), .Z(n1250) );
NOR2_X1 U931 ( .A1(n1177), .A2(n1251), .ZN(n1092) );
AND2_X1 U932 ( .A1(n1252), .A2(n1178), .ZN(n1251) );
XOR2_X1 U933 ( .A(n1173), .B(n1253), .Z(n1252) );
XOR2_X1 U934 ( .A(n1254), .B(n1255), .Z(n1253) );
NAND2_X1 U935 ( .A1(KEYINPUT30), .A2(n1208), .ZN(n1255) );
AND2_X1 U936 ( .A1(G224), .A2(n1124), .ZN(n1208) );
NAND2_X1 U937 ( .A1(n1211), .A2(n1212), .ZN(n1254) );
NAND2_X1 U938 ( .A1(n1256), .A2(n1160), .ZN(n1212) );
XNOR2_X1 U939 ( .A(KEYINPUT9), .B(G125), .ZN(n1256) );
NAND2_X1 U940 ( .A1(n1257), .A2(n1258), .ZN(n1211) );
XOR2_X1 U941 ( .A(KEYINPUT9), .B(G125), .Z(n1258) );
XNOR2_X1 U942 ( .A(n1132), .B(n1259), .ZN(n1173) );
NOR2_X1 U943 ( .A1(KEYINPUT45), .A2(n1133), .ZN(n1259) );
NAND2_X1 U944 ( .A1(n1260), .A2(n1261), .ZN(n1133) );
NAND2_X1 U945 ( .A1(KEYINPUT21), .A2(n1262), .ZN(n1261) );
NAND2_X1 U946 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
NAND2_X1 U947 ( .A1(n1265), .A2(n1242), .ZN(n1264) );
NAND2_X1 U948 ( .A1(n1266), .A2(n1267), .ZN(n1260) );
INV_X1 U949 ( .A(KEYINPUT21), .ZN(n1267) );
XNOR2_X1 U950 ( .A(n1242), .B(n1268), .ZN(n1266) );
XOR2_X1 U951 ( .A(n1269), .B(n1270), .Z(n1132) );
XNOR2_X1 U952 ( .A(G110), .B(n1271), .ZN(n1270) );
XOR2_X1 U953 ( .A(n1272), .B(n1273), .Z(n1269) );
NAND2_X1 U954 ( .A1(KEYINPUT18), .A2(G101), .ZN(n1272) );
NAND2_X1 U955 ( .A1(G210), .A2(n1274), .ZN(n1177) );
INV_X1 U956 ( .A(n1050), .ZN(n1076) );
NAND2_X1 U957 ( .A1(G214), .A2(n1274), .ZN(n1050) );
NAND2_X1 U958 ( .A1(n1275), .A2(n1178), .ZN(n1274) );
NAND2_X1 U959 ( .A1(n1276), .A2(n1073), .ZN(n1203) );
NAND3_X1 U960 ( .A1(n1277), .A2(n1233), .A3(G952), .ZN(n1073) );
INV_X1 U961 ( .A(n1044), .ZN(n1277) );
XOR2_X1 U962 ( .A(G953), .B(KEYINPUT51), .Z(n1044) );
NAND4_X1 U963 ( .A1(G902), .A2(G953), .A3(n1233), .A4(n1278), .ZN(n1276) );
INV_X1 U964 ( .A(G898), .ZN(n1278) );
NAND2_X1 U965 ( .A1(G237), .A2(G234), .ZN(n1233) );
NOR2_X1 U966 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
AND2_X1 U967 ( .A1(G221), .A2(n1279), .ZN(n1059) );
XOR2_X1 U968 ( .A(n1280), .B(G469), .Z(n1058) );
NAND2_X1 U969 ( .A1(n1281), .A2(n1178), .ZN(n1280) );
XNOR2_X1 U970 ( .A(n1282), .B(n1283), .ZN(n1281) );
INV_X1 U971 ( .A(n1169), .ZN(n1283) );
XNOR2_X1 U972 ( .A(n1284), .B(n1285), .ZN(n1169) );
XOR2_X1 U973 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U974 ( .A(n1288), .B(n1289), .Z(n1287) );
NAND2_X1 U975 ( .A1(G227), .A2(n1124), .ZN(n1289) );
NAND3_X1 U976 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1288) );
NAND2_X1 U977 ( .A1(G104), .A2(n1271), .ZN(n1292) );
INV_X1 U978 ( .A(G107), .ZN(n1271) );
NAND2_X1 U979 ( .A1(KEYINPUT24), .A2(n1293), .ZN(n1291) );
NAND2_X1 U980 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XNOR2_X1 U981 ( .A(KEYINPUT38), .B(G107), .ZN(n1294) );
NAND2_X1 U982 ( .A1(n1296), .A2(n1297), .ZN(n1290) );
INV_X1 U983 ( .A(KEYINPUT24), .ZN(n1297) );
NAND2_X1 U984 ( .A1(n1298), .A2(n1299), .ZN(n1296) );
OR2_X1 U985 ( .A1(G107), .A2(KEYINPUT38), .ZN(n1299) );
NAND3_X1 U986 ( .A1(G107), .A2(n1295), .A3(KEYINPUT38), .ZN(n1298) );
XNOR2_X1 U987 ( .A(G110), .B(n1300), .ZN(n1284) );
XOR2_X1 U988 ( .A(KEYINPUT57), .B(G140), .Z(n1300) );
NOR2_X1 U989 ( .A1(KEYINPUT37), .A2(n1170), .ZN(n1282) );
XNOR2_X1 U990 ( .A(n1301), .B(n1302), .ZN(n1170) );
NAND3_X1 U991 ( .A1(n1220), .A2(n1067), .A3(n1219), .ZN(n1064) );
XNOR2_X1 U992 ( .A(n1082), .B(KEYINPUT0), .ZN(n1219) );
XNOR2_X1 U993 ( .A(n1303), .B(n1145), .ZN(n1082) );
AND2_X1 U994 ( .A1(G217), .A2(n1279), .ZN(n1145) );
NAND2_X1 U995 ( .A1(G234), .A2(n1178), .ZN(n1279) );
NAND2_X1 U996 ( .A1(n1143), .A2(n1178), .ZN(n1303) );
XOR2_X1 U997 ( .A(n1304), .B(n1305), .Z(n1143) );
NOR3_X1 U998 ( .A1(n1306), .A2(KEYINPUT15), .A3(n1307), .ZN(n1305) );
INV_X1 U999 ( .A(G221), .ZN(n1306) );
XNOR2_X1 U1000 ( .A(G137), .B(n1308), .ZN(n1304) );
NOR2_X1 U1001 ( .A1(KEYINPUT48), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1002 ( .A(n1113), .B(n1310), .Z(n1309) );
XNOR2_X1 U1003 ( .A(G146), .B(n1311), .ZN(n1310) );
NAND2_X1 U1004 ( .A1(KEYINPUT39), .A2(n1312), .ZN(n1311) );
XOR2_X1 U1005 ( .A(G110), .B(n1313), .Z(n1312) );
XNOR2_X1 U1006 ( .A(n1302), .B(G119), .ZN(n1313) );
NAND2_X1 U1007 ( .A1(n1314), .A2(n1315), .ZN(n1067) );
OR3_X1 U1008 ( .A1(n1236), .A2(n1235), .A3(KEYINPUT36), .ZN(n1315) );
NAND2_X1 U1009 ( .A1(KEYINPUT36), .A2(n1070), .ZN(n1314) );
NOR2_X1 U1010 ( .A1(n1235), .A2(n1217), .ZN(n1070) );
INV_X1 U1011 ( .A(n1236), .ZN(n1217) );
NAND2_X1 U1012 ( .A1(n1085), .A2(n1316), .ZN(n1236) );
OR2_X1 U1013 ( .A1(n1087), .A2(n1086), .ZN(n1316) );
NAND2_X1 U1014 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
INV_X1 U1015 ( .A(G478), .ZN(n1087) );
NOR2_X1 U1016 ( .A1(n1147), .A2(G902), .ZN(n1086) );
XOR2_X1 U1017 ( .A(n1317), .B(n1318), .Z(n1147) );
XOR2_X1 U1018 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1019 ( .A(n1321), .B(n1322), .ZN(n1320) );
NOR3_X1 U1020 ( .A1(n1323), .A2(KEYINPUT22), .A3(n1307), .ZN(n1322) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1124), .ZN(n1307) );
INV_X1 U1022 ( .A(G217), .ZN(n1323) );
NAND2_X1 U1023 ( .A1(n1324), .A2(KEYINPUT44), .ZN(n1321) );
XNOR2_X1 U1024 ( .A(G116), .B(G122), .ZN(n1324) );
XNOR2_X1 U1025 ( .A(G107), .B(n1325), .ZN(n1317) );
XNOR2_X1 U1026 ( .A(n1117), .B(G128), .ZN(n1325) );
INV_X1 U1027 ( .A(G134), .ZN(n1117) );
INV_X1 U1028 ( .A(n1218), .ZN(n1235) );
XOR2_X1 U1029 ( .A(n1096), .B(n1097), .Z(n1218) );
INV_X1 U1030 ( .A(G475), .ZN(n1097) );
NOR2_X1 U1031 ( .A1(n1154), .A2(G902), .ZN(n1096) );
INV_X1 U1032 ( .A(n1153), .ZN(n1154) );
NAND3_X1 U1033 ( .A1(n1326), .A2(n1327), .A3(n1328), .ZN(n1153) );
NAND2_X1 U1034 ( .A1(KEYINPUT47), .A2(n1329), .ZN(n1328) );
OR3_X1 U1035 ( .A1(n1329), .A2(KEYINPUT47), .A3(n1330), .ZN(n1327) );
NAND2_X1 U1036 ( .A1(n1330), .A2(n1331), .ZN(n1326) );
NAND2_X1 U1037 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
INV_X1 U1038 ( .A(KEYINPUT47), .ZN(n1333) );
XOR2_X1 U1039 ( .A(KEYINPUT12), .B(n1329), .Z(n1332) );
XNOR2_X1 U1040 ( .A(n1334), .B(n1335), .ZN(n1329) );
XNOR2_X1 U1041 ( .A(G131), .B(n1336), .ZN(n1335) );
NAND3_X1 U1042 ( .A1(n1275), .A2(n1124), .A3(n1337), .ZN(n1336) );
XOR2_X1 U1043 ( .A(KEYINPUT2), .B(G214), .Z(n1337) );
XNOR2_X1 U1044 ( .A(n1301), .B(n1113), .ZN(n1334) );
XOR2_X1 U1045 ( .A(G140), .B(G125), .Z(n1113) );
XNOR2_X1 U1046 ( .A(n1273), .B(n1338), .ZN(n1330) );
XNOR2_X1 U1047 ( .A(n1339), .B(KEYINPUT59), .ZN(n1338) );
NAND2_X1 U1048 ( .A1(KEYINPUT50), .A2(n1242), .ZN(n1339) );
XNOR2_X1 U1049 ( .A(G122), .B(n1295), .ZN(n1273) );
INV_X1 U1050 ( .A(G104), .ZN(n1295) );
INV_X1 U1051 ( .A(n1237), .ZN(n1220) );
NAND3_X1 U1052 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1237) );
NAND2_X1 U1053 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NAND3_X1 U1054 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1343) );
NAND2_X1 U1055 ( .A1(KEYINPUT23), .A2(n1348), .ZN(n1347) );
OR2_X1 U1056 ( .A1(G472), .A2(KEYINPUT58), .ZN(n1346) );
NAND2_X1 U1057 ( .A1(KEYINPUT58), .A2(n1349), .ZN(n1345) );
NAND2_X1 U1058 ( .A1(n1164), .A2(n1350), .ZN(n1349) );
NAND2_X1 U1059 ( .A1(KEYINPUT1), .A2(n1351), .ZN(n1350) );
NAND4_X1 U1060 ( .A1(n1093), .A2(n1164), .A3(KEYINPUT23), .A4(KEYINPUT1), .ZN(n1341) );
NAND2_X1 U1061 ( .A1(n1352), .A2(n1348), .ZN(n1340) );
INV_X1 U1062 ( .A(KEYINPUT1), .ZN(n1348) );
NAND2_X1 U1063 ( .A1(n1164), .A2(n1353), .ZN(n1352) );
NAND2_X1 U1064 ( .A1(n1093), .A2(n1351), .ZN(n1353) );
INV_X1 U1065 ( .A(KEYINPUT23), .ZN(n1351) );
INV_X1 U1066 ( .A(n1344), .ZN(n1093) );
NAND3_X1 U1067 ( .A1(n1354), .A2(n1355), .A3(n1178), .ZN(n1344) );
INV_X1 U1068 ( .A(G902), .ZN(n1178) );
NAND3_X1 U1069 ( .A1(n1356), .A2(n1357), .A3(n1358), .ZN(n1355) );
INV_X1 U1070 ( .A(KEYINPUT14), .ZN(n1358) );
XNOR2_X1 U1071 ( .A(G101), .B(n1359), .ZN(n1357) );
XOR2_X1 U1072 ( .A(n1360), .B(n1361), .Z(n1356) );
NAND2_X1 U1073 ( .A1(n1362), .A2(KEYINPUT14), .ZN(n1354) );
XOR2_X1 U1074 ( .A(n1361), .B(n1161), .Z(n1362) );
XOR2_X1 U1075 ( .A(n1359), .B(n1286), .Z(n1161) );
XNOR2_X1 U1076 ( .A(n1360), .B(G101), .ZN(n1286) );
NAND2_X1 U1077 ( .A1(n1363), .A2(n1364), .ZN(n1360) );
NAND2_X1 U1078 ( .A1(n1365), .A2(G131), .ZN(n1364) );
XOR2_X1 U1079 ( .A(KEYINPUT49), .B(n1366), .Z(n1363) );
NOR2_X1 U1080 ( .A1(G131), .A2(n1365), .ZN(n1366) );
XNOR2_X1 U1081 ( .A(G134), .B(n1367), .ZN(n1365) );
NOR2_X1 U1082 ( .A1(G137), .A2(KEYINPUT27), .ZN(n1367) );
NAND3_X1 U1083 ( .A1(n1275), .A2(n1124), .A3(G210), .ZN(n1359) );
INV_X1 U1084 ( .A(G953), .ZN(n1124) );
INV_X1 U1085 ( .A(G237), .ZN(n1275) );
XNOR2_X1 U1086 ( .A(n1368), .B(n1257), .ZN(n1361) );
INV_X1 U1087 ( .A(n1160), .ZN(n1257) );
XOR2_X1 U1088 ( .A(n1369), .B(n1370), .Z(n1160) );
INV_X1 U1089 ( .A(n1301), .ZN(n1370) );
XOR2_X1 U1090 ( .A(G146), .B(n1319), .Z(n1301) );
XOR2_X1 U1091 ( .A(G143), .B(KEYINPUT35), .Z(n1319) );
NAND2_X1 U1092 ( .A1(KEYINPUT61), .A2(n1302), .ZN(n1369) );
INV_X1 U1093 ( .A(G128), .ZN(n1302) );
XNOR2_X1 U1094 ( .A(n1165), .B(KEYINPUT7), .ZN(n1368) );
AND2_X1 U1095 ( .A1(n1371), .A2(n1372), .ZN(n1165) );
NAND2_X1 U1096 ( .A1(n1265), .A2(n1373), .ZN(n1372) );
XNOR2_X1 U1097 ( .A(KEYINPUT56), .B(n1242), .ZN(n1373) );
INV_X1 U1098 ( .A(G113), .ZN(n1242) );
INV_X1 U1099 ( .A(n1268), .ZN(n1265) );
XOR2_X1 U1100 ( .A(n1263), .B(KEYINPUT32), .Z(n1371) );
NAND2_X1 U1101 ( .A1(G113), .A2(n1268), .ZN(n1263) );
XOR2_X1 U1102 ( .A(G116), .B(G119), .Z(n1268) );
INV_X1 U1103 ( .A(G472), .ZN(n1164) );
endmodule


