//Key = 1011100011000011010111000011010110000010110000101111010100101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;

XOR2_X1 U726 ( .A(G107), .B(n998), .Z(G9) );
NAND4_X1 U727 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(G75) );
NAND4_X1 U728 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1001) );
NOR4_X1 U729 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
XOR2_X1 U730 ( .A(n1011), .B(KEYINPUT47), .Z(n1008) );
NAND2_X1 U731 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND2_X1 U732 ( .A1(G478), .A2(n1014), .ZN(n1013) );
XOR2_X1 U733 ( .A(n1015), .B(n1016), .Z(n1005) );
NAND2_X1 U734 ( .A1(KEYINPUT14), .A2(n1017), .ZN(n1015) );
XNOR2_X1 U735 ( .A(KEYINPUT28), .B(n1018), .ZN(n1017) );
XNOR2_X1 U736 ( .A(n1019), .B(KEYINPUT22), .ZN(n1004) );
XNOR2_X1 U737 ( .A(n1020), .B(n1021), .ZN(n1003) );
XNOR2_X1 U738 ( .A(n1022), .B(KEYINPUT10), .ZN(n1020) );
NAND2_X1 U739 ( .A1(n1023), .A2(n1024), .ZN(n1000) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND3_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
NAND3_X1 U742 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1028) );
NAND2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND3_X1 U744 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1031) );
XOR2_X1 U745 ( .A(n1038), .B(KEYINPUT3), .Z(n1037) );
XNOR2_X1 U746 ( .A(n1033), .B(KEYINPUT2), .ZN(n1035) );
NAND2_X1 U747 ( .A1(n1039), .A2(n1040), .ZN(n1030) );
NAND2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND4_X1 U749 ( .A1(n1043), .A2(n1044), .A3(n1039), .A4(n1045), .ZN(n1025) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U751 ( .A1(n1029), .A2(n1027), .ZN(n1046) );
NAND4_X1 U752 ( .A1(n1048), .A2(n1049), .A3(n1027), .A4(n1050), .ZN(n1044) );
NAND2_X1 U753 ( .A1(n1007), .A2(n1051), .ZN(n1043) );
INV_X1 U754 ( .A(n1052), .ZN(n1023) );
XOR2_X1 U755 ( .A(n1053), .B(n1054), .Z(G72) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U757 ( .A1(n1057), .A2(n1002), .ZN(n1055) );
AND2_X1 U758 ( .A1(G227), .A2(G900), .ZN(n1057) );
NAND2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1053) );
NAND2_X1 U760 ( .A1(G953), .A2(n1060), .ZN(n1059) );
XNOR2_X1 U761 ( .A(n1061), .B(n1062), .ZN(n1058) );
XNOR2_X1 U762 ( .A(n1063), .B(n1064), .ZN(n1062) );
NOR2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
XOR2_X1 U764 ( .A(KEYINPUT13), .B(n1067), .Z(n1066) );
NAND2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(G69) );
NAND2_X1 U766 ( .A1(n1070), .A2(n1002), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U768 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NAND2_X1 U769 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1075), .A2(n1074), .ZN(n1077) );
XNOR2_X1 U771 ( .A(n1078), .B(KEYINPUT59), .ZN(n1074) );
XOR2_X1 U772 ( .A(n1079), .B(KEYINPUT62), .Z(n1076) );
NAND2_X1 U773 ( .A1(n1080), .A2(G953), .ZN(n1068) );
XNOR2_X1 U774 ( .A(n1073), .B(n1081), .ZN(n1080) );
NOR2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U776 ( .A(n1079), .B(KEYINPUT57), .ZN(n1073) );
NAND2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
NAND2_X1 U778 ( .A1(G953), .A2(n1083), .ZN(n1085) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(n1084) );
NAND2_X1 U780 ( .A1(KEYINPUT21), .A2(n1088), .ZN(n1086) );
NOR2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(G66) );
NOR3_X1 U782 ( .A1(n1022), .A2(n1091), .A3(n1092), .ZN(n1090) );
AND3_X1 U783 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NOR2_X1 U784 ( .A1(n1096), .A2(n1093), .ZN(n1091) );
NOR2_X1 U785 ( .A1(n999), .A2(n1021), .ZN(n1096) );
NOR2_X1 U786 ( .A1(n1089), .A2(n1097), .ZN(G63) );
XOR2_X1 U787 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U788 ( .A1(n1100), .A2(KEYINPUT43), .ZN(n1099) );
NAND2_X1 U789 ( .A1(n1095), .A2(G478), .ZN(n1098) );
NOR2_X1 U790 ( .A1(n1089), .A2(n1101), .ZN(G60) );
NOR3_X1 U791 ( .A1(n1016), .A2(n1102), .A3(n1103), .ZN(n1101) );
AND3_X1 U792 ( .A1(n1104), .A2(G475), .A3(n1095), .ZN(n1103) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1104), .ZN(n1102) );
NOR2_X1 U794 ( .A1(n999), .A2(n1018), .ZN(n1105) );
XOR2_X1 U795 ( .A(G104), .B(n1106), .Z(G6) );
NOR2_X1 U796 ( .A1(n1089), .A2(n1107), .ZN(G57) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U799 ( .A(n1112), .B(n1113), .Z(n1108) );
NOR2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U803 ( .A1(n1120), .A2(n1121), .ZN(n1116) );
AND2_X1 U804 ( .A1(n1118), .A2(KEYINPUT16), .ZN(n1120) );
NOR4_X1 U805 ( .A1(KEYINPUT16), .A2(n1121), .A3(n1118), .A4(n1119), .ZN(n1114) );
INV_X1 U806 ( .A(KEYINPUT53), .ZN(n1119) );
NAND2_X1 U807 ( .A1(n1095), .A2(G472), .ZN(n1112) );
NOR2_X1 U808 ( .A1(n1089), .A2(n1122), .ZN(G54) );
XOR2_X1 U809 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U810 ( .A1(n1095), .A2(G469), .ZN(n1124) );
NAND2_X1 U811 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U813 ( .A(n1129), .B(KEYINPUT42), .Z(n1125) );
OR2_X1 U814 ( .A1(n1128), .A2(n1127), .ZN(n1129) );
AND2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
NAND2_X1 U816 ( .A1(n1132), .A2(n1118), .ZN(n1131) );
XOR2_X1 U817 ( .A(KEYINPUT49), .B(n1133), .Z(n1132) );
NAND2_X1 U818 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
XNOR2_X1 U819 ( .A(n1135), .B(n1063), .ZN(n1133) );
XNOR2_X1 U820 ( .A(n1136), .B(KEYINPUT50), .ZN(n1135) );
XOR2_X1 U821 ( .A(n1137), .B(KEYINPUT27), .Z(n1128) );
NOR2_X1 U822 ( .A1(n1089), .A2(n1138), .ZN(G51) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1139) );
NAND2_X1 U825 ( .A1(n1095), .A2(n1143), .ZN(n1141) );
NOR2_X1 U826 ( .A1(n1144), .A2(n999), .ZN(n1095) );
NOR3_X1 U827 ( .A1(n1078), .A2(n1056), .A3(n1145), .ZN(n999) );
INV_X1 U828 ( .A(n1075), .ZN(n1145) );
NOR4_X1 U829 ( .A1(n1146), .A2(n1106), .A3(n1147), .A4(n998), .ZN(n1075) );
NOR3_X1 U830 ( .A1(n1047), .A2(n1148), .A3(n1048), .ZN(n998) );
NOR3_X1 U831 ( .A1(n1047), .A2(n1148), .A3(n1049), .ZN(n1106) );
INV_X1 U832 ( .A(n1033), .ZN(n1047) );
NOR3_X1 U833 ( .A1(n1051), .A2(n1148), .A3(n1041), .ZN(n1146) );
NAND4_X1 U834 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1056) );
AND3_X1 U835 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
NAND2_X1 U836 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
NAND2_X1 U837 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U838 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U839 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U841 ( .A(n1034), .B(KEYINPUT60), .ZN(n1164) );
NAND2_X1 U842 ( .A1(n1039), .A2(n1166), .ZN(n1162) );
INV_X1 U843 ( .A(n1167), .ZN(n1158) );
NAND4_X1 U844 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1078) );
AND2_X1 U845 ( .A1(G953), .A2(n1172), .ZN(n1089) );
XOR2_X1 U846 ( .A(KEYINPUT46), .B(G952), .Z(n1172) );
XOR2_X1 U847 ( .A(G146), .B(n1173), .Z(G48) );
NOR3_X1 U848 ( .A1(n1174), .A2(n1175), .A3(n1049), .ZN(n1173) );
XNOR2_X1 U849 ( .A(n1165), .B(KEYINPUT7), .ZN(n1175) );
INV_X1 U850 ( .A(n1176), .ZN(n1174) );
XNOR2_X1 U851 ( .A(G143), .B(n1149), .ZN(G45) );
NAND4_X1 U852 ( .A1(n1176), .A2(n1166), .A3(n1177), .A4(n1178), .ZN(n1149) );
XNOR2_X1 U853 ( .A(G140), .B(n1150), .ZN(G42) );
OR4_X1 U854 ( .A1(n1009), .A2(n1179), .A3(n1049), .A4(n1042), .ZN(n1150) );
NAND3_X1 U855 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(G39) );
NAND4_X1 U856 ( .A1(n1019), .A2(n1183), .A3(n1165), .A4(n1184), .ZN(n1182) );
NOR3_X1 U857 ( .A1(n1185), .A2(n1009), .A3(n1186), .ZN(n1184) );
INV_X1 U858 ( .A(n1029), .ZN(n1186) );
NOR2_X1 U859 ( .A1(n1051), .A2(n1007), .ZN(n1029) );
XNOR2_X1 U860 ( .A(KEYINPUT1), .B(n1187), .ZN(n1185) );
NAND2_X1 U861 ( .A1(n1188), .A2(KEYINPUT26), .ZN(n1183) );
XNOR2_X1 U862 ( .A(G137), .B(KEYINPUT29), .ZN(n1188) );
OR2_X1 U863 ( .A1(G137), .A2(KEYINPUT26), .ZN(n1181) );
NAND3_X1 U864 ( .A1(G137), .A2(n1189), .A3(KEYINPUT26), .ZN(n1180) );
NAND3_X1 U865 ( .A1(n1190), .A2(n1191), .A3(n1167), .ZN(n1189) );
NOR3_X1 U866 ( .A1(n1192), .A2(n1051), .A3(n1009), .ZN(n1167) );
INV_X1 U867 ( .A(n1165), .ZN(n1192) );
OR2_X1 U868 ( .A1(n1156), .A2(KEYINPUT1), .ZN(n1191) );
NAND2_X1 U869 ( .A1(KEYINPUT1), .A2(n1193), .ZN(n1190) );
OR3_X1 U870 ( .A1(n1027), .A2(n1007), .A3(n1187), .ZN(n1193) );
INV_X1 U871 ( .A(n1050), .ZN(n1007) );
XOR2_X1 U872 ( .A(n1153), .B(n1194), .Z(G36) );
XNOR2_X1 U873 ( .A(G134), .B(KEYINPUT45), .ZN(n1194) );
NAND4_X1 U874 ( .A1(n1039), .A2(n1156), .A3(n1166), .A4(n1195), .ZN(n1153) );
INV_X1 U875 ( .A(n1179), .ZN(n1156) );
INV_X1 U876 ( .A(n1009), .ZN(n1039) );
XOR2_X1 U877 ( .A(G131), .B(n1196), .Z(G33) );
NOR4_X1 U878 ( .A1(n1049), .A2(n1041), .A3(n1179), .A4(n1197), .ZN(n1196) );
XNOR2_X1 U879 ( .A(KEYINPUT17), .B(n1009), .ZN(n1197) );
NAND2_X1 U880 ( .A1(n1036), .A2(n1038), .ZN(n1009) );
XNOR2_X1 U881 ( .A(G128), .B(n1155), .ZN(G30) );
NAND3_X1 U882 ( .A1(n1165), .A2(n1195), .A3(n1176), .ZN(n1155) );
NOR2_X1 U883 ( .A1(n1179), .A2(n1198), .ZN(n1176) );
NAND3_X1 U884 ( .A1(n1050), .A2(n1187), .A3(n1019), .ZN(n1179) );
XNOR2_X1 U885 ( .A(n1199), .B(n1200), .ZN(G3) );
NOR3_X1 U886 ( .A1(n1201), .A2(n1148), .A3(n1041), .ZN(n1200) );
INV_X1 U887 ( .A(n1166), .ZN(n1041) );
XNOR2_X1 U888 ( .A(KEYINPUT55), .B(n1051), .ZN(n1201) );
XNOR2_X1 U889 ( .A(G125), .B(n1154), .ZN(G27) );
NAND4_X1 U890 ( .A1(n1050), .A2(n1187), .A3(n1034), .A4(n1202), .ZN(n1154) );
NOR3_X1 U891 ( .A1(n1019), .A2(n1042), .A3(n1049), .ZN(n1202) );
NAND2_X1 U892 ( .A1(n1203), .A2(n1052), .ZN(n1187) );
NAND4_X1 U893 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1060), .ZN(n1203) );
INV_X1 U894 ( .A(G900), .ZN(n1060) );
XNOR2_X1 U895 ( .A(G122), .B(n1168), .ZN(G24) );
NAND4_X1 U896 ( .A1(n1205), .A2(n1033), .A3(n1177), .A4(n1178), .ZN(n1168) );
NOR2_X1 U897 ( .A1(n1010), .A2(n1206), .ZN(n1033) );
XNOR2_X1 U898 ( .A(G119), .B(n1169), .ZN(G21) );
NAND3_X1 U899 ( .A1(n1205), .A2(n1207), .A3(n1165), .ZN(n1169) );
NOR2_X1 U900 ( .A1(n1208), .A2(n1209), .ZN(n1165) );
INV_X1 U901 ( .A(n1206), .ZN(n1208) );
XOR2_X1 U902 ( .A(n1170), .B(n1210), .Z(G18) );
NAND2_X1 U903 ( .A1(KEYINPUT63), .A2(G116), .ZN(n1210) );
NAND3_X1 U904 ( .A1(n1166), .A2(n1195), .A3(n1205), .ZN(n1170) );
INV_X1 U905 ( .A(n1048), .ZN(n1195) );
NAND2_X1 U906 ( .A1(n1211), .A2(n1178), .ZN(n1048) );
INV_X1 U907 ( .A(n1177), .ZN(n1211) );
XNOR2_X1 U908 ( .A(G113), .B(n1171), .ZN(G15) );
NAND3_X1 U909 ( .A1(n1166), .A2(n1160), .A3(n1205), .ZN(n1171) );
AND4_X1 U910 ( .A1(n1027), .A2(n1034), .A3(n1212), .A4(n1050), .ZN(n1205) );
INV_X1 U911 ( .A(n1019), .ZN(n1027) );
INV_X1 U912 ( .A(n1049), .ZN(n1160) );
NAND2_X1 U913 ( .A1(n1213), .A2(n1177), .ZN(n1049) );
XOR2_X1 U914 ( .A(n1178), .B(KEYINPUT32), .Z(n1213) );
NOR2_X1 U915 ( .A1(n1206), .A2(n1209), .ZN(n1166) );
XNOR2_X1 U916 ( .A(n1214), .B(n1147), .ZN(G12) );
NOR3_X1 U917 ( .A1(n1042), .A2(n1148), .A3(n1051), .ZN(n1147) );
INV_X1 U918 ( .A(n1207), .ZN(n1051) );
NOR2_X1 U919 ( .A1(n1178), .A2(n1177), .ZN(n1207) );
XNOR2_X1 U920 ( .A(n1016), .B(n1018), .ZN(n1177) );
INV_X1 U921 ( .A(G475), .ZN(n1018) );
NOR2_X1 U922 ( .A1(n1104), .A2(G902), .ZN(n1016) );
XOR2_X1 U923 ( .A(n1215), .B(n1216), .Z(n1104) );
XNOR2_X1 U924 ( .A(n1217), .B(n1218), .ZN(n1216) );
INV_X1 U925 ( .A(n1061), .ZN(n1218) );
XOR2_X1 U926 ( .A(G125), .B(n1219), .Z(n1061) );
XOR2_X1 U927 ( .A(G140), .B(G131), .Z(n1219) );
XOR2_X1 U928 ( .A(n1220), .B(n1221), .Z(n1215) );
AND3_X1 U929 ( .A1(G214), .A2(n1222), .A3(n1223), .ZN(n1221) );
INV_X1 U930 ( .A(KEYINPUT25), .ZN(n1222) );
NAND2_X1 U931 ( .A1(n1224), .A2(n1225), .ZN(n1220) );
OR2_X1 U932 ( .A1(n1226), .A2(G104), .ZN(n1225) );
XOR2_X1 U933 ( .A(n1227), .B(KEYINPUT12), .Z(n1224) );
NAND2_X1 U934 ( .A1(G104), .A2(n1226), .ZN(n1227) );
XNOR2_X1 U935 ( .A(G113), .B(n1228), .ZN(n1226) );
INV_X1 U936 ( .A(G122), .ZN(n1228) );
NAND3_X1 U937 ( .A1(n1229), .A2(n1230), .A3(n1012), .ZN(n1178) );
OR2_X1 U938 ( .A1(n1014), .A2(G478), .ZN(n1012) );
OR2_X1 U939 ( .A1(G478), .A2(KEYINPUT0), .ZN(n1230) );
NAND3_X1 U940 ( .A1(G478), .A2(n1014), .A3(KEYINPUT0), .ZN(n1229) );
OR2_X1 U941 ( .A1(G902), .A2(n1100), .ZN(n1014) );
AND2_X1 U942 ( .A1(n1231), .A2(n1232), .ZN(n1100) );
NAND4_X1 U943 ( .A1(n1233), .A2(G234), .A3(G217), .A4(n1002), .ZN(n1232) );
XOR2_X1 U944 ( .A(n1234), .B(KEYINPUT40), .Z(n1233) );
NAND2_X1 U945 ( .A1(n1234), .A2(n1235), .ZN(n1231) );
NAND3_X1 U946 ( .A1(G217), .A2(n1002), .A3(G234), .ZN(n1235) );
XOR2_X1 U947 ( .A(n1236), .B(n1237), .Z(n1234) );
NOR3_X1 U948 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1237) );
NOR2_X1 U949 ( .A1(KEYINPUT35), .A2(n1241), .ZN(n1240) );
NOR2_X1 U950 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
AND3_X1 U951 ( .A1(KEYINPUT48), .A2(n1244), .A3(G134), .ZN(n1243) );
NOR2_X1 U952 ( .A1(KEYINPUT48), .A2(G134), .ZN(n1242) );
NOR2_X1 U953 ( .A1(n1245), .A2(n1246), .ZN(n1239) );
INV_X1 U954 ( .A(KEYINPUT35), .ZN(n1246) );
NOR2_X1 U955 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
XNOR2_X1 U956 ( .A(KEYINPUT48), .B(n1249), .ZN(n1248) );
INV_X1 U957 ( .A(n1244), .ZN(n1247) );
NOR2_X1 U958 ( .A1(G134), .A2(n1244), .ZN(n1238) );
XOR2_X1 U959 ( .A(G128), .B(G143), .Z(n1244) );
XOR2_X1 U960 ( .A(n1250), .B(G107), .Z(n1236) );
NAND2_X1 U961 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
OR2_X1 U962 ( .A1(n1253), .A2(G116), .ZN(n1252) );
XOR2_X1 U963 ( .A(n1254), .B(KEYINPUT54), .Z(n1251) );
NAND2_X1 U964 ( .A1(G116), .A2(n1253), .ZN(n1254) );
XOR2_X1 U965 ( .A(G122), .B(KEYINPUT15), .Z(n1253) );
NAND4_X1 U966 ( .A1(n1034), .A2(n1019), .A3(n1212), .A4(n1050), .ZN(n1148) );
NAND2_X1 U967 ( .A1(G221), .A2(n1255), .ZN(n1050) );
NAND2_X1 U968 ( .A1(n1052), .A2(n1256), .ZN(n1212) );
NAND4_X1 U969 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1083), .ZN(n1256) );
INV_X1 U970 ( .A(G898), .ZN(n1083) );
NAND3_X1 U971 ( .A1(n1204), .A2(n1002), .A3(G952), .ZN(n1052) );
NAND2_X1 U972 ( .A1(G237), .A2(n1257), .ZN(n1204) );
XNOR2_X1 U973 ( .A(n1258), .B(G469), .ZN(n1019) );
NAND2_X1 U974 ( .A1(n1259), .A2(n1144), .ZN(n1258) );
XOR2_X1 U975 ( .A(n1260), .B(n1261), .Z(n1259) );
XNOR2_X1 U976 ( .A(n1118), .B(n1063), .ZN(n1261) );
XOR2_X1 U977 ( .A(G128), .B(n1217), .Z(n1063) );
XOR2_X1 U978 ( .A(G143), .B(G146), .Z(n1217) );
INV_X1 U979 ( .A(n1134), .ZN(n1118) );
XOR2_X1 U980 ( .A(n1262), .B(n1263), .Z(n1260) );
XNOR2_X1 U981 ( .A(KEYINPUT23), .B(n1264), .ZN(n1263) );
NOR2_X1 U982 ( .A1(KEYINPUT36), .A2(n1136), .ZN(n1264) );
NAND2_X1 U983 ( .A1(KEYINPUT4), .A2(n1137), .ZN(n1262) );
XNOR2_X1 U984 ( .A(n1265), .B(n1266), .ZN(n1137) );
XNOR2_X1 U985 ( .A(G140), .B(n1214), .ZN(n1266) );
NAND2_X1 U986 ( .A1(G227), .A2(n1002), .ZN(n1265) );
INV_X1 U987 ( .A(n1198), .ZN(n1034) );
NAND2_X1 U988 ( .A1(n1267), .A2(n1038), .ZN(n1198) );
NAND2_X1 U989 ( .A1(G214), .A2(n1268), .ZN(n1038) );
XNOR2_X1 U990 ( .A(KEYINPUT61), .B(n1036), .ZN(n1267) );
XOR2_X1 U991 ( .A(n1269), .B(n1143), .Z(n1036) );
AND2_X1 U992 ( .A1(G210), .A2(n1268), .ZN(n1143) );
NAND2_X1 U993 ( .A1(n1270), .A2(n1144), .ZN(n1268) );
XOR2_X1 U994 ( .A(KEYINPUT20), .B(G237), .Z(n1270) );
NAND2_X1 U995 ( .A1(n1271), .A2(n1144), .ZN(n1269) );
XOR2_X1 U996 ( .A(n1142), .B(n1272), .Z(n1271) );
XNOR2_X1 U997 ( .A(n1273), .B(KEYINPUT18), .ZN(n1272) );
NAND2_X1 U998 ( .A1(KEYINPUT9), .A2(n1140), .ZN(n1273) );
XOR2_X1 U999 ( .A(n1088), .B(n1274), .Z(n1140) );
XOR2_X1 U1000 ( .A(KEYINPUT34), .B(n1087), .Z(n1274) );
XNOR2_X1 U1001 ( .A(n1275), .B(G122), .ZN(n1087) );
NAND2_X1 U1002 ( .A1(KEYINPUT31), .A2(n1214), .ZN(n1275) );
XNOR2_X1 U1003 ( .A(n1276), .B(n1110), .ZN(n1088) );
XNOR2_X1 U1004 ( .A(n1136), .B(KEYINPUT5), .ZN(n1276) );
XOR2_X1 U1005 ( .A(G101), .B(n1277), .Z(n1136) );
XOR2_X1 U1006 ( .A(G107), .B(G104), .Z(n1277) );
XNOR2_X1 U1007 ( .A(n1121), .B(n1278), .ZN(n1142) );
XOR2_X1 U1008 ( .A(G125), .B(n1279), .Z(n1278) );
NOR2_X1 U1009 ( .A1(G953), .A2(n1082), .ZN(n1279) );
INV_X1 U1010 ( .A(G224), .ZN(n1082) );
NAND2_X1 U1011 ( .A1(n1209), .A2(n1206), .ZN(n1042) );
XNOR2_X1 U1012 ( .A(n1280), .B(n1022), .ZN(n1206) );
NOR2_X1 U1013 ( .A1(n1093), .A2(G902), .ZN(n1022) );
XNOR2_X1 U1014 ( .A(n1281), .B(n1282), .ZN(n1093) );
NOR2_X1 U1015 ( .A1(KEYINPUT56), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U1016 ( .A(n1284), .B(n1285), .ZN(n1283) );
AND3_X1 U1017 ( .A1(G221), .A2(n1002), .A3(G234), .ZN(n1285) );
INV_X1 U1018 ( .A(G953), .ZN(n1002) );
NAND3_X1 U1019 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1281) );
NAND2_X1 U1020 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
OR3_X1 U1021 ( .A1(n1290), .A2(n1289), .A3(KEYINPUT39), .ZN(n1287) );
AND3_X1 U1022 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1289) );
NAND2_X1 U1023 ( .A1(G110), .A2(n1294), .ZN(n1293) );
OR3_X1 U1024 ( .A1(n1294), .A2(G110), .A3(KEYINPUT52), .ZN(n1292) );
OR2_X1 U1025 ( .A1(KEYINPUT30), .A2(n1295), .ZN(n1294) );
NAND2_X1 U1026 ( .A1(KEYINPUT52), .A2(n1295), .ZN(n1291) );
XNOR2_X1 U1027 ( .A(G119), .B(G128), .ZN(n1295) );
OR2_X1 U1028 ( .A1(KEYINPUT44), .A2(n1296), .ZN(n1290) );
NAND2_X1 U1029 ( .A1(n1296), .A2(KEYINPUT39), .ZN(n1286) );
XNOR2_X1 U1030 ( .A(n1297), .B(n1298), .ZN(n1296) );
NOR2_X1 U1031 ( .A1(KEYINPUT11), .A2(G125), .ZN(n1298) );
XNOR2_X1 U1032 ( .A(G140), .B(G146), .ZN(n1297) );
NAND2_X1 U1033 ( .A1(KEYINPUT19), .A2(n1094), .ZN(n1280) );
INV_X1 U1034 ( .A(n1021), .ZN(n1094) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1255), .ZN(n1021) );
NAND2_X1 U1036 ( .A1(n1257), .A2(n1144), .ZN(n1255) );
XOR2_X1 U1037 ( .A(G234), .B(KEYINPUT24), .Z(n1257) );
INV_X1 U1038 ( .A(n1010), .ZN(n1209) );
XNOR2_X1 U1039 ( .A(n1299), .B(G472), .ZN(n1010) );
NAND2_X1 U1040 ( .A1(n1300), .A2(n1144), .ZN(n1299) );
INV_X1 U1041 ( .A(G902), .ZN(n1144) );
XNOR2_X1 U1042 ( .A(n1301), .B(n1111), .ZN(n1300) );
XOR2_X1 U1043 ( .A(n1302), .B(n1199), .Z(n1111) );
INV_X1 U1044 ( .A(G101), .ZN(n1199) );
NAND2_X1 U1045 ( .A1(G210), .A2(n1223), .ZN(n1302) );
NOR2_X1 U1046 ( .A1(G953), .A2(G237), .ZN(n1223) );
NAND2_X1 U1047 ( .A1(KEYINPUT58), .A2(n1303), .ZN(n1301) );
XOR2_X1 U1048 ( .A(n1304), .B(n1305), .Z(n1303) );
XNOR2_X1 U1049 ( .A(n1110), .B(n1134), .ZN(n1305) );
XNOR2_X1 U1050 ( .A(n1306), .B(n1307), .ZN(n1134) );
NOR2_X1 U1051 ( .A1(n1067), .A2(n1065), .ZN(n1307) );
NOR2_X1 U1052 ( .A1(n1249), .A2(G137), .ZN(n1065) );
INV_X1 U1053 ( .A(G134), .ZN(n1249) );
NOR2_X1 U1054 ( .A1(n1284), .A2(G134), .ZN(n1067) );
INV_X1 U1055 ( .A(G137), .ZN(n1284) );
NAND2_X1 U1056 ( .A1(KEYINPUT41), .A2(G131), .ZN(n1306) );
XNOR2_X1 U1057 ( .A(n1308), .B(n1309), .ZN(n1110) );
XOR2_X1 U1058 ( .A(KEYINPUT51), .B(G119), .Z(n1309) );
XNOR2_X1 U1059 ( .A(G113), .B(G116), .ZN(n1308) );
XNOR2_X1 U1060 ( .A(KEYINPUT37), .B(n1310), .ZN(n1304) );
NOR2_X1 U1061 ( .A1(KEYINPUT6), .A2(n1121), .ZN(n1310) );
XOR2_X1 U1062 ( .A(n1311), .B(n1312), .Z(n1121) );
NOR2_X1 U1063 ( .A1(G143), .A2(KEYINPUT33), .ZN(n1312) );
XOR2_X1 U1064 ( .A(n1313), .B(G146), .Z(n1311) );
NAND2_X1 U1065 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
INV_X1 U1066 ( .A(G128), .ZN(n1315) );
XNOR2_X1 U1067 ( .A(KEYINPUT8), .B(KEYINPUT38), .ZN(n1314) );
INV_X1 U1068 ( .A(G110), .ZN(n1214) );
endmodule


