//Key = 1100101010000010111000001001001110100001111000111000001101111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323;

XNOR2_X1 U727 ( .A(G107), .B(n997), .ZN(G9) );
NAND3_X1 U728 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
XNOR2_X1 U729 ( .A(KEYINPUT7), .B(n1001), .ZN(n999) );
NOR2_X1 U730 ( .A1(n1002), .A2(n1003), .ZN(G75) );
NOR4_X1 U731 ( .A1(G953), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1003) );
XOR2_X1 U732 ( .A(KEYINPUT2), .B(n1007), .Z(n1006) );
NOR3_X1 U733 ( .A1(n1008), .A2(KEYINPUT20), .A3(n1009), .ZN(n1007) );
INV_X1 U734 ( .A(n1010), .ZN(n1009) );
NOR2_X1 U735 ( .A1(n1011), .A2(n1012), .ZN(n1008) );
NOR2_X1 U736 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U737 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U738 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR2_X1 U739 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U740 ( .A1(n1021), .A2(n1001), .ZN(n1020) );
NOR2_X1 U741 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR2_X1 U742 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U743 ( .A1(n1026), .A2(n1027), .ZN(n1019) );
NOR2_X1 U744 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
AND4_X1 U745 ( .A1(n1001), .A2(n998), .A3(n1030), .A4(KEYINPUT3), .ZN(n1015) );
NOR3_X1 U746 ( .A1(n1027), .A2(n1031), .A3(n1001), .ZN(n1011) );
NOR2_X1 U747 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U748 ( .A1(n1034), .A2(n1018), .ZN(n1033) );
NOR2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U751 ( .A1(n1039), .A2(n1014), .ZN(n1032) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U753 ( .A1(KEYINPUT3), .A2(n1042), .ZN(n1040) );
INV_X1 U754 ( .A(n1030), .ZN(n1027) );
NOR3_X1 U755 ( .A1(n1004), .A2(G953), .A3(G952), .ZN(n1002) );
AND4_X1 U756 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1004) );
NOR4_X1 U757 ( .A1(n1047), .A2(n1048), .A3(n1014), .A4(n1049), .ZN(n1046) );
XOR2_X1 U758 ( .A(n1050), .B(KEYINPUT40), .Z(n1047) );
NOR3_X1 U759 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1045) );
NAND2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1044) );
XOR2_X1 U761 ( .A(KEYINPUT53), .B(n1056), .Z(n1054) );
XOR2_X1 U762 ( .A(KEYINPUT62), .B(n1057), .Z(n1043) );
XOR2_X1 U763 ( .A(n1058), .B(n1059), .Z(G72) );
XOR2_X1 U764 ( .A(n1060), .B(n1061), .Z(n1059) );
NAND2_X1 U765 ( .A1(G953), .A2(n1062), .ZN(n1061) );
NAND2_X1 U766 ( .A1(G900), .A2(G227), .ZN(n1062) );
NAND2_X1 U767 ( .A1(n1063), .A2(n1064), .ZN(n1060) );
NAND2_X1 U768 ( .A1(G953), .A2(n1065), .ZN(n1064) );
XOR2_X1 U769 ( .A(n1066), .B(n1067), .Z(n1063) );
XOR2_X1 U770 ( .A(n1068), .B(n1069), .Z(n1067) );
XOR2_X1 U771 ( .A(n1070), .B(KEYINPUT6), .Z(n1066) );
NOR2_X1 U772 ( .A1(n1071), .A2(G953), .ZN(n1058) );
XOR2_X1 U773 ( .A(n1072), .B(n1073), .Z(G69) );
XOR2_X1 U774 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U775 ( .A1(n1076), .A2(G953), .ZN(n1075) );
NOR2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U777 ( .A(KEYINPUT30), .B(n1079), .Z(n1078) );
NOR2_X1 U778 ( .A1(n1080), .A2(n1081), .ZN(n1074) );
XOR2_X1 U779 ( .A(n1082), .B(n1083), .Z(n1081) );
XOR2_X1 U780 ( .A(n1084), .B(KEYINPUT29), .Z(n1083) );
NAND3_X1 U781 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NAND2_X1 U782 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U783 ( .A1(KEYINPUT51), .A2(n1090), .ZN(n1086) );
NAND2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U785 ( .A(n1093), .B(KEYINPUT34), .ZN(n1091) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1085) );
INV_X1 U787 ( .A(KEYINPUT51), .ZN(n1095) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
OR2_X1 U789 ( .A1(n1093), .A2(KEYINPUT34), .ZN(n1097) );
NAND3_X1 U790 ( .A1(n1093), .A2(n1092), .A3(KEYINPUT34), .ZN(n1096) );
XOR2_X1 U791 ( .A(KEYINPUT28), .B(n1098), .Z(n1080) );
NOR2_X1 U792 ( .A1(G898), .A2(n1099), .ZN(n1098) );
NOR2_X1 U793 ( .A1(n1100), .A2(n1099), .ZN(n1072) );
NOR2_X1 U794 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U795 ( .A1(n1103), .A2(n1104), .ZN(G66) );
XNOR2_X1 U796 ( .A(n1105), .B(n1106), .ZN(n1104) );
NOR3_X1 U797 ( .A1(n1107), .A2(KEYINPUT45), .A3(n1108), .ZN(n1106) );
NOR2_X1 U798 ( .A1(n1103), .A2(n1109), .ZN(G63) );
XNOR2_X1 U799 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U800 ( .A1(n1112), .A2(n1107), .ZN(n1111) );
NOR2_X1 U801 ( .A1(n1103), .A2(n1113), .ZN(G60) );
XNOR2_X1 U802 ( .A(n1114), .B(n1115), .ZN(n1113) );
NOR2_X1 U803 ( .A1(n1116), .A2(n1107), .ZN(n1115) );
XNOR2_X1 U804 ( .A(G104), .B(n1117), .ZN(G6) );
NOR2_X1 U805 ( .A1(n1103), .A2(n1118), .ZN(G57) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U807 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1107), .ZN(n1122) );
NOR2_X1 U809 ( .A1(n1103), .A2(n1124), .ZN(G54) );
XOR2_X1 U810 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U811 ( .A(G146), .B(n1127), .ZN(n1126) );
NAND3_X1 U812 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(n1127) );
OR2_X1 U813 ( .A1(n1131), .A2(KEYINPUT60), .ZN(n1130) );
OR3_X1 U814 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1129) );
INV_X1 U815 ( .A(KEYINPUT60), .ZN(n1132) );
NAND2_X1 U816 ( .A1(n1133), .A2(n1134), .ZN(n1128) );
NAND2_X1 U817 ( .A1(KEYINPUT16), .A2(n1131), .ZN(n1133) );
XOR2_X1 U818 ( .A(G140), .B(G110), .Z(n1131) );
XOR2_X1 U819 ( .A(n1135), .B(n1136), .Z(n1125) );
NOR3_X1 U820 ( .A1(n1107), .A2(KEYINPUT15), .A3(n1137), .ZN(n1136) );
XNOR2_X1 U821 ( .A(G469), .B(KEYINPUT19), .ZN(n1137) );
NOR2_X1 U822 ( .A1(n1103), .A2(n1138), .ZN(G51) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U824 ( .A(n1141), .B(n1142), .ZN(n1140) );
OR3_X1 U825 ( .A1(n1107), .A2(n1055), .A3(n1143), .ZN(n1141) );
INV_X1 U826 ( .A(KEYINPUT14), .ZN(n1143) );
NAND2_X1 U827 ( .A1(G902), .A2(n1005), .ZN(n1107) );
NAND3_X1 U828 ( .A1(n1071), .A2(n1144), .A3(n1079), .ZN(n1005) );
AND4_X1 U829 ( .A1(n1145), .A2(n1117), .A3(n1146), .A4(n1147), .ZN(n1079) );
NAND3_X1 U830 ( .A1(n1000), .A2(n1148), .A3(n1041), .ZN(n1117) );
NAND3_X1 U831 ( .A1(n998), .A2(n1148), .A3(n1000), .ZN(n1145) );
INV_X1 U832 ( .A(n1042), .ZN(n998) );
INV_X1 U833 ( .A(n1077), .ZN(n1144) );
NAND2_X1 U834 ( .A1(n1149), .A2(n1150), .ZN(n1077) );
NAND2_X1 U835 ( .A1(n1151), .A2(n1023), .ZN(n1150) );
XOR2_X1 U836 ( .A(n1152), .B(KEYINPUT0), .Z(n1151) );
NAND3_X1 U837 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
XNOR2_X1 U838 ( .A(n1156), .B(KEYINPUT27), .ZN(n1155) );
NAND2_X1 U839 ( .A1(n1157), .A2(n1158), .ZN(n1149) );
NAND4_X1 U840 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1158) );
OR3_X1 U841 ( .A1(n1042), .A2(n1028), .A3(KEYINPUT1), .ZN(n1162) );
NAND2_X1 U842 ( .A1(KEYINPUT1), .A2(n1163), .ZN(n1161) );
NAND2_X1 U843 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
NAND2_X1 U844 ( .A1(n1041), .A2(n1028), .ZN(n1159) );
AND4_X1 U845 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1071) );
AND4_X1 U846 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
NOR2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(n1168) );
NOR4_X1 U848 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
XOR2_X1 U849 ( .A(KEYINPUT17), .B(n1041), .Z(n1179) );
NOR2_X1 U850 ( .A1(n1036), .A2(n1180), .ZN(n1174) );
NAND4_X1 U851 ( .A1(n1163), .A2(n1030), .A3(n1181), .A4(n1182), .ZN(n1180) );
INV_X1 U852 ( .A(KEYINPUT42), .ZN(n1182) );
NAND2_X1 U853 ( .A1(n1183), .A2(n1184), .ZN(n1167) );
NAND2_X1 U854 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XNOR2_X1 U855 ( .A(KEYINPUT41), .B(n1187), .ZN(n1185) );
NAND2_X1 U856 ( .A1(KEYINPUT42), .A2(n1188), .ZN(n1166) );
XNOR2_X1 U857 ( .A(n1189), .B(n1190), .ZN(n1139) );
NOR2_X1 U858 ( .A1(KEYINPUT52), .A2(n1191), .ZN(n1190) );
NOR3_X1 U859 ( .A1(n1101), .A2(KEYINPUT33), .A3(n1192), .ZN(n1189) );
NOR2_X1 U860 ( .A1(n1099), .A2(G952), .ZN(n1103) );
XOR2_X1 U861 ( .A(n1193), .B(n1194), .Z(G48) );
NOR4_X1 U862 ( .A1(n1195), .A2(n1196), .A3(n1176), .A4(n1197), .ZN(n1194) );
XOR2_X1 U863 ( .A(n1181), .B(KEYINPUT59), .Z(n1197) );
INV_X1 U864 ( .A(n1036), .ZN(n1176) );
NAND2_X1 U865 ( .A1(n1164), .A2(n1041), .ZN(n1195) );
NAND2_X1 U866 ( .A1(KEYINPUT46), .A2(n1198), .ZN(n1193) );
XNOR2_X1 U867 ( .A(G143), .B(n1173), .ZN(G45) );
NAND4_X1 U868 ( .A1(n1036), .A2(n1199), .A3(n1028), .A4(n1200), .ZN(n1173) );
NOR2_X1 U869 ( .A1(n1178), .A2(n1201), .ZN(n1200) );
XOR2_X1 U870 ( .A(n1202), .B(n1203), .Z(G42) );
NOR2_X1 U871 ( .A1(n1187), .A2(n1204), .ZN(n1203) );
NAND2_X1 U872 ( .A1(KEYINPUT8), .A2(n1205), .ZN(n1202) );
NAND3_X1 U873 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(G39) );
NAND2_X1 U874 ( .A1(KEYINPUT11), .A2(n1209), .ZN(n1208) );
NAND3_X1 U875 ( .A1(G137), .A2(n1210), .A3(n1172), .ZN(n1207) );
NAND2_X1 U876 ( .A1(n1211), .A2(n1212), .ZN(n1206) );
NAND2_X1 U877 ( .A1(n1213), .A2(n1210), .ZN(n1212) );
INV_X1 U878 ( .A(KEYINPUT11), .ZN(n1210) );
XNOR2_X1 U879 ( .A(G137), .B(KEYINPUT39), .ZN(n1213) );
INV_X1 U880 ( .A(n1172), .ZN(n1211) );
NAND3_X1 U881 ( .A1(n1164), .A2(n1165), .A3(n1214), .ZN(n1172) );
INV_X1 U882 ( .A(n1177), .ZN(n1164) );
XOR2_X1 U883 ( .A(G134), .B(n1188), .Z(G36) );
AND2_X1 U884 ( .A1(n1163), .A2(n1214), .ZN(n1188) );
XNOR2_X1 U885 ( .A(G131), .B(n1215), .ZN(G33) );
NAND2_X1 U886 ( .A1(n1183), .A2(n1028), .ZN(n1215) );
INV_X1 U887 ( .A(n1204), .ZN(n1183) );
NAND2_X1 U888 ( .A1(n1214), .A2(n1041), .ZN(n1204) );
AND3_X1 U889 ( .A1(n1036), .A2(n1181), .A3(n1030), .ZN(n1214) );
NOR2_X1 U890 ( .A1(n1024), .A2(n1051), .ZN(n1030) );
INV_X1 U891 ( .A(n1216), .ZN(n1024) );
XNOR2_X1 U892 ( .A(n1217), .B(KEYINPUT22), .ZN(n1036) );
XNOR2_X1 U893 ( .A(G128), .B(n1171), .ZN(G30) );
OR4_X1 U894 ( .A1(n1177), .A2(n1178), .A3(n1042), .A4(n1217), .ZN(n1171) );
XNOR2_X1 U895 ( .A(G101), .B(n1146), .ZN(G3) );
NAND3_X1 U896 ( .A1(n1165), .A2(n1000), .A3(n1028), .ZN(n1146) );
XNOR2_X1 U897 ( .A(G125), .B(n1170), .ZN(G27) );
NAND4_X1 U898 ( .A1(n1218), .A2(n1041), .A3(n1029), .A4(n1154), .ZN(n1170) );
INV_X1 U899 ( .A(n1014), .ZN(n1154) );
INV_X1 U900 ( .A(n1178), .ZN(n1218) );
NAND2_X1 U901 ( .A1(n1023), .A2(n1181), .ZN(n1178) );
NAND2_X1 U902 ( .A1(n1219), .A2(n1220), .ZN(n1181) );
NAND3_X1 U903 ( .A1(n1010), .A2(n1099), .A3(G952), .ZN(n1220) );
INV_X1 U904 ( .A(G953), .ZN(n1099) );
XOR2_X1 U905 ( .A(n1221), .B(KEYINPUT25), .Z(n1219) );
NAND4_X1 U906 ( .A1(G953), .A2(G902), .A3(n1010), .A4(n1065), .ZN(n1221) );
INV_X1 U907 ( .A(G900), .ZN(n1065) );
XOR2_X1 U908 ( .A(G122), .B(n1222), .Z(G24) );
AND2_X1 U909 ( .A1(n1153), .A2(n1157), .ZN(n1222) );
NOR3_X1 U910 ( .A1(n1001), .A2(n1223), .A3(n1201), .ZN(n1153) );
INV_X1 U911 ( .A(n1148), .ZN(n1001) );
NOR2_X1 U912 ( .A1(n1224), .A2(n1049), .ZN(n1148) );
XNOR2_X1 U913 ( .A(G119), .B(n1225), .ZN(G21) );
NAND4_X1 U914 ( .A1(n1023), .A2(n1226), .A3(n1156), .A4(n1227), .ZN(n1225) );
NOR2_X1 U915 ( .A1(n1018), .A2(n1177), .ZN(n1227) );
NAND2_X1 U916 ( .A1(n1049), .A2(n1224), .ZN(n1177) );
INV_X1 U917 ( .A(n1228), .ZN(n1156) );
XNOR2_X1 U918 ( .A(KEYINPUT35), .B(n1014), .ZN(n1226) );
XOR2_X1 U919 ( .A(G116), .B(n1229), .Z(G18) );
AND2_X1 U920 ( .A1(n1163), .A2(n1157), .ZN(n1229) );
NOR2_X1 U921 ( .A1(n1186), .A2(n1042), .ZN(n1163) );
NAND2_X1 U922 ( .A1(n1199), .A2(n1201), .ZN(n1042) );
INV_X1 U923 ( .A(n1028), .ZN(n1186) );
XNOR2_X1 U924 ( .A(G113), .B(n1230), .ZN(G15) );
NAND3_X1 U925 ( .A1(n1157), .A2(n1041), .A3(n1231), .ZN(n1230) );
XNOR2_X1 U926 ( .A(n1028), .B(KEYINPUT48), .ZN(n1231) );
NOR2_X1 U927 ( .A1(n1224), .A2(n1232), .ZN(n1028) );
NOR2_X1 U928 ( .A1(n1201), .A2(n1199), .ZN(n1041) );
NOR3_X1 U929 ( .A1(n1228), .A2(n1196), .A3(n1014), .ZN(n1157) );
NAND2_X1 U930 ( .A1(n1233), .A2(n1038), .ZN(n1014) );
INV_X1 U931 ( .A(n1037), .ZN(n1233) );
XOR2_X1 U932 ( .A(n1147), .B(n1234), .Z(G12) );
NOR2_X1 U933 ( .A1(G110), .A2(KEYINPUT26), .ZN(n1234) );
NAND3_X1 U934 ( .A1(n1165), .A2(n1000), .A3(n1029), .ZN(n1147) );
INV_X1 U935 ( .A(n1187), .ZN(n1029) );
NAND2_X1 U936 ( .A1(n1232), .A2(n1224), .ZN(n1187) );
NAND2_X1 U937 ( .A1(n1050), .A2(n1235), .ZN(n1224) );
INV_X1 U938 ( .A(n1052), .ZN(n1235) );
NOR2_X1 U939 ( .A1(n1236), .A2(n1237), .ZN(n1052) );
AND2_X1 U940 ( .A1(G217), .A2(n1238), .ZN(n1237) );
NAND3_X1 U941 ( .A1(n1238), .A2(n1236), .A3(G217), .ZN(n1050) );
NAND2_X1 U942 ( .A1(n1105), .A2(n1239), .ZN(n1236) );
XNOR2_X1 U943 ( .A(n1240), .B(n1241), .ZN(n1105) );
XNOR2_X1 U944 ( .A(n1068), .B(n1242), .ZN(n1241) );
XOR2_X1 U945 ( .A(n1243), .B(n1244), .Z(n1242) );
NOR2_X1 U946 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
INV_X1 U947 ( .A(G221), .ZN(n1245) );
NAND3_X1 U948 ( .A1(n1247), .A2(n1248), .A3(KEYINPUT58), .ZN(n1243) );
NAND2_X1 U949 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
INV_X1 U950 ( .A(KEYINPUT23), .ZN(n1250) );
XNOR2_X1 U951 ( .A(G119), .B(G128), .ZN(n1249) );
NAND3_X1 U952 ( .A1(G128), .A2(n1251), .A3(KEYINPUT23), .ZN(n1247) );
XOR2_X1 U953 ( .A(n1252), .B(n1253), .Z(n1240) );
XNOR2_X1 U954 ( .A(n1209), .B(G110), .ZN(n1253) );
INV_X1 U955 ( .A(G137), .ZN(n1209) );
XNOR2_X1 U956 ( .A(KEYINPUT63), .B(KEYINPUT36), .ZN(n1252) );
INV_X1 U957 ( .A(n1049), .ZN(n1232) );
XOR2_X1 U958 ( .A(n1254), .B(n1123), .Z(n1049) );
INV_X1 U959 ( .A(G472), .ZN(n1123) );
NAND2_X1 U960 ( .A1(n1255), .A2(n1239), .ZN(n1254) );
XOR2_X1 U961 ( .A(n1256), .B(n1257), .Z(n1255) );
XOR2_X1 U962 ( .A(KEYINPUT61), .B(KEYINPUT4), .Z(n1257) );
XOR2_X1 U963 ( .A(n1119), .B(n1258), .Z(n1256) );
NOR2_X1 U964 ( .A1(KEYINPUT13), .A2(n1121), .ZN(n1258) );
NAND2_X1 U965 ( .A1(n1259), .A2(G210), .ZN(n1121) );
XOR2_X1 U966 ( .A(n1260), .B(n1261), .Z(n1119) );
XOR2_X1 U967 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U968 ( .A(n1264), .B(G101), .ZN(n1263) );
INV_X1 U969 ( .A(G113), .ZN(n1264) );
XOR2_X1 U970 ( .A(n1265), .B(n1266), .Z(n1260) );
NOR3_X1 U971 ( .A1(n1196), .A2(n1217), .A3(n1228), .ZN(n1000) );
NAND3_X1 U972 ( .A1(n1267), .A2(n1268), .A3(n1010), .ZN(n1228) );
NAND2_X1 U973 ( .A1(G237), .A2(G234), .ZN(n1010) );
OR2_X1 U974 ( .A1(G952), .A2(G953), .ZN(n1268) );
NAND2_X1 U975 ( .A1(G953), .A2(n1269), .ZN(n1267) );
NAND2_X1 U976 ( .A1(G902), .A2(n1102), .ZN(n1269) );
INV_X1 U977 ( .A(G898), .ZN(n1102) );
NAND2_X1 U978 ( .A1(n1037), .A2(n1038), .ZN(n1217) );
NAND2_X1 U979 ( .A1(G221), .A2(n1238), .ZN(n1038) );
NAND2_X1 U980 ( .A1(G234), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U981 ( .A(n1270), .B(G469), .ZN(n1037) );
NAND2_X1 U982 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XNOR2_X1 U983 ( .A(KEYINPUT57), .B(n1239), .ZN(n1272) );
XOR2_X1 U984 ( .A(n1273), .B(n1274), .Z(n1271) );
XNOR2_X1 U985 ( .A(G110), .B(n1275), .ZN(n1274) );
XNOR2_X1 U986 ( .A(KEYINPUT37), .B(KEYINPUT31), .ZN(n1275) );
XOR2_X1 U987 ( .A(n1135), .B(n1276), .Z(n1273) );
XOR2_X1 U988 ( .A(n1134), .B(n1277), .Z(n1276) );
NAND2_X1 U989 ( .A1(G227), .A2(n1278), .ZN(n1134) );
XOR2_X1 U990 ( .A(n1279), .B(n1280), .Z(n1135) );
XNOR2_X1 U991 ( .A(n1088), .B(n1069), .ZN(n1280) );
XNOR2_X1 U992 ( .A(n1281), .B(KEYINPUT18), .ZN(n1069) );
XOR2_X1 U993 ( .A(n1265), .B(KEYINPUT49), .Z(n1279) );
XOR2_X1 U994 ( .A(n1070), .B(KEYINPUT54), .Z(n1265) );
XOR2_X1 U995 ( .A(n1282), .B(n1283), .Z(n1070) );
XNOR2_X1 U996 ( .A(G137), .B(n1284), .ZN(n1282) );
INV_X1 U997 ( .A(n1023), .ZN(n1196) );
NOR2_X1 U998 ( .A1(n1216), .A2(n1051), .ZN(n1023) );
INV_X1 U999 ( .A(n1025), .ZN(n1051) );
NAND2_X1 U1000 ( .A1(n1285), .A2(n1286), .ZN(n1025) );
XOR2_X1 U1001 ( .A(KEYINPUT50), .B(G214), .Z(n1285) );
NOR2_X1 U1002 ( .A1(n1053), .A2(n1287), .ZN(n1216) );
AND2_X1 U1003 ( .A1(n1056), .A2(n1055), .ZN(n1287) );
NOR2_X1 U1004 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
AND2_X1 U1005 ( .A1(n1288), .A2(n1239), .ZN(n1056) );
XNOR2_X1 U1006 ( .A(n1289), .B(n1290), .ZN(n1288) );
INV_X1 U1007 ( .A(n1142), .ZN(n1290) );
XNOR2_X1 U1008 ( .A(n1291), .B(n1292), .ZN(n1142) );
XNOR2_X1 U1009 ( .A(n1093), .B(n1088), .ZN(n1292) );
INV_X1 U1010 ( .A(n1092), .ZN(n1088) );
XOR2_X1 U1011 ( .A(G101), .B(n1293), .Z(n1092) );
XOR2_X1 U1012 ( .A(G107), .B(G104), .Z(n1293) );
INV_X1 U1013 ( .A(n1089), .ZN(n1093) );
NAND2_X1 U1014 ( .A1(n1294), .A2(n1295), .ZN(n1089) );
NAND2_X1 U1015 ( .A1(G113), .A2(n1262), .ZN(n1295) );
XOR2_X1 U1016 ( .A(n1296), .B(KEYINPUT56), .Z(n1294) );
OR2_X1 U1017 ( .A1(n1262), .A2(G113), .ZN(n1296) );
XNOR2_X1 U1018 ( .A(G116), .B(n1251), .ZN(n1262) );
INV_X1 U1019 ( .A(G119), .ZN(n1251) );
XNOR2_X1 U1020 ( .A(n1297), .B(n1298), .ZN(n1291) );
INV_X1 U1021 ( .A(G125), .ZN(n1298) );
NAND2_X1 U1022 ( .A1(KEYINPUT32), .A2(n1082), .ZN(n1297) );
XNOR2_X1 U1023 ( .A(G110), .B(G122), .ZN(n1082) );
XNOR2_X1 U1024 ( .A(n1191), .B(n1299), .ZN(n1289) );
NOR2_X1 U1025 ( .A1(n1192), .A2(n1101), .ZN(n1299) );
INV_X1 U1026 ( .A(G224), .ZN(n1101) );
XOR2_X1 U1027 ( .A(n1266), .B(G128), .Z(n1191) );
XNOR2_X1 U1028 ( .A(n1300), .B(KEYINPUT38), .ZN(n1266) );
NAND3_X1 U1029 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1300) );
NAND2_X1 U1030 ( .A1(KEYINPUT21), .A2(G143), .ZN(n1303) );
NAND3_X1 U1031 ( .A1(n1304), .A2(n1305), .A3(n1198), .ZN(n1302) );
INV_X1 U1032 ( .A(KEYINPUT21), .ZN(n1305) );
OR2_X1 U1033 ( .A1(n1198), .A2(n1304), .ZN(n1301) );
NOR2_X1 U1034 ( .A1(G143), .A2(KEYINPUT12), .ZN(n1304) );
NAND2_X1 U1035 ( .A1(G210), .A2(n1286), .ZN(n1055) );
NAND2_X1 U1036 ( .A1(n1306), .A2(n1239), .ZN(n1286) );
INV_X1 U1037 ( .A(G237), .ZN(n1306) );
INV_X1 U1038 ( .A(n1018), .ZN(n1165) );
NAND2_X1 U1039 ( .A1(n1223), .A2(n1201), .ZN(n1018) );
XOR2_X1 U1040 ( .A(n1048), .B(KEYINPUT24), .Z(n1201) );
XOR2_X1 U1041 ( .A(n1307), .B(n1116), .Z(n1048) );
INV_X1 U1042 ( .A(G475), .ZN(n1116) );
NAND2_X1 U1043 ( .A1(n1114), .A2(n1239), .ZN(n1307) );
XNOR2_X1 U1044 ( .A(n1308), .B(n1309), .ZN(n1114) );
XNOR2_X1 U1045 ( .A(n1068), .B(n1310), .ZN(n1309) );
XNOR2_X1 U1046 ( .A(n1283), .B(n1311), .ZN(n1310) );
AND2_X1 U1047 ( .A1(G214), .A2(n1259), .ZN(n1311) );
NOR2_X1 U1048 ( .A1(n1192), .A2(G237), .ZN(n1259) );
INV_X1 U1049 ( .A(n1278), .ZN(n1192) );
XOR2_X1 U1050 ( .A(G131), .B(KEYINPUT43), .Z(n1283) );
XNOR2_X1 U1051 ( .A(G125), .B(n1277), .ZN(n1068) );
XNOR2_X1 U1052 ( .A(n1205), .B(n1198), .ZN(n1277) );
INV_X1 U1053 ( .A(G146), .ZN(n1198) );
INV_X1 U1054 ( .A(G140), .ZN(n1205) );
XOR2_X1 U1055 ( .A(n1312), .B(n1313), .Z(n1308) );
NOR2_X1 U1056 ( .A1(KEYINPUT44), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1057 ( .A(n1315), .B(n1316), .Z(n1314) );
NOR2_X1 U1058 ( .A1(KEYINPUT9), .A2(G104), .ZN(n1316) );
XNOR2_X1 U1059 ( .A(G113), .B(G122), .ZN(n1315) );
XNOR2_X1 U1060 ( .A(G143), .B(KEYINPUT47), .ZN(n1312) );
INV_X1 U1061 ( .A(n1199), .ZN(n1223) );
XOR2_X1 U1062 ( .A(n1057), .B(KEYINPUT5), .Z(n1199) );
XOR2_X1 U1063 ( .A(n1317), .B(n1112), .Z(n1057) );
INV_X1 U1064 ( .A(G478), .ZN(n1112) );
NAND2_X1 U1065 ( .A1(n1110), .A2(n1239), .ZN(n1317) );
INV_X1 U1066 ( .A(G902), .ZN(n1239) );
XNOR2_X1 U1067 ( .A(n1318), .B(n1319), .ZN(n1110) );
XOR2_X1 U1068 ( .A(n1320), .B(n1321), .Z(n1319) );
XNOR2_X1 U1069 ( .A(n1281), .B(G107), .ZN(n1321) );
INV_X1 U1070 ( .A(G143), .ZN(n1281) );
NOR2_X1 U1071 ( .A1(KEYINPUT10), .A2(n1322), .ZN(n1320) );
XNOR2_X1 U1072 ( .A(G116), .B(G122), .ZN(n1322) );
XNOR2_X1 U1073 ( .A(n1284), .B(n1323), .ZN(n1318) );
NOR2_X1 U1074 ( .A1(n1246), .A2(n1108), .ZN(n1323) );
INV_X1 U1075 ( .A(G217), .ZN(n1108) );
NAND2_X1 U1076 ( .A1(G234), .A2(n1278), .ZN(n1246) );
XOR2_X1 U1077 ( .A(G953), .B(KEYINPUT55), .Z(n1278) );
XOR2_X1 U1078 ( .A(G134), .B(G128), .Z(n1284) );
endmodule


