//Key = 1000101010010010010110011110000011011111011001010100110101000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407;

XNOR2_X1 U774 ( .A(G107), .B(n1069), .ZN(G9) );
NAND4_X1 U775 ( .A1(KEYINPUT61), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1069) );
NAND4_X1 U776 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(G75) );
NAND4_X1 U777 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1075) );
NOR3_X1 U778 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
INV_X1 U779 ( .A(n1084), .ZN(n1079) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1078) );
NAND2_X1 U781 ( .A1(n1070), .A2(n1087), .ZN(n1086) );
NAND3_X1 U782 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1077) );
NAND2_X1 U783 ( .A1(n1087), .A2(n1091), .ZN(n1089) );
NAND2_X1 U784 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U785 ( .A1(n1070), .A2(n1094), .ZN(n1088) );
NAND2_X1 U786 ( .A1(n1095), .A2(n1090), .ZN(n1074) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND4_X1 U788 ( .A1(n1098), .A2(n1087), .A3(n1070), .A4(n1099), .ZN(n1097) );
NOR3_X1 U789 ( .A1(n1084), .A2(n1100), .A3(n1101), .ZN(n1099) );
NOR4_X1 U790 ( .A1(n1081), .A2(n1072), .A3(n1102), .A4(n1082), .ZN(n1101) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND2_X1 U792 ( .A1(n1082), .A2(n1105), .ZN(n1098) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1103), .ZN(n1105) );
NAND4_X1 U794 ( .A1(n1106), .A2(n1070), .A3(n1107), .A4(n1108), .ZN(n1096) );
NOR4_X1 U795 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
XNOR2_X1 U796 ( .A(KEYINPUT46), .B(n1113), .ZN(n1112) );
XNOR2_X1 U797 ( .A(G469), .B(n1114), .ZN(n1111) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1110) );
INV_X1 U799 ( .A(KEYINPUT26), .ZN(n1115) );
NOR2_X1 U800 ( .A1(KEYINPUT26), .A2(n1117), .ZN(n1109) );
AND2_X1 U801 ( .A1(n1118), .A2(n1119), .ZN(n1107) );
XOR2_X1 U802 ( .A(n1120), .B(KEYINPUT33), .Z(n1106) );
NAND2_X1 U803 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U804 ( .A1(G478), .A2(n1123), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(G72) );
NAND2_X1 U806 ( .A1(G953), .A2(n1126), .ZN(n1125) );
NAND2_X1 U807 ( .A1(G900), .A2(n1127), .ZN(n1126) );
NAND2_X1 U808 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U809 ( .A(n1130), .B(KEYINPUT16), .Z(n1124) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U811 ( .A1(G953), .A2(n1129), .ZN(n1132) );
INV_X1 U812 ( .A(G227), .ZN(n1129) );
XNOR2_X1 U813 ( .A(n1133), .B(n1128), .ZN(n1131) );
NAND2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(n1128) );
NAND2_X1 U815 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XNOR2_X1 U816 ( .A(n1138), .B(n1139), .ZN(n1136) );
XOR2_X1 U817 ( .A(n1140), .B(KEYINPUT28), .Z(n1134) );
NAND2_X1 U818 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XNOR2_X1 U819 ( .A(n1139), .B(n1143), .ZN(n1142) );
INV_X1 U820 ( .A(n1138), .ZN(n1143) );
XOR2_X1 U821 ( .A(G137), .B(n1144), .Z(n1138) );
NOR2_X1 U822 ( .A1(KEYINPUT13), .A2(n1145), .ZN(n1144) );
XOR2_X1 U823 ( .A(n1146), .B(n1147), .Z(G69) );
NOR2_X1 U824 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U825 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U826 ( .A(KEYINPUT47), .B(n1152), .Z(n1151) );
NOR2_X1 U827 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
NOR3_X1 U828 ( .A1(n1154), .A2(n1153), .A3(n1152), .ZN(n1148) );
AND2_X1 U829 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
NAND2_X1 U830 ( .A1(G953), .A2(n1157), .ZN(n1156) );
INV_X1 U831 ( .A(n1158), .ZN(n1153) );
XNOR2_X1 U832 ( .A(G953), .B(KEYINPUT55), .ZN(n1154) );
NAND2_X1 U833 ( .A1(G953), .A2(n1159), .ZN(n1146) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1159) );
NOR2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(G66) );
XNOR2_X1 U836 ( .A(n1162), .B(n1163), .ZN(n1161) );
NOR2_X1 U837 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NOR2_X1 U838 ( .A1(n1160), .A2(n1166), .ZN(G63) );
XOR2_X1 U839 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U840 ( .A1(n1169), .A2(n1165), .ZN(n1167) );
NOR2_X1 U841 ( .A1(n1160), .A2(n1170), .ZN(G60) );
XOR2_X1 U842 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1165), .ZN(n1171) );
XNOR2_X1 U844 ( .A(G104), .B(n1174), .ZN(G6) );
NOR3_X1 U845 ( .A1(n1175), .A2(n1160), .A3(n1176), .ZN(G57) );
NOR4_X1 U846 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
NOR2_X1 U847 ( .A1(n1181), .A2(n1182), .ZN(n1178) );
NOR2_X1 U848 ( .A1(G101), .A2(n1183), .ZN(n1177) );
NOR3_X1 U849 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1175) );
NOR2_X1 U850 ( .A1(G101), .A2(n1182), .ZN(n1186) );
XOR2_X1 U851 ( .A(n1183), .B(n1187), .Z(n1182) );
XOR2_X1 U852 ( .A(KEYINPUT34), .B(KEYINPUT20), .Z(n1187) );
NOR2_X1 U853 ( .A1(n1181), .A2(n1183), .ZN(n1185) );
XOR2_X1 U854 ( .A(n1188), .B(n1189), .Z(n1183) );
NOR2_X1 U855 ( .A1(n1190), .A2(n1165), .ZN(n1189) );
NAND2_X1 U856 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
NAND2_X1 U857 ( .A1(n1193), .A2(n1145), .ZN(n1192) );
XOR2_X1 U858 ( .A(KEYINPUT44), .B(n1194), .Z(n1193) );
NAND2_X1 U859 ( .A1(n1195), .A2(n1196), .ZN(n1191) );
XOR2_X1 U860 ( .A(KEYINPUT57), .B(n1194), .Z(n1195) );
NOR2_X1 U861 ( .A1(n1179), .A2(n1180), .ZN(n1184) );
INV_X1 U862 ( .A(KEYINPUT17), .ZN(n1180) );
NOR2_X1 U863 ( .A1(n1160), .A2(n1197), .ZN(G54) );
XOR2_X1 U864 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U865 ( .A(n1200), .B(n1201), .ZN(n1199) );
NAND2_X1 U866 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
NAND3_X1 U867 ( .A1(KEYINPUT0), .A2(n1196), .A3(n1204), .ZN(n1203) );
XNOR2_X1 U868 ( .A(n1205), .B(n1206), .ZN(n1204) );
NOR2_X1 U869 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
INV_X1 U870 ( .A(KEYINPUT52), .ZN(n1208) );
NAND2_X1 U871 ( .A1(n1209), .A2(n1210), .ZN(n1202) );
NAND2_X1 U872 ( .A1(KEYINPUT0), .A2(n1196), .ZN(n1210) );
XNOR2_X1 U873 ( .A(n1211), .B(n1212), .ZN(n1209) );
INV_X1 U874 ( .A(n1205), .ZN(n1212) );
XOR2_X1 U875 ( .A(n1213), .B(KEYINPUT50), .Z(n1205) );
NAND2_X1 U876 ( .A1(KEYINPUT52), .A2(n1207), .ZN(n1211) );
XOR2_X1 U877 ( .A(KEYINPUT8), .B(n1214), .Z(n1198) );
NOR2_X1 U878 ( .A1(n1215), .A2(n1165), .ZN(n1214) );
NOR3_X1 U879 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(G51) );
NOR3_X1 U880 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1218) );
NOR2_X1 U881 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
XNOR2_X1 U882 ( .A(KEYINPUT53), .B(n1224), .ZN(n1223) );
NOR2_X1 U883 ( .A1(n1225), .A2(n1226), .ZN(n1217) );
NOR2_X1 U884 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
AND2_X1 U885 ( .A1(KEYINPUT53), .A2(n1221), .ZN(n1228) );
AND2_X1 U886 ( .A1(n1224), .A2(n1222), .ZN(n1221) );
NOR2_X1 U887 ( .A1(n1229), .A2(n1224), .ZN(n1227) );
XNOR2_X1 U888 ( .A(n1230), .B(n1231), .ZN(n1224) );
NOR3_X1 U889 ( .A1(n1232), .A2(n1233), .A3(n1165), .ZN(n1231) );
OR2_X1 U890 ( .A1(n1234), .A2(n1073), .ZN(n1165) );
NOR2_X1 U891 ( .A1(n1158), .A2(n1133), .ZN(n1073) );
NAND2_X1 U892 ( .A1(n1235), .A2(n1236), .ZN(n1133) );
AND4_X1 U893 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1236) );
NOR4_X1 U894 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1235) );
NOR3_X1 U895 ( .A1(n1245), .A2(n1246), .A3(n1092), .ZN(n1244) );
INV_X1 U896 ( .A(n1247), .ZN(n1243) );
NAND4_X1 U897 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1158) );
AND4_X1 U898 ( .A1(n1174), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1251) );
NAND3_X1 U899 ( .A1(n1070), .A2(n1071), .A3(n1102), .ZN(n1174) );
NOR2_X1 U900 ( .A1(n1255), .A2(n1256), .ZN(n1250) );
NOR3_X1 U901 ( .A1(n1257), .A2(n1246), .A3(n1258), .ZN(n1256) );
XOR2_X1 U902 ( .A(KEYINPUT45), .B(n1070), .Z(n1257) );
INV_X1 U903 ( .A(G210), .ZN(n1233) );
XNOR2_X1 U904 ( .A(KEYINPUT30), .B(n1259), .ZN(n1232) );
AND2_X1 U905 ( .A1(n1222), .A2(KEYINPUT53), .ZN(n1229) );
XOR2_X1 U906 ( .A(KEYINPUT58), .B(n1160), .Z(n1216) );
NOR2_X1 U907 ( .A1(n1260), .A2(G952), .ZN(n1160) );
XNOR2_X1 U908 ( .A(KEYINPUT54), .B(G953), .ZN(n1260) );
XNOR2_X1 U909 ( .A(G146), .B(n1240), .ZN(G48) );
NAND3_X1 U910 ( .A1(n1102), .A2(n1261), .A3(n1262), .ZN(n1240) );
NAND2_X1 U911 ( .A1(n1263), .A2(n1264), .ZN(G45) );
OR2_X1 U912 ( .A1(n1247), .A2(G143), .ZN(n1264) );
XOR2_X1 U913 ( .A(n1265), .B(KEYINPUT62), .Z(n1263) );
NAND2_X1 U914 ( .A1(G143), .A2(n1247), .ZN(n1265) );
NAND3_X1 U915 ( .A1(n1266), .A2(n1261), .A3(n1267), .ZN(n1247) );
NOR3_X1 U916 ( .A1(n1119), .A2(n1268), .A3(n1269), .ZN(n1267) );
XNOR2_X1 U917 ( .A(G140), .B(n1239), .ZN(G42) );
OR3_X1 U918 ( .A1(n1093), .A2(n1270), .A3(n1245), .ZN(n1239) );
INV_X1 U919 ( .A(n1271), .ZN(n1093) );
XNOR2_X1 U920 ( .A(n1272), .B(n1242), .ZN(G39) );
NOR3_X1 U921 ( .A1(n1273), .A2(n1274), .A3(n1245), .ZN(n1242) );
XNOR2_X1 U922 ( .A(n1275), .B(n1276), .ZN(G36) );
NOR3_X1 U923 ( .A1(n1277), .A2(n1246), .A3(n1245), .ZN(n1276) );
INV_X1 U924 ( .A(n1072), .ZN(n1246) );
XNOR2_X1 U925 ( .A(KEYINPUT24), .B(n1092), .ZN(n1277) );
XOR2_X1 U926 ( .A(G131), .B(n1241), .Z(G33) );
NOR3_X1 U927 ( .A1(n1092), .A2(n1270), .A3(n1245), .ZN(n1241) );
NAND3_X1 U928 ( .A1(n1081), .A2(n1087), .A3(n1278), .ZN(n1245) );
NOR3_X1 U929 ( .A1(n1269), .A2(n1085), .A3(n1082), .ZN(n1278) );
INV_X1 U930 ( .A(n1113), .ZN(n1082) );
INV_X1 U931 ( .A(n1090), .ZN(n1085) );
XNOR2_X1 U932 ( .A(n1094), .B(KEYINPUT31), .ZN(n1087) );
XNOR2_X1 U933 ( .A(G128), .B(n1238), .ZN(G30) );
NAND3_X1 U934 ( .A1(n1072), .A2(n1261), .A3(n1262), .ZN(n1238) );
NOR3_X1 U935 ( .A1(n1279), .A2(n1269), .A3(n1273), .ZN(n1262) );
XNOR2_X1 U936 ( .A(n1181), .B(n1255), .ZN(G3) );
NOR3_X1 U937 ( .A1(n1083), .A2(n1258), .A3(n1092), .ZN(n1255) );
INV_X1 U938 ( .A(n1266), .ZN(n1092) );
INV_X1 U939 ( .A(n1103), .ZN(n1083) );
XNOR2_X1 U940 ( .A(G125), .B(n1237), .ZN(G27) );
NAND3_X1 U941 ( .A1(n1104), .A2(n1271), .A3(n1280), .ZN(n1237) );
NOR3_X1 U942 ( .A1(n1270), .A2(n1269), .A3(n1281), .ZN(n1280) );
AND2_X1 U943 ( .A1(n1084), .A2(n1282), .ZN(n1269) );
NAND4_X1 U944 ( .A1(G953), .A2(G902), .A3(n1283), .A4(n1284), .ZN(n1282) );
INV_X1 U945 ( .A(G900), .ZN(n1284) );
INV_X1 U946 ( .A(n1102), .ZN(n1270) );
NOR2_X1 U947 ( .A1(n1285), .A2(n1279), .ZN(n1271) );
INV_X1 U948 ( .A(n1286), .ZN(n1279) );
XOR2_X1 U949 ( .A(n1248), .B(n1287), .Z(G24) );
NAND2_X1 U950 ( .A1(KEYINPUT4), .A2(G122), .ZN(n1287) );
NAND4_X1 U951 ( .A1(n1288), .A2(n1070), .A3(n1289), .A4(n1290), .ZN(n1248) );
NOR2_X1 U952 ( .A1(n1286), .A2(n1285), .ZN(n1070) );
NAND2_X1 U953 ( .A1(n1291), .A2(n1292), .ZN(G21) );
NAND2_X1 U954 ( .A1(G119), .A2(n1249), .ZN(n1292) );
XOR2_X1 U955 ( .A(n1293), .B(KEYINPUT22), .Z(n1291) );
OR2_X1 U956 ( .A1(n1249), .A2(G119), .ZN(n1293) );
NAND3_X1 U957 ( .A1(n1285), .A2(n1294), .A3(n1288), .ZN(n1249) );
INV_X1 U958 ( .A(n1273), .ZN(n1285) );
XNOR2_X1 U959 ( .A(G116), .B(n1254), .ZN(G18) );
NAND3_X1 U960 ( .A1(n1288), .A2(n1072), .A3(n1266), .ZN(n1254) );
NOR2_X1 U961 ( .A1(n1289), .A2(n1268), .ZN(n1072) );
INV_X1 U962 ( .A(n1290), .ZN(n1268) );
NAND2_X1 U963 ( .A1(n1295), .A2(n1296), .ZN(G15) );
NAND2_X1 U964 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XNOR2_X1 U965 ( .A(KEYINPUT21), .B(n1253), .ZN(n1297) );
NAND2_X1 U966 ( .A1(n1299), .A2(G113), .ZN(n1295) );
XNOR2_X1 U967 ( .A(KEYINPUT11), .B(n1253), .ZN(n1299) );
NAND3_X1 U968 ( .A1(n1288), .A2(n1102), .A3(n1266), .ZN(n1253) );
NOR2_X1 U969 ( .A1(n1273), .A2(n1286), .ZN(n1266) );
NOR2_X1 U970 ( .A1(n1290), .A2(n1119), .ZN(n1102) );
INV_X1 U971 ( .A(n1289), .ZN(n1119) );
NOR3_X1 U972 ( .A1(n1281), .A2(n1300), .A3(n1081), .ZN(n1288) );
INV_X1 U973 ( .A(n1104), .ZN(n1081) );
INV_X1 U974 ( .A(n1301), .ZN(n1300) );
XNOR2_X1 U975 ( .A(G110), .B(n1252), .ZN(G12) );
NAND3_X1 U976 ( .A1(n1071), .A2(n1273), .A3(n1294), .ZN(n1252) );
INV_X1 U977 ( .A(n1274), .ZN(n1294) );
NAND2_X1 U978 ( .A1(n1103), .A2(n1286), .ZN(n1274) );
XOR2_X1 U979 ( .A(n1302), .B(n1164), .Z(n1286) );
NAND2_X1 U980 ( .A1(G217), .A2(n1303), .ZN(n1164) );
NAND2_X1 U981 ( .A1(n1162), .A2(n1234), .ZN(n1302) );
XNOR2_X1 U982 ( .A(n1304), .B(n1305), .ZN(n1162) );
XOR2_X1 U983 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U984 ( .A(n1308), .B(G128), .ZN(n1307) );
XOR2_X1 U985 ( .A(KEYINPUT59), .B(KEYINPUT42), .Z(n1306) );
XOR2_X1 U986 ( .A(n1309), .B(n1310), .Z(n1304) );
XOR2_X1 U987 ( .A(n1311), .B(n1312), .Z(n1310) );
NOR2_X1 U988 ( .A1(G137), .A2(KEYINPUT43), .ZN(n1312) );
AND3_X1 U989 ( .A1(G221), .A2(n1076), .A3(G234), .ZN(n1311) );
XNOR2_X1 U990 ( .A(n1313), .B(n1141), .ZN(n1309) );
NOR2_X1 U991 ( .A1(n1290), .A2(n1289), .ZN(n1103) );
XNOR2_X1 U992 ( .A(n1314), .B(n1315), .ZN(n1289) );
XNOR2_X1 U993 ( .A(KEYINPUT48), .B(n1173), .ZN(n1315) );
INV_X1 U994 ( .A(G475), .ZN(n1173) );
OR2_X1 U995 ( .A1(n1172), .A2(G902), .ZN(n1314) );
XNOR2_X1 U996 ( .A(n1316), .B(n1317), .ZN(n1172) );
XOR2_X1 U997 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U998 ( .A(n1320), .B(n1321), .Z(n1319) );
NOR2_X1 U999 ( .A1(KEYINPUT3), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1000 ( .A(n1323), .B(n1324), .Z(n1322) );
NAND2_X1 U1001 ( .A1(KEYINPUT19), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1002 ( .A1(n1326), .A2(n1327), .ZN(n1320) );
NAND2_X1 U1003 ( .A1(n1137), .A2(n1328), .ZN(n1327) );
NAND2_X1 U1004 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U1005 ( .A1(n1308), .A2(n1331), .ZN(n1330) );
INV_X1 U1006 ( .A(G146), .ZN(n1308) );
INV_X1 U1007 ( .A(n1141), .ZN(n1137) );
NAND2_X1 U1008 ( .A1(G146), .A2(n1332), .ZN(n1326) );
NAND2_X1 U1009 ( .A1(n1331), .A2(n1333), .ZN(n1332) );
NAND2_X1 U1010 ( .A1(n1141), .A2(n1329), .ZN(n1333) );
INV_X1 U1011 ( .A(KEYINPUT51), .ZN(n1329) );
XNOR2_X1 U1012 ( .A(G140), .B(G125), .ZN(n1141) );
INV_X1 U1013 ( .A(KEYINPUT56), .ZN(n1331) );
NAND2_X1 U1014 ( .A1(G214), .A2(n1334), .ZN(n1318) );
XNOR2_X1 U1015 ( .A(G131), .B(n1335), .ZN(n1316) );
XOR2_X1 U1016 ( .A(KEYINPUT23), .B(G143), .Z(n1335) );
NAND3_X1 U1017 ( .A1(n1336), .A2(n1337), .A3(n1121), .ZN(n1290) );
NAND2_X1 U1018 ( .A1(n1338), .A2(n1169), .ZN(n1121) );
INV_X1 U1019 ( .A(G478), .ZN(n1169) );
OR2_X1 U1020 ( .A1(G478), .A2(KEYINPUT39), .ZN(n1337) );
NAND3_X1 U1021 ( .A1(G478), .A2(n1123), .A3(KEYINPUT39), .ZN(n1336) );
INV_X1 U1022 ( .A(n1338), .ZN(n1123) );
NOR2_X1 U1023 ( .A1(n1168), .A2(G902), .ZN(n1338) );
XNOR2_X1 U1024 ( .A(n1339), .B(n1340), .ZN(n1168) );
XNOR2_X1 U1025 ( .A(G134), .B(n1341), .ZN(n1340) );
NAND3_X1 U1026 ( .A1(G234), .A2(n1076), .A3(G217), .ZN(n1341) );
XNOR2_X1 U1027 ( .A(n1342), .B(n1343), .ZN(n1339) );
NOR2_X1 U1028 ( .A1(KEYINPUT12), .A2(n1344), .ZN(n1343) );
XNOR2_X1 U1029 ( .A(n1345), .B(n1346), .ZN(n1273) );
XNOR2_X1 U1030 ( .A(KEYINPUT38), .B(n1190), .ZN(n1346) );
INV_X1 U1031 ( .A(G472), .ZN(n1190) );
NAND2_X1 U1032 ( .A1(n1347), .A2(n1234), .ZN(n1345) );
XOR2_X1 U1033 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1034 ( .A(n1350), .B(n1194), .Z(n1349) );
XNOR2_X1 U1035 ( .A(n1351), .B(n1352), .ZN(n1194) );
XNOR2_X1 U1036 ( .A(G113), .B(n1353), .ZN(n1352) );
NAND2_X1 U1037 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NAND2_X1 U1038 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1039 ( .A(n1358), .B(KEYINPUT40), .Z(n1354) );
OR2_X1 U1040 ( .A1(n1357), .A2(n1356), .ZN(n1358) );
XOR2_X1 U1041 ( .A(n1359), .B(KEYINPUT10), .Z(n1356) );
INV_X1 U1042 ( .A(G116), .ZN(n1357) );
NOR2_X1 U1043 ( .A1(n1360), .A2(n1361), .ZN(n1350) );
XOR2_X1 U1044 ( .A(n1362), .B(KEYINPUT36), .Z(n1361) );
NAND2_X1 U1045 ( .A1(n1181), .A2(n1179), .ZN(n1362) );
NOR2_X1 U1046 ( .A1(n1179), .A2(n1181), .ZN(n1360) );
NAND2_X1 U1047 ( .A1(G210), .A2(n1334), .ZN(n1179) );
NOR2_X1 U1048 ( .A1(G953), .A2(G237), .ZN(n1334) );
XNOR2_X1 U1049 ( .A(n1363), .B(KEYINPUT63), .ZN(n1348) );
NAND2_X1 U1050 ( .A1(n1364), .A2(KEYINPUT49), .ZN(n1363) );
XNOR2_X1 U1051 ( .A(n1196), .B(KEYINPUT9), .ZN(n1364) );
INV_X1 U1052 ( .A(n1258), .ZN(n1071) );
NAND2_X1 U1053 ( .A1(n1261), .A2(n1301), .ZN(n1258) );
NAND2_X1 U1054 ( .A1(n1084), .A2(n1365), .ZN(n1301) );
NAND4_X1 U1055 ( .A1(G953), .A2(G902), .A3(n1283), .A4(n1157), .ZN(n1365) );
INV_X1 U1056 ( .A(G898), .ZN(n1157) );
NAND3_X1 U1057 ( .A1(n1283), .A2(n1076), .A3(G952), .ZN(n1084) );
NAND2_X1 U1058 ( .A1(G237), .A2(n1366), .ZN(n1283) );
NOR2_X1 U1059 ( .A1(n1281), .A2(n1104), .ZN(n1261) );
XOR2_X1 U1060 ( .A(n1367), .B(n1215), .Z(n1104) );
INV_X1 U1061 ( .A(G469), .ZN(n1215) );
NAND2_X1 U1062 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
NAND2_X1 U1063 ( .A1(KEYINPUT35), .A2(n1370), .ZN(n1369) );
OR2_X1 U1064 ( .A1(KEYINPUT37), .A2(n1370), .ZN(n1368) );
INV_X1 U1065 ( .A(n1114), .ZN(n1370) );
NAND3_X1 U1066 ( .A1(n1371), .A2(n1372), .A3(n1234), .ZN(n1114) );
NAND2_X1 U1067 ( .A1(n1213), .A2(n1373), .ZN(n1372) );
NAND2_X1 U1068 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U1069 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
XNOR2_X1 U1070 ( .A(KEYINPUT60), .B(n1378), .ZN(n1377) );
XNOR2_X1 U1071 ( .A(n1201), .B(KEYINPUT7), .ZN(n1376) );
NAND2_X1 U1072 ( .A1(n1379), .A2(n1201), .ZN(n1374) );
XOR2_X1 U1073 ( .A(n1378), .B(KEYINPUT60), .Z(n1379) );
NAND2_X1 U1074 ( .A1(n1380), .A2(n1351), .ZN(n1371) );
INV_X1 U1075 ( .A(n1213), .ZN(n1351) );
XOR2_X1 U1076 ( .A(n1139), .B(n1381), .Z(n1213) );
XNOR2_X1 U1077 ( .A(n1382), .B(KEYINPUT5), .ZN(n1381) );
NAND2_X1 U1078 ( .A1(KEYINPUT32), .A2(n1272), .ZN(n1382) );
INV_X1 U1079 ( .A(G137), .ZN(n1272) );
XNOR2_X1 U1080 ( .A(G131), .B(n1275), .ZN(n1139) );
INV_X1 U1081 ( .A(G134), .ZN(n1275) );
XNOR2_X1 U1082 ( .A(n1383), .B(n1201), .ZN(n1380) );
XNOR2_X1 U1083 ( .A(n1384), .B(n1385), .ZN(n1201) );
XNOR2_X1 U1084 ( .A(G140), .B(n1386), .ZN(n1385) );
INV_X1 U1085 ( .A(G110), .ZN(n1386) );
NAND2_X1 U1086 ( .A1(G227), .A2(n1076), .ZN(n1384) );
NAND2_X1 U1087 ( .A1(n1378), .A2(n1387), .ZN(n1383) );
INV_X1 U1088 ( .A(KEYINPUT7), .ZN(n1387) );
XOR2_X1 U1089 ( .A(n1388), .B(n1389), .Z(n1378) );
XOR2_X1 U1090 ( .A(KEYINPUT6), .B(KEYINPUT29), .Z(n1389) );
XNOR2_X1 U1091 ( .A(n1207), .B(n1145), .ZN(n1388) );
NAND2_X1 U1092 ( .A1(n1390), .A2(n1391), .ZN(n1207) );
NAND2_X1 U1093 ( .A1(n1392), .A2(n1181), .ZN(n1391) );
XOR2_X1 U1094 ( .A(n1393), .B(KEYINPUT15), .Z(n1390) );
OR2_X1 U1095 ( .A1(n1392), .A2(n1181), .ZN(n1393) );
XOR2_X1 U1096 ( .A(G104), .B(n1394), .Z(n1392) );
XOR2_X1 U1097 ( .A(KEYINPUT14), .B(G107), .Z(n1394) );
NAND3_X1 U1098 ( .A1(n1113), .A2(n1090), .A3(n1094), .ZN(n1281) );
NAND2_X1 U1099 ( .A1(n1116), .A2(n1118), .ZN(n1094) );
NAND3_X1 U1100 ( .A1(n1395), .A2(n1259), .A3(G210), .ZN(n1118) );
NAND2_X1 U1101 ( .A1(n1117), .A2(n1396), .ZN(n1116) );
NAND2_X1 U1102 ( .A1(G210), .A2(n1259), .ZN(n1396) );
INV_X1 U1103 ( .A(n1395), .ZN(n1117) );
NAND2_X1 U1104 ( .A1(n1397), .A2(n1234), .ZN(n1395) );
XNOR2_X1 U1105 ( .A(n1155), .B(n1398), .ZN(n1397) );
XNOR2_X1 U1106 ( .A(n1219), .B(n1399), .ZN(n1398) );
NAND3_X1 U1107 ( .A1(n1400), .A2(n1401), .A3(KEYINPUT41), .ZN(n1399) );
OR2_X1 U1108 ( .A1(n1222), .A2(KEYINPUT18), .ZN(n1401) );
XNOR2_X1 U1109 ( .A(G125), .B(n1145), .ZN(n1222) );
NAND3_X1 U1110 ( .A1(G125), .A2(n1145), .A3(KEYINPUT18), .ZN(n1400) );
INV_X1 U1111 ( .A(n1196), .ZN(n1145) );
XOR2_X1 U1112 ( .A(G146), .B(n1342), .Z(n1196) );
XOR2_X1 U1113 ( .A(G128), .B(G143), .Z(n1342) );
INV_X1 U1114 ( .A(n1226), .ZN(n1219) );
NAND2_X1 U1115 ( .A1(G224), .A2(n1076), .ZN(n1226) );
INV_X1 U1116 ( .A(G953), .ZN(n1076) );
INV_X1 U1117 ( .A(n1230), .ZN(n1155) );
XNOR2_X1 U1118 ( .A(n1402), .B(n1403), .ZN(n1230) );
XOR2_X1 U1119 ( .A(n1344), .B(n1404), .Z(n1403) );
XNOR2_X1 U1120 ( .A(KEYINPUT2), .B(n1181), .ZN(n1404) );
INV_X1 U1121 ( .A(G101), .ZN(n1181) );
XOR2_X1 U1122 ( .A(G107), .B(n1405), .Z(n1344) );
XNOR2_X1 U1123 ( .A(n1325), .B(G116), .ZN(n1405) );
INV_X1 U1124 ( .A(G122), .ZN(n1325) );
XOR2_X1 U1125 ( .A(n1313), .B(n1324), .Z(n1402) );
XNOR2_X1 U1126 ( .A(G104), .B(n1298), .ZN(n1324) );
INV_X1 U1127 ( .A(G113), .ZN(n1298) );
XNOR2_X1 U1128 ( .A(G110), .B(n1359), .ZN(n1313) );
XOR2_X1 U1129 ( .A(G119), .B(KEYINPUT1), .Z(n1359) );
NAND2_X1 U1130 ( .A1(G214), .A2(n1259), .ZN(n1090) );
NAND2_X1 U1131 ( .A1(n1406), .A2(n1407), .ZN(n1259) );
INV_X1 U1132 ( .A(G237), .ZN(n1407) );
NAND2_X1 U1133 ( .A1(G221), .A2(n1303), .ZN(n1113) );
NAND2_X1 U1134 ( .A1(n1366), .A2(n1406), .ZN(n1303) );
XNOR2_X1 U1135 ( .A(n1234), .B(KEYINPUT25), .ZN(n1406) );
INV_X1 U1136 ( .A(G902), .ZN(n1234) );
XOR2_X1 U1137 ( .A(G234), .B(KEYINPUT27), .Z(n1366) );
endmodule


