//Key = 1111001101010110110101101111001001111101011100100011011010011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316;

XOR2_X1 U720 ( .A(G107), .B(n994), .Z(G9) );
NOR2_X1 U721 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR3_X1 U722 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
XOR2_X1 U723 ( .A(n1000), .B(KEYINPUT21), .Z(n998) );
NAND2_X1 U724 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NAND2_X1 U725 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND3_X1 U726 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
NAND2_X1 U727 ( .A1(n1008), .A2(n1009), .ZN(n1003) );
NAND2_X1 U728 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U729 ( .A1(n1006), .A2(n1012), .ZN(n1011) );
NAND2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U731 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U732 ( .A1(n1017), .A2(n1018), .ZN(n1013) );
NAND2_X1 U733 ( .A1(n1007), .A2(n1019), .ZN(n1010) );
NAND3_X1 U734 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n997) );
NAND2_X1 U735 ( .A1(n1001), .A2(n1023), .ZN(n1022) );
NAND2_X1 U736 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND4_X1 U737 ( .A1(n1026), .A2(n1007), .A3(n1027), .A4(n1028), .ZN(n1025) );
XOR2_X1 U738 ( .A(KEYINPUT23), .B(n1008), .Z(n1028) );
NAND2_X1 U739 ( .A1(n1006), .A2(n1029), .ZN(n1024) );
NAND2_X1 U740 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U741 ( .A1(n1007), .A2(n1032), .ZN(n1031) );
NOR2_X1 U742 ( .A1(n1033), .A2(n1034), .ZN(n1007) );
NAND2_X1 U743 ( .A1(n1008), .A2(n1035), .ZN(n1030) );
NAND2_X1 U744 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U745 ( .A1(n1017), .A2(n1038), .A3(n1039), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1016), .A2(n1040), .ZN(n1036) );
INV_X1 U747 ( .A(n1041), .ZN(n1001) );
AND3_X1 U748 ( .A1(n1020), .A2(n1021), .A3(n1042), .ZN(n995) );
NAND4_X1 U749 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1020) );
NOR4_X1 U750 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
XOR2_X1 U751 ( .A(KEYINPUT13), .B(n1051), .Z(n1050) );
NOR2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U753 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U754 ( .A(KEYINPUT50), .B(n1056), .Z(n1055) );
NOR2_X1 U755 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
INV_X1 U756 ( .A(n1054), .ZN(n1057) );
XOR2_X1 U757 ( .A(n1058), .B(KEYINPUT40), .Z(n1056) );
XNOR2_X1 U758 ( .A(G469), .B(n1059), .ZN(n1049) );
XNOR2_X1 U759 ( .A(n1060), .B(n1061), .ZN(n1048) );
XOR2_X1 U760 ( .A(KEYINPUT52), .B(KEYINPUT25), .Z(n1061) );
XOR2_X1 U761 ( .A(n1062), .B(n1063), .Z(n1047) );
NOR2_X1 U762 ( .A1(G472), .A2(KEYINPUT45), .ZN(n1063) );
NOR3_X1 U763 ( .A1(n1064), .A2(n1065), .A3(n1026), .ZN(n1045) );
INV_X1 U764 ( .A(n1066), .ZN(n1064) );
XOR2_X1 U765 ( .A(n1067), .B(n1068), .Z(n1043) );
NAND2_X1 U766 ( .A1(KEYINPUT17), .A2(n1069), .ZN(n1068) );
XOR2_X1 U767 ( .A(n1070), .B(n1071), .Z(G72) );
XOR2_X1 U768 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U770 ( .A(n1076), .B(n1077), .Z(n1075) );
XNOR2_X1 U771 ( .A(n1078), .B(n1079), .ZN(n1077) );
XOR2_X1 U772 ( .A(n1080), .B(n1081), .Z(n1076) );
XNOR2_X1 U773 ( .A(G131), .B(G125), .ZN(n1081) );
NAND2_X1 U774 ( .A1(n1082), .A2(KEYINPUT39), .ZN(n1080) );
XNOR2_X1 U775 ( .A(n1083), .B(KEYINPUT12), .ZN(n1082) );
NOR2_X1 U776 ( .A1(G900), .A2(n1021), .ZN(n1074) );
NOR2_X1 U777 ( .A1(G953), .A2(n1084), .ZN(n1072) );
NOR2_X1 U778 ( .A1(n1085), .A2(n1021), .ZN(n1070) );
NOR2_X1 U779 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U780 ( .A(n1088), .B(n1089), .Z(G69) );
NOR2_X1 U781 ( .A1(KEYINPUT31), .A2(n1090), .ZN(n1089) );
XOR2_X1 U782 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U783 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U784 ( .A1(G953), .A2(n1095), .ZN(n1094) );
XOR2_X1 U785 ( .A(n1096), .B(n1097), .Z(n1093) );
NAND3_X1 U786 ( .A1(n1098), .A2(n1021), .A3(KEYINPUT22), .ZN(n1091) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U788 ( .A(KEYINPUT6), .B(n1101), .ZN(n1100) );
NAND2_X1 U789 ( .A1(G953), .A2(n1102), .ZN(n1088) );
NAND2_X1 U790 ( .A1(G898), .A2(G224), .ZN(n1102) );
NOR2_X1 U791 ( .A1(n1103), .A2(n1104), .ZN(G66) );
NOR3_X1 U792 ( .A1(n1054), .A2(n1105), .A3(n1106), .ZN(n1104) );
AND3_X1 U793 ( .A1(n1107), .A2(n1058), .A3(n1108), .ZN(n1106) );
NOR2_X1 U794 ( .A1(n1109), .A2(n1107), .ZN(n1105) );
AND2_X1 U795 ( .A1(n999), .A2(n1058), .ZN(n1109) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1110), .ZN(G63) );
XNOR2_X1 U797 ( .A(n1111), .B(n1112), .ZN(n1110) );
AND2_X1 U798 ( .A1(G478), .A2(n1108), .ZN(n1112) );
NOR3_X1 U799 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(G60) );
AND2_X1 U800 ( .A1(KEYINPUT11), .A2(n1103), .ZN(n1115) );
NOR3_X1 U801 ( .A1(KEYINPUT11), .A2(n1021), .A3(n1042), .ZN(n1114) );
INV_X1 U802 ( .A(G952), .ZN(n1042) );
XOR2_X1 U803 ( .A(n1116), .B(n1117), .Z(n1113) );
XOR2_X1 U804 ( .A(KEYINPUT27), .B(n1118), .Z(n1117) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U806 ( .A(G104), .B(n1121), .ZN(G6) );
NOR2_X1 U807 ( .A1(n1122), .A2(n1123), .ZN(G57) );
XOR2_X1 U808 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U809 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U810 ( .A(n1128), .B(n1129), .ZN(n1127) );
AND2_X1 U811 ( .A1(G472), .A2(n1108), .ZN(n1126) );
XNOR2_X1 U812 ( .A(n1130), .B(n1131), .ZN(n1124) );
NAND3_X1 U813 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1130) );
OR2_X1 U814 ( .A1(n1135), .A2(n1078), .ZN(n1134) );
NAND2_X1 U815 ( .A1(KEYINPUT55), .A2(n1136), .ZN(n1133) );
NAND2_X1 U816 ( .A1(n1135), .A2(n1137), .ZN(n1136) );
XNOR2_X1 U817 ( .A(KEYINPUT60), .B(n1078), .ZN(n1137) );
NAND2_X1 U818 ( .A1(n1138), .A2(n1139), .ZN(n1132) );
INV_X1 U819 ( .A(KEYINPUT55), .ZN(n1139) );
NAND2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NAND3_X1 U821 ( .A1(KEYINPUT60), .A2(n1135), .A3(n1078), .ZN(n1141) );
OR2_X1 U822 ( .A1(n1078), .A2(KEYINPUT60), .ZN(n1140) );
NOR2_X1 U823 ( .A1(G952), .A2(n1142), .ZN(n1122) );
XNOR2_X1 U824 ( .A(G953), .B(KEYINPUT18), .ZN(n1142) );
NOR2_X1 U825 ( .A1(n1103), .A2(n1143), .ZN(G54) );
XOR2_X1 U826 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U827 ( .A(n1146), .B(n1147), .ZN(n1145) );
AND2_X1 U828 ( .A1(G469), .A2(n1108), .ZN(n1146) );
INV_X1 U829 ( .A(n1120), .ZN(n1108) );
NAND2_X1 U830 ( .A1(n1148), .A2(n1149), .ZN(n1144) );
NAND2_X1 U831 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U832 ( .A(n1152), .B(n1153), .Z(n1150) );
NOR2_X1 U833 ( .A1(G110), .A2(n1154), .ZN(n1153) );
OR2_X1 U834 ( .A1(n1155), .A2(n1151), .ZN(n1148) );
INV_X1 U835 ( .A(KEYINPUT53), .ZN(n1151) );
NOR2_X1 U836 ( .A1(n1103), .A2(n1156), .ZN(G51) );
XOR2_X1 U837 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U838 ( .A(n1159), .B(n1160), .ZN(n1158) );
NAND2_X1 U839 ( .A1(KEYINPUT26), .A2(n1161), .ZN(n1159) );
OR2_X1 U840 ( .A1(n1120), .A2(n1069), .ZN(n1161) );
NAND2_X1 U841 ( .A1(G902), .A2(n999), .ZN(n1120) );
NAND3_X1 U842 ( .A1(n1099), .A2(n1101), .A3(n1084), .ZN(n999) );
AND4_X1 U843 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1084) );
AND4_X1 U844 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
NAND2_X1 U845 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
NAND2_X1 U846 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U847 ( .A(KEYINPUT33), .B(n1040), .Z(n1172) );
NAND3_X1 U848 ( .A1(n1174), .A2(n1016), .A3(n1175), .ZN(n1162) );
NAND2_X1 U849 ( .A1(n1176), .A2(n1177), .ZN(n1101) );
XNOR2_X1 U850 ( .A(KEYINPUT16), .B(n1178), .ZN(n1177) );
AND4_X1 U851 ( .A1(n1121), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1099) );
NOR3_X1 U852 ( .A1(n994), .A2(n1182), .A3(n1183), .ZN(n1181) );
NOR3_X1 U853 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1183) );
NAND3_X1 U854 ( .A1(n1187), .A2(n1188), .A3(n1017), .ZN(n1184) );
OR2_X1 U855 ( .A1(n1189), .A2(KEYINPUT47), .ZN(n1188) );
NAND2_X1 U856 ( .A1(KEYINPUT47), .A2(n1190), .ZN(n1187) );
NAND3_X1 U857 ( .A1(n1191), .A2(n1192), .A3(n1006), .ZN(n1190) );
AND2_X1 U858 ( .A1(n1032), .A2(n1193), .ZN(n994) );
NAND2_X1 U859 ( .A1(n1189), .A2(n1194), .ZN(n1180) );
NAND2_X1 U860 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U861 ( .A1(n1197), .A2(n1015), .ZN(n1195) );
XNOR2_X1 U862 ( .A(n1032), .B(KEYINPUT7), .ZN(n1197) );
NAND2_X1 U863 ( .A1(n1005), .A2(n1193), .ZN(n1121) );
AND3_X1 U864 ( .A1(n1178), .A2(n1017), .A3(n1198), .ZN(n1193) );
XNOR2_X1 U865 ( .A(G125), .B(n1199), .ZN(n1157) );
NOR2_X1 U866 ( .A1(n1021), .A2(G952), .ZN(n1103) );
XNOR2_X1 U867 ( .A(G146), .B(n1163), .ZN(G48) );
NAND3_X1 U868 ( .A1(n1200), .A2(n1005), .A3(n1174), .ZN(n1163) );
XNOR2_X1 U869 ( .A(G143), .B(n1169), .ZN(G45) );
NAND3_X1 U870 ( .A1(n1015), .A2(n1174), .A3(n1201), .ZN(n1169) );
NOR3_X1 U871 ( .A1(n1192), .A2(n1185), .A3(n1186), .ZN(n1201) );
INV_X1 U872 ( .A(n1018), .ZN(n1192) );
XOR2_X1 U873 ( .A(G140), .B(n1202), .Z(G42) );
AND2_X1 U874 ( .A1(n1040), .A2(n1170), .ZN(n1202) );
INV_X1 U875 ( .A(n1203), .ZN(n1170) );
XOR2_X1 U876 ( .A(n1204), .B(G137), .Z(G39) );
NAND2_X1 U877 ( .A1(KEYINPUT36), .A2(n1205), .ZN(n1204) );
NAND3_X1 U878 ( .A1(n1175), .A2(n1174), .A3(n1206), .ZN(n1205) );
XNOR2_X1 U879 ( .A(n1016), .B(KEYINPUT14), .ZN(n1206) );
XNOR2_X1 U880 ( .A(G134), .B(n1168), .ZN(G36) );
NAND4_X1 U881 ( .A1(n1015), .A2(n1174), .A3(n1016), .A4(n1032), .ZN(n1168) );
XNOR2_X1 U882 ( .A(n1207), .B(n1208), .ZN(G33) );
NOR2_X1 U883 ( .A1(n1173), .A2(n1203), .ZN(n1208) );
NAND3_X1 U884 ( .A1(n1016), .A2(n1005), .A3(n1174), .ZN(n1203) );
AND2_X1 U885 ( .A1(n1019), .A2(n1209), .ZN(n1174) );
INV_X1 U886 ( .A(n1033), .ZN(n1016) );
NAND2_X1 U887 ( .A1(n1038), .A2(n1044), .ZN(n1033) );
NAND2_X1 U888 ( .A1(n1210), .A2(n1211), .ZN(G30) );
OR2_X1 U889 ( .A1(n1167), .A2(G128), .ZN(n1211) );
XOR2_X1 U890 ( .A(n1212), .B(KEYINPUT4), .Z(n1210) );
NAND2_X1 U891 ( .A1(G128), .A2(n1167), .ZN(n1212) );
NAND4_X1 U892 ( .A1(n1200), .A2(n1032), .A3(n1178), .A4(n1209), .ZN(n1167) );
AND3_X1 U893 ( .A1(n1018), .A2(n1213), .A3(n1214), .ZN(n1200) );
NAND2_X1 U894 ( .A1(n1215), .A2(n1216), .ZN(G3) );
NAND2_X1 U895 ( .A1(n1217), .A2(n1128), .ZN(n1216) );
XOR2_X1 U896 ( .A(KEYINPUT61), .B(n1218), .Z(n1215) );
NOR2_X1 U897 ( .A1(n1217), .A2(n1128), .ZN(n1218) );
INV_X1 U898 ( .A(G101), .ZN(n1128) );
INV_X1 U899 ( .A(n1179), .ZN(n1217) );
NAND4_X1 U900 ( .A1(n1015), .A2(n1008), .A3(n1178), .A4(n1198), .ZN(n1179) );
XNOR2_X1 U901 ( .A(G125), .B(n1166), .ZN(G27) );
NAND3_X1 U902 ( .A1(n1005), .A2(n1006), .A3(n1219), .ZN(n1166) );
AND3_X1 U903 ( .A1(n1040), .A2(n1209), .A3(n1018), .ZN(n1219) );
NAND2_X1 U904 ( .A1(n1041), .A2(n1220), .ZN(n1209) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1087), .ZN(n1220) );
INV_X1 U906 ( .A(G900), .ZN(n1087) );
XOR2_X1 U907 ( .A(G122), .B(n1222), .Z(G24) );
NOR4_X1 U908 ( .A1(n1185), .A2(n1186), .A3(n1034), .A4(n1223), .ZN(n1222) );
INV_X1 U909 ( .A(n1017), .ZN(n1034) );
NOR2_X1 U910 ( .A1(n1213), .A2(n1214), .ZN(n1017) );
XNOR2_X1 U911 ( .A(G119), .B(n1224), .ZN(G21) );
NAND4_X1 U912 ( .A1(n1225), .A2(n1175), .A3(n1006), .A4(n1191), .ZN(n1224) );
INV_X1 U913 ( .A(n1196), .ZN(n1175) );
NAND3_X1 U914 ( .A1(n1214), .A2(n1213), .A3(n1008), .ZN(n1196) );
INV_X1 U915 ( .A(n1226), .ZN(n1214) );
XNOR2_X1 U916 ( .A(n1018), .B(KEYINPUT0), .ZN(n1225) );
XNOR2_X1 U917 ( .A(G116), .B(n1227), .ZN(G18) );
NAND4_X1 U918 ( .A1(KEYINPUT30), .A2(n1189), .A3(n1015), .A4(n1032), .ZN(n1227) );
NOR2_X1 U919 ( .A1(n1228), .A2(n1186), .ZN(n1032) );
INV_X1 U920 ( .A(n1060), .ZN(n1186) );
XOR2_X1 U921 ( .A(G113), .B(n1182), .Z(G15) );
AND3_X1 U922 ( .A1(n1015), .A2(n1005), .A3(n1189), .ZN(n1182) );
INV_X1 U923 ( .A(n1223), .ZN(n1189) );
NAND2_X1 U924 ( .A1(n1006), .A2(n1198), .ZN(n1223) );
NOR2_X1 U925 ( .A1(n1229), .A2(n1026), .ZN(n1006) );
NOR2_X1 U926 ( .A1(n1060), .A2(n1185), .ZN(n1005) );
INV_X1 U927 ( .A(n1228), .ZN(n1185) );
INV_X1 U928 ( .A(n1173), .ZN(n1015) );
NAND2_X1 U929 ( .A1(n1226), .A2(n1213), .ZN(n1173) );
XNOR2_X1 U930 ( .A(G110), .B(n1230), .ZN(G12) );
NAND2_X1 U931 ( .A1(n1176), .A2(n1178), .ZN(n1230) );
XNOR2_X1 U932 ( .A(n1019), .B(KEYINPUT51), .ZN(n1178) );
NOR2_X1 U933 ( .A1(n1027), .A2(n1026), .ZN(n1019) );
AND2_X1 U934 ( .A1(G221), .A2(n1231), .ZN(n1026) );
INV_X1 U935 ( .A(n1229), .ZN(n1027) );
NAND2_X1 U936 ( .A1(n1232), .A2(n1233), .ZN(n1229) );
NAND2_X1 U937 ( .A1(G469), .A2(n1059), .ZN(n1233) );
XOR2_X1 U938 ( .A(KEYINPUT37), .B(n1234), .Z(n1232) );
NOR2_X1 U939 ( .A1(G469), .A2(n1059), .ZN(n1234) );
NAND3_X1 U940 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1059) );
NAND2_X1 U941 ( .A1(n1238), .A2(n1239), .ZN(n1236) );
INV_X1 U942 ( .A(KEYINPUT10), .ZN(n1239) );
XOR2_X1 U943 ( .A(n1155), .B(n1147), .Z(n1238) );
NAND3_X1 U944 ( .A1(n1147), .A2(n1155), .A3(KEYINPUT10), .ZN(n1235) );
XOR2_X1 U945 ( .A(n1240), .B(n1154), .Z(n1155) );
XNOR2_X1 U946 ( .A(n1241), .B(KEYINPUT2), .ZN(n1154) );
XNOR2_X1 U947 ( .A(G110), .B(n1152), .ZN(n1240) );
NOR2_X1 U948 ( .A1(n1086), .A2(G953), .ZN(n1152) );
INV_X1 U949 ( .A(G227), .ZN(n1086) );
XNOR2_X1 U950 ( .A(n1242), .B(n1135), .ZN(n1147) );
XNOR2_X1 U951 ( .A(n1243), .B(KEYINPUT57), .ZN(n1242) );
AND3_X1 U952 ( .A1(n1040), .A2(n1198), .A3(n1008), .ZN(n1176) );
NOR2_X1 U953 ( .A1(n1060), .A2(n1228), .ZN(n1008) );
NAND2_X1 U954 ( .A1(n1244), .A2(n1066), .ZN(n1228) );
NAND3_X1 U955 ( .A1(n1119), .A2(n1237), .A3(n1116), .ZN(n1066) );
INV_X1 U956 ( .A(G475), .ZN(n1119) );
XOR2_X1 U957 ( .A(KEYINPUT41), .B(n1065), .Z(n1244) );
AND2_X1 U958 ( .A1(G475), .A2(n1245), .ZN(n1065) );
NAND2_X1 U959 ( .A1(n1116), .A2(n1237), .ZN(n1245) );
XNOR2_X1 U960 ( .A(n1246), .B(n1247), .ZN(n1116) );
XNOR2_X1 U961 ( .A(n1248), .B(n1249), .ZN(n1247) );
XOR2_X1 U962 ( .A(n1250), .B(n1251), .Z(n1249) );
AND3_X1 U963 ( .A1(G214), .A2(n1021), .A3(n1252), .ZN(n1251) );
NAND2_X1 U964 ( .A1(KEYINPUT54), .A2(n1207), .ZN(n1250) );
INV_X1 U965 ( .A(G131), .ZN(n1207) );
XOR2_X1 U966 ( .A(n1253), .B(n1254), .Z(n1246) );
XOR2_X1 U967 ( .A(G122), .B(G113), .Z(n1254) );
XOR2_X1 U968 ( .A(n1255), .B(G104), .Z(n1253) );
NAND2_X1 U969 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U970 ( .A1(G125), .A2(n1241), .ZN(n1257) );
XOR2_X1 U971 ( .A(KEYINPUT34), .B(n1258), .Z(n1256) );
NOR2_X1 U972 ( .A1(G125), .A2(n1241), .ZN(n1258) );
XNOR2_X1 U973 ( .A(n1259), .B(G478), .ZN(n1060) );
NAND2_X1 U974 ( .A1(n1111), .A2(n1237), .ZN(n1259) );
XNOR2_X1 U975 ( .A(n1260), .B(n1261), .ZN(n1111) );
XOR2_X1 U976 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U977 ( .A(n1264), .B(n1265), .ZN(n1263) );
AND4_X1 U978 ( .A1(n1266), .A2(n1021), .A3(G217), .A4(G234), .ZN(n1265) );
INV_X1 U979 ( .A(KEYINPUT29), .ZN(n1266) );
NAND2_X1 U980 ( .A1(KEYINPUT43), .A2(G116), .ZN(n1264) );
XOR2_X1 U981 ( .A(n1267), .B(n1268), .Z(n1260) );
XNOR2_X1 U982 ( .A(n1269), .B(G128), .ZN(n1268) );
INV_X1 U983 ( .A(G143), .ZN(n1269) );
XNOR2_X1 U984 ( .A(G107), .B(G122), .ZN(n1267) );
AND2_X1 U985 ( .A1(n1018), .A2(n1191), .ZN(n1198) );
NAND2_X1 U986 ( .A1(n1041), .A2(n1270), .ZN(n1191) );
NAND4_X1 U987 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1095), .ZN(n1270) );
INV_X1 U988 ( .A(G898), .ZN(n1095) );
NAND3_X1 U989 ( .A1(n1221), .A2(n1021), .A3(G952), .ZN(n1041) );
NAND2_X1 U990 ( .A1(G237), .A2(G234), .ZN(n1221) );
NOR2_X1 U991 ( .A1(n1038), .A2(n1039), .ZN(n1018) );
INV_X1 U992 ( .A(n1044), .ZN(n1039) );
NAND2_X1 U993 ( .A1(G214), .A2(n1271), .ZN(n1044) );
XOR2_X1 U994 ( .A(n1272), .B(n1067), .Z(n1038) );
NAND2_X1 U995 ( .A1(n1273), .A2(n1237), .ZN(n1067) );
XOR2_X1 U996 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U997 ( .A(n1276), .B(n1277), .ZN(n1275) );
INV_X1 U998 ( .A(n1160), .ZN(n1277) );
XOR2_X1 U999 ( .A(n1097), .B(n1243), .Z(n1160) );
XNOR2_X1 U1000 ( .A(n1096), .B(n1078), .ZN(n1243) );
INV_X1 U1001 ( .A(n1278), .ZN(n1078) );
XOR2_X1 U1002 ( .A(G101), .B(n1279), .Z(n1096) );
XOR2_X1 U1003 ( .A(G107), .B(G104), .Z(n1279) );
XNOR2_X1 U1004 ( .A(n1280), .B(n1281), .ZN(n1097) );
XOR2_X1 U1005 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U1006 ( .A(G119), .B(n1284), .ZN(n1283) );
XOR2_X1 U1007 ( .A(n1285), .B(n1286), .Z(n1280) );
XOR2_X1 U1008 ( .A(KEYINPUT24), .B(G122), .Z(n1286) );
XNOR2_X1 U1009 ( .A(KEYINPUT56), .B(KEYINPUT46), .ZN(n1285) );
NOR2_X1 U1010 ( .A1(G125), .A2(KEYINPUT28), .ZN(n1276) );
XOR2_X1 U1011 ( .A(n1287), .B(KEYINPUT59), .Z(n1274) );
NAND2_X1 U1012 ( .A1(KEYINPUT42), .A2(n1199), .ZN(n1287) );
NAND2_X1 U1013 ( .A1(G224), .A2(n1021), .ZN(n1199) );
NAND2_X1 U1014 ( .A1(n1288), .A2(KEYINPUT9), .ZN(n1272) );
XOR2_X1 U1015 ( .A(n1069), .B(KEYINPUT58), .Z(n1288) );
NAND2_X1 U1016 ( .A1(G210), .A2(n1271), .ZN(n1069) );
NAND2_X1 U1017 ( .A1(n1252), .A2(n1237), .ZN(n1271) );
NOR2_X1 U1018 ( .A1(n1226), .A2(n1213), .ZN(n1040) );
XNOR2_X1 U1019 ( .A(n1062), .B(G472), .ZN(n1213) );
NAND2_X1 U1020 ( .A1(n1289), .A2(n1237), .ZN(n1062) );
XOR2_X1 U1021 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U1022 ( .A(n1278), .B(n1135), .ZN(n1291) );
XNOR2_X1 U1023 ( .A(G131), .B(n1292), .ZN(n1135) );
NOR2_X1 U1024 ( .A1(KEYINPUT49), .A2(n1293), .ZN(n1292) );
XOR2_X1 U1025 ( .A(KEYINPUT38), .B(n1079), .Z(n1293) );
XOR2_X1 U1026 ( .A(G137), .B(n1262), .Z(n1079) );
XOR2_X1 U1027 ( .A(G134), .B(KEYINPUT48), .Z(n1262) );
XNOR2_X1 U1028 ( .A(n1294), .B(n1248), .ZN(n1278) );
XNOR2_X1 U1029 ( .A(G143), .B(n1295), .ZN(n1248) );
XNOR2_X1 U1030 ( .A(G128), .B(KEYINPUT62), .ZN(n1294) );
XOR2_X1 U1031 ( .A(n1296), .B(n1297), .Z(n1290) );
XNOR2_X1 U1032 ( .A(G101), .B(n1298), .ZN(n1297) );
NOR2_X1 U1033 ( .A1(KEYINPUT20), .A2(n1131), .ZN(n1298) );
XNOR2_X1 U1034 ( .A(n1282), .B(n1299), .ZN(n1131) );
NOR2_X1 U1035 ( .A1(KEYINPUT5), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1036 ( .A(KEYINPUT19), .B(G119), .Z(n1300) );
XOR2_X1 U1037 ( .A(G113), .B(G116), .Z(n1282) );
NAND2_X1 U1038 ( .A1(KEYINPUT35), .A2(n1129), .ZN(n1296) );
AND3_X1 U1039 ( .A1(n1252), .A2(n1021), .A3(G210), .ZN(n1129) );
INV_X1 U1040 ( .A(G237), .ZN(n1252) );
XNOR2_X1 U1041 ( .A(n1301), .B(n1302), .ZN(n1226) );
NOR2_X1 U1042 ( .A1(KEYINPUT44), .A2(n1058), .ZN(n1302) );
AND2_X1 U1043 ( .A1(G217), .A2(n1231), .ZN(n1058) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1237), .ZN(n1231) );
INV_X1 U1045 ( .A(G902), .ZN(n1237) );
XNOR2_X1 U1046 ( .A(n1054), .B(KEYINPUT15), .ZN(n1301) );
NOR2_X1 U1047 ( .A1(n1107), .A2(G902), .ZN(n1054) );
XNOR2_X1 U1048 ( .A(n1303), .B(n1304), .ZN(n1107) );
XOR2_X1 U1049 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1050 ( .A(G137), .B(n1284), .ZN(n1306) );
INV_X1 U1051 ( .A(G110), .ZN(n1284) );
NOR2_X1 U1052 ( .A1(KEYINPUT32), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1053 ( .A(G128), .B(G119), .Z(n1307) );
XOR2_X1 U1054 ( .A(n1308), .B(n1309), .Z(n1303) );
AND3_X1 U1055 ( .A1(G221), .A2(n1021), .A3(G234), .ZN(n1309) );
INV_X1 U1056 ( .A(G953), .ZN(n1021) );
NAND2_X1 U1057 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
NAND2_X1 U1058 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
XOR2_X1 U1059 ( .A(KEYINPUT3), .B(n1314), .Z(n1310) );
NOR2_X1 U1060 ( .A1(n1312), .A2(n1313), .ZN(n1314) );
XNOR2_X1 U1061 ( .A(KEYINPUT63), .B(n1295), .ZN(n1313) );
INV_X1 U1062 ( .A(G146), .ZN(n1295) );
XNOR2_X1 U1063 ( .A(n1315), .B(n1241), .ZN(n1312) );
INV_X1 U1064 ( .A(n1083), .ZN(n1241) );
XOR2_X1 U1065 ( .A(G140), .B(KEYINPUT8), .Z(n1083) );
NAND2_X1 U1066 ( .A1(KEYINPUT1), .A2(n1316), .ZN(n1315) );
INV_X1 U1067 ( .A(G125), .ZN(n1316) );
endmodule


