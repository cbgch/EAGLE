//Key = 1011011000000000010011000101001110101100001000100111010100110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344;

XNOR2_X1 U732 ( .A(G107), .B(n1021), .ZN(G9) );
NOR2_X1 U733 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U734 ( .A1(n1024), .A2(n1025), .A3(KEYINPUT41), .A4(G953), .ZN(n1023) );
NAND2_X1 U735 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NAND2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND3_X1 U738 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND2_X1 U739 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NAND2_X1 U740 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U742 ( .A1(n1041), .A2(n1042), .ZN(n1035) );
NAND2_X1 U743 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U744 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U745 ( .A1(n1037), .A2(n1047), .A3(n1041), .ZN(n1030) );
NAND2_X1 U746 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U747 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
OR2_X1 U748 ( .A1(n1053), .A2(n1032), .ZN(n1051) );
OR3_X1 U749 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1050) );
NAND2_X1 U750 ( .A1(n1057), .A2(n1032), .ZN(n1048) );
INV_X1 U751 ( .A(n1058), .ZN(n1028) );
NOR3_X1 U752 ( .A1(n1025), .A2(G953), .A3(G952), .ZN(n1022) );
AND4_X1 U753 ( .A1(n1059), .A2(n1037), .A3(n1034), .A4(n1060), .ZN(n1025) );
NOR4_X1 U754 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
XOR2_X1 U755 ( .A(n1065), .B(G478), .Z(n1064) );
NAND2_X1 U756 ( .A1(n1066), .A2(KEYINPUT55), .ZN(n1065) );
XNOR2_X1 U757 ( .A(n1067), .B(KEYINPUT12), .ZN(n1066) );
XOR2_X1 U758 ( .A(n1068), .B(G472), .Z(n1063) );
NAND2_X1 U759 ( .A1(n1069), .A2(KEYINPUT5), .ZN(n1068) );
XOR2_X1 U760 ( .A(n1070), .B(KEYINPUT22), .Z(n1069) );
NOR2_X1 U761 ( .A1(n1071), .A2(n1072), .ZN(n1062) );
XOR2_X1 U762 ( .A(KEYINPUT53), .B(n1073), .Z(n1072) );
NOR2_X1 U763 ( .A1(G902), .A2(n1074), .ZN(n1071) );
NAND2_X1 U764 ( .A1(n1075), .A2(n1076), .ZN(G72) );
NAND3_X1 U765 ( .A1(KEYINPUT21), .A2(n1077), .A3(n1078), .ZN(n1076) );
NAND2_X1 U766 ( .A1(n1079), .A2(n1080), .ZN(n1075) );
NAND2_X1 U767 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U768 ( .A1(n1077), .A2(n1083), .ZN(n1082) );
INV_X1 U769 ( .A(KEYINPUT59), .ZN(n1083) );
NAND2_X1 U770 ( .A1(KEYINPUT59), .A2(n1084), .ZN(n1081) );
NAND2_X1 U771 ( .A1(KEYINPUT21), .A2(n1077), .ZN(n1084) );
AND2_X1 U772 ( .A1(n1085), .A2(n1086), .ZN(n1077) );
NAND2_X1 U773 ( .A1(G900), .A2(G227), .ZN(n1086) );
XOR2_X1 U774 ( .A(KEYINPUT57), .B(G953), .Z(n1085) );
INV_X1 U775 ( .A(n1078), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1087), .A2(n1088), .ZN(n1078) );
NAND2_X1 U777 ( .A1(G953), .A2(n1089), .ZN(n1088) );
XOR2_X1 U778 ( .A(n1090), .B(n1091), .Z(n1087) );
XOR2_X1 U779 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U780 ( .A(KEYINPUT0), .B(G131), .Z(n1093) );
NOR2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
XNOR2_X1 U782 ( .A(n1096), .B(n1097), .ZN(n1090) );
XNOR2_X1 U783 ( .A(n1098), .B(n1099), .ZN(n1096) );
NOR2_X1 U784 ( .A1(KEYINPUT11), .A2(n1100), .ZN(n1099) );
XOR2_X1 U785 ( .A(n1101), .B(n1102), .Z(G69) );
NAND2_X1 U786 ( .A1(G953), .A2(n1103), .ZN(n1102) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1103) );
NAND2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
OR2_X1 U791 ( .A1(n1110), .A2(KEYINPUT38), .ZN(n1109) );
INV_X1 U792 ( .A(n1111), .ZN(n1106) );
NAND2_X1 U793 ( .A1(n1112), .A2(n1110), .ZN(n1104) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NAND2_X1 U795 ( .A1(G953), .A2(n1115), .ZN(n1114) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1113) );
NAND2_X1 U797 ( .A1(KEYINPUT3), .A2(n1118), .ZN(n1116) );
NAND2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1112) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1108), .ZN(n1120) );
INV_X1 U800 ( .A(KEYINPUT35), .ZN(n1108) );
NAND2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1111) );
NAND3_X1 U802 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
XNOR2_X1 U803 ( .A(n1126), .B(KEYINPUT33), .ZN(n1125) );
INV_X1 U804 ( .A(n1127), .ZN(n1123) );
INV_X1 U805 ( .A(KEYINPUT38), .ZN(n1119) );
NOR2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XNOR2_X1 U807 ( .A(n1074), .B(n1130), .ZN(n1129) );
XOR2_X1 U808 ( .A(KEYINPUT17), .B(n1131), .Z(n1130) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U810 ( .A1(n1128), .A2(n1134), .ZN(G63) );
NOR3_X1 U811 ( .A1(n1067), .A2(n1135), .A3(n1136), .ZN(n1134) );
NOR3_X1 U812 ( .A1(n1137), .A2(n1138), .A3(n1133), .ZN(n1136) );
NOR2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1026), .A2(n1138), .ZN(n1139) );
INV_X1 U815 ( .A(G478), .ZN(n1138) );
INV_X1 U816 ( .A(n1141), .ZN(n1026) );
NOR2_X1 U817 ( .A1(n1142), .A2(n1143), .ZN(G60) );
XOR2_X1 U818 ( .A(KEYINPUT45), .B(n1128), .Z(n1143) );
NOR2_X1 U819 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U821 ( .A1(n1148), .A2(n1133), .ZN(n1147) );
INV_X1 U822 ( .A(G475), .ZN(n1148) );
NOR2_X1 U823 ( .A1(KEYINPUT15), .A2(n1149), .ZN(n1146) );
AND2_X1 U824 ( .A1(n1149), .A2(KEYINPUT15), .ZN(n1144) );
XNOR2_X1 U825 ( .A(G104), .B(n1150), .ZN(G6) );
NOR2_X1 U826 ( .A1(n1128), .A2(n1151), .ZN(G57) );
XOR2_X1 U827 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U828 ( .A(n1154), .B(n1155), .ZN(n1153) );
XOR2_X1 U829 ( .A(n1156), .B(n1157), .Z(n1152) );
XNOR2_X1 U830 ( .A(G101), .B(n1158), .ZN(n1157) );
NOR2_X1 U831 ( .A1(n1159), .A2(KEYINPUT52), .ZN(n1158) );
NOR2_X1 U832 ( .A1(n1160), .A2(n1133), .ZN(n1159) );
NAND2_X1 U833 ( .A1(KEYINPUT62), .A2(n1161), .ZN(n1156) );
NOR2_X1 U834 ( .A1(n1128), .A2(n1162), .ZN(G54) );
XOR2_X1 U835 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U836 ( .A(n1097), .B(n1165), .ZN(n1164) );
XOR2_X1 U837 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U838 ( .A(n1168), .B(n1169), .Z(n1163) );
XOR2_X1 U839 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XNOR2_X1 U841 ( .A(n1174), .B(KEYINPUT9), .ZN(n1172) );
NOR2_X1 U842 ( .A1(n1175), .A2(n1133), .ZN(n1168) );
NOR2_X1 U843 ( .A1(n1128), .A2(n1176), .ZN(G51) );
XOR2_X1 U844 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U845 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U846 ( .A(G125), .B(n1181), .Z(n1180) );
NOR2_X1 U847 ( .A1(n1182), .A2(n1133), .ZN(n1179) );
NAND2_X1 U848 ( .A1(G902), .A2(n1141), .ZN(n1133) );
NAND4_X1 U849 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1141) );
INV_X1 U850 ( .A(n1095), .ZN(n1186) );
NAND4_X1 U851 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1095) );
NAND3_X1 U852 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1187) );
NOR2_X1 U853 ( .A1(n1126), .A2(n1127), .ZN(n1185) );
NAND4_X1 U854 ( .A1(n1150), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1127) );
AND3_X1 U855 ( .A1(n1197), .A2(n1021), .A3(n1198), .ZN(n1196) );
NAND3_X1 U856 ( .A1(n1199), .A2(n1032), .A3(n1200), .ZN(n1021) );
NAND3_X1 U857 ( .A1(n1201), .A2(n1054), .A3(n1191), .ZN(n1195) );
NAND3_X1 U858 ( .A1(n1200), .A2(n1032), .A3(n1191), .ZN(n1150) );
XOR2_X1 U859 ( .A(n1094), .B(KEYINPUT49), .Z(n1184) );
NAND4_X1 U860 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1094) );
NAND2_X1 U861 ( .A1(n1206), .A2(n1037), .ZN(n1202) );
INV_X1 U862 ( .A(n1207), .ZN(n1206) );
XOR2_X1 U863 ( .A(n1124), .B(KEYINPUT24), .Z(n1183) );
XOR2_X1 U864 ( .A(n1208), .B(n1209), .Z(n1177) );
NOR2_X1 U865 ( .A1(KEYINPUT43), .A2(n1210), .ZN(n1209) );
NOR2_X1 U866 ( .A1(n1211), .A2(G952), .ZN(n1128) );
XOR2_X1 U867 ( .A(G953), .B(KEYINPUT6), .Z(n1211) );
XOR2_X1 U868 ( .A(n1212), .B(n1213), .Z(G48) );
NAND4_X1 U869 ( .A1(n1214), .A2(n1191), .A3(n1215), .A4(n1192), .ZN(n1213) );
NOR2_X1 U870 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U871 ( .A(n1218), .B(KEYINPUT39), .Z(n1217) );
XOR2_X1 U872 ( .A(n1043), .B(KEYINPUT50), .Z(n1214) );
XNOR2_X1 U873 ( .A(G143), .B(n1188), .ZN(G45) );
NAND4_X1 U874 ( .A1(n1193), .A2(n1054), .A3(n1219), .A4(n1220), .ZN(n1188) );
NAND2_X1 U875 ( .A1(n1221), .A2(n1222), .ZN(G42) );
NAND2_X1 U876 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XNOR2_X1 U877 ( .A(KEYINPUT29), .B(n1189), .ZN(n1224) );
XOR2_X1 U878 ( .A(KEYINPUT51), .B(G140), .Z(n1223) );
XOR2_X1 U879 ( .A(n1225), .B(KEYINPUT60), .Z(n1221) );
NAND2_X1 U880 ( .A1(G140), .A2(n1189), .ZN(n1225) );
NAND3_X1 U881 ( .A1(n1226), .A2(n1055), .A3(n1191), .ZN(n1189) );
XNOR2_X1 U882 ( .A(G137), .B(n1190), .ZN(G39) );
NAND3_X1 U883 ( .A1(n1226), .A2(n1192), .A3(n1041), .ZN(n1190) );
XNOR2_X1 U884 ( .A(G134), .B(n1203), .ZN(G36) );
NAND3_X1 U885 ( .A1(n1054), .A2(n1199), .A3(n1226), .ZN(n1203) );
XOR2_X1 U886 ( .A(n1227), .B(n1204), .Z(G33) );
NAND3_X1 U887 ( .A1(n1226), .A2(n1054), .A3(n1191), .ZN(n1204) );
AND3_X1 U888 ( .A1(n1228), .A2(n1229), .A3(n1034), .ZN(n1226) );
AND2_X1 U889 ( .A1(n1052), .A2(n1053), .ZN(n1034) );
XOR2_X1 U890 ( .A(n1205), .B(n1230), .Z(G30) );
XOR2_X1 U891 ( .A(KEYINPUT2), .B(G128), .Z(n1230) );
NAND3_X1 U892 ( .A1(n1192), .A2(n1199), .A3(n1193), .ZN(n1205) );
NOR3_X1 U893 ( .A1(n1218), .A2(n1216), .A3(n1043), .ZN(n1193) );
INV_X1 U894 ( .A(n1228), .ZN(n1043) );
INV_X1 U895 ( .A(n1229), .ZN(n1216) );
XNOR2_X1 U896 ( .A(G101), .B(n1124), .ZN(G3) );
NAND3_X1 U897 ( .A1(n1054), .A2(n1200), .A3(n1041), .ZN(n1124) );
XOR2_X1 U898 ( .A(G125), .B(n1231), .Z(G27) );
NOR2_X1 U899 ( .A1(n1232), .A2(n1207), .ZN(n1231) );
NAND4_X1 U900 ( .A1(n1191), .A2(n1055), .A3(n1057), .A4(n1229), .ZN(n1207) );
NAND2_X1 U901 ( .A1(n1058), .A2(n1233), .ZN(n1229) );
NAND4_X1 U902 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1089), .ZN(n1233) );
INV_X1 U903 ( .A(G900), .ZN(n1089) );
XNOR2_X1 U904 ( .A(n1037), .B(KEYINPUT16), .ZN(n1232) );
XNOR2_X1 U905 ( .A(G122), .B(n1194), .ZN(G24) );
NAND4_X1 U906 ( .A1(n1201), .A2(n1032), .A3(n1219), .A4(n1220), .ZN(n1194) );
NAND2_X1 U907 ( .A1(n1235), .A2(n1236), .ZN(n1032) );
NAND3_X1 U908 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1236) );
INV_X1 U909 ( .A(KEYINPUT56), .ZN(n1239) );
NAND2_X1 U910 ( .A1(KEYINPUT56), .A2(n1055), .ZN(n1235) );
XOR2_X1 U911 ( .A(n1240), .B(n1197), .Z(G21) );
NAND3_X1 U912 ( .A1(n1192), .A2(n1201), .A3(n1041), .ZN(n1197) );
INV_X1 U913 ( .A(n1241), .ZN(n1201) );
NOR2_X1 U914 ( .A1(n1238), .A2(n1237), .ZN(n1192) );
XOR2_X1 U915 ( .A(n1242), .B(n1243), .Z(G18) );
NOR2_X1 U916 ( .A1(n1126), .A2(KEYINPUT23), .ZN(n1243) );
NOR3_X1 U917 ( .A1(n1244), .A2(n1040), .A3(n1241), .ZN(n1126) );
INV_X1 U918 ( .A(n1199), .ZN(n1040) );
NOR2_X1 U919 ( .A1(n1220), .A2(n1245), .ZN(n1199) );
XNOR2_X1 U920 ( .A(G113), .B(n1246), .ZN(G15) );
NAND4_X1 U921 ( .A1(n1191), .A2(n1054), .A3(n1247), .A4(n1248), .ZN(n1246) );
NAND2_X1 U922 ( .A1(KEYINPUT46), .A2(n1241), .ZN(n1248) );
NAND3_X1 U923 ( .A1(n1057), .A2(n1249), .A3(n1037), .ZN(n1241) );
NAND2_X1 U924 ( .A1(n1250), .A2(n1251), .ZN(n1247) );
INV_X1 U925 ( .A(KEYINPUT46), .ZN(n1251) );
NAND3_X1 U926 ( .A1(n1249), .A2(n1218), .A3(n1037), .ZN(n1250) );
NOR2_X1 U927 ( .A1(n1252), .A2(n1045), .ZN(n1037) );
INV_X1 U928 ( .A(n1046), .ZN(n1252) );
INV_X1 U929 ( .A(n1057), .ZN(n1218) );
INV_X1 U930 ( .A(n1244), .ZN(n1054) );
NAND2_X1 U931 ( .A1(n1253), .A2(n1254), .ZN(n1244) );
XOR2_X1 U932 ( .A(KEYINPUT56), .B(n1237), .Z(n1254) );
INV_X1 U933 ( .A(n1039), .ZN(n1191) );
NAND2_X1 U934 ( .A1(n1245), .A2(n1220), .ZN(n1039) );
INV_X1 U935 ( .A(n1219), .ZN(n1245) );
XNOR2_X1 U936 ( .A(n1198), .B(n1255), .ZN(G12) );
NOR2_X1 U937 ( .A1(KEYINPUT28), .A2(n1256), .ZN(n1255) );
NAND3_X1 U938 ( .A1(n1200), .A2(n1055), .A3(n1041), .ZN(n1198) );
NOR2_X1 U939 ( .A1(n1219), .A2(n1220), .ZN(n1041) );
XNOR2_X1 U940 ( .A(n1059), .B(KEYINPUT40), .ZN(n1220) );
XOR2_X1 U941 ( .A(n1257), .B(G475), .Z(n1059) );
OR2_X1 U942 ( .A1(n1149), .A2(G902), .ZN(n1257) );
XOR2_X1 U943 ( .A(n1258), .B(n1259), .Z(n1149) );
XOR2_X1 U944 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U945 ( .A1(KEYINPUT19), .A2(n1262), .ZN(n1260) );
NOR2_X1 U946 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U947 ( .A(n1265), .B(KEYINPUT42), .Z(n1264) );
NAND2_X1 U948 ( .A1(n1266), .A2(n1227), .ZN(n1265) );
NOR2_X1 U949 ( .A1(n1227), .A2(n1266), .ZN(n1263) );
XNOR2_X1 U950 ( .A(n1267), .B(G143), .ZN(n1266) );
NAND3_X1 U951 ( .A1(n1268), .A2(n1121), .A3(G214), .ZN(n1267) );
XOR2_X1 U952 ( .A(KEYINPUT27), .B(G237), .Z(n1268) );
XNOR2_X1 U953 ( .A(G104), .B(n1269), .ZN(n1258) );
XOR2_X1 U954 ( .A(G122), .B(G113), .Z(n1269) );
XOR2_X1 U955 ( .A(n1067), .B(G478), .Z(n1219) );
NOR2_X1 U956 ( .A1(n1140), .A2(G902), .ZN(n1067) );
INV_X1 U957 ( .A(n1137), .ZN(n1140) );
XOR2_X1 U958 ( .A(n1270), .B(n1271), .Z(n1137) );
XOR2_X1 U959 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U960 ( .A(n1274), .B(n1275), .Z(n1270) );
NOR2_X1 U961 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
INV_X1 U962 ( .A(G217), .ZN(n1277) );
XOR2_X1 U963 ( .A(n1278), .B(G107), .Z(n1274) );
NAND3_X1 U964 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1278) );
OR2_X1 U965 ( .A1(G122), .A2(KEYINPUT30), .ZN(n1281) );
NAND3_X1 U966 ( .A1(KEYINPUT30), .A2(G122), .A3(n1242), .ZN(n1280) );
INV_X1 U967 ( .A(G116), .ZN(n1242) );
NAND2_X1 U968 ( .A1(G116), .A2(n1282), .ZN(n1279) );
NAND2_X1 U969 ( .A1(n1283), .A2(KEYINPUT30), .ZN(n1282) );
XNOR2_X1 U970 ( .A(G122), .B(KEYINPUT58), .ZN(n1283) );
NOR2_X1 U971 ( .A1(n1253), .A2(n1237), .ZN(n1055) );
NOR2_X1 U972 ( .A1(n1061), .A2(n1284), .ZN(n1237) );
AND2_X1 U973 ( .A1(n1073), .A2(n1285), .ZN(n1284) );
OR2_X1 U974 ( .A1(n1074), .A2(G902), .ZN(n1285) );
NOR3_X1 U975 ( .A1(n1073), .A2(G902), .A3(n1074), .ZN(n1061) );
XOR2_X1 U976 ( .A(n1286), .B(n1287), .Z(n1074) );
XOR2_X1 U977 ( .A(G137), .B(n1288), .Z(n1287) );
NOR3_X1 U978 ( .A1(KEYINPUT54), .A2(n1289), .A3(n1290), .ZN(n1288) );
NOR3_X1 U979 ( .A1(G110), .A2(n1291), .A3(n1292), .ZN(n1290) );
NOR2_X1 U980 ( .A1(n1293), .A2(n1256), .ZN(n1289) );
NOR2_X1 U981 ( .A1(n1291), .A2(n1292), .ZN(n1293) );
XNOR2_X1 U982 ( .A(n1294), .B(KEYINPUT14), .ZN(n1292) );
NAND2_X1 U983 ( .A1(G128), .A2(n1240), .ZN(n1294) );
NOR2_X1 U984 ( .A1(n1240), .A2(G128), .ZN(n1291) );
INV_X1 U985 ( .A(G119), .ZN(n1240) );
XNOR2_X1 U986 ( .A(n1261), .B(n1295), .ZN(n1286) );
NOR2_X1 U987 ( .A1(n1296), .A2(n1276), .ZN(n1295) );
NAND2_X1 U988 ( .A1(G234), .A2(n1121), .ZN(n1276) );
INV_X1 U989 ( .A(G221), .ZN(n1296) );
XNOR2_X1 U990 ( .A(n1212), .B(n1098), .ZN(n1261) );
XOR2_X1 U991 ( .A(G125), .B(G140), .Z(n1098) );
INV_X1 U992 ( .A(n1132), .ZN(n1073) );
NAND2_X1 U993 ( .A1(G217), .A2(n1297), .ZN(n1132) );
INV_X1 U994 ( .A(n1238), .ZN(n1253) );
NAND3_X1 U995 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1238) );
NAND2_X1 U996 ( .A1(KEYINPUT44), .A2(G472), .ZN(n1300) );
NAND3_X1 U997 ( .A1(n1301), .A2(n1302), .A3(n1070), .ZN(n1299) );
INV_X1 U998 ( .A(KEYINPUT44), .ZN(n1302) );
OR2_X1 U999 ( .A1(n1070), .A2(n1301), .ZN(n1298) );
AND2_X1 U1000 ( .A1(n1303), .A2(n1160), .ZN(n1301) );
INV_X1 U1001 ( .A(G472), .ZN(n1160) );
XNOR2_X1 U1002 ( .A(KEYINPUT36), .B(KEYINPUT32), .ZN(n1303) );
NAND2_X1 U1003 ( .A1(n1304), .A2(n1305), .ZN(n1070) );
XOR2_X1 U1004 ( .A(n1306), .B(n1307), .Z(n1304) );
XNOR2_X1 U1005 ( .A(n1308), .B(n1154), .ZN(n1307) );
XNOR2_X1 U1006 ( .A(n1309), .B(KEYINPUT63), .ZN(n1154) );
NAND2_X1 U1007 ( .A1(KEYINPUT20), .A2(n1155), .ZN(n1308) );
XOR2_X1 U1008 ( .A(n1210), .B(n1310), .Z(n1155) );
INV_X1 U1009 ( .A(n1166), .ZN(n1310) );
XOR2_X1 U1010 ( .A(n1161), .B(n1311), .Z(n1306) );
XNOR2_X1 U1011 ( .A(G101), .B(KEYINPUT26), .ZN(n1311) );
NAND3_X1 U1012 ( .A1(n1312), .A2(n1121), .A3(G210), .ZN(n1161) );
AND3_X1 U1013 ( .A1(n1057), .A2(n1249), .A3(n1228), .ZN(n1200) );
NOR2_X1 U1014 ( .A1(n1046), .A2(n1045), .ZN(n1228) );
AND2_X1 U1015 ( .A1(G221), .A2(n1297), .ZN(n1045) );
NAND2_X1 U1016 ( .A1(G234), .A2(n1305), .ZN(n1297) );
XOR2_X1 U1017 ( .A(n1175), .B(n1313), .Z(n1046) );
NOR2_X1 U1018 ( .A1(G902), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1019 ( .A(n1315), .B(n1316), .Z(n1314) );
NOR3_X1 U1020 ( .A1(n1317), .A2(KEYINPUT1), .A3(n1318), .ZN(n1316) );
AND2_X1 U1021 ( .A1(n1319), .A2(n1166), .ZN(n1318) );
XOR2_X1 U1022 ( .A(KEYINPUT18), .B(n1320), .Z(n1317) );
NOR2_X1 U1023 ( .A1(n1166), .A2(n1319), .ZN(n1320) );
XNOR2_X1 U1024 ( .A(n1321), .B(n1322), .ZN(n1319) );
NOR2_X1 U1025 ( .A1(KEYINPUT48), .A2(n1097), .ZN(n1322) );
XOR2_X1 U1026 ( .A(n1323), .B(n1324), .Z(n1097) );
NOR2_X1 U1027 ( .A1(KEYINPUT7), .A2(n1212), .ZN(n1324) );
XOR2_X1 U1028 ( .A(n1227), .B(n1100), .Z(n1166) );
XNOR2_X1 U1029 ( .A(G137), .B(n1273), .ZN(n1100) );
XOR2_X1 U1030 ( .A(G134), .B(KEYINPUT13), .Z(n1273) );
INV_X1 U1031 ( .A(G131), .ZN(n1227) );
NOR2_X1 U1032 ( .A1(n1325), .A2(n1326), .ZN(n1315) );
XOR2_X1 U1033 ( .A(KEYINPUT8), .B(n1327), .Z(n1326) );
NOR3_X1 U1034 ( .A1(n1170), .A2(n1174), .A3(n1328), .ZN(n1327) );
NOR2_X1 U1035 ( .A1(n1329), .A2(n1330), .ZN(n1325) );
INV_X1 U1036 ( .A(n1170), .ZN(n1330) );
NAND2_X1 U1037 ( .A1(G227), .A2(n1121), .ZN(n1170) );
NOR2_X1 U1038 ( .A1(n1174), .A2(n1328), .ZN(n1329) );
INV_X1 U1039 ( .A(n1173), .ZN(n1328) );
NAND2_X1 U1040 ( .A1(G140), .A2(n1256), .ZN(n1173) );
NOR2_X1 U1041 ( .A1(n1256), .A2(G140), .ZN(n1174) );
INV_X1 U1042 ( .A(G110), .ZN(n1256) );
INV_X1 U1043 ( .A(G469), .ZN(n1175) );
NAND2_X1 U1044 ( .A1(n1331), .A2(n1058), .ZN(n1249) );
NAND3_X1 U1045 ( .A1(n1234), .A2(n1121), .A3(G952), .ZN(n1058) );
NAND4_X1 U1046 ( .A1(G953), .A2(G902), .A3(n1115), .A4(n1234), .ZN(n1331) );
NAND2_X1 U1047 ( .A1(G237), .A2(G234), .ZN(n1234) );
XOR2_X1 U1048 ( .A(KEYINPUT34), .B(G898), .Z(n1115) );
NOR2_X1 U1049 ( .A1(n1052), .A2(n1056), .ZN(n1057) );
INV_X1 U1050 ( .A(n1053), .ZN(n1056) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1332), .ZN(n1053) );
XNOR2_X1 U1052 ( .A(n1333), .B(n1182), .ZN(n1052) );
NAND2_X1 U1053 ( .A1(G210), .A2(n1332), .ZN(n1182) );
NAND2_X1 U1054 ( .A1(n1312), .A2(n1305), .ZN(n1332) );
INV_X1 U1055 ( .A(G237), .ZN(n1312) );
NAND2_X1 U1056 ( .A1(n1334), .A2(n1305), .ZN(n1333) );
INV_X1 U1057 ( .A(G902), .ZN(n1305) );
XOR2_X1 U1058 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U1059 ( .A(n1208), .B(n1337), .Z(n1336) );
XNOR2_X1 U1060 ( .A(n1210), .B(n1181), .ZN(n1337) );
AND2_X1 U1061 ( .A1(G224), .A2(n1121), .ZN(n1181) );
INV_X1 U1062 ( .A(G953), .ZN(n1121) );
XOR2_X1 U1063 ( .A(n1212), .B(n1323), .Z(n1210) );
XNOR2_X1 U1064 ( .A(n1272), .B(KEYINPUT10), .ZN(n1323) );
XOR2_X1 U1065 ( .A(G143), .B(G128), .Z(n1272) );
INV_X1 U1066 ( .A(G146), .ZN(n1212) );
XOR2_X1 U1067 ( .A(n1117), .B(n1118), .Z(n1208) );
XNOR2_X1 U1068 ( .A(n1309), .B(KEYINPUT37), .ZN(n1118) );
XNOR2_X1 U1069 ( .A(G113), .B(n1338), .ZN(n1309) );
XOR2_X1 U1070 ( .A(G119), .B(G116), .Z(n1338) );
XOR2_X1 U1071 ( .A(n1339), .B(n1340), .Z(n1117) );
XOR2_X1 U1072 ( .A(KEYINPUT31), .B(G110), .Z(n1340) );
XOR2_X1 U1073 ( .A(n1341), .B(n1167), .Z(n1339) );
INV_X1 U1074 ( .A(n1321), .ZN(n1167) );
XNOR2_X1 U1075 ( .A(G101), .B(n1342), .ZN(n1321) );
XOR2_X1 U1076 ( .A(G107), .B(G104), .Z(n1342) );
NAND2_X1 U1077 ( .A1(n1343), .A2(KEYINPUT25), .ZN(n1341) );
XNOR2_X1 U1078 ( .A(G122), .B(KEYINPUT4), .ZN(n1343) );
XNOR2_X1 U1079 ( .A(G125), .B(n1344), .ZN(n1335) );
XNOR2_X1 U1080 ( .A(KEYINPUT61), .B(KEYINPUT47), .ZN(n1344) );
endmodule


