//Key = 1011010111111010100000110001010010010011100101011110011111000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;

XNOR2_X1 U758 ( .A(n1038), .B(n1039), .ZN(G9) );
NOR2_X1 U759 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U760 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U761 ( .A1(G953), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1043) );
INV_X1 U762 ( .A(n1047), .ZN(n1046) );
NOR2_X1 U763 ( .A1(n1048), .A2(n1049), .ZN(n1045) );
NOR2_X1 U764 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR3_X1 U765 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
NOR3_X1 U766 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR2_X1 U767 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U768 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U769 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U770 ( .A1(n1064), .A2(n1065), .ZN(n1056) );
NOR2_X1 U771 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U772 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U773 ( .A1(n1070), .A2(n1071), .ZN(n1053) );
NOR3_X1 U774 ( .A1(n1065), .A2(n1072), .A3(n1059), .ZN(n1071) );
NOR4_X1 U775 ( .A1(n1073), .A2(n1055), .A3(n1059), .A4(n1065), .ZN(n1050) );
NOR2_X1 U776 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR3_X1 U777 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n1042) );
AND4_X1 U778 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1044) );
NOR3_X1 U779 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
XOR2_X1 U780 ( .A(n1083), .B(n1084), .Z(n1081) );
NOR2_X1 U781 ( .A1(KEYINPUT52), .A2(n1085), .ZN(n1084) );
XNOR2_X1 U782 ( .A(G469), .B(KEYINPUT48), .ZN(n1085) );
NAND3_X1 U783 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1080) );
XOR2_X1 U784 ( .A(n1089), .B(n1090), .Z(n1088) );
XNOR2_X1 U785 ( .A(n1091), .B(n1092), .ZN(n1090) );
XNOR2_X1 U786 ( .A(KEYINPUT24), .B(KEYINPUT18), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1093), .A2(n1094), .ZN(n1087) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
OR2_X1 U789 ( .A1(n1097), .A2(KEYINPUT6), .ZN(n1096) );
NAND2_X1 U790 ( .A1(n1098), .A2(n1097), .ZN(n1095) );
NAND2_X1 U791 ( .A1(KEYINPUT12), .A2(n1099), .ZN(n1098) );
INV_X1 U792 ( .A(KEYINPUT6), .ZN(n1099) );
NAND3_X1 U793 ( .A1(KEYINPUT12), .A2(n1097), .A3(n1100), .ZN(n1086) );
NOR3_X1 U794 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1078) );
NAND2_X1 U795 ( .A1(n1104), .A2(G478), .ZN(n1077) );
XOR2_X1 U796 ( .A(n1105), .B(KEYINPUT37), .Z(n1104) );
XOR2_X1 U797 ( .A(n1106), .B(n1107), .Z(n1076) );
XNOR2_X1 U798 ( .A(KEYINPUT63), .B(KEYINPUT58), .ZN(n1107) );
NAND2_X1 U799 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NAND2_X1 U800 ( .A1(G472), .A2(n1110), .ZN(n1109) );
XOR2_X1 U801 ( .A(KEYINPUT29), .B(n1111), .Z(n1108) );
NOR2_X1 U802 ( .A1(G472), .A2(n1110), .ZN(n1111) );
XOR2_X1 U803 ( .A(n1112), .B(n1113), .Z(G72) );
NOR2_X1 U804 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NAND2_X1 U806 ( .A1(n1118), .A2(n1119), .ZN(n1112) );
OR2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND3_X1 U808 ( .A1(n1122), .A2(n1120), .A3(n1121), .ZN(n1118) );
XNOR2_X1 U809 ( .A(n1123), .B(n1124), .ZN(n1121) );
XOR2_X1 U810 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U811 ( .A(n1127), .B(n1128), .ZN(n1126) );
XOR2_X1 U812 ( .A(n1129), .B(n1130), .Z(n1123) );
XOR2_X1 U813 ( .A(KEYINPUT34), .B(KEYINPUT10), .Z(n1130) );
NAND2_X1 U814 ( .A1(KEYINPUT55), .A2(n1131), .ZN(n1129) );
NAND2_X1 U815 ( .A1(n1115), .A2(n1132), .ZN(n1120) );
NAND2_X1 U816 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
INV_X1 U817 ( .A(n1135), .ZN(n1134) );
XOR2_X1 U818 ( .A(n1136), .B(KEYINPUT56), .Z(n1133) );
NAND2_X1 U819 ( .A1(G953), .A2(n1117), .ZN(n1122) );
NAND2_X1 U820 ( .A1(n1137), .A2(n1138), .ZN(G69) );
NAND2_X1 U821 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XOR2_X1 U822 ( .A(KEYINPUT11), .B(n1141), .Z(n1137) );
NOR2_X1 U823 ( .A1(n1139), .A2(n1140), .ZN(n1141) );
NAND2_X1 U824 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NAND2_X1 U825 ( .A1(G953), .A2(n1144), .ZN(n1143) );
AND2_X1 U826 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
NAND3_X1 U827 ( .A1(n1147), .A2(n1142), .A3(n1148), .ZN(n1146) );
XNOR2_X1 U828 ( .A(n1149), .B(n1150), .ZN(n1148) );
INV_X1 U829 ( .A(n1151), .ZN(n1142) );
NAND2_X1 U830 ( .A1(n1152), .A2(n1115), .ZN(n1147) );
XOR2_X1 U831 ( .A(n1153), .B(KEYINPUT28), .Z(n1145) );
NAND3_X1 U832 ( .A1(n1152), .A2(n1115), .A3(n1154), .ZN(n1153) );
XNOR2_X1 U833 ( .A(n1149), .B(n1155), .ZN(n1154) );
INV_X1 U834 ( .A(n1150), .ZN(n1155) );
NAND2_X1 U835 ( .A1(KEYINPUT0), .A2(n1156), .ZN(n1149) );
NOR2_X1 U836 ( .A1(n1157), .A2(n1158), .ZN(G66) );
NOR3_X1 U837 ( .A1(n1091), .A2(n1159), .A3(n1160), .ZN(n1158) );
NOR2_X1 U838 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1047), .A2(n1092), .ZN(n1161) );
NOR3_X1 U840 ( .A1(n1163), .A2(n1092), .A3(n1164), .ZN(n1159) );
INV_X1 U841 ( .A(n1162), .ZN(n1163) );
NOR2_X1 U842 ( .A1(n1157), .A2(n1165), .ZN(G63) );
XNOR2_X1 U843 ( .A(n1166), .B(n1167), .ZN(n1165) );
AND2_X1 U844 ( .A1(G478), .A2(n1168), .ZN(n1167) );
NOR2_X1 U845 ( .A1(n1157), .A2(n1169), .ZN(G60) );
XOR2_X1 U846 ( .A(n1170), .B(n1171), .Z(n1169) );
AND2_X1 U847 ( .A1(G475), .A2(n1168), .ZN(n1170) );
XOR2_X1 U848 ( .A(G104), .B(n1172), .Z(G6) );
NOR2_X1 U849 ( .A1(n1157), .A2(n1173), .ZN(G57) );
XOR2_X1 U850 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U851 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U852 ( .A1(KEYINPUT21), .A2(n1178), .ZN(n1176) );
XOR2_X1 U853 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U854 ( .A(n1181), .B(n1182), .Z(n1179) );
AND2_X1 U855 ( .A1(G472), .A2(n1168), .ZN(n1182) );
XNOR2_X1 U856 ( .A(n1183), .B(KEYINPUT59), .ZN(n1174) );
NOR2_X1 U857 ( .A1(n1157), .A2(n1184), .ZN(G54) );
XOR2_X1 U858 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U859 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U860 ( .A(KEYINPUT26), .B(n1189), .Z(n1188) );
NOR2_X1 U861 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U862 ( .A1(n1192), .A2(n1193), .ZN(n1187) );
XOR2_X1 U863 ( .A(KEYINPUT43), .B(n1190), .Z(n1193) );
XNOR2_X1 U864 ( .A(n1194), .B(n1195), .ZN(n1190) );
NAND2_X1 U865 ( .A1(KEYINPUT2), .A2(n1196), .ZN(n1194) );
INV_X1 U866 ( .A(n1191), .ZN(n1192) );
XOR2_X1 U867 ( .A(n1197), .B(n1198), .Z(n1191) );
NOR2_X1 U868 ( .A1(KEYINPUT44), .A2(n1199), .ZN(n1198) );
XOR2_X1 U869 ( .A(n1125), .B(n1200), .Z(n1199) );
NOR4_X1 U870 ( .A1(n1201), .A2(n1202), .A3(KEYINPUT25), .A4(n1203), .ZN(n1185) );
INV_X1 U871 ( .A(G469), .ZN(n1203) );
NOR2_X1 U872 ( .A1(n1204), .A2(n1205), .ZN(n1202) );
INV_X1 U873 ( .A(KEYINPUT1), .ZN(n1205) );
NOR2_X1 U874 ( .A1(G902), .A2(n1047), .ZN(n1204) );
NOR2_X1 U875 ( .A1(KEYINPUT1), .A2(n1168), .ZN(n1201) );
NOR2_X1 U876 ( .A1(n1115), .A2(G952), .ZN(n1157) );
NOR2_X1 U877 ( .A1(n1206), .A2(n1207), .ZN(G51) );
XOR2_X1 U878 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U879 ( .A(KEYINPUT40), .B(n1210), .Z(n1209) );
NOR2_X1 U880 ( .A1(KEYINPUT36), .A2(n1211), .ZN(n1210) );
XOR2_X1 U881 ( .A(n1212), .B(n1213), .Z(n1208) );
NOR2_X1 U882 ( .A1(n1097), .A2(n1164), .ZN(n1213) );
INV_X1 U883 ( .A(n1168), .ZN(n1164) );
NOR2_X1 U884 ( .A1(n1214), .A2(n1047), .ZN(n1168) );
NOR3_X1 U885 ( .A1(n1152), .A2(n1136), .A3(n1135), .ZN(n1047) );
NAND4_X1 U886 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1135) );
NAND4_X1 U887 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1136) );
NAND3_X1 U888 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1219) );
NAND4_X1 U889 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1152) );
NOR4_X1 U890 ( .A1(n1230), .A2(n1231), .A3(n1172), .A4(n1232), .ZN(n1229) );
INV_X1 U891 ( .A(n1233), .ZN(n1232) );
AND4_X1 U892 ( .A1(n1234), .A2(n1075), .A3(n1067), .A4(n1070), .ZN(n1172) );
NOR3_X1 U893 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1228) );
NOR2_X1 U894 ( .A1(n1041), .A2(n1238), .ZN(n1237) );
XOR2_X1 U895 ( .A(n1040), .B(KEYINPUT17), .Z(n1238) );
NAND4_X1 U896 ( .A1(n1067), .A2(n1074), .A3(n1070), .A4(n1239), .ZN(n1040) );
AND4_X1 U897 ( .A1(n1041), .A2(KEYINPUT60), .A3(n1239), .A4(n1240), .ZN(n1236) );
INV_X1 U898 ( .A(n1061), .ZN(n1041) );
NOR2_X1 U899 ( .A1(KEYINPUT60), .A2(n1241), .ZN(n1235) );
NAND2_X1 U900 ( .A1(n1242), .A2(n1243), .ZN(n1226) );
NOR2_X1 U901 ( .A1(G952), .A2(n1244), .ZN(n1206) );
XNOR2_X1 U902 ( .A(KEYINPUT47), .B(n1115), .ZN(n1244) );
XOR2_X1 U903 ( .A(n1220), .B(n1245), .Z(G48) );
XOR2_X1 U904 ( .A(KEYINPUT35), .B(G146), .Z(n1245) );
NAND3_X1 U905 ( .A1(n1075), .A2(n1061), .A3(n1224), .ZN(n1220) );
XNOR2_X1 U906 ( .A(G143), .B(n1221), .ZN(G45) );
NAND4_X1 U907 ( .A1(n1246), .A2(n1061), .A3(n1082), .A4(n1247), .ZN(n1221) );
XNOR2_X1 U908 ( .A(n1248), .B(n1222), .ZN(G42) );
NAND3_X1 U909 ( .A1(n1249), .A2(n1067), .A3(n1223), .ZN(n1222) );
NAND2_X1 U910 ( .A1(KEYINPUT27), .A2(n1250), .ZN(n1248) );
XNOR2_X1 U911 ( .A(n1131), .B(n1251), .ZN(G39) );
NOR4_X1 U912 ( .A1(KEYINPUT62), .A2(n1252), .A3(n1065), .A4(n1052), .ZN(n1251) );
INV_X1 U913 ( .A(n1225), .ZN(n1052) );
INV_X1 U914 ( .A(n1223), .ZN(n1065) );
XNOR2_X1 U915 ( .A(G134), .B(n1215), .ZN(G36) );
NAND3_X1 U916 ( .A1(n1223), .A2(n1074), .A3(n1246), .ZN(n1215) );
XNOR2_X1 U917 ( .A(G131), .B(n1216), .ZN(G33) );
NAND3_X1 U918 ( .A1(n1223), .A2(n1075), .A3(n1246), .ZN(n1216) );
AND2_X1 U919 ( .A1(n1243), .A2(n1253), .ZN(n1246) );
NOR2_X1 U920 ( .A1(n1062), .A2(n1103), .ZN(n1223) );
XNOR2_X1 U921 ( .A(G128), .B(n1217), .ZN(G30) );
NAND3_X1 U922 ( .A1(n1061), .A2(n1074), .A3(n1224), .ZN(n1217) );
INV_X1 U923 ( .A(n1252), .ZN(n1224) );
NAND3_X1 U924 ( .A1(n1067), .A2(n1253), .A3(n1072), .ZN(n1252) );
XNOR2_X1 U925 ( .A(G101), .B(n1254), .ZN(G3) );
NAND3_X1 U926 ( .A1(n1242), .A2(n1243), .A3(KEYINPUT57), .ZN(n1254) );
AND3_X1 U927 ( .A1(n1255), .A2(n1256), .A3(n1067), .ZN(n1243) );
XNOR2_X1 U928 ( .A(G125), .B(n1218), .ZN(G27) );
NAND3_X1 U929 ( .A1(n1249), .A2(n1061), .A3(n1257), .ZN(n1218) );
AND4_X1 U930 ( .A1(n1258), .A2(n1075), .A3(n1259), .A4(n1253), .ZN(n1249) );
NAND2_X1 U931 ( .A1(n1049), .A2(n1260), .ZN(n1253) );
NAND4_X1 U932 ( .A1(G902), .A2(G953), .A3(n1261), .A4(n1117), .ZN(n1260) );
INV_X1 U933 ( .A(G900), .ZN(n1117) );
XNOR2_X1 U934 ( .A(G122), .B(n1241), .ZN(G24) );
NAND2_X1 U935 ( .A1(n1240), .A2(n1234), .ZN(n1241) );
NOR4_X1 U936 ( .A1(n1059), .A2(n1055), .A3(n1262), .A4(n1263), .ZN(n1240) );
INV_X1 U937 ( .A(n1070), .ZN(n1055) );
NOR2_X1 U938 ( .A1(n1259), .A2(n1256), .ZN(n1070) );
INV_X1 U939 ( .A(n1257), .ZN(n1059) );
XNOR2_X1 U940 ( .A(G119), .B(n1227), .ZN(G21) );
NAND3_X1 U941 ( .A1(n1072), .A2(n1257), .A3(n1242), .ZN(n1227) );
NOR2_X1 U942 ( .A1(n1258), .A2(n1255), .ZN(n1072) );
XOR2_X1 U943 ( .A(G116), .B(n1231), .Z(G18) );
AND2_X1 U944 ( .A1(n1264), .A2(n1074), .ZN(n1231) );
NOR2_X1 U945 ( .A1(n1082), .A2(n1263), .ZN(n1074) );
XNOR2_X1 U946 ( .A(n1265), .B(n1230), .ZN(G15) );
AND2_X1 U947 ( .A1(n1264), .A2(n1075), .ZN(n1230) );
NOR2_X1 U948 ( .A1(n1247), .A2(n1262), .ZN(n1075) );
INV_X1 U949 ( .A(n1082), .ZN(n1262) );
AND4_X1 U950 ( .A1(n1234), .A2(n1257), .A3(n1255), .A4(n1256), .ZN(n1264) );
INV_X1 U951 ( .A(n1259), .ZN(n1255) );
NOR2_X1 U952 ( .A1(n1068), .A2(n1101), .ZN(n1257) );
INV_X1 U953 ( .A(n1069), .ZN(n1101) );
XNOR2_X1 U954 ( .A(G110), .B(n1233), .ZN(G12) );
NAND4_X1 U955 ( .A1(n1242), .A2(n1067), .A3(n1258), .A4(n1259), .ZN(n1233) );
XNOR2_X1 U956 ( .A(n1092), .B(n1266), .ZN(n1259) );
NOR2_X1 U957 ( .A1(KEYINPUT13), .A2(n1267), .ZN(n1266) );
INV_X1 U958 ( .A(n1091), .ZN(n1267) );
NOR2_X1 U959 ( .A1(n1162), .A2(G902), .ZN(n1091) );
XNOR2_X1 U960 ( .A(n1268), .B(n1269), .ZN(n1162) );
NOR2_X1 U961 ( .A1(KEYINPUT33), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U962 ( .A(G110), .B(n1271), .ZN(n1270) );
NAND2_X1 U963 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
OR2_X1 U964 ( .A1(n1274), .A2(G119), .ZN(n1273) );
XOR2_X1 U965 ( .A(n1275), .B(KEYINPUT42), .Z(n1272) );
NAND2_X1 U966 ( .A1(G119), .A2(n1274), .ZN(n1275) );
NAND2_X1 U967 ( .A1(n1276), .A2(n1277), .ZN(n1268) );
NAND2_X1 U968 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
INV_X1 U969 ( .A(KEYINPUT38), .ZN(n1279) );
XOR2_X1 U970 ( .A(n1280), .B(n1281), .Z(n1278) );
NAND2_X1 U971 ( .A1(G146), .A2(n1127), .ZN(n1280) );
NAND2_X1 U972 ( .A1(n1282), .A2(KEYINPUT38), .ZN(n1276) );
XNOR2_X1 U973 ( .A(n1281), .B(n1283), .ZN(n1282) );
XNOR2_X1 U974 ( .A(n1284), .B(n1131), .ZN(n1281) );
INV_X1 U975 ( .A(G137), .ZN(n1131) );
NAND3_X1 U976 ( .A1(n1285), .A2(G221), .A3(KEYINPUT14), .ZN(n1284) );
NAND2_X1 U977 ( .A1(G217), .A2(n1286), .ZN(n1092) );
INV_X1 U978 ( .A(n1256), .ZN(n1258) );
XNOR2_X1 U979 ( .A(n1110), .B(n1287), .ZN(n1256) );
XOR2_X1 U980 ( .A(KEYINPUT30), .B(G472), .Z(n1287) );
NAND2_X1 U981 ( .A1(n1288), .A2(n1214), .ZN(n1110) );
XOR2_X1 U982 ( .A(n1289), .B(n1290), .Z(n1288) );
XNOR2_X1 U983 ( .A(n1177), .B(n1291), .ZN(n1290) );
NAND2_X1 U984 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
OR2_X1 U985 ( .A1(n1180), .A2(KEYINPUT4), .ZN(n1293) );
XOR2_X1 U986 ( .A(n1197), .B(n1294), .Z(n1180) );
NAND3_X1 U987 ( .A1(n1294), .A2(n1295), .A3(KEYINPUT4), .ZN(n1292) );
XOR2_X1 U988 ( .A(n1296), .B(n1181), .Z(n1289) );
XOR2_X1 U989 ( .A(n1297), .B(n1298), .Z(n1181) );
NAND2_X1 U990 ( .A1(KEYINPUT50), .A2(G113), .ZN(n1297) );
NAND2_X1 U991 ( .A1(KEYINPUT8), .A2(n1183), .ZN(n1296) );
AND3_X1 U992 ( .A1(n1299), .A2(n1115), .A3(G210), .ZN(n1183) );
AND2_X1 U993 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U994 ( .A1(G221), .A2(n1286), .ZN(n1069) );
NAND2_X1 U995 ( .A1(G234), .A2(n1214), .ZN(n1286) );
XOR2_X1 U996 ( .A(n1083), .B(n1300), .Z(n1068) );
NOR2_X1 U997 ( .A1(G469), .A2(KEYINPUT15), .ZN(n1300) );
NAND2_X1 U998 ( .A1(n1301), .A2(n1214), .ZN(n1083) );
XOR2_X1 U999 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U1000 ( .A(n1295), .B(n1195), .ZN(n1303) );
XNOR2_X1 U1001 ( .A(n1250), .B(n1304), .ZN(n1195) );
NOR2_X1 U1002 ( .A1(G953), .A2(n1116), .ZN(n1304) );
INV_X1 U1003 ( .A(G227), .ZN(n1116) );
INV_X1 U1004 ( .A(G140), .ZN(n1250) );
INV_X1 U1005 ( .A(n1197), .ZN(n1295) );
XNOR2_X1 U1006 ( .A(n1305), .B(n1128), .ZN(n1197) );
XOR2_X1 U1007 ( .A(G131), .B(G134), .Z(n1128) );
XNOR2_X1 U1008 ( .A(G137), .B(KEYINPUT16), .ZN(n1305) );
XOR2_X1 U1009 ( .A(n1306), .B(n1307), .Z(n1302) );
XNOR2_X1 U1010 ( .A(KEYINPUT61), .B(n1196), .ZN(n1307) );
INV_X1 U1011 ( .A(G110), .ZN(n1196) );
NAND2_X1 U1012 ( .A1(KEYINPUT5), .A2(n1308), .ZN(n1306) );
XOR2_X1 U1013 ( .A(n1309), .B(n1125), .Z(n1308) );
XOR2_X1 U1014 ( .A(n1310), .B(n1311), .Z(n1125) );
NOR2_X1 U1015 ( .A1(KEYINPUT31), .A2(n1312), .ZN(n1311) );
XNOR2_X1 U1016 ( .A(G128), .B(KEYINPUT45), .ZN(n1312) );
XNOR2_X1 U1017 ( .A(G143), .B(G146), .ZN(n1310) );
NAND2_X1 U1018 ( .A1(KEYINPUT23), .A2(n1200), .ZN(n1309) );
XNOR2_X1 U1019 ( .A(n1313), .B(n1177), .ZN(n1200) );
XOR2_X1 U1020 ( .A(n1314), .B(G104), .Z(n1313) );
NAND2_X1 U1021 ( .A1(KEYINPUT22), .A2(n1038), .ZN(n1314) );
AND2_X1 U1022 ( .A1(n1225), .A2(n1234), .ZN(n1242) );
AND2_X1 U1023 ( .A1(n1061), .A2(n1239), .ZN(n1234) );
NAND2_X1 U1024 ( .A1(n1049), .A2(n1315), .ZN(n1239) );
NAND3_X1 U1025 ( .A1(n1151), .A2(n1261), .A3(G902), .ZN(n1315) );
NOR2_X1 U1026 ( .A1(G898), .A2(n1115), .ZN(n1151) );
NAND3_X1 U1027 ( .A1(n1261), .A2(n1115), .A3(G952), .ZN(n1049) );
NAND2_X1 U1028 ( .A1(G237), .A2(G234), .ZN(n1261) );
NOR2_X1 U1029 ( .A1(n1316), .A2(n1103), .ZN(n1061) );
INV_X1 U1030 ( .A(n1063), .ZN(n1103) );
NAND2_X1 U1031 ( .A1(G214), .A2(n1317), .ZN(n1063) );
INV_X1 U1032 ( .A(n1062), .ZN(n1316) );
XOR2_X1 U1033 ( .A(n1318), .B(n1097), .Z(n1062) );
NAND2_X1 U1034 ( .A1(G210), .A2(n1317), .ZN(n1097) );
NAND2_X1 U1035 ( .A1(n1299), .A2(n1214), .ZN(n1317) );
XNOR2_X1 U1036 ( .A(n1100), .B(KEYINPUT46), .ZN(n1318) );
INV_X1 U1037 ( .A(n1094), .ZN(n1100) );
NAND2_X1 U1038 ( .A1(n1319), .A2(n1214), .ZN(n1094) );
XOR2_X1 U1039 ( .A(n1212), .B(n1320), .Z(n1319) );
XNOR2_X1 U1040 ( .A(KEYINPUT19), .B(n1211), .ZN(n1320) );
INV_X1 U1041 ( .A(G125), .ZN(n1211) );
XOR2_X1 U1042 ( .A(n1321), .B(n1322), .Z(n1212) );
XOR2_X1 U1043 ( .A(n1323), .B(n1294), .Z(n1322) );
XNOR2_X1 U1044 ( .A(n1274), .B(n1324), .ZN(n1294) );
NOR2_X1 U1045 ( .A1(KEYINPUT51), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1046 ( .A(n1326), .B(G146), .Z(n1325) );
NAND2_X1 U1047 ( .A1(KEYINPUT32), .A2(G143), .ZN(n1326) );
NOR2_X1 U1048 ( .A1(G953), .A2(n1144), .ZN(n1323) );
INV_X1 U1049 ( .A(G224), .ZN(n1144) );
XNOR2_X1 U1050 ( .A(n1156), .B(n1150), .ZN(n1321) );
XNOR2_X1 U1051 ( .A(G110), .B(n1327), .ZN(n1150) );
INV_X1 U1052 ( .A(G122), .ZN(n1327) );
XNOR2_X1 U1053 ( .A(n1328), .B(n1329), .ZN(n1156) );
XNOR2_X1 U1054 ( .A(n1038), .B(n1330), .ZN(n1329) );
XNOR2_X1 U1055 ( .A(KEYINPUT41), .B(n1265), .ZN(n1330) );
XOR2_X1 U1056 ( .A(n1331), .B(n1298), .Z(n1328) );
XOR2_X1 U1057 ( .A(G116), .B(G119), .Z(n1298) );
XOR2_X1 U1058 ( .A(n1332), .B(G104), .Z(n1331) );
NAND2_X1 U1059 ( .A1(KEYINPUT3), .A2(n1177), .ZN(n1332) );
XOR2_X1 U1060 ( .A(G101), .B(KEYINPUT39), .Z(n1177) );
NOR2_X1 U1061 ( .A1(n1247), .A2(n1082), .ZN(n1225) );
XNOR2_X1 U1062 ( .A(n1333), .B(G475), .ZN(n1082) );
NAND2_X1 U1063 ( .A1(n1334), .A2(n1214), .ZN(n1333) );
XOR2_X1 U1064 ( .A(KEYINPUT9), .B(n1171), .Z(n1334) );
XNOR2_X1 U1065 ( .A(n1335), .B(n1336), .ZN(n1171) );
XOR2_X1 U1066 ( .A(G104), .B(n1337), .Z(n1336) );
XNOR2_X1 U1067 ( .A(n1338), .B(G131), .ZN(n1337) );
XOR2_X1 U1068 ( .A(n1339), .B(n1283), .Z(n1335) );
XOR2_X1 U1069 ( .A(G146), .B(n1127), .Z(n1283) );
XOR2_X1 U1070 ( .A(G140), .B(G125), .Z(n1127) );
XOR2_X1 U1071 ( .A(n1340), .B(n1341), .Z(n1339) );
AND3_X1 U1072 ( .A1(G214), .A2(n1115), .A3(n1299), .ZN(n1341) );
INV_X1 U1073 ( .A(G237), .ZN(n1299) );
NAND2_X1 U1074 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1075 ( .A1(G122), .A2(n1265), .ZN(n1343) );
XOR2_X1 U1076 ( .A(KEYINPUT53), .B(n1344), .Z(n1342) );
NOR2_X1 U1077 ( .A1(G122), .A2(n1265), .ZN(n1344) );
INV_X1 U1078 ( .A(G113), .ZN(n1265) );
INV_X1 U1079 ( .A(n1263), .ZN(n1247) );
NOR2_X1 U1080 ( .A1(n1345), .A2(n1102), .ZN(n1263) );
NOR2_X1 U1081 ( .A1(n1105), .A2(G478), .ZN(n1102) );
AND2_X1 U1082 ( .A1(n1346), .A2(n1105), .ZN(n1345) );
NAND2_X1 U1083 ( .A1(n1166), .A2(n1214), .ZN(n1105) );
INV_X1 U1084 ( .A(G902), .ZN(n1214) );
XNOR2_X1 U1085 ( .A(n1347), .B(n1348), .ZN(n1166) );
AND2_X1 U1086 ( .A1(n1285), .A2(G217), .ZN(n1348) );
AND2_X1 U1087 ( .A1(G234), .A2(n1115), .ZN(n1285) );
INV_X1 U1088 ( .A(G953), .ZN(n1115) );
NAND2_X1 U1089 ( .A1(n1349), .A2(KEYINPUT54), .ZN(n1347) );
XOR2_X1 U1090 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1091 ( .A(n1038), .B(n1352), .ZN(n1351) );
NOR2_X1 U1092 ( .A1(KEYINPUT20), .A2(n1353), .ZN(n1352) );
XOR2_X1 U1093 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1094 ( .A(G134), .B(n1274), .ZN(n1355) );
INV_X1 U1095 ( .A(G128), .ZN(n1274) );
NAND2_X1 U1096 ( .A1(KEYINPUT49), .A2(n1338), .ZN(n1354) );
INV_X1 U1097 ( .A(G143), .ZN(n1338) );
INV_X1 U1098 ( .A(G107), .ZN(n1038) );
XNOR2_X1 U1099 ( .A(G116), .B(G122), .ZN(n1350) );
XNOR2_X1 U1100 ( .A(G478), .B(KEYINPUT7), .ZN(n1346) );
endmodule


