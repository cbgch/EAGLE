//Key = 0001100001101110110000010001001100101100101101010011000010110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350;

XOR2_X1 U754 ( .A(G107), .B(n1037), .Z(G9) );
NOR2_X1 U755 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NOR2_X1 U757 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND4_X1 U758 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
INV_X1 U759 ( .A(KEYINPUT59), .ZN(n1049) );
INV_X1 U760 ( .A(n1050), .ZN(n1044) );
NOR2_X1 U761 ( .A1(n1051), .A2(n1050), .ZN(n1042) );
NOR2_X1 U762 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U763 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
INV_X1 U764 ( .A(n1048), .ZN(n1055) );
NOR2_X1 U765 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U766 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR3_X1 U767 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1058) );
NOR2_X1 U768 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U769 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR3_X1 U771 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1061) );
XNOR2_X1 U772 ( .A(KEYINPUT42), .B(n1072), .ZN(n1069) );
AND2_X1 U773 ( .A1(n1046), .A2(KEYINPUT59), .ZN(n1060) );
AND3_X1 U774 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1056) );
NOR3_X1 U775 ( .A1(n1064), .A2(n1076), .A3(n1072), .ZN(n1052) );
NOR2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
AND2_X1 U777 ( .A1(n1048), .A2(n1079), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1080), .A2(n1059), .ZN(n1077) );
INV_X1 U779 ( .A(n1047), .ZN(n1059) );
NOR2_X1 U780 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XNOR2_X1 U781 ( .A(n1083), .B(KEYINPUT34), .ZN(n1082) );
NAND3_X1 U782 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1040) );
NOR3_X1 U783 ( .A1(n1087), .A2(G953), .A3(G952), .ZN(n1038) );
INV_X1 U784 ( .A(n1084), .ZN(n1087) );
NAND4_X1 U785 ( .A1(n1088), .A2(n1074), .A3(n1089), .A4(n1090), .ZN(n1084) );
NOR4_X1 U786 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
XOR2_X1 U787 ( .A(n1095), .B(G478), .Z(n1089) );
INV_X1 U788 ( .A(n1072), .ZN(n1074) );
XOR2_X1 U789 ( .A(n1096), .B(n1097), .Z(G72) );
XOR2_X1 U790 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U791 ( .A1(G953), .A2(n1100), .ZN(n1099) );
NAND2_X1 U792 ( .A1(G900), .A2(G227), .ZN(n1100) );
NAND2_X1 U793 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U794 ( .A1(G953), .A2(n1103), .ZN(n1102) );
XOR2_X1 U795 ( .A(n1104), .B(n1105), .Z(n1101) );
NAND3_X1 U796 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1104) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U799 ( .A(n1113), .ZN(n1111) );
OR3_X1 U800 ( .A1(n1112), .A2(n1113), .A3(KEYINPUT25), .ZN(n1107) );
XNOR2_X1 U801 ( .A(n1109), .B(n1114), .ZN(n1112) );
XOR2_X1 U802 ( .A(KEYINPUT9), .B(KEYINPUT35), .Z(n1114) );
NAND2_X1 U803 ( .A1(n1113), .A2(KEYINPUT25), .ZN(n1106) );
XOR2_X1 U804 ( .A(G131), .B(n1115), .Z(n1113) );
NOR2_X1 U805 ( .A1(KEYINPUT39), .A2(n1116), .ZN(n1115) );
NOR2_X1 U806 ( .A1(n1086), .A2(G953), .ZN(n1096) );
NAND3_X1 U807 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(G69) );
NAND3_X1 U808 ( .A1(n1120), .A2(n1121), .A3(G953), .ZN(n1119) );
NAND3_X1 U809 ( .A1(G224), .A2(n1122), .A3(G898), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1123), .A2(n1122), .ZN(n1118) );
INV_X1 U811 ( .A(KEYINPUT6), .ZN(n1122) );
NAND2_X1 U812 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U813 ( .A1(n1126), .A2(n1085), .ZN(n1125) );
XNOR2_X1 U814 ( .A(n1127), .B(n1128), .ZN(n1126) );
NAND3_X1 U815 ( .A1(n1128), .A2(G224), .A3(G953), .ZN(n1124) );
NAND2_X1 U816 ( .A1(KEYINPUT6), .A2(n1129), .ZN(n1117) );
NAND2_X1 U817 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U818 ( .A1(n1127), .A2(n1121), .ZN(n1131) );
NAND3_X1 U819 ( .A1(n1041), .A2(n1085), .A3(n1128), .ZN(n1130) );
INV_X1 U820 ( .A(n1121), .ZN(n1128) );
NAND2_X1 U821 ( .A1(n1132), .A2(n1133), .ZN(n1121) );
NAND2_X1 U822 ( .A1(G953), .A2(n1134), .ZN(n1133) );
XNOR2_X1 U823 ( .A(n1135), .B(n1136), .ZN(n1132) );
NAND2_X1 U824 ( .A1(KEYINPUT4), .A2(n1137), .ZN(n1135) );
XOR2_X1 U825 ( .A(KEYINPUT43), .B(n1138), .Z(n1137) );
NOR2_X1 U826 ( .A1(n1139), .A2(n1140), .ZN(G66) );
XOR2_X1 U827 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U828 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NOR2_X1 U829 ( .A1(n1139), .A2(n1145), .ZN(G63) );
XOR2_X1 U830 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U831 ( .A1(KEYINPUT57), .A2(n1148), .ZN(n1147) );
INV_X1 U832 ( .A(n1149), .ZN(n1148) );
NAND2_X1 U833 ( .A1(n1143), .A2(n1150), .ZN(n1146) );
XOR2_X1 U834 ( .A(KEYINPUT28), .B(G478), .Z(n1150) );
NOR2_X1 U835 ( .A1(n1139), .A2(n1151), .ZN(G60) );
XOR2_X1 U836 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U837 ( .A1(n1143), .A2(n1154), .ZN(n1152) );
XOR2_X1 U838 ( .A(KEYINPUT0), .B(G475), .Z(n1154) );
XOR2_X1 U839 ( .A(G104), .B(n1155), .Z(G6) );
NOR2_X1 U840 ( .A1(n1139), .A2(n1156), .ZN(G57) );
NOR2_X1 U841 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U842 ( .A(KEYINPUT61), .B(n1159), .Z(n1158) );
NOR2_X1 U843 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
AND2_X1 U844 ( .A1(n1161), .A2(n1160), .ZN(n1157) );
AND3_X1 U845 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1160) );
NAND2_X1 U846 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
OR4_X1 U847 ( .A1(n1165), .A2(KEYINPUT1), .A3(n1166), .A4(n1167), .ZN(n1163) );
INV_X1 U848 ( .A(KEYINPUT51), .ZN(n1166) );
NAND2_X1 U849 ( .A1(n1143), .A2(G472), .ZN(n1165) );
NAND2_X1 U850 ( .A1(n1167), .A2(n1168), .ZN(n1162) );
NAND3_X1 U851 ( .A1(G472), .A2(n1169), .A3(n1143), .ZN(n1168) );
INV_X1 U852 ( .A(KEYINPUT1), .ZN(n1169) );
XOR2_X1 U853 ( .A(n1170), .B(n1171), .Z(n1167) );
NOR2_X1 U854 ( .A1(KEYINPUT32), .A2(n1172), .ZN(n1171) );
NOR2_X1 U855 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U856 ( .A1(n1139), .A2(n1175), .ZN(G54) );
XOR2_X1 U857 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U858 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U859 ( .A(n1180), .B(n1181), .ZN(n1179) );
XOR2_X1 U860 ( .A(n1182), .B(n1183), .Z(n1176) );
XNOR2_X1 U861 ( .A(KEYINPUT62), .B(n1184), .ZN(n1183) );
NOR2_X1 U862 ( .A1(KEYINPUT21), .A2(n1185), .ZN(n1184) );
XOR2_X1 U863 ( .A(n1186), .B(n1187), .Z(n1185) );
XNOR2_X1 U864 ( .A(n1188), .B(n1189), .ZN(n1187) );
NOR2_X1 U865 ( .A1(G110), .A2(KEYINPUT52), .ZN(n1188) );
XOR2_X1 U866 ( .A(KEYINPUT44), .B(n1190), .Z(n1186) );
NAND2_X1 U867 ( .A1(n1143), .A2(G469), .ZN(n1182) );
NOR2_X1 U868 ( .A1(n1139), .A2(n1191), .ZN(G51) );
XOR2_X1 U869 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U870 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U871 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NOR3_X1 U872 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1197) );
INV_X1 U873 ( .A(KEYINPUT38), .ZN(n1198) );
NOR2_X1 U874 ( .A1(KEYINPUT38), .A2(n1201), .ZN(n1196) );
XNOR2_X1 U875 ( .A(n1202), .B(n1203), .ZN(n1192) );
NAND2_X1 U876 ( .A1(n1143), .A2(n1204), .ZN(n1202) );
AND2_X1 U877 ( .A1(G902), .A2(n1205), .ZN(n1143) );
NAND2_X1 U878 ( .A1(n1127), .A2(n1206), .ZN(n1205) );
XOR2_X1 U879 ( .A(KEYINPUT48), .B(n1086), .Z(n1206) );
AND4_X1 U880 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1086) );
AND4_X1 U881 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
NOR2_X1 U882 ( .A1(n1215), .A2(n1216), .ZN(n1209) );
INV_X1 U883 ( .A(n1041), .ZN(n1127) );
NAND4_X1 U884 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1041) );
NOR4_X1 U885 ( .A1(n1037), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1220) );
AND3_X1 U886 ( .A1(n1079), .A2(n1048), .A3(n1224), .ZN(n1037) );
NOR2_X1 U887 ( .A1(n1155), .A2(n1225), .ZN(n1219) );
NOR2_X1 U888 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U889 ( .A(n1228), .B(KEYINPUT18), .Z(n1226) );
AND3_X1 U890 ( .A1(n1224), .A2(n1048), .A3(n1075), .ZN(n1155) );
NOR2_X1 U891 ( .A1(n1085), .A2(G952), .ZN(n1139) );
XOR2_X1 U892 ( .A(G146), .B(n1229), .Z(G48) );
NOR2_X1 U893 ( .A1(KEYINPUT8), .A2(n1214), .ZN(n1229) );
NAND3_X1 U894 ( .A1(n1230), .A2(n1075), .A3(n1231), .ZN(n1214) );
XNOR2_X1 U895 ( .A(G143), .B(n1213), .ZN(G45) );
NAND3_X1 U896 ( .A1(n1232), .A2(n1081), .A3(n1231), .ZN(n1213) );
XNOR2_X1 U897 ( .A(G140), .B(n1212), .ZN(G42) );
NAND3_X1 U898 ( .A1(n1075), .A2(n1083), .A3(n1233), .ZN(n1212) );
XNOR2_X1 U899 ( .A(G137), .B(n1211), .ZN(G39) );
NAND3_X1 U900 ( .A1(n1230), .A2(n1047), .A3(n1233), .ZN(n1211) );
XOR2_X1 U901 ( .A(G134), .B(n1216), .Z(G36) );
AND3_X1 U902 ( .A1(n1081), .A2(n1079), .A3(n1233), .ZN(n1216) );
NAND2_X1 U903 ( .A1(n1234), .A2(n1235), .ZN(G33) );
NAND2_X1 U904 ( .A1(n1215), .A2(n1236), .ZN(n1235) );
XOR2_X1 U905 ( .A(KEYINPUT14), .B(n1237), .Z(n1234) );
NOR2_X1 U906 ( .A1(n1215), .A2(n1236), .ZN(n1237) );
INV_X1 U907 ( .A(G131), .ZN(n1236) );
AND3_X1 U908 ( .A1(n1081), .A2(n1075), .A3(n1233), .ZN(n1215) );
AND2_X1 U909 ( .A1(n1046), .A2(n1238), .ZN(n1233) );
NOR3_X1 U910 ( .A1(n1088), .A2(n1091), .A3(n1072), .ZN(n1046) );
NAND2_X1 U911 ( .A1(n1239), .A2(n1068), .ZN(n1072) );
INV_X1 U912 ( .A(n1067), .ZN(n1239) );
XNOR2_X1 U913 ( .A(G128), .B(n1207), .ZN(G30) );
NAND3_X1 U914 ( .A1(n1230), .A2(n1079), .A3(n1231), .ZN(n1207) );
AND3_X1 U915 ( .A1(n1071), .A2(n1070), .A3(n1240), .ZN(n1231) );
NAND2_X1 U916 ( .A1(n1241), .A2(n1242), .ZN(G3) );
OR2_X1 U917 ( .A1(n1243), .A2(G101), .ZN(n1242) );
NAND2_X1 U918 ( .A1(G101), .A2(n1244), .ZN(n1241) );
NAND2_X1 U919 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
OR2_X1 U920 ( .A1(n1217), .A2(KEYINPUT17), .ZN(n1246) );
NAND2_X1 U921 ( .A1(KEYINPUT17), .A2(n1243), .ZN(n1245) );
NAND2_X1 U922 ( .A1(KEYINPUT63), .A2(n1247), .ZN(n1243) );
INV_X1 U923 ( .A(n1217), .ZN(n1247) );
NAND3_X1 U924 ( .A1(n1224), .A2(n1047), .A3(n1081), .ZN(n1217) );
XNOR2_X1 U925 ( .A(G125), .B(n1208), .ZN(G27) );
NAND4_X1 U926 ( .A1(n1240), .A2(n1073), .A3(n1075), .A4(n1083), .ZN(n1208) );
AND2_X1 U927 ( .A1(n1066), .A2(n1238), .ZN(n1240) );
NAND2_X1 U928 ( .A1(n1050), .A2(n1248), .ZN(n1238) );
NAND4_X1 U929 ( .A1(G953), .A2(G902), .A3(n1103), .A4(n1249), .ZN(n1248) );
XOR2_X1 U930 ( .A(KEYINPUT3), .B(G900), .Z(n1103) );
XOR2_X1 U931 ( .A(G122), .B(n1250), .Z(G24) );
NOR2_X1 U932 ( .A1(n1227), .A2(n1228), .ZN(n1250) );
NAND4_X1 U933 ( .A1(n1232), .A2(n1073), .A3(n1048), .A4(n1251), .ZN(n1228) );
NAND2_X1 U934 ( .A1(n1252), .A2(n1253), .ZN(n1048) );
NAND2_X1 U935 ( .A1(n1083), .A2(n1254), .ZN(n1253) );
OR3_X1 U936 ( .A1(n1094), .A2(n1093), .A3(n1254), .ZN(n1252) );
AND2_X1 U937 ( .A1(n1255), .A2(n1092), .ZN(n1232) );
XNOR2_X1 U938 ( .A(KEYINPUT46), .B(n1256), .ZN(n1255) );
XNOR2_X1 U939 ( .A(G119), .B(n1218), .ZN(G21) );
NAND3_X1 U940 ( .A1(n1257), .A2(n1047), .A3(n1230), .ZN(n1218) );
AND2_X1 U941 ( .A1(n1093), .A2(n1094), .ZN(n1230) );
XOR2_X1 U942 ( .A(G116), .B(n1223), .Z(G18) );
AND3_X1 U943 ( .A1(n1257), .A2(n1079), .A3(n1081), .ZN(n1223) );
NOR2_X1 U944 ( .A1(n1092), .A2(n1256), .ZN(n1079) );
XOR2_X1 U945 ( .A(G113), .B(n1222), .Z(G15) );
AND3_X1 U946 ( .A1(n1257), .A2(n1075), .A3(n1081), .ZN(n1222) );
AND2_X1 U947 ( .A1(n1258), .A2(n1094), .ZN(n1081) );
XNOR2_X1 U948 ( .A(n1254), .B(n1093), .ZN(n1258) );
INV_X1 U949 ( .A(KEYINPUT12), .ZN(n1254) );
AND3_X1 U950 ( .A1(n1066), .A2(n1251), .A3(n1073), .ZN(n1257) );
INV_X1 U951 ( .A(n1064), .ZN(n1073) );
NAND2_X1 U952 ( .A1(n1259), .A2(n1088), .ZN(n1064) );
INV_X1 U953 ( .A(n1071), .ZN(n1088) );
XNOR2_X1 U954 ( .A(n1091), .B(KEYINPUT5), .ZN(n1259) );
INV_X1 U955 ( .A(n1070), .ZN(n1091) );
XOR2_X1 U956 ( .A(G110), .B(n1221), .Z(G12) );
AND3_X1 U957 ( .A1(n1083), .A2(n1047), .A3(n1224), .ZN(n1221) );
AND4_X1 U958 ( .A1(n1066), .A2(n1071), .A3(n1251), .A4(n1070), .ZN(n1224) );
NAND2_X1 U959 ( .A1(G221), .A2(n1260), .ZN(n1070) );
NAND2_X1 U960 ( .A1(n1050), .A2(n1261), .ZN(n1251) );
NAND4_X1 U961 ( .A1(G953), .A2(G902), .A3(n1249), .A4(n1134), .ZN(n1261) );
INV_X1 U962 ( .A(G898), .ZN(n1134) );
NAND3_X1 U963 ( .A1(n1249), .A2(n1085), .A3(G952), .ZN(n1050) );
NAND2_X1 U964 ( .A1(G237), .A2(G234), .ZN(n1249) );
XNOR2_X1 U965 ( .A(n1262), .B(G469), .ZN(n1071) );
NAND2_X1 U966 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U967 ( .A(n1265), .B(n1190), .Z(n1263) );
AND2_X1 U968 ( .A1(G227), .A2(n1085), .ZN(n1190) );
XOR2_X1 U969 ( .A(n1266), .B(n1267), .Z(n1265) );
NOR2_X1 U970 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XOR2_X1 U971 ( .A(KEYINPUT49), .B(n1270), .Z(n1269) );
NOR2_X1 U972 ( .A1(G110), .A2(n1189), .ZN(n1270) );
AND2_X1 U973 ( .A1(G110), .A2(n1189), .ZN(n1268) );
XNOR2_X1 U974 ( .A(G140), .B(KEYINPUT55), .ZN(n1189) );
NAND3_X1 U975 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1266) );
NAND2_X1 U976 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
NAND2_X1 U977 ( .A1(n1276), .A2(KEYINPUT56), .ZN(n1275) );
XNOR2_X1 U978 ( .A(n1180), .B(KEYINPUT58), .ZN(n1276) );
INV_X1 U979 ( .A(n1277), .ZN(n1274) );
NAND3_X1 U980 ( .A1(KEYINPUT56), .A2(n1277), .A3(n1180), .ZN(n1272) );
XOR2_X1 U981 ( .A(n1278), .B(n1181), .Z(n1277) );
INV_X1 U982 ( .A(n1109), .ZN(n1181) );
XOR2_X1 U983 ( .A(n1279), .B(n1280), .Z(n1109) );
NOR2_X1 U984 ( .A1(KEYINPUT2), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U985 ( .A(G143), .B(KEYINPUT37), .ZN(n1281) );
XNOR2_X1 U986 ( .A(KEYINPUT19), .B(n1282), .ZN(n1278) );
NOR2_X1 U987 ( .A1(KEYINPUT11), .A2(n1178), .ZN(n1282) );
XOR2_X1 U988 ( .A(G101), .B(n1283), .Z(n1178) );
OR2_X1 U989 ( .A1(n1180), .A2(KEYINPUT56), .ZN(n1271) );
INV_X1 U990 ( .A(n1227), .ZN(n1066) );
NAND2_X1 U991 ( .A1(n1067), .A2(n1068), .ZN(n1227) );
NAND2_X1 U992 ( .A1(G214), .A2(n1284), .ZN(n1068) );
XNOR2_X1 U993 ( .A(n1285), .B(n1204), .ZN(n1067) );
AND2_X1 U994 ( .A1(G210), .A2(n1284), .ZN(n1204) );
NAND2_X1 U995 ( .A1(n1264), .A2(n1286), .ZN(n1284) );
NAND3_X1 U996 ( .A1(n1287), .A2(n1264), .A3(n1288), .ZN(n1285) );
XOR2_X1 U997 ( .A(KEYINPUT30), .B(n1289), .Z(n1288) );
NOR2_X1 U998 ( .A1(n1290), .A2(n1194), .ZN(n1289) );
NAND2_X1 U999 ( .A1(n1290), .A2(n1194), .ZN(n1287) );
XOR2_X1 U1000 ( .A(n1138), .B(n1136), .Z(n1194) );
XNOR2_X1 U1001 ( .A(n1291), .B(n1292), .ZN(n1136) );
XOR2_X1 U1002 ( .A(n1293), .B(n1283), .Z(n1292) );
XOR2_X1 U1003 ( .A(G104), .B(G107), .Z(n1283) );
NOR2_X1 U1004 ( .A1(G101), .A2(KEYINPUT7), .ZN(n1293) );
XNOR2_X1 U1005 ( .A(G110), .B(n1294), .ZN(n1291) );
NOR2_X1 U1006 ( .A1(KEYINPUT41), .A2(n1295), .ZN(n1294) );
XOR2_X1 U1007 ( .A(G119), .B(n1296), .Z(n1138) );
XNOR2_X1 U1008 ( .A(n1297), .B(n1201), .ZN(n1290) );
XNOR2_X1 U1009 ( .A(n1200), .B(n1199), .ZN(n1201) );
INV_X1 U1010 ( .A(G125), .ZN(n1200) );
XOR2_X1 U1011 ( .A(n1203), .B(KEYINPUT24), .Z(n1297) );
NAND2_X1 U1012 ( .A1(G224), .A2(n1085), .ZN(n1203) );
NAND2_X1 U1013 ( .A1(n1298), .A2(n1299), .ZN(n1047) );
OR3_X1 U1014 ( .A1(n1300), .A2(n1092), .A3(KEYINPUT33), .ZN(n1299) );
NAND2_X1 U1015 ( .A1(KEYINPUT33), .A2(n1075), .ZN(n1298) );
NOR2_X1 U1016 ( .A1(n1300), .A2(n1301), .ZN(n1075) );
INV_X1 U1017 ( .A(n1092), .ZN(n1301) );
XNOR2_X1 U1018 ( .A(n1302), .B(G475), .ZN(n1092) );
NAND2_X1 U1019 ( .A1(n1153), .A2(n1264), .ZN(n1302) );
XOR2_X1 U1020 ( .A(n1303), .B(n1304), .Z(n1153) );
XOR2_X1 U1021 ( .A(n1295), .B(n1305), .Z(n1304) );
XNOR2_X1 U1022 ( .A(n1306), .B(n1307), .ZN(n1305) );
NAND2_X1 U1023 ( .A1(KEYINPUT31), .A2(n1308), .ZN(n1307) );
NAND2_X1 U1024 ( .A1(KEYINPUT16), .A2(n1309), .ZN(n1306) );
XNOR2_X1 U1025 ( .A(G131), .B(n1310), .ZN(n1309) );
NAND2_X1 U1026 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND4_X1 U1027 ( .A1(G143), .A2(G214), .A3(n1286), .A4(n1085), .ZN(n1312) );
XOR2_X1 U1028 ( .A(n1313), .B(KEYINPUT26), .Z(n1311) );
NAND2_X1 U1029 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND3_X1 U1030 ( .A1(n1286), .A2(n1085), .A3(G214), .ZN(n1315) );
XNOR2_X1 U1031 ( .A(G104), .B(n1316), .ZN(n1303) );
XOR2_X1 U1032 ( .A(G146), .B(G113), .Z(n1316) );
XNOR2_X1 U1033 ( .A(n1256), .B(KEYINPUT15), .ZN(n1300) );
XNOR2_X1 U1034 ( .A(n1317), .B(n1095), .ZN(n1256) );
NAND2_X1 U1035 ( .A1(n1318), .A2(n1149), .ZN(n1095) );
XNOR2_X1 U1036 ( .A(n1319), .B(n1320), .ZN(n1149) );
XOR2_X1 U1037 ( .A(n1295), .B(n1321), .Z(n1320) );
XOR2_X1 U1038 ( .A(n1322), .B(n1323), .Z(n1321) );
NAND2_X1 U1039 ( .A1(KEYINPUT10), .A2(n1324), .ZN(n1322) );
XNOR2_X1 U1040 ( .A(G122), .B(KEYINPUT50), .ZN(n1295) );
XOR2_X1 U1041 ( .A(n1325), .B(n1326), .Z(n1319) );
XNOR2_X1 U1042 ( .A(n1314), .B(G116), .ZN(n1326) );
XOR2_X1 U1043 ( .A(n1327), .B(G107), .Z(n1325) );
NAND3_X1 U1044 ( .A1(G217), .A2(n1328), .A3(KEYINPUT36), .ZN(n1327) );
XNOR2_X1 U1045 ( .A(G902), .B(KEYINPUT54), .ZN(n1318) );
NAND2_X1 U1046 ( .A1(KEYINPUT47), .A2(G478), .ZN(n1317) );
NOR2_X1 U1047 ( .A1(n1094), .A2(n1329), .ZN(n1083) );
INV_X1 U1048 ( .A(n1093), .ZN(n1329) );
XNOR2_X1 U1049 ( .A(n1330), .B(n1144), .ZN(n1093) );
AND2_X1 U1050 ( .A1(G217), .A2(n1260), .ZN(n1144) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1264), .ZN(n1260) );
NAND2_X1 U1052 ( .A1(n1331), .A2(n1142), .ZN(n1330) );
XNOR2_X1 U1053 ( .A(n1332), .B(n1333), .ZN(n1142) );
XOR2_X1 U1054 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1055 ( .A(G137), .B(G110), .Z(n1335) );
XOR2_X1 U1056 ( .A(KEYINPUT27), .B(G146), .Z(n1334) );
XOR2_X1 U1057 ( .A(n1336), .B(n1337), .Z(n1332) );
AND2_X1 U1058 ( .A1(G221), .A2(n1328), .ZN(n1337) );
AND2_X1 U1059 ( .A1(G234), .A2(n1085), .ZN(n1328) );
XOR2_X1 U1060 ( .A(n1338), .B(n1339), .Z(n1336) );
NOR2_X1 U1061 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
XOR2_X1 U1062 ( .A(KEYINPUT60), .B(n1342), .Z(n1341) );
NOR2_X1 U1063 ( .A1(G119), .A2(n1324), .ZN(n1342) );
AND2_X1 U1064 ( .A1(n1324), .A2(G119), .ZN(n1340) );
INV_X1 U1065 ( .A(G128), .ZN(n1324) );
NAND2_X1 U1066 ( .A1(KEYINPUT40), .A2(n1308), .ZN(n1338) );
XOR2_X1 U1067 ( .A(n1105), .B(KEYINPUT13), .Z(n1308) );
XNOR2_X1 U1068 ( .A(G140), .B(G125), .ZN(n1105) );
XNOR2_X1 U1069 ( .A(KEYINPUT23), .B(n1264), .ZN(n1331) );
XNOR2_X1 U1070 ( .A(n1343), .B(G472), .ZN(n1094) );
NAND2_X1 U1071 ( .A1(n1344), .A2(n1264), .ZN(n1343) );
INV_X1 U1072 ( .A(G902), .ZN(n1264) );
XOR2_X1 U1073 ( .A(n1345), .B(n1346), .Z(n1344) );
XNOR2_X1 U1074 ( .A(n1161), .B(n1170), .ZN(n1346) );
XOR2_X1 U1075 ( .A(n1296), .B(n1347), .Z(n1170) );
NOR2_X1 U1076 ( .A1(G119), .A2(KEYINPUT22), .ZN(n1347) );
XOR2_X1 U1077 ( .A(G113), .B(G116), .Z(n1296) );
XOR2_X1 U1078 ( .A(G101), .B(n1348), .Z(n1161) );
AND3_X1 U1079 ( .A1(G210), .A2(n1085), .A3(n1286), .ZN(n1348) );
INV_X1 U1080 ( .A(G237), .ZN(n1286) );
INV_X1 U1081 ( .A(G953), .ZN(n1085) );
XNOR2_X1 U1082 ( .A(KEYINPUT45), .B(n1349), .ZN(n1345) );
NOR3_X1 U1083 ( .A1(n1350), .A2(KEYINPUT53), .A3(n1174), .ZN(n1349) );
AND2_X1 U1084 ( .A1(n1199), .A2(n1180), .ZN(n1174) );
XOR2_X1 U1085 ( .A(KEYINPUT29), .B(n1173), .Z(n1350) );
NOR2_X1 U1086 ( .A1(n1199), .A2(n1180), .ZN(n1173) );
XNOR2_X1 U1087 ( .A(G131), .B(n1116), .ZN(n1180) );
XNOR2_X1 U1088 ( .A(G137), .B(n1323), .ZN(n1116) );
XOR2_X1 U1089 ( .A(G134), .B(KEYINPUT20), .Z(n1323) );
XNOR2_X1 U1090 ( .A(n1314), .B(n1279), .ZN(n1199) );
XOR2_X1 U1091 ( .A(G128), .B(G146), .Z(n1279) );
INV_X1 U1092 ( .A(G143), .ZN(n1314) );
endmodule


