//Key = 1110110011001010011011001001100000000110010110100000111000101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286;

XNOR2_X1 U709 ( .A(G107), .B(n981), .ZN(G9) );
NOR2_X1 U710 ( .A1(n982), .A2(n983), .ZN(G75) );
NOR4_X1 U711 ( .A1(n984), .A2(n985), .A3(n986), .A4(n987), .ZN(n983) );
XOR2_X1 U712 ( .A(n988), .B(KEYINPUT42), .Z(n987) );
NAND2_X1 U713 ( .A1(n989), .A2(n990), .ZN(n988) );
NOR2_X1 U714 ( .A1(n991), .A2(n992), .ZN(n986) );
INV_X1 U715 ( .A(n993), .ZN(n992) );
NOR2_X1 U716 ( .A1(n994), .A2(n995), .ZN(n991) );
NOR3_X1 U717 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n995) );
NOR3_X1 U718 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n998) );
NOR2_X1 U719 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U720 ( .A1(n1004), .A2(n1005), .ZN(n997) );
NOR2_X1 U721 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NOR2_X1 U722 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR3_X1 U723 ( .A1(n1007), .A2(n1010), .A3(n999), .ZN(n994) );
NOR2_X1 U724 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U725 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR2_X1 U726 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U727 ( .A1(n1017), .A2(n1018), .ZN(n1011) );
NOR2_X1 U728 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
AND3_X1 U729 ( .A1(n1021), .A2(n1022), .A3(G221), .ZN(n1019) );
INV_X1 U730 ( .A(n1023), .ZN(n1007) );
NAND4_X1 U731 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n984) );
AND3_X1 U732 ( .A1(n1025), .A2(n1027), .A3(n1028), .ZN(n982) );
NAND4_X1 U733 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1025) );
NOR4_X1 U734 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
XOR2_X1 U735 ( .A(n1037), .B(KEYINPUT46), .Z(n1035) );
NOR3_X1 U736 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1034) );
NOR2_X1 U737 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR3_X1 U738 ( .A1(G478), .A2(KEYINPUT49), .A3(n1043), .ZN(n1039) );
INV_X1 U739 ( .A(n1041), .ZN(n1043) );
NOR2_X1 U740 ( .A1(n1044), .A2(KEYINPUT35), .ZN(n1041) );
AND2_X1 U741 ( .A1(n1044), .A2(KEYINPUT49), .ZN(n1038) );
XOR2_X1 U742 ( .A(n1045), .B(n1046), .Z(n1031) );
XNOR2_X1 U743 ( .A(n1047), .B(G475), .ZN(n1029) );
XOR2_X1 U744 ( .A(n1048), .B(n1049), .Z(G72) );
NOR2_X1 U745 ( .A1(n1050), .A2(n1027), .ZN(n1049) );
NOR2_X1 U746 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U747 ( .A1(KEYINPUT31), .A2(n1053), .ZN(n1048) );
XOR2_X1 U748 ( .A(n1054), .B(n1055), .Z(n1053) );
NOR2_X1 U749 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XOR2_X1 U750 ( .A(n1058), .B(KEYINPUT4), .Z(n1057) );
NAND2_X1 U751 ( .A1(n1059), .A2(n1052), .ZN(n1058) );
XOR2_X1 U752 ( .A(n1027), .B(KEYINPUT63), .Z(n1059) );
XOR2_X1 U753 ( .A(n1060), .B(n1061), .Z(n1056) );
XNOR2_X1 U754 ( .A(n1062), .B(n1063), .ZN(n1061) );
NOR3_X1 U755 ( .A1(KEYINPUT33), .A2(n1064), .A3(n1065), .ZN(n1062) );
AND2_X1 U756 ( .A1(KEYINPUT52), .A2(n1066), .ZN(n1065) );
NOR3_X1 U757 ( .A1(KEYINPUT52), .A2(G131), .A3(n1067), .ZN(n1064) );
NAND2_X1 U758 ( .A1(n1068), .A2(n1027), .ZN(n1054) );
NAND3_X1 U759 ( .A1(n1069), .A2(n1024), .A3(n1070), .ZN(n1068) );
XNOR2_X1 U760 ( .A(KEYINPUT27), .B(n1026), .ZN(n1069) );
XOR2_X1 U761 ( .A(n1071), .B(n1072), .Z(G69) );
NOR2_X1 U762 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND3_X1 U763 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1071) );
INV_X1 U764 ( .A(n1073), .ZN(n1077) );
NAND2_X1 U765 ( .A1(G953), .A2(n1078), .ZN(n1076) );
NAND2_X1 U766 ( .A1(n1079), .A2(n1027), .ZN(n1075) );
NAND2_X1 U767 ( .A1(n1080), .A2(n989), .ZN(n1079) );
XOR2_X1 U768 ( .A(n990), .B(KEYINPUT59), .Z(n1080) );
NOR2_X1 U769 ( .A1(n1081), .A2(n1082), .ZN(G66) );
XNOR2_X1 U770 ( .A(n1083), .B(n1084), .ZN(n1082) );
NAND3_X1 U771 ( .A1(n1085), .A2(G217), .A3(KEYINPUT44), .ZN(n1084) );
NAND2_X1 U772 ( .A1(KEYINPUT0), .A2(n1086), .ZN(n1083) );
NOR2_X1 U773 ( .A1(n1081), .A2(n1087), .ZN(G63) );
XOR2_X1 U774 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U775 ( .A1(KEYINPUT47), .A2(n1090), .ZN(n1089) );
NAND3_X1 U776 ( .A1(n1091), .A2(n1092), .A3(G478), .ZN(n1088) );
XOR2_X1 U777 ( .A(KEYINPUT13), .B(G902), .Z(n1091) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1093), .ZN(G60) );
NOR3_X1 U779 ( .A1(n1047), .A2(n1094), .A3(n1095), .ZN(n1093) );
NOR3_X1 U780 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
INV_X1 U781 ( .A(n1099), .ZN(n1096) );
NOR2_X1 U782 ( .A1(n1100), .A2(n1099), .ZN(n1094) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1097), .ZN(n1100) );
XNOR2_X1 U784 ( .A(G475), .B(KEYINPUT25), .ZN(n1097) );
INV_X1 U785 ( .A(n1092), .ZN(n1101) );
XOR2_X1 U786 ( .A(n1102), .B(n1103), .Z(G6) );
NAND2_X1 U787 ( .A1(KEYINPUT37), .A2(G104), .ZN(n1103) );
NOR2_X1 U788 ( .A1(n1081), .A2(n1104), .ZN(G57) );
NOR2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U790 ( .A(n1107), .B(KEYINPUT17), .Z(n1106) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
XNOR2_X1 U793 ( .A(n1110), .B(n1111), .ZN(n1109) );
NOR2_X1 U794 ( .A1(G101), .A2(KEYINPUT39), .ZN(n1111) );
AND2_X1 U795 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
NAND3_X1 U796 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(n1112) );
NAND2_X1 U798 ( .A1(n1116), .A2(n1115), .ZN(n1118) );
NAND2_X1 U799 ( .A1(n1119), .A2(n1120), .ZN(n1115) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U801 ( .A(n1123), .B(n1124), .Z(n1119) );
XOR2_X1 U802 ( .A(n1125), .B(KEYINPUT61), .Z(n1116) );
NAND2_X1 U803 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U804 ( .A(n1066), .B(n1122), .Z(n1127) );
XNOR2_X1 U805 ( .A(n1128), .B(KEYINPUT24), .ZN(n1122) );
NAND2_X1 U806 ( .A1(KEYINPUT60), .A2(n1129), .ZN(n1128) );
XNOR2_X1 U807 ( .A(n1123), .B(n1124), .ZN(n1126) );
XOR2_X1 U808 ( .A(KEYINPUT12), .B(n1114), .Z(n1117) );
AND2_X1 U809 ( .A1(n1085), .A2(G472), .ZN(n1114) );
NOR2_X1 U810 ( .A1(n1081), .A2(n1130), .ZN(G54) );
XOR2_X1 U811 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U812 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U813 ( .A(n1063), .B(n1135), .ZN(n1134) );
XOR2_X1 U814 ( .A(n1136), .B(n1137), .Z(n1131) );
XNOR2_X1 U815 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR3_X1 U816 ( .A1(n1051), .A2(KEYINPUT56), .A3(G953), .ZN(n1139) );
INV_X1 U817 ( .A(G227), .ZN(n1051) );
NAND3_X1 U818 ( .A1(n1085), .A2(G469), .A3(KEYINPUT1), .ZN(n1138) );
XNOR2_X1 U819 ( .A(KEYINPUT28), .B(KEYINPUT14), .ZN(n1136) );
NOR2_X1 U820 ( .A1(n1081), .A2(n1140), .ZN(G51) );
XOR2_X1 U821 ( .A(n1141), .B(KEYINPUT2), .Z(n1140) );
NAND3_X1 U822 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
NAND2_X1 U823 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
OR3_X1 U824 ( .A1(n1146), .A2(n1145), .A3(KEYINPUT40), .ZN(n1143) );
AND2_X1 U825 ( .A1(KEYINPUT54), .A2(n1147), .ZN(n1145) );
NAND2_X1 U826 ( .A1(KEYINPUT40), .A2(n1148), .ZN(n1142) );
OR2_X1 U827 ( .A1(n1147), .A2(n1146), .ZN(n1148) );
XNOR2_X1 U828 ( .A(n1074), .B(n1149), .ZN(n1146) );
NAND2_X1 U829 ( .A1(n1085), .A2(n1046), .ZN(n1147) );
INV_X1 U830 ( .A(n1098), .ZN(n1085) );
NAND2_X1 U831 ( .A1(G902), .A2(n1092), .ZN(n1098) );
NAND3_X1 U832 ( .A1(n1070), .A2(n989), .A3(n1150), .ZN(n1092) );
AND3_X1 U833 ( .A1(n990), .A2(n1026), .A3(n1024), .ZN(n1150) );
AND4_X1 U834 ( .A1(n1151), .A2(n1152), .A3(n1102), .A4(n1153), .ZN(n989) );
AND4_X1 U835 ( .A1(n1154), .A2(n1155), .A3(n981), .A4(n1156), .ZN(n1153) );
NAND3_X1 U836 ( .A1(n1004), .A2(n1157), .A3(n1015), .ZN(n981) );
NAND3_X1 U837 ( .A1(n1004), .A2(n1157), .A3(n1016), .ZN(n1102) );
INV_X1 U838 ( .A(n985), .ZN(n1070) );
NAND4_X1 U839 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n985) );
NOR3_X1 U840 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1161) );
NAND3_X1 U841 ( .A1(n1016), .A2(n1165), .A3(n1023), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1027), .A2(G952), .ZN(n1081) );
XOR2_X1 U843 ( .A(n1166), .B(G146), .Z(G48) );
NAND2_X1 U844 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND3_X1 U845 ( .A1(n1000), .A2(n1169), .A3(n1170), .ZN(n1168) );
NAND2_X1 U846 ( .A1(n1016), .A2(n1171), .ZN(n1169) );
OR2_X1 U847 ( .A1(n1024), .A2(n1170), .ZN(n1167) );
INV_X1 U848 ( .A(KEYINPUT62), .ZN(n1170) );
NAND3_X1 U849 ( .A1(n1171), .A2(n1000), .A3(n1016), .ZN(n1024) );
XOR2_X1 U850 ( .A(n1172), .B(n1026), .Z(G45) );
NAND4_X1 U851 ( .A1(n1173), .A2(n1165), .A3(n1000), .A4(n1174), .ZN(n1026) );
XNOR2_X1 U852 ( .A(n1158), .B(n1175), .ZN(G42) );
XOR2_X1 U853 ( .A(KEYINPUT32), .B(G140), .Z(n1175) );
NAND3_X1 U854 ( .A1(n1176), .A2(n1020), .A3(n1023), .ZN(n1158) );
XNOR2_X1 U855 ( .A(G137), .B(n1159), .ZN(G39) );
NAND3_X1 U856 ( .A1(n1023), .A2(n1171), .A3(n1177), .ZN(n1159) );
XOR2_X1 U857 ( .A(G134), .B(n1162), .Z(G36) );
AND3_X1 U858 ( .A1(n1165), .A2(n1015), .A3(n1023), .ZN(n1162) );
XNOR2_X1 U859 ( .A(G131), .B(n1178), .ZN(G33) );
NAND4_X1 U860 ( .A1(KEYINPUT20), .A2(n1023), .A3(n1016), .A4(n1165), .ZN(n1178) );
AND4_X1 U861 ( .A1(n1179), .A2(n1020), .A3(n1009), .A4(n1036), .ZN(n1165) );
NOR2_X1 U862 ( .A1(n1002), .A2(n1033), .ZN(n1023) );
INV_X1 U863 ( .A(n1003), .ZN(n1033) );
XOR2_X1 U864 ( .A(G128), .B(n1164), .Z(G30) );
AND3_X1 U865 ( .A1(n1015), .A2(n1000), .A3(n1171), .ZN(n1164) );
AND4_X1 U866 ( .A1(n1180), .A2(n1179), .A3(n1020), .A4(n1181), .ZN(n1171) );
XOR2_X1 U867 ( .A(n990), .B(n1182), .Z(G3) );
XNOR2_X1 U868 ( .A(G101), .B(KEYINPUT50), .ZN(n1182) );
NAND4_X1 U869 ( .A1(n1177), .A2(n1157), .A3(n1009), .A4(n1036), .ZN(n990) );
INV_X1 U870 ( .A(n1008), .ZN(n1036) );
XOR2_X1 U871 ( .A(G125), .B(n1163), .Z(G27) );
AND3_X1 U872 ( .A1(n1030), .A2(n1000), .A3(n1176), .ZN(n1163) );
AND4_X1 U873 ( .A1(n1016), .A2(n1179), .A3(n1008), .A4(n1181), .ZN(n1176) );
AND3_X1 U874 ( .A1(n1183), .A2(n1184), .A3(n993), .ZN(n1179) );
NAND2_X1 U875 ( .A1(n1028), .A2(n1027), .ZN(n1184) );
INV_X1 U876 ( .A(G952), .ZN(n1028) );
NAND2_X1 U877 ( .A1(G953), .A2(n1185), .ZN(n1183) );
NAND2_X1 U878 ( .A1(G902), .A2(n1052), .ZN(n1185) );
INV_X1 U879 ( .A(G900), .ZN(n1052) );
XOR2_X1 U880 ( .A(n1151), .B(n1186), .Z(G24) );
NOR2_X1 U881 ( .A1(G122), .A2(KEYINPUT16), .ZN(n1186) );
NAND4_X1 U882 ( .A1(n1187), .A2(n1174), .A3(n1004), .A4(n1188), .ZN(n1151) );
NOR2_X1 U883 ( .A1(n1014), .A2(n1189), .ZN(n1188) );
INV_X1 U884 ( .A(n999), .ZN(n1004) );
NAND2_X1 U885 ( .A1(n1008), .A2(n1009), .ZN(n999) );
XNOR2_X1 U886 ( .A(G119), .B(n1152), .ZN(G21) );
NAND4_X1 U887 ( .A1(n1180), .A2(n1190), .A3(n1187), .A4(n1181), .ZN(n1152) );
INV_X1 U888 ( .A(n996), .ZN(n1190) );
NAND2_X1 U889 ( .A1(n1177), .A2(n1030), .ZN(n996) );
XOR2_X1 U890 ( .A(n1008), .B(KEYINPUT8), .Z(n1180) );
XOR2_X1 U891 ( .A(n1191), .B(n1155), .Z(G18) );
NAND3_X1 U892 ( .A1(n1015), .A2(n1187), .A3(n1192), .ZN(n1155) );
NOR2_X1 U893 ( .A1(n1193), .A2(n1173), .ZN(n1015) );
XNOR2_X1 U894 ( .A(G113), .B(n1154), .ZN(G15) );
NAND3_X1 U895 ( .A1(n1016), .A2(n1187), .A3(n1192), .ZN(n1154) );
NOR3_X1 U896 ( .A1(n1181), .A2(n1008), .A3(n1014), .ZN(n1192) );
INV_X1 U897 ( .A(n1030), .ZN(n1014) );
NOR2_X1 U898 ( .A1(n1194), .A2(n1195), .ZN(n1030) );
AND2_X1 U899 ( .A1(G221), .A2(n1022), .ZN(n1195) );
NOR2_X1 U900 ( .A1(n1189), .A2(n1174), .ZN(n1016) );
INV_X1 U901 ( .A(n1193), .ZN(n1174) );
XOR2_X1 U902 ( .A(n1196), .B(n1156), .Z(G12) );
NAND4_X1 U903 ( .A1(n1177), .A2(n1157), .A3(n1008), .A4(n1181), .ZN(n1156) );
INV_X1 U904 ( .A(n1009), .ZN(n1181) );
XOR2_X1 U905 ( .A(n1037), .B(KEYINPUT15), .Z(n1009) );
XOR2_X1 U906 ( .A(n1197), .B(n1198), .Z(n1037) );
AND2_X1 U907 ( .A1(n1022), .A2(G217), .ZN(n1198) );
NAND2_X1 U908 ( .A1(n1086), .A2(n1199), .ZN(n1197) );
XOR2_X1 U909 ( .A(n1200), .B(n1201), .Z(n1086) );
XOR2_X1 U910 ( .A(n1202), .B(n1203), .Z(n1201) );
XOR2_X1 U911 ( .A(G137), .B(G119), .Z(n1203) );
NOR2_X1 U912 ( .A1(G125), .A2(KEYINPUT6), .ZN(n1202) );
XOR2_X1 U913 ( .A(n1204), .B(n1205), .Z(n1200) );
INV_X1 U914 ( .A(n1133), .ZN(n1205) );
XOR2_X1 U915 ( .A(n1196), .B(G140), .Z(n1133) );
XOR2_X1 U916 ( .A(n1206), .B(n1207), .Z(n1204) );
NAND2_X1 U917 ( .A1(G221), .A2(n1208), .ZN(n1206) );
XOR2_X1 U918 ( .A(n1209), .B(G472), .Z(n1008) );
NAND2_X1 U919 ( .A1(n1210), .A2(n1199), .ZN(n1209) );
XOR2_X1 U920 ( .A(n1211), .B(n1212), .Z(n1210) );
XNOR2_X1 U921 ( .A(n1123), .B(n1213), .ZN(n1212) );
XNOR2_X1 U922 ( .A(KEYINPUT9), .B(n1110), .ZN(n1213) );
NAND3_X1 U923 ( .A1(n1214), .A2(n1027), .A3(G210), .ZN(n1110) );
NAND2_X1 U924 ( .A1(n1215), .A2(n1191), .ZN(n1123) );
INV_X1 U925 ( .A(G116), .ZN(n1191) );
XNOR2_X1 U926 ( .A(KEYINPUT5), .B(KEYINPUT38), .ZN(n1215) );
XOR2_X1 U927 ( .A(n1216), .B(n1217), .Z(n1211) );
XOR2_X1 U928 ( .A(n1129), .B(n1066), .Z(n1216) );
AND2_X1 U929 ( .A1(n1187), .A2(n1020), .ZN(n1157) );
AND2_X1 U930 ( .A1(n1194), .A2(n1218), .ZN(n1020) );
NAND2_X1 U931 ( .A1(G221), .A2(n1022), .ZN(n1218) );
NAND2_X1 U932 ( .A1(n1219), .A2(n1199), .ZN(n1022) );
INV_X1 U933 ( .A(n1021), .ZN(n1194) );
XOR2_X1 U934 ( .A(n1220), .B(G469), .Z(n1021) );
NAND2_X1 U935 ( .A1(n1221), .A2(n1199), .ZN(n1220) );
XOR2_X1 U936 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U937 ( .A(n1224), .B(n1135), .Z(n1223) );
XOR2_X1 U938 ( .A(n1066), .B(n1225), .Z(n1135) );
XOR2_X1 U939 ( .A(G101), .B(n1226), .Z(n1225) );
NOR2_X1 U940 ( .A1(KEYINPUT29), .A2(n1227), .ZN(n1226) );
XOR2_X1 U941 ( .A(KEYINPUT7), .B(n1228), .Z(n1227) );
INV_X1 U942 ( .A(n1121), .ZN(n1066) );
XNOR2_X1 U943 ( .A(G131), .B(n1067), .ZN(n1121) );
XOR2_X1 U944 ( .A(G134), .B(G137), .Z(n1067) );
NOR2_X1 U945 ( .A1(KEYINPUT51), .A2(n1063), .ZN(n1224) );
XNOR2_X1 U946 ( .A(G143), .B(n1207), .ZN(n1063) );
XOR2_X1 U947 ( .A(G128), .B(G146), .Z(n1207) );
XOR2_X1 U948 ( .A(n1229), .B(n1230), .Z(n1222) );
XOR2_X1 U949 ( .A(G227), .B(G110), .Z(n1230) );
NOR2_X1 U950 ( .A1(G140), .A2(KEYINPUT22), .ZN(n1229) );
AND3_X1 U951 ( .A1(n1231), .A2(n993), .A3(n1000), .ZN(n1187) );
AND2_X1 U952 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NAND2_X1 U953 ( .A1(G214), .A2(n1232), .ZN(n1003) );
XOR2_X1 U954 ( .A(n1045), .B(n1233), .Z(n1002) );
NOR2_X1 U955 ( .A1(n1046), .A2(KEYINPUT34), .ZN(n1233) );
AND2_X1 U956 ( .A1(G210), .A2(n1232), .ZN(n1046) );
NAND2_X1 U957 ( .A1(n1214), .A2(n1199), .ZN(n1232) );
NAND3_X1 U958 ( .A1(n1234), .A2(n1199), .A3(n1235), .ZN(n1045) );
NAND2_X1 U959 ( .A1(n1236), .A2(n1149), .ZN(n1235) );
XOR2_X1 U960 ( .A(KEYINPUT23), .B(n1237), .Z(n1236) );
INV_X1 U961 ( .A(n1074), .ZN(n1237) );
INV_X1 U962 ( .A(G902), .ZN(n1199) );
NAND2_X1 U963 ( .A1(n1238), .A2(n1239), .ZN(n1234) );
XNOR2_X1 U964 ( .A(n1149), .B(KEYINPUT19), .ZN(n1239) );
XNOR2_X1 U965 ( .A(n1129), .B(n1240), .ZN(n1149) );
XOR2_X1 U966 ( .A(G125), .B(n1241), .Z(n1240) );
NOR2_X1 U967 ( .A1(G953), .A2(n1078), .ZN(n1241) );
INV_X1 U968 ( .A(G224), .ZN(n1078) );
XOR2_X1 U969 ( .A(n1242), .B(G128), .Z(n1129) );
NAND2_X1 U970 ( .A1(n1243), .A2(KEYINPUT21), .ZN(n1242) );
XOR2_X1 U971 ( .A(n1244), .B(G143), .Z(n1243) );
XOR2_X1 U972 ( .A(n1074), .B(KEYINPUT30), .Z(n1238) );
XOR2_X1 U973 ( .A(n1245), .B(n1246), .Z(n1074) );
XNOR2_X1 U974 ( .A(n1217), .B(n1247), .ZN(n1246) );
XOR2_X1 U975 ( .A(G101), .B(n1124), .Z(n1217) );
XOR2_X1 U976 ( .A(G119), .B(G113), .Z(n1124) );
XOR2_X1 U977 ( .A(n1248), .B(n1228), .Z(n1245) );
XOR2_X1 U978 ( .A(G107), .B(G104), .Z(n1228) );
NAND2_X1 U979 ( .A1(KEYINPUT43), .A2(n1196), .ZN(n1248) );
NAND2_X1 U980 ( .A1(G237), .A2(n1219), .ZN(n993) );
XNOR2_X1 U981 ( .A(G234), .B(KEYINPUT53), .ZN(n1219) );
NAND2_X1 U982 ( .A1(n1249), .A2(n1250), .ZN(n1231) );
NAND2_X1 U983 ( .A1(G902), .A2(n1073), .ZN(n1250) );
NOR2_X1 U984 ( .A1(G898), .A2(n1027), .ZN(n1073) );
NAND2_X1 U985 ( .A1(G952), .A2(n1027), .ZN(n1249) );
INV_X1 U986 ( .A(n1018), .ZN(n1177) );
NAND2_X1 U987 ( .A1(n1189), .A2(n1193), .ZN(n1018) );
NAND2_X1 U988 ( .A1(n1251), .A2(n1252), .ZN(n1193) );
NAND2_X1 U989 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
INV_X1 U990 ( .A(n1044), .ZN(n1254) );
NAND2_X1 U991 ( .A1(KEYINPUT58), .A2(n1255), .ZN(n1253) );
NAND2_X1 U992 ( .A1(KEYINPUT18), .A2(n1042), .ZN(n1255) );
INV_X1 U993 ( .A(G478), .ZN(n1042) );
NAND2_X1 U994 ( .A1(G478), .A2(n1256), .ZN(n1251) );
NAND2_X1 U995 ( .A1(KEYINPUT18), .A2(n1257), .ZN(n1256) );
NAND2_X1 U996 ( .A1(n1044), .A2(KEYINPUT58), .ZN(n1257) );
NOR2_X1 U997 ( .A1(n1090), .A2(G902), .ZN(n1044) );
XNOR2_X1 U998 ( .A(n1258), .B(n1259), .ZN(n1090) );
XOR2_X1 U999 ( .A(G107), .B(n1260), .Z(n1259) );
NOR2_X1 U1000 ( .A1(KEYINPUT3), .A2(n1247), .ZN(n1260) );
XNOR2_X1 U1001 ( .A(G116), .B(G122), .ZN(n1247) );
XOR2_X1 U1002 ( .A(n1261), .B(n1262), .Z(n1258) );
NOR2_X1 U1003 ( .A1(KEYINPUT36), .A2(n1263), .ZN(n1262) );
XOR2_X1 U1004 ( .A(n1264), .B(G134), .Z(n1263) );
NAND2_X1 U1005 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U1006 ( .A1(G128), .A2(n1172), .ZN(n1266) );
INV_X1 U1007 ( .A(G143), .ZN(n1172) );
XOR2_X1 U1008 ( .A(n1267), .B(KEYINPUT11), .Z(n1265) );
NAND2_X1 U1009 ( .A1(G143), .A2(n1268), .ZN(n1267) );
INV_X1 U1010 ( .A(G128), .ZN(n1268) );
NAND2_X1 U1011 ( .A1(G217), .A2(n1208), .ZN(n1261) );
AND2_X1 U1012 ( .A1(G234), .A2(n1027), .ZN(n1208) );
INV_X1 U1013 ( .A(n1173), .ZN(n1189) );
XNOR2_X1 U1014 ( .A(n1047), .B(n1269), .ZN(n1173) );
NOR2_X1 U1015 ( .A1(G475), .A2(KEYINPUT10), .ZN(n1269) );
NOR2_X1 U1016 ( .A1(n1099), .A2(G902), .ZN(n1047) );
XOR2_X1 U1017 ( .A(n1270), .B(n1271), .Z(n1099) );
XOR2_X1 U1018 ( .A(n1060), .B(n1272), .Z(n1271) );
XOR2_X1 U1019 ( .A(n1273), .B(n1274), .Z(n1272) );
AND3_X1 U1020 ( .A1(G214), .A2(n1027), .A3(n1214), .ZN(n1274) );
INV_X1 U1021 ( .A(G237), .ZN(n1214) );
INV_X1 U1022 ( .A(G953), .ZN(n1027) );
NAND2_X1 U1023 ( .A1(KEYINPUT41), .A2(n1244), .ZN(n1273) );
INV_X1 U1024 ( .A(G146), .ZN(n1244) );
XOR2_X1 U1025 ( .A(n1275), .B(G140), .Z(n1060) );
INV_X1 U1026 ( .A(G125), .ZN(n1275) );
XOR2_X1 U1027 ( .A(n1276), .B(n1277), .Z(n1270) );
XOR2_X1 U1028 ( .A(KEYINPUT57), .B(G143), .Z(n1277) );
XNOR2_X1 U1029 ( .A(G131), .B(n1278), .ZN(n1276) );
NOR2_X1 U1030 ( .A1(KEYINPUT45), .A2(n1279), .ZN(n1278) );
NOR2_X1 U1031 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
XOR2_X1 U1032 ( .A(KEYINPUT55), .B(n1282), .Z(n1281) );
AND2_X1 U1033 ( .A1(n1283), .A2(G104), .ZN(n1282) );
NOR2_X1 U1034 ( .A1(G104), .A2(n1283), .ZN(n1280) );
XOR2_X1 U1035 ( .A(G122), .B(n1284), .Z(n1283) );
NOR2_X1 U1036 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NOR2_X1 U1037 ( .A1(KEYINPUT48), .A2(G113), .ZN(n1286) );
AND2_X1 U1038 ( .A1(KEYINPUT26), .A2(G113), .ZN(n1285) );
INV_X1 U1039 ( .A(G110), .ZN(n1196) );
endmodule


