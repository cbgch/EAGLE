//Key = 1000010011011101001000010010001000011100101010000011000110001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;

XNOR2_X1 U729 ( .A(n1000), .B(n1001), .ZN(G9) );
NAND4_X1 U730 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(G75) );
INV_X1 U731 ( .A(n1006), .ZN(n1005) );
NAND3_X1 U732 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1004) );
NAND2_X1 U733 ( .A1(n1010), .A2(n1011), .ZN(n1007) );
NAND4_X1 U734 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
NOR2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
XNOR2_X1 U736 ( .A(KEYINPUT57), .B(n1018), .ZN(n1017) );
XNOR2_X1 U737 ( .A(G469), .B(n1019), .ZN(n1016) );
NAND4_X1 U738 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1010) );
NAND2_X1 U739 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND2_X1 U740 ( .A1(G952), .A2(n1026), .ZN(n1003) );
NAND4_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
NAND3_X1 U742 ( .A1(n1021), .A2(n1031), .A3(n1032), .ZN(n1030) );
NAND3_X1 U743 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1031) );
NAND3_X1 U744 ( .A1(n1036), .A2(n1008), .A3(n1022), .ZN(n1035) );
NAND3_X1 U745 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1020), .ZN(n1039) );
NAND3_X1 U747 ( .A1(n1009), .A2(n1041), .A3(n1042), .ZN(n1037) );
NAND2_X1 U748 ( .A1(n1009), .A2(n1043), .ZN(n1034) );
NAND2_X1 U749 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U750 ( .A1(n1046), .A2(n1020), .ZN(n1045) );
XNOR2_X1 U751 ( .A(n1022), .B(n1047), .ZN(n1046) );
NAND2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1044) );
INV_X1 U753 ( .A(KEYINPUT22), .ZN(n1049) );
NAND3_X1 U754 ( .A1(KEYINPUT22), .A2(n1048), .A3(n1050), .ZN(n1033) );
INV_X1 U755 ( .A(n1009), .ZN(n1050) );
INV_X1 U756 ( .A(n1051), .ZN(n1021) );
NAND2_X1 U757 ( .A1(KEYINPUT17), .A2(n1052), .ZN(n1029) );
OR2_X1 U758 ( .A1(n1052), .A2(KEYINPUT17), .ZN(n1002) );
XOR2_X1 U759 ( .A(n1053), .B(n1054), .Z(G72) );
NOR2_X1 U760 ( .A1(n1052), .A2(n1055), .ZN(n1054) );
XOR2_X1 U761 ( .A(KEYINPUT31), .B(n1056), .Z(n1055) );
NOR2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1053) );
NAND2_X1 U764 ( .A1(n1061), .A2(n1052), .ZN(n1060) );
XNOR2_X1 U765 ( .A(n1062), .B(n1028), .ZN(n1061) );
NAND3_X1 U766 ( .A1(G900), .A2(n1062), .A3(G953), .ZN(n1059) );
XNOR2_X1 U767 ( .A(n1063), .B(n1064), .ZN(n1062) );
XOR2_X1 U768 ( .A(G131), .B(n1065), .Z(n1064) );
XNOR2_X1 U769 ( .A(KEYINPUT43), .B(n1066), .ZN(n1065) );
XNOR2_X1 U770 ( .A(n1067), .B(n1068), .ZN(n1063) );
XOR2_X1 U771 ( .A(n1069), .B(n1070), .Z(n1068) );
NAND2_X1 U772 ( .A1(KEYINPUT44), .A2(n1071), .ZN(n1070) );
NAND2_X1 U773 ( .A1(KEYINPUT18), .A2(n1072), .ZN(n1069) );
XOR2_X1 U774 ( .A(n1073), .B(n1074), .Z(G69) );
XOR2_X1 U775 ( .A(n1075), .B(n1076), .Z(n1074) );
NAND2_X1 U776 ( .A1(G953), .A2(n1077), .ZN(n1076) );
NAND2_X1 U777 ( .A1(G898), .A2(G224), .ZN(n1077) );
NAND2_X1 U778 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
NAND2_X1 U779 ( .A1(n1080), .A2(G953), .ZN(n1079) );
XOR2_X1 U780 ( .A(n1081), .B(n1082), .Z(n1078) );
NAND2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
XNOR2_X1 U782 ( .A(KEYINPUT46), .B(KEYINPUT34), .ZN(n1083) );
NOR2_X1 U783 ( .A1(n1027), .A2(G953), .ZN(n1073) );
NOR2_X1 U784 ( .A1(n1006), .A2(n1085), .ZN(G66) );
XNOR2_X1 U785 ( .A(n1086), .B(n1087), .ZN(n1085) );
NOR2_X1 U786 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U787 ( .A1(n1006), .A2(n1090), .ZN(G63) );
XNOR2_X1 U788 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR2_X1 U789 ( .A1(n1093), .A2(n1089), .ZN(n1092) );
NOR2_X1 U790 ( .A1(n1006), .A2(n1094), .ZN(G60) );
XOR2_X1 U791 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U792 ( .A1(n1097), .A2(n1089), .ZN(n1095) );
XNOR2_X1 U793 ( .A(G104), .B(n1098), .ZN(G6) );
NOR2_X1 U794 ( .A1(n1099), .A2(KEYINPUT45), .ZN(n1098) );
NOR2_X1 U795 ( .A1(n1006), .A2(n1100), .ZN(G57) );
XOR2_X1 U796 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U797 ( .A(n1103), .B(n1104), .ZN(n1102) );
NAND2_X1 U798 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U799 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U800 ( .A(n1109), .B(KEYINPUT2), .ZN(n1107) );
NAND2_X1 U801 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
XNOR2_X1 U802 ( .A(KEYINPUT32), .B(n1112), .ZN(n1110) );
XOR2_X1 U803 ( .A(n1113), .B(n1114), .Z(n1101) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1089), .ZN(n1114) );
NAND2_X1 U805 ( .A1(KEYINPUT56), .A2(n1116), .ZN(n1113) );
NOR2_X1 U806 ( .A1(n1117), .A2(n1118), .ZN(G54) );
XOR2_X1 U807 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U808 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U809 ( .A1(n1123), .A2(n1089), .ZN(n1122) );
INV_X1 U810 ( .A(G469), .ZN(n1123) );
XOR2_X1 U811 ( .A(n1124), .B(n1125), .Z(n1119) );
NOR2_X1 U812 ( .A1(KEYINPUT19), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U813 ( .A(n1127), .B(n1108), .ZN(n1126) );
NAND2_X1 U814 ( .A1(n1128), .A2(KEYINPUT12), .ZN(n1127) );
XOR2_X1 U815 ( .A(n1129), .B(n1067), .Z(n1128) );
NAND2_X1 U816 ( .A1(KEYINPUT51), .A2(n1130), .ZN(n1129) );
XNOR2_X1 U817 ( .A(G140), .B(KEYINPUT52), .ZN(n1124) );
NOR2_X1 U818 ( .A1(n1052), .A2(n1131), .ZN(n1117) );
XOR2_X1 U819 ( .A(KEYINPUT7), .B(G952), .Z(n1131) );
NOR2_X1 U820 ( .A1(n1006), .A2(n1132), .ZN(G51) );
XOR2_X1 U821 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U822 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND2_X1 U823 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
OR2_X1 U824 ( .A1(KEYINPUT24), .A2(n1139), .ZN(n1138) );
NAND2_X1 U825 ( .A1(KEYINPUT53), .A2(n1139), .ZN(n1137) );
XOR2_X1 U826 ( .A(n1140), .B(n1141), .Z(n1133) );
NOR2_X1 U827 ( .A1(n1142), .A2(n1089), .ZN(n1141) );
NAND2_X1 U828 ( .A1(G902), .A2(n1143), .ZN(n1089) );
NAND2_X1 U829 ( .A1(n1027), .A2(n1028), .ZN(n1143) );
AND4_X1 U830 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1028) );
NOR4_X1 U831 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1147) );
INV_X1 U832 ( .A(n1152), .ZN(n1151) );
NAND2_X1 U833 ( .A1(n1020), .A2(n1153), .ZN(n1146) );
NAND2_X1 U834 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U835 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
AND4_X1 U836 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1027) );
NOR4_X1 U837 ( .A1(n1099), .A2(n1001), .A3(n1162), .A4(n1163), .ZN(n1161) );
AND3_X1 U838 ( .A1(n1009), .A2(n1164), .A3(n1165), .ZN(n1001) );
AND3_X1 U839 ( .A1(n1165), .A2(n1009), .A3(n1166), .ZN(n1099) );
NOR2_X1 U840 ( .A1(n1167), .A2(n1168), .ZN(n1160) );
NOR2_X1 U841 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U842 ( .A(KEYINPUT5), .B(n1171), .Z(n1170) );
NOR4_X1 U843 ( .A1(n1172), .A2(n1173), .A3(n1025), .A4(n1174), .ZN(n1171) );
NAND2_X1 U844 ( .A1(n1008), .A2(n1175), .ZN(n1173) );
NOR2_X1 U845 ( .A1(n1052), .A2(G952), .ZN(n1006) );
XNOR2_X1 U846 ( .A(G146), .B(n1144), .ZN(G48) );
NAND2_X1 U847 ( .A1(n1176), .A2(n1166), .ZN(n1144) );
XNOR2_X1 U848 ( .A(G143), .B(n1145), .ZN(G45) );
NAND3_X1 U849 ( .A1(n1156), .A2(n1040), .A3(n1177), .ZN(n1145) );
NOR3_X1 U850 ( .A1(n1169), .A2(n1018), .A3(n1014), .ZN(n1177) );
NAND2_X1 U851 ( .A1(n1178), .A2(n1179), .ZN(G42) );
NAND2_X1 U852 ( .A1(n1180), .A2(n1066), .ZN(n1179) );
XNOR2_X1 U853 ( .A(n1150), .B(KEYINPUT26), .ZN(n1180) );
NAND2_X1 U854 ( .A1(n1181), .A2(G140), .ZN(n1178) );
XNOR2_X1 U855 ( .A(n1150), .B(KEYINPUT54), .ZN(n1181) );
NOR3_X1 U856 ( .A1(n1182), .A2(n1024), .A3(n1038), .ZN(n1150) );
NAND3_X1 U857 ( .A1(n1183), .A2(n1184), .A3(n1020), .ZN(n1038) );
INV_X1 U858 ( .A(n1166), .ZN(n1024) );
XOR2_X1 U859 ( .A(G137), .B(n1185), .Z(G39) );
NOR3_X1 U860 ( .A1(n1182), .A2(n1186), .A3(n1187), .ZN(n1185) );
XNOR2_X1 U861 ( .A(n1020), .B(KEYINPUT3), .ZN(n1186) );
XOR2_X1 U862 ( .A(G134), .B(n1149), .Z(G36) );
NOR4_X1 U863 ( .A1(n1182), .A2(n1174), .A3(n1188), .A4(n1025), .ZN(n1149) );
INV_X1 U864 ( .A(n1164), .ZN(n1025) );
INV_X1 U865 ( .A(n1040), .ZN(n1174) );
NAND2_X1 U866 ( .A1(n1189), .A2(n1190), .ZN(G33) );
NAND2_X1 U867 ( .A1(G131), .A2(n1191), .ZN(n1190) );
XOR2_X1 U868 ( .A(KEYINPUT23), .B(n1192), .Z(n1189) );
NOR2_X1 U869 ( .A1(G131), .A2(n1191), .ZN(n1192) );
NAND2_X1 U870 ( .A1(n1193), .A2(n1020), .ZN(n1191) );
INV_X1 U871 ( .A(n1188), .ZN(n1020) );
NAND2_X1 U872 ( .A1(n1041), .A2(n1013), .ZN(n1188) );
XOR2_X1 U873 ( .A(n1155), .B(KEYINPUT0), .Z(n1193) );
NAND3_X1 U874 ( .A1(n1040), .A2(n1166), .A3(n1156), .ZN(n1155) );
XOR2_X1 U875 ( .A(G128), .B(n1148), .Z(G30) );
AND2_X1 U876 ( .A1(n1176), .A2(n1164), .ZN(n1148) );
NOR4_X1 U877 ( .A1(n1182), .A2(n1169), .A3(n1183), .A4(n1194), .ZN(n1176) );
INV_X1 U878 ( .A(n1156), .ZN(n1182) );
NOR3_X1 U879 ( .A1(n1195), .A2(n1047), .A3(n1022), .ZN(n1156) );
XOR2_X1 U880 ( .A(G101), .B(n1196), .Z(G3) );
NOR2_X1 U881 ( .A1(KEYINPUT48), .A2(n1158), .ZN(n1196) );
NAND3_X1 U882 ( .A1(n1032), .A2(n1165), .A3(n1040), .ZN(n1158) );
XNOR2_X1 U883 ( .A(n1071), .B(n1197), .ZN(G27) );
NOR2_X1 U884 ( .A1(KEYINPUT10), .A2(n1152), .ZN(n1197) );
NAND3_X1 U885 ( .A1(n1048), .A2(n1166), .A3(n1198), .ZN(n1152) );
NOR3_X1 U886 ( .A1(n1199), .A2(n1195), .A3(n1194), .ZN(n1198) );
INV_X1 U887 ( .A(n1184), .ZN(n1194) );
AND2_X1 U888 ( .A1(n1051), .A2(n1200), .ZN(n1195) );
NAND4_X1 U889 ( .A1(G902), .A2(G953), .A3(n1201), .A4(n1058), .ZN(n1200) );
INV_X1 U890 ( .A(G900), .ZN(n1058) );
XNOR2_X1 U891 ( .A(G122), .B(n1159), .ZN(G24) );
NAND4_X1 U892 ( .A1(n1202), .A2(n1009), .A3(n1203), .A4(n1204), .ZN(n1159) );
NOR2_X1 U893 ( .A1(n1184), .A2(n1199), .ZN(n1009) );
XOR2_X1 U894 ( .A(n1205), .B(G119), .Z(G21) );
NAND2_X1 U895 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U896 ( .A1(n1167), .A2(n1208), .ZN(n1207) );
INV_X1 U897 ( .A(KEYINPUT29), .ZN(n1208) );
AND2_X1 U898 ( .A1(n1157), .A2(n1202), .ZN(n1167) );
NAND4_X1 U899 ( .A1(n1157), .A2(n1048), .A3(n1209), .A4(KEYINPUT29), .ZN(n1206) );
INV_X1 U900 ( .A(n1187), .ZN(n1157) );
NAND3_X1 U901 ( .A1(n1199), .A2(n1184), .A3(n1032), .ZN(n1187) );
XNOR2_X1 U902 ( .A(G116), .B(n1210), .ZN(G18) );
NAND4_X1 U903 ( .A1(n1040), .A2(n1048), .A3(n1164), .A4(n1211), .ZN(n1210) );
XNOR2_X1 U904 ( .A(KEYINPUT40), .B(n1175), .ZN(n1211) );
NOR2_X1 U905 ( .A1(n1203), .A2(n1018), .ZN(n1164) );
INV_X1 U906 ( .A(n1204), .ZN(n1018) );
XOR2_X1 U907 ( .A(G113), .B(n1163), .Z(G15) );
AND3_X1 U908 ( .A1(n1202), .A2(n1166), .A3(n1040), .ZN(n1163) );
NOR2_X1 U909 ( .A1(n1184), .A2(n1183), .ZN(n1040) );
NOR2_X1 U910 ( .A1(n1204), .A2(n1014), .ZN(n1166) );
INV_X1 U911 ( .A(n1203), .ZN(n1014) );
AND2_X1 U912 ( .A1(n1048), .A2(n1175), .ZN(n1202) );
NOR3_X1 U913 ( .A1(n1172), .A2(n1047), .A3(n1169), .ZN(n1048) );
INV_X1 U914 ( .A(n1022), .ZN(n1172) );
XOR2_X1 U915 ( .A(G110), .B(n1162), .Z(G12) );
AND4_X1 U916 ( .A1(n1032), .A2(n1165), .A3(n1183), .A4(n1184), .ZN(n1162) );
XOR2_X1 U917 ( .A(n1212), .B(n1088), .Z(n1184) );
NAND2_X1 U918 ( .A1(G217), .A2(n1213), .ZN(n1088) );
NAND2_X1 U919 ( .A1(n1086), .A2(n1214), .ZN(n1212) );
XNOR2_X1 U920 ( .A(n1215), .B(n1216), .ZN(n1086) );
XNOR2_X1 U921 ( .A(n1217), .B(n1218), .ZN(n1216) );
XOR2_X1 U922 ( .A(n1219), .B(n1220), .Z(n1215) );
XNOR2_X1 U923 ( .A(G137), .B(n1221), .ZN(n1220) );
NAND3_X1 U924 ( .A1(n1222), .A2(n1223), .A3(KEYINPUT15), .ZN(n1221) );
NAND2_X1 U925 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
XOR2_X1 U926 ( .A(KEYINPUT11), .B(n1226), .Z(n1222) );
NOR2_X1 U927 ( .A1(n1225), .A2(n1224), .ZN(n1226) );
XOR2_X1 U928 ( .A(KEYINPUT21), .B(G110), .Z(n1224) );
XOR2_X1 U929 ( .A(G119), .B(G128), .Z(n1225) );
NAND3_X1 U930 ( .A1(n1227), .A2(G221), .A3(KEYINPUT36), .ZN(n1219) );
INV_X1 U931 ( .A(n1199), .ZN(n1183) );
XOR2_X1 U932 ( .A(n1228), .B(n1115), .Z(n1199) );
INV_X1 U933 ( .A(G472), .ZN(n1115) );
NAND2_X1 U934 ( .A1(n1229), .A2(n1214), .ZN(n1228) );
XOR2_X1 U935 ( .A(n1230), .B(n1231), .Z(n1229) );
XNOR2_X1 U936 ( .A(n1232), .B(n1233), .ZN(n1231) );
XNOR2_X1 U937 ( .A(n1116), .B(n1111), .ZN(n1233) );
XOR2_X1 U938 ( .A(n1234), .B(G101), .Z(n1116) );
NAND2_X1 U939 ( .A1(n1235), .A2(G210), .ZN(n1234) );
INV_X1 U940 ( .A(n1103), .ZN(n1232) );
XOR2_X1 U941 ( .A(G116), .B(n1236), .Z(n1103) );
XNOR2_X1 U942 ( .A(n1109), .B(n1237), .ZN(n1230) );
XOR2_X1 U943 ( .A(KEYINPUT59), .B(KEYINPUT49), .Z(n1237) );
NOR4_X1 U944 ( .A1(n1022), .A2(n1169), .A3(n1047), .A4(n1209), .ZN(n1165) );
INV_X1 U945 ( .A(n1175), .ZN(n1209) );
NAND2_X1 U946 ( .A1(n1238), .A2(n1239), .ZN(n1175) );
NAND4_X1 U947 ( .A1(n1080), .A2(G902), .A3(G953), .A4(n1201), .ZN(n1239) );
XNOR2_X1 U948 ( .A(G898), .B(KEYINPUT14), .ZN(n1080) );
XNOR2_X1 U949 ( .A(KEYINPUT35), .B(n1051), .ZN(n1238) );
NAND3_X1 U950 ( .A1(n1201), .A2(n1052), .A3(G952), .ZN(n1051) );
INV_X1 U951 ( .A(G953), .ZN(n1052) );
NAND2_X1 U952 ( .A1(G237), .A2(G234), .ZN(n1201) );
INV_X1 U953 ( .A(n1008), .ZN(n1047) );
NAND2_X1 U954 ( .A1(G221), .A2(n1213), .ZN(n1008) );
NAND2_X1 U955 ( .A1(G234), .A2(n1214), .ZN(n1213) );
OR2_X1 U956 ( .A1(n1041), .A2(n1042), .ZN(n1169) );
INV_X1 U957 ( .A(n1013), .ZN(n1042) );
NAND2_X1 U958 ( .A1(G214), .A2(n1240), .ZN(n1013) );
XNOR2_X1 U959 ( .A(n1012), .B(KEYINPUT37), .ZN(n1041) );
XNOR2_X1 U960 ( .A(n1241), .B(n1142), .ZN(n1012) );
NAND2_X1 U961 ( .A1(G210), .A2(n1240), .ZN(n1142) );
NAND2_X1 U962 ( .A1(n1242), .A2(n1214), .ZN(n1240) );
INV_X1 U963 ( .A(G237), .ZN(n1242) );
NAND2_X1 U964 ( .A1(n1243), .A2(n1214), .ZN(n1241) );
XOR2_X1 U965 ( .A(n1140), .B(n1244), .Z(n1243) );
XOR2_X1 U966 ( .A(n1139), .B(n1245), .Z(n1244) );
NOR3_X1 U967 ( .A1(KEYINPUT41), .A2(n1246), .A3(n1247), .ZN(n1245) );
NOR2_X1 U968 ( .A1(n1248), .A2(n1135), .ZN(n1247) );
XNOR2_X1 U969 ( .A(n1109), .B(G125), .ZN(n1135) );
INV_X1 U970 ( .A(KEYINPUT9), .ZN(n1248) );
NOR3_X1 U971 ( .A1(KEYINPUT9), .A2(n1112), .A3(n1071), .ZN(n1246) );
INV_X1 U972 ( .A(n1109), .ZN(n1112) );
XOR2_X1 U973 ( .A(n1249), .B(n1250), .Z(n1109) );
XOR2_X1 U974 ( .A(KEYINPUT1), .B(n1251), .Z(n1250) );
NAND2_X1 U975 ( .A1(G224), .A2(n1252), .ZN(n1139) );
XNOR2_X1 U976 ( .A(n1084), .B(n1082), .ZN(n1140) );
XNOR2_X1 U977 ( .A(n1253), .B(n1254), .ZN(n1082) );
NOR2_X1 U978 ( .A1(G110), .A2(KEYINPUT39), .ZN(n1254) );
XNOR2_X1 U979 ( .A(G122), .B(n1255), .ZN(n1253) );
NOR2_X1 U980 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U981 ( .A(KEYINPUT47), .B(n1258), .Z(n1257) );
NOR2_X1 U982 ( .A1(G101), .A2(n1259), .ZN(n1258) );
AND2_X1 U983 ( .A1(n1259), .A2(G101), .ZN(n1256) );
XNOR2_X1 U984 ( .A(G104), .B(n1000), .ZN(n1259) );
XNOR2_X1 U985 ( .A(n1260), .B(n1236), .ZN(n1084) );
XOR2_X1 U986 ( .A(G113), .B(G119), .Z(n1236) );
NAND2_X1 U987 ( .A1(KEYINPUT62), .A2(n1261), .ZN(n1260) );
XNOR2_X1 U988 ( .A(n1019), .B(n1262), .ZN(n1022) );
NOR2_X1 U989 ( .A1(G469), .A2(KEYINPUT4), .ZN(n1262) );
NAND3_X1 U990 ( .A1(n1263), .A2(n1214), .A3(n1264), .ZN(n1019) );
NAND3_X1 U991 ( .A1(n1108), .A2(KEYINPUT8), .A3(n1265), .ZN(n1264) );
XOR2_X1 U992 ( .A(n1266), .B(n1267), .Z(n1265) );
NAND2_X1 U993 ( .A1(n1268), .A2(KEYINPUT42), .ZN(n1266) );
INV_X1 U994 ( .A(n1269), .ZN(n1268) );
NAND2_X1 U995 ( .A1(n1270), .A2(n1271), .ZN(n1263) );
NAND2_X1 U996 ( .A1(KEYINPUT8), .A2(n1108), .ZN(n1271) );
INV_X1 U997 ( .A(n1111), .ZN(n1108) );
XNOR2_X1 U998 ( .A(G131), .B(n1072), .ZN(n1111) );
XNOR2_X1 U999 ( .A(G134), .B(G137), .ZN(n1072) );
XOR2_X1 U1000 ( .A(n1272), .B(n1267), .Z(n1270) );
XNOR2_X1 U1001 ( .A(n1121), .B(n1273), .ZN(n1267) );
NOR2_X1 U1002 ( .A1(KEYINPUT6), .A2(n1066), .ZN(n1273) );
INV_X1 U1003 ( .A(G140), .ZN(n1066) );
XNOR2_X1 U1004 ( .A(G110), .B(n1274), .ZN(n1121) );
NOR2_X1 U1005 ( .A1(n1275), .A2(n1057), .ZN(n1274) );
INV_X1 U1006 ( .A(G227), .ZN(n1057) );
NAND2_X1 U1007 ( .A1(KEYINPUT42), .A2(n1269), .ZN(n1272) );
XNOR2_X1 U1008 ( .A(n1067), .B(n1130), .ZN(n1269) );
XOR2_X1 U1009 ( .A(n1276), .B(n1277), .Z(n1130) );
NOR2_X1 U1010 ( .A1(G101), .A2(KEYINPUT38), .ZN(n1277) );
NAND2_X1 U1011 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
OR2_X1 U1012 ( .A1(n1000), .A2(G104), .ZN(n1279) );
XOR2_X1 U1013 ( .A(n1280), .B(KEYINPUT20), .Z(n1278) );
NAND2_X1 U1014 ( .A1(G104), .A2(n1000), .ZN(n1280) );
XNOR2_X1 U1015 ( .A(n1281), .B(n1282), .ZN(n1067) );
XOR2_X1 U1016 ( .A(KEYINPUT61), .B(G128), .Z(n1282) );
NAND2_X1 U1017 ( .A1(KEYINPUT50), .A2(n1283), .ZN(n1281) );
NAND2_X1 U1018 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U1019 ( .A1(n1217), .A2(n1286), .ZN(n1285) );
XNOR2_X1 U1020 ( .A(KEYINPUT60), .B(n1287), .ZN(n1286) );
INV_X1 U1021 ( .A(n1249), .ZN(n1217) );
XOR2_X1 U1022 ( .A(n1288), .B(KEYINPUT16), .Z(n1284) );
NAND2_X1 U1023 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XNOR2_X1 U1024 ( .A(n1249), .B(KEYINPUT63), .ZN(n1290) );
XNOR2_X1 U1025 ( .A(n1291), .B(KEYINPUT55), .ZN(n1289) );
NOR2_X1 U1026 ( .A1(n1204), .A2(n1203), .ZN(n1032) );
XOR2_X1 U1027 ( .A(n1292), .B(n1097), .Z(n1203) );
INV_X1 U1028 ( .A(G475), .ZN(n1097) );
OR2_X1 U1029 ( .A1(n1096), .A2(G902), .ZN(n1292) );
XNOR2_X1 U1030 ( .A(n1293), .B(n1294), .ZN(n1096) );
XOR2_X1 U1031 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1032 ( .A(G104), .B(n1297), .Z(n1296) );
NOR2_X1 U1033 ( .A1(KEYINPUT28), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U1034 ( .A(n1299), .B(n1249), .ZN(n1298) );
XOR2_X1 U1035 ( .A(G146), .B(KEYINPUT25), .Z(n1249) );
NAND2_X1 U1036 ( .A1(KEYINPUT30), .A2(n1218), .ZN(n1299) );
XNOR2_X1 U1037 ( .A(n1071), .B(G140), .ZN(n1218) );
INV_X1 U1038 ( .A(G125), .ZN(n1071) );
XOR2_X1 U1039 ( .A(G131), .B(G122), .Z(n1295) );
XNOR2_X1 U1040 ( .A(n1300), .B(n1287), .ZN(n1293) );
INV_X1 U1041 ( .A(n1291), .ZN(n1287) );
XOR2_X1 U1042 ( .A(n1301), .B(n1302), .Z(n1300) );
NOR2_X1 U1043 ( .A1(G113), .A2(KEYINPUT58), .ZN(n1302) );
NAND2_X1 U1044 ( .A1(n1235), .A2(G214), .ZN(n1301) );
NOR2_X1 U1045 ( .A1(n1275), .A2(G237), .ZN(n1235) );
XOR2_X1 U1046 ( .A(n1303), .B(n1093), .Z(n1204) );
INV_X1 U1047 ( .A(G478), .ZN(n1093) );
NAND2_X1 U1048 ( .A1(n1091), .A2(n1214), .ZN(n1303) );
INV_X1 U1049 ( .A(G902), .ZN(n1214) );
XNOR2_X1 U1050 ( .A(n1304), .B(n1305), .ZN(n1091) );
XNOR2_X1 U1051 ( .A(n1000), .B(n1306), .ZN(n1305) );
XNOR2_X1 U1052 ( .A(G122), .B(n1261), .ZN(n1306) );
INV_X1 U1053 ( .A(G116), .ZN(n1261) );
INV_X1 U1054 ( .A(G107), .ZN(n1000) );
XOR2_X1 U1055 ( .A(n1307), .B(n1251), .Z(n1304) );
XOR2_X1 U1056 ( .A(G128), .B(n1291), .Z(n1251) );
XOR2_X1 U1057 ( .A(G143), .B(KEYINPUT13), .Z(n1291) );
XOR2_X1 U1058 ( .A(n1308), .B(n1309), .Z(n1307) );
NOR2_X1 U1059 ( .A1(KEYINPUT27), .A2(G134), .ZN(n1309) );
NAND2_X1 U1060 ( .A1(n1227), .A2(G217), .ZN(n1308) );
AND2_X1 U1061 ( .A1(G234), .A2(n1252), .ZN(n1227) );
INV_X1 U1062 ( .A(n1275), .ZN(n1252) );
XOR2_X1 U1063 ( .A(G953), .B(KEYINPUT33), .Z(n1275) );
endmodule


