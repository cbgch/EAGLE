//Key = 0010011000011101001001100010100111100111101011000111010100111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345;

XOR2_X1 U733 ( .A(n1029), .B(n1030), .Z(G9) );
NAND2_X1 U734 ( .A1(KEYINPUT58), .A2(G107), .ZN(n1030) );
NOR2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(G75) );
NOR3_X1 U736 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
NOR2_X1 U737 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR3_X1 U738 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1036) );
XOR2_X1 U739 ( .A(n1041), .B(KEYINPUT39), .Z(n1040) );
NAND4_X1 U740 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
NOR3_X1 U741 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1039) );
NOR2_X1 U742 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
AND2_X1 U743 ( .A1(n1043), .A2(n1051), .ZN(n1050) );
AND3_X1 U744 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1049) );
XOR2_X1 U745 ( .A(KEYINPUT7), .B(n1055), .Z(n1038) );
NOR4_X1 U746 ( .A1(n1056), .A2(n1054), .A3(n1057), .A4(n1048), .ZN(n1055) );
INV_X1 U747 ( .A(n1052), .ZN(n1057) );
NAND2_X1 U748 ( .A1(n1058), .A2(n1042), .ZN(n1056) );
NAND3_X1 U749 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1033) );
NAND4_X1 U750 ( .A1(n1042), .A2(n1043), .A3(n1052), .A4(n1062), .ZN(n1061) );
NAND3_X1 U751 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NAND2_X1 U752 ( .A1(n1045), .A2(n1066), .ZN(n1065) );
NAND3_X1 U753 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1064) );
XOR2_X1 U754 ( .A(KEYINPUT23), .B(n1045), .Z(n1068) );
NAND2_X1 U755 ( .A1(n1070), .A2(n1071), .ZN(n1063) );
NAND2_X1 U756 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
INV_X1 U757 ( .A(n1046), .ZN(n1042) );
NOR3_X1 U758 ( .A1(n1074), .A2(G953), .A3(G952), .ZN(n1031) );
INV_X1 U759 ( .A(n1059), .ZN(n1074) );
NAND4_X1 U760 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1059) );
NOR4_X1 U761 ( .A1(n1058), .A2(n1069), .A3(n1079), .A4(n1080), .ZN(n1078) );
XOR2_X1 U762 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U763 ( .A1(KEYINPUT33), .A2(n1083), .ZN(n1082) );
XOR2_X1 U764 ( .A(n1084), .B(n1085), .Z(n1079) );
NAND2_X1 U765 ( .A1(KEYINPUT40), .A2(n1086), .ZN(n1084) );
XNOR2_X1 U766 ( .A(KEYINPUT44), .B(n1087), .ZN(n1086) );
INV_X1 U767 ( .A(n1088), .ZN(n1069) );
NOR3_X1 U768 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1077) );
AND2_X1 U769 ( .A1(G469), .A2(n1092), .ZN(n1091) );
NOR2_X1 U770 ( .A1(G469), .A2(n1093), .ZN(n1090) );
NOR2_X1 U771 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR2_X1 U772 ( .A1(KEYINPUT25), .A2(n1092), .ZN(n1095) );
NOR2_X1 U773 ( .A1(n1096), .A2(KEYINPUT16), .ZN(n1092) );
INV_X1 U774 ( .A(n1097), .ZN(n1096) );
AND2_X1 U775 ( .A1(n1097), .A2(KEYINPUT25), .ZN(n1094) );
XOR2_X1 U776 ( .A(G478), .B(n1098), .Z(n1089) );
XOR2_X1 U777 ( .A(n1099), .B(n1100), .Z(n1076) );
NOR2_X1 U778 ( .A1(n1101), .A2(KEYINPUT36), .ZN(n1100) );
XOR2_X1 U779 ( .A(n1102), .B(KEYINPUT62), .Z(n1099) );
XOR2_X1 U780 ( .A(n1103), .B(KEYINPUT29), .Z(n1075) );
XOR2_X1 U781 ( .A(n1104), .B(n1105), .Z(G72) );
NOR2_X1 U782 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U783 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U784 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U785 ( .A1(KEYINPUT21), .A2(n1112), .ZN(n1110) );
XOR2_X1 U786 ( .A(G140), .B(G125), .Z(n1112) );
XOR2_X1 U787 ( .A(n1113), .B(n1114), .Z(n1108) );
XOR2_X1 U788 ( .A(G146), .B(G131), .Z(n1114) );
NOR2_X1 U789 ( .A1(KEYINPUT46), .A2(n1115), .ZN(n1113) );
XOR2_X1 U790 ( .A(G137), .B(G134), .Z(n1115) );
NAND3_X1 U791 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1104) );
INV_X1 U792 ( .A(n1106), .ZN(n1117) );
NAND2_X1 U793 ( .A1(G953), .A2(n1119), .ZN(n1116) );
XOR2_X1 U794 ( .A(n1120), .B(n1121), .Z(G69) );
XOR2_X1 U795 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U796 ( .A1(n1124), .A2(n1060), .ZN(n1123) );
AND2_X1 U797 ( .A1(G224), .A2(G898), .ZN(n1124) );
NAND2_X1 U798 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
INV_X1 U799 ( .A(n1127), .ZN(n1126) );
NAND2_X1 U800 ( .A1(n1060), .A2(n1128), .ZN(n1120) );
NAND2_X1 U801 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U802 ( .A1(n1131), .A2(n1132), .ZN(G66) );
NOR3_X1 U803 ( .A1(n1085), .A2(n1133), .A3(n1134), .ZN(n1132) );
NOR3_X1 U804 ( .A1(n1135), .A2(n1087), .A3(n1136), .ZN(n1134) );
NOR2_X1 U805 ( .A1(n1137), .A2(n1138), .ZN(n1133) );
NOR2_X1 U806 ( .A1(n1139), .A2(n1087), .ZN(n1138) );
NOR2_X1 U807 ( .A1(n1131), .A2(n1140), .ZN(G63) );
NOR3_X1 U808 ( .A1(n1098), .A2(n1141), .A3(n1142), .ZN(n1140) );
NOR3_X1 U809 ( .A1(n1143), .A2(n1144), .A3(n1136), .ZN(n1142) );
NOR2_X1 U810 ( .A1(n1145), .A2(n1146), .ZN(n1141) );
NOR2_X1 U811 ( .A1(n1139), .A2(n1144), .ZN(n1145) );
INV_X1 U812 ( .A(n1035), .ZN(n1139) );
NOR2_X1 U813 ( .A1(n1131), .A2(n1147), .ZN(G60) );
XOR2_X1 U814 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U815 ( .A1(n1150), .A2(n1136), .ZN(n1148) );
INV_X1 U816 ( .A(G475), .ZN(n1150) );
XNOR2_X1 U817 ( .A(G104), .B(n1130), .ZN(G6) );
NOR2_X1 U818 ( .A1(n1151), .A2(n1152), .ZN(G57) );
XOR2_X1 U819 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U820 ( .A(n1155), .B(n1156), .Z(n1154) );
NAND2_X1 U821 ( .A1(KEYINPUT60), .A2(n1157), .ZN(n1155) );
XOR2_X1 U822 ( .A(n1158), .B(n1159), .Z(n1153) );
NOR2_X1 U823 ( .A1(n1160), .A2(KEYINPUT35), .ZN(n1159) );
NOR2_X1 U824 ( .A1(n1102), .A2(n1136), .ZN(n1160) );
INV_X1 U825 ( .A(G472), .ZN(n1102) );
XOR2_X1 U826 ( .A(n1161), .B(KEYINPUT48), .Z(n1151) );
NAND2_X1 U827 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U828 ( .A1(n1131), .A2(n1164), .ZN(n1163) );
INV_X1 U829 ( .A(KEYINPUT63), .ZN(n1164) );
NAND3_X1 U830 ( .A1(G952), .A2(G953), .A3(KEYINPUT63), .ZN(n1162) );
NOR2_X1 U831 ( .A1(n1131), .A2(n1165), .ZN(G54) );
XOR2_X1 U832 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U833 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U834 ( .A1(KEYINPUT28), .A2(n1170), .ZN(n1169) );
NAND2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
NAND2_X1 U836 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U837 ( .A(KEYINPUT18), .B(n1175), .Z(n1171) );
NOR2_X1 U838 ( .A1(n1176), .A2(n1174), .ZN(n1175) );
XNOR2_X1 U839 ( .A(n1173), .B(KEYINPUT32), .ZN(n1176) );
XNOR2_X1 U840 ( .A(n1177), .B(G146), .ZN(n1173) );
XOR2_X1 U841 ( .A(n1178), .B(n1179), .Z(n1166) );
NOR2_X1 U842 ( .A1(n1180), .A2(n1136), .ZN(n1179) );
XNOR2_X1 U843 ( .A(G110), .B(n1181), .ZN(n1178) );
NOR2_X1 U844 ( .A1(KEYINPUT0), .A2(n1182), .ZN(n1181) );
NOR2_X1 U845 ( .A1(n1131), .A2(n1183), .ZN(G51) );
XOR2_X1 U846 ( .A(n1184), .B(n1125), .Z(n1183) );
XOR2_X1 U847 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U848 ( .A1(n1187), .A2(n1136), .ZN(n1186) );
NAND2_X1 U849 ( .A1(G902), .A2(n1035), .ZN(n1136) );
NAND3_X1 U850 ( .A1(n1118), .A2(n1129), .A3(n1188), .ZN(n1035) );
XOR2_X1 U851 ( .A(n1130), .B(KEYINPUT8), .Z(n1188) );
NAND3_X1 U852 ( .A1(n1189), .A2(n1052), .A3(n1190), .ZN(n1130) );
AND4_X1 U853 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1129) );
AND4_X1 U854 ( .A1(n1029), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1194) );
NAND3_X1 U855 ( .A1(n1198), .A2(n1052), .A3(n1189), .ZN(n1029) );
AND4_X1 U856 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1118) );
AND4_X1 U857 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
NOR2_X1 U858 ( .A1(n1207), .A2(n1208), .ZN(n1201) );
NOR3_X1 U859 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
XOR2_X1 U860 ( .A(n1073), .B(KEYINPUT61), .Z(n1210) );
NAND2_X1 U861 ( .A1(n1212), .A2(n1213), .ZN(n1185) );
NAND2_X1 U862 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U863 ( .A(n1216), .B(n1217), .Z(n1214) );
XOR2_X1 U864 ( .A(n1218), .B(KEYINPUT54), .Z(n1212) );
NAND2_X1 U865 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
XNOR2_X1 U866 ( .A(n1217), .B(n1216), .ZN(n1219) );
NOR2_X1 U867 ( .A1(G125), .A2(KEYINPUT27), .ZN(n1216) );
NOR2_X1 U868 ( .A1(n1060), .A2(G952), .ZN(n1131) );
XNOR2_X1 U869 ( .A(n1207), .B(n1221), .ZN(G48) );
NAND2_X1 U870 ( .A1(KEYINPUT53), .A2(G146), .ZN(n1221) );
NOR3_X1 U871 ( .A1(n1209), .A2(n1211), .A3(n1072), .ZN(n1207) );
INV_X1 U872 ( .A(n1190), .ZN(n1072) );
XNOR2_X1 U873 ( .A(G143), .B(n1199), .ZN(G45) );
NAND4_X1 U874 ( .A1(n1222), .A2(n1066), .A3(n1223), .A4(n1224), .ZN(n1199) );
XOR2_X1 U875 ( .A(n1170), .B(n1200), .Z(G42) );
NAND4_X1 U876 ( .A1(n1190), .A2(n1044), .A3(n1070), .A4(n1225), .ZN(n1200) );
XNOR2_X1 U877 ( .A(G137), .B(n1203), .ZN(G39) );
OR3_X1 U878 ( .A1(n1037), .A2(n1209), .A3(n1048), .ZN(n1203) );
INV_X1 U879 ( .A(n1045), .ZN(n1048) );
XOR2_X1 U880 ( .A(n1226), .B(n1206), .Z(G36) );
NAND3_X1 U881 ( .A1(n1070), .A2(n1198), .A3(n1222), .ZN(n1206) );
NAND2_X1 U882 ( .A1(n1227), .A2(n1228), .ZN(G33) );
NAND2_X1 U883 ( .A1(G131), .A2(n1205), .ZN(n1228) );
XOR2_X1 U884 ( .A(n1229), .B(KEYINPUT3), .Z(n1227) );
OR2_X1 U885 ( .A1(n1205), .A2(G131), .ZN(n1229) );
NAND3_X1 U886 ( .A1(n1190), .A2(n1070), .A3(n1222), .ZN(n1205) );
AND2_X1 U887 ( .A1(n1051), .A2(n1225), .ZN(n1222) );
INV_X1 U888 ( .A(n1037), .ZN(n1070) );
NAND2_X1 U889 ( .A1(n1230), .A2(n1088), .ZN(n1037) );
XOR2_X1 U890 ( .A(n1067), .B(KEYINPUT43), .Z(n1230) );
XOR2_X1 U891 ( .A(G128), .B(n1231), .Z(G30) );
NOR3_X1 U892 ( .A1(n1209), .A2(n1232), .A3(n1073), .ZN(n1231) );
XOR2_X1 U893 ( .A(n1211), .B(KEYINPUT9), .Z(n1232) );
NAND3_X1 U894 ( .A1(n1233), .A2(n1234), .A3(n1225), .ZN(n1209) );
AND3_X1 U895 ( .A1(n1235), .A2(n1053), .A3(n1054), .ZN(n1225) );
XOR2_X1 U896 ( .A(n1157), .B(n1193), .Z(G3) );
NAND3_X1 U897 ( .A1(n1045), .A2(n1189), .A3(n1051), .ZN(n1193) );
XNOR2_X1 U898 ( .A(G125), .B(n1204), .ZN(G27) );
NAND4_X1 U899 ( .A1(n1190), .A2(n1043), .A3(n1236), .A4(n1044), .ZN(n1204) );
AND2_X1 U900 ( .A1(n1235), .A2(n1066), .ZN(n1236) );
NAND2_X1 U901 ( .A1(n1046), .A2(n1237), .ZN(n1235) );
NAND3_X1 U902 ( .A1(G902), .A2(n1238), .A3(n1106), .ZN(n1237) );
NOR2_X1 U903 ( .A1(G900), .A2(n1060), .ZN(n1106) );
XOR2_X1 U904 ( .A(n1191), .B(n1239), .Z(G24) );
NAND2_X1 U905 ( .A1(KEYINPUT6), .A2(G122), .ZN(n1239) );
NAND4_X1 U906 ( .A1(n1240), .A2(n1052), .A3(n1223), .A4(n1224), .ZN(n1191) );
NOR2_X1 U907 ( .A1(n1234), .A2(n1233), .ZN(n1052) );
XOR2_X1 U908 ( .A(n1241), .B(G119), .Z(G21) );
NAND2_X1 U909 ( .A1(KEYINPUT5), .A2(n1192), .ZN(n1241) );
NAND4_X1 U910 ( .A1(n1240), .A2(n1045), .A3(n1233), .A4(n1234), .ZN(n1192) );
XOR2_X1 U911 ( .A(G116), .B(n1242), .Z(G18) );
NOR2_X1 U912 ( .A1(KEYINPUT10), .A2(n1197), .ZN(n1242) );
NAND3_X1 U913 ( .A1(n1051), .A2(n1198), .A3(n1240), .ZN(n1197) );
INV_X1 U914 ( .A(n1073), .ZN(n1198) );
NAND2_X1 U915 ( .A1(n1243), .A2(n1224), .ZN(n1073) );
XNOR2_X1 U916 ( .A(G113), .B(n1196), .ZN(G15) );
NAND3_X1 U917 ( .A1(n1051), .A2(n1190), .A3(n1240), .ZN(n1196) );
AND2_X1 U918 ( .A1(n1043), .A2(n1244), .ZN(n1240) );
NOR2_X1 U919 ( .A1(n1054), .A2(n1058), .ZN(n1043) );
INV_X1 U920 ( .A(n1053), .ZN(n1058) );
NOR2_X1 U921 ( .A1(n1224), .A2(n1243), .ZN(n1190) );
NOR2_X1 U922 ( .A1(n1233), .A2(n1245), .ZN(n1051) );
XNOR2_X1 U923 ( .A(G110), .B(n1195), .ZN(G12) );
NAND3_X1 U924 ( .A1(n1045), .A2(n1189), .A3(n1044), .ZN(n1195) );
AND2_X1 U925 ( .A1(n1245), .A2(n1233), .ZN(n1044) );
XNOR2_X1 U926 ( .A(n1085), .B(n1087), .ZN(n1233) );
NAND2_X1 U927 ( .A1(G217), .A2(n1246), .ZN(n1087) );
NOR2_X1 U928 ( .A1(n1137), .A2(G902), .ZN(n1085) );
INV_X1 U929 ( .A(n1135), .ZN(n1137) );
NAND2_X1 U930 ( .A1(n1247), .A2(n1248), .ZN(n1135) );
NAND2_X1 U931 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
XOR2_X1 U932 ( .A(KEYINPUT38), .B(n1251), .Z(n1247) );
NOR2_X1 U933 ( .A1(n1250), .A2(n1249), .ZN(n1251) );
XOR2_X1 U934 ( .A(n1252), .B(n1253), .Z(n1249) );
XOR2_X1 U935 ( .A(n1254), .B(n1255), .Z(n1253) );
NAND2_X1 U936 ( .A1(KEYINPUT2), .A2(n1256), .ZN(n1252) );
XOR2_X1 U937 ( .A(G125), .B(n1257), .Z(n1256) );
XOR2_X1 U938 ( .A(G137), .B(n1258), .Z(n1250) );
NOR2_X1 U939 ( .A1(n1259), .A2(KEYINPUT47), .ZN(n1258) );
AND3_X1 U940 ( .A1(G221), .A2(n1060), .A3(G234), .ZN(n1259) );
INV_X1 U941 ( .A(n1234), .ZN(n1245) );
XOR2_X1 U942 ( .A(n1101), .B(G472), .Z(n1234) );
AND2_X1 U943 ( .A1(n1260), .A2(n1261), .ZN(n1101) );
XOR2_X1 U944 ( .A(n1262), .B(n1263), .Z(n1260) );
NOR2_X1 U945 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NOR2_X1 U946 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
INV_X1 U947 ( .A(n1158), .ZN(n1267) );
NOR2_X1 U948 ( .A1(n1268), .A2(n1269), .ZN(n1266) );
NOR2_X1 U949 ( .A1(n1270), .A2(n1271), .ZN(n1264) );
XOR2_X1 U950 ( .A(n1157), .B(KEYINPUT59), .Z(n1271) );
NOR2_X1 U951 ( .A1(n1272), .A2(n1268), .ZN(n1270) );
XOR2_X1 U952 ( .A(n1157), .B(KEYINPUT12), .Z(n1268) );
INV_X1 U953 ( .A(G101), .ZN(n1157) );
NOR2_X1 U954 ( .A1(n1158), .A2(n1269), .ZN(n1272) );
INV_X1 U955 ( .A(KEYINPUT34), .ZN(n1269) );
NAND2_X1 U956 ( .A1(n1273), .A2(G210), .ZN(n1158) );
NAND2_X1 U957 ( .A1(n1274), .A2(KEYINPUT45), .ZN(n1262) );
XNOR2_X1 U958 ( .A(n1156), .B(n1275), .ZN(n1274) );
XOR2_X1 U959 ( .A(KEYINPUT14), .B(KEYINPUT1), .Z(n1275) );
XNOR2_X1 U960 ( .A(n1276), .B(n1277), .ZN(n1156) );
XOR2_X1 U961 ( .A(n1278), .B(n1279), .Z(n1277) );
XNOR2_X1 U962 ( .A(G113), .B(KEYINPUT37), .ZN(n1279) );
NAND2_X1 U963 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
NAND2_X1 U964 ( .A1(G116), .A2(n1282), .ZN(n1281) );
XOR2_X1 U965 ( .A(n1283), .B(KEYINPUT4), .Z(n1280) );
OR2_X1 U966 ( .A1(n1282), .A2(G116), .ZN(n1283) );
INV_X1 U967 ( .A(G119), .ZN(n1282) );
XNOR2_X1 U968 ( .A(n1217), .B(n1174), .ZN(n1276) );
AND3_X1 U969 ( .A1(n1054), .A2(n1053), .A3(n1244), .ZN(n1189) );
AND2_X1 U970 ( .A1(n1066), .A2(n1284), .ZN(n1244) );
NAND2_X1 U971 ( .A1(n1046), .A2(n1285), .ZN(n1284) );
NAND3_X1 U972 ( .A1(n1127), .A2(n1286), .A3(G902), .ZN(n1285) );
XNOR2_X1 U973 ( .A(KEYINPUT49), .B(n1238), .ZN(n1286) );
NOR2_X1 U974 ( .A1(n1060), .A2(G898), .ZN(n1127) );
NAND3_X1 U975 ( .A1(n1238), .A2(n1060), .A3(G952), .ZN(n1046) );
NAND2_X1 U976 ( .A1(G237), .A2(G234), .ZN(n1238) );
INV_X1 U977 ( .A(n1211), .ZN(n1066) );
NAND2_X1 U978 ( .A1(n1287), .A2(n1088), .ZN(n1211) );
NAND2_X1 U979 ( .A1(G214), .A2(n1288), .ZN(n1088) );
INV_X1 U980 ( .A(n1067), .ZN(n1287) );
XOR2_X1 U981 ( .A(n1081), .B(n1083), .Z(n1067) );
INV_X1 U982 ( .A(n1187), .ZN(n1083) );
NAND2_X1 U983 ( .A1(G210), .A2(n1288), .ZN(n1187) );
NAND2_X1 U984 ( .A1(n1289), .A2(n1261), .ZN(n1288) );
INV_X1 U985 ( .A(G237), .ZN(n1289) );
NAND2_X1 U986 ( .A1(n1290), .A2(n1261), .ZN(n1081) );
XOR2_X1 U987 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U988 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U989 ( .A(G125), .B(KEYINPUT26), .ZN(n1294) );
NAND2_X1 U990 ( .A1(KEYINPUT11), .A2(n1220), .ZN(n1293) );
INV_X1 U991 ( .A(n1215), .ZN(n1220) );
NAND2_X1 U992 ( .A1(G224), .A2(n1060), .ZN(n1215) );
XNOR2_X1 U993 ( .A(n1217), .B(n1125), .ZN(n1291) );
XNOR2_X1 U994 ( .A(n1295), .B(n1296), .ZN(n1125) );
XOR2_X1 U995 ( .A(n1255), .B(n1297), .Z(n1296) );
XOR2_X1 U996 ( .A(KEYINPUT31), .B(G101), .Z(n1297) );
XOR2_X1 U997 ( .A(G110), .B(G119), .Z(n1255) );
XOR2_X1 U998 ( .A(n1298), .B(n1299), .Z(n1295) );
XNOR2_X1 U999 ( .A(n1300), .B(G128), .ZN(n1217) );
NAND2_X1 U1000 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1001 ( .A1(G146), .A2(n1303), .ZN(n1302) );
XOR2_X1 U1002 ( .A(KEYINPUT55), .B(n1304), .Z(n1301) );
NOR2_X1 U1003 ( .A1(G146), .A2(n1303), .ZN(n1304) );
XOR2_X1 U1004 ( .A(KEYINPUT57), .B(n1305), .Z(n1303) );
NAND2_X1 U1005 ( .A1(G221), .A2(n1246), .ZN(n1053) );
NAND2_X1 U1006 ( .A1(G234), .A2(n1261), .ZN(n1246) );
XOR2_X1 U1007 ( .A(n1097), .B(n1180), .Z(n1054) );
INV_X1 U1008 ( .A(G469), .ZN(n1180) );
NAND2_X1 U1009 ( .A1(n1306), .A2(n1261), .ZN(n1097) );
INV_X1 U1010 ( .A(G902), .ZN(n1261) );
XOR2_X1 U1011 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1012 ( .A(n1177), .B(n1309), .Z(n1308) );
XOR2_X1 U1013 ( .A(n1310), .B(n1174), .Z(n1309) );
XNOR2_X1 U1014 ( .A(n1311), .B(n1312), .ZN(n1174) );
XOR2_X1 U1015 ( .A(G131), .B(n1313), .Z(n1312) );
NOR2_X1 U1016 ( .A1(G137), .A2(KEYINPUT30), .ZN(n1313) );
XOR2_X1 U1017 ( .A(n1226), .B(KEYINPUT15), .Z(n1311) );
INV_X1 U1018 ( .A(G134), .ZN(n1226) );
XOR2_X1 U1019 ( .A(n1314), .B(n1315), .Z(n1177) );
XOR2_X1 U1020 ( .A(KEYINPUT51), .B(G101), .Z(n1315) );
XOR2_X1 U1021 ( .A(n1111), .B(n1316), .Z(n1314) );
NOR2_X1 U1022 ( .A1(KEYINPUT56), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1023 ( .A(G104), .B(G107), .ZN(n1317) );
XOR2_X1 U1024 ( .A(n1254), .B(n1305), .Z(n1111) );
XOR2_X1 U1025 ( .A(G143), .B(KEYINPUT13), .Z(n1305) );
INV_X1 U1026 ( .A(G128), .ZN(n1254) );
XOR2_X1 U1027 ( .A(n1182), .B(n1318), .Z(n1307) );
XOR2_X1 U1028 ( .A(KEYINPUT24), .B(G110), .Z(n1318) );
NOR2_X1 U1029 ( .A1(n1119), .A2(G953), .ZN(n1182) );
INV_X1 U1030 ( .A(G227), .ZN(n1119) );
NOR2_X1 U1031 ( .A1(n1224), .A2(n1223), .ZN(n1045) );
INV_X1 U1032 ( .A(n1243), .ZN(n1223) );
XOR2_X1 U1033 ( .A(n1103), .B(KEYINPUT17), .Z(n1243) );
XOR2_X1 U1034 ( .A(n1319), .B(G475), .Z(n1103) );
OR2_X1 U1035 ( .A1(n1149), .A2(G902), .ZN(n1319) );
XNOR2_X1 U1036 ( .A(n1298), .B(n1320), .ZN(n1149) );
NOR2_X1 U1037 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
NOR2_X1 U1038 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NOR2_X1 U1039 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
INV_X1 U1040 ( .A(KEYINPUT42), .ZN(n1326) );
AND2_X1 U1041 ( .A1(n1327), .A2(KEYINPUT50), .ZN(n1325) );
NOR2_X1 U1042 ( .A1(n1328), .A2(n1327), .ZN(n1321) );
XNOR2_X1 U1043 ( .A(n1329), .B(n1330), .ZN(n1327) );
XOR2_X1 U1044 ( .A(G143), .B(G131), .Z(n1330) );
NAND2_X1 U1045 ( .A1(n1273), .A2(G214), .ZN(n1329) );
NOR2_X1 U1046 ( .A1(G953), .A2(G237), .ZN(n1273) );
NOR2_X1 U1047 ( .A1(n1331), .A2(n1332), .ZN(n1328) );
INV_X1 U1048 ( .A(KEYINPUT50), .ZN(n1332) );
AND2_X1 U1049 ( .A1(n1324), .A2(KEYINPUT42), .ZN(n1331) );
XNOR2_X1 U1050 ( .A(n1333), .B(n1257), .ZN(n1324) );
INV_X1 U1051 ( .A(n1310), .ZN(n1257) );
XOR2_X1 U1052 ( .A(n1170), .B(G146), .Z(n1310) );
INV_X1 U1053 ( .A(G140), .ZN(n1170) );
NAND2_X1 U1054 ( .A1(KEYINPUT22), .A2(G125), .ZN(n1333) );
XNOR2_X1 U1055 ( .A(G104), .B(n1334), .ZN(n1298) );
XOR2_X1 U1056 ( .A(G122), .B(G113), .Z(n1334) );
NAND2_X1 U1057 ( .A1(n1335), .A2(n1336), .ZN(n1224) );
NAND2_X1 U1058 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1059 ( .A(KEYINPUT41), .B(G478), .Z(n1338) );
XNOR2_X1 U1060 ( .A(n1098), .B(KEYINPUT52), .ZN(n1337) );
XOR2_X1 U1061 ( .A(n1339), .B(KEYINPUT19), .Z(n1335) );
NAND2_X1 U1062 ( .A1(n1098), .A2(n1144), .ZN(n1339) );
INV_X1 U1063 ( .A(G478), .ZN(n1144) );
NOR2_X1 U1064 ( .A1(n1146), .A2(G902), .ZN(n1098) );
INV_X1 U1065 ( .A(n1143), .ZN(n1146) );
XOR2_X1 U1066 ( .A(n1340), .B(n1341), .Z(n1143) );
XOR2_X1 U1067 ( .A(G122), .B(n1342), .Z(n1341) );
XOR2_X1 U1068 ( .A(G143), .B(G134), .Z(n1342) );
XOR2_X1 U1069 ( .A(n1343), .B(n1299), .Z(n1340) );
XOR2_X1 U1070 ( .A(G107), .B(G116), .Z(n1299) );
XOR2_X1 U1071 ( .A(n1344), .B(n1345), .Z(n1343) );
NOR2_X1 U1072 ( .A1(G128), .A2(KEYINPUT20), .ZN(n1345) );
NAND3_X1 U1073 ( .A1(G234), .A2(n1060), .A3(G217), .ZN(n1344) );
INV_X1 U1074 ( .A(G953), .ZN(n1060) );
endmodule


