//Key = 0101110100100110111110001101100101000111110001111110111000001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369;

NAND2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(G9) );
OR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
XOR2_X1 U756 ( .A(n1053), .B(KEYINPUT35), .Z(n1049) );
NAND2_X1 U757 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
NOR3_X1 U758 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1052) );
NOR2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(G75) );
NOR4_X1 U760 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U763 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
INV_X1 U764 ( .A(n1069), .ZN(n1068) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1067) );
NOR3_X1 U766 ( .A1(n1072), .A2(n1073), .A3(n1054), .ZN(n1065) );
NOR2_X1 U767 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR2_X1 U770 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1074) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
XOR2_X1 U774 ( .A(KEYINPUT39), .B(n1088), .Z(n1087) );
NAND3_X1 U775 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1059) );
NAND3_X1 U776 ( .A1(n1092), .A2(n1093), .A3(n1069), .ZN(n1091) );
NOR3_X1 U777 ( .A1(n1077), .A2(n1083), .A3(n1072), .ZN(n1069) );
INV_X1 U778 ( .A(n1094), .ZN(n1077) );
NAND2_X1 U779 ( .A1(n1095), .A2(n1055), .ZN(n1093) );
NOR3_X1 U780 ( .A1(n1096), .A2(G953), .A3(G952), .ZN(n1057) );
INV_X1 U781 ( .A(n1089), .ZN(n1096) );
NAND4_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1089) );
NOR4_X1 U783 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
XOR2_X1 U784 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U785 ( .A(KEYINPUT34), .B(n1107), .ZN(n1103) );
XOR2_X1 U786 ( .A(n1108), .B(n1109), .Z(n1102) );
XOR2_X1 U787 ( .A(n1110), .B(G469), .Z(n1109) );
XNOR2_X1 U788 ( .A(KEYINPUT47), .B(KEYINPUT40), .ZN(n1108) );
NOR3_X1 U789 ( .A1(n1111), .A2(n1112), .A3(n1088), .ZN(n1099) );
NAND2_X1 U790 ( .A1(G478), .A2(n1113), .ZN(n1098) );
XNOR2_X1 U791 ( .A(KEYINPUT5), .B(n1114), .ZN(n1113) );
XOR2_X1 U792 ( .A(n1115), .B(n1116), .Z(G72) );
NOR2_X1 U793 ( .A1(n1117), .A2(n1090), .ZN(n1116) );
AND2_X1 U794 ( .A1(G227), .A2(G900), .ZN(n1117) );
NAND2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1115) );
NAND2_X1 U796 ( .A1(n1120), .A2(n1090), .ZN(n1119) );
XOR2_X1 U797 ( .A(n1121), .B(n1060), .Z(n1120) );
NAND3_X1 U798 ( .A1(G900), .A2(n1121), .A3(G953), .ZN(n1118) );
XNOR2_X1 U799 ( .A(n1122), .B(n1123), .ZN(n1121) );
XOR2_X1 U800 ( .A(n1124), .B(n1125), .Z(n1123) );
XNOR2_X1 U801 ( .A(n1126), .B(n1127), .ZN(n1122) );
NAND2_X1 U802 ( .A1(KEYINPUT45), .A2(n1128), .ZN(n1126) );
XOR2_X1 U803 ( .A(n1129), .B(n1130), .Z(G69) );
XOR2_X1 U804 ( .A(n1131), .B(n1132), .Z(n1130) );
AND2_X1 U805 ( .A1(n1062), .A2(n1090), .ZN(n1132) );
NOR2_X1 U806 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
XOR2_X1 U807 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U808 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U809 ( .A1(KEYINPUT52), .A2(n1139), .ZN(n1137) );
XOR2_X1 U810 ( .A(n1140), .B(KEYINPUT61), .Z(n1135) );
NOR2_X1 U811 ( .A1(G898), .A2(n1090), .ZN(n1133) );
NOR2_X1 U812 ( .A1(n1141), .A2(n1090), .ZN(n1129) );
AND2_X1 U813 ( .A1(G224), .A2(G898), .ZN(n1141) );
NOR2_X1 U814 ( .A1(n1142), .A2(n1143), .ZN(G66) );
XNOR2_X1 U815 ( .A(n1144), .B(n1145), .ZN(n1143) );
NAND3_X1 U816 ( .A1(n1146), .A2(G217), .A3(KEYINPUT48), .ZN(n1144) );
NOR3_X1 U817 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(G63) );
AND2_X1 U818 ( .A1(KEYINPUT18), .A2(n1142), .ZN(n1149) );
NOR3_X1 U819 ( .A1(KEYINPUT18), .A2(G953), .A3(G952), .ZN(n1148) );
XOR2_X1 U820 ( .A(n1150), .B(n1151), .Z(n1147) );
AND2_X1 U821 ( .A1(G478), .A2(n1146), .ZN(n1151) );
NAND2_X1 U822 ( .A1(KEYINPUT7), .A2(n1152), .ZN(n1150) );
NOR2_X1 U823 ( .A1(n1142), .A2(n1153), .ZN(G60) );
XNOR2_X1 U824 ( .A(n1154), .B(n1155), .ZN(n1153) );
AND2_X1 U825 ( .A1(G475), .A2(n1146), .ZN(n1155) );
XNOR2_X1 U826 ( .A(G104), .B(n1156), .ZN(G6) );
NOR2_X1 U827 ( .A1(n1142), .A2(n1157), .ZN(G57) );
XNOR2_X1 U828 ( .A(n1158), .B(n1159), .ZN(n1157) );
NAND2_X1 U829 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND2_X1 U830 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U831 ( .A1(KEYINPUT62), .A2(n1164), .ZN(n1162) );
NAND2_X1 U832 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NAND2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1160) );
NAND2_X1 U834 ( .A1(n1166), .A2(n1169), .ZN(n1168) );
NAND2_X1 U835 ( .A1(n1170), .A2(KEYINPUT62), .ZN(n1169) );
INV_X1 U836 ( .A(n1163), .ZN(n1170) );
NAND2_X1 U837 ( .A1(n1146), .A2(G472), .ZN(n1163) );
INV_X1 U838 ( .A(KEYINPUT21), .ZN(n1166) );
NOR2_X1 U839 ( .A1(n1142), .A2(n1171), .ZN(G54) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U842 ( .A(n1176), .B(n1177), .Z(n1175) );
AND2_X1 U843 ( .A1(G469), .A2(n1146), .ZN(n1176) );
INV_X1 U844 ( .A(n1178), .ZN(n1146) );
XOR2_X1 U845 ( .A(n1179), .B(n1180), .Z(n1172) );
XOR2_X1 U846 ( .A(KEYINPUT41), .B(n1181), .Z(n1180) );
NOR2_X1 U847 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XOR2_X1 U848 ( .A(KEYINPUT63), .B(n1184), .Z(n1183) );
AND2_X1 U849 ( .A1(n1125), .A2(n1185), .ZN(n1184) );
NOR2_X1 U850 ( .A1(n1125), .A2(n1185), .ZN(n1182) );
XOR2_X1 U851 ( .A(n1139), .B(KEYINPUT20), .Z(n1185) );
NOR2_X1 U852 ( .A1(n1186), .A2(KEYINPUT56), .ZN(n1179) );
INV_X1 U853 ( .A(n1187), .ZN(n1186) );
NOR2_X1 U854 ( .A1(n1142), .A2(n1188), .ZN(G51) );
XOR2_X1 U855 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U856 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U857 ( .A(KEYINPUT55), .B(n1193), .Z(n1192) );
AND2_X1 U858 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U859 ( .A1(n1195), .A2(n1194), .ZN(n1191) );
NAND2_X1 U860 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
NAND2_X1 U861 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XOR2_X1 U862 ( .A(n1200), .B(KEYINPUT30), .Z(n1196) );
OR2_X1 U863 ( .A1(n1199), .A2(n1198), .ZN(n1200) );
XOR2_X1 U864 ( .A(n1201), .B(G125), .Z(n1198) );
NAND2_X1 U865 ( .A1(KEYINPUT33), .A2(n1202), .ZN(n1201) );
NOR2_X1 U866 ( .A1(n1105), .A2(n1178), .ZN(n1189) );
NAND2_X1 U867 ( .A1(G902), .A2(n1203), .ZN(n1178) );
OR2_X1 U868 ( .A1(n1060), .A2(n1062), .ZN(n1203) );
NAND4_X1 U869 ( .A1(n1204), .A2(n1156), .A3(n1205), .A4(n1206), .ZN(n1062) );
AND4_X1 U870 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
NAND2_X1 U871 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
NAND2_X1 U872 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND3_X1 U873 ( .A1(n1215), .A2(n1216), .A3(n1092), .ZN(n1214) );
NAND2_X1 U874 ( .A1(KEYINPUT50), .A2(n1056), .ZN(n1216) );
NAND2_X1 U875 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
INV_X1 U876 ( .A(KEYINPUT50), .ZN(n1218) );
NAND2_X1 U877 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
NAND2_X1 U878 ( .A1(n1221), .A2(n1071), .ZN(n1213) );
NAND3_X1 U879 ( .A1(n1222), .A2(n1092), .A3(n1223), .ZN(n1156) );
NAND3_X1 U880 ( .A1(n1224), .A2(n1092), .A3(n1221), .ZN(n1204) );
NAND2_X1 U881 ( .A1(n1225), .A2(n1226), .ZN(n1060) );
NOR4_X1 U882 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1226) );
NOR4_X1 U883 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1225) );
NOR3_X1 U884 ( .A1(n1235), .A2(n1236), .A3(n1064), .ZN(n1233) );
XOR2_X1 U885 ( .A(KEYINPUT53), .B(n1237), .Z(n1235) );
NOR4_X1 U886 ( .A1(n1238), .A2(n1239), .A3(n1055), .A4(n1240), .ZN(n1232) );
NOR2_X1 U887 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
INV_X1 U888 ( .A(KEYINPUT15), .ZN(n1242) );
NOR2_X1 U889 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
NOR2_X1 U890 ( .A1(KEYINPUT15), .A2(n1245), .ZN(n1238) );
NOR2_X1 U891 ( .A1(n1090), .A2(G952), .ZN(n1142) );
XNOR2_X1 U892 ( .A(G146), .B(n1246), .ZN(G48) );
NOR2_X1 U893 ( .A1(n1231), .A2(KEYINPUT0), .ZN(n1246) );
AND2_X1 U894 ( .A1(n1223), .A2(n1247), .ZN(n1231) );
XOR2_X1 U895 ( .A(G143), .B(n1230), .Z(G45) );
AND4_X1 U896 ( .A1(n1224), .A2(n1071), .A3(n1248), .A4(n1079), .ZN(n1230) );
XOR2_X1 U897 ( .A(G140), .B(n1229), .Z(G42) );
AND3_X1 U898 ( .A1(n1223), .A2(n1245), .A3(n1070), .ZN(n1229) );
XNOR2_X1 U899 ( .A(G137), .B(n1249), .ZN(G39) );
NAND3_X1 U900 ( .A1(n1245), .A2(n1237), .A3(n1250), .ZN(n1249) );
XOR2_X1 U901 ( .A(n1251), .B(n1252), .Z(G36) );
NOR2_X1 U902 ( .A1(KEYINPUT8), .A2(n1253), .ZN(n1252) );
XNOR2_X1 U903 ( .A(G134), .B(KEYINPUT37), .ZN(n1253) );
NAND3_X1 U904 ( .A1(n1245), .A2(n1211), .A3(n1071), .ZN(n1251) );
XOR2_X1 U905 ( .A(n1228), .B(n1254), .Z(G33) );
NOR2_X1 U906 ( .A1(KEYINPUT43), .A2(n1127), .ZN(n1254) );
NOR3_X1 U907 ( .A1(n1240), .A2(n1236), .A3(n1095), .ZN(n1228) );
INV_X1 U908 ( .A(n1245), .ZN(n1236) );
NOR2_X1 U909 ( .A1(n1083), .A2(n1244), .ZN(n1245) );
INV_X1 U910 ( .A(n1243), .ZN(n1083) );
NOR2_X1 U911 ( .A1(n1080), .A2(n1111), .ZN(n1243) );
INV_X1 U912 ( .A(n1081), .ZN(n1111) );
XNOR2_X1 U913 ( .A(G128), .B(n1255), .ZN(G30) );
NAND2_X1 U914 ( .A1(KEYINPUT24), .A2(n1227), .ZN(n1255) );
AND2_X1 U915 ( .A1(n1247), .A2(n1211), .ZN(n1227) );
INV_X1 U916 ( .A(n1055), .ZN(n1211) );
AND3_X1 U917 ( .A1(n1248), .A2(n1079), .A3(n1237), .ZN(n1247) );
INV_X1 U918 ( .A(n1244), .ZN(n1248) );
NAND2_X1 U919 ( .A1(n1085), .A2(n1256), .ZN(n1244) );
XNOR2_X1 U920 ( .A(G101), .B(n1210), .ZN(G3) );
NAND3_X1 U921 ( .A1(n1071), .A2(n1222), .A3(n1250), .ZN(n1210) );
XNOR2_X1 U922 ( .A(n1257), .B(n1258), .ZN(G27) );
NAND2_X1 U923 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND3_X1 U924 ( .A1(n1079), .A2(n1261), .A3(n1262), .ZN(n1260) );
INV_X1 U925 ( .A(KEYINPUT49), .ZN(n1262) );
NAND2_X1 U926 ( .A1(n1234), .A2(KEYINPUT49), .ZN(n1259) );
NOR2_X1 U927 ( .A1(n1261), .A2(n1263), .ZN(n1234) );
INV_X1 U928 ( .A(n1079), .ZN(n1263) );
NAND4_X1 U929 ( .A1(n1094), .A2(n1070), .A3(n1223), .A4(n1256), .ZN(n1261) );
NAND2_X1 U930 ( .A1(n1264), .A2(n1072), .ZN(n1256) );
NAND4_X1 U931 ( .A1(G902), .A2(G953), .A3(n1265), .A4(n1266), .ZN(n1264) );
INV_X1 U932 ( .A(G900), .ZN(n1266) );
XOR2_X1 U933 ( .A(n1267), .B(n1268), .Z(G24) );
XNOR2_X1 U934 ( .A(G122), .B(KEYINPUT2), .ZN(n1268) );
NAND3_X1 U935 ( .A1(n1092), .A2(n1269), .A3(n1221), .ZN(n1267) );
XOR2_X1 U936 ( .A(KEYINPUT26), .B(n1224), .Z(n1269) );
AND2_X1 U937 ( .A1(n1101), .A2(n1270), .ZN(n1224) );
INV_X1 U938 ( .A(n1054), .ZN(n1092) );
NAND2_X1 U939 ( .A1(n1097), .A2(n1107), .ZN(n1054) );
XOR2_X1 U940 ( .A(n1208), .B(n1271), .Z(G21) );
NAND2_X1 U941 ( .A1(KEYINPUT14), .A2(G119), .ZN(n1271) );
NAND3_X1 U942 ( .A1(n1250), .A2(n1237), .A3(n1221), .ZN(n1208) );
NOR2_X1 U943 ( .A1(n1107), .A2(n1097), .ZN(n1237) );
INV_X1 U944 ( .A(n1272), .ZN(n1107) );
XNOR2_X1 U945 ( .A(G116), .B(n1273), .ZN(G18) );
NAND3_X1 U946 ( .A1(n1071), .A2(n1274), .A3(n1221), .ZN(n1273) );
AND3_X1 U947 ( .A1(n1079), .A2(n1275), .A3(n1094), .ZN(n1221) );
XOR2_X1 U948 ( .A(n1276), .B(KEYINPUT51), .Z(n1079) );
XNOR2_X1 U949 ( .A(KEYINPUT11), .B(n1055), .ZN(n1274) );
NAND2_X1 U950 ( .A1(n1277), .A2(n1270), .ZN(n1055) );
INV_X1 U951 ( .A(n1278), .ZN(n1270) );
XOR2_X1 U952 ( .A(n1207), .B(n1279), .Z(G15) );
NAND2_X1 U953 ( .A1(KEYINPUT27), .A2(G113), .ZN(n1279) );
NAND4_X1 U954 ( .A1(n1094), .A2(n1223), .A3(n1071), .A4(n1219), .ZN(n1207) );
INV_X1 U955 ( .A(n1240), .ZN(n1071) );
NAND2_X1 U956 ( .A1(n1097), .A2(n1272), .ZN(n1240) );
INV_X1 U957 ( .A(n1095), .ZN(n1223) );
NAND2_X1 U958 ( .A1(n1278), .A2(n1101), .ZN(n1095) );
NOR2_X1 U959 ( .A1(n1280), .A2(n1086), .ZN(n1094) );
XNOR2_X1 U960 ( .A(G110), .B(n1209), .ZN(G12) );
NAND3_X1 U961 ( .A1(n1070), .A2(n1222), .A3(n1250), .ZN(n1209) );
INV_X1 U962 ( .A(n1064), .ZN(n1250) );
NAND2_X1 U963 ( .A1(n1278), .A2(n1277), .ZN(n1064) );
XNOR2_X1 U964 ( .A(n1101), .B(KEYINPUT44), .ZN(n1277) );
XNOR2_X1 U965 ( .A(n1281), .B(G475), .ZN(n1101) );
NAND2_X1 U966 ( .A1(n1154), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U967 ( .A(n1283), .B(n1284), .ZN(n1154) );
XNOR2_X1 U968 ( .A(n1285), .B(n1286), .ZN(n1284) );
XOR2_X1 U969 ( .A(n1287), .B(n1128), .Z(n1286) );
XNOR2_X1 U970 ( .A(n1258), .B(G140), .ZN(n1128) );
INV_X1 U971 ( .A(G125), .ZN(n1258) );
NAND2_X1 U972 ( .A1(n1288), .A2(G214), .ZN(n1287) );
XOR2_X1 U973 ( .A(n1289), .B(n1290), .Z(n1283) );
XNOR2_X1 U974 ( .A(KEYINPUT6), .B(n1127), .ZN(n1290) );
NAND2_X1 U975 ( .A1(n1291), .A2(n1292), .ZN(n1289) );
OR2_X1 U976 ( .A1(n1293), .A2(G104), .ZN(n1292) );
XOR2_X1 U977 ( .A(n1294), .B(KEYINPUT32), .Z(n1291) );
NAND2_X1 U978 ( .A1(G104), .A2(n1293), .ZN(n1294) );
XOR2_X1 U979 ( .A(G113), .B(G122), .Z(n1293) );
NOR2_X1 U980 ( .A1(n1112), .A2(n1295), .ZN(n1278) );
AND2_X1 U981 ( .A1(G478), .A2(n1114), .ZN(n1295) );
NOR2_X1 U982 ( .A1(n1114), .A2(G478), .ZN(n1112) );
NAND2_X1 U983 ( .A1(n1296), .A2(n1282), .ZN(n1114) );
XOR2_X1 U984 ( .A(n1152), .B(KEYINPUT58), .Z(n1296) );
NAND2_X1 U985 ( .A1(n1297), .A2(n1298), .ZN(n1152) );
NAND2_X1 U986 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U987 ( .A(KEYINPUT28), .B(n1301), .Z(n1297) );
NOR2_X1 U988 ( .A1(n1299), .A2(n1300), .ZN(n1301) );
NAND3_X1 U989 ( .A1(G234), .A2(n1090), .A3(G217), .ZN(n1300) );
XNOR2_X1 U990 ( .A(n1302), .B(n1303), .ZN(n1299) );
XOR2_X1 U991 ( .A(G122), .B(n1304), .Z(n1303) );
XOR2_X1 U992 ( .A(G143), .B(G134), .Z(n1304) );
XOR2_X1 U993 ( .A(n1305), .B(n1306), .Z(n1302) );
XNOR2_X1 U994 ( .A(n1051), .B(n1307), .ZN(n1306) );
NOR2_X1 U995 ( .A1(G116), .A2(KEYINPUT9), .ZN(n1307) );
NAND2_X1 U996 ( .A1(KEYINPUT3), .A2(n1308), .ZN(n1305) );
INV_X1 U997 ( .A(n1056), .ZN(n1222) );
NAND2_X1 U998 ( .A1(n1085), .A2(n1219), .ZN(n1056) );
AND2_X1 U999 ( .A1(n1276), .A2(n1275), .ZN(n1219) );
NAND2_X1 U1000 ( .A1(n1072), .A2(n1309), .ZN(n1275) );
NAND4_X1 U1001 ( .A1(G902), .A2(G953), .A3(n1265), .A4(n1310), .ZN(n1309) );
INV_X1 U1002 ( .A(G898), .ZN(n1310) );
NAND3_X1 U1003 ( .A1(n1265), .A2(n1090), .A3(n1311), .ZN(n1072) );
XOR2_X1 U1004 ( .A(KEYINPUT12), .B(G952), .Z(n1311) );
NAND2_X1 U1005 ( .A1(G237), .A2(G234), .ZN(n1265) );
AND2_X1 U1006 ( .A1(n1080), .A2(n1081), .ZN(n1276) );
NAND2_X1 U1007 ( .A1(G214), .A2(n1312), .ZN(n1081) );
XNOR2_X1 U1008 ( .A(n1313), .B(n1105), .ZN(n1080) );
NAND2_X1 U1009 ( .A1(G210), .A2(n1312), .ZN(n1105) );
NAND2_X1 U1010 ( .A1(n1314), .A2(n1282), .ZN(n1312) );
INV_X1 U1011 ( .A(G237), .ZN(n1314) );
NAND2_X1 U1012 ( .A1(KEYINPUT13), .A2(n1106), .ZN(n1313) );
NAND2_X1 U1013 ( .A1(n1315), .A2(n1282), .ZN(n1106) );
XOR2_X1 U1014 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1015 ( .A(n1318), .B(n1195), .ZN(n1317) );
XOR2_X1 U1016 ( .A(n1138), .B(n1319), .Z(n1195) );
XNOR2_X1 U1017 ( .A(n1320), .B(n1139), .ZN(n1319) );
NAND2_X1 U1018 ( .A1(KEYINPUT16), .A2(n1140), .ZN(n1320) );
NAND2_X1 U1019 ( .A1(n1321), .A2(n1322), .ZN(n1140) );
NAND2_X1 U1020 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1021 ( .A(KEYINPUT4), .B(n1325), .Z(n1323) );
XOR2_X1 U1022 ( .A(G110), .B(G122), .Z(n1138) );
NAND2_X1 U1023 ( .A1(KEYINPUT46), .A2(n1326), .ZN(n1318) );
XNOR2_X1 U1024 ( .A(G125), .B(n1327), .ZN(n1326) );
XNOR2_X1 U1025 ( .A(KEYINPUT23), .B(n1199), .ZN(n1316) );
NAND2_X1 U1026 ( .A1(G224), .A2(n1328), .ZN(n1199) );
XNOR2_X1 U1027 ( .A(KEYINPUT25), .B(n1090), .ZN(n1328) );
INV_X1 U1028 ( .A(n1220), .ZN(n1085) );
NAND2_X1 U1029 ( .A1(n1086), .A2(n1329), .ZN(n1220) );
INV_X1 U1030 ( .A(n1280), .ZN(n1329) );
XNOR2_X1 U1031 ( .A(n1088), .B(KEYINPUT31), .ZN(n1280) );
AND2_X1 U1032 ( .A1(G221), .A2(n1330), .ZN(n1088) );
NAND2_X1 U1033 ( .A1(G234), .A2(n1282), .ZN(n1330) );
XOR2_X1 U1034 ( .A(n1331), .B(n1332), .Z(n1086) );
XOR2_X1 U1035 ( .A(KEYINPUT22), .B(G469), .Z(n1332) );
NAND2_X1 U1036 ( .A1(KEYINPUT1), .A2(n1110), .ZN(n1331) );
NAND2_X1 U1037 ( .A1(n1333), .A2(n1282), .ZN(n1110) );
XOR2_X1 U1038 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1039 ( .A(n1336), .B(n1125), .ZN(n1335) );
XOR2_X1 U1040 ( .A(n1285), .B(n1308), .Z(n1125) );
INV_X1 U1041 ( .A(n1139), .ZN(n1336) );
XOR2_X1 U1042 ( .A(G101), .B(n1337), .Z(n1139) );
XNOR2_X1 U1043 ( .A(n1051), .B(G104), .ZN(n1337) );
INV_X1 U1044 ( .A(G107), .ZN(n1051) );
XNOR2_X1 U1045 ( .A(n1338), .B(n1177), .ZN(n1334) );
NAND2_X1 U1046 ( .A1(KEYINPUT60), .A2(n1339), .ZN(n1338) );
XNOR2_X1 U1047 ( .A(n1174), .B(n1340), .ZN(n1339) );
NOR2_X1 U1048 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
AND2_X1 U1049 ( .A1(KEYINPUT29), .A2(n1187), .ZN(n1342) );
NOR2_X1 U1050 ( .A1(KEYINPUT42), .A2(n1187), .ZN(n1341) );
NAND2_X1 U1051 ( .A1(G227), .A2(n1090), .ZN(n1187) );
XOR2_X1 U1052 ( .A(G110), .B(n1343), .Z(n1174) );
XOR2_X1 U1053 ( .A(KEYINPUT59), .B(G140), .Z(n1343) );
NOR2_X1 U1054 ( .A1(n1272), .A2(n1097), .ZN(n1070) );
AND3_X1 U1055 ( .A1(n1344), .A2(n1345), .A3(n1346), .ZN(n1097) );
NAND2_X1 U1056 ( .A1(n1347), .A2(n1145), .ZN(n1346) );
OR3_X1 U1057 ( .A1(n1145), .A2(n1347), .A3(G902), .ZN(n1345) );
NOR2_X1 U1058 ( .A1(n1348), .A2(G234), .ZN(n1347) );
INV_X1 U1059 ( .A(G217), .ZN(n1348) );
XOR2_X1 U1060 ( .A(n1349), .B(n1350), .Z(n1145) );
XOR2_X1 U1061 ( .A(n1351), .B(n1352), .Z(n1350) );
XNOR2_X1 U1062 ( .A(n1324), .B(G110), .ZN(n1352) );
XOR2_X1 U1063 ( .A(G146), .B(G137), .Z(n1351) );
XNOR2_X1 U1064 ( .A(n1308), .B(n1353), .ZN(n1349) );
XOR2_X1 U1065 ( .A(n1354), .B(n1355), .Z(n1353) );
AND3_X1 U1066 ( .A1(G221), .A2(n1090), .A3(G234), .ZN(n1355) );
INV_X1 U1067 ( .A(G953), .ZN(n1090) );
NOR2_X1 U1068 ( .A1(KEYINPUT57), .A2(n1356), .ZN(n1354) );
XNOR2_X1 U1069 ( .A(G125), .B(n1357), .ZN(n1356) );
NOR2_X1 U1070 ( .A1(G140), .A2(KEYINPUT36), .ZN(n1357) );
NAND2_X1 U1071 ( .A1(G217), .A2(G902), .ZN(n1344) );
XNOR2_X1 U1072 ( .A(n1358), .B(G472), .ZN(n1272) );
NAND2_X1 U1073 ( .A1(n1359), .A2(n1282), .ZN(n1358) );
INV_X1 U1074 ( .A(G902), .ZN(n1282) );
XNOR2_X1 U1075 ( .A(n1167), .B(n1159), .ZN(n1359) );
XNOR2_X1 U1076 ( .A(n1360), .B(G101), .ZN(n1159) );
NAND2_X1 U1077 ( .A1(n1288), .A2(G210), .ZN(n1360) );
NOR2_X1 U1078 ( .A1(G953), .A2(G237), .ZN(n1288) );
INV_X1 U1079 ( .A(n1165), .ZN(n1167) );
XOR2_X1 U1080 ( .A(n1177), .B(n1361), .Z(n1165) );
XNOR2_X1 U1081 ( .A(n1202), .B(n1362), .ZN(n1361) );
NAND2_X1 U1082 ( .A1(n1321), .A2(n1363), .ZN(n1362) );
NAND2_X1 U1083 ( .A1(n1364), .A2(n1324), .ZN(n1363) );
INV_X1 U1084 ( .A(G119), .ZN(n1324) );
XOR2_X1 U1085 ( .A(KEYINPUT38), .B(n1325), .Z(n1364) );
NAND2_X1 U1086 ( .A1(G119), .A2(n1325), .ZN(n1321) );
XOR2_X1 U1087 ( .A(G113), .B(G116), .Z(n1325) );
INV_X1 U1088 ( .A(n1327), .ZN(n1202) );
NAND3_X1 U1089 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1327) );
OR2_X1 U1090 ( .A1(n1308), .A2(n1368), .ZN(n1367) );
NAND3_X1 U1091 ( .A1(n1368), .A2(n1308), .A3(KEYINPUT17), .ZN(n1366) );
XOR2_X1 U1092 ( .A(G128), .B(KEYINPUT10), .Z(n1308) );
AND2_X1 U1093 ( .A1(KEYINPUT54), .A2(n1285), .ZN(n1368) );
OR2_X1 U1094 ( .A1(n1285), .A2(KEYINPUT17), .ZN(n1365) );
XOR2_X1 U1095 ( .A(G143), .B(G146), .Z(n1285) );
XNOR2_X1 U1096 ( .A(n1369), .B(n1124), .ZN(n1177) );
XOR2_X1 U1097 ( .A(G134), .B(G137), .Z(n1124) );
NAND2_X1 U1098 ( .A1(KEYINPUT19), .A2(n1127), .ZN(n1369) );
INV_X1 U1099 ( .A(G131), .ZN(n1127) );
endmodule


