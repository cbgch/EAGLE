//Key = 1111000100101111110101111010001001000101010100001011111110111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284;

XOR2_X1 U704 ( .A(n971), .B(n972), .Z(G9) );
NAND4_X1 U705 ( .A1(n973), .A2(n974), .A3(n975), .A4(n976), .ZN(n972) );
NOR2_X1 U706 ( .A1(n977), .A2(n978), .ZN(n976) );
XNOR2_X1 U707 ( .A(KEYINPUT47), .B(n979), .ZN(n978) );
NOR2_X1 U708 ( .A1(n980), .A2(n981), .ZN(G75) );
NOR4_X1 U709 ( .A1(n982), .A2(n983), .A3(n984), .A4(n985), .ZN(n981) );
INV_X1 U710 ( .A(G952), .ZN(n985) );
NOR4_X1 U711 ( .A1(n986), .A2(n987), .A3(n988), .A4(n989), .ZN(n984) );
NOR2_X1 U712 ( .A1(n990), .A2(n991), .ZN(n986) );
NOR2_X1 U713 ( .A1(n992), .A2(n993), .ZN(n991) );
INV_X1 U714 ( .A(n994), .ZN(n993) );
NOR2_X1 U715 ( .A1(n995), .A2(n996), .ZN(n992) );
NOR2_X1 U716 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR2_X1 U717 ( .A1(n999), .A2(n1000), .ZN(n990) );
NOR2_X1 U718 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U719 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NAND4_X1 U720 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n982) );
NAND3_X1 U721 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1006) );
XOR2_X1 U722 ( .A(n1012), .B(KEYINPUT48), .Z(n1011) );
NAND4_X1 U723 ( .A1(n1013), .A2(n1014), .A3(n974), .A4(n994), .ZN(n1012) );
NAND4_X1 U724 ( .A1(n974), .A2(n994), .A3(n1015), .A4(n1016), .ZN(n1005) );
NAND2_X1 U725 ( .A1(n1017), .A2(n989), .ZN(n1016) );
NAND3_X1 U726 ( .A1(n1014), .A2(n1018), .A3(KEYINPUT40), .ZN(n1017) );
NAND3_X1 U727 ( .A1(n1019), .A2(n1020), .A3(n1013), .ZN(n1015) );
INV_X1 U728 ( .A(n989), .ZN(n1013) );
OR3_X1 U729 ( .A1(n1021), .A2(KEYINPUT40), .A3(n988), .ZN(n1020) );
NAND2_X1 U730 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
OR2_X1 U731 ( .A1(n1024), .A2(n975), .ZN(n1023) );
NOR3_X1 U732 ( .A1(n1025), .A2(G953), .A3(n1026), .ZN(n980) );
INV_X1 U733 ( .A(n1007), .ZN(n1026) );
NAND4_X1 U734 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1007) );
NOR4_X1 U735 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
XOR2_X1 U736 ( .A(n1035), .B(n1036), .Z(n1034) );
XOR2_X1 U737 ( .A(KEYINPUT58), .B(KEYINPUT27), .Z(n1036) );
XOR2_X1 U738 ( .A(n1037), .B(n1038), .Z(n1035) );
AND2_X1 U739 ( .A1(n1039), .A2(G475), .ZN(n1033) );
INV_X1 U740 ( .A(n1004), .ZN(n1032) );
NOR2_X1 U741 ( .A1(n987), .A2(n997), .ZN(n1029) );
XOR2_X1 U742 ( .A(n1040), .B(n1041), .Z(n1028) );
XOR2_X1 U743 ( .A(n1042), .B(KEYINPUT32), .Z(n1027) );
XOR2_X1 U744 ( .A(KEYINPUT57), .B(G952), .Z(n1025) );
XOR2_X1 U745 ( .A(n1043), .B(n1044), .Z(G72) );
NOR2_X1 U746 ( .A1(n1045), .A2(n1008), .ZN(n1044) );
NOR2_X1 U747 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1043) );
NAND2_X1 U749 ( .A1(n1050), .A2(n1008), .ZN(n1049) );
XOR2_X1 U750 ( .A(n1051), .B(n1052), .Z(n1050) );
NAND3_X1 U751 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1051) );
AND3_X1 U752 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
XOR2_X1 U753 ( .A(KEYINPUT63), .B(n1059), .Z(n1054) );
XOR2_X1 U754 ( .A(KEYINPUT35), .B(n1060), .Z(n1053) );
NAND3_X1 U755 ( .A1(G900), .A2(n1052), .A3(G953), .ZN(n1048) );
XOR2_X1 U756 ( .A(n1061), .B(n1062), .Z(n1052) );
XOR2_X1 U757 ( .A(n1063), .B(n1064), .Z(n1062) );
XNOR2_X1 U758 ( .A(G143), .B(KEYINPUT42), .ZN(n1064) );
NAND3_X1 U759 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1063) );
NAND2_X1 U760 ( .A1(KEYINPUT5), .A2(n1068), .ZN(n1067) );
OR3_X1 U761 ( .A1(n1068), .A2(KEYINPUT5), .A3(n1069), .ZN(n1066) );
NAND2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NAND2_X1 U763 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
INV_X1 U764 ( .A(KEYINPUT5), .ZN(n1072) );
XOR2_X1 U765 ( .A(n1068), .B(KEYINPUT53), .Z(n1071) );
XNOR2_X1 U766 ( .A(G134), .B(G137), .ZN(n1069) );
XOR2_X1 U767 ( .A(n1073), .B(n1074), .Z(n1061) );
XOR2_X1 U768 ( .A(n1075), .B(n1076), .Z(G69) );
NOR2_X1 U769 ( .A1(n1077), .A2(n1008), .ZN(n1076) );
NOR2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1075) );
NAND3_X1 U772 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NAND2_X1 U773 ( .A1(G953), .A2(n1079), .ZN(n1083) );
OR2_X1 U774 ( .A1(n1082), .A2(n1084), .ZN(n1080) );
NAND2_X1 U775 ( .A1(n1008), .A2(n1085), .ZN(n1084) );
NAND3_X1 U776 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
AND3_X1 U777 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
XNOR2_X1 U778 ( .A(n1092), .B(KEYINPUT37), .ZN(n1086) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1082) );
NOR2_X1 U780 ( .A1(n1095), .A2(n1096), .ZN(G66) );
NOR3_X1 U781 ( .A1(n1037), .A2(n1097), .A3(n1098), .ZN(n1096) );
NOR2_X1 U782 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR2_X1 U783 ( .A1(n1101), .A2(n1038), .ZN(n1099) );
INV_X1 U784 ( .A(n983), .ZN(n1101) );
NOR3_X1 U785 ( .A1(n1102), .A2(n1038), .A3(n1103), .ZN(n1097) );
INV_X1 U786 ( .A(n1100), .ZN(n1102) );
NOR2_X1 U787 ( .A1(n1095), .A2(n1104), .ZN(G63) );
XOR2_X1 U788 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U789 ( .A1(n1041), .A2(n1103), .ZN(n1105) );
INV_X1 U790 ( .A(G478), .ZN(n1041) );
NOR2_X1 U791 ( .A1(n1095), .A2(n1107), .ZN(G60) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND3_X1 U793 ( .A1(G475), .A2(n983), .A3(n1110), .ZN(n1108) );
XOR2_X1 U794 ( .A(n1111), .B(KEYINPUT13), .Z(n1110) );
XOR2_X1 U795 ( .A(G104), .B(n1112), .Z(G6) );
NOR2_X1 U796 ( .A1(n1095), .A2(n1113), .ZN(G57) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1113) );
XNOR2_X1 U798 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U799 ( .A1(KEYINPUT12), .A2(n1118), .ZN(n1116) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(n1120) );
NAND2_X1 U802 ( .A1(KEYINPUT39), .A2(n1123), .ZN(n1121) );
XOR2_X1 U803 ( .A(G113), .B(n1124), .Z(n1119) );
NOR2_X1 U804 ( .A1(n1125), .A2(n1103), .ZN(n1124) );
INV_X1 U805 ( .A(G472), .ZN(n1125) );
NAND2_X1 U806 ( .A1(KEYINPUT24), .A2(G101), .ZN(n1114) );
NOR2_X1 U807 ( .A1(n1095), .A2(n1126), .ZN(G54) );
XOR2_X1 U808 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U809 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1103), .ZN(n1130) );
INV_X1 U811 ( .A(G469), .ZN(n1131) );
XOR2_X1 U812 ( .A(n1132), .B(n1133), .Z(n1127) );
NOR2_X1 U813 ( .A1(KEYINPUT11), .A2(n1134), .ZN(n1133) );
XNOR2_X1 U814 ( .A(n1135), .B(n1136), .ZN(n1134) );
NOR2_X1 U815 ( .A1(n1095), .A2(n1137), .ZN(G51) );
XOR2_X1 U816 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1103), .ZN(n1138) );
NAND2_X1 U818 ( .A1(G902), .A2(n983), .ZN(n1103) );
NAND4_X1 U819 ( .A1(n1092), .A2(n1060), .A3(n1141), .A4(n1142), .ZN(n983) );
AND4_X1 U820 ( .A1(n1143), .A2(n1057), .A3(n1091), .A4(n1089), .ZN(n1142) );
AND2_X1 U821 ( .A1(n1056), .A2(n1058), .ZN(n1143) );
NOR3_X1 U822 ( .A1(n1144), .A2(n1059), .A3(n1145), .ZN(n1141) );
INV_X1 U823 ( .A(n1087), .ZN(n1145) );
NAND4_X1 U824 ( .A1(n1146), .A2(n1147), .A3(n975), .A4(n1148), .ZN(n1087) );
XOR2_X1 U825 ( .A(KEYINPUT38), .B(n1018), .Z(n1148) );
XOR2_X1 U826 ( .A(n1149), .B(KEYINPUT10), .Z(n1146) );
AND2_X1 U827 ( .A1(n1150), .A2(n1018), .ZN(n1059) );
XNOR2_X1 U828 ( .A(n1151), .B(KEYINPUT50), .ZN(n1150) );
XOR2_X1 U829 ( .A(n1090), .B(KEYINPUT19), .Z(n1144) );
AND4_X1 U830 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1060) );
NOR3_X1 U831 ( .A1(n1112), .A2(n1156), .A3(n1157), .ZN(n1092) );
AND2_X1 U832 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U833 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U834 ( .A1(n975), .A2(n974), .ZN(n1161) );
NAND2_X1 U835 ( .A1(n996), .A2(n1014), .ZN(n1160) );
AND3_X1 U836 ( .A1(n1024), .A2(n974), .A3(n1158), .ZN(n1112) );
INV_X1 U837 ( .A(n1162), .ZN(n1158) );
NOR2_X1 U838 ( .A1(n1008), .A2(G952), .ZN(n1095) );
XNOR2_X1 U839 ( .A(G146), .B(n1152), .ZN(G48) );
NAND3_X1 U840 ( .A1(n1163), .A2(n1018), .A3(n1024), .ZN(n1152) );
XNOR2_X1 U841 ( .A(G143), .B(n1153), .ZN(G45) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1165), .ZN(n1153) );
XNOR2_X1 U843 ( .A(n1154), .B(n1166), .ZN(G42) );
XOR2_X1 U844 ( .A(KEYINPUT8), .B(G140), .Z(n1166) );
NAND3_X1 U845 ( .A1(n1022), .A2(n1002), .A3(n1167), .ZN(n1154) );
XNOR2_X1 U846 ( .A(G137), .B(n1155), .ZN(G39) );
NAND3_X1 U847 ( .A1(n1014), .A2(n1022), .A3(n1163), .ZN(n1155) );
XNOR2_X1 U848 ( .A(G134), .B(n1056), .ZN(G36) );
NAND3_X1 U849 ( .A1(n1022), .A2(n975), .A3(n1164), .ZN(n1056) );
XNOR2_X1 U850 ( .A(n1058), .B(n1168), .ZN(G33) );
NOR2_X1 U851 ( .A1(KEYINPUT49), .A2(n1068), .ZN(n1168) );
NAND3_X1 U852 ( .A1(n1164), .A2(n1022), .A3(n1024), .ZN(n1058) );
INV_X1 U853 ( .A(n987), .ZN(n1022) );
NAND2_X1 U854 ( .A1(n1009), .A2(n1169), .ZN(n987) );
AND3_X1 U855 ( .A1(n1002), .A2(n1170), .A3(n996), .ZN(n1164) );
XNOR2_X1 U856 ( .A(G128), .B(n1057), .ZN(G30) );
NAND3_X1 U857 ( .A1(n975), .A2(n1018), .A3(n1163), .ZN(n1057) );
AND4_X1 U858 ( .A1(n1171), .A2(n1002), .A3(n1172), .A4(n1170), .ZN(n1163) );
XOR2_X1 U859 ( .A(G101), .B(n1173), .Z(G3) );
NOR4_X1 U860 ( .A1(KEYINPUT45), .A2(n988), .A3(n1149), .A4(n1162), .ZN(n1173) );
XOR2_X1 U861 ( .A(n1174), .B(n1175), .Z(G27) );
NAND2_X1 U862 ( .A1(n1151), .A2(n1018), .ZN(n1175) );
AND2_X1 U863 ( .A1(n1167), .A2(n994), .ZN(n1151) );
AND4_X1 U864 ( .A1(n1024), .A2(n1171), .A3(n1176), .A4(n1170), .ZN(n1167) );
NAND2_X1 U865 ( .A1(n989), .A2(n1177), .ZN(n1170) );
NAND4_X1 U866 ( .A1(G953), .A2(G902), .A3(n1178), .A4(n1047), .ZN(n1177) );
INV_X1 U867 ( .A(G900), .ZN(n1047) );
XOR2_X1 U868 ( .A(n1179), .B(n1089), .Z(G24) );
NAND3_X1 U869 ( .A1(n1147), .A2(n974), .A3(n1165), .ZN(n1089) );
NOR3_X1 U870 ( .A1(n1180), .A2(n1181), .A3(n1021), .ZN(n1165) );
INV_X1 U871 ( .A(n1000), .ZN(n974) );
NAND2_X1 U872 ( .A1(n1176), .A2(n998), .ZN(n1000) );
XNOR2_X1 U873 ( .A(G119), .B(n1091), .ZN(G21) );
NAND4_X1 U874 ( .A1(n1014), .A2(n1171), .A3(n1182), .A4(n1147), .ZN(n1091) );
NOR2_X1 U875 ( .A1(n1183), .A2(n1021), .ZN(n1182) );
INV_X1 U876 ( .A(n998), .ZN(n1171) );
INV_X1 U877 ( .A(n988), .ZN(n1014) );
XNOR2_X1 U878 ( .A(G116), .B(n1184), .ZN(G18) );
NAND4_X1 U879 ( .A1(n996), .A2(n1147), .A3(n975), .A4(n1018), .ZN(n1184) );
NOR2_X1 U880 ( .A1(n1185), .A2(n1180), .ZN(n975) );
XOR2_X1 U881 ( .A(n1186), .B(n1187), .Z(G15) );
XOR2_X1 U882 ( .A(KEYINPUT18), .B(G113), .Z(n1187) );
NAND2_X1 U883 ( .A1(KEYINPUT3), .A2(n1090), .ZN(n1186) );
NAND4_X1 U884 ( .A1(n1024), .A2(n996), .A3(n973), .A4(n1147), .ZN(n1090) );
AND2_X1 U885 ( .A1(n994), .A2(n979), .ZN(n1147) );
NAND2_X1 U886 ( .A1(n1188), .A2(n1189), .ZN(n994) );
OR2_X1 U887 ( .A1(n977), .A2(KEYINPUT15), .ZN(n1189) );
NAND3_X1 U888 ( .A1(n1042), .A2(n1004), .A3(KEYINPUT15), .ZN(n1188) );
INV_X1 U889 ( .A(n1149), .ZN(n996) );
NAND2_X1 U890 ( .A1(n1172), .A2(n998), .ZN(n1149) );
INV_X1 U891 ( .A(n1183), .ZN(n1172) );
XOR2_X1 U892 ( .A(n1176), .B(KEYINPUT6), .Z(n1183) );
NOR2_X1 U893 ( .A1(n1190), .A2(n1181), .ZN(n1024) );
INV_X1 U894 ( .A(n1180), .ZN(n1190) );
XOR2_X1 U895 ( .A(n1191), .B(n1156), .Z(G12) );
NOR4_X1 U896 ( .A1(n1162), .A2(n988), .A3(n997), .A4(n998), .ZN(n1156) );
NAND3_X1 U897 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n998) );
NAND2_X1 U898 ( .A1(n1037), .A2(n1195), .ZN(n1194) );
INV_X1 U899 ( .A(KEYINPUT59), .ZN(n1195) );
NAND3_X1 U900 ( .A1(KEYINPUT59), .A2(n1196), .A3(n1038), .ZN(n1193) );
OR2_X1 U901 ( .A1(n1038), .A2(n1196), .ZN(n1192) );
NOR2_X1 U902 ( .A1(n1037), .A2(KEYINPUT61), .ZN(n1196) );
NOR2_X1 U903 ( .A1(n1100), .A2(G902), .ZN(n1037) );
XOR2_X1 U904 ( .A(n1197), .B(n1198), .Z(n1100) );
XNOR2_X1 U905 ( .A(n1135), .B(n1199), .ZN(n1198) );
NAND2_X1 U906 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U907 ( .A1(KEYINPUT1), .A2(n1202), .ZN(n1201) );
XOR2_X1 U908 ( .A(n1174), .B(G140), .Z(n1202) );
OR3_X1 U909 ( .A1(n1132), .A2(G125), .A3(KEYINPUT1), .ZN(n1200) );
XOR2_X1 U910 ( .A(n1203), .B(n1204), .Z(n1197) );
AND2_X1 U911 ( .A1(G221), .A2(n1205), .ZN(n1204) );
XOR2_X1 U912 ( .A(n1206), .B(G137), .Z(n1203) );
NAND2_X1 U913 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U914 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U915 ( .A(KEYINPUT7), .B(n1211), .Z(n1207) );
NOR2_X1 U916 ( .A1(n1209), .A2(n1210), .ZN(n1211) );
XOR2_X1 U917 ( .A(n1212), .B(G128), .Z(n1209) );
NAND2_X1 U918 ( .A1(KEYINPUT21), .A2(G119), .ZN(n1212) );
NAND2_X1 U919 ( .A1(G217), .A2(n1213), .ZN(n1038) );
INV_X1 U920 ( .A(n1176), .ZN(n997) );
XOR2_X1 U921 ( .A(n1214), .B(G472), .Z(n1176) );
NAND2_X1 U922 ( .A1(n1215), .A2(n1111), .ZN(n1214) );
XOR2_X1 U923 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U924 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U925 ( .A(n1122), .B(n1123), .Z(n1219) );
XOR2_X1 U926 ( .A(n1220), .B(n1221), .Z(n1123) );
XNOR2_X1 U927 ( .A(n1222), .B(n1223), .ZN(n1220) );
XOR2_X1 U928 ( .A(n1224), .B(KEYINPUT31), .Z(n1122) );
NAND2_X1 U929 ( .A1(KEYINPUT52), .A2(n1225), .ZN(n1224) );
XOR2_X1 U930 ( .A(n1117), .B(n1226), .Z(n1218) );
NAND2_X1 U931 ( .A1(G210), .A2(n1227), .ZN(n1117) );
XOR2_X1 U932 ( .A(n1228), .B(n1229), .Z(n1216) );
XNOR2_X1 U933 ( .A(KEYINPUT29), .B(KEYINPUT16), .ZN(n1229) );
XNOR2_X1 U934 ( .A(KEYINPUT60), .B(KEYINPUT44), .ZN(n1228) );
NAND2_X1 U935 ( .A1(n1180), .A2(n1181), .ZN(n988) );
INV_X1 U936 ( .A(n1185), .ZN(n1181) );
NAND2_X1 U937 ( .A1(n1230), .A2(n1231), .ZN(n1185) );
NAND2_X1 U938 ( .A1(G475), .A2(n1039), .ZN(n1231) );
XOR2_X1 U939 ( .A(KEYINPUT30), .B(n1031), .Z(n1230) );
NOR2_X1 U940 ( .A1(n1039), .A2(G475), .ZN(n1031) );
NAND2_X1 U941 ( .A1(n1109), .A2(n1111), .ZN(n1039) );
XOR2_X1 U942 ( .A(n1232), .B(n1233), .Z(n1109) );
XOR2_X1 U943 ( .A(G104), .B(n1234), .Z(n1233) );
NOR2_X1 U944 ( .A1(KEYINPUT36), .A2(n1235), .ZN(n1234) );
XOR2_X1 U945 ( .A(n1073), .B(n1236), .Z(n1235) );
XOR2_X1 U946 ( .A(n1237), .B(G125), .Z(n1236) );
NAND2_X1 U947 ( .A1(KEYINPUT23), .A2(n1238), .ZN(n1237) );
XOR2_X1 U948 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U949 ( .A(G143), .B(n1068), .Z(n1240) );
INV_X1 U950 ( .A(G131), .ZN(n1068) );
NAND2_X1 U951 ( .A1(G214), .A2(n1227), .ZN(n1239) );
NOR2_X1 U952 ( .A1(G953), .A2(G237), .ZN(n1227) );
XOR2_X1 U953 ( .A(G113), .B(n1179), .Z(n1232) );
XOR2_X1 U954 ( .A(n1241), .B(G478), .Z(n1180) );
NAND2_X1 U955 ( .A1(KEYINPUT41), .A2(n1040), .ZN(n1241) );
NOR2_X1 U956 ( .A1(n1106), .A2(G902), .ZN(n1040) );
XNOR2_X1 U957 ( .A(n1242), .B(n1243), .ZN(n1106) );
XOR2_X1 U958 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND2_X1 U959 ( .A1(G217), .A2(n1205), .ZN(n1245) );
AND2_X1 U960 ( .A1(G234), .A2(n1008), .ZN(n1205) );
NAND2_X1 U961 ( .A1(KEYINPUT62), .A2(n1246), .ZN(n1244) );
XNOR2_X1 U962 ( .A(n1247), .B(n1248), .ZN(n1246) );
XOR2_X1 U963 ( .A(n1249), .B(G107), .Z(n1248) );
NAND2_X1 U964 ( .A1(KEYINPUT0), .A2(n1179), .ZN(n1249) );
INV_X1 U965 ( .A(G122), .ZN(n1179) );
NAND3_X1 U966 ( .A1(n973), .A2(n979), .A3(n1002), .ZN(n1162) );
INV_X1 U967 ( .A(n977), .ZN(n1002) );
NAND2_X1 U968 ( .A1(n1003), .A2(n1004), .ZN(n977) );
NAND2_X1 U969 ( .A1(G221), .A2(n1213), .ZN(n1004) );
NAND2_X1 U970 ( .A1(G234), .A2(n1111), .ZN(n1213) );
INV_X1 U971 ( .A(n1042), .ZN(n1003) );
XOR2_X1 U972 ( .A(n1250), .B(G469), .Z(n1042) );
NAND2_X1 U973 ( .A1(n1251), .A2(n1111), .ZN(n1250) );
XOR2_X1 U974 ( .A(n1252), .B(n1136), .Z(n1251) );
XNOR2_X1 U975 ( .A(n1253), .B(n1254), .ZN(n1136) );
XOR2_X1 U976 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U977 ( .A(KEYINPUT43), .B(G101), .Z(n1256) );
NOR4_X1 U978 ( .A1(n1257), .A2(n1258), .A3(KEYINPUT28), .A4(n1259), .ZN(n1255) );
AND2_X1 U979 ( .A1(n1260), .A2(KEYINPUT46), .ZN(n1259) );
NOR2_X1 U980 ( .A1(n1261), .A2(n971), .ZN(n1258) );
INV_X1 U981 ( .A(G107), .ZN(n971) );
NOR2_X1 U982 ( .A1(n1260), .A2(n1262), .ZN(n1261) );
NOR4_X1 U983 ( .A1(G107), .A2(n1262), .A3(KEYINPUT46), .A4(n1260), .ZN(n1257) );
XNOR2_X1 U984 ( .A(G104), .B(KEYINPUT33), .ZN(n1260) );
INV_X1 U985 ( .A(KEYINPUT26), .ZN(n1262) );
XOR2_X1 U986 ( .A(n1242), .B(n1222), .Z(n1253) );
XOR2_X1 U987 ( .A(G137), .B(G131), .Z(n1222) );
XNOR2_X1 U988 ( .A(G143), .B(n1221), .ZN(n1242) );
XOR2_X1 U989 ( .A(G134), .B(G128), .Z(n1221) );
XOR2_X1 U990 ( .A(n1073), .B(n1263), .Z(n1252) );
INV_X1 U991 ( .A(n1129), .ZN(n1263) );
XOR2_X1 U992 ( .A(n1210), .B(n1264), .Z(n1129) );
NOR2_X1 U993 ( .A1(G953), .A2(n1046), .ZN(n1264) );
INV_X1 U994 ( .A(G227), .ZN(n1046) );
XOR2_X1 U995 ( .A(n1132), .B(n1135), .Z(n1073) );
INV_X1 U996 ( .A(G140), .ZN(n1132) );
NAND2_X1 U997 ( .A1(n989), .A2(n1265), .ZN(n979) );
NAND4_X1 U998 ( .A1(G953), .A2(G902), .A3(n1178), .A4(n1079), .ZN(n1265) );
INV_X1 U999 ( .A(G898), .ZN(n1079) );
NAND3_X1 U1000 ( .A1(n1178), .A2(n1008), .A3(G952), .ZN(n989) );
INV_X1 U1001 ( .A(G953), .ZN(n1008) );
NAND2_X1 U1002 ( .A1(G237), .A2(G234), .ZN(n1178) );
XOR2_X1 U1003 ( .A(n1021), .B(KEYINPUT2), .Z(n973) );
INV_X1 U1004 ( .A(n1018), .ZN(n1021) );
NOR2_X1 U1005 ( .A1(n1009), .A2(n1010), .ZN(n1018) );
INV_X1 U1006 ( .A(n1169), .ZN(n1010) );
NAND2_X1 U1007 ( .A1(G214), .A2(n1266), .ZN(n1169) );
XNOR2_X1 U1008 ( .A(n1267), .B(n1140), .ZN(n1009) );
NAND2_X1 U1009 ( .A1(G210), .A2(n1266), .ZN(n1140) );
NAND2_X1 U1010 ( .A1(n1111), .A2(n1268), .ZN(n1266) );
INV_X1 U1011 ( .A(G237), .ZN(n1268) );
NAND2_X1 U1012 ( .A1(n1269), .A2(n1111), .ZN(n1267) );
INV_X1 U1013 ( .A(G902), .ZN(n1111) );
XOR2_X1 U1014 ( .A(KEYINPUT22), .B(n1139), .Z(n1269) );
XNOR2_X1 U1015 ( .A(n1270), .B(n1271), .ZN(n1139) );
XNOR2_X1 U1016 ( .A(n1093), .B(n1074), .ZN(n1271) );
XNOR2_X1 U1017 ( .A(n1174), .B(G128), .ZN(n1074) );
INV_X1 U1018 ( .A(G125), .ZN(n1174) );
XOR2_X1 U1019 ( .A(n1272), .B(n1273), .Z(n1093) );
XOR2_X1 U1020 ( .A(G107), .B(n1274), .Z(n1273) );
NOR2_X1 U1021 ( .A1(KEYINPUT25), .A2(n1225), .ZN(n1274) );
XOR2_X1 U1022 ( .A(G119), .B(n1247), .Z(n1225) );
XOR2_X1 U1023 ( .A(G116), .B(KEYINPUT20), .Z(n1247) );
XNOR2_X1 U1024 ( .A(n1275), .B(n1226), .ZN(n1272) );
XNOR2_X1 U1025 ( .A(G101), .B(G113), .ZN(n1226) );
NAND2_X1 U1026 ( .A1(KEYINPUT14), .A2(n1276), .ZN(n1275) );
INV_X1 U1027 ( .A(G104), .ZN(n1276) );
XOR2_X1 U1028 ( .A(n1277), .B(n1278), .Z(n1270) );
NOR2_X1 U1029 ( .A1(G953), .A2(n1078), .ZN(n1278) );
INV_X1 U1030 ( .A(G224), .ZN(n1078) );
XOR2_X1 U1031 ( .A(n1279), .B(n1223), .Z(n1277) );
NOR2_X1 U1032 ( .A1(KEYINPUT34), .A2(n1280), .ZN(n1223) );
XNOR2_X1 U1033 ( .A(G143), .B(n1135), .ZN(n1280) );
XOR2_X1 U1034 ( .A(G146), .B(KEYINPUT9), .Z(n1135) );
NAND2_X1 U1035 ( .A1(n1281), .A2(KEYINPUT17), .ZN(n1279) );
XNOR2_X1 U1036 ( .A(n1094), .B(KEYINPUT4), .ZN(n1281) );
XNOR2_X1 U1037 ( .A(n1282), .B(n1283), .ZN(n1094) );
XOR2_X1 U1038 ( .A(KEYINPUT51), .B(G110), .Z(n1283) );
NAND2_X1 U1039 ( .A1(KEYINPUT54), .A2(n1284), .ZN(n1282) );
XOR2_X1 U1040 ( .A(KEYINPUT55), .B(G122), .Z(n1284) );
NAND2_X1 U1041 ( .A1(KEYINPUT56), .A2(n1210), .ZN(n1191) );
INV_X1 U1042 ( .A(G110), .ZN(n1210) );
endmodule


