//Key = 0000010111000011010101111001010111111101011001000111101100111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321;

XOR2_X1 U736 ( .A(G107), .B(n1010), .Z(G9) );
NOR2_X1 U737 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
XNOR2_X1 U738 ( .A(n1013), .B(KEYINPUT1), .ZN(n1011) );
NOR2_X1 U739 ( .A1(n1014), .A2(n1015), .ZN(G75) );
NOR4_X1 U740 ( .A1(G953), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1015) );
NOR2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NOR2_X1 U742 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NOR2_X1 U743 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U744 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U745 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U746 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U747 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1029) );
NOR2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR3_X1 U752 ( .A1(n1038), .A2(n1041), .A3(n1032), .ZN(n1025) );
NOR3_X1 U753 ( .A1(n1038), .A2(n1042), .A3(n1032), .ZN(n1021) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1045), .A2(n1028), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR3_X1 U758 ( .A1(n1016), .A2(G953), .A3(G952), .ZN(n1014) );
AND2_X1 U759 ( .A1(n1050), .A2(n1051), .ZN(n1016) );
NOR4_X1 U760 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
INV_X1 U761 ( .A(n1036), .ZN(n1053) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
XOR2_X1 U763 ( .A(n1058), .B(KEYINPUT3), .Z(n1057) );
NOR4_X1 U764 ( .A1(n1059), .A2(n1060), .A3(n1028), .A4(n1061), .ZN(n1050) );
XOR2_X1 U765 ( .A(KEYINPUT12), .B(n1048), .Z(n1061) );
INV_X1 U766 ( .A(n1062), .ZN(n1048) );
XOR2_X1 U767 ( .A(n1063), .B(n1064), .Z(n1059) );
XOR2_X1 U768 ( .A(n1065), .B(KEYINPUT21), .Z(n1063) );
XOR2_X1 U769 ( .A(n1066), .B(n1067), .Z(G72) );
XNOR2_X1 U770 ( .A(n1068), .B(n1069), .ZN(n1067) );
NOR2_X1 U771 ( .A1(KEYINPUT48), .A2(n1070), .ZN(n1069) );
NOR2_X1 U772 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U773 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
XNOR2_X1 U774 ( .A(G227), .B(KEYINPUT38), .ZN(n1073) );
NAND3_X1 U775 ( .A1(KEYINPUT32), .A2(n1075), .A3(n1076), .ZN(n1068) );
XOR2_X1 U776 ( .A(n1077), .B(n1078), .Z(n1076) );
XOR2_X1 U777 ( .A(n1079), .B(n1080), .Z(n1078) );
OR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U779 ( .A(n1083), .B(n1084), .Z(n1077) );
NAND2_X1 U780 ( .A1(n1085), .A2(n1074), .ZN(n1075) );
NAND2_X1 U781 ( .A1(n1086), .A2(n1087), .ZN(n1066) );
XOR2_X1 U782 ( .A(n1088), .B(n1089), .Z(G69) );
XOR2_X1 U783 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U784 ( .A1(G953), .A2(n1092), .ZN(n1091) );
NOR2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U786 ( .A1(n1095), .A2(n1096), .ZN(n1090) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1096) );
INV_X1 U788 ( .A(n1072), .ZN(n1095) );
XOR2_X1 U789 ( .A(n1086), .B(KEYINPUT63), .Z(n1072) );
NAND2_X1 U790 ( .A1(n1097), .A2(n1098), .ZN(n1088) );
NAND2_X1 U791 ( .A1(n1085), .A2(n1099), .ZN(n1098) );
XOR2_X1 U792 ( .A(n1100), .B(n1101), .Z(n1097) );
NOR2_X1 U793 ( .A1(KEYINPUT44), .A2(n1102), .ZN(n1100) );
NOR2_X1 U794 ( .A1(n1103), .A2(n1104), .ZN(G66) );
XOR2_X1 U795 ( .A(KEYINPUT40), .B(n1105), .Z(n1104) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(n1103) );
NAND4_X1 U797 ( .A1(KEYINPUT27), .A2(G902), .A3(G217), .A4(n1108), .ZN(n1106) );
XNOR2_X1 U798 ( .A(KEYINPUT22), .B(n1018), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1105), .A2(n1109), .ZN(G63) );
XOR2_X1 U800 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U801 ( .A(KEYINPUT9), .B(n1112), .Z(n1111) );
NOR2_X1 U802 ( .A1(KEYINPUT13), .A2(n1113), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(n1110) );
INV_X1 U804 ( .A(G478), .ZN(n1114) );
NOR2_X1 U805 ( .A1(n1105), .A2(n1116), .ZN(G60) );
XNOR2_X1 U806 ( .A(n1117), .B(n1118), .ZN(n1116) );
NOR2_X1 U807 ( .A1(n1119), .A2(n1115), .ZN(n1118) );
INV_X1 U808 ( .A(G475), .ZN(n1119) );
XNOR2_X1 U809 ( .A(G104), .B(n1120), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1105), .A2(n1121), .ZN(G57) );
XOR2_X1 U811 ( .A(n1122), .B(n1123), .Z(n1121) );
XNOR2_X1 U812 ( .A(n1124), .B(KEYINPUT39), .ZN(n1123) );
NAND2_X1 U813 ( .A1(n1125), .A2(KEYINPUT41), .ZN(n1124) );
XOR2_X1 U814 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U815 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U816 ( .A1(n1065), .A2(n1115), .ZN(n1128) );
XOR2_X1 U817 ( .A(n1130), .B(KEYINPUT55), .Z(n1126) );
NAND2_X1 U818 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U819 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U820 ( .A(n1135), .B(KEYINPUT25), .Z(n1131) );
NAND2_X1 U821 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NOR2_X1 U822 ( .A1(n1105), .A2(n1138), .ZN(G54) );
XOR2_X1 U823 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U824 ( .A1(n1141), .A2(n1115), .ZN(n1140) );
INV_X1 U825 ( .A(G469), .ZN(n1141) );
NAND2_X1 U826 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
XOR2_X1 U827 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U828 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U829 ( .A1(G110), .A2(KEYINPUT47), .ZN(n1147) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1144) );
NOR2_X1 U831 ( .A1(KEYINPUT26), .A2(n1133), .ZN(n1149) );
XOR2_X1 U832 ( .A(KEYINPUT37), .B(KEYINPUT2), .Z(n1142) );
NOR2_X1 U833 ( .A1(n1105), .A2(n1150), .ZN(G51) );
XOR2_X1 U834 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U835 ( .A1(n1058), .A2(n1115), .ZN(n1152) );
NAND2_X1 U836 ( .A1(G902), .A2(n1018), .ZN(n1115) );
OR3_X1 U837 ( .A1(n1087), .A2(n1094), .A3(n1153), .ZN(n1018) );
XNOR2_X1 U838 ( .A(n1093), .B(KEYINPUT33), .ZN(n1153) );
NAND4_X1 U839 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1093) );
NAND4_X1 U840 ( .A1(n1158), .A2(n1120), .A3(n1159), .A4(n1160), .ZN(n1094) );
NAND3_X1 U841 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1120) );
NAND2_X1 U842 ( .A1(n1164), .A2(n1013), .ZN(n1158) );
AND4_X1 U843 ( .A1(n1047), .A2(n1162), .A3(n1165), .A4(n1166), .ZN(n1013) );
NAND4_X1 U844 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1087) );
AND3_X1 U845 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
NAND2_X1 U846 ( .A1(n1174), .A2(n1175), .ZN(n1169) );
NAND3_X1 U847 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1175) );
XOR2_X1 U848 ( .A(KEYINPUT31), .B(n1179), .Z(n1178) );
NOR3_X1 U849 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1179) );
XOR2_X1 U850 ( .A(KEYINPUT60), .B(n1047), .Z(n1180) );
NAND2_X1 U851 ( .A1(n1040), .A2(n1183), .ZN(n1177) );
NAND2_X1 U852 ( .A1(n1184), .A2(n1185), .ZN(n1176) );
NAND2_X1 U853 ( .A1(KEYINPUT19), .A2(n1186), .ZN(n1151) );
XOR2_X1 U854 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U855 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
AND3_X1 U856 ( .A1(KEYINPUT57), .A2(n1136), .A3(G125), .ZN(n1190) );
INV_X1 U857 ( .A(n1134), .ZN(n1136) );
NOR2_X1 U858 ( .A1(KEYINPUT57), .A2(n1191), .ZN(n1189) );
NOR2_X1 U859 ( .A1(n1086), .A2(G952), .ZN(n1105) );
NAND2_X1 U860 ( .A1(n1192), .A2(n1193), .ZN(G48) );
NAND2_X1 U861 ( .A1(G146), .A2(n1167), .ZN(n1193) );
XOR2_X1 U862 ( .A(KEYINPUT24), .B(n1194), .Z(n1192) );
NOR2_X1 U863 ( .A1(G146), .A2(n1167), .ZN(n1194) );
NAND3_X1 U864 ( .A1(n1184), .A2(n1034), .A3(n1161), .ZN(n1167) );
XNOR2_X1 U865 ( .A(G143), .B(n1168), .ZN(G45) );
NAND4_X1 U866 ( .A1(n1040), .A2(n1195), .A3(n1196), .A4(n1034), .ZN(n1168) );
XOR2_X1 U867 ( .A(n1148), .B(n1173), .Z(G42) );
NAND3_X1 U868 ( .A1(n1183), .A2(n1039), .A3(n1174), .ZN(n1173) );
INV_X1 U869 ( .A(n1197), .ZN(n1183) );
XNOR2_X1 U870 ( .A(G137), .B(n1198), .ZN(G39) );
NAND3_X1 U871 ( .A1(n1174), .A2(n1184), .A3(n1199), .ZN(n1198) );
XOR2_X1 U872 ( .A(n1028), .B(KEYINPUT50), .Z(n1199) );
INV_X1 U873 ( .A(n1185), .ZN(n1028) );
XNOR2_X1 U874 ( .A(G134), .B(n1200), .ZN(G36) );
NAND4_X1 U875 ( .A1(n1201), .A2(n1174), .A3(n1047), .A4(n1202), .ZN(n1200) );
XOR2_X1 U876 ( .A(KEYINPUT36), .B(n1181), .Z(n1202) );
INV_X1 U877 ( .A(n1203), .ZN(n1181) );
INV_X1 U878 ( .A(n1038), .ZN(n1174) );
XOR2_X1 U879 ( .A(G131), .B(n1204), .Z(G33) );
NOR4_X1 U880 ( .A1(KEYINPUT62), .A2(n1197), .A3(n1038), .A4(n1205), .ZN(n1204) );
NAND2_X1 U881 ( .A1(n1206), .A2(n1036), .ZN(n1038) );
NAND2_X1 U882 ( .A1(n1161), .A2(n1196), .ZN(n1197) );
XOR2_X1 U883 ( .A(n1207), .B(n1172), .Z(G30) );
NAND3_X1 U884 ( .A1(n1165), .A2(n1034), .A3(n1184), .ZN(n1172) );
AND3_X1 U885 ( .A1(n1208), .A2(n1060), .A3(n1196), .ZN(n1184) );
AND2_X1 U886 ( .A1(n1047), .A2(n1203), .ZN(n1196) );
XOR2_X1 U887 ( .A(n1159), .B(n1209), .Z(G3) );
NAND2_X1 U888 ( .A1(KEYINPUT8), .A2(G101), .ZN(n1209) );
NAND3_X1 U889 ( .A1(n1040), .A2(n1185), .A3(n1163), .ZN(n1159) );
XOR2_X1 U890 ( .A(n1210), .B(n1171), .Z(G27) );
NAND4_X1 U891 ( .A1(n1044), .A2(n1039), .A3(n1034), .A4(n1203), .ZN(n1171) );
NAND2_X1 U892 ( .A1(n1020), .A2(n1211), .ZN(n1203) );
NAND4_X1 U893 ( .A1(n1085), .A2(G902), .A3(n1212), .A4(n1074), .ZN(n1211) );
INV_X1 U894 ( .A(G900), .ZN(n1074) );
XNOR2_X1 U895 ( .A(G122), .B(n1154), .ZN(G24) );
NAND3_X1 U896 ( .A1(n1195), .A2(n1162), .A3(n1213), .ZN(n1154) );
INV_X1 U897 ( .A(n1032), .ZN(n1162) );
NAND2_X1 U898 ( .A1(n1214), .A2(n1215), .ZN(n1032) );
INV_X1 U899 ( .A(n1208), .ZN(n1215) );
AND2_X1 U900 ( .A1(n1216), .A2(n1217), .ZN(n1195) );
XOR2_X1 U901 ( .A(n1218), .B(KEYINPUT49), .Z(n1216) );
NAND2_X1 U902 ( .A1(n1219), .A2(n1220), .ZN(G21) );
NAND2_X1 U903 ( .A1(G119), .A2(n1155), .ZN(n1220) );
XOR2_X1 U904 ( .A(n1221), .B(KEYINPUT16), .Z(n1219) );
OR2_X1 U905 ( .A1(n1155), .A2(G119), .ZN(n1221) );
NAND4_X1 U906 ( .A1(n1208), .A2(n1213), .A3(n1185), .A4(n1060), .ZN(n1155) );
XNOR2_X1 U907 ( .A(G116), .B(n1156), .ZN(G18) );
NAND2_X1 U908 ( .A1(n1213), .A2(n1201), .ZN(n1156) );
INV_X1 U909 ( .A(n1182), .ZN(n1201) );
NAND2_X1 U910 ( .A1(n1040), .A2(n1165), .ZN(n1182) );
INV_X1 U911 ( .A(n1041), .ZN(n1165) );
NAND2_X1 U912 ( .A1(n1222), .A2(n1217), .ZN(n1041) );
AND3_X1 U913 ( .A1(n1034), .A2(n1166), .A3(n1223), .ZN(n1213) );
XOR2_X1 U914 ( .A(n1164), .B(KEYINPUT4), .Z(n1034) );
NAND2_X1 U915 ( .A1(n1224), .A2(n1225), .ZN(G15) );
OR2_X1 U916 ( .A1(n1157), .A2(G113), .ZN(n1225) );
XOR2_X1 U917 ( .A(n1226), .B(KEYINPUT56), .Z(n1224) );
NAND2_X1 U918 ( .A1(G113), .A2(n1157), .ZN(n1226) );
NAND4_X1 U919 ( .A1(n1040), .A2(n1044), .A3(n1164), .A4(n1166), .ZN(n1157) );
AND2_X1 U920 ( .A1(n1223), .A2(n1161), .ZN(n1044) );
NOR2_X1 U921 ( .A1(n1217), .A2(n1218), .ZN(n1161) );
XOR2_X1 U922 ( .A(n1222), .B(KEYINPUT53), .Z(n1218) );
INV_X1 U923 ( .A(n1024), .ZN(n1223) );
NAND2_X1 U924 ( .A1(n1062), .A2(n1049), .ZN(n1024) );
INV_X1 U925 ( .A(n1205), .ZN(n1040) );
NAND2_X1 U926 ( .A1(n1208), .A2(n1214), .ZN(n1205) );
XOR2_X1 U927 ( .A(n1227), .B(n1160), .Z(G12) );
NAND3_X1 U928 ( .A1(n1039), .A2(n1185), .A3(n1163), .ZN(n1160) );
AND3_X1 U929 ( .A1(n1047), .A2(n1166), .A3(n1164), .ZN(n1163) );
INV_X1 U930 ( .A(n1012), .ZN(n1164) );
NAND2_X1 U931 ( .A1(n1036), .A2(n1035), .ZN(n1012) );
INV_X1 U932 ( .A(n1206), .ZN(n1035) );
NOR2_X1 U933 ( .A1(n1054), .A2(n1228), .ZN(n1206) );
NOR2_X1 U934 ( .A1(n1058), .A2(n1056), .ZN(n1228) );
AND2_X1 U935 ( .A1(n1056), .A2(n1058), .ZN(n1054) );
NAND2_X1 U936 ( .A1(G210), .A2(n1229), .ZN(n1058) );
AND2_X1 U937 ( .A1(n1230), .A2(n1231), .ZN(n1056) );
XOR2_X1 U938 ( .A(n1187), .B(n1232), .Z(n1230) );
XOR2_X1 U939 ( .A(KEYINPUT18), .B(n1191), .Z(n1232) );
XOR2_X1 U940 ( .A(G125), .B(n1134), .Z(n1191) );
XOR2_X1 U941 ( .A(n1233), .B(n1234), .Z(n1187) );
XOR2_X1 U942 ( .A(KEYINPUT59), .B(n1235), .Z(n1234) );
AND2_X1 U943 ( .A1(n1086), .A2(G224), .ZN(n1235) );
XNOR2_X1 U944 ( .A(n1101), .B(n1102), .ZN(n1233) );
XNOR2_X1 U945 ( .A(n1236), .B(n1237), .ZN(n1102) );
XOR2_X1 U946 ( .A(n1238), .B(KEYINPUT6), .Z(n1236) );
XNOR2_X1 U947 ( .A(n1239), .B(n1240), .ZN(n1101) );
XOR2_X1 U948 ( .A(n1241), .B(n1242), .Z(n1239) );
NAND2_X1 U949 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
NAND2_X1 U950 ( .A1(n1245), .A2(n1227), .ZN(n1244) );
XOR2_X1 U951 ( .A(KEYINPUT29), .B(n1246), .Z(n1243) );
NOR2_X1 U952 ( .A1(n1245), .A2(n1227), .ZN(n1246) );
NAND2_X1 U953 ( .A1(G214), .A2(n1229), .ZN(n1036) );
NAND2_X1 U954 ( .A1(n1247), .A2(n1231), .ZN(n1229) );
INV_X1 U955 ( .A(G237), .ZN(n1247) );
NAND2_X1 U956 ( .A1(n1020), .A2(n1248), .ZN(n1166) );
NAND4_X1 U957 ( .A1(n1085), .A2(G902), .A3(n1212), .A4(n1099), .ZN(n1248) );
INV_X1 U958 ( .A(G898), .ZN(n1099) );
XOR2_X1 U959 ( .A(n1086), .B(KEYINPUT34), .Z(n1085) );
NAND3_X1 U960 ( .A1(n1212), .A2(n1086), .A3(G952), .ZN(n1020) );
NAND2_X1 U961 ( .A1(G237), .A2(G234), .ZN(n1212) );
NOR2_X1 U962 ( .A1(n1062), .A2(n1055), .ZN(n1047) );
INV_X1 U963 ( .A(n1049), .ZN(n1055) );
NAND2_X1 U964 ( .A1(G221), .A2(n1249), .ZN(n1049) );
NAND2_X1 U965 ( .A1(G234), .A2(n1231), .ZN(n1249) );
XOR2_X1 U966 ( .A(n1250), .B(G469), .Z(n1062) );
NAND2_X1 U967 ( .A1(n1251), .A2(n1231), .ZN(n1250) );
XOR2_X1 U968 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U969 ( .A(G140), .B(G110), .Z(n1253) );
XOR2_X1 U970 ( .A(n1146), .B(n1137), .Z(n1252) );
XOR2_X1 U971 ( .A(n1254), .B(n1255), .Z(n1146) );
XOR2_X1 U972 ( .A(n1256), .B(n1257), .Z(n1255) );
NAND2_X1 U973 ( .A1(KEYINPUT35), .A2(n1238), .ZN(n1257) );
INV_X1 U974 ( .A(G101), .ZN(n1238) );
NAND2_X1 U975 ( .A1(G227), .A2(n1086), .ZN(n1256) );
INV_X1 U976 ( .A(G953), .ZN(n1086) );
XNOR2_X1 U977 ( .A(n1237), .B(n1084), .ZN(n1254) );
XOR2_X1 U978 ( .A(n1258), .B(n1259), .Z(n1084) );
NOR2_X1 U979 ( .A1(G143), .A2(KEYINPUT30), .ZN(n1259) );
XOR2_X1 U980 ( .A(G104), .B(G107), .Z(n1237) );
NOR2_X1 U981 ( .A1(n1217), .A2(n1260), .ZN(n1185) );
INV_X1 U982 ( .A(n1222), .ZN(n1260) );
XOR2_X1 U983 ( .A(n1261), .B(G475), .Z(n1222) );
NAND2_X1 U984 ( .A1(n1262), .A2(n1117), .ZN(n1261) );
XNOR2_X1 U985 ( .A(n1263), .B(n1264), .ZN(n1117) );
XOR2_X1 U986 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U987 ( .A(n1267), .B(n1268), .Z(n1266) );
AND2_X1 U988 ( .A1(G214), .A2(n1269), .ZN(n1268) );
NAND4_X1 U989 ( .A1(n1270), .A2(n1271), .A3(n1272), .A4(n1273), .ZN(n1267) );
NAND3_X1 U990 ( .A1(n1082), .A2(n1274), .A3(KEYINPUT51), .ZN(n1273) );
INV_X1 U991 ( .A(KEYINPUT11), .ZN(n1274) );
OR2_X1 U992 ( .A1(n1210), .A2(KEYINPUT51), .ZN(n1272) );
INV_X1 U993 ( .A(G125), .ZN(n1210) );
NAND2_X1 U994 ( .A1(KEYINPUT11), .A2(G140), .ZN(n1270) );
XOR2_X1 U995 ( .A(n1275), .B(n1276), .Z(n1263) );
XOR2_X1 U996 ( .A(G146), .B(G131), .Z(n1276) );
XNOR2_X1 U997 ( .A(G104), .B(G113), .ZN(n1275) );
XOR2_X1 U998 ( .A(KEYINPUT54), .B(G902), .Z(n1262) );
XNOR2_X1 U999 ( .A(n1277), .B(G478), .ZN(n1217) );
OR2_X1 U1000 ( .A1(n1113), .A2(G902), .ZN(n1277) );
XNOR2_X1 U1001 ( .A(n1278), .B(n1279), .ZN(n1113) );
XOR2_X1 U1002 ( .A(G107), .B(n1280), .Z(n1279) );
XOR2_X1 U1003 ( .A(G128), .B(G116), .Z(n1280) );
XOR2_X1 U1004 ( .A(n1281), .B(n1282), .Z(n1278) );
XOR2_X1 U1005 ( .A(n1265), .B(n1283), .Z(n1281) );
AND2_X1 U1006 ( .A1(n1284), .A2(G217), .ZN(n1283) );
XNOR2_X1 U1007 ( .A(G143), .B(n1245), .ZN(n1265) );
XOR2_X1 U1008 ( .A(G122), .B(KEYINPUT10), .Z(n1245) );
NOR2_X1 U1009 ( .A1(n1208), .A2(n1214), .ZN(n1039) );
INV_X1 U1010 ( .A(n1060), .ZN(n1214) );
NAND2_X1 U1011 ( .A1(n1285), .A2(n1286), .ZN(n1060) );
NAND2_X1 U1012 ( .A1(G217), .A2(n1287), .ZN(n1286) );
NAND2_X1 U1013 ( .A1(n1231), .A2(n1288), .ZN(n1287) );
OR2_X1 U1014 ( .A1(n1289), .A2(G234), .ZN(n1288) );
NAND3_X1 U1015 ( .A1(n1290), .A2(n1231), .A3(n1289), .ZN(n1285) );
XNOR2_X1 U1016 ( .A(n1107), .B(KEYINPUT58), .ZN(n1289) );
XNOR2_X1 U1017 ( .A(n1291), .B(n1292), .ZN(n1107) );
XOR2_X1 U1018 ( .A(n1293), .B(n1294), .Z(n1292) );
XOR2_X1 U1019 ( .A(n1295), .B(n1296), .Z(n1294) );
NOR3_X1 U1020 ( .A1(n1081), .A2(n1297), .A3(n1298), .ZN(n1296) );
AND2_X1 U1021 ( .A1(n1082), .A2(KEYINPUT15), .ZN(n1298) );
NOR2_X1 U1022 ( .A1(G140), .A2(G125), .ZN(n1082) );
NOR2_X1 U1023 ( .A1(KEYINPUT15), .A2(n1148), .ZN(n1297) );
INV_X1 U1024 ( .A(G140), .ZN(n1148) );
INV_X1 U1025 ( .A(n1271), .ZN(n1081) );
NAND2_X1 U1026 ( .A1(G140), .A2(G125), .ZN(n1271) );
NAND2_X1 U1027 ( .A1(n1299), .A2(n1300), .ZN(n1295) );
XNOR2_X1 U1028 ( .A(G137), .B(n1301), .ZN(n1300) );
NAND2_X1 U1029 ( .A1(n1284), .A2(G221), .ZN(n1301) );
NOR2_X1 U1030 ( .A1(n1302), .A2(G953), .ZN(n1284) );
XNOR2_X1 U1031 ( .A(KEYINPUT42), .B(KEYINPUT23), .ZN(n1299) );
XOR2_X1 U1032 ( .A(n1227), .B(n1303), .Z(n1291) );
XOR2_X1 U1033 ( .A(KEYINPUT0), .B(G119), .Z(n1303) );
NAND2_X1 U1034 ( .A1(G217), .A2(n1302), .ZN(n1290) );
INV_X1 U1035 ( .A(G234), .ZN(n1302) );
XOR2_X1 U1036 ( .A(n1065), .B(n1304), .Z(n1208) );
NOR2_X1 U1037 ( .A1(n1064), .A2(KEYINPUT61), .ZN(n1304) );
AND2_X1 U1038 ( .A1(n1305), .A2(n1231), .ZN(n1064) );
INV_X1 U1039 ( .A(G902), .ZN(n1231) );
XOR2_X1 U1040 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1041 ( .A(n1308), .B(n1309), .Z(n1307) );
NOR2_X1 U1042 ( .A1(KEYINPUT20), .A2(n1129), .ZN(n1309) );
XNOR2_X1 U1043 ( .A(n1310), .B(n1242), .ZN(n1129) );
XOR2_X1 U1044 ( .A(G113), .B(KEYINPUT17), .Z(n1242) );
NAND2_X1 U1045 ( .A1(KEYINPUT45), .A2(n1240), .ZN(n1310) );
XOR2_X1 U1046 ( .A(G116), .B(G119), .Z(n1240) );
NOR3_X1 U1047 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1308) );
NOR2_X1 U1048 ( .A1(n1314), .A2(n1137), .ZN(n1313) );
AND3_X1 U1049 ( .A1(n1137), .A2(n1314), .A3(KEYINPUT52), .ZN(n1312) );
AND2_X1 U1050 ( .A1(KEYINPUT7), .A2(n1315), .ZN(n1314) );
INV_X1 U1051 ( .A(n1133), .ZN(n1137) );
XOR2_X1 U1052 ( .A(n1316), .B(n1317), .Z(n1133) );
INV_X1 U1053 ( .A(n1083), .ZN(n1317) );
XNOR2_X1 U1054 ( .A(G137), .B(n1282), .ZN(n1083) );
XOR2_X1 U1055 ( .A(G134), .B(KEYINPUT5), .Z(n1282) );
XOR2_X1 U1056 ( .A(n1079), .B(KEYINPUT43), .Z(n1316) );
INV_X1 U1057 ( .A(G131), .ZN(n1079) );
NOR2_X1 U1058 ( .A1(KEYINPUT52), .A2(n1315), .ZN(n1311) );
XOR2_X1 U1059 ( .A(n1134), .B(KEYINPUT46), .Z(n1315) );
XOR2_X1 U1060 ( .A(G143), .B(n1258), .Z(n1134) );
INV_X1 U1061 ( .A(n1293), .ZN(n1258) );
XOR2_X1 U1062 ( .A(n1207), .B(G146), .Z(n1293) );
INV_X1 U1063 ( .A(G128), .ZN(n1207) );
NOR2_X1 U1064 ( .A1(n1318), .A2(n1319), .ZN(n1306) );
NOR2_X1 U1065 ( .A1(KEYINPUT14), .A2(n1320), .ZN(n1319) );
INV_X1 U1066 ( .A(n1122), .ZN(n1320) );
NOR2_X1 U1067 ( .A1(KEYINPUT28), .A2(n1122), .ZN(n1318) );
XOR2_X1 U1068 ( .A(n1321), .B(G101), .Z(n1122) );
NAND2_X1 U1069 ( .A1(n1269), .A2(G210), .ZN(n1321) );
NOR2_X1 U1070 ( .A1(G953), .A2(G237), .ZN(n1269) );
INV_X1 U1071 ( .A(G472), .ZN(n1065) );
INV_X1 U1072 ( .A(G110), .ZN(n1227) );
endmodule


