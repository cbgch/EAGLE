//Key = 1110111110011000111000000011110110000010010000000101110001111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;

XNOR2_X1 U733 ( .A(G107), .B(n1018), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1021), .A2(n1022), .A3(G953), .A4(n1023), .ZN(n1020) );
NOR3_X1 U736 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1022) );
NOR2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR3_X1 U738 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1027) );
INV_X1 U739 ( .A(KEYINPUT62), .ZN(n1029) );
NAND3_X1 U740 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1021) );
NAND2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NAND3_X1 U742 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
XOR2_X1 U743 ( .A(KEYINPUT58), .B(n1040), .Z(n1039) );
NOR2_X1 U744 ( .A1(n1041), .A2(n1024), .ZN(n1040) );
NAND3_X1 U745 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1038) );
NAND2_X1 U746 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
OR2_X1 U747 ( .A1(n1047), .A2(KEYINPUT6), .ZN(n1045) );
NAND4_X1 U748 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1042) );
NAND2_X1 U749 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NAND3_X1 U750 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND2_X1 U751 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U752 ( .A1(KEYINPUT62), .A2(n1059), .ZN(n1058) );
NAND4_X1 U753 ( .A1(n1060), .A2(n1061), .A3(n1057), .A4(n1059), .ZN(n1049) );
INV_X1 U754 ( .A(KEYINPUT13), .ZN(n1059) );
NAND2_X1 U755 ( .A1(KEYINPUT6), .A2(n1062), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1063), .A2(n1064), .ZN(n1037) );
INV_X1 U757 ( .A(n1024), .ZN(n1063) );
NAND3_X1 U758 ( .A1(n1052), .A2(n1057), .A3(n1051), .ZN(n1024) );
INV_X1 U759 ( .A(n1046), .ZN(n1051) );
NOR3_X1 U760 ( .A1(n1023), .A2(G953), .A3(G952), .ZN(n1019) );
AND4_X1 U761 ( .A1(n1065), .A2(n1052), .A3(n1066), .A4(n1067), .ZN(n1023) );
NOR4_X1 U762 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1067) );
NOR2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
NOR2_X1 U764 ( .A1(G902), .A2(n1074), .ZN(n1072) );
XOR2_X1 U765 ( .A(n1075), .B(G472), .Z(n1066) );
XNOR2_X1 U766 ( .A(n1076), .B(n1077), .ZN(n1065) );
NAND2_X1 U767 ( .A1(KEYINPUT57), .A2(n1078), .ZN(n1076) );
XOR2_X1 U768 ( .A(n1079), .B(n1080), .Z(G72) );
NOR2_X1 U769 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U770 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
XOR2_X1 U771 ( .A(n1085), .B(n1086), .Z(n1079) );
NOR2_X1 U772 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U773 ( .A(n1089), .B(n1090), .Z(n1088) );
XOR2_X1 U774 ( .A(n1091), .B(n1092), .Z(n1090) );
XNOR2_X1 U775 ( .A(n1093), .B(n1094), .ZN(n1092) );
NAND2_X1 U776 ( .A1(KEYINPUT53), .A2(n1095), .ZN(n1091) );
XNOR2_X1 U777 ( .A(KEYINPUT61), .B(n1096), .ZN(n1095) );
XOR2_X1 U778 ( .A(n1097), .B(n1098), .Z(n1089) );
XOR2_X1 U779 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U780 ( .A1(KEYINPUT30), .A2(n1101), .ZN(n1099) );
NOR2_X1 U781 ( .A1(G900), .A2(n1082), .ZN(n1087) );
NAND2_X1 U782 ( .A1(KEYINPUT0), .A2(n1102), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1103), .A2(n1082), .ZN(n1102) );
NAND2_X1 U784 ( .A1(n1104), .A2(n1105), .ZN(G69) );
NAND2_X1 U785 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U786 ( .A1(G953), .A2(n1108), .ZN(n1107) );
NAND3_X1 U787 ( .A1(G953), .A2(n1109), .A3(n1110), .ZN(n1104) );
XNOR2_X1 U788 ( .A(n1106), .B(KEYINPUT55), .ZN(n1110) );
XNOR2_X1 U789 ( .A(n1111), .B(n1112), .ZN(n1106) );
NOR2_X1 U790 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U791 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U792 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U793 ( .A1(KEYINPUT44), .A2(n1119), .ZN(n1118) );
NAND3_X1 U794 ( .A1(n1120), .A2(n1082), .A3(KEYINPUT16), .ZN(n1111) );
NAND2_X1 U795 ( .A1(G898), .A2(G224), .ZN(n1109) );
NOR3_X1 U796 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(G66) );
NOR3_X1 U797 ( .A1(n1124), .A2(G953), .A3(n1125), .ZN(n1123) );
AND2_X1 U798 ( .A1(n1124), .A2(n1126), .ZN(n1122) );
INV_X1 U799 ( .A(KEYINPUT24), .ZN(n1124) );
XNOR2_X1 U800 ( .A(n1127), .B(n1128), .ZN(n1121) );
NOR2_X1 U801 ( .A1(n1073), .A2(n1129), .ZN(n1128) );
NOR2_X1 U802 ( .A1(n1126), .A2(n1130), .ZN(G63) );
NOR3_X1 U803 ( .A1(n1078), .A2(n1131), .A3(n1132), .ZN(n1130) );
NOR3_X1 U804 ( .A1(n1133), .A2(n1077), .A3(n1129), .ZN(n1132) );
NOR2_X1 U805 ( .A1(n1134), .A2(n1135), .ZN(n1131) );
NOR2_X1 U806 ( .A1(n1136), .A2(n1077), .ZN(n1134) );
NOR2_X1 U807 ( .A1(n1103), .A2(n1120), .ZN(n1136) );
NOR2_X1 U808 ( .A1(n1126), .A2(n1137), .ZN(G60) );
XOR2_X1 U809 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U810 ( .A1(n1140), .A2(n1129), .ZN(n1138) );
XOR2_X1 U811 ( .A(n1141), .B(n1142), .Z(G6) );
NOR4_X1 U812 ( .A1(n1143), .A2(n1144), .A3(n1041), .A4(n1145), .ZN(n1142) );
XOR2_X1 U813 ( .A(KEYINPUT49), .B(n1146), .Z(n1145) );
NAND2_X1 U814 ( .A1(KEYINPUT17), .A2(n1147), .ZN(n1141) );
NOR2_X1 U815 ( .A1(n1126), .A2(n1148), .ZN(G57) );
XOR2_X1 U816 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U817 ( .A1(n1129), .A2(n1151), .ZN(n1149) );
XOR2_X1 U818 ( .A(KEYINPUT38), .B(G472), .Z(n1151) );
NOR2_X1 U819 ( .A1(n1126), .A2(n1152), .ZN(G54) );
XOR2_X1 U820 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U821 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U822 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U823 ( .A1(n1159), .A2(n1129), .ZN(n1158) );
NOR2_X1 U824 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NOR2_X1 U825 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U826 ( .A(KEYINPUT37), .B(n1164), .Z(n1153) );
XOR2_X1 U827 ( .A(KEYINPUT54), .B(KEYINPUT40), .Z(n1164) );
NOR2_X1 U828 ( .A1(n1126), .A2(n1165), .ZN(G51) );
XOR2_X1 U829 ( .A(n1166), .B(n1167), .Z(n1165) );
XNOR2_X1 U830 ( .A(n1168), .B(n1169), .ZN(n1167) );
XOR2_X1 U831 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U832 ( .A(n1172), .B(n1173), .Z(n1166) );
XOR2_X1 U833 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U834 ( .A1(n1176), .A2(n1129), .ZN(n1175) );
NAND2_X1 U835 ( .A1(G902), .A2(n1177), .ZN(n1129) );
NAND2_X1 U836 ( .A1(n1034), .A2(n1032), .ZN(n1177) );
INV_X1 U837 ( .A(n1103), .ZN(n1032) );
NAND4_X1 U838 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1103) );
AND4_X1 U839 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
NOR2_X1 U840 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
NOR2_X1 U841 ( .A1(n1041), .A2(n1188), .ZN(n1187) );
NOR3_X1 U842 ( .A1(n1189), .A2(n1070), .A3(n1026), .ZN(n1186) );
INV_X1 U843 ( .A(n1120), .ZN(n1034) );
NAND2_X1 U844 ( .A1(n1190), .A2(n1191), .ZN(n1120) );
AND4_X1 U845 ( .A1(n1018), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1191) );
NAND3_X1 U846 ( .A1(n1062), .A2(n1195), .A3(n1064), .ZN(n1018) );
INV_X1 U847 ( .A(n1047), .ZN(n1062) );
NOR4_X1 U848 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1190) );
NOR3_X1 U849 ( .A1(n1041), .A2(n1144), .A3(n1047), .ZN(n1199) );
NAND2_X1 U850 ( .A1(n1146), .A2(n1057), .ZN(n1047) );
NOR2_X1 U851 ( .A1(G125), .A2(KEYINPUT35), .ZN(n1172) );
NOR2_X1 U852 ( .A1(n1082), .A2(n1125), .ZN(n1126) );
XNOR2_X1 U853 ( .A(G952), .B(KEYINPUT7), .ZN(n1125) );
XNOR2_X1 U854 ( .A(G146), .B(n1178), .ZN(G48) );
NAND3_X1 U855 ( .A1(n1200), .A2(n1028), .A3(n1201), .ZN(n1178) );
XNOR2_X1 U856 ( .A(G143), .B(n1179), .ZN(G45) );
NAND4_X1 U857 ( .A1(n1028), .A2(n1146), .A3(n1202), .A4(n1203), .ZN(n1179) );
AND3_X1 U858 ( .A1(n1071), .A2(n1204), .A3(n1205), .ZN(n1203) );
XNOR2_X1 U859 ( .A(G140), .B(n1185), .ZN(G42) );
NAND3_X1 U860 ( .A1(n1200), .A2(n1206), .A3(n1207), .ZN(n1185) );
XNOR2_X1 U861 ( .A(n1096), .B(n1208), .ZN(G39) );
NOR3_X1 U862 ( .A1(n1209), .A2(n1026), .A3(n1189), .ZN(n1208) );
INV_X1 U863 ( .A(n1044), .ZN(n1026) );
XNOR2_X1 U864 ( .A(KEYINPUT4), .B(n1070), .ZN(n1209) );
XNOR2_X1 U865 ( .A(G134), .B(n1184), .ZN(G36) );
NAND3_X1 U866 ( .A1(n1202), .A2(n1064), .A3(n1207), .ZN(n1184) );
XNOR2_X1 U867 ( .A(G131), .B(n1183), .ZN(G33) );
NAND3_X1 U868 ( .A1(n1200), .A2(n1202), .A3(n1207), .ZN(n1183) );
AND3_X1 U869 ( .A1(n1146), .A2(n1205), .A3(n1035), .ZN(n1207) );
INV_X1 U870 ( .A(n1070), .ZN(n1035) );
NAND2_X1 U871 ( .A1(n1210), .A2(n1030), .ZN(n1070) );
INV_X1 U872 ( .A(n1031), .ZN(n1210) );
XNOR2_X1 U873 ( .A(G128), .B(n1182), .ZN(G30) );
NAND3_X1 U874 ( .A1(n1064), .A2(n1028), .A3(n1201), .ZN(n1182) );
INV_X1 U875 ( .A(n1189), .ZN(n1201) );
NAND4_X1 U876 ( .A1(n1211), .A2(n1146), .A3(n1205), .A4(n1212), .ZN(n1189) );
NAND2_X1 U877 ( .A1(n1213), .A2(n1214), .ZN(G3) );
NAND2_X1 U878 ( .A1(n1198), .A2(n1215), .ZN(n1214) );
XOR2_X1 U879 ( .A(KEYINPUT5), .B(n1216), .Z(n1213) );
NOR2_X1 U880 ( .A1(n1198), .A2(n1215), .ZN(n1216) );
AND2_X1 U881 ( .A1(n1202), .A2(n1217), .ZN(n1198) );
XNOR2_X1 U882 ( .A(n1218), .B(n1219), .ZN(G27) );
NOR2_X1 U883 ( .A1(n1188), .A2(n1220), .ZN(n1219) );
XNOR2_X1 U884 ( .A(KEYINPUT8), .B(n1041), .ZN(n1220) );
INV_X1 U885 ( .A(n1200), .ZN(n1041) );
NAND4_X1 U886 ( .A1(n1206), .A2(n1052), .A3(n1028), .A4(n1205), .ZN(n1188) );
NAND2_X1 U887 ( .A1(n1046), .A2(n1221), .ZN(n1205) );
NAND4_X1 U888 ( .A1(G902), .A2(G953), .A3(n1222), .A4(n1084), .ZN(n1221) );
INV_X1 U889 ( .A(G900), .ZN(n1084) );
NAND2_X1 U890 ( .A1(n1223), .A2(n1224), .ZN(G24) );
NAND2_X1 U891 ( .A1(G122), .A2(n1225), .ZN(n1224) );
XOR2_X1 U892 ( .A(n1226), .B(KEYINPUT50), .Z(n1223) );
NAND2_X1 U893 ( .A1(n1197), .A2(n1227), .ZN(n1226) );
INV_X1 U894 ( .A(n1225), .ZN(n1197) );
NAND4_X1 U895 ( .A1(n1228), .A2(n1057), .A3(n1071), .A4(n1204), .ZN(n1225) );
INV_X1 U896 ( .A(n1143), .ZN(n1057) );
NAND2_X1 U897 ( .A1(n1229), .A2(n1230), .ZN(n1143) );
XOR2_X1 U898 ( .A(G119), .B(n1196), .Z(G21) );
AND4_X1 U899 ( .A1(n1211), .A2(n1228), .A3(n1044), .A4(n1212), .ZN(n1196) );
XNOR2_X1 U900 ( .A(G116), .B(n1194), .ZN(G18) );
NAND3_X1 U901 ( .A1(n1228), .A2(n1064), .A3(n1202), .ZN(n1194) );
AND2_X1 U902 ( .A1(n1231), .A2(n1204), .ZN(n1064) );
XOR2_X1 U903 ( .A(KEYINPUT45), .B(n1232), .Z(n1231) );
XOR2_X1 U904 ( .A(n1193), .B(n1233), .Z(G15) );
NAND2_X1 U905 ( .A1(KEYINPUT26), .A2(G113), .ZN(n1233) );
NAND3_X1 U906 ( .A1(n1202), .A2(n1228), .A3(n1200), .ZN(n1193) );
NOR2_X1 U907 ( .A1(n1204), .A2(n1232), .ZN(n1200) );
INV_X1 U908 ( .A(n1071), .ZN(n1232) );
AND2_X1 U909 ( .A1(n1052), .A2(n1195), .ZN(n1228) );
NOR2_X1 U910 ( .A1(n1234), .A2(n1061), .ZN(n1052) );
INV_X1 U911 ( .A(n1054), .ZN(n1202) );
NAND2_X1 U912 ( .A1(n1211), .A2(n1229), .ZN(n1054) );
XOR2_X1 U913 ( .A(n1212), .B(KEYINPUT2), .Z(n1229) );
INV_X1 U914 ( .A(n1230), .ZN(n1211) );
NAND2_X1 U915 ( .A1(n1235), .A2(n1236), .ZN(G12) );
NAND2_X1 U916 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U917 ( .A(KEYINPUT47), .B(n1192), .ZN(n1237) );
NAND2_X1 U918 ( .A1(G110), .A2(n1239), .ZN(n1235) );
XOR2_X1 U919 ( .A(n1192), .B(KEYINPUT10), .Z(n1239) );
NAND2_X1 U920 ( .A1(n1206), .A2(n1217), .ZN(n1192) );
AND3_X1 U921 ( .A1(n1195), .A2(n1146), .A3(n1044), .ZN(n1217) );
NOR2_X1 U922 ( .A1(n1240), .A2(n1204), .ZN(n1044) );
NAND3_X1 U923 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1204) );
OR2_X1 U924 ( .A1(n1077), .A2(KEYINPUT1), .ZN(n1243) );
NAND3_X1 U925 ( .A1(KEYINPUT1), .A2(n1077), .A3(n1078), .ZN(n1242) );
NAND2_X1 U926 ( .A1(n1244), .A2(n1245), .ZN(n1241) );
INV_X1 U927 ( .A(n1078), .ZN(n1245) );
NOR2_X1 U928 ( .A1(n1135), .A2(G902), .ZN(n1078) );
INV_X1 U929 ( .A(n1133), .ZN(n1135) );
XNOR2_X1 U930 ( .A(n1246), .B(n1247), .ZN(n1133) );
XOR2_X1 U931 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U932 ( .A(n1094), .B(G128), .ZN(n1249) );
XNOR2_X1 U933 ( .A(KEYINPUT14), .B(n1250), .ZN(n1248) );
XOR2_X1 U934 ( .A(n1251), .B(n1252), .Z(n1246) );
XNOR2_X1 U935 ( .A(n1227), .B(G116), .ZN(n1252) );
INV_X1 U936 ( .A(G122), .ZN(n1227) );
XNOR2_X1 U937 ( .A(n1253), .B(n1254), .ZN(n1251) );
INV_X1 U938 ( .A(G107), .ZN(n1254) );
NAND2_X1 U939 ( .A1(G217), .A2(n1255), .ZN(n1253) );
NAND2_X1 U940 ( .A1(KEYINPUT1), .A2(n1256), .ZN(n1244) );
XNOR2_X1 U941 ( .A(KEYINPUT28), .B(n1077), .ZN(n1256) );
INV_X1 U942 ( .A(G478), .ZN(n1077) );
XOR2_X1 U943 ( .A(KEYINPUT45), .B(n1071), .Z(n1240) );
XOR2_X1 U944 ( .A(n1257), .B(n1140), .Z(n1071) );
INV_X1 U945 ( .A(G475), .ZN(n1140) );
OR2_X1 U946 ( .A1(n1139), .A2(G902), .ZN(n1257) );
XNOR2_X1 U947 ( .A(n1258), .B(n1259), .ZN(n1139) );
XOR2_X1 U948 ( .A(n1097), .B(n1260), .Z(n1259) );
NAND2_X1 U949 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
OR2_X1 U950 ( .A1(n1263), .A2(G104), .ZN(n1262) );
NAND2_X1 U951 ( .A1(n1264), .A2(n1263), .ZN(n1261) );
XOR2_X1 U952 ( .A(n1265), .B(n1266), .Z(n1263) );
NOR2_X1 U953 ( .A1(KEYINPUT34), .A2(G122), .ZN(n1266) );
XNOR2_X1 U954 ( .A(G113), .B(KEYINPUT42), .ZN(n1265) );
XNOR2_X1 U955 ( .A(G104), .B(KEYINPUT27), .ZN(n1264) );
XNOR2_X1 U956 ( .A(G125), .B(G140), .ZN(n1097) );
XNOR2_X1 U957 ( .A(n1267), .B(n1268), .ZN(n1258) );
XNOR2_X1 U958 ( .A(n1269), .B(n1101), .ZN(n1267) );
NAND2_X1 U959 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND4_X1 U960 ( .A1(n1272), .A2(G214), .A3(n1273), .A4(n1082), .ZN(n1271) );
XNOR2_X1 U961 ( .A(G143), .B(KEYINPUT59), .ZN(n1272) );
XOR2_X1 U962 ( .A(n1274), .B(KEYINPUT36), .Z(n1270) );
NAND2_X1 U963 ( .A1(n1250), .A2(n1275), .ZN(n1274) );
NAND3_X1 U964 ( .A1(n1273), .A2(n1082), .A3(G214), .ZN(n1275) );
NOR2_X1 U965 ( .A1(n1060), .A2(n1061), .ZN(n1146) );
AND2_X1 U966 ( .A1(G221), .A2(n1276), .ZN(n1061) );
XNOR2_X1 U967 ( .A(KEYINPUT29), .B(n1277), .ZN(n1276) );
INV_X1 U968 ( .A(n1234), .ZN(n1060) );
XOR2_X1 U969 ( .A(n1278), .B(n1159), .Z(n1234) );
INV_X1 U970 ( .A(G469), .ZN(n1159) );
NAND2_X1 U971 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U972 ( .A(n1155), .B(n1281), .ZN(n1279) );
NOR3_X1 U973 ( .A1(n1160), .A2(n1282), .A3(n1283), .ZN(n1281) );
NOR3_X1 U974 ( .A1(n1163), .A2(KEYINPUT43), .A3(n1162), .ZN(n1283) );
AND2_X1 U975 ( .A1(n1163), .A2(KEYINPUT43), .ZN(n1282) );
AND2_X1 U976 ( .A1(n1162), .A2(n1163), .ZN(n1160) );
XNOR2_X1 U977 ( .A(G140), .B(n1284), .ZN(n1163) );
NOR2_X1 U978 ( .A1(n1083), .A2(G953), .ZN(n1162) );
INV_X1 U979 ( .A(G227), .ZN(n1083) );
XNOR2_X1 U980 ( .A(n1285), .B(n1286), .ZN(n1155) );
XOR2_X1 U981 ( .A(n1287), .B(n1288), .Z(n1286) );
NAND2_X1 U982 ( .A1(KEYINPUT60), .A2(n1289), .ZN(n1287) );
XOR2_X1 U983 ( .A(n1093), .B(KEYINPUT3), .Z(n1285) );
NAND2_X1 U984 ( .A1(KEYINPUT32), .A2(n1250), .ZN(n1093) );
INV_X1 U985 ( .A(n1144), .ZN(n1195) );
NAND2_X1 U986 ( .A1(n1028), .A2(n1290), .ZN(n1144) );
NAND2_X1 U987 ( .A1(n1291), .A2(n1046), .ZN(n1290) );
NAND3_X1 U988 ( .A1(n1222), .A2(n1082), .A3(G952), .ZN(n1046) );
NAND3_X1 U989 ( .A1(G902), .A2(n1113), .A3(n1292), .ZN(n1291) );
XOR2_X1 U990 ( .A(n1222), .B(KEYINPUT15), .Z(n1292) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1222) );
NOR2_X1 U992 ( .A1(n1082), .A2(G898), .ZN(n1113) );
AND2_X1 U993 ( .A1(n1031), .A2(n1030), .ZN(n1028) );
NAND2_X1 U994 ( .A1(G214), .A2(n1293), .ZN(n1030) );
XOR2_X1 U995 ( .A(n1294), .B(n1176), .Z(n1031) );
NAND2_X1 U996 ( .A1(G210), .A2(n1293), .ZN(n1176) );
NAND2_X1 U997 ( .A1(n1273), .A2(n1280), .ZN(n1293) );
NAND3_X1 U998 ( .A1(n1295), .A2(n1280), .A3(n1296), .ZN(n1294) );
XOR2_X1 U999 ( .A(n1297), .B(KEYINPUT56), .Z(n1296) );
OR2_X1 U1000 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U1001 ( .A1(n1299), .A2(n1298), .ZN(n1295) );
XOR2_X1 U1002 ( .A(n1119), .B(n1171), .Z(n1298) );
XOR2_X1 U1003 ( .A(n1300), .B(n1117), .Z(n1171) );
NAND2_X1 U1004 ( .A1(n1301), .A2(n1302), .ZN(n1117) );
OR2_X1 U1005 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XOR2_X1 U1006 ( .A(n1305), .B(KEYINPUT9), .Z(n1301) );
NAND2_X1 U1007 ( .A1(n1304), .A2(n1303), .ZN(n1305) );
INV_X1 U1008 ( .A(n1306), .ZN(n1303) );
XOR2_X1 U1009 ( .A(G113), .B(KEYINPUT46), .Z(n1304) );
XNOR2_X1 U1010 ( .A(KEYINPUT12), .B(n1307), .ZN(n1300) );
NOR2_X1 U1011 ( .A1(KEYINPUT33), .A2(n1115), .ZN(n1307) );
XNOR2_X1 U1012 ( .A(G122), .B(n1284), .ZN(n1115) );
XNOR2_X1 U1013 ( .A(n1174), .B(n1215), .ZN(n1119) );
INV_X1 U1014 ( .A(G101), .ZN(n1215) );
NOR2_X1 U1015 ( .A1(n1308), .A2(n1289), .ZN(n1174) );
XNOR2_X1 U1016 ( .A(G107), .B(n1147), .ZN(n1289) );
INV_X1 U1017 ( .A(G104), .ZN(n1147) );
INV_X1 U1018 ( .A(KEYINPUT41), .ZN(n1308) );
XNOR2_X1 U1019 ( .A(n1309), .B(n1310), .ZN(n1299) );
XNOR2_X1 U1020 ( .A(n1100), .B(n1170), .ZN(n1310) );
XNOR2_X1 U1021 ( .A(G143), .B(n1311), .ZN(n1170) );
NOR2_X1 U1022 ( .A1(G953), .A2(n1108), .ZN(n1311) );
INV_X1 U1023 ( .A(G224), .ZN(n1108) );
XNOR2_X1 U1024 ( .A(G125), .B(KEYINPUT20), .ZN(n1309) );
INV_X1 U1025 ( .A(n1055), .ZN(n1206) );
NAND2_X1 U1026 ( .A1(n1230), .A2(n1212), .ZN(n1055) );
NAND2_X1 U1027 ( .A1(n1312), .A2(n1313), .ZN(n1212) );
NAND2_X1 U1028 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND3_X1 U1029 ( .A1(n1280), .A2(n1316), .A3(n1127), .ZN(n1315) );
NAND2_X1 U1030 ( .A1(n1068), .A2(n1316), .ZN(n1312) );
INV_X1 U1031 ( .A(KEYINPUT19), .ZN(n1316) );
NOR3_X1 U1032 ( .A1(n1314), .A2(G902), .A3(n1074), .ZN(n1068) );
INV_X1 U1033 ( .A(n1127), .ZN(n1074) );
XNOR2_X1 U1034 ( .A(n1317), .B(n1318), .ZN(n1127) );
XNOR2_X1 U1035 ( .A(G137), .B(n1319), .ZN(n1318) );
NAND2_X1 U1036 ( .A1(n1320), .A2(KEYINPUT18), .ZN(n1319) );
XOR2_X1 U1037 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1038 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR2_X1 U1039 ( .A1(KEYINPUT48), .A2(n1218), .ZN(n1324) );
INV_X1 U1040 ( .A(G125), .ZN(n1218) );
NOR2_X1 U1041 ( .A1(KEYINPUT21), .A2(n1268), .ZN(n1323) );
XNOR2_X1 U1042 ( .A(G146), .B(KEYINPUT51), .ZN(n1268) );
XOR2_X1 U1043 ( .A(n1325), .B(G140), .Z(n1321) );
NAND2_X1 U1044 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND2_X1 U1045 ( .A1(n1328), .A2(n1284), .ZN(n1327) );
XOR2_X1 U1046 ( .A(KEYINPUT11), .B(n1329), .Z(n1326) );
NOR2_X1 U1047 ( .A1(n1284), .A2(n1328), .ZN(n1329) );
XOR2_X1 U1048 ( .A(G128), .B(G119), .Z(n1328) );
XNOR2_X1 U1049 ( .A(n1238), .B(KEYINPUT63), .ZN(n1284) );
INV_X1 U1050 ( .A(G110), .ZN(n1238) );
NAND2_X1 U1051 ( .A1(G221), .A2(n1255), .ZN(n1317) );
AND2_X1 U1052 ( .A1(G234), .A2(n1082), .ZN(n1255) );
INV_X1 U1053 ( .A(n1073), .ZN(n1314) );
NAND2_X1 U1054 ( .A1(G217), .A2(n1277), .ZN(n1073) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1280), .ZN(n1277) );
XNOR2_X1 U1056 ( .A(n1075), .B(n1330), .ZN(n1230) );
NOR2_X1 U1057 ( .A1(G472), .A2(KEYINPUT22), .ZN(n1330) );
NAND2_X1 U1058 ( .A1(n1331), .A2(n1280), .ZN(n1075) );
INV_X1 U1059 ( .A(G902), .ZN(n1280) );
XOR2_X1 U1060 ( .A(KEYINPUT31), .B(n1150), .Z(n1331) );
XNOR2_X1 U1061 ( .A(n1332), .B(n1333), .ZN(n1150) );
XOR2_X1 U1062 ( .A(n1288), .B(n1334), .Z(n1333) );
XOR2_X1 U1063 ( .A(n1335), .B(n1336), .Z(n1334) );
NOR2_X1 U1064 ( .A1(KEYINPUT39), .A2(n1306), .ZN(n1336) );
XNOR2_X1 U1065 ( .A(G116), .B(G119), .ZN(n1306) );
NAND3_X1 U1066 ( .A1(n1273), .A2(n1082), .A3(G210), .ZN(n1335) );
INV_X1 U1067 ( .A(G953), .ZN(n1082) );
INV_X1 U1068 ( .A(G237), .ZN(n1273) );
XOR2_X1 U1069 ( .A(n1337), .B(n1168), .Z(n1288) );
XOR2_X1 U1070 ( .A(G101), .B(n1100), .Z(n1168) );
XOR2_X1 U1071 ( .A(G146), .B(G128), .Z(n1100) );
XNOR2_X1 U1072 ( .A(n1338), .B(n1101), .ZN(n1337) );
INV_X1 U1073 ( .A(G131), .ZN(n1101) );
NAND3_X1 U1074 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1338) );
NAND2_X1 U1075 ( .A1(KEYINPUT25), .A2(G134), .ZN(n1341) );
NAND3_X1 U1076 ( .A1(n1094), .A2(n1342), .A3(G137), .ZN(n1340) );
NAND2_X1 U1077 ( .A1(n1343), .A2(n1096), .ZN(n1339) );
INV_X1 U1078 ( .A(G137), .ZN(n1096) );
NAND2_X1 U1079 ( .A1(n1344), .A2(n1342), .ZN(n1343) );
INV_X1 U1080 ( .A(KEYINPUT25), .ZN(n1342) );
XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(n1094), .ZN(n1344) );
INV_X1 U1082 ( .A(G134), .ZN(n1094) );
XNOR2_X1 U1083 ( .A(G113), .B(n1345), .ZN(n1332) );
XNOR2_X1 U1084 ( .A(KEYINPUT23), .B(n1250), .ZN(n1345) );
INV_X1 U1085 ( .A(G143), .ZN(n1250) );
endmodule


