//Key = 1011001100101111110001001111001101111110000101001011011101110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;

XNOR2_X1 U736 ( .A(n1015), .B(n1016), .ZN(G9) );
NOR2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1019), .A2(n1020), .A3(G953), .A4(n1021), .ZN(n1018) );
NOR3_X1 U739 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1020) );
NAND3_X1 U740 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1022) );
NAND2_X1 U741 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND3_X1 U742 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1028) );
INV_X1 U743 ( .A(KEYINPUT16), .ZN(n1031) );
NAND3_X1 U744 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1025) );
NAND2_X1 U745 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NAND2_X1 U746 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U747 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U748 ( .A1(n1030), .A2(n1042), .ZN(n1033) );
NAND2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U750 ( .A1(KEYINPUT16), .A2(n1032), .ZN(n1044) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1019) );
NAND4_X1 U752 ( .A1(n1035), .A2(n1036), .A3(n1030), .A4(n1047), .ZN(n1046) );
NAND2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U754 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
NAND2_X1 U755 ( .A1(n1023), .A2(n1053), .ZN(n1051) );
NAND3_X1 U756 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
NAND2_X1 U758 ( .A1(n1059), .A2(n1027), .ZN(n1048) );
INV_X1 U759 ( .A(n1029), .ZN(n1035) );
NOR3_X1 U760 ( .A1(n1021), .A2(G953), .A3(G952), .ZN(n1017) );
AND4_X1 U761 ( .A1(n1052), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1021) );
NOR4_X1 U762 ( .A1(n1063), .A2(n1040), .A3(n1064), .A4(n1065), .ZN(n1062) );
XNOR2_X1 U763 ( .A(n1066), .B(n1067), .ZN(n1065) );
NAND2_X1 U764 ( .A1(KEYINPUT58), .A2(n1068), .ZN(n1066) );
NOR2_X1 U765 ( .A1(n1069), .A2(n1070), .ZN(n1064) );
XOR2_X1 U766 ( .A(KEYINPUT51), .B(G478), .Z(n1070) );
INV_X1 U767 ( .A(n1071), .ZN(n1069) );
NOR2_X1 U768 ( .A1(n1053), .A2(n1072), .ZN(n1061) );
XOR2_X1 U769 ( .A(KEYINPUT55), .B(n1073), .Z(n1072) );
NOR2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U771 ( .A(n1076), .B(KEYINPUT26), .Z(n1075) );
NAND2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XNOR2_X1 U773 ( .A(n1079), .B(KEYINPUT43), .ZN(n1077) );
XNOR2_X1 U774 ( .A(KEYINPUT33), .B(n1056), .ZN(n1060) );
XOR2_X1 U775 ( .A(n1080), .B(n1081), .Z(G72) );
NOR2_X1 U776 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NAND2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1080) );
NAND3_X1 U779 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
NAND2_X1 U780 ( .A1(G953), .A2(n1091), .ZN(n1089) );
NAND2_X1 U781 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U782 ( .A1(G900), .A2(n1094), .ZN(n1092) );
NAND2_X1 U783 ( .A1(n1095), .A2(n1083), .ZN(n1088) );
OR2_X1 U784 ( .A1(n1093), .A2(n1094), .ZN(n1095) );
INV_X1 U785 ( .A(KEYINPUT25), .ZN(n1093) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1096), .ZN(n1086) );
NAND2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U788 ( .A1(G900), .A2(n1099), .ZN(n1098) );
NAND2_X1 U789 ( .A1(n1090), .A2(n1100), .ZN(n1099) );
NAND2_X1 U790 ( .A1(KEYINPUT25), .A2(G953), .ZN(n1100) );
NAND2_X1 U791 ( .A1(n1101), .A2(n1083), .ZN(n1097) );
NAND2_X1 U792 ( .A1(KEYINPUT25), .A2(n1090), .ZN(n1101) );
XNOR2_X1 U793 ( .A(n1102), .B(n1103), .ZN(n1094) );
XOR2_X1 U794 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U795 ( .A1(KEYINPUT45), .A2(n1106), .ZN(n1105) );
XNOR2_X1 U796 ( .A(KEYINPUT11), .B(n1107), .ZN(n1106) );
NAND2_X1 U797 ( .A1(n1108), .A2(n1109), .ZN(n1104) );
NAND2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XNOR2_X1 U799 ( .A(G125), .B(KEYINPUT1), .ZN(n1110) );
XOR2_X1 U800 ( .A(KEYINPUT37), .B(n1112), .Z(n1108) );
NOR2_X1 U801 ( .A1(n1111), .A2(n1113), .ZN(n1112) );
XNOR2_X1 U802 ( .A(G140), .B(KEYINPUT36), .ZN(n1111) );
XNOR2_X1 U803 ( .A(n1114), .B(n1115), .ZN(n1102) );
XOR2_X1 U804 ( .A(n1116), .B(n1117), .Z(G69) );
XOR2_X1 U805 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U806 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
INV_X1 U807 ( .A(n1122), .ZN(n1121) );
XOR2_X1 U808 ( .A(n1123), .B(n1124), .Z(n1120) );
NAND2_X1 U809 ( .A1(KEYINPUT61), .A2(n1125), .ZN(n1123) );
NAND2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1118) );
XNOR2_X1 U811 ( .A(KEYINPUT0), .B(n1083), .ZN(n1126) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1083), .ZN(n1116) );
AND2_X1 U813 ( .A1(G224), .A2(G898), .ZN(n1128) );
NOR2_X1 U814 ( .A1(n1129), .A2(n1130), .ZN(G66) );
NOR2_X1 U815 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U816 ( .A(KEYINPUT19), .B(n1133), .Z(n1132) );
NOR2_X1 U817 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U818 ( .A(n1136), .B(KEYINPUT6), .Z(n1135) );
INV_X1 U819 ( .A(n1137), .ZN(n1134) );
NOR2_X1 U820 ( .A1(n1136), .A2(n1137), .ZN(n1131) );
NAND2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NOR2_X1 U822 ( .A1(n1129), .A2(n1140), .ZN(G63) );
XOR2_X1 U823 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U824 ( .A1(n1138), .A2(G478), .ZN(n1141) );
NOR2_X1 U825 ( .A1(n1129), .A2(n1143), .ZN(G60) );
NOR3_X1 U826 ( .A1(n1079), .A2(n1144), .A3(n1145), .ZN(n1143) );
NOR4_X1 U827 ( .A1(n1146), .A2(n1147), .A3(KEYINPUT20), .A4(n1078), .ZN(n1145) );
INV_X1 U828 ( .A(n1138), .ZN(n1147) );
NOR2_X1 U829 ( .A1(n1148), .A2(n1149), .ZN(n1144) );
NOR3_X1 U830 ( .A1(n1078), .A2(KEYINPUT20), .A3(n1045), .ZN(n1149) );
XOR2_X1 U831 ( .A(G104), .B(n1150), .Z(G6) );
NOR2_X1 U832 ( .A1(n1129), .A2(n1151), .ZN(G57) );
XOR2_X1 U833 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U834 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U835 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U836 ( .A(n1158), .B(KEYINPUT2), .Z(n1157) );
NAND2_X1 U837 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U838 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
XNOR2_X1 U839 ( .A(KEYINPUT60), .B(G101), .ZN(n1159) );
NOR2_X1 U840 ( .A1(n1161), .A2(n1162), .ZN(n1154) );
XOR2_X1 U841 ( .A(n1163), .B(KEYINPUT27), .Z(n1162) );
NAND3_X1 U842 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1163) );
XNOR2_X1 U843 ( .A(KEYINPUT34), .B(n1167), .ZN(n1166) );
NAND2_X1 U844 ( .A1(n1168), .A2(n1169), .ZN(n1164) );
NOR2_X1 U845 ( .A1(n1170), .A2(n1171), .ZN(n1161) );
NOR2_X1 U846 ( .A1(n1172), .A2(n1168), .ZN(n1170) );
XNOR2_X1 U847 ( .A(n1173), .B(KEYINPUT46), .ZN(n1168) );
NAND2_X1 U848 ( .A1(n1138), .A2(G472), .ZN(n1152) );
NOR2_X1 U849 ( .A1(n1174), .A2(n1175), .ZN(G54) );
XOR2_X1 U850 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR3_X1 U851 ( .A1(n1067), .A2(n1178), .A3(n1179), .ZN(n1177) );
NOR2_X1 U852 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
INV_X1 U853 ( .A(KEYINPUT9), .ZN(n1181) );
NOR2_X1 U854 ( .A1(G902), .A2(n1045), .ZN(n1180) );
NOR2_X1 U855 ( .A1(KEYINPUT9), .A2(n1138), .ZN(n1178) );
NAND3_X1 U856 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1176) );
NAND2_X1 U857 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U858 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U859 ( .A(n1189), .B(n1190), .Z(n1185) );
NAND4_X1 U860 ( .A1(n1191), .A2(n1188), .A3(n1187), .A4(n1192), .ZN(n1183) );
INV_X1 U861 ( .A(KEYINPUT8), .ZN(n1188) );
XNOR2_X1 U862 ( .A(n1189), .B(n1190), .ZN(n1191) );
OR2_X1 U863 ( .A1(n1192), .A2(n1187), .ZN(n1182) );
XOR2_X1 U864 ( .A(n1193), .B(n1169), .Z(n1187) );
INV_X1 U865 ( .A(KEYINPUT18), .ZN(n1192) );
NOR2_X1 U866 ( .A1(n1194), .A2(n1195), .ZN(n1174) );
XNOR2_X1 U867 ( .A(G952), .B(KEYINPUT63), .ZN(n1194) );
NOR2_X1 U868 ( .A1(n1129), .A2(n1196), .ZN(G51) );
XOR2_X1 U869 ( .A(n1197), .B(n1198), .Z(n1196) );
XNOR2_X1 U870 ( .A(n1199), .B(n1200), .ZN(n1198) );
NAND2_X1 U871 ( .A1(n1138), .A2(n1201), .ZN(n1199) );
NOR2_X1 U872 ( .A1(n1202), .A2(n1045), .ZN(n1138) );
NOR2_X1 U873 ( .A1(n1127), .A2(n1090), .ZN(n1045) );
NAND4_X1 U874 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1090) );
NOR4_X1 U875 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
NAND2_X1 U876 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
NAND2_X1 U877 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
OR2_X1 U878 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U879 ( .A(KEYINPUT17), .B(n1217), .Z(n1213) );
NAND4_X1 U880 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1127) );
NOR4_X1 U881 ( .A1(n1016), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1221) );
AND3_X1 U882 ( .A1(n1056), .A2(n1032), .A3(n1225), .ZN(n1016) );
NOR2_X1 U883 ( .A1(n1226), .A2(n1150), .ZN(n1220) );
AND3_X1 U884 ( .A1(n1056), .A2(n1225), .A3(n1227), .ZN(n1150) );
XOR2_X1 U885 ( .A(n1228), .B(KEYINPUT38), .Z(n1197) );
NAND3_X1 U886 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1228) );
NAND2_X1 U887 ( .A1(KEYINPUT56), .A2(n1232), .ZN(n1231) );
OR3_X1 U888 ( .A1(n1232), .A2(KEYINPUT56), .A3(n1233), .ZN(n1230) );
NAND2_X1 U889 ( .A1(n1233), .A2(n1234), .ZN(n1229) );
NAND2_X1 U890 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
INV_X1 U891 ( .A(KEYINPUT56), .ZN(n1236) );
XNOR2_X1 U892 ( .A(n1232), .B(KEYINPUT22), .ZN(n1235) );
XNOR2_X1 U893 ( .A(n1237), .B(KEYINPUT24), .ZN(n1233) );
NOR2_X1 U894 ( .A1(n1195), .A2(G952), .ZN(n1129) );
XNOR2_X1 U895 ( .A(KEYINPUT10), .B(n1083), .ZN(n1195) );
XNOR2_X1 U896 ( .A(G146), .B(n1203), .ZN(G48) );
NAND3_X1 U897 ( .A1(n1227), .A2(n1211), .A3(n1238), .ZN(n1203) );
XNOR2_X1 U898 ( .A(G143), .B(n1204), .ZN(G45) );
NAND4_X1 U899 ( .A1(n1211), .A2(n1239), .A3(n1059), .A4(n1240), .ZN(n1204) );
NOR3_X1 U900 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1240) );
XOR2_X1 U901 ( .A(n1210), .B(n1244), .Z(G42) );
NOR2_X1 U902 ( .A1(KEYINPUT47), .A2(n1245), .ZN(n1244) );
NOR3_X1 U903 ( .A1(n1053), .A2(n1038), .A3(n1215), .ZN(n1210) );
XOR2_X1 U904 ( .A(n1246), .B(n1209), .Z(G39) );
AND3_X1 U905 ( .A1(n1036), .A2(n1027), .A3(n1238), .ZN(n1209) );
XNOR2_X1 U906 ( .A(G137), .B(KEYINPUT15), .ZN(n1246) );
XNOR2_X1 U907 ( .A(n1107), .B(n1208), .ZN(G36) );
AND2_X1 U908 ( .A1(n1247), .A2(n1032), .ZN(n1208) );
XOR2_X1 U909 ( .A(G131), .B(n1207), .Z(G33) );
AND2_X1 U910 ( .A1(n1247), .A2(n1227), .ZN(n1207) );
AND4_X1 U911 ( .A1(n1059), .A2(n1027), .A3(n1239), .A4(n1248), .ZN(n1247) );
INV_X1 U912 ( .A(n1053), .ZN(n1027) );
NAND2_X1 U913 ( .A1(n1058), .A2(n1249), .ZN(n1053) );
XOR2_X1 U914 ( .A(G128), .B(n1250), .Z(G30) );
NOR2_X1 U915 ( .A1(n1055), .A2(n1251), .ZN(n1250) );
XOR2_X1 U916 ( .A(KEYINPUT48), .B(n1217), .Z(n1251) );
AND2_X1 U917 ( .A1(n1238), .A2(n1032), .ZN(n1217) );
NOR4_X1 U918 ( .A1(n1056), .A2(n1052), .A3(n1038), .A4(n1241), .ZN(n1238) );
INV_X1 U919 ( .A(n1248), .ZN(n1241) );
INV_X1 U920 ( .A(n1239), .ZN(n1038) );
INV_X1 U921 ( .A(n1211), .ZN(n1055) );
XOR2_X1 U922 ( .A(G101), .B(n1226), .Z(G3) );
AND3_X1 U923 ( .A1(n1036), .A2(n1239), .A3(n1252), .ZN(n1226) );
XNOR2_X1 U924 ( .A(n1113), .B(n1253), .ZN(G27) );
NOR4_X1 U925 ( .A1(KEYINPUT49), .A2(n1254), .A3(n1216), .A4(n1215), .ZN(n1253) );
NAND4_X1 U926 ( .A1(n1052), .A2(n1227), .A3(n1023), .A4(n1248), .ZN(n1215) );
NAND2_X1 U927 ( .A1(n1029), .A2(n1255), .ZN(n1248) );
NAND4_X1 U928 ( .A1(G902), .A2(G953), .A3(n1256), .A4(n1085), .ZN(n1255) );
INV_X1 U929 ( .A(G900), .ZN(n1085) );
XNOR2_X1 U930 ( .A(n1211), .B(KEYINPUT52), .ZN(n1254) );
XNOR2_X1 U931 ( .A(G122), .B(n1218), .ZN(G24) );
NAND3_X1 U932 ( .A1(n1056), .A2(n1257), .A3(n1258), .ZN(n1218) );
NOR3_X1 U933 ( .A1(n1024), .A2(n1242), .A3(n1243), .ZN(n1258) );
INV_X1 U934 ( .A(n1023), .ZN(n1056) );
XNOR2_X1 U935 ( .A(G119), .B(n1259), .ZN(G21) );
NOR2_X1 U936 ( .A1(n1260), .A2(KEYINPUT4), .ZN(n1259) );
INV_X1 U937 ( .A(n1219), .ZN(n1260) );
NAND4_X1 U938 ( .A1(n1257), .A2(n1036), .A3(n1023), .A4(n1024), .ZN(n1219) );
XOR2_X1 U939 ( .A(G116), .B(n1224), .Z(G18) );
AND3_X1 U940 ( .A1(n1059), .A2(n1032), .A3(n1257), .ZN(n1224) );
AND3_X1 U941 ( .A1(n1030), .A2(n1261), .A3(n1211), .ZN(n1257) );
NOR2_X1 U942 ( .A1(n1262), .A2(n1242), .ZN(n1032) );
XOR2_X1 U943 ( .A(G113), .B(n1223), .Z(G15) );
AND3_X1 U944 ( .A1(n1252), .A2(n1030), .A3(n1227), .ZN(n1223) );
INV_X1 U945 ( .A(n1043), .ZN(n1227) );
NAND2_X1 U946 ( .A1(n1242), .A2(n1262), .ZN(n1043) );
AND3_X1 U947 ( .A1(n1263), .A2(n1261), .A3(n1059), .ZN(n1252) );
NOR2_X1 U948 ( .A1(n1023), .A2(n1052), .ZN(n1059) );
XOR2_X1 U949 ( .A(G110), .B(n1222), .Z(G12) );
AND3_X1 U950 ( .A1(n1225), .A2(n1023), .A3(n1036), .ZN(n1222) );
AND2_X1 U951 ( .A1(n1242), .A2(n1243), .ZN(n1036) );
INV_X1 U952 ( .A(n1262), .ZN(n1243) );
NAND2_X1 U953 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
NAND2_X1 U954 ( .A1(n1266), .A2(n1078), .ZN(n1265) );
NAND2_X1 U955 ( .A1(KEYINPUT53), .A2(n1267), .ZN(n1266) );
INV_X1 U956 ( .A(n1079), .ZN(n1267) );
NAND2_X1 U957 ( .A1(n1074), .A2(KEYINPUT53), .ZN(n1264) );
NOR2_X1 U958 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
NOR2_X1 U959 ( .A1(G902), .A2(n1148), .ZN(n1079) );
INV_X1 U960 ( .A(n1146), .ZN(n1148) );
NAND3_X1 U961 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1146) );
NAND2_X1 U962 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NAND3_X1 U963 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1272) );
NAND2_X1 U964 ( .A1(KEYINPUT28), .A2(n1276), .ZN(n1275) );
NAND2_X1 U965 ( .A1(n1277), .A2(n1278), .ZN(n1274) );
INV_X1 U966 ( .A(KEYINPUT3), .ZN(n1278) );
NAND2_X1 U967 ( .A1(KEYINPUT3), .A2(n1279), .ZN(n1273) );
NAND2_X1 U968 ( .A1(n1277), .A2(n1280), .ZN(n1279) );
NAND2_X1 U969 ( .A1(KEYINPUT41), .A2(n1281), .ZN(n1280) );
INV_X1 U970 ( .A(n1282), .ZN(n1271) );
NAND4_X1 U971 ( .A1(n1277), .A2(n1276), .A3(n1282), .A4(n1281), .ZN(n1269) );
INV_X1 U972 ( .A(KEYINPUT28), .ZN(n1281) );
INV_X1 U973 ( .A(KEYINPUT41), .ZN(n1276) );
NAND2_X1 U974 ( .A1(KEYINPUT28), .A2(n1283), .ZN(n1268) );
NAND2_X1 U975 ( .A1(n1277), .A2(n1284), .ZN(n1283) );
NAND2_X1 U976 ( .A1(KEYINPUT41), .A2(n1282), .ZN(n1284) );
XNOR2_X1 U977 ( .A(n1285), .B(n1286), .ZN(n1282) );
XNOR2_X1 U978 ( .A(G122), .B(n1287), .ZN(n1285) );
NAND2_X1 U979 ( .A1(n1288), .A2(n1289), .ZN(n1277) );
NAND2_X1 U980 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U981 ( .A(KEYINPUT59), .B(n1292), .Z(n1288) );
NOR2_X1 U982 ( .A1(n1290), .A2(n1291), .ZN(n1292) );
XNOR2_X1 U983 ( .A(n1293), .B(n1294), .ZN(n1291) );
XOR2_X1 U984 ( .A(G143), .B(G131), .Z(n1294) );
NAND2_X1 U985 ( .A1(G214), .A2(n1295), .ZN(n1293) );
XNOR2_X1 U986 ( .A(n1113), .B(n1296), .ZN(n1290) );
XNOR2_X1 U987 ( .A(G146), .B(n1245), .ZN(n1296) );
INV_X1 U988 ( .A(G475), .ZN(n1078) );
NOR2_X1 U989 ( .A1(n1297), .A2(n1063), .ZN(n1242) );
NOR2_X1 U990 ( .A1(n1071), .A2(G478), .ZN(n1063) );
AND2_X1 U991 ( .A1(G478), .A2(n1071), .ZN(n1297) );
NAND2_X1 U992 ( .A1(n1142), .A2(n1202), .ZN(n1071) );
XNOR2_X1 U993 ( .A(n1298), .B(n1299), .ZN(n1142) );
XOR2_X1 U994 ( .A(n1300), .B(n1301), .Z(n1299) );
XNOR2_X1 U995 ( .A(n1015), .B(n1302), .ZN(n1301) );
AND4_X1 U996 ( .A1(n1303), .A2(n1083), .A3(G234), .A4(G217), .ZN(n1302) );
INV_X1 U997 ( .A(KEYINPUT44), .ZN(n1303) );
INV_X1 U998 ( .A(G107), .ZN(n1015) );
XNOR2_X1 U999 ( .A(G116), .B(n1304), .ZN(n1298) );
XNOR2_X1 U1000 ( .A(n1107), .B(G122), .ZN(n1304) );
INV_X1 U1001 ( .A(G134), .ZN(n1107) );
XNOR2_X1 U1002 ( .A(n1305), .B(n1139), .ZN(n1023) );
AND2_X1 U1003 ( .A1(G217), .A2(n1306), .ZN(n1139) );
NAND2_X1 U1004 ( .A1(n1136), .A2(n1202), .ZN(n1305) );
XOR2_X1 U1005 ( .A(n1307), .B(n1308), .Z(n1136) );
XNOR2_X1 U1006 ( .A(n1190), .B(n1309), .ZN(n1308) );
XOR2_X1 U1007 ( .A(n1310), .B(n1311), .Z(n1309) );
AND3_X1 U1008 ( .A1(G221), .A2(n1083), .A3(G234), .ZN(n1311) );
NAND2_X1 U1009 ( .A1(KEYINPUT54), .A2(n1113), .ZN(n1310) );
INV_X1 U1010 ( .A(G125), .ZN(n1113) );
XNOR2_X1 U1011 ( .A(G110), .B(n1245), .ZN(n1190) );
INV_X1 U1012 ( .A(G140), .ZN(n1245) );
XOR2_X1 U1013 ( .A(n1312), .B(n1313), .Z(n1307) );
NOR2_X1 U1014 ( .A1(KEYINPUT32), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U1015 ( .A(G119), .B(G128), .ZN(n1314) );
XNOR2_X1 U1016 ( .A(G137), .B(G146), .ZN(n1312) );
AND4_X1 U1017 ( .A1(n1052), .A2(n1263), .A3(n1239), .A4(n1261), .ZN(n1225) );
NAND2_X1 U1018 ( .A1(n1029), .A2(n1315), .ZN(n1261) );
NAND3_X1 U1019 ( .A1(n1122), .A2(n1256), .A3(G902), .ZN(n1315) );
NOR2_X1 U1020 ( .A1(n1083), .A2(G898), .ZN(n1122) );
NAND3_X1 U1021 ( .A1(n1256), .A2(n1083), .A3(G952), .ZN(n1029) );
NAND2_X1 U1022 ( .A1(G237), .A2(G234), .ZN(n1256) );
NAND2_X1 U1023 ( .A1(n1316), .A2(n1317), .ZN(n1239) );
NAND2_X1 U1024 ( .A1(n1030), .A2(n1318), .ZN(n1317) );
INV_X1 U1025 ( .A(n1216), .ZN(n1030) );
NAND2_X1 U1026 ( .A1(n1041), .A2(n1319), .ZN(n1216) );
OR3_X1 U1027 ( .A1(n1041), .A2(n1040), .A3(n1318), .ZN(n1316) );
INV_X1 U1028 ( .A(KEYINPUT62), .ZN(n1318) );
INV_X1 U1029 ( .A(n1319), .ZN(n1040) );
NAND2_X1 U1030 ( .A1(G221), .A2(n1306), .ZN(n1319) );
NAND2_X1 U1031 ( .A1(G234), .A2(n1202), .ZN(n1306) );
XOR2_X1 U1032 ( .A(n1320), .B(n1068), .Z(n1041) );
NAND2_X1 U1033 ( .A1(n1321), .A2(n1202), .ZN(n1068) );
XOR2_X1 U1034 ( .A(n1169), .B(n1322), .Z(n1321) );
XNOR2_X1 U1035 ( .A(n1323), .B(n1324), .ZN(n1322) );
NOR2_X1 U1036 ( .A1(KEYINPUT29), .A2(n1193), .ZN(n1324) );
XOR2_X1 U1037 ( .A(n1325), .B(n1326), .Z(n1193) );
XNOR2_X1 U1038 ( .A(G101), .B(n1173), .ZN(n1326) );
INV_X1 U1039 ( .A(n1115), .ZN(n1173) );
NAND2_X1 U1040 ( .A1(KEYINPUT31), .A2(n1327), .ZN(n1323) );
XOR2_X1 U1041 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U1042 ( .A(G140), .B(n1189), .ZN(n1329) );
NOR2_X1 U1043 ( .A1(n1084), .A2(G953), .ZN(n1189) );
INV_X1 U1044 ( .A(G227), .ZN(n1084) );
NAND2_X1 U1045 ( .A1(KEYINPUT12), .A2(G110), .ZN(n1328) );
NAND2_X1 U1046 ( .A1(KEYINPUT21), .A2(n1067), .ZN(n1320) );
INV_X1 U1047 ( .A(G469), .ZN(n1067) );
XNOR2_X1 U1048 ( .A(n1211), .B(KEYINPUT57), .ZN(n1263) );
NOR2_X1 U1049 ( .A1(n1058), .A2(n1057), .ZN(n1211) );
INV_X1 U1050 ( .A(n1249), .ZN(n1057) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1330), .ZN(n1249) );
XOR2_X1 U1052 ( .A(n1331), .B(n1201), .Z(n1058) );
AND2_X1 U1053 ( .A1(G210), .A2(n1330), .ZN(n1201) );
NAND2_X1 U1054 ( .A1(n1332), .A2(n1202), .ZN(n1330) );
INV_X1 U1055 ( .A(G237), .ZN(n1332) );
NAND2_X1 U1056 ( .A1(n1333), .A2(n1202), .ZN(n1331) );
XNOR2_X1 U1057 ( .A(n1334), .B(n1335), .ZN(n1333) );
INV_X1 U1058 ( .A(n1200), .ZN(n1335) );
XOR2_X1 U1059 ( .A(n1124), .B(n1125), .Z(n1200) );
XNOR2_X1 U1060 ( .A(G110), .B(n1336), .ZN(n1125) );
XNOR2_X1 U1061 ( .A(KEYINPUT30), .B(n1337), .ZN(n1336) );
INV_X1 U1062 ( .A(G122), .ZN(n1337) );
XNOR2_X1 U1063 ( .A(n1338), .B(n1167), .ZN(n1124) );
NAND3_X1 U1064 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1338) );
NAND2_X1 U1065 ( .A1(KEYINPUT5), .A2(n1342), .ZN(n1341) );
OR3_X1 U1066 ( .A1(n1342), .A2(KEYINPUT5), .A3(G101), .ZN(n1340) );
NAND2_X1 U1067 ( .A1(G101), .A2(n1343), .ZN(n1339) );
NAND2_X1 U1068 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
INV_X1 U1069 ( .A(KEYINPUT5), .ZN(n1345) );
XNOR2_X1 U1070 ( .A(KEYINPUT23), .B(n1342), .ZN(n1344) );
INV_X1 U1071 ( .A(n1325), .ZN(n1342) );
XOR2_X1 U1072 ( .A(G107), .B(n1287), .Z(n1325) );
XOR2_X1 U1073 ( .A(G104), .B(KEYINPUT7), .Z(n1287) );
NAND2_X1 U1074 ( .A1(n1346), .A2(KEYINPUT35), .ZN(n1334) );
XOR2_X1 U1075 ( .A(n1347), .B(n1232), .Z(n1346) );
XOR2_X1 U1076 ( .A(G125), .B(n1115), .Z(n1232) );
XOR2_X1 U1077 ( .A(n1237), .B(KEYINPUT42), .Z(n1347) );
NAND2_X1 U1078 ( .A1(G224), .A2(n1083), .ZN(n1237) );
INV_X1 U1079 ( .A(G953), .ZN(n1083) );
INV_X1 U1080 ( .A(n1024), .ZN(n1052) );
XNOR2_X1 U1081 ( .A(n1348), .B(G472), .ZN(n1024) );
NAND2_X1 U1082 ( .A1(n1349), .A2(n1202), .ZN(n1348) );
INV_X1 U1083 ( .A(G902), .ZN(n1202) );
XOR2_X1 U1084 ( .A(n1350), .B(n1351), .Z(n1349) );
NOR2_X1 U1085 ( .A1(KEYINPUT40), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1086 ( .A(n1160), .B(n1353), .Z(n1352) );
XNOR2_X1 U1087 ( .A(G101), .B(KEYINPUT50), .ZN(n1353) );
NAND2_X1 U1088 ( .A1(G210), .A2(n1295), .ZN(n1160) );
NOR2_X1 U1089 ( .A1(G953), .A2(G237), .ZN(n1295) );
NOR2_X1 U1090 ( .A1(n1354), .A2(n1355), .ZN(n1350) );
XOR2_X1 U1091 ( .A(n1356), .B(KEYINPUT14), .Z(n1355) );
NAND3_X1 U1092 ( .A1(n1357), .A2(n1165), .A3(n1167), .ZN(n1356) );
INV_X1 U1093 ( .A(n1358), .ZN(n1167) );
INV_X1 U1094 ( .A(n1172), .ZN(n1165) );
NAND2_X1 U1095 ( .A1(n1115), .A2(n1169), .ZN(n1357) );
NOR2_X1 U1096 ( .A1(n1359), .A2(n1171), .ZN(n1354) );
NAND2_X1 U1097 ( .A1(n1358), .A2(n1360), .ZN(n1171) );
OR2_X1 U1098 ( .A1(n1169), .A2(n1172), .ZN(n1360) );
XNOR2_X1 U1099 ( .A(n1361), .B(n1286), .ZN(n1358) );
XOR2_X1 U1100 ( .A(G113), .B(KEYINPUT13), .Z(n1286) );
XNOR2_X1 U1101 ( .A(G116), .B(G119), .ZN(n1361) );
NOR2_X1 U1102 ( .A1(n1172), .A2(n1115), .ZN(n1359) );
NOR2_X1 U1103 ( .A1(n1169), .A2(n1115), .ZN(n1172) );
XOR2_X1 U1104 ( .A(G146), .B(n1300), .Z(n1115) );
XOR2_X1 U1105 ( .A(G128), .B(G143), .Z(n1300) );
XNOR2_X1 U1106 ( .A(n1362), .B(n1114), .ZN(n1169) );
XNOR2_X1 U1107 ( .A(G131), .B(n1363), .ZN(n1114) );
INV_X1 U1108 ( .A(G137), .ZN(n1363) );
XNOR2_X1 U1109 ( .A(G134), .B(KEYINPUT39), .ZN(n1362) );
endmodule


