//Key = 1100011110101111111000011100001010011100010001111010000100010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351;

XNOR2_X1 U740 ( .A(G107), .B(n1019), .ZN(G9) );
NOR2_X1 U741 ( .A1(n1020), .A2(n1021), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
XNOR2_X1 U743 ( .A(n1026), .B(KEYINPUT37), .ZN(n1024) );
NAND3_X1 U744 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1022) );
NAND4_X1 U745 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
NAND2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U747 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1034) );
INV_X1 U748 ( .A(KEYINPUT12), .ZN(n1037) );
NAND4_X1 U749 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1032) );
NAND2_X1 U750 ( .A1(n1038), .A2(n1043), .ZN(n1041) );
NAND2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U752 ( .A1(KEYINPUT12), .A2(n1036), .ZN(n1045) );
NAND3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1040) );
INV_X1 U754 ( .A(KEYINPUT38), .ZN(n1047) );
NAND2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1039) );
XOR2_X1 U756 ( .A(KEYINPUT21), .B(n1046), .Z(n1050) );
NAND3_X1 U757 ( .A1(n1046), .A2(n1051), .A3(n1042), .ZN(n1027) );
INV_X1 U758 ( .A(n1035), .ZN(n1042) );
NAND2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND4_X1 U760 ( .A1(n1048), .A2(KEYINPUT38), .A3(n1031), .A4(n1054), .ZN(n1053) );
INV_X1 U761 ( .A(n1030), .ZN(n1054) );
XOR2_X1 U762 ( .A(n1055), .B(KEYINPUT36), .Z(n1048) );
NAND2_X1 U763 ( .A1(n1038), .A2(n1056), .ZN(n1052) );
NAND2_X1 U764 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U765 ( .A1(n1030), .A2(n1059), .ZN(n1058) );
NAND2_X1 U766 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U767 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U768 ( .A1(n1031), .A2(n1064), .ZN(n1057) );
NAND2_X1 U769 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR3_X1 U771 ( .A1(n1069), .A2(G953), .A3(n1026), .ZN(n1020) );
AND4_X1 U772 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1026) );
NOR4_X1 U773 ( .A1(n1074), .A2(n1062), .A3(n1075), .A4(n1067), .ZN(n1073) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
AND2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NAND3_X1 U776 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1074) );
NOR3_X1 U777 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1072) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U779 ( .A(KEYINPUT47), .B(G478), .Z(n1087) );
AND2_X1 U780 ( .A1(n1088), .A2(n1086), .ZN(n1084) );
XOR2_X1 U781 ( .A(n1089), .B(n1090), .Z(n1083) );
XOR2_X1 U782 ( .A(n1091), .B(KEYINPUT9), .Z(n1071) );
NAND2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U784 ( .A(n1094), .B(KEYINPUT18), .Z(n1092) );
NOR2_X1 U785 ( .A1(n1095), .A2(n1096), .ZN(n1070) );
XOR2_X1 U786 ( .A(n1097), .B(n1098), .Z(n1096) );
XNOR2_X1 U787 ( .A(n1099), .B(KEYINPUT13), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1100), .A2(n1101), .ZN(n1095) );
XOR2_X1 U789 ( .A(KEYINPUT16), .B(G475), .Z(n1101) );
XOR2_X1 U790 ( .A(n1025), .B(KEYINPUT61), .Z(n1069) );
INV_X1 U791 ( .A(G952), .ZN(n1025) );
XOR2_X1 U792 ( .A(n1102), .B(n1103), .Z(G72) );
NOR2_X1 U793 ( .A1(n1104), .A2(n1028), .ZN(n1103) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U795 ( .A1(n1107), .A2(n1108), .ZN(n1102) );
NAND2_X1 U796 ( .A1(n1109), .A2(n1028), .ZN(n1108) );
XOR2_X1 U797 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XNOR2_X1 U799 ( .A(n1114), .B(KEYINPUT56), .ZN(n1110) );
NAND3_X1 U800 ( .A1(n1114), .A2(G900), .A3(G953), .ZN(n1107) );
NOR2_X1 U801 ( .A1(KEYINPUT63), .A2(n1115), .ZN(n1114) );
XOR2_X1 U802 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U803 ( .A(G125), .B(n1118), .Z(n1117) );
NOR2_X1 U804 ( .A1(KEYINPUT29), .A2(n1119), .ZN(n1118) );
XOR2_X1 U805 ( .A(n1120), .B(n1121), .Z(G69) );
XOR2_X1 U806 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND2_X1 U807 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U808 ( .A1(G953), .A2(n1126), .ZN(n1125) );
XNOR2_X1 U809 ( .A(n1127), .B(n1128), .ZN(n1124) );
XOR2_X1 U810 ( .A(n1129), .B(KEYINPUT0), .Z(n1127) );
NAND2_X1 U811 ( .A1(n1130), .A2(n1028), .ZN(n1122) );
XOR2_X1 U812 ( .A(n1131), .B(KEYINPUT53), .Z(n1130) );
NAND2_X1 U813 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U814 ( .A1(n1134), .A2(n1028), .ZN(n1120) );
NOR2_X1 U815 ( .A1(n1135), .A2(n1126), .ZN(n1134) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(G66) );
NOR3_X1 U817 ( .A1(n1099), .A2(n1138), .A3(n1139), .ZN(n1137) );
NOR3_X1 U818 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1139) );
INV_X1 U819 ( .A(n1143), .ZN(n1140) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1143), .ZN(n1138) );
AND2_X1 U821 ( .A1(n1023), .A2(G217), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1136), .A2(n1145), .ZN(G63) );
XNOR2_X1 U823 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U824 ( .A1(n1088), .A2(n1142), .ZN(n1147) );
INV_X1 U825 ( .A(G478), .ZN(n1088) );
NOR2_X1 U826 ( .A1(n1136), .A2(n1148), .ZN(G60) );
XOR2_X1 U827 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR2_X1 U828 ( .A1(n1151), .A2(n1142), .ZN(n1149) );
NAND2_X1 U829 ( .A1(n1152), .A2(n1153), .ZN(G6) );
NAND2_X1 U830 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U831 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NAND2_X1 U832 ( .A1(KEYINPUT57), .A2(KEYINPUT10), .ZN(n1157) );
INV_X1 U833 ( .A(G104), .ZN(n1156) );
NAND3_X1 U834 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1152) );
INV_X1 U835 ( .A(KEYINPUT57), .ZN(n1160) );
OR2_X1 U836 ( .A1(G104), .A2(KEYINPUT10), .ZN(n1159) );
NAND2_X1 U837 ( .A1(KEYINPUT10), .A2(n1161), .ZN(n1158) );
OR2_X1 U838 ( .A1(n1155), .A2(G104), .ZN(n1161) );
NOR2_X1 U839 ( .A1(n1136), .A2(n1162), .ZN(G57) );
XOR2_X1 U840 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U841 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U842 ( .A1(n1089), .A2(n1142), .ZN(n1165) );
XOR2_X1 U843 ( .A(n1167), .B(n1168), .Z(n1163) );
NOR2_X1 U844 ( .A1(n1136), .A2(n1169), .ZN(G54) );
XOR2_X1 U845 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U846 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U847 ( .A1(n1077), .A2(n1142), .ZN(n1172) );
XOR2_X1 U848 ( .A(n1174), .B(n1175), .Z(n1170) );
XNOR2_X1 U849 ( .A(G101), .B(n1176), .ZN(n1175) );
NAND3_X1 U850 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
NAND2_X1 U851 ( .A1(KEYINPUT4), .A2(G110), .ZN(n1179) );
OR3_X1 U852 ( .A1(n1180), .A2(KEYINPUT4), .A3(G140), .ZN(n1178) );
NAND2_X1 U853 ( .A1(G140), .A2(n1180), .ZN(n1177) );
NAND2_X1 U854 ( .A1(KEYINPUT23), .A2(n1181), .ZN(n1180) );
NOR2_X1 U855 ( .A1(KEYINPUT11), .A2(n1166), .ZN(n1174) );
NOR2_X1 U856 ( .A1(n1136), .A2(n1182), .ZN(G51) );
XOR2_X1 U857 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U858 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U859 ( .A1(n1094), .A2(n1142), .ZN(n1186) );
NAND2_X1 U860 ( .A1(G902), .A2(n1023), .ZN(n1142) );
NAND4_X1 U861 ( .A1(n1187), .A2(n1132), .A3(n1188), .A4(n1189), .ZN(n1023) );
XOR2_X1 U862 ( .A(KEYINPUT49), .B(n1133), .Z(n1189) );
AND3_X1 U863 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1133) );
NAND4_X1 U864 ( .A1(n1193), .A2(n1031), .A3(n1194), .A4(n1195), .ZN(n1192) );
OR2_X1 U865 ( .A1(n1196), .A2(n1049), .ZN(n1195) );
NAND2_X1 U866 ( .A1(n1197), .A2(n1198), .ZN(n1190) );
XNOR2_X1 U867 ( .A(KEYINPUT2), .B(n1199), .ZN(n1198) );
XNOR2_X1 U868 ( .A(KEYINPUT52), .B(n1112), .ZN(n1188) );
NAND3_X1 U869 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1112) );
NAND2_X1 U870 ( .A1(n1197), .A2(n1203), .ZN(n1202) );
NAND2_X1 U871 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NAND2_X1 U872 ( .A1(n1206), .A2(n1049), .ZN(n1204) );
AND4_X1 U873 ( .A1(n1155), .A2(n1207), .A3(n1208), .A4(n1019), .ZN(n1132) );
NAND3_X1 U874 ( .A1(n1046), .A2(n1209), .A3(n1196), .ZN(n1019) );
NAND3_X1 U875 ( .A1(n1046), .A2(n1209), .A3(n1049), .ZN(n1155) );
INV_X1 U876 ( .A(n1113), .ZN(n1187) );
NAND4_X1 U877 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1113) );
NAND4_X1 U878 ( .A1(n1030), .A2(n1214), .A3(n1049), .A4(n1215), .ZN(n1211) );
NAND2_X1 U879 ( .A1(n1216), .A2(n1197), .ZN(n1210) );
XNOR2_X1 U880 ( .A(n1217), .B(KEYINPUT6), .ZN(n1216) );
NAND3_X1 U881 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1185) );
NAND2_X1 U882 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
OR3_X1 U883 ( .A1(n1222), .A2(n1223), .A3(G125), .ZN(n1219) );
INV_X1 U884 ( .A(KEYINPUT1), .ZN(n1222) );
NAND2_X1 U885 ( .A1(G125), .A2(n1223), .ZN(n1218) );
NAND2_X1 U886 ( .A1(KEYINPUT14), .A2(n1168), .ZN(n1223) );
NOR2_X1 U887 ( .A1(n1028), .A2(G952), .ZN(n1136) );
XNOR2_X1 U888 ( .A(G146), .B(n1224), .ZN(G48) );
NAND3_X1 U889 ( .A1(n1049), .A2(n1225), .A3(n1206), .ZN(n1224) );
XOR2_X1 U890 ( .A(KEYINPUT60), .B(n1197), .Z(n1225) );
XOR2_X1 U891 ( .A(G143), .B(n1226), .Z(G45) );
NOR2_X1 U892 ( .A1(n1205), .A2(n1227), .ZN(n1226) );
XOR2_X1 U893 ( .A(KEYINPUT55), .B(n1197), .Z(n1227) );
NAND4_X1 U894 ( .A1(n1214), .A2(n1228), .A3(n1215), .A4(n1229), .ZN(n1205) );
XNOR2_X1 U895 ( .A(G140), .B(n1200), .ZN(G42) );
NAND3_X1 U896 ( .A1(n1230), .A2(n1231), .A3(n1030), .ZN(n1200) );
XNOR2_X1 U897 ( .A(G137), .B(n1201), .ZN(G39) );
NAND3_X1 U898 ( .A1(n1206), .A2(n1030), .A3(n1038), .ZN(n1201) );
XNOR2_X1 U899 ( .A(G134), .B(n1232), .ZN(G36) );
NOR2_X1 U900 ( .A1(n1233), .A2(KEYINPUT34), .ZN(n1232) );
INV_X1 U901 ( .A(n1212), .ZN(n1233) );
NAND4_X1 U902 ( .A1(n1030), .A2(n1214), .A3(n1196), .A4(n1215), .ZN(n1212) );
XNOR2_X1 U903 ( .A(G131), .B(n1234), .ZN(G33) );
NAND4_X1 U904 ( .A1(n1235), .A2(n1030), .A3(n1214), .A4(n1049), .ZN(n1234) );
NOR2_X1 U905 ( .A1(n1044), .A2(n1060), .ZN(n1214) );
NOR2_X1 U906 ( .A1(n1236), .A2(n1067), .ZN(n1030) );
XOR2_X1 U907 ( .A(n1215), .B(KEYINPUT39), .Z(n1235) );
XNOR2_X1 U908 ( .A(G128), .B(n1237), .ZN(G30) );
NAND2_X1 U909 ( .A1(n1217), .A2(n1197), .ZN(n1237) );
AND2_X1 U910 ( .A1(n1206), .A2(n1196), .ZN(n1217) );
INV_X1 U911 ( .A(n1055), .ZN(n1196) );
AND4_X1 U912 ( .A1(n1238), .A2(n1239), .A3(n1231), .A4(n1215), .ZN(n1206) );
XNOR2_X1 U913 ( .A(G101), .B(n1207), .ZN(G3) );
NAND3_X1 U914 ( .A1(n1193), .A2(n1209), .A3(n1038), .ZN(n1207) );
XNOR2_X1 U915 ( .A(G125), .B(n1213), .ZN(G27) );
NAND3_X1 U916 ( .A1(n1230), .A2(n1197), .A3(n1031), .ZN(n1213) );
AND3_X1 U917 ( .A1(n1036), .A2(n1215), .A3(n1049), .ZN(n1230) );
NAND2_X1 U918 ( .A1(n1035), .A2(n1240), .ZN(n1215) );
NAND4_X1 U919 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1106), .ZN(n1240) );
INV_X1 U920 ( .A(G900), .ZN(n1106) );
XNOR2_X1 U921 ( .A(G122), .B(n1191), .ZN(G24) );
NAND4_X1 U922 ( .A1(n1031), .A2(n1046), .A3(n1242), .A4(n1194), .ZN(n1191) );
AND2_X1 U923 ( .A1(n1229), .A2(n1228), .ZN(n1242) );
NOR2_X1 U924 ( .A1(n1238), .A2(n1239), .ZN(n1046) );
XOR2_X1 U925 ( .A(G119), .B(n1243), .Z(G21) );
NOR2_X1 U926 ( .A1(n1065), .A2(n1199), .ZN(n1243) );
NAND3_X1 U927 ( .A1(n1238), .A2(n1038), .A3(n1244), .ZN(n1199) );
NOR3_X1 U928 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
XOR2_X1 U929 ( .A(n1248), .B(n1249), .Z(G18) );
NOR4_X1 U930 ( .A1(n1250), .A2(n1055), .A3(n1245), .A4(n1251), .ZN(n1249) );
XOR2_X1 U931 ( .A(KEYINPUT24), .B(n1193), .Z(n1251) );
INV_X1 U932 ( .A(n1031), .ZN(n1245) );
NAND2_X1 U933 ( .A1(n1252), .A2(n1228), .ZN(n1055) );
NAND2_X1 U934 ( .A1(KEYINPUT59), .A2(n1253), .ZN(n1248) );
INV_X1 U935 ( .A(G116), .ZN(n1253) );
XNOR2_X1 U936 ( .A(G113), .B(n1254), .ZN(G15) );
NAND4_X1 U937 ( .A1(n1193), .A2(n1049), .A3(n1194), .A4(n1255), .ZN(n1254) );
XOR2_X1 U938 ( .A(KEYINPUT27), .B(n1031), .Z(n1255) );
NOR2_X1 U939 ( .A1(n1256), .A2(n1062), .ZN(n1031) );
NOR2_X1 U940 ( .A1(n1228), .A2(n1252), .ZN(n1049) );
INV_X1 U941 ( .A(n1229), .ZN(n1252) );
INV_X1 U942 ( .A(n1044), .ZN(n1193) );
NAND2_X1 U943 ( .A1(n1238), .A2(n1247), .ZN(n1044) );
XNOR2_X1 U944 ( .A(n1208), .B(n1257), .ZN(G12) );
NOR2_X1 U945 ( .A1(KEYINPUT31), .A2(n1181), .ZN(n1257) );
INV_X1 U946 ( .A(G110), .ZN(n1181) );
NAND3_X1 U947 ( .A1(n1036), .A2(n1209), .A3(n1038), .ZN(n1208) );
NOR2_X1 U948 ( .A1(n1228), .A2(n1229), .ZN(n1038) );
NAND2_X1 U949 ( .A1(n1258), .A2(n1081), .ZN(n1229) );
NAND2_X1 U950 ( .A1(n1100), .A2(n1151), .ZN(n1081) );
OR2_X1 U951 ( .A1(n1151), .A2(n1100), .ZN(n1258) );
NOR2_X1 U952 ( .A1(n1150), .A2(G902), .ZN(n1100) );
XNOR2_X1 U953 ( .A(n1259), .B(n1260), .ZN(n1150) );
XOR2_X1 U954 ( .A(G122), .B(G104), .Z(n1260) );
XOR2_X1 U955 ( .A(n1261), .B(n1262), .Z(n1259) );
NOR2_X1 U956 ( .A1(G113), .A2(KEYINPUT28), .ZN(n1262) );
NAND3_X1 U957 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1261) );
NAND2_X1 U958 ( .A1(KEYINPUT33), .A2(n1266), .ZN(n1265) );
OR3_X1 U959 ( .A1(n1266), .A2(KEYINPUT33), .A3(n1267), .ZN(n1264) );
NAND2_X1 U960 ( .A1(n1267), .A2(n1268), .ZN(n1263) );
NAND2_X1 U961 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
INV_X1 U962 ( .A(KEYINPUT33), .ZN(n1270) );
XOR2_X1 U963 ( .A(KEYINPUT7), .B(n1266), .Z(n1269) );
XNOR2_X1 U964 ( .A(n1271), .B(G131), .ZN(n1266) );
NAND2_X1 U965 ( .A1(n1272), .A2(KEYINPUT45), .ZN(n1271) );
XOR2_X1 U966 ( .A(n1273), .B(G143), .Z(n1272) );
NAND3_X1 U967 ( .A1(n1274), .A2(n1028), .A3(G214), .ZN(n1273) );
XOR2_X1 U968 ( .A(KEYINPUT17), .B(G237), .Z(n1274) );
XNOR2_X1 U969 ( .A(n1275), .B(G125), .ZN(n1267) );
INV_X1 U970 ( .A(G475), .ZN(n1151) );
XOR2_X1 U971 ( .A(n1086), .B(G478), .Z(n1228) );
AND2_X1 U972 ( .A1(n1146), .A2(n1078), .ZN(n1086) );
NAND3_X1 U973 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1146) );
OR2_X1 U974 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U975 ( .A1(KEYINPUT26), .A2(n1281), .ZN(n1277) );
NAND2_X1 U976 ( .A1(n1280), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U977 ( .A(KEYINPUT48), .B(n1279), .ZN(n1282) );
NAND2_X1 U978 ( .A1(n1283), .A2(n1284), .ZN(n1276) );
INV_X1 U979 ( .A(KEYINPUT26), .ZN(n1284) );
NAND2_X1 U980 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
OR2_X1 U981 ( .A1(n1279), .A2(KEYINPUT48), .ZN(n1286) );
NAND3_X1 U982 ( .A1(n1280), .A2(n1279), .A3(KEYINPUT48), .ZN(n1285) );
OR2_X1 U983 ( .A1(n1141), .A2(n1287), .ZN(n1279) );
INV_X1 U984 ( .A(G217), .ZN(n1141) );
XOR2_X1 U985 ( .A(n1288), .B(n1289), .Z(n1280) );
XOR2_X1 U986 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U987 ( .A(G116), .B(G107), .Z(n1291) );
NOR2_X1 U988 ( .A1(G143), .A2(KEYINPUT44), .ZN(n1290) );
XNOR2_X1 U989 ( .A(G122), .B(n1292), .ZN(n1288) );
XOR2_X1 U990 ( .A(G134), .B(G128), .Z(n1292) );
NOR2_X1 U991 ( .A1(n1250), .A2(n1060), .ZN(n1209) );
INV_X1 U992 ( .A(n1231), .ZN(n1060) );
NOR2_X1 U993 ( .A1(n1062), .A2(n1063), .ZN(n1231) );
INV_X1 U994 ( .A(n1256), .ZN(n1063) );
NAND2_X1 U995 ( .A1(n1293), .A2(n1080), .ZN(n1256) );
NAND3_X1 U996 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1080) );
INV_X1 U997 ( .A(G469), .ZN(n1077) );
NAND2_X1 U998 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NAND2_X1 U999 ( .A1(n1079), .A2(n1078), .ZN(n1295) );
XOR2_X1 U1000 ( .A(n1296), .B(n1297), .Z(n1079) );
XNOR2_X1 U1001 ( .A(n1173), .B(n1116), .ZN(n1296) );
XNOR2_X1 U1002 ( .A(n1166), .B(G140), .ZN(n1116) );
XNOR2_X1 U1003 ( .A(n1298), .B(n1299), .ZN(n1173) );
XOR2_X1 U1004 ( .A(KEYINPUT22), .B(n1300), .Z(n1299) );
NOR2_X1 U1005 ( .A1(G953), .A2(n1105), .ZN(n1300) );
INV_X1 U1006 ( .A(G227), .ZN(n1105) );
XNOR2_X1 U1007 ( .A(n1301), .B(n1119), .ZN(n1298) );
XNOR2_X1 U1008 ( .A(n1302), .B(n1303), .ZN(n1119) );
XOR2_X1 U1009 ( .A(n1304), .B(KEYINPUT32), .Z(n1302) );
XOR2_X1 U1010 ( .A(KEYINPUT3), .B(G469), .Z(n1294) );
AND2_X1 U1011 ( .A1(G221), .A2(n1305), .ZN(n1062) );
INV_X1 U1012 ( .A(n1194), .ZN(n1250) );
NOR2_X1 U1013 ( .A1(n1065), .A2(n1246), .ZN(n1194) );
AND2_X1 U1014 ( .A1(n1306), .A2(n1035), .ZN(n1246) );
NAND3_X1 U1015 ( .A1(n1241), .A2(n1028), .A3(G952), .ZN(n1035) );
NAND4_X1 U1016 ( .A1(G953), .A2(G902), .A3(n1241), .A4(n1126), .ZN(n1306) );
INV_X1 U1017 ( .A(G898), .ZN(n1126) );
NAND2_X1 U1018 ( .A1(G234), .A2(G237), .ZN(n1241) );
INV_X1 U1019 ( .A(n1197), .ZN(n1065) );
NOR2_X1 U1020 ( .A1(n1068), .A2(n1067), .ZN(n1197) );
AND2_X1 U1021 ( .A1(G214), .A2(n1307), .ZN(n1067) );
INV_X1 U1022 ( .A(n1236), .ZN(n1068) );
NAND3_X1 U1023 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1236) );
XOR2_X1 U1024 ( .A(KEYINPUT15), .B(n1311), .Z(n1310) );
NOR2_X1 U1025 ( .A1(n1312), .A2(n1094), .ZN(n1311) );
OR2_X1 U1026 ( .A1(n1082), .A2(KEYINPUT51), .ZN(n1309) );
NAND2_X1 U1027 ( .A1(n1312), .A2(n1094), .ZN(n1082) );
INV_X1 U1028 ( .A(n1093), .ZN(n1312) );
NAND3_X1 U1029 ( .A1(n1094), .A2(n1093), .A3(KEYINPUT51), .ZN(n1308) );
NAND2_X1 U1030 ( .A1(n1313), .A2(n1078), .ZN(n1093) );
XOR2_X1 U1031 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1032 ( .A(KEYINPUT5), .B(G125), .Z(n1315) );
XOR2_X1 U1033 ( .A(n1183), .B(n1168), .Z(n1314) );
XOR2_X1 U1034 ( .A(n1129), .B(n1316), .Z(n1183) );
XOR2_X1 U1035 ( .A(n1317), .B(n1318), .Z(n1316) );
NOR2_X1 U1036 ( .A1(KEYINPUT40), .A2(n1128), .ZN(n1318) );
XOR2_X1 U1037 ( .A(n1319), .B(n1320), .Z(n1128) );
XNOR2_X1 U1038 ( .A(G119), .B(KEYINPUT8), .ZN(n1319) );
NOR2_X1 U1039 ( .A1(G953), .A2(n1135), .ZN(n1317) );
INV_X1 U1040 ( .A(G224), .ZN(n1135) );
XOR2_X1 U1041 ( .A(n1321), .B(n1297), .Z(n1129) );
XOR2_X1 U1042 ( .A(G101), .B(G110), .Z(n1297) );
XOR2_X1 U1043 ( .A(n1322), .B(G122), .Z(n1321) );
NAND2_X1 U1044 ( .A1(KEYINPUT35), .A2(n1301), .ZN(n1322) );
XOR2_X1 U1045 ( .A(G107), .B(G104), .Z(n1301) );
NAND2_X1 U1046 ( .A1(G210), .A2(n1307), .ZN(n1094) );
NAND2_X1 U1047 ( .A1(n1323), .A2(n1078), .ZN(n1307) );
NOR2_X1 U1048 ( .A1(n1247), .A2(n1238), .ZN(n1036) );
AND2_X1 U1049 ( .A1(n1324), .A2(n1325), .ZN(n1238) );
NAND2_X1 U1050 ( .A1(n1326), .A2(n1089), .ZN(n1325) );
INV_X1 U1051 ( .A(G472), .ZN(n1089) );
XOR2_X1 U1052 ( .A(n1090), .B(KEYINPUT20), .Z(n1326) );
NAND2_X1 U1053 ( .A1(n1327), .A2(G472), .ZN(n1324) );
XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n1090), .ZN(n1327) );
NAND2_X1 U1055 ( .A1(n1328), .A2(n1078), .ZN(n1090) );
XOR2_X1 U1056 ( .A(n1329), .B(n1330), .Z(n1328) );
INV_X1 U1057 ( .A(n1167), .ZN(n1330) );
XOR2_X1 U1058 ( .A(n1331), .B(n1332), .Z(n1167) );
XOR2_X1 U1059 ( .A(G101), .B(n1333), .Z(n1332) );
NOR2_X1 U1060 ( .A1(KEYINPUT42), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1061 ( .A(G119), .B(KEYINPUT25), .ZN(n1334) );
XOR2_X1 U1062 ( .A(n1335), .B(n1320), .Z(n1331) );
XOR2_X1 U1063 ( .A(G113), .B(G116), .Z(n1320) );
NAND3_X1 U1064 ( .A1(n1323), .A2(n1028), .A3(G210), .ZN(n1335) );
INV_X1 U1065 ( .A(G237), .ZN(n1323) );
NAND2_X1 U1066 ( .A1(n1336), .A2(KEYINPUT46), .ZN(n1329) );
XNOR2_X1 U1067 ( .A(n1337), .B(n1166), .ZN(n1336) );
XNOR2_X1 U1068 ( .A(G131), .B(n1338), .ZN(n1166) );
XOR2_X1 U1069 ( .A(G137), .B(G134), .Z(n1338) );
NAND2_X1 U1070 ( .A1(KEYINPUT41), .A2(n1168), .ZN(n1337) );
INV_X1 U1071 ( .A(n1221), .ZN(n1168) );
XOR2_X1 U1072 ( .A(n1339), .B(n1303), .Z(n1221) );
XOR2_X1 U1073 ( .A(G146), .B(G128), .Z(n1303) );
NAND2_X1 U1074 ( .A1(KEYINPUT30), .A2(n1304), .ZN(n1339) );
INV_X1 U1075 ( .A(G143), .ZN(n1304) );
INV_X1 U1076 ( .A(n1239), .ZN(n1247) );
XNOR2_X1 U1077 ( .A(n1099), .B(n1340), .ZN(n1239) );
NOR2_X1 U1078 ( .A1(n1098), .A2(KEYINPUT58), .ZN(n1340) );
AND2_X1 U1079 ( .A1(n1341), .A2(G217), .ZN(n1098) );
XOR2_X1 U1080 ( .A(n1305), .B(KEYINPUT43), .Z(n1341) );
NAND2_X1 U1081 ( .A1(G234), .A2(n1078), .ZN(n1305) );
INV_X1 U1082 ( .A(G902), .ZN(n1078) );
NOR2_X1 U1083 ( .A1(n1143), .A2(G902), .ZN(n1099) );
XOR2_X1 U1084 ( .A(n1342), .B(n1343), .Z(n1143) );
XOR2_X1 U1085 ( .A(n1344), .B(n1345), .Z(n1343) );
XOR2_X1 U1086 ( .A(G110), .B(n1346), .Z(n1345) );
NOR2_X1 U1087 ( .A1(KEYINPUT62), .A2(n1347), .ZN(n1346) );
XOR2_X1 U1088 ( .A(n1275), .B(n1348), .Z(n1347) );
NOR2_X1 U1089 ( .A1(G125), .A2(KEYINPUT19), .ZN(n1348) );
XNOR2_X1 U1090 ( .A(G140), .B(n1349), .ZN(n1275) );
XOR2_X1 U1091 ( .A(KEYINPUT50), .B(G146), .Z(n1349) );
NOR2_X1 U1092 ( .A1(n1287), .A2(n1350), .ZN(n1344) );
INV_X1 U1093 ( .A(G221), .ZN(n1350) );
NAND2_X1 U1094 ( .A1(G234), .A2(n1028), .ZN(n1287) );
INV_X1 U1095 ( .A(G953), .ZN(n1028) );
XNOR2_X1 U1096 ( .A(G119), .B(n1351), .ZN(n1342) );
XOR2_X1 U1097 ( .A(G137), .B(G128), .Z(n1351) );
endmodule


