//Key = 0000111000011110010001011010000000100010111000000110010010111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;

XNOR2_X1 U740 ( .A(G107), .B(n1027), .ZN(G9) );
NAND3_X1 U741 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(G75) );
NAND2_X1 U742 ( .A1(G952), .A2(n1031), .ZN(n1030) );
NAND3_X1 U743 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NAND4_X1 U744 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1033) );
NAND2_X1 U745 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U747 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1042) );
OR3_X1 U748 ( .A1(n1046), .A2(n1047), .A3(KEYINPUT0), .ZN(n1044) );
NAND2_X1 U749 ( .A1(KEYINPUT0), .A2(n1048), .ZN(n1043) );
NAND2_X1 U750 ( .A1(n1048), .A2(n1049), .ZN(n1039) );
NAND2_X1 U751 ( .A1(n1048), .A2(n1050), .ZN(n1032) );
NAND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U753 ( .A1(n1053), .A2(n1038), .A3(n1041), .ZN(n1052) );
NAND2_X1 U754 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND3_X1 U755 ( .A1(n1056), .A2(n1057), .A3(n1036), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1035), .A2(n1058), .ZN(n1054) );
OR2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U758 ( .A(KEYINPUT34), .B(n1061), .Z(n1051) );
NOR3_X1 U759 ( .A1(n1062), .A2(n1057), .A3(n1056), .ZN(n1061) );
NAND3_X1 U760 ( .A1(n1041), .A2(n1038), .A3(n1036), .ZN(n1062) );
NAND4_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1028) );
NOR4_X1 U762 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
NOR3_X1 U763 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
INV_X1 U764 ( .A(KEYINPUT17), .ZN(n1071) );
NOR2_X1 U765 ( .A1(KEYINPUT17), .A2(n1074), .ZN(n1069) );
XNOR2_X1 U766 ( .A(G478), .B(n1075), .ZN(n1068) );
NAND4_X1 U767 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1067) );
OR2_X1 U768 ( .A1(G475), .A2(KEYINPUT38), .ZN(n1079) );
NAND3_X1 U769 ( .A1(G475), .A2(n1080), .A3(KEYINPUT38), .ZN(n1078) );
OR2_X1 U770 ( .A1(n1035), .A2(KEYINPUT63), .ZN(n1077) );
NAND2_X1 U771 ( .A1(KEYINPUT63), .A2(n1081), .ZN(n1076) );
NAND3_X1 U772 ( .A1(n1082), .A2(n1057), .A3(G469), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1065) );
XNOR2_X1 U774 ( .A(G472), .B(n1085), .ZN(n1083) );
NOR2_X1 U775 ( .A1(n1086), .A2(KEYINPUT35), .ZN(n1085) );
XOR2_X1 U776 ( .A(n1087), .B(n1088), .Z(G72) );
NOR2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR2_X1 U778 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U779 ( .A(KEYINPUT18), .B(n1093), .ZN(n1091) );
NOR2_X1 U780 ( .A1(n1094), .A2(n1093), .ZN(n1089) );
NAND2_X1 U781 ( .A1(n1029), .A2(n1095), .ZN(n1093) );
INV_X1 U782 ( .A(n1092), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
NAND2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U785 ( .A(G953), .B(KEYINPUT59), .ZN(n1098) );
XOR2_X1 U786 ( .A(n1100), .B(n1101), .Z(n1096) );
XNOR2_X1 U787 ( .A(G125), .B(n1102), .ZN(n1101) );
NOR2_X1 U788 ( .A1(KEYINPUT52), .A2(n1103), .ZN(n1102) );
XNOR2_X1 U789 ( .A(n1104), .B(n1105), .ZN(n1103) );
NOR2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR3_X1 U791 ( .A1(KEYINPUT40), .A2(G137), .A3(n1108), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
INV_X1 U793 ( .A(KEYINPUT40), .ZN(n1110) );
NAND2_X1 U794 ( .A1(G953), .A2(n1111), .ZN(n1087) );
NAND2_X1 U795 ( .A1(G900), .A2(G227), .ZN(n1111) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(G69) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U798 ( .A(KEYINPUT19), .B(n1116), .Z(n1115) );
NOR2_X1 U799 ( .A1(n1117), .A2(n1029), .ZN(n1116) );
AND2_X1 U800 ( .A1(G224), .A2(G898), .ZN(n1117) );
NOR2_X1 U801 ( .A1(n1118), .A2(G953), .ZN(n1114) );
NOR3_X1 U802 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
NAND2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(n1112) );
NAND2_X1 U804 ( .A1(G953), .A2(n1124), .ZN(n1123) );
XOR2_X1 U805 ( .A(n1125), .B(n1126), .Z(n1122) );
NAND2_X1 U806 ( .A1(KEYINPUT23), .A2(n1127), .ZN(n1125) );
NOR2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U809 ( .A1(KEYINPUT12), .A2(n1132), .ZN(n1131) );
NAND2_X1 U810 ( .A1(n1133), .A2(n1074), .ZN(n1130) );
INV_X1 U811 ( .A(n1073), .ZN(n1074) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1134), .ZN(G63) );
NOR3_X1 U813 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
NOR3_X1 U814 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
NOR2_X1 U815 ( .A1(n1141), .A2(n1142), .ZN(n1136) );
NOR2_X1 U816 ( .A1(n1034), .A2(n1139), .ZN(n1141) );
NOR2_X1 U817 ( .A1(n1128), .A2(n1143), .ZN(G60) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND3_X1 U819 ( .A1(n1133), .A2(G475), .A3(KEYINPUT42), .ZN(n1144) );
XNOR2_X1 U820 ( .A(G104), .B(n1146), .ZN(G6) );
NOR2_X1 U821 ( .A1(n1128), .A2(n1147), .ZN(G57) );
XNOR2_X1 U822 ( .A(n1148), .B(n1149), .ZN(n1147) );
NOR2_X1 U823 ( .A1(KEYINPUT37), .A2(n1150), .ZN(n1148) );
XNOR2_X1 U824 ( .A(n1151), .B(n1152), .ZN(n1150) );
XOR2_X1 U825 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U826 ( .A1(KEYINPUT25), .A2(n1155), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1156), .A2(n1140), .ZN(n1153) );
NOR2_X1 U828 ( .A1(n1128), .A2(n1157), .ZN(G54) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U830 ( .A(n1100), .B(n1160), .Z(n1159) );
XNOR2_X1 U831 ( .A(n1161), .B(n1162), .ZN(n1160) );
XNOR2_X1 U832 ( .A(n1163), .B(n1164), .ZN(n1100) );
XOR2_X1 U833 ( .A(n1165), .B(n1166), .Z(n1158) );
XOR2_X1 U834 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR3_X1 U835 ( .A1(n1140), .A2(KEYINPUT45), .A3(n1169), .ZN(n1168) );
NAND2_X1 U836 ( .A1(KEYINPUT56), .A2(n1170), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1128), .A2(n1171), .ZN(G51) );
XOR2_X1 U838 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U839 ( .A(n1155), .B(n1174), .Z(n1173) );
XOR2_X1 U840 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U841 ( .A1(n1177), .A2(n1140), .ZN(n1176) );
INV_X1 U842 ( .A(n1133), .ZN(n1140) );
NOR2_X1 U843 ( .A1(n1178), .A2(n1034), .ZN(n1133) );
NOR4_X1 U844 ( .A1(n1179), .A2(n1119), .A3(n1095), .A4(n1120), .ZN(n1034) );
AND4_X1 U845 ( .A1(n1180), .A2(n1035), .A3(n1181), .A4(n1041), .ZN(n1120) );
NOR2_X1 U846 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U847 ( .A(n1184), .B(KEYINPUT30), .ZN(n1183) );
INV_X1 U848 ( .A(n1185), .ZN(n1182) );
XNOR2_X1 U849 ( .A(n1186), .B(KEYINPUT50), .ZN(n1180) );
NAND4_X1 U850 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1095) );
NOR4_X1 U851 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190) );
NOR2_X1 U852 ( .A1(n1195), .A2(n1196), .ZN(n1189) );
NAND3_X1 U853 ( .A1(n1197), .A2(n1059), .A3(n1198), .ZN(n1187) );
XNOR2_X1 U854 ( .A(KEYINPUT47), .B(n1084), .ZN(n1197) );
NAND3_X1 U855 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1119) );
XNOR2_X1 U856 ( .A(n1121), .B(KEYINPUT60), .ZN(n1179) );
NAND3_X1 U857 ( .A1(n1146), .A2(n1027), .A3(n1202), .ZN(n1121) );
NAND3_X1 U858 ( .A1(n1184), .A2(n1049), .A3(n1203), .ZN(n1202) );
INV_X1 U859 ( .A(n1204), .ZN(n1203) );
NAND2_X1 U860 ( .A1(n1205), .A2(n1206), .ZN(n1049) );
NAND2_X1 U861 ( .A1(n1207), .A2(n1059), .ZN(n1027) );
NAND2_X1 U862 ( .A1(n1060), .A2(n1207), .ZN(n1146) );
AND3_X1 U863 ( .A1(n1041), .A2(n1184), .A3(n1208), .ZN(n1207) );
NAND2_X1 U864 ( .A1(KEYINPUT21), .A2(n1209), .ZN(n1175) );
XOR2_X1 U865 ( .A(n1210), .B(n1211), .Z(n1172) );
XNOR2_X1 U866 ( .A(KEYINPUT55), .B(n1212), .ZN(n1211) );
NOR2_X1 U867 ( .A1(n1029), .A2(G952), .ZN(n1128) );
XNOR2_X1 U868 ( .A(n1213), .B(n1214), .ZN(G48) );
NOR2_X1 U869 ( .A1(KEYINPUT27), .A2(n1188), .ZN(n1214) );
NAND3_X1 U870 ( .A1(n1060), .A2(n1184), .A3(n1215), .ZN(n1188) );
XOR2_X1 U871 ( .A(G143), .B(n1193), .Z(G45) );
AND3_X1 U872 ( .A1(n1186), .A2(n1184), .A3(n1198), .ZN(n1193) );
XOR2_X1 U873 ( .A(n1192), .B(n1216), .Z(G42) );
NOR2_X1 U874 ( .A1(KEYINPUT32), .A2(n1164), .ZN(n1216) );
INV_X1 U875 ( .A(G140), .ZN(n1164) );
AND4_X1 U876 ( .A1(n1217), .A2(n1218), .A3(n1060), .A4(n1048), .ZN(n1192) );
XOR2_X1 U877 ( .A(G137), .B(n1196), .Z(G39) );
AND3_X1 U878 ( .A1(n1048), .A2(n1036), .A3(n1215), .ZN(n1196) );
XNOR2_X1 U879 ( .A(G134), .B(n1219), .ZN(G36) );
NAND4_X1 U880 ( .A1(n1220), .A2(n1218), .A3(n1048), .A4(n1059), .ZN(n1219) );
XNOR2_X1 U881 ( .A(n1221), .B(KEYINPUT53), .ZN(n1220) );
XNOR2_X1 U882 ( .A(n1104), .B(n1191), .ZN(G33) );
AND3_X1 U883 ( .A1(n1060), .A2(n1048), .A3(n1198), .ZN(n1191) );
AND2_X1 U884 ( .A1(n1218), .A2(n1221), .ZN(n1198) );
INV_X1 U885 ( .A(n1084), .ZN(n1048) );
NAND2_X1 U886 ( .A1(n1222), .A2(n1046), .ZN(n1084) );
XOR2_X1 U887 ( .A(G128), .B(n1195), .Z(G30) );
AND3_X1 U888 ( .A1(n1184), .A2(n1059), .A3(n1215), .ZN(n1195) );
AND3_X1 U889 ( .A1(n1223), .A2(n1224), .A3(n1218), .ZN(n1215) );
AND3_X1 U890 ( .A1(n1225), .A2(n1057), .A3(n1056), .ZN(n1218) );
NAND2_X1 U891 ( .A1(KEYINPUT39), .A2(n1205), .ZN(n1224) );
NAND2_X1 U892 ( .A1(n1226), .A2(n1227), .ZN(n1223) );
INV_X1 U893 ( .A(KEYINPUT39), .ZN(n1227) );
NAND2_X1 U894 ( .A1(n1228), .A2(n1229), .ZN(n1226) );
XNOR2_X1 U895 ( .A(G101), .B(n1230), .ZN(G3) );
NAND2_X1 U896 ( .A1(n1184), .A2(n1231), .ZN(n1230) );
XOR2_X1 U897 ( .A(KEYINPUT16), .B(n1232), .Z(n1231) );
NOR2_X1 U898 ( .A1(n1206), .A2(n1204), .ZN(n1232) );
INV_X1 U899 ( .A(n1221), .ZN(n1206) );
NAND2_X1 U900 ( .A1(n1233), .A2(n1234), .ZN(G27) );
NAND2_X1 U901 ( .A1(n1194), .A2(n1212), .ZN(n1234) );
INV_X1 U902 ( .A(n1235), .ZN(n1194) );
XOR2_X1 U903 ( .A(n1236), .B(KEYINPUT22), .Z(n1233) );
NAND2_X1 U904 ( .A1(G125), .A2(n1235), .ZN(n1236) );
NAND4_X1 U905 ( .A1(n1217), .A2(n1060), .A3(n1237), .A4(n1035), .ZN(n1235) );
AND2_X1 U906 ( .A1(n1225), .A2(n1184), .ZN(n1237) );
NAND2_X1 U907 ( .A1(n1238), .A2(n1239), .ZN(n1225) );
NAND4_X1 U908 ( .A1(G953), .A2(G902), .A3(n1038), .A4(n1099), .ZN(n1239) );
INV_X1 U909 ( .A(G900), .ZN(n1099) );
INV_X1 U910 ( .A(n1205), .ZN(n1217) );
XNOR2_X1 U911 ( .A(G122), .B(n1240), .ZN(G24) );
NAND3_X1 U912 ( .A1(n1186), .A2(n1041), .A3(n1241), .ZN(n1240) );
NOR2_X1 U913 ( .A1(n1229), .A2(n1228), .ZN(n1041) );
AND2_X1 U914 ( .A1(n1242), .A2(n1243), .ZN(n1186) );
XNOR2_X1 U915 ( .A(n1244), .B(n1245), .ZN(n1242) );
XNOR2_X1 U916 ( .A(G119), .B(n1201), .ZN(G21) );
NAND4_X1 U917 ( .A1(n1241), .A2(n1036), .A3(n1246), .A4(n1229), .ZN(n1201) );
XNOR2_X1 U918 ( .A(KEYINPUT39), .B(n1247), .ZN(n1246) );
XNOR2_X1 U919 ( .A(G116), .B(n1199), .ZN(G18) );
NAND3_X1 U920 ( .A1(n1221), .A2(n1059), .A3(n1241), .ZN(n1199) );
NAND2_X1 U921 ( .A1(n1248), .A2(n1249), .ZN(n1059) );
NAND2_X1 U922 ( .A1(n1036), .A2(n1244), .ZN(n1249) );
OR3_X1 U923 ( .A1(n1243), .A2(n1245), .A3(n1244), .ZN(n1248) );
INV_X1 U924 ( .A(KEYINPUT14), .ZN(n1244) );
XOR2_X1 U925 ( .A(n1200), .B(n1250), .Z(G15) );
NOR2_X1 U926 ( .A1(G113), .A2(KEYINPUT51), .ZN(n1250) );
NAND3_X1 U927 ( .A1(n1060), .A2(n1221), .A3(n1241), .ZN(n1200) );
AND3_X1 U928 ( .A1(n1184), .A2(n1185), .A3(n1035), .ZN(n1241) );
NOR2_X1 U929 ( .A1(n1056), .A2(n1251), .ZN(n1035) );
INV_X1 U930 ( .A(n1057), .ZN(n1251) );
NOR2_X1 U931 ( .A1(n1229), .A2(n1252), .ZN(n1221) );
XNOR2_X1 U932 ( .A(KEYINPUT57), .B(n1228), .ZN(n1252) );
INV_X1 U933 ( .A(n1247), .ZN(n1228) );
AND2_X1 U934 ( .A1(n1253), .A2(n1245), .ZN(n1060) );
XOR2_X1 U935 ( .A(n1243), .B(KEYINPUT10), .Z(n1253) );
XNOR2_X1 U936 ( .A(G110), .B(n1254), .ZN(G12) );
NOR2_X1 U937 ( .A1(KEYINPUT43), .A2(n1255), .ZN(n1254) );
NOR3_X1 U938 ( .A1(n1204), .A2(n1256), .A3(n1205), .ZN(n1255) );
NAND2_X1 U939 ( .A1(n1247), .A2(n1229), .ZN(n1205) );
NAND2_X1 U940 ( .A1(n1257), .A2(n1064), .ZN(n1229) );
NAND2_X1 U941 ( .A1(n1072), .A2(n1073), .ZN(n1064) );
OR2_X1 U942 ( .A1(n1073), .A2(n1072), .ZN(n1257) );
NOR2_X1 U943 ( .A1(G902), .A2(n1132), .ZN(n1072) );
AND2_X1 U944 ( .A1(n1258), .A2(n1259), .ZN(n1132) );
NAND2_X1 U945 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
XOR2_X1 U946 ( .A(n1262), .B(KEYINPUT33), .Z(n1258) );
OR2_X1 U947 ( .A1(n1261), .A2(n1260), .ZN(n1262) );
XOR2_X1 U948 ( .A(n1263), .B(n1264), .Z(n1260) );
XNOR2_X1 U949 ( .A(n1170), .B(n1265), .ZN(n1264) );
XNOR2_X1 U950 ( .A(KEYINPUT49), .B(n1212), .ZN(n1265) );
XOR2_X1 U951 ( .A(n1266), .B(n1267), .Z(n1263) );
NAND2_X1 U952 ( .A1(n1268), .A2(n1269), .ZN(n1266) );
OR2_X1 U953 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XOR2_X1 U954 ( .A(n1272), .B(KEYINPUT48), .Z(n1268) );
NAND2_X1 U955 ( .A1(n1271), .A2(n1270), .ZN(n1272) );
XOR2_X1 U956 ( .A(G128), .B(KEYINPUT44), .Z(n1271) );
XNOR2_X1 U957 ( .A(n1273), .B(G137), .ZN(n1261) );
NAND2_X1 U958 ( .A1(n1274), .A2(G221), .ZN(n1273) );
NAND2_X1 U959 ( .A1(G217), .A2(n1275), .ZN(n1073) );
XOR2_X1 U960 ( .A(n1086), .B(n1156), .Z(n1247) );
INV_X1 U961 ( .A(G472), .ZN(n1156) );
AND2_X1 U962 ( .A1(n1276), .A2(n1178), .ZN(n1086) );
XNOR2_X1 U963 ( .A(n1277), .B(n1278), .ZN(n1276) );
INV_X1 U964 ( .A(n1151), .ZN(n1278) );
XOR2_X1 U965 ( .A(n1109), .B(n1279), .Z(n1151) );
XOR2_X1 U966 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U967 ( .A(n1282), .B(n1283), .ZN(n1277) );
NOR2_X1 U968 ( .A1(KEYINPUT8), .A2(n1155), .ZN(n1283) );
NOR2_X1 U969 ( .A1(KEYINPUT2), .A2(n1149), .ZN(n1282) );
XOR2_X1 U970 ( .A(n1284), .B(G101), .Z(n1149) );
NAND2_X1 U971 ( .A1(G210), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U972 ( .A(n1184), .B(KEYINPUT9), .ZN(n1256) );
INV_X1 U973 ( .A(n1045), .ZN(n1184) );
NAND2_X1 U974 ( .A1(n1047), .A2(n1046), .ZN(n1045) );
NAND2_X1 U975 ( .A1(G214), .A2(n1286), .ZN(n1046) );
INV_X1 U976 ( .A(n1222), .ZN(n1047) );
XNOR2_X1 U977 ( .A(n1287), .B(n1177), .ZN(n1222) );
NAND2_X1 U978 ( .A1(G210), .A2(n1286), .ZN(n1177) );
NAND2_X1 U979 ( .A1(n1288), .A2(n1178), .ZN(n1286) );
INV_X1 U980 ( .A(G237), .ZN(n1288) );
NAND2_X1 U981 ( .A1(n1289), .A2(n1178), .ZN(n1287) );
XOR2_X1 U982 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U983 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U984 ( .A(n1210), .B(KEYINPUT1), .Z(n1293) );
NAND2_X1 U985 ( .A1(G224), .A2(n1029), .ZN(n1210) );
NAND2_X1 U986 ( .A1(KEYINPUT6), .A2(n1212), .ZN(n1292) );
XOR2_X1 U987 ( .A(n1209), .B(n1155), .Z(n1290) );
XNOR2_X1 U988 ( .A(n1294), .B(n1213), .ZN(n1155) );
XNOR2_X1 U989 ( .A(n1126), .B(n1127), .ZN(n1209) );
XNOR2_X1 U990 ( .A(n1170), .B(G122), .ZN(n1127) );
XOR2_X1 U991 ( .A(n1295), .B(n1296), .Z(n1126) );
XNOR2_X1 U992 ( .A(G101), .B(n1297), .ZN(n1296) );
NAND2_X1 U993 ( .A1(KEYINPUT62), .A2(n1298), .ZN(n1297) );
XOR2_X1 U994 ( .A(KEYINPUT29), .B(n1299), .Z(n1298) );
NAND2_X1 U995 ( .A1(n1300), .A2(n1301), .ZN(n1295) );
NAND2_X1 U996 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
INV_X1 U997 ( .A(KEYINPUT61), .ZN(n1303) );
XOR2_X1 U998 ( .A(G113), .B(n1281), .Z(n1302) );
NAND3_X1 U999 ( .A1(G113), .A2(n1281), .A3(KEYINPUT61), .ZN(n1300) );
XNOR2_X1 U1000 ( .A(G116), .B(n1270), .ZN(n1281) );
INV_X1 U1001 ( .A(G119), .ZN(n1270) );
NAND2_X1 U1002 ( .A1(n1036), .A2(n1208), .ZN(n1204) );
AND3_X1 U1003 ( .A1(n1185), .A2(n1057), .A3(n1056), .ZN(n1208) );
XOR2_X1 U1004 ( .A(n1082), .B(n1169), .Z(n1056) );
INV_X1 U1005 ( .A(G469), .ZN(n1169) );
NAND2_X1 U1006 ( .A1(n1304), .A2(n1178), .ZN(n1082) );
XOR2_X1 U1007 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U1008 ( .A(n1163), .B(n1307), .Z(n1306) );
XNOR2_X1 U1009 ( .A(n1308), .B(n1167), .ZN(n1307) );
NAND2_X1 U1010 ( .A1(n1309), .A2(G227), .ZN(n1167) );
XNOR2_X1 U1011 ( .A(G953), .B(KEYINPUT28), .ZN(n1309) );
NAND2_X1 U1012 ( .A1(KEYINPUT58), .A2(n1161), .ZN(n1308) );
XOR2_X1 U1013 ( .A(G131), .B(n1109), .Z(n1161) );
XNOR2_X1 U1014 ( .A(n1108), .B(G137), .ZN(n1109) );
NAND2_X1 U1015 ( .A1(n1310), .A2(n1311), .ZN(n1163) );
NAND2_X1 U1016 ( .A1(G146), .A2(n1294), .ZN(n1311) );
NAND2_X1 U1017 ( .A1(n1312), .A2(n1213), .ZN(n1310) );
INV_X1 U1018 ( .A(G146), .ZN(n1213) );
XOR2_X1 U1019 ( .A(n1294), .B(KEYINPUT4), .Z(n1312) );
XNOR2_X1 U1020 ( .A(G128), .B(n1313), .ZN(n1294) );
XOR2_X1 U1021 ( .A(KEYINPUT26), .B(G143), .Z(n1313) );
XOR2_X1 U1022 ( .A(n1314), .B(n1315), .Z(n1305) );
XNOR2_X1 U1023 ( .A(n1170), .B(n1316), .ZN(n1315) );
NOR2_X1 U1024 ( .A1(KEYINPUT36), .A2(G140), .ZN(n1316) );
INV_X1 U1025 ( .A(G110), .ZN(n1170) );
NOR2_X1 U1026 ( .A1(KEYINPUT20), .A2(n1162), .ZN(n1314) );
XNOR2_X1 U1027 ( .A(n1317), .B(n1299), .ZN(n1162) );
XOR2_X1 U1028 ( .A(G104), .B(G107), .Z(n1299) );
INV_X1 U1029 ( .A(G101), .ZN(n1317) );
NAND2_X1 U1030 ( .A1(n1318), .A2(G221), .ZN(n1057) );
XOR2_X1 U1031 ( .A(n1275), .B(KEYINPUT54), .Z(n1318) );
NAND2_X1 U1032 ( .A1(G234), .A2(n1178), .ZN(n1275) );
NAND2_X1 U1033 ( .A1(n1238), .A2(n1319), .ZN(n1185) );
NAND4_X1 U1034 ( .A1(n1320), .A2(G953), .A3(G902), .A4(n1124), .ZN(n1319) );
INV_X1 U1035 ( .A(G898), .ZN(n1124) );
XOR2_X1 U1036 ( .A(n1038), .B(KEYINPUT3), .Z(n1320) );
NAND3_X1 U1037 ( .A1(G952), .A2(n1029), .A3(n1321), .ZN(n1238) );
XOR2_X1 U1038 ( .A(n1038), .B(KEYINPUT7), .Z(n1321) );
NAND2_X1 U1039 ( .A1(n1322), .A2(G234), .ZN(n1038) );
XNOR2_X1 U1040 ( .A(G237), .B(KEYINPUT5), .ZN(n1322) );
NOR2_X1 U1041 ( .A1(n1243), .A2(n1323), .ZN(n1036) );
INV_X1 U1042 ( .A(n1245), .ZN(n1323) );
XOR2_X1 U1043 ( .A(n1324), .B(n1075), .Z(n1245) );
INV_X1 U1044 ( .A(n1135), .ZN(n1075) );
NOR2_X1 U1045 ( .A1(n1142), .A2(G902), .ZN(n1135) );
INV_X1 U1046 ( .A(n1138), .ZN(n1142) );
XNOR2_X1 U1047 ( .A(n1325), .B(n1326), .ZN(n1138) );
XOR2_X1 U1048 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1049 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U1050 ( .A1(KEYINPUT31), .A2(n1331), .ZN(n1330) );
XNOR2_X1 U1051 ( .A(G107), .B(KEYINPUT13), .ZN(n1331) );
NAND2_X1 U1052 ( .A1(n1332), .A2(KEYINPUT41), .ZN(n1329) );
XNOR2_X1 U1053 ( .A(G128), .B(G143), .ZN(n1332) );
AND2_X1 U1054 ( .A1(G217), .A2(n1274), .ZN(n1327) );
AND2_X1 U1055 ( .A1(G234), .A2(n1029), .ZN(n1274) );
INV_X1 U1056 ( .A(G953), .ZN(n1029) );
XNOR2_X1 U1057 ( .A(G116), .B(n1333), .ZN(n1325) );
XNOR2_X1 U1058 ( .A(n1108), .B(G122), .ZN(n1333) );
INV_X1 U1059 ( .A(G134), .ZN(n1108) );
NAND2_X1 U1060 ( .A1(KEYINPUT24), .A2(n1139), .ZN(n1324) );
INV_X1 U1061 ( .A(G478), .ZN(n1139) );
NAND3_X1 U1062 ( .A1(n1334), .A2(n1335), .A3(n1063), .ZN(n1243) );
NAND2_X1 U1063 ( .A1(n1336), .A2(n1337), .ZN(n1063) );
OR3_X1 U1064 ( .A1(n1337), .A2(n1336), .A3(KEYINPUT46), .ZN(n1335) );
INV_X1 U1065 ( .A(G475), .ZN(n1337) );
NAND2_X1 U1066 ( .A1(KEYINPUT46), .A2(n1336), .ZN(n1334) );
INV_X1 U1067 ( .A(n1080), .ZN(n1336) );
NAND2_X1 U1068 ( .A1(n1145), .A2(n1178), .ZN(n1080) );
INV_X1 U1069 ( .A(G902), .ZN(n1178) );
XOR2_X1 U1070 ( .A(n1338), .B(n1339), .Z(n1145) );
XNOR2_X1 U1071 ( .A(n1280), .B(n1340), .ZN(n1339) );
XNOR2_X1 U1072 ( .A(n1267), .B(n1341), .ZN(n1340) );
AND3_X1 U1073 ( .A1(G214), .A2(n1342), .A3(n1285), .ZN(n1341) );
NOR2_X1 U1074 ( .A1(G953), .A2(G237), .ZN(n1285) );
INV_X1 U1075 ( .A(KEYINPUT15), .ZN(n1342) );
XOR2_X1 U1076 ( .A(G140), .B(G146), .Z(n1267) );
XNOR2_X1 U1077 ( .A(G113), .B(n1104), .ZN(n1280) );
INV_X1 U1078 ( .A(G131), .ZN(n1104) );
XOR2_X1 U1079 ( .A(n1343), .B(n1344), .Z(n1338) );
XOR2_X1 U1080 ( .A(G143), .B(G122), .Z(n1344) );
XOR2_X1 U1081 ( .A(n1345), .B(G104), .Z(n1343) );
NAND2_X1 U1082 ( .A1(KEYINPUT11), .A2(n1212), .ZN(n1345) );
INV_X1 U1083 ( .A(G125), .ZN(n1212) );
endmodule


