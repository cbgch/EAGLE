//Key = 1010100000010111001111001010101101101111110100000000001100000001


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185;

OR2_X1 U1232 ( .A1(n1703), .A2(STATO_REG_0__SCAN_IN), .ZN(n1647) );
INV_X2 U1233 ( .A(n1647), .ZN(n1648) );
INV_X2 U1234 ( .A(U280), .ZN(n1800) );
NAND2_X1 U1235 ( .A1(n1649), .A2(n1650), .ZN(U344) );
NAND2_X1 U1236 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1651), .ZN(n1650) );
NAND2_X1 U1237 ( .A1(n1652), .A2(DATA_IN_7_), .ZN(n1649) );
NAND2_X1 U1238 ( .A1(n1653), .A2(n1654), .ZN(U343) );
NAND2_X1 U1239 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1651), .ZN(n1654) );
NAND2_X1 U1240 ( .A1(n1652), .A2(DATA_IN_6_), .ZN(n1653) );
NAND2_X1 U1241 ( .A1(n1655), .A2(n1656), .ZN(U342) );
NAND2_X1 U1242 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1651), .ZN(n1656) );
NAND2_X1 U1243 ( .A1(n1652), .A2(DATA_IN_5_), .ZN(n1655) );
NAND2_X1 U1244 ( .A1(n1657), .A2(n1658), .ZN(U341) );
NAND2_X1 U1245 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1651), .ZN(n1658) );
NAND2_X1 U1246 ( .A1(n1652), .A2(DATA_IN_4_), .ZN(n1657) );
NAND2_X1 U1247 ( .A1(n1659), .A2(n1660), .ZN(U340) );
NAND2_X1 U1248 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1651), .ZN(n1660) );
NAND2_X1 U1249 ( .A1(n1652), .A2(DATA_IN_3_), .ZN(n1659) );
NAND3_X1 U1250 ( .A1(n1661), .A2(n1662), .A3(n1663), .ZN(U339) );
NAND2_X1 U1251 ( .A1(KEYINPUT6), .A2(n1664), .ZN(n1663) );
NAND3_X1 U1252 ( .A1(DATA_IN_2_), .A2(n1665), .A3(n1652), .ZN(n1662) );
NAND2_X1 U1253 ( .A1(n1666), .A2(n1651), .ZN(n1661) );
NAND2_X1 U1254 ( .A1(n1667), .A2(n1665), .ZN(n1666) );
INV_X1 U1255 ( .A(KEYINPUT6), .ZN(n1665) );
XNOR2_X1 U1256 ( .A(RMAX_REG_2__SCAN_IN), .B(KEYINPUT8), .ZN(n1667) );
NAND2_X1 U1257 ( .A1(n1668), .A2(n1669), .ZN(U338) );
NAND2_X1 U1258 ( .A1(n1670), .A2(RMAX_REG_1__SCAN_IN), .ZN(n1669) );
XNOR2_X1 U1259 ( .A(n1652), .B(KEYINPUT44), .ZN(n1670) );
NAND2_X1 U1260 ( .A1(n1652), .A2(DATA_IN_1_), .ZN(n1668) );
NAND2_X1 U1261 ( .A1(n1671), .A2(n1672), .ZN(U337) );
NAND2_X1 U1262 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1651), .ZN(n1672) );
NAND2_X1 U1263 ( .A1(n1652), .A2(DATA_IN_0_), .ZN(n1671) );
INV_X1 U1264 ( .A(n1651), .ZN(n1652) );
NAND2_X1 U1265 ( .A1(n1673), .A2(n1674), .ZN(n1651) );
NAND3_X1 U1266 ( .A1(n1675), .A2(n1676), .A3(n1677), .ZN(n1674) );
NAND2_X1 U1267 ( .A1(n1678), .A2(n1679), .ZN(U336) );
NAND2_X1 U1268 ( .A1(n1680), .A2(RMIN_REG_7__SCAN_IN), .ZN(n1679) );
XOR2_X1 U1269 ( .A(n1681), .B(KEYINPUT50), .Z(n1680) );
NAND2_X1 U1270 ( .A1(DATA_IN_7_), .A2(n1682), .ZN(n1678) );
NAND2_X1 U1271 ( .A1(n1683), .A2(n1684), .ZN(U335) );
NAND2_X1 U1272 ( .A1(DATA_IN_6_), .A2(n1682), .ZN(n1684) );
NAND2_X1 U1273 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1681), .ZN(n1683) );
NAND2_X1 U1274 ( .A1(n1685), .A2(n1686), .ZN(U334) );
NAND2_X1 U1275 ( .A1(DATA_IN_5_), .A2(n1682), .ZN(n1686) );
NAND2_X1 U1276 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1681), .ZN(n1685) );
NAND2_X1 U1277 ( .A1(n1687), .A2(n1688), .ZN(U333) );
NAND2_X1 U1278 ( .A1(DATA_IN_4_), .A2(n1682), .ZN(n1688) );
NAND2_X1 U1279 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1681), .ZN(n1687) );
NAND2_X1 U1280 ( .A1(n1689), .A2(n1690), .ZN(U332) );
NAND2_X1 U1281 ( .A1(n1691), .A2(n1681), .ZN(n1690) );
XNOR2_X1 U1282 ( .A(n1692), .B(KEYINPUT59), .ZN(n1691) );
NAND2_X1 U1283 ( .A1(DATA_IN_3_), .A2(n1682), .ZN(n1689) );
NAND2_X1 U1284 ( .A1(n1693), .A2(n1694), .ZN(U331) );
NAND2_X1 U1285 ( .A1(DATA_IN_2_), .A2(n1682), .ZN(n1694) );
NAND2_X1 U1286 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1681), .ZN(n1693) );
NAND2_X1 U1287 ( .A1(n1695), .A2(n1696), .ZN(U330) );
NAND2_X1 U1288 ( .A1(DATA_IN_1_), .A2(n1682), .ZN(n1696) );
NAND2_X1 U1289 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1681), .ZN(n1695) );
NAND2_X1 U1290 ( .A1(n1697), .A2(n1698), .ZN(U329) );
NAND2_X1 U1291 ( .A1(DATA_IN_0_), .A2(n1699), .ZN(n1698) );
XNOR2_X1 U1292 ( .A(KEYINPUT30), .B(n1682), .ZN(n1699) );
NAND2_X1 U1293 ( .A1(n1676), .A2(n1700), .ZN(n1682) );
NAND2_X1 U1294 ( .A1(n1701), .A2(n1702), .ZN(n1700) );
XNOR2_X1 U1295 ( .A(n1703), .B(KEYINPUT48), .ZN(n1702) );
INV_X1 U1296 ( .A(n1704), .ZN(n1701) );
NAND2_X1 U1297 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1681), .ZN(n1697) );
NAND2_X1 U1298 ( .A1(n1673), .A2(n1705), .ZN(n1681) );
NAND2_X1 U1299 ( .A1(n1704), .A2(n1676), .ZN(n1705) );
NAND3_X1 U1300 ( .A1(n1677), .A2(n1675), .A3(n1706), .ZN(n1704) );
NAND2_X1 U1301 ( .A1(n1707), .A2(n1708), .ZN(n1706) );
NAND3_X1 U1302 ( .A1(n1709), .A2(n1710), .A3(n1711), .ZN(n1708) );
XOR2_X1 U1303 ( .A(KEYINPUT55), .B(n1712), .Z(n1711) );
NOR2_X1 U1304 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1713), .ZN(n1712) );
XNOR2_X1 U1305 ( .A(DATA_IN_6_), .B(KEYINPUT56), .ZN(n1713) );
NAND3_X1 U1306 ( .A1(n1714), .A2(n1715), .A3(n1716), .ZN(n1710) );
NAND2_X1 U1307 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1717), .ZN(n1716) );
NAND3_X1 U1308 ( .A1(n1718), .A2(n1719), .A3(n1720), .ZN(n1715) );
NAND2_X1 U1309 ( .A1(DATA_IN_4_), .A2(n1721), .ZN(n1720) );
NAND3_X1 U1310 ( .A1(n1722), .A2(n1723), .A3(n1724), .ZN(n1719) );
NAND2_X1 U1311 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1725), .ZN(n1724) );
NAND3_X1 U1312 ( .A1(n1726), .A2(n1727), .A3(n1728), .ZN(n1723) );
NAND2_X1 U1313 ( .A1(DATA_IN_3_), .A2(n1692), .ZN(n1728) );
NAND3_X1 U1314 ( .A1(n1729), .A2(n1730), .A3(n1731), .ZN(n1727) );
NAND2_X1 U1315 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1664), .ZN(n1731) );
NAND3_X1 U1316 ( .A1(n1732), .A2(n1733), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1730) );
NAND2_X1 U1317 ( .A1(DATA_IN_1_), .A2(n1734), .ZN(n1732) );
NAND2_X1 U1318 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1735), .ZN(n1729) );
NAND2_X1 U1319 ( .A1(DATA_IN_2_), .A2(n1736), .ZN(n1726) );
NAND2_X1 U1320 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1737), .ZN(n1722) );
NAND2_X1 U1321 ( .A1(DATA_IN_5_), .A2(n1738), .ZN(n1718) );
XNOR2_X1 U1322 ( .A(n1739), .B(KEYINPUT13), .ZN(n1738) );
NAND2_X1 U1323 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1740), .ZN(n1714) );
OR2_X1 U1324 ( .A1(n1741), .A2(DATA_IN_7_), .ZN(n1709) );
NAND2_X1 U1325 ( .A1(DATA_IN_7_), .A2(n1741), .ZN(n1707) );
NAND2_X1 U1326 ( .A1(n1742), .A2(RMAX_REG_7__SCAN_IN), .ZN(n1675) );
XNOR2_X1 U1327 ( .A(DATA_IN_7_), .B(KEYINPUT46), .ZN(n1742) );
NAND3_X1 U1328 ( .A1(n1743), .A2(n1744), .A3(n1745), .ZN(n1677) );
XOR2_X1 U1329 ( .A(n1746), .B(KEYINPUT1), .Z(n1745) );
NAND2_X1 U1330 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1717), .ZN(n1746) );
NAND3_X1 U1331 ( .A1(n1747), .A2(n1748), .A3(n1749), .ZN(n1744) );
XOR2_X1 U1332 ( .A(KEYINPUT54), .B(n1750), .Z(n1749) );
NOR3_X1 U1333 ( .A1(n1751), .A2(n1752), .A3(n1753), .ZN(n1750) );
NOR2_X1 U1334 ( .A1(DATA_IN_5_), .A2(n1754), .ZN(n1753) );
NOR3_X1 U1335 ( .A1(n1755), .A2(n1756), .A3(n1757), .ZN(n1752) );
NOR2_X1 U1336 ( .A1(n1758), .A2(n1759), .ZN(n1757) );
XNOR2_X1 U1337 ( .A(n1760), .B(KEYINPUT3), .ZN(n1759) );
XNOR2_X1 U1338 ( .A(KEYINPUT26), .B(n1737), .ZN(n1758) );
NOR2_X1 U1339 ( .A1(n1725), .A2(n1761), .ZN(n1756) );
XNOR2_X1 U1340 ( .A(n1762), .B(KEYINPUT61), .ZN(n1761) );
NOR3_X1 U1341 ( .A1(n1763), .A2(n1764), .A3(n1765), .ZN(n1755) );
NOR2_X1 U1342 ( .A1(DATA_IN_2_), .A2(n1766), .ZN(n1765) );
NOR2_X1 U1343 ( .A1(n1767), .A2(n1768), .ZN(n1764) );
AND2_X1 U1344 ( .A1(n1766), .A2(DATA_IN_2_), .ZN(n1767) );
NAND2_X1 U1345 ( .A1(n1769), .A2(n1770), .ZN(n1766) );
NAND3_X1 U1346 ( .A1(n1771), .A2(n1772), .A3(DATA_IN_0_), .ZN(n1770) );
INV_X1 U1347 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1772) );
NAND2_X1 U1348 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1735), .ZN(n1771) );
INV_X1 U1349 ( .A(DATA_IN_1_), .ZN(n1735) );
NAND2_X1 U1350 ( .A1(DATA_IN_1_), .A2(n1773), .ZN(n1769) );
NOR2_X1 U1351 ( .A1(DATA_IN_3_), .A2(n1760), .ZN(n1763) );
NOR2_X1 U1352 ( .A1(n1774), .A2(n1762), .ZN(n1751) );
XNOR2_X1 U1353 ( .A(DATA_IN_4_), .B(KEYINPUT0), .ZN(n1774) );
NAND2_X1 U1354 ( .A1(DATA_IN_5_), .A2(n1754), .ZN(n1748) );
OR2_X1 U1355 ( .A1(n1717), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1747) );
NAND2_X1 U1356 ( .A1(DATA_IN_7_), .A2(n1775), .ZN(n1743) );
NAND2_X1 U1357 ( .A1(n1776), .A2(n1777), .ZN(U328) );
NAND2_X1 U1358 ( .A1(n1778), .A2(DATA_IN_7_), .ZN(n1777) );
NAND2_X1 U1359 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1779), .ZN(n1776) );
NAND2_X1 U1360 ( .A1(n1780), .A2(n1781), .ZN(U327) );
NAND2_X1 U1361 ( .A1(n1778), .A2(DATA_IN_6_), .ZN(n1781) );
NAND2_X1 U1362 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1779), .ZN(n1780) );
NAND2_X1 U1363 ( .A1(n1782), .A2(n1783), .ZN(U326) );
NAND2_X1 U1364 ( .A1(n1778), .A2(DATA_IN_5_), .ZN(n1783) );
NAND2_X1 U1365 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1779), .ZN(n1782) );
NAND2_X1 U1366 ( .A1(n1784), .A2(n1785), .ZN(U325) );
NAND2_X1 U1367 ( .A1(n1778), .A2(n1786), .ZN(n1785) );
XNOR2_X1 U1368 ( .A(KEYINPUT27), .B(n1725), .ZN(n1786) );
NAND2_X1 U1369 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1779), .ZN(n1784) );
NAND2_X1 U1370 ( .A1(n1787), .A2(n1788), .ZN(U324) );
NAND2_X1 U1371 ( .A1(n1778), .A2(DATA_IN_3_), .ZN(n1788) );
NAND2_X1 U1372 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1779), .ZN(n1787) );
NAND2_X1 U1373 ( .A1(n1789), .A2(n1790), .ZN(U323) );
NAND2_X1 U1374 ( .A1(n1778), .A2(DATA_IN_2_), .ZN(n1790) );
XOR2_X1 U1375 ( .A(n1791), .B(KEYINPUT35), .Z(n1789) );
NAND2_X1 U1376 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1779), .ZN(n1791) );
NAND2_X1 U1377 ( .A1(n1792), .A2(n1793), .ZN(U322) );
NAND2_X1 U1378 ( .A1(n1778), .A2(DATA_IN_1_), .ZN(n1793) );
NAND2_X1 U1379 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1779), .ZN(n1792) );
NAND2_X1 U1380 ( .A1(n1794), .A2(n1795), .ZN(U321) );
NAND2_X1 U1381 ( .A1(n1778), .A2(DATA_IN_0_), .ZN(n1795) );
AND2_X1 U1382 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1796), .ZN(n1778) );
NAND2_X1 U1383 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1779), .ZN(n1794) );
NAND2_X1 U1384 ( .A1(n1673), .A2(n1796), .ZN(n1779) );
NAND2_X1 U1385 ( .A1(n1676), .A2(n1797), .ZN(n1796) );
INV_X1 U1386 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1676) );
INV_X1 U1387 ( .A(U375), .ZN(n1673) );
NOR2_X1 U1388 ( .A1(STATO_REG_0__SCAN_IN), .A2(STATO_REG_1__SCAN_IN), .ZN(U375) );
NAND2_X1 U1389 ( .A1(n1798), .A2(n1799), .ZN(U320) );
NAND2_X1 U1390 ( .A1(n1648), .A2(DATA_IN_7_), .ZN(n1799) );
NAND2_X1 U1391 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1800), .ZN(n1798) );
NAND2_X1 U1392 ( .A1(n1801), .A2(n1802), .ZN(U319) );
NAND2_X1 U1393 ( .A1(n1648), .A2(DATA_IN_6_), .ZN(n1802) );
NAND2_X1 U1394 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1800), .ZN(n1801) );
NAND2_X1 U1395 ( .A1(n1803), .A2(n1804), .ZN(U318) );
NAND2_X1 U1396 ( .A1(n1648), .A2(DATA_IN_5_), .ZN(n1804) );
NAND2_X1 U1397 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1800), .ZN(n1803) );
NAND2_X1 U1398 ( .A1(n1805), .A2(n1806), .ZN(U317) );
NAND2_X1 U1399 ( .A1(n1648), .A2(DATA_IN_4_), .ZN(n1806) );
NAND2_X1 U1400 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1800), .ZN(n1805) );
NAND2_X1 U1401 ( .A1(n1807), .A2(n1808), .ZN(U316) );
NAND2_X1 U1402 ( .A1(n1809), .A2(n1648), .ZN(n1808) );
XNOR2_X1 U1403 ( .A(DATA_IN_3_), .B(KEYINPUT21), .ZN(n1809) );
NAND2_X1 U1404 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1800), .ZN(n1807) );
NAND2_X1 U1405 ( .A1(n1810), .A2(n1811), .ZN(U315) );
NAND2_X1 U1406 ( .A1(DATA_IN_2_), .A2(n1812), .ZN(n1811) );
XNOR2_X1 U1407 ( .A(KEYINPUT29), .B(n1647), .ZN(n1812) );
NAND2_X1 U1408 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1800), .ZN(n1810) );
NAND2_X1 U1409 ( .A1(n1813), .A2(n1814), .ZN(U314) );
NAND2_X1 U1410 ( .A1(n1648), .A2(DATA_IN_1_), .ZN(n1814) );
NAND2_X1 U1411 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1800), .ZN(n1813) );
NAND2_X1 U1412 ( .A1(n1815), .A2(n1816), .ZN(U313) );
NAND2_X1 U1413 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1800), .ZN(n1816) );
XOR2_X1 U1414 ( .A(KEYINPUT43), .B(n1817), .Z(n1815) );
NOR2_X1 U1415 ( .A1(n1733), .A2(n1647), .ZN(n1817) );
NAND2_X1 U1416 ( .A1(n1818), .A2(n1819), .ZN(U312) );
NAND2_X1 U1417 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1648), .ZN(n1819) );
NAND2_X1 U1418 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1800), .ZN(n1818) );
NAND2_X1 U1419 ( .A1(n1820), .A2(n1821), .ZN(U311) );
NAND2_X1 U1420 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1648), .ZN(n1821) );
NAND2_X1 U1421 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1800), .ZN(n1820) );
NAND2_X1 U1422 ( .A1(n1822), .A2(n1823), .ZN(U310) );
NAND2_X1 U1423 ( .A1(n1824), .A2(n1800), .ZN(n1823) );
XNOR2_X1 U1424 ( .A(REG2_REG_5__SCAN_IN), .B(KEYINPUT15), .ZN(n1824) );
NAND2_X1 U1425 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1648), .ZN(n1822) );
NAND2_X1 U1426 ( .A1(n1825), .A2(n1826), .ZN(U309) );
NAND2_X1 U1427 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1648), .ZN(n1826) );
NAND2_X1 U1428 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1800), .ZN(n1825) );
NAND2_X1 U1429 ( .A1(n1827), .A2(n1828), .ZN(U308) );
NAND2_X1 U1430 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1648), .ZN(n1828) );
XOR2_X1 U1431 ( .A(n1829), .B(KEYINPUT53), .Z(n1827) );
NAND2_X1 U1432 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1800), .ZN(n1829) );
NAND2_X1 U1433 ( .A1(n1830), .A2(n1831), .ZN(U307) );
NAND2_X1 U1434 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1648), .ZN(n1831) );
NAND2_X1 U1435 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1800), .ZN(n1830) );
NAND2_X1 U1436 ( .A1(n1832), .A2(n1833), .ZN(U306) );
NAND2_X1 U1437 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1800), .ZN(n1833) );
XOR2_X1 U1438 ( .A(KEYINPUT31), .B(n1834), .Z(n1832) );
AND2_X1 U1439 ( .A1(n1648), .A2(REG1_REG_1__SCAN_IN), .ZN(n1834) );
NAND2_X1 U1440 ( .A1(n1835), .A2(n1836), .ZN(U305) );
NAND2_X1 U1441 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1800), .ZN(n1836) );
XOR2_X1 U1442 ( .A(n1837), .B(KEYINPUT58), .Z(n1835) );
NAND2_X1 U1443 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1648), .ZN(n1837) );
NAND2_X1 U1444 ( .A1(n1838), .A2(n1839), .ZN(U304) );
NAND2_X1 U1445 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1648), .ZN(n1839) );
NAND2_X1 U1446 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1800), .ZN(n1838) );
NAND2_X1 U1447 ( .A1(n1840), .A2(n1841), .ZN(U303) );
NAND2_X1 U1448 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1648), .ZN(n1841) );
NAND2_X1 U1449 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1800), .ZN(n1840) );
NAND2_X1 U1450 ( .A1(n1842), .A2(n1843), .ZN(U302) );
NAND2_X1 U1451 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1648), .ZN(n1843) );
NAND2_X1 U1452 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1800), .ZN(n1842) );
NAND2_X1 U1453 ( .A1(n1844), .A2(n1845), .ZN(U301) );
NAND2_X1 U1454 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1648), .ZN(n1845) );
NAND2_X1 U1455 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1800), .ZN(n1844) );
NAND2_X1 U1456 ( .A1(n1846), .A2(n1847), .ZN(U300) );
NAND2_X1 U1457 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1648), .ZN(n1847) );
NAND2_X1 U1458 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1800), .ZN(n1846) );
NAND2_X1 U1459 ( .A1(n1848), .A2(n1849), .ZN(U299) );
NAND2_X1 U1460 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1648), .ZN(n1849) );
NAND2_X1 U1461 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1800), .ZN(n1848) );
NAND2_X1 U1462 ( .A1(n1850), .A2(n1851), .ZN(U298) );
NAND2_X1 U1463 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1648), .ZN(n1851) );
NAND2_X1 U1464 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1800), .ZN(n1850) );
NAND2_X1 U1465 ( .A1(n1852), .A2(n1853), .ZN(U297) );
NAND2_X1 U1466 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1648), .ZN(n1853) );
NAND2_X1 U1467 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1800), .ZN(n1852) );
NAND2_X1 U1468 ( .A1(n1854), .A2(n1855), .ZN(U296) );
NAND2_X1 U1469 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1648), .ZN(n1855) );
NAND2_X1 U1470 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1800), .ZN(n1854) );
NAND2_X1 U1471 ( .A1(n1856), .A2(n1857), .ZN(U295) );
NAND2_X1 U1472 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1648), .ZN(n1857) );
NAND2_X1 U1473 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1800), .ZN(n1856) );
NAND2_X1 U1474 ( .A1(n1858), .A2(n1859), .ZN(U294) );
NAND2_X1 U1475 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1648), .ZN(n1859) );
NAND2_X1 U1476 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1800), .ZN(n1858) );
NAND2_X1 U1477 ( .A1(n1860), .A2(n1861), .ZN(U293) );
NAND2_X1 U1478 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1648), .ZN(n1861) );
NAND2_X1 U1479 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1800), .ZN(n1860) );
NAND2_X1 U1480 ( .A1(n1862), .A2(n1863), .ZN(U292) );
NAND2_X1 U1481 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1648), .ZN(n1863) );
NAND2_X1 U1482 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1800), .ZN(n1862) );
NAND2_X1 U1483 ( .A1(n1864), .A2(n1865), .ZN(U291) );
NAND2_X1 U1484 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1648), .ZN(n1865) );
NAND2_X1 U1485 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1800), .ZN(n1864) );
NAND2_X1 U1486 ( .A1(n1866), .A2(n1867), .ZN(U290) );
NAND2_X1 U1487 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1648), .ZN(n1867) );
NAND2_X1 U1488 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1800), .ZN(n1866) );
NAND2_X1 U1489 ( .A1(n1868), .A2(n1869), .ZN(U289) );
NAND2_X1 U1490 ( .A1(n1648), .A2(n1870), .ZN(n1869) );
XOR2_X1 U1491 ( .A(REG3_REG_0__SCAN_IN), .B(KEYINPUT10), .Z(n1870) );
XOR2_X1 U1492 ( .A(n1871), .B(KEYINPUT7), .Z(n1868) );
NAND2_X1 U1493 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1800), .ZN(n1871) );
NAND4_X1 U1494 ( .A1(n1872), .A2(n1873), .A3(n1874), .A4(n1875), .ZN(U288));
NAND2_X1 U1495 ( .A1(n1876), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1874) );
NAND2_X1 U1496 ( .A1(n1877), .A2(REG4_REG_7__SCAN_IN), .ZN(n1873) );
NAND2_X1 U1497 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1800), .ZN(n1872) );
NAND4_X1 U1498 ( .A1(n1878), .A2(n1879), .A3(n1880), .A4(n1881), .ZN(U287));
NOR3_X1 U1499 ( .A1(n1882), .A2(n1883), .A3(n1884), .ZN(n1881) );
NOR4_X1 U1500 ( .A1(n1885), .A2(n1886), .A3(n1887), .A4(n1888), .ZN(n1884));
INV_X1 U1501 ( .A(n1889), .ZN(n1888) );
INV_X1 U1502 ( .A(n1875), .ZN(n1883) );
NAND2_X1 U1503 ( .A1(n1885), .A2(n1890), .ZN(n1875) );
NOR4_X1 U1504 ( .A1(n1891), .A2(n1892), .A3(n1893), .A4(n1894), .ZN(n1882));
NAND2_X1 U1505 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1800), .ZN(n1880) );
NAND2_X1 U1506 ( .A1(n1876), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1879) );
NAND2_X1 U1507 ( .A1(n1877), .A2(REG4_REG_6__SCAN_IN), .ZN(n1878) );
NAND4_X1 U1508 ( .A1(n1895), .A2(n1896), .A3(n1897), .A4(n1898), .ZN(U286));
AND4_X1 U1509 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .ZN(n1898));
NAND2_X1 U1510 ( .A1(n1890), .A2(n1903), .ZN(n1902) );
INV_X1 U1511 ( .A(n1886), .ZN(n1903) );
NAND3_X1 U1512 ( .A1(n1889), .A2(n1904), .A3(n1886), .ZN(n1901) );
NOR2_X1 U1513 ( .A1(n1905), .A2(n1885), .ZN(n1886) );
NOR2_X1 U1514 ( .A1(n1906), .A2(n1907), .ZN(n1885) );
AND2_X1 U1515 ( .A1(n1907), .A2(n1906), .ZN(n1905) );
NAND2_X1 U1516 ( .A1(n1877), .A2(REG4_REG_5__SCAN_IN), .ZN(n1900) );
NAND2_X1 U1517 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1800), .ZN(n1899) );
NAND2_X1 U1518 ( .A1(n1876), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1897) );
NAND2_X1 U1519 ( .A1(n1908), .A2(n1909), .ZN(n1896) );
XOR2_X1 U1520 ( .A(n1893), .B(n1892), .Z(n1909) );
XNOR2_X1 U1521 ( .A(n1891), .B(n1907), .ZN(n1892) );
NAND2_X1 U1522 ( .A1(n1910), .A2(n1907), .ZN(n1895) );
AND2_X1 U1523 ( .A1(n1911), .A2(n1912), .ZN(n1907) );
NAND4_X1 U1524 ( .A1(n1913), .A2(n1914), .A3(n1915), .A4(n1916), .ZN(n1912));
NAND2_X1 U1525 ( .A1(n1917), .A2(n1918), .ZN(n1916) );
XNOR2_X1 U1526 ( .A(n1919), .B(DATA_IN_6_), .ZN(n1917) );
NAND2_X1 U1527 ( .A1(n1920), .A2(RESTART), .ZN(n1915) );
XNOR2_X1 U1528 ( .A(n1921), .B(RMAX_REG_6__SCAN_IN), .ZN(n1920) );
NAND2_X1 U1529 ( .A1(n1922), .A2(n1923), .ZN(n1914) );
NAND4_X1 U1530 ( .A1(n1923), .A2(n1924), .A3(n1925), .A4(n1926), .ZN(n1911));
NAND2_X1 U1531 ( .A1(n1927), .A2(n1918), .ZN(n1926) );
XNOR2_X1 U1532 ( .A(REG4_REG_6__SCAN_IN), .B(DATA_IN_6_), .ZN(n1927) );
NAND2_X1 U1533 ( .A1(n1928), .A2(RESTART), .ZN(n1925) );
XNOR2_X1 U1534 ( .A(RMAX_REG_6__SCAN_IN), .B(RMIN_REG_6__SCAN_IN), .ZN(n1928) );
NAND2_X1 U1535 ( .A1(n1913), .A2(n1929), .ZN(n1924) );
NAND2_X1 U1536 ( .A1(n1930), .A2(n1931), .ZN(n1913) );
INV_X1 U1537 ( .A(n1932), .ZN(n1930) );
NAND2_X1 U1538 ( .A1(n1933), .A2(n1932), .ZN(n1923) );
NAND4_X1 U1539 ( .A1(n1934), .A2(n1935), .A3(n1936), .A4(n1937), .ZN(U285));
NOR3_X1 U1540 ( .A1(n1938), .A2(n1939), .A3(n1940), .ZN(n1937) );
NOR2_X1 U1541 ( .A1(n1941), .A2(n1942), .ZN(n1940) );
NOR2_X1 U1542 ( .A1(n1943), .A2(n1944), .ZN(n1939) );
XNOR2_X1 U1543 ( .A(n1877), .B(KEYINPUT23), .ZN(n1943) );
AND2_X1 U1544 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1876), .ZN(n1938) );
NAND2_X1 U1545 ( .A1(n1945), .A2(n1800), .ZN(n1936) );
XNOR2_X1 U1546 ( .A(KEYINPUT24), .B(DATA_OUT_REG_4__SCAN_IN), .ZN(n1945) );
NAND3_X1 U1547 ( .A1(n1946), .A2(n1893), .A3(n1908), .ZN(n1935) );
NAND3_X1 U1548 ( .A1(n1947), .A2(n1948), .A3(n1949), .ZN(n1893) );
NAND2_X1 U1549 ( .A1(n1950), .A2(n1951), .ZN(n1948) );
INV_X1 U1550 ( .A(n1891), .ZN(n1951) );
NOR3_X1 U1551 ( .A1(n1952), .A2(n1953), .A3(n1954), .ZN(n1891) );
XNOR2_X1 U1552 ( .A(n1955), .B(n1941), .ZN(n1954) );
XNOR2_X1 U1553 ( .A(KEYINPUT62), .B(KEYINPUT11), .ZN(n1955) );
NAND2_X1 U1554 ( .A1(n1952), .A2(n1956), .ZN(n1950) );
NAND2_X1 U1555 ( .A1(n1941), .A2(n1957), .ZN(n1946) );
NAND2_X1 U1556 ( .A1(n1949), .A2(n1947), .ZN(n1957) );
INV_X1 U1557 ( .A(n1956), .ZN(n1941) );
NAND2_X1 U1558 ( .A1(n1890), .A2(n1958), .ZN(n1934) );
NAND2_X1 U1559 ( .A1(n1959), .A2(n1960), .ZN(n1958) );
NOR2_X1 U1560 ( .A1(n1887), .A2(n1889), .ZN(n1890) );
NOR2_X1 U1561 ( .A1(n1960), .A2(n1959), .ZN(n1889) );
AND2_X1 U1562 ( .A1(n1906), .A2(n1961), .ZN(n1959) );
NAND2_X1 U1563 ( .A1(n1956), .A2(n1962), .ZN(n1961) );
OR2_X1 U1564 ( .A1(n1962), .A2(n1956), .ZN(n1906) );
NAND2_X1 U1565 ( .A1(n1963), .A2(n1964), .ZN(n1956) );
NAND2_X1 U1566 ( .A1(n1965), .A2(n1922), .ZN(n1964) );
XOR2_X1 U1567 ( .A(KEYINPUT18), .B(n1966), .Z(n1963) );
NOR2_X1 U1568 ( .A1(n1922), .A2(n1965), .ZN(n1966) );
XNOR2_X1 U1569 ( .A(n1933), .B(n1932), .ZN(n1965) );
NAND2_X1 U1570 ( .A1(n1967), .A2(n1968), .ZN(n1932) );
NAND2_X1 U1571 ( .A1(RESTART), .A2(n1754), .ZN(n1968) );
NAND2_X1 U1572 ( .A1(n1740), .A2(n1918), .ZN(n1967) );
INV_X1 U1573 ( .A(n1931), .ZN(n1933) );
NAND3_X1 U1574 ( .A1(n1969), .A2(n1970), .A3(n1971), .ZN(n1931) );
OR2_X1 U1575 ( .A1(KEYINPUT36), .A2(RMIN_REG_5__SCAN_IN), .ZN(n1971) );
NAND3_X1 U1576 ( .A1(KEYINPUT36), .A2(RMIN_REG_5__SCAN_IN), .A3(RESTART),
.ZN(n1970) );
NAND2_X1 U1577 ( .A1(n1972), .A2(n1918), .ZN(n1969) );
NAND2_X1 U1578 ( .A1(KEYINPUT36), .A2(n1973), .ZN(n1972) );
INV_X1 U1579 ( .A(n1929), .ZN(n1922) );
NAND2_X1 U1580 ( .A1(n1974), .A2(n1975), .ZN(n1929) );
NAND2_X1 U1581 ( .A1(n1976), .A2(n1977), .ZN(n1975) );
NAND2_X1 U1582 ( .A1(n1978), .A2(n1979), .ZN(n1977) );
XNOR2_X1 U1583 ( .A(KEYINPUT51), .B(n1980), .ZN(n1978) );
NAND2_X1 U1584 ( .A1(n1980), .A2(n1981), .ZN(n1974) );
NAND4_X1 U1585 ( .A1(n1982), .A2(n1983), .A3(n1984), .A4(n1985), .ZN(U284));
NAND3_X1 U1586 ( .A1(n1986), .A2(n1987), .A3(n1904), .ZN(n1985) );
NAND3_X1 U1587 ( .A1(n1988), .A2(n1962), .A3(n1989), .ZN(n1987) );
XNOR2_X1 U1588 ( .A(KEYINPUT41), .B(n1960), .ZN(n1986) );
NAND2_X1 U1589 ( .A1(n1990), .A2(n1991), .ZN(n1960) );
NAND2_X1 U1590 ( .A1(n1989), .A2(n1962), .ZN(n1991) );
NAND2_X1 U1591 ( .A1(n1992), .A2(n1993), .ZN(n1962) );
XOR2_X1 U1592 ( .A(n1952), .B(KEYINPUT33), .Z(n1993) );
XNOR2_X1 U1593 ( .A(n1994), .B(KEYINPUT2), .ZN(n1989) );
NAND2_X1 U1594 ( .A1(n1995), .A2(n1952), .ZN(n1994) );
XNOR2_X1 U1595 ( .A(n1992), .B(KEYINPUT5), .ZN(n1995) );
NAND2_X1 U1596 ( .A1(n1908), .A2(n1996), .ZN(n1984) );
XOR2_X1 U1597 ( .A(n1949), .B(n1947), .Z(n1996) );
XNOR2_X1 U1598 ( .A(n1952), .B(n1953), .ZN(n1947) );
NAND2_X1 U1599 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1800), .ZN(n1983) );
XOR2_X1 U1600 ( .A(n1997), .B(KEYINPUT37), .Z(n1982) );
NAND3_X1 U1601 ( .A1(n1998), .A2(n1999), .A3(n2000), .ZN(n1997) );
NAND2_X1 U1602 ( .A1(n1877), .A2(REG4_REG_3__SCAN_IN), .ZN(n2000) );
NAND2_X1 U1603 ( .A1(n1910), .A2(n1952), .ZN(n1999) );
XNOR2_X1 U1604 ( .A(n2001), .B(n1980), .ZN(n1952) );
NAND2_X1 U1605 ( .A1(n2002), .A2(n2003), .ZN(n1980) );
NAND2_X1 U1606 ( .A1(RESTART), .A2(n1762), .ZN(n2003) );
NAND2_X1 U1607 ( .A1(n1725), .A2(n1918), .ZN(n2002) );
XNOR2_X1 U1608 ( .A(n1979), .B(n1976), .ZN(n2001) );
AND3_X1 U1609 ( .A1(n2004), .A2(n2005), .A3(n2006), .ZN(n1976) );
NAND2_X1 U1610 ( .A1(KEYINPUT42), .A2(n1721), .ZN(n2006) );
NAND3_X1 U1611 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n2007), .A3(RESTART), .ZN(n2005) );
NAND2_X1 U1612 ( .A1(n2008), .A2(n1918), .ZN(n2004) );
NAND2_X1 U1613 ( .A1(n2007), .A2(n1944), .ZN(n2008) );
INV_X1 U1614 ( .A(KEYINPUT42), .ZN(n2007) );
INV_X1 U1615 ( .A(n1981), .ZN(n1979) );
NAND2_X1 U1616 ( .A1(n2009), .A2(n2010), .ZN(n1981) );
NAND2_X1 U1617 ( .A1(n2011), .A2(n2012), .ZN(n2010) );
OR2_X1 U1618 ( .A1(n2013), .A2(n2014), .ZN(n2011) );
NAND2_X1 U1619 ( .A1(n2014), .A2(n2013), .ZN(n2009) );
NAND2_X1 U1620 ( .A1(n1876), .A2(RLAST_REG_3__SCAN_IN), .ZN(n1998) );
NAND4_X1 U1621 ( .A1(n2015), .A2(n2016), .A3(n2017), .A4(n2018), .ZN(U283));
NOR3_X1 U1622 ( .A1(n2019), .A2(n2020), .A3(n2021), .ZN(n2018) );
NOR3_X1 U1623 ( .A1(n1894), .A2(n1949), .A3(n2022), .ZN(n2021) );
NOR2_X1 U1624 ( .A1(n2023), .A2(n2024), .ZN(n2022) );
NOR2_X1 U1625 ( .A1(n2025), .A2(n2026), .ZN(n2023) );
AND3_X1 U1626 ( .A1(n2027), .A2(n2028), .A3(n2029), .ZN(n1949) );
NAND2_X1 U1627 ( .A1(n1953), .A2(n2030), .ZN(n2029) );
NAND2_X1 U1628 ( .A1(n2024), .A2(n2031), .ZN(n2030) );
NAND2_X1 U1629 ( .A1(n2032), .A2(n2033), .ZN(n1953) );
XNOR2_X1 U1630 ( .A(n2024), .B(KEYINPUT16), .ZN(n2032) );
NOR3_X1 U1631 ( .A1(n1887), .A2(n1990), .A3(n2034), .ZN(n2020) );
NOR2_X1 U1632 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
AND2_X1 U1633 ( .A1(n2037), .A2(n2038), .ZN(n2035) );
INV_X1 U1634 ( .A(n1988), .ZN(n1990) );
NAND3_X1 U1635 ( .A1(n2038), .A2(n2037), .A3(n2036), .ZN(n1988) );
NAND2_X1 U1636 ( .A1(n2039), .A2(n2040), .ZN(n2036) );
NAND2_X1 U1637 ( .A1(n2024), .A2(n2041), .ZN(n2040) );
NAND2_X1 U1638 ( .A1(n2033), .A2(n2042), .ZN(n2041) );
NAND2_X1 U1639 ( .A1(n1992), .A2(n2042), .ZN(n2039) );
INV_X1 U1640 ( .A(KEYINPUT47), .ZN(n2042) );
NOR2_X1 U1641 ( .A1(n2031), .A2(n2024), .ZN(n1992) );
NOR2_X1 U1642 ( .A1(n2043), .A2(n2044), .ZN(n2019) );
XNOR2_X1 U1643 ( .A(n2045), .B(KEYINPUT19), .ZN(n2044) );
NAND2_X1 U1644 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1800), .ZN(n2017) );
NAND2_X1 U1645 ( .A1(n1910), .A2(n2024), .ZN(n2016) );
XNOR2_X1 U1646 ( .A(n2012), .B(n2046), .ZN(n2024) );
NOR2_X1 U1647 ( .A1(KEYINPUT25), .A2(n2047), .ZN(n2046) );
XNOR2_X1 U1648 ( .A(n2014), .B(n2013), .ZN(n2047) );
NAND2_X1 U1649 ( .A1(n2048), .A2(n2049), .ZN(n2013) );
NAND2_X1 U1650 ( .A1(RESTART), .A2(n1760), .ZN(n2049) );
NAND2_X1 U1651 ( .A1(n1737), .A2(n1918), .ZN(n2048) );
INV_X1 U1652 ( .A(DATA_IN_3_), .ZN(n1737) );
NAND2_X1 U1653 ( .A1(n2050), .A2(n2051), .ZN(n2014) );
NAND2_X1 U1654 ( .A1(RESTART), .A2(n1692), .ZN(n2051) );
NAND2_X1 U1655 ( .A1(n2052), .A2(n1918), .ZN(n2050) );
NAND2_X1 U1656 ( .A1(n2053), .A2(n2054), .ZN(n2012) );
NAND2_X1 U1657 ( .A1(n2055), .A2(n2056), .ZN(n2054) );
OR2_X1 U1658 ( .A1(n2057), .A2(n2058), .ZN(n2056) );
NAND2_X1 U1659 ( .A1(n2058), .A2(n2057), .ZN(n2053) );
INV_X1 U1660 ( .A(n1942), .ZN(n1910) );
NAND2_X1 U1661 ( .A1(n1876), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2015) );
NAND4_X1 U1662 ( .A1(n2059), .A2(n2060), .A3(n2061), .A4(n2062), .ZN(U282));
NOR3_X1 U1663 ( .A1(n2063), .A2(n2064), .A3(n2065), .ZN(n2062) );
NOR2_X1 U1664 ( .A1(n2066), .A2(n1887), .ZN(n2065) );
XNOR2_X1 U1665 ( .A(n2038), .B(n2037), .ZN(n2066) );
NAND2_X1 U1666 ( .A1(n2031), .A2(n2067), .ZN(n2038) );
NAND2_X1 U1667 ( .A1(n2068), .A2(n2069), .ZN(n2067) );
NOR3_X1 U1668 ( .A1(n1894), .A2(n2070), .A3(n2071), .ZN(n2064) );
NOR2_X1 U1669 ( .A1(n2028), .A2(n2072), .ZN(n2071) );
NOR2_X1 U1670 ( .A1(n2073), .A2(n2074), .ZN(n2072) );
AND3_X1 U1671 ( .A1(KEYINPUT39), .A2(n2026), .A3(KEYINPUT20), .ZN(n2074) );
NOR2_X1 U1672 ( .A1(KEYINPUT39), .A2(n2026), .ZN(n2073) );
NOR2_X1 U1673 ( .A1(n2025), .A2(n2075), .ZN(n2070) );
AND2_X1 U1674 ( .A1(n2026), .A2(KEYINPUT20), .ZN(n2075) );
INV_X1 U1675 ( .A(n2027), .ZN(n2026) );
NAND2_X1 U1676 ( .A1(n2076), .A2(n2031), .ZN(n2027) );
INV_X1 U1677 ( .A(n2033), .ZN(n2031) );
NOR2_X1 U1678 ( .A1(n2069), .A2(n2068), .ZN(n2033) );
INV_X1 U1679 ( .A(n2077), .ZN(n2068) );
XOR2_X1 U1680 ( .A(KEYINPUT28), .B(n2078), .Z(n2076) );
NOR2_X1 U1681 ( .A1(n2079), .A2(n2077), .ZN(n2078) );
XOR2_X1 U1682 ( .A(n2069), .B(KEYINPUT14), .Z(n2079) );
INV_X1 U1683 ( .A(n1908), .ZN(n1894) );
NOR2_X1 U1684 ( .A1(n2077), .A2(n1942), .ZN(n2063) );
XNOR2_X1 U1685 ( .A(n2055), .B(n2080), .ZN(n2077) );
XNOR2_X1 U1686 ( .A(n2081), .B(n2058), .ZN(n2080) );
NAND2_X1 U1687 ( .A1(n2082), .A2(n2083), .ZN(n2058) );
NAND2_X1 U1688 ( .A1(RESTART), .A2(n1736), .ZN(n2083) );
NAND2_X1 U1689 ( .A1(n2045), .A2(n1918), .ZN(n2082) );
NOR2_X1 U1690 ( .A1(KEYINPUT60), .A2(n2084), .ZN(n2081) );
INV_X1 U1691 ( .A(n2057), .ZN(n2084) );
NAND2_X1 U1692 ( .A1(n2085), .A2(n2086), .ZN(n2057) );
NAND2_X1 U1693 ( .A1(n2087), .A2(n2088), .ZN(n2086) );
XNOR2_X1 U1694 ( .A(n2089), .B(KEYINPUT32), .ZN(n2087) );
OR2_X1 U1695 ( .A1(n2090), .A2(n2091), .ZN(n2085) );
NAND2_X1 U1696 ( .A1(n2092), .A2(n2093), .ZN(n2055) );
NAND2_X1 U1697 ( .A1(RESTART), .A2(n1768), .ZN(n2093) );
NAND2_X1 U1698 ( .A1(n1664), .A2(n1918), .ZN(n2092) );
NAND2_X1 U1699 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1800), .ZN(n2061) );
NAND2_X1 U1700 ( .A1(n1876), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2060) );
NAND2_X1 U1701 ( .A1(n1877), .A2(REG4_REG_1__SCAN_IN), .ZN(n2059) );
NAND4_X1 U1702 ( .A1(n2094), .A2(n2095), .A3(n2096), .A4(n2097), .ZN(U281));
NOR3_X1 U1703 ( .A1(n2098), .A2(n2099), .A3(n2100), .ZN(n2097) );
AND2_X1 U1704 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1876), .ZN(n2100) );
NOR2_X1 U1705 ( .A1(n2101), .A2(ENABLE), .ZN(n1876) );
NOR2_X1 U1706 ( .A1(n1942), .A2(n2102), .ZN(n2099) );
XOR2_X1 U1707 ( .A(KEYINPUT45), .B(n2103), .Z(n2102) );
NAND4_X1 U1708 ( .A1(n2104), .A2(STATO_REG_1__SCAN_IN), .A3(n2105), .A4(U280), .ZN(n1942) );
NAND2_X1 U1709 ( .A1(n2106), .A2(n1918), .ZN(n2105) );
NAND3_X1 U1710 ( .A1(n2107), .A2(n2108), .A3(ENABLE), .ZN(n2106) );
XOR2_X1 U1711 ( .A(n2109), .B(KEYINPUT12), .Z(n2104) );
NOR2_X1 U1712 ( .A1(n1887), .A2(n2037), .ZN(n2098) );
NAND2_X1 U1713 ( .A1(n2069), .A2(n2110), .ZN(n2037) );
OR2_X1 U1714 ( .A1(n2111), .A2(n2103), .ZN(n2110) );
INV_X1 U1715 ( .A(n1904), .ZN(n1887) );
NOR3_X1 U1716 ( .A1(n1703), .A2(n1800), .A3(n2109), .ZN(n1904) );
NAND3_X1 U1717 ( .A1(n2112), .A2(n2113), .A3(RESTART), .ZN(n2109) );
NAND2_X1 U1718 ( .A1(n2114), .A2(n1741), .ZN(n2113) );
INV_X1 U1719 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1741) );
OR2_X1 U1720 ( .A1(n2115), .A2(n1775), .ZN(n2114) );
NAND2_X1 U1721 ( .A1(n2115), .A2(n1775), .ZN(n2112) );
INV_X1 U1722 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1775) );
NAND2_X1 U1723 ( .A1(n2116), .A2(n2117), .ZN(n2115) );
NAND2_X1 U1724 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n2118), .ZN(n2117) );
NAND2_X1 U1725 ( .A1(n2119), .A2(n1921), .ZN(n2118) );
INV_X1 U1726 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1921) );
XOR2_X1 U1727 ( .A(KEYINPUT63), .B(n2120), .Z(n2119) );
NAND2_X1 U1728 ( .A1(n2120), .A2(RMIN_REG_6__SCAN_IN), .ZN(n2116) );
AND2_X1 U1729 ( .A1(n2121), .A2(n2122), .ZN(n2120) );
NAND3_X1 U1730 ( .A1(n2123), .A2(n2124), .A3(n2125), .ZN(n2122) );
NAND2_X1 U1731 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2125) );
NAND3_X1 U1732 ( .A1(n2126), .A2(n2127), .A3(n2128), .ZN(n2124) );
NAND2_X1 U1733 ( .A1(n1762), .A2(n1721), .ZN(n2128) );
INV_X1 U1734 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1721) );
INV_X1 U1735 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1762) );
NAND3_X1 U1736 ( .A1(n2129), .A2(n2130), .A3(n2131), .ZN(n2127) );
NAND2_X1 U1737 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2131) );
NAND3_X1 U1738 ( .A1(n2132), .A2(n2133), .A3(n2134), .ZN(n2130) );
NAND2_X1 U1739 ( .A1(n1768), .A2(n1736), .ZN(n2134) );
INV_X1 U1740 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1736) );
INV_X1 U1741 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1768) );
NAND2_X1 U1742 ( .A1(n2135), .A2(n1734), .ZN(n2133) );
INV_X1 U1743 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1734) );
OR2_X1 U1744 ( .A1(n2136), .A2(n1773), .ZN(n2135) );
NAND2_X1 U1745 ( .A1(n2136), .A2(n1773), .ZN(n2132) );
NAND2_X1 U1746 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2129) );
NAND2_X1 U1747 ( .A1(n1760), .A2(n1692), .ZN(n2126) );
INV_X1 U1748 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1692) );
INV_X1 U1749 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1760) );
NAND2_X1 U1750 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n2137), .ZN(n2123) );
XNOR2_X1 U1751 ( .A(n1739), .B(KEYINPUT52), .ZN(n2137) );
NAND2_X1 U1752 ( .A1(n1739), .A2(n1754), .ZN(n2121) );
INV_X1 U1753 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1754) );
INV_X1 U1754 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1739) );
XOR2_X1 U1755 ( .A(KEYINPUT4), .B(n2138), .Z(n2096) );
NOR2_X1 U1756 ( .A1(n2139), .A2(n2043), .ZN(n2138) );
INV_X1 U1757 ( .A(n1877), .ZN(n2043) );
NOR3_X1 U1758 ( .A1(n2108), .A2(n2101), .A3(n1797), .ZN(n1877) );
INV_X1 U1759 ( .A(AVERAGE), .ZN(n2108) );
NAND2_X1 U1760 ( .A1(n2025), .A2(n1908), .ZN(n2095) );
NOR4_X1 U1761 ( .A1(n2107), .A2(n1797), .A3(n2101), .A4(AVERAGE), .ZN(n1908));
NAND3_X1 U1762 ( .A1(U280), .A2(n1918), .A3(STATO_REG_1__SCAN_IN), .ZN(n2101) );
INV_X1 U1763 ( .A(ENABLE), .ZN(n1797) );
NAND2_X1 U1764 ( .A1(n2140), .A2(n2141), .ZN(n2107) );
NAND2_X1 U1765 ( .A1(n2142), .A2(n2143), .ZN(n2141) );
NAND2_X1 U1766 ( .A1(REG4_REG_7__SCAN_IN), .A2(DATA_IN_7_), .ZN(n2143) );
NAND2_X1 U1767 ( .A1(n2144), .A2(n2145), .ZN(n2142) );
NAND2_X1 U1768 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2145) );
NAND3_X1 U1769 ( .A1(n2146), .A2(n2147), .A3(n2148), .ZN(n2144) );
NAND2_X1 U1770 ( .A1(n1717), .A2(n1919), .ZN(n2148) );
INV_X1 U1771 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1919) );
INV_X1 U1772 ( .A(DATA_IN_6_), .ZN(n1717) );
NAND3_X1 U1773 ( .A1(n2149), .A2(n2150), .A3(n2151), .ZN(n2147) );
NAND2_X1 U1774 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2151) );
NAND3_X1 U1775 ( .A1(n2152), .A2(n2153), .A3(n2154), .ZN(n2150) );
NAND2_X1 U1776 ( .A1(n2155), .A2(n2052), .ZN(n2154) );
INV_X1 U1777 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2052) );
XNOR2_X1 U1778 ( .A(DATA_IN_3_), .B(KEYINPUT49), .ZN(n2155) );
NAND3_X1 U1779 ( .A1(n2156), .A2(n2157), .A3(n2158), .ZN(n2153) );
NAND2_X1 U1780 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2158) );
NAND3_X1 U1781 ( .A1(n2159), .A2(n2160), .A3(n2161), .ZN(n2157) );
OR2_X1 U1782 ( .A1(DATA_IN_1_), .A2(REG4_REG_1__SCAN_IN), .ZN(n2161) );
NAND2_X1 U1783 ( .A1(n2162), .A2(n2163), .ZN(n2160) );
NAND2_X1 U1784 ( .A1(n2164), .A2(REG4_REG_1__SCAN_IN), .ZN(n2163) );
XNOR2_X1 U1785 ( .A(DATA_IN_1_), .B(KEYINPUT38), .ZN(n2164) );
NAND2_X1 U1786 ( .A1(n2165), .A2(n1664), .ZN(n2159) );
INV_X1 U1787 ( .A(DATA_IN_2_), .ZN(n1664) );
XNOR2_X1 U1788 ( .A(REG4_REG_2__SCAN_IN), .B(KEYINPUT9), .ZN(n2165) );
NAND2_X1 U1789 ( .A1(DATA_IN_2_), .A2(n2166), .ZN(n2156) );
XNOR2_X1 U1790 ( .A(n2045), .B(KEYINPUT57), .ZN(n2166) );
INV_X1 U1791 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2045) );
NAND2_X1 U1792 ( .A1(n2167), .A2(n1725), .ZN(n2152) );
INV_X1 U1793 ( .A(DATA_IN_4_), .ZN(n1725) );
XNOR2_X1 U1794 ( .A(n1944), .B(KEYINPUT40), .ZN(n2167) );
INV_X1 U1795 ( .A(REG4_REG_4__SCAN_IN), .ZN(n1944) );
NAND2_X1 U1796 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2149) );
NAND2_X1 U1797 ( .A1(n1740), .A2(n1973), .ZN(n2146) );
INV_X1 U1798 ( .A(REG4_REG_5__SCAN_IN), .ZN(n1973) );
INV_X1 U1799 ( .A(DATA_IN_5_), .ZN(n1740) );
OR2_X1 U1800 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2140) );
INV_X1 U1801 ( .A(n2028), .ZN(n2025) );
NAND3_X1 U1802 ( .A1(n2168), .A2(n2169), .A3(n2069), .ZN(n2028) );
NAND2_X1 U1803 ( .A1(n2103), .A2(n2111), .ZN(n2069) );
OR3_X1 U1804 ( .A1(n2111), .A2(n2103), .A3(KEYINPUT22), .ZN(n2169) );
NAND3_X1 U1805 ( .A1(n2170), .A2(n2171), .A3(n2172), .ZN(n2111) );
NAND3_X1 U1806 ( .A1(n1733), .A2(n2139), .A3(n1918), .ZN(n2171) );
INV_X1 U1807 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2139) );
INV_X1 U1808 ( .A(DATA_IN_0_), .ZN(n1733) );
OR3_X1 U1809 ( .A1(RMAX_REG_0__SCAN_IN), .A2(RMIN_REG_0__SCAN_IN), .A3(n1918), .ZN(n2170) );
NAND2_X1 U1810 ( .A1(KEYINPUT22), .A2(n2103), .ZN(n2168) );
AND3_X1 U1811 ( .A1(n2173), .A2(n2174), .A3(n2175), .ZN(n2103) );
NAND2_X1 U1812 ( .A1(n2091), .A2(n2090), .ZN(n2175) );
NOR2_X1 U1813 ( .A1(n2088), .A2(n2172), .ZN(n2091) );
OR3_X1 U1814 ( .A1(n2089), .A2(n2090), .A3(n2088), .ZN(n2174) );
NAND2_X1 U1815 ( .A1(n2176), .A2(n2088), .ZN(n2173) );
NAND2_X1 U1816 ( .A1(n2177), .A2(n2178), .ZN(n2088) );
NAND2_X1 U1817 ( .A1(RESTART), .A2(n1773), .ZN(n2178) );
INV_X1 U1818 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1773) );
NAND2_X1 U1819 ( .A1(n2179), .A2(n1918), .ZN(n2177) );
XNOR2_X1 U1820 ( .A(DATA_IN_1_), .B(KEYINPUT17), .ZN(n2179) );
XOR2_X1 U1821 ( .A(n2090), .B(n2180), .Z(n2176) );
XNOR2_X1 U1822 ( .A(n2089), .B(KEYINPUT34), .ZN(n2180) );
INV_X1 U1823 ( .A(n2172), .ZN(n2089) );
NAND2_X1 U1824 ( .A1(n2181), .A2(n2182), .ZN(n2172) );
NAND2_X1 U1825 ( .A1(RESTART), .A2(n2136), .ZN(n2182) );
NAND2_X1 U1826 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2136) );
NAND2_X1 U1827 ( .A1(n2162), .A2(n1918), .ZN(n2181) );
NAND2_X1 U1828 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2162) );
NAND2_X1 U1829 ( .A1(n2183), .A2(n2184), .ZN(n2090) );
NAND2_X1 U1830 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1918), .ZN(n2184) );
INV_X1 U1831 ( .A(RESTART), .ZN(n1918) );
NAND2_X1 U1832 ( .A1(RESTART), .A2(RMIN_REG_1__SCAN_IN), .ZN(n2183) );
NAND2_X1 U1833 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1800), .ZN(n2094) );
NAND2_X1 U1834 ( .A1(n1647), .A2(n2185), .ZN(U280) );
NAND2_X1 U1835 ( .A1(STATO_REG_0__SCAN_IN), .A2(n1703), .ZN(n2185) );
INV_X1 U1836 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1703) );
endmodule


