//Key = 1000000001011001000011010011101100000010111001110010000000100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;

XOR2_X1 U773 ( .A(G107), .B(n1066), .Z(G9) );
NOR2_X1 U774 ( .A1(n1067), .A2(n1068), .ZN(G75) );
NOR4_X1 U775 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1068) );
INV_X1 U776 ( .A(n1073), .ZN(n1071) );
NOR3_X1 U777 ( .A1(n1074), .A2(KEYINPUT44), .A3(n1075), .ZN(n1070) );
INV_X1 U778 ( .A(n1076), .ZN(n1075) );
NOR2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
NOR3_X1 U780 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NOR2_X1 U781 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR2_X1 U782 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U784 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1082) );
NOR2_X1 U786 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR3_X1 U787 ( .A1(n1091), .A2(n1094), .A3(n1085), .ZN(n1077) );
NOR2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U789 ( .A1(n1097), .A2(n1081), .ZN(n1096) );
NOR2_X1 U790 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U791 ( .A1(n1100), .A2(n1079), .ZN(n1095) );
NOR2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR3_X1 U794 ( .A1(n1072), .A2(G952), .A3(n1069), .ZN(n1067) );
AND4_X1 U795 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1069) );
NOR4_X1 U796 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
INV_X1 U797 ( .A(n1089), .ZN(n1110) );
NOR2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1107) );
XNOR2_X1 U799 ( .A(KEYINPUT18), .B(n1115), .ZN(n1114) );
XNOR2_X1 U800 ( .A(G469), .B(n1116), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1117), .B(n1118), .Z(n1106) );
XNOR2_X1 U802 ( .A(n1119), .B(n1120), .ZN(n1118) );
NOR2_X1 U803 ( .A1(KEYINPUT4), .A2(n1121), .ZN(n1119) );
XOR2_X1 U804 ( .A(KEYINPUT37), .B(n1122), .Z(n1121) );
XNOR2_X1 U805 ( .A(KEYINPUT30), .B(KEYINPUT2), .ZN(n1117) );
XNOR2_X1 U806 ( .A(n1123), .B(n1124), .ZN(n1105) );
NOR2_X1 U807 ( .A1(KEYINPUT7), .A2(n1125), .ZN(n1124) );
XOR2_X1 U808 ( .A(n1126), .B(n1127), .Z(G72) );
XOR2_X1 U809 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U810 ( .A1(G953), .A2(n1130), .ZN(n1129) );
XNOR2_X1 U811 ( .A(KEYINPUT43), .B(n1131), .ZN(n1130) );
NAND2_X1 U812 ( .A1(n1132), .A2(n1133), .ZN(n1128) );
INV_X1 U813 ( .A(n1134), .ZN(n1133) );
XOR2_X1 U814 ( .A(n1135), .B(n1136), .Z(n1132) );
XNOR2_X1 U815 ( .A(n1137), .B(n1138), .ZN(n1136) );
XNOR2_X1 U816 ( .A(G125), .B(G140), .ZN(n1135) );
NAND2_X1 U817 ( .A1(G953), .A2(n1139), .ZN(n1126) );
NAND2_X1 U818 ( .A1(G900), .A2(G227), .ZN(n1139) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(G69) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U822 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
NAND3_X1 U823 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1142) );
XOR2_X1 U824 ( .A(n1151), .B(KEYINPUT5), .Z(n1150) );
NAND2_X1 U825 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
OR2_X1 U826 ( .A1(n1153), .A2(n1152), .ZN(n1149) );
XNOR2_X1 U827 ( .A(n1154), .B(n1155), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1156), .B(KEYINPUT45), .Z(n1154) );
NAND2_X1 U829 ( .A1(G953), .A2(n1147), .ZN(n1148) );
NAND2_X1 U830 ( .A1(n1145), .A2(n1157), .ZN(n1140) );
NOR2_X1 U831 ( .A1(n1158), .A2(n1159), .ZN(G66) );
NOR3_X1 U832 ( .A1(n1123), .A2(n1160), .A3(n1161), .ZN(n1159) );
NOR3_X1 U833 ( .A1(n1162), .A2(n1125), .A3(n1163), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
NOR2_X1 U835 ( .A1(n1073), .A2(n1125), .ZN(n1164) );
NOR3_X1 U836 ( .A1(n1158), .A2(n1166), .A3(n1167), .ZN(G63) );
NOR3_X1 U837 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
INV_X1 U839 ( .A(KEYINPUT8), .ZN(n1172) );
NOR2_X1 U840 ( .A1(n1173), .A2(n1174), .ZN(n1166) );
NOR2_X1 U841 ( .A1(KEYINPUT8), .A2(n1171), .ZN(n1173) );
XOR2_X1 U842 ( .A(n1169), .B(KEYINPUT13), .Z(n1171) );
AND2_X1 U843 ( .A1(n1175), .A2(G478), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1158), .A2(n1176), .ZN(G60) );
XNOR2_X1 U845 ( .A(n1177), .B(n1178), .ZN(n1176) );
AND2_X1 U846 ( .A1(G475), .A2(n1175), .ZN(n1178) );
XOR2_X1 U847 ( .A(G104), .B(n1179), .Z(G6) );
NOR2_X1 U848 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NOR2_X1 U849 ( .A1(n1182), .A2(n1183), .ZN(G57) );
XNOR2_X1 U850 ( .A(n1158), .B(KEYINPUT61), .ZN(n1183) );
XOR2_X1 U851 ( .A(n1184), .B(n1185), .Z(n1182) );
AND2_X1 U852 ( .A1(G472), .A2(n1175), .ZN(n1184) );
NOR2_X1 U853 ( .A1(n1158), .A2(n1186), .ZN(G54) );
XOR2_X1 U854 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U855 ( .A(n1138), .B(n1189), .ZN(n1188) );
XNOR2_X1 U856 ( .A(n1190), .B(n1191), .ZN(n1189) );
NOR2_X1 U857 ( .A1(KEYINPUT24), .A2(n1192), .ZN(n1191) );
NAND3_X1 U858 ( .A1(n1175), .A2(G469), .A3(KEYINPUT26), .ZN(n1190) );
XNOR2_X1 U859 ( .A(n1193), .B(n1194), .ZN(n1187) );
XNOR2_X1 U860 ( .A(n1195), .B(n1196), .ZN(n1194) );
NOR2_X1 U861 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XOR2_X1 U862 ( .A(n1199), .B(KEYINPUT50), .Z(n1198) );
NAND2_X1 U863 ( .A1(n1137), .A2(n1200), .ZN(n1199) );
NOR2_X1 U864 ( .A1(n1137), .A2(n1200), .ZN(n1197) );
NOR2_X1 U865 ( .A1(n1158), .A2(n1201), .ZN(G51) );
XOR2_X1 U866 ( .A(n1202), .B(n1203), .Z(n1201) );
XNOR2_X1 U867 ( .A(n1204), .B(n1205), .ZN(n1203) );
XNOR2_X1 U868 ( .A(n1206), .B(n1207), .ZN(n1202) );
NOR2_X1 U869 ( .A1(n1120), .A2(n1163), .ZN(n1207) );
INV_X1 U870 ( .A(n1175), .ZN(n1163) );
NOR2_X1 U871 ( .A1(n1208), .A2(n1073), .ZN(n1175) );
NOR2_X1 U872 ( .A1(n1157), .A2(n1131), .ZN(n1073) );
NAND4_X1 U873 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1131) );
AND4_X1 U874 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1212) );
NOR3_X1 U875 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1211) );
NOR2_X1 U876 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
XOR2_X1 U877 ( .A(n1222), .B(KEYINPUT29), .Z(n1221) );
NOR4_X1 U878 ( .A1(n1087), .A2(n1223), .A3(n1081), .A4(n1224), .ZN(n1218) );
AND2_X1 U879 ( .A1(n1223), .A2(n1225), .ZN(n1217) );
INV_X1 U880 ( .A(KEYINPUT56), .ZN(n1223) );
NAND4_X1 U881 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1157) );
NOR2_X1 U882 ( .A1(n1230), .A2(n1066), .ZN(n1228) );
NOR2_X1 U883 ( .A1(n1231), .A2(n1180), .ZN(n1066) );
OR3_X1 U884 ( .A1(n1232), .A2(n1085), .A3(n1233), .ZN(n1180) );
NOR2_X1 U885 ( .A1(n1234), .A2(n1232), .ZN(n1230) );
INV_X1 U886 ( .A(n1235), .ZN(n1232) );
NOR3_X1 U887 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1234) );
NOR3_X1 U888 ( .A1(n1239), .A2(n1231), .A3(n1081), .ZN(n1238) );
INV_X1 U889 ( .A(n1098), .ZN(n1231) );
NOR3_X1 U890 ( .A1(n1181), .A2(n1240), .A3(n1085), .ZN(n1237) );
XNOR2_X1 U891 ( .A(n1102), .B(KEYINPUT34), .ZN(n1240) );
NOR2_X1 U892 ( .A1(n1241), .A2(n1079), .ZN(n1236) );
INV_X1 U893 ( .A(n1242), .ZN(n1079) );
NOR2_X1 U894 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
NOR2_X1 U895 ( .A1(n1239), .A2(n1245), .ZN(n1243) );
XNOR2_X1 U896 ( .A(KEYINPUT42), .B(n1233), .ZN(n1245) );
NAND3_X1 U897 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(n1226) );
XNOR2_X1 U898 ( .A(n1087), .B(KEYINPUT15), .ZN(n1248) );
INV_X1 U899 ( .A(n1249), .ZN(n1247) );
NOR2_X1 U900 ( .A1(n1145), .A2(G952), .ZN(n1158) );
NAND2_X1 U901 ( .A1(n1250), .A2(n1251), .ZN(G48) );
OR2_X1 U902 ( .A1(n1209), .A2(G146), .ZN(n1251) );
XOR2_X1 U903 ( .A(n1252), .B(KEYINPUT49), .Z(n1250) );
NAND2_X1 U904 ( .A1(G146), .A2(n1209), .ZN(n1252) );
NAND3_X1 U905 ( .A1(n1099), .A2(n1087), .A3(n1253), .ZN(n1209) );
XNOR2_X1 U906 ( .A(n1254), .B(n1255), .ZN(G45) );
NOR2_X1 U907 ( .A1(n1220), .A2(n1222), .ZN(n1255) );
NAND3_X1 U908 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1222) );
XNOR2_X1 U909 ( .A(G140), .B(n1210), .ZN(G42) );
OR3_X1 U910 ( .A1(n1091), .A2(n1233), .A3(n1224), .ZN(n1210) );
XNOR2_X1 U911 ( .A(G137), .B(n1216), .ZN(G39) );
NAND3_X1 U912 ( .A1(n1253), .A2(n1242), .A3(n1259), .ZN(n1216) );
XNOR2_X1 U913 ( .A(G134), .B(n1215), .ZN(G36) );
NAND3_X1 U914 ( .A1(n1258), .A2(n1098), .A3(n1259), .ZN(n1215) );
XNOR2_X1 U915 ( .A(G131), .B(n1214), .ZN(G33) );
NAND3_X1 U916 ( .A1(n1258), .A2(n1099), .A3(n1259), .ZN(n1214) );
INV_X1 U917 ( .A(n1091), .ZN(n1259) );
NAND2_X1 U918 ( .A1(n1260), .A2(n1089), .ZN(n1091) );
XNOR2_X1 U919 ( .A(KEYINPUT22), .B(n1088), .ZN(n1260) );
AND3_X1 U920 ( .A1(n1093), .A2(n1102), .A3(n1261), .ZN(n1258) );
NAND2_X1 U921 ( .A1(n1262), .A2(n1263), .ZN(G30) );
NAND2_X1 U922 ( .A1(G128), .A2(n1213), .ZN(n1263) );
XOR2_X1 U923 ( .A(n1264), .B(KEYINPUT32), .Z(n1262) );
OR2_X1 U924 ( .A1(n1213), .A2(G128), .ZN(n1264) );
NAND3_X1 U925 ( .A1(n1098), .A2(n1087), .A3(n1253), .ZN(n1213) );
AND4_X1 U926 ( .A1(n1265), .A2(n1261), .A3(n1102), .A4(n1111), .ZN(n1253) );
XNOR2_X1 U927 ( .A(G101), .B(n1266), .ZN(G3) );
NAND4_X1 U928 ( .A1(n1267), .A2(n1268), .A3(n1242), .A4(n1269), .ZN(n1266) );
NOR2_X1 U929 ( .A1(n1233), .A2(n1239), .ZN(n1269) );
INV_X1 U930 ( .A(n1102), .ZN(n1233) );
OR2_X1 U931 ( .A1(n1235), .A2(KEYINPUT52), .ZN(n1268) );
NAND2_X1 U932 ( .A1(KEYINPUT52), .A2(n1270), .ZN(n1267) );
NAND2_X1 U933 ( .A1(n1087), .A2(n1249), .ZN(n1270) );
XNOR2_X1 U934 ( .A(n1271), .B(n1225), .ZN(G27) );
NOR3_X1 U935 ( .A1(n1081), .A2(n1220), .A3(n1224), .ZN(n1225) );
NAND4_X1 U936 ( .A1(n1261), .A2(n1099), .A3(n1272), .A4(n1273), .ZN(n1224) );
AND2_X1 U937 ( .A1(n1274), .A2(n1076), .ZN(n1261) );
NAND2_X1 U938 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND2_X1 U939 ( .A1(n1134), .A2(G902), .ZN(n1276) );
NOR2_X1 U940 ( .A1(n1145), .A2(G900), .ZN(n1134) );
XNOR2_X1 U941 ( .A(G122), .B(n1227), .ZN(G24) );
NAND4_X1 U942 ( .A1(n1256), .A2(n1277), .A3(n1278), .A4(n1235), .ZN(n1227) );
NOR2_X1 U943 ( .A1(n1115), .A2(n1085), .ZN(n1278) );
NAND2_X1 U944 ( .A1(n1279), .A2(n1273), .ZN(n1085) );
XNOR2_X1 U945 ( .A(KEYINPUT20), .B(n1280), .ZN(n1279) );
XNOR2_X1 U946 ( .A(G119), .B(n1281), .ZN(G21) );
NAND4_X1 U947 ( .A1(KEYINPUT28), .A2(n1244), .A3(n1242), .A4(n1235), .ZN(n1281) );
AND3_X1 U948 ( .A1(n1277), .A2(n1111), .A3(n1265), .ZN(n1244) );
XNOR2_X1 U949 ( .A(n1272), .B(KEYINPUT31), .ZN(n1265) );
XNOR2_X1 U950 ( .A(G116), .B(n1282), .ZN(G18) );
NAND4_X1 U951 ( .A1(n1093), .A2(n1277), .A3(n1283), .A4(n1098), .ZN(n1282) );
NOR2_X1 U952 ( .A1(n1256), .A2(n1115), .ZN(n1098) );
INV_X1 U953 ( .A(n1257), .ZN(n1115) );
NOR2_X1 U954 ( .A1(n1284), .A2(n1249), .ZN(n1283) );
XNOR2_X1 U955 ( .A(n1087), .B(KEYINPUT51), .ZN(n1284) );
INV_X1 U956 ( .A(n1220), .ZN(n1087) );
INV_X1 U957 ( .A(n1239), .ZN(n1093) );
XNOR2_X1 U958 ( .A(G113), .B(n1285), .ZN(G15) );
NAND2_X1 U959 ( .A1(n1246), .A2(n1235), .ZN(n1285) );
NOR3_X1 U960 ( .A1(n1081), .A2(n1181), .A3(n1239), .ZN(n1246) );
NAND2_X1 U961 ( .A1(n1280), .A2(n1111), .ZN(n1239) );
INV_X1 U962 ( .A(n1099), .ZN(n1181) );
NOR2_X1 U963 ( .A1(n1286), .A2(n1257), .ZN(n1099) );
INV_X1 U964 ( .A(n1277), .ZN(n1081) );
NOR2_X1 U965 ( .A1(n1103), .A2(n1109), .ZN(n1277) );
XNOR2_X1 U966 ( .A(G110), .B(n1229), .ZN(G12) );
NAND4_X1 U967 ( .A1(n1242), .A2(n1102), .A3(n1092), .A4(n1235), .ZN(n1229) );
NOR2_X1 U968 ( .A1(n1249), .A2(n1220), .ZN(n1235) );
NAND2_X1 U969 ( .A1(n1089), .A2(n1088), .ZN(n1220) );
NAND2_X1 U970 ( .A1(n1287), .A2(n1288), .ZN(n1088) );
NAND2_X1 U971 ( .A1(n1122), .A2(n1120), .ZN(n1288) );
XOR2_X1 U972 ( .A(n1289), .B(KEYINPUT14), .Z(n1287) );
OR2_X1 U973 ( .A1(n1120), .A2(n1122), .ZN(n1289) );
AND2_X1 U974 ( .A1(n1290), .A2(n1208), .ZN(n1122) );
XOR2_X1 U975 ( .A(n1291), .B(n1205), .Z(n1290) );
XNOR2_X1 U976 ( .A(n1271), .B(n1292), .ZN(n1205) );
XNOR2_X1 U977 ( .A(n1293), .B(n1294), .ZN(n1291) );
INV_X1 U978 ( .A(n1204), .ZN(n1294) );
XNOR2_X1 U979 ( .A(n1153), .B(n1295), .ZN(n1204) );
NOR2_X1 U980 ( .A1(n1296), .A2(KEYINPUT1), .ZN(n1295) );
NOR2_X1 U981 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U982 ( .A(KEYINPUT60), .B(n1299), .Z(n1298) );
AND2_X1 U983 ( .A1(n1300), .A2(n1155), .ZN(n1299) );
NOR2_X1 U984 ( .A1(n1155), .A2(n1300), .ZN(n1297) );
XNOR2_X1 U985 ( .A(n1156), .B(KEYINPUT33), .ZN(n1300) );
NAND3_X1 U986 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1156) );
NAND2_X1 U987 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
OR3_X1 U988 ( .A1(n1305), .A2(n1304), .A3(KEYINPUT25), .ZN(n1302) );
XNOR2_X1 U989 ( .A(n1306), .B(KEYINPUT35), .ZN(n1304) );
NAND2_X1 U990 ( .A1(KEYINPUT27), .A2(n1307), .ZN(n1305) );
NAND2_X1 U991 ( .A1(G101), .A2(KEYINPUT25), .ZN(n1301) );
AND2_X1 U992 ( .A1(n1308), .A2(n1309), .ZN(n1155) );
NAND3_X1 U993 ( .A1(G113), .A2(n1310), .A3(n1311), .ZN(n1309) );
INV_X1 U994 ( .A(KEYINPUT41), .ZN(n1311) );
NAND2_X1 U995 ( .A1(n1312), .A2(KEYINPUT41), .ZN(n1308) );
NAND2_X1 U996 ( .A1(n1313), .A2(n1314), .ZN(n1153) );
NAND2_X1 U997 ( .A1(G110), .A2(n1315), .ZN(n1314) );
XOR2_X1 U998 ( .A(KEYINPUT40), .B(n1316), .Z(n1313) );
NOR2_X1 U999 ( .A1(G110), .A2(n1315), .ZN(n1316) );
NAND2_X1 U1000 ( .A1(KEYINPUT58), .A2(n1206), .ZN(n1293) );
NOR2_X1 U1001 ( .A1(n1146), .A2(G953), .ZN(n1206) );
INV_X1 U1002 ( .A(G224), .ZN(n1146) );
NAND2_X1 U1003 ( .A1(G210), .A2(n1317), .ZN(n1120) );
NAND2_X1 U1004 ( .A1(G214), .A2(n1317), .ZN(n1089) );
NAND2_X1 U1005 ( .A1(n1318), .A2(n1208), .ZN(n1317) );
NAND2_X1 U1006 ( .A1(n1319), .A2(n1076), .ZN(n1249) );
NAND2_X1 U1007 ( .A1(G237), .A2(G234), .ZN(n1076) );
NAND2_X1 U1008 ( .A1(n1275), .A2(n1320), .ZN(n1319) );
NAND3_X1 U1009 ( .A1(G902), .A2(n1147), .A3(G953), .ZN(n1320) );
INV_X1 U1010 ( .A(G898), .ZN(n1147) );
NAND2_X1 U1011 ( .A1(G952), .A2(n1321), .ZN(n1275) );
INV_X1 U1012 ( .A(n1072), .ZN(n1321) );
XOR2_X1 U1013 ( .A(G953), .B(KEYINPUT10), .Z(n1072) );
NOR2_X1 U1014 ( .A1(n1322), .A2(n1280), .ZN(n1092) );
INV_X1 U1015 ( .A(n1272), .ZN(n1280) );
XNOR2_X1 U1016 ( .A(n1123), .B(n1125), .ZN(n1272) );
NAND2_X1 U1017 ( .A1(G217), .A2(n1323), .ZN(n1125) );
NOR2_X1 U1018 ( .A1(n1165), .A2(G902), .ZN(n1123) );
INV_X1 U1019 ( .A(n1162), .ZN(n1165) );
XNOR2_X1 U1020 ( .A(n1324), .B(n1325), .ZN(n1162) );
XOR2_X1 U1021 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1022 ( .A(G137), .B(n1195), .ZN(n1327) );
NOR3_X1 U1023 ( .A1(KEYINPUT16), .A2(n1328), .A3(n1329), .ZN(n1326) );
NOR2_X1 U1024 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
XNOR2_X1 U1025 ( .A(n1332), .B(n1333), .ZN(n1331) );
NAND2_X1 U1026 ( .A1(n1334), .A2(n1271), .ZN(n1332) );
INV_X1 U1027 ( .A(KEYINPUT48), .ZN(n1330) );
NOR2_X1 U1028 ( .A1(KEYINPUT48), .A2(n1335), .ZN(n1328) );
XNOR2_X1 U1029 ( .A(n1333), .B(n1336), .ZN(n1335) );
XOR2_X1 U1030 ( .A(n1337), .B(n1338), .Z(n1324) );
NOR2_X1 U1031 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
INV_X1 U1032 ( .A(G221), .ZN(n1340) );
NAND2_X1 U1033 ( .A1(n1341), .A2(KEYINPUT0), .ZN(n1337) );
XOR2_X1 U1034 ( .A(n1342), .B(G128), .Z(n1341) );
NAND2_X1 U1035 ( .A1(KEYINPUT21), .A2(n1343), .ZN(n1342) );
INV_X1 U1036 ( .A(G119), .ZN(n1343) );
INV_X1 U1037 ( .A(n1273), .ZN(n1322) );
XOR2_X1 U1038 ( .A(n1111), .B(KEYINPUT11), .Z(n1273) );
XNOR2_X1 U1039 ( .A(n1344), .B(G472), .ZN(n1111) );
NAND3_X1 U1040 ( .A1(n1345), .A2(n1346), .A3(n1208), .ZN(n1344) );
NAND2_X1 U1041 ( .A1(n1185), .A2(n1347), .ZN(n1346) );
INV_X1 U1042 ( .A(KEYINPUT19), .ZN(n1347) );
XOR2_X1 U1043 ( .A(n1348), .B(n1349), .Z(n1185) );
NAND3_X1 U1044 ( .A1(n1348), .A2(n1349), .A3(KEYINPUT19), .ZN(n1345) );
XNOR2_X1 U1045 ( .A(n1312), .B(n1350), .ZN(n1349) );
XNOR2_X1 U1046 ( .A(n1292), .B(n1138), .ZN(n1350) );
INV_X1 U1047 ( .A(n1351), .ZN(n1138) );
XOR2_X1 U1048 ( .A(G128), .B(n1352), .Z(n1292) );
NOR2_X1 U1049 ( .A1(n1353), .A2(n1354), .ZN(n1352) );
NOR2_X1 U1050 ( .A1(KEYINPUT12), .A2(n1355), .ZN(n1354) );
AND2_X1 U1051 ( .A1(KEYINPUT46), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1052 ( .A(G113), .B(n1310), .Z(n1312) );
XNOR2_X1 U1053 ( .A(n1356), .B(G119), .ZN(n1310) );
INV_X1 U1054 ( .A(G116), .ZN(n1356) );
XNOR2_X1 U1055 ( .A(n1357), .B(n1307), .ZN(n1348) );
INV_X1 U1056 ( .A(G101), .ZN(n1307) );
NAND3_X1 U1057 ( .A1(n1318), .A2(n1145), .A3(G210), .ZN(n1357) );
NOR2_X1 U1058 ( .A1(n1358), .A2(n1109), .ZN(n1102) );
INV_X1 U1059 ( .A(n1104), .ZN(n1109) );
NAND2_X1 U1060 ( .A1(G221), .A2(n1323), .ZN(n1104) );
NAND2_X1 U1061 ( .A1(G234), .A2(n1208), .ZN(n1323) );
INV_X1 U1062 ( .A(n1103), .ZN(n1358) );
XOR2_X1 U1063 ( .A(G469), .B(n1359), .Z(n1103) );
NOR2_X1 U1064 ( .A1(KEYINPUT53), .A2(n1116), .ZN(n1359) );
NAND2_X1 U1065 ( .A1(n1360), .A2(n1208), .ZN(n1116) );
XOR2_X1 U1066 ( .A(n1361), .B(n1362), .Z(n1360) );
XNOR2_X1 U1067 ( .A(n1137), .B(n1200), .ZN(n1362) );
XOR2_X1 U1068 ( .A(G101), .B(n1306), .Z(n1200) );
XOR2_X1 U1069 ( .A(G104), .B(G107), .Z(n1306) );
XOR2_X1 U1070 ( .A(n1363), .B(G128), .Z(n1137) );
NAND2_X1 U1071 ( .A1(KEYINPUT47), .A2(n1364), .ZN(n1363) );
INV_X1 U1072 ( .A(n1355), .ZN(n1364) );
XNOR2_X1 U1073 ( .A(G143), .B(n1333), .ZN(n1355) );
XNOR2_X1 U1074 ( .A(n1351), .B(n1365), .ZN(n1361) );
XOR2_X1 U1075 ( .A(n1193), .B(n1366), .Z(n1365) );
NOR2_X1 U1076 ( .A1(KEYINPUT54), .A2(n1367), .ZN(n1366) );
XOR2_X1 U1077 ( .A(n1368), .B(n1192), .Z(n1367) );
XOR2_X1 U1078 ( .A(G140), .B(KEYINPUT39), .Z(n1192) );
NOR2_X1 U1079 ( .A1(KEYINPUT59), .A2(n1195), .ZN(n1368) );
INV_X1 U1080 ( .A(G110), .ZN(n1195) );
NAND2_X1 U1081 ( .A1(G227), .A2(n1145), .ZN(n1193) );
XOR2_X1 U1082 ( .A(G131), .B(n1369), .Z(n1351) );
XOR2_X1 U1083 ( .A(G137), .B(G134), .Z(n1369) );
NOR2_X1 U1084 ( .A1(n1257), .A2(n1256), .ZN(n1242) );
INV_X1 U1085 ( .A(n1286), .ZN(n1256) );
XOR2_X1 U1086 ( .A(n1112), .B(KEYINPUT9), .Z(n1286) );
XNOR2_X1 U1087 ( .A(n1370), .B(G475), .ZN(n1112) );
NAND2_X1 U1088 ( .A1(n1177), .A2(n1208), .ZN(n1370) );
XNOR2_X1 U1089 ( .A(n1371), .B(n1372), .ZN(n1177) );
XNOR2_X1 U1090 ( .A(n1315), .B(G104), .ZN(n1372) );
XOR2_X1 U1091 ( .A(n1373), .B(n1374), .Z(n1371) );
NOR2_X1 U1092 ( .A1(KEYINPUT63), .A2(n1375), .ZN(n1374) );
XNOR2_X1 U1093 ( .A(G113), .B(KEYINPUT23), .ZN(n1375) );
NAND2_X1 U1094 ( .A1(n1376), .A2(n1377), .ZN(n1373) );
NAND2_X1 U1095 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
INV_X1 U1096 ( .A(n1380), .ZN(n1379) );
NAND2_X1 U1097 ( .A1(n1381), .A2(n1382), .ZN(n1378) );
NAND2_X1 U1098 ( .A1(n1383), .A2(n1333), .ZN(n1382) );
NAND2_X1 U1099 ( .A1(n1384), .A2(G146), .ZN(n1381) );
NAND2_X1 U1100 ( .A1(n1380), .A2(n1385), .ZN(n1376) );
NAND2_X1 U1101 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
NAND2_X1 U1102 ( .A1(n1383), .A2(G146), .ZN(n1387) );
NAND2_X1 U1103 ( .A1(n1384), .A2(n1333), .ZN(n1386) );
INV_X1 U1104 ( .A(G146), .ZN(n1333) );
XNOR2_X1 U1105 ( .A(n1383), .B(n1388), .ZN(n1384) );
XOR2_X1 U1106 ( .A(KEYINPUT55), .B(KEYINPUT17), .Z(n1388) );
XNOR2_X1 U1107 ( .A(G131), .B(n1389), .ZN(n1383) );
NOR2_X1 U1108 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
XOR2_X1 U1109 ( .A(KEYINPUT57), .B(n1392), .Z(n1391) );
NOR2_X1 U1110 ( .A1(n1393), .A2(n1394), .ZN(n1392) );
XNOR2_X1 U1111 ( .A(G143), .B(KEYINPUT6), .ZN(n1393) );
AND2_X1 U1112 ( .A1(n1254), .A2(n1394), .ZN(n1390) );
NAND3_X1 U1113 ( .A1(n1318), .A2(n1145), .A3(n1395), .ZN(n1394) );
XNOR2_X1 U1114 ( .A(G214), .B(KEYINPUT38), .ZN(n1395) );
INV_X1 U1115 ( .A(G237), .ZN(n1318) );
NOR2_X1 U1116 ( .A1(KEYINPUT62), .A2(n1336), .ZN(n1380) );
XNOR2_X1 U1117 ( .A(n1271), .B(n1334), .ZN(n1336) );
XOR2_X1 U1118 ( .A(G140), .B(KEYINPUT36), .Z(n1334) );
INV_X1 U1119 ( .A(G125), .ZN(n1271) );
XNOR2_X1 U1120 ( .A(n1396), .B(G478), .ZN(n1257) );
NAND2_X1 U1121 ( .A1(n1168), .A2(n1208), .ZN(n1396) );
INV_X1 U1122 ( .A(G902), .ZN(n1208) );
INV_X1 U1123 ( .A(n1174), .ZN(n1168) );
XNOR2_X1 U1124 ( .A(n1397), .B(n1398), .ZN(n1174) );
XOR2_X1 U1125 ( .A(n1399), .B(n1400), .Z(n1398) );
XOR2_X1 U1126 ( .A(G107), .B(n1401), .Z(n1400) );
NOR2_X1 U1127 ( .A1(KEYINPUT3), .A2(n1402), .ZN(n1401) );
XNOR2_X1 U1128 ( .A(n1254), .B(G128), .ZN(n1402) );
INV_X1 U1129 ( .A(G143), .ZN(n1254) );
NOR2_X1 U1130 ( .A1(n1339), .A2(n1403), .ZN(n1399) );
INV_X1 U1131 ( .A(G217), .ZN(n1403) );
NAND2_X1 U1132 ( .A1(G234), .A2(n1145), .ZN(n1339) );
INV_X1 U1133 ( .A(G953), .ZN(n1145) );
XNOR2_X1 U1134 ( .A(G116), .B(n1404), .ZN(n1397) );
XNOR2_X1 U1135 ( .A(G134), .B(n1315), .ZN(n1404) );
INV_X1 U1136 ( .A(G122), .ZN(n1315) );
endmodule


