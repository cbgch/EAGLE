//Key = 0010010000010100010100111000000110101001100010001011111101000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280;

XOR2_X1 U700 ( .A(n973), .B(n974), .Z(G9) );
NOR2_X1 U701 ( .A1(KEYINPUT4), .A2(n975), .ZN(n974) );
NOR2_X1 U702 ( .A1(n976), .A2(n977), .ZN(G75) );
NOR3_X1 U703 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n977) );
NOR3_X1 U704 ( .A1(n981), .A2(n982), .A3(n983), .ZN(n979) );
NOR2_X1 U705 ( .A1(n984), .A2(n985), .ZN(n983) );
NOR2_X1 U706 ( .A1(n986), .A2(n987), .ZN(n985) );
NOR2_X1 U707 ( .A1(n988), .A2(n989), .ZN(n986) );
XOR2_X1 U708 ( .A(KEYINPUT61), .B(n990), .Z(n989) );
NOR2_X1 U709 ( .A1(n991), .A2(n992), .ZN(n990) );
XOR2_X1 U710 ( .A(n993), .B(n994), .Z(n992) );
XOR2_X1 U711 ( .A(n995), .B(KEYINPUT63), .Z(n991) );
NOR3_X1 U712 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n984) );
NOR4_X1 U713 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(n998) );
NOR2_X1 U714 ( .A1(KEYINPUT8), .A2(n1003), .ZN(n1002) );
AND3_X1 U715 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1001) );
NOR2_X1 U716 ( .A1(n1007), .A2(n1008), .ZN(n1000) );
NOR2_X1 U717 ( .A1(n1009), .A2(n1010), .ZN(n997) );
NOR2_X1 U718 ( .A1(n1003), .A2(n1011), .ZN(n1010) );
INV_X1 U719 ( .A(KEYINPUT8), .ZN(n1011) );
NAND3_X1 U720 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n978) );
NAND3_X1 U721 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
INV_X1 U722 ( .A(n987), .ZN(n1017) );
NAND3_X1 U723 ( .A1(n1009), .A2(n1018), .A3(n1004), .ZN(n987) );
INV_X1 U724 ( .A(n999), .ZN(n1009) );
NAND2_X1 U725 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
NAND2_X1 U726 ( .A1(n982), .A2(n1021), .ZN(n1020) );
AND3_X1 U727 ( .A1(n1012), .A2(n1013), .A3(n1022), .ZN(n976) );
NAND4_X1 U728 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1012) );
NOR4_X1 U729 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
XOR2_X1 U730 ( .A(n1031), .B(n1032), .Z(n1030) );
XOR2_X1 U731 ( .A(G475), .B(n1033), .Z(n1029) );
XOR2_X1 U732 ( .A(n1034), .B(n1035), .Z(n1028) );
NOR3_X1 U733 ( .A1(n1036), .A2(n1037), .A3(n982), .ZN(n1025) );
XOR2_X1 U734 ( .A(KEYINPUT23), .B(n981), .Z(n1024) );
XOR2_X1 U735 ( .A(n1038), .B(n1039), .Z(G72) );
XOR2_X1 U736 ( .A(n1040), .B(n1041), .Z(n1039) );
NOR3_X1 U737 ( .A1(n1042), .A2(KEYINPUT43), .A3(n1043), .ZN(n1041) );
NOR2_X1 U738 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
XOR2_X1 U739 ( .A(n1046), .B(KEYINPUT17), .Z(n1044) );
XOR2_X1 U740 ( .A(KEYINPUT45), .B(G953), .Z(n1042) );
NOR2_X1 U741 ( .A1(n1047), .A2(n1048), .ZN(n1040) );
XNOR2_X1 U742 ( .A(n1049), .B(n1050), .ZN(n1048) );
XOR2_X1 U743 ( .A(n1051), .B(KEYINPUT28), .Z(n1050) );
NAND2_X1 U744 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U745 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U746 ( .A(n1056), .B(KEYINPUT15), .Z(n1052) );
OR2_X1 U747 ( .A1(n1054), .A2(n1055), .ZN(n1056) );
XNOR2_X1 U748 ( .A(n1057), .B(n1058), .ZN(n1054) );
XNOR2_X1 U749 ( .A(n1059), .B(KEYINPUT36), .ZN(n1058) );
NAND2_X1 U750 ( .A1(KEYINPUT54), .A2(n1060), .ZN(n1059) );
XNOR2_X1 U751 ( .A(n1061), .B(KEYINPUT40), .ZN(n1047) );
NOR2_X1 U752 ( .A1(n1062), .A2(n1013), .ZN(n1038) );
AND2_X1 U753 ( .A1(G227), .A2(G900), .ZN(n1062) );
XOR2_X1 U754 ( .A(n1063), .B(n1064), .Z(G69) );
XOR2_X1 U755 ( .A(n1065), .B(n1066), .Z(n1064) );
NOR2_X1 U756 ( .A1(n1067), .A2(G953), .ZN(n1066) );
NOR2_X1 U757 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XOR2_X1 U758 ( .A(n1070), .B(KEYINPUT22), .Z(n1068) );
NAND2_X1 U759 ( .A1(n1071), .A2(n1072), .ZN(n1065) );
NAND2_X1 U760 ( .A1(G953), .A2(n1073), .ZN(n1072) );
XOR2_X1 U761 ( .A(n1074), .B(n1075), .Z(n1071) );
XOR2_X1 U762 ( .A(n1076), .B(n1077), .Z(n1075) );
NOR2_X1 U763 ( .A1(KEYINPUT7), .A2(n1078), .ZN(n1076) );
NAND2_X1 U764 ( .A1(G953), .A2(n1079), .ZN(n1063) );
NAND2_X1 U765 ( .A1(G898), .A2(G224), .ZN(n1079) );
NOR2_X1 U766 ( .A1(n1080), .A2(n1081), .ZN(G66) );
XOR2_X1 U767 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U769 ( .A1(n1080), .A2(n1086), .ZN(G63) );
XOR2_X1 U770 ( .A(n1087), .B(n1088), .Z(n1086) );
XOR2_X1 U771 ( .A(KEYINPUT5), .B(n1089), .Z(n1088) );
NOR2_X1 U772 ( .A1(n1090), .A2(n1085), .ZN(n1089) );
INV_X1 U773 ( .A(G478), .ZN(n1090) );
NOR2_X1 U774 ( .A1(n1080), .A2(n1091), .ZN(G60) );
XOR2_X1 U775 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR2_X1 U776 ( .A1(n1094), .A2(n1085), .ZN(n1092) );
XNOR2_X1 U777 ( .A(G104), .B(n1095), .ZN(G6) );
NAND4_X1 U778 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1018), .ZN(n1095) );
AND2_X1 U779 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U780 ( .A(n1101), .B(KEYINPUT57), .Z(n1096) );
NOR2_X1 U781 ( .A1(n1080), .A2(n1102), .ZN(G57) );
XOR2_X1 U782 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U783 ( .A(G101), .B(n1105), .Z(n1104) );
NOR2_X1 U784 ( .A1(n1031), .A2(n1085), .ZN(n1105) );
INV_X1 U785 ( .A(G472), .ZN(n1031) );
NOR2_X1 U786 ( .A1(n1080), .A2(n1106), .ZN(G54) );
XOR2_X1 U787 ( .A(n1107), .B(n1108), .Z(n1106) );
NOR2_X1 U788 ( .A1(n1109), .A2(n1085), .ZN(n1107) );
INV_X1 U789 ( .A(G469), .ZN(n1109) );
NOR2_X1 U790 ( .A1(n1080), .A2(n1110), .ZN(G51) );
XOR2_X1 U791 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U792 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U793 ( .A1(n1115), .A2(n1085), .ZN(n1113) );
NAND2_X1 U794 ( .A1(G902), .A2(n980), .ZN(n1085) );
NAND4_X1 U795 ( .A1(n1116), .A2(n1117), .A3(n1046), .A4(n1070), .ZN(n980) );
INV_X1 U796 ( .A(n1045), .ZN(n1117) );
NAND4_X1 U797 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1045) );
NOR3_X1 U798 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
OR2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(n1120) );
NAND2_X1 U800 ( .A1(n1127), .A2(n1015), .ZN(n1119) );
XOR2_X1 U801 ( .A(KEYINPUT33), .B(n1128), .Z(n1127) );
NOR4_X1 U802 ( .A1(n1129), .A2(n1019), .A3(n1130), .A4(n1131), .ZN(n1128) );
XNOR2_X1 U803 ( .A(KEYINPUT56), .B(n1132), .ZN(n1131) );
INV_X1 U804 ( .A(n1100), .ZN(n1019) );
OR2_X1 U805 ( .A1(n1133), .A2(n1007), .ZN(n1118) );
INV_X1 U806 ( .A(n1134), .ZN(n1007) );
INV_X1 U807 ( .A(n1069), .ZN(n1116) );
NAND4_X1 U808 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1069) );
NOR2_X1 U809 ( .A1(n973), .A2(n1139), .ZN(n1137) );
NOR3_X1 U810 ( .A1(n1126), .A2(n1140), .A3(n1008), .ZN(n973) );
NAND3_X1 U811 ( .A1(n1141), .A2(n1134), .A3(n1142), .ZN(n1136) );
NAND2_X1 U812 ( .A1(n1130), .A2(n1126), .ZN(n1134) );
NAND2_X1 U813 ( .A1(n1143), .A2(n1144), .ZN(n1135) );
NAND2_X1 U814 ( .A1(n1003), .A2(n1145), .ZN(n1144) );
NAND2_X1 U815 ( .A1(n1097), .A2(n1018), .ZN(n1145) );
AND2_X1 U816 ( .A1(n1146), .A2(n1022), .ZN(n1080) );
INV_X1 U817 ( .A(G952), .ZN(n1022) );
XOR2_X1 U818 ( .A(n1013), .B(KEYINPUT32), .Z(n1146) );
XOR2_X1 U819 ( .A(G146), .B(n1147), .Z(G48) );
NOR2_X1 U820 ( .A1(n1130), .A2(n1133), .ZN(n1147) );
NAND2_X1 U821 ( .A1(n1148), .A2(n1149), .ZN(G45) );
NAND2_X1 U822 ( .A1(n1122), .A2(n1150), .ZN(n1149) );
INV_X1 U823 ( .A(n1151), .ZN(n1122) );
XOR2_X1 U824 ( .A(n1152), .B(KEYINPUT10), .Z(n1148) );
NAND2_X1 U825 ( .A1(G143), .A2(n1151), .ZN(n1152) );
NAND4_X1 U826 ( .A1(n1141), .A2(n1153), .A3(n988), .A4(n1154), .ZN(n1151) );
NOR2_X1 U827 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U828 ( .A(G140), .B(n1124), .Z(G42) );
AND2_X1 U829 ( .A1(n1157), .A2(n1158), .ZN(n1124) );
XOR2_X1 U830 ( .A(n1060), .B(n1046), .Z(G39) );
NAND3_X1 U831 ( .A1(n1158), .A2(n1004), .A3(n1159), .ZN(n1046) );
XOR2_X1 U832 ( .A(G134), .B(n1160), .Z(G36) );
NOR2_X1 U833 ( .A1(n1161), .A2(n1125), .ZN(n1160) );
XOR2_X1 U834 ( .A(n1126), .B(KEYINPUT18), .Z(n1161) );
XOR2_X1 U835 ( .A(G131), .B(n1162), .Z(G33) );
NOR2_X1 U836 ( .A1(n1130), .A2(n1125), .ZN(n1162) );
NAND2_X1 U837 ( .A1(n1158), .A2(n1141), .ZN(n1125) );
NOR2_X1 U838 ( .A1(n1155), .A2(n996), .ZN(n1158) );
INV_X1 U839 ( .A(n1015), .ZN(n996) );
NAND2_X1 U840 ( .A1(n1163), .A2(n1164), .ZN(n1015) );
NAND3_X1 U841 ( .A1(n994), .A2(n995), .A3(n993), .ZN(n1164) );
INV_X1 U842 ( .A(KEYINPUT35), .ZN(n993) );
NAND2_X1 U843 ( .A1(KEYINPUT35), .A2(n988), .ZN(n1163) );
XOR2_X1 U844 ( .A(G128), .B(n1165), .Z(G30) );
NOR2_X1 U845 ( .A1(n1133), .A2(n1166), .ZN(n1165) );
XNOR2_X1 U846 ( .A(KEYINPUT34), .B(n1126), .ZN(n1166) );
NAND3_X1 U847 ( .A1(n1167), .A2(n988), .A3(n1159), .ZN(n1133) );
INV_X1 U848 ( .A(n1155), .ZN(n1167) );
NAND2_X1 U849 ( .A1(n1100), .A2(n1132), .ZN(n1155) );
XOR2_X1 U850 ( .A(G101), .B(n1168), .Z(G3) );
NOR3_X1 U851 ( .A1(n1003), .A2(KEYINPUT62), .A3(n1140), .ZN(n1168) );
NAND2_X1 U852 ( .A1(n1004), .A2(n1141), .ZN(n1003) );
XNOR2_X1 U853 ( .A(n1123), .B(n1169), .ZN(G27) );
XOR2_X1 U854 ( .A(KEYINPUT39), .B(G125), .Z(n1169) );
AND3_X1 U855 ( .A1(n1170), .A2(n1132), .A3(n1157), .ZN(n1123) );
NOR3_X1 U856 ( .A1(n1171), .A2(n1172), .A3(n1130), .ZN(n1157) );
INV_X1 U857 ( .A(n1097), .ZN(n1130) );
NAND2_X1 U858 ( .A1(n999), .A2(n1173), .ZN(n1132) );
NAND3_X1 U859 ( .A1(G902), .A2(n1174), .A3(n1061), .ZN(n1173) );
NOR2_X1 U860 ( .A1(n1013), .A2(G900), .ZN(n1061) );
XOR2_X1 U861 ( .A(n1175), .B(n1138), .Z(G24) );
NAND4_X1 U862 ( .A1(n1176), .A2(n1142), .A3(n1018), .A4(n1153), .ZN(n1138) );
XOR2_X1 U863 ( .A(G119), .B(n1139), .Z(G21) );
AND3_X1 U864 ( .A1(n1159), .A2(n1004), .A3(n1142), .ZN(n1139) );
AND2_X1 U865 ( .A1(n1177), .A2(n1005), .ZN(n1159) );
XOR2_X1 U866 ( .A(n1171), .B(KEYINPUT3), .Z(n1177) );
XOR2_X1 U867 ( .A(G116), .B(n1178), .Z(G18) );
NOR4_X1 U868 ( .A1(KEYINPUT21), .A2(n1129), .A3(n1126), .A4(n1179), .ZN(n1178) );
NAND2_X1 U869 ( .A1(n1156), .A2(n1153), .ZN(n1126) );
INV_X1 U870 ( .A(n1141), .ZN(n1129) );
XOR2_X1 U871 ( .A(n1180), .B(n1181), .Z(G15) );
XOR2_X1 U872 ( .A(KEYINPUT24), .B(G113), .Z(n1181) );
NAND3_X1 U873 ( .A1(n1182), .A2(n1142), .A3(n1097), .ZN(n1180) );
NOR2_X1 U874 ( .A1(n1156), .A2(n1153), .ZN(n1097) );
INV_X1 U875 ( .A(n1176), .ZN(n1156) );
INV_X1 U876 ( .A(n1179), .ZN(n1142) );
NAND2_X1 U877 ( .A1(n1170), .A2(n1099), .ZN(n1179) );
NOR3_X1 U878 ( .A1(n1101), .A2(n982), .A3(n981), .ZN(n1170) );
INV_X1 U879 ( .A(n1021), .ZN(n981) );
INV_X1 U880 ( .A(n988), .ZN(n1101) );
XOR2_X1 U881 ( .A(n1141), .B(KEYINPUT37), .Z(n1182) );
NAND2_X1 U882 ( .A1(n1183), .A2(n1184), .ZN(n1141) );
OR3_X1 U883 ( .A1(n1005), .A2(n1006), .A3(KEYINPUT3), .ZN(n1184) );
NAND2_X1 U884 ( .A1(KEYINPUT3), .A2(n1018), .ZN(n1183) );
INV_X1 U885 ( .A(n1008), .ZN(n1018) );
NAND2_X1 U886 ( .A1(n1006), .A2(n1172), .ZN(n1008) );
XOR2_X1 U887 ( .A(n1185), .B(n1070), .Z(G12) );
NAND4_X1 U888 ( .A1(n1004), .A2(n1143), .A3(n1006), .A4(n1005), .ZN(n1070) );
INV_X1 U889 ( .A(n1172), .ZN(n1005) );
NOR2_X1 U890 ( .A1(n1186), .A2(n1037), .ZN(n1172) );
NOR3_X1 U891 ( .A1(n1187), .A2(G902), .A3(n1082), .ZN(n1037) );
XNOR2_X1 U892 ( .A(KEYINPUT47), .B(n1023), .ZN(n1186) );
AND2_X1 U893 ( .A1(n1188), .A2(n1189), .ZN(n1023) );
NAND2_X1 U894 ( .A1(n1187), .A2(n1082), .ZN(n1189) );
XOR2_X1 U895 ( .A(n1190), .B(n1191), .Z(n1082) );
XOR2_X1 U896 ( .A(n1192), .B(n1193), .Z(n1191) );
AND2_X1 U897 ( .A1(n1194), .A2(G221), .ZN(n1192) );
XOR2_X1 U898 ( .A(n1195), .B(n1196), .Z(n1190) );
XOR2_X1 U899 ( .A(n1060), .B(n1197), .Z(n1196) );
NAND3_X1 U900 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1197) );
NAND2_X1 U901 ( .A1(KEYINPUT29), .A2(n1201), .ZN(n1200) );
NAND3_X1 U902 ( .A1(n1202), .A2(n1203), .A3(G128), .ZN(n1199) );
NAND2_X1 U903 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NAND2_X1 U904 ( .A1(n1206), .A2(n1203), .ZN(n1204) );
INV_X1 U905 ( .A(KEYINPUT29), .ZN(n1203) );
XOR2_X1 U906 ( .A(n1202), .B(KEYINPUT0), .Z(n1206) );
INV_X1 U907 ( .A(G137), .ZN(n1060) );
NAND2_X1 U908 ( .A1(KEYINPUT50), .A2(n1185), .ZN(n1195) );
NOR2_X1 U909 ( .A1(n1084), .A2(G234), .ZN(n1187) );
INV_X1 U910 ( .A(G217), .ZN(n1084) );
NAND2_X1 U911 ( .A1(G902), .A2(G217), .ZN(n1188) );
INV_X1 U912 ( .A(n1171), .ZN(n1006) );
NAND2_X1 U913 ( .A1(n1207), .A2(n1208), .ZN(n1171) );
NAND2_X1 U914 ( .A1(G472), .A2(n1032), .ZN(n1208) );
XOR2_X1 U915 ( .A(n1209), .B(KEYINPUT49), .Z(n1207) );
OR2_X1 U916 ( .A1(n1032), .A2(G472), .ZN(n1209) );
NAND2_X1 U917 ( .A1(n1210), .A2(n1211), .ZN(n1032) );
XOR2_X1 U918 ( .A(n1103), .B(n1212), .Z(n1210) );
XOR2_X1 U919 ( .A(KEYINPUT16), .B(n1213), .Z(n1212) );
NOR2_X1 U920 ( .A1(G101), .A2(KEYINPUT46), .ZN(n1213) );
XNOR2_X1 U921 ( .A(n1214), .B(n1215), .ZN(n1103) );
XOR2_X1 U922 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U923 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR3_X1 U924 ( .A1(n1115), .A2(G953), .A3(G237), .ZN(n1219) );
INV_X1 U925 ( .A(G210), .ZN(n1115) );
XOR2_X1 U926 ( .A(n1220), .B(n1201), .Z(n1214) );
INV_X1 U927 ( .A(n1202), .ZN(n1201) );
INV_X1 U928 ( .A(n1140), .ZN(n1143) );
NAND3_X1 U929 ( .A1(n988), .A2(n1099), .A3(n1100), .ZN(n1140) );
NOR2_X1 U930 ( .A1(n1021), .A2(n982), .ZN(n1100) );
AND2_X1 U931 ( .A1(G221), .A2(n1221), .ZN(n982) );
NAND2_X1 U932 ( .A1(G234), .A2(n1211), .ZN(n1221) );
XOR2_X1 U933 ( .A(n1222), .B(G469), .Z(n1021) );
NAND2_X1 U934 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XNOR2_X1 U935 ( .A(n1108), .B(KEYINPUT27), .ZN(n1224) );
XNOR2_X1 U936 ( .A(n1225), .B(n1226), .ZN(n1108) );
XOR2_X1 U937 ( .A(n1227), .B(n1228), .Z(n1226) );
XOR2_X1 U938 ( .A(G110), .B(n1229), .Z(n1228) );
AND2_X1 U939 ( .A1(n1013), .A2(G227), .ZN(n1229) );
XOR2_X1 U940 ( .A(KEYINPUT2), .B(G140), .Z(n1227) );
XOR2_X1 U941 ( .A(n1220), .B(n1230), .Z(n1225) );
XOR2_X1 U942 ( .A(n1078), .B(n1055), .Z(n1230) );
XOR2_X1 U943 ( .A(n1231), .B(n1232), .Z(n1055) );
NOR2_X1 U944 ( .A1(G128), .A2(KEYINPUT30), .ZN(n1232) );
XOR2_X1 U945 ( .A(n1057), .B(G137), .Z(n1220) );
XNOR2_X1 U946 ( .A(G131), .B(n1233), .ZN(n1057) );
XOR2_X1 U947 ( .A(n1211), .B(KEYINPUT42), .Z(n1223) );
NAND2_X1 U948 ( .A1(n999), .A2(n1234), .ZN(n1099) );
NAND4_X1 U949 ( .A1(G953), .A2(G902), .A3(n1174), .A4(n1073), .ZN(n1234) );
INV_X1 U950 ( .A(G898), .ZN(n1073) );
NAND3_X1 U951 ( .A1(n1174), .A2(n1013), .A3(G952), .ZN(n999) );
NAND2_X1 U952 ( .A1(G237), .A2(G234), .ZN(n1174) );
NOR2_X1 U953 ( .A1(n994), .A2(n1036), .ZN(n988) );
INV_X1 U954 ( .A(n995), .ZN(n1036) );
NAND2_X1 U955 ( .A1(G214), .A2(n1235), .ZN(n995) );
XOR2_X1 U956 ( .A(n1236), .B(n1035), .Z(n994) );
NAND2_X1 U957 ( .A1(n1237), .A2(n1211), .ZN(n1035) );
XOR2_X1 U958 ( .A(n1238), .B(n1114), .Z(n1237) );
XNOR2_X1 U959 ( .A(n1218), .B(n1239), .ZN(n1114) );
XOR2_X1 U960 ( .A(G125), .B(n1240), .Z(n1239) );
AND2_X1 U961 ( .A1(n1013), .A2(G224), .ZN(n1240) );
XOR2_X1 U962 ( .A(n1205), .B(n1231), .Z(n1218) );
XOR2_X1 U963 ( .A(n1241), .B(n1150), .Z(n1231) );
INV_X1 U964 ( .A(G143), .ZN(n1150) );
INV_X1 U965 ( .A(G146), .ZN(n1241) );
NAND2_X1 U966 ( .A1(KEYINPUT11), .A2(n1111), .ZN(n1238) );
NAND2_X1 U967 ( .A1(n1242), .A2(n1243), .ZN(n1111) );
NAND2_X1 U968 ( .A1(n1244), .A2(n1074), .ZN(n1243) );
XOR2_X1 U969 ( .A(KEYINPUT12), .B(n1245), .Z(n1244) );
NAND2_X1 U970 ( .A1(n1246), .A2(n1247), .ZN(n1242) );
INV_X1 U971 ( .A(n1074), .ZN(n1247) );
XOR2_X1 U972 ( .A(n1248), .B(n1249), .Z(n1074) );
INV_X1 U973 ( .A(n1216), .ZN(n1249) );
XNOR2_X1 U974 ( .A(G113), .B(G116), .ZN(n1216) );
NAND2_X1 U975 ( .A1(n1250), .A2(KEYINPUT55), .ZN(n1248) );
XOR2_X1 U976 ( .A(n1202), .B(KEYINPUT60), .Z(n1250) );
XNOR2_X1 U977 ( .A(G119), .B(KEYINPUT1), .ZN(n1202) );
XOR2_X1 U978 ( .A(n1245), .B(n1251), .Z(n1246) );
XOR2_X1 U979 ( .A(KEYINPUT38), .B(KEYINPUT31), .Z(n1251) );
XOR2_X1 U980 ( .A(n1078), .B(n1077), .Z(n1245) );
XOR2_X1 U981 ( .A(G110), .B(G122), .Z(n1077) );
XOR2_X1 U982 ( .A(G101), .B(n1252), .Z(n1078) );
XOR2_X1 U983 ( .A(G107), .B(G104), .Z(n1252) );
NAND2_X1 U984 ( .A1(KEYINPUT51), .A2(n1253), .ZN(n1236) );
XNOR2_X1 U985 ( .A(KEYINPUT44), .B(n1034), .ZN(n1253) );
NAND2_X1 U986 ( .A1(n1254), .A2(G210), .ZN(n1034) );
XOR2_X1 U987 ( .A(n1235), .B(KEYINPUT58), .Z(n1254) );
OR2_X1 U988 ( .A1(G902), .A2(G237), .ZN(n1235) );
NOR2_X1 U989 ( .A1(n1153), .A2(n1176), .ZN(n1004) );
XOR2_X1 U990 ( .A(n1255), .B(n1256), .Z(n1176) );
NOR2_X1 U991 ( .A1(KEYINPUT20), .A2(n1033), .ZN(n1256) );
NOR2_X1 U992 ( .A1(n1257), .A2(n1093), .ZN(n1033) );
XNOR2_X1 U993 ( .A(n1258), .B(n1259), .ZN(n1093) );
XOR2_X1 U994 ( .A(n1260), .B(n1261), .Z(n1259) );
XNOR2_X1 U995 ( .A(G104), .B(G131), .ZN(n1261) );
NAND2_X1 U996 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
XOR2_X1 U997 ( .A(G122), .B(G113), .Z(n1263) );
XNOR2_X1 U998 ( .A(KEYINPUT53), .B(KEYINPUT48), .ZN(n1262) );
XOR2_X1 U999 ( .A(n1264), .B(n1193), .Z(n1258) );
XOR2_X1 U1000 ( .A(G146), .B(n1049), .Z(n1193) );
XOR2_X1 U1001 ( .A(G125), .B(G140), .Z(n1049) );
XOR2_X1 U1002 ( .A(n1265), .B(n1266), .Z(n1264) );
NOR2_X1 U1003 ( .A1(G143), .A2(KEYINPUT14), .ZN(n1266) );
NAND3_X1 U1004 ( .A1(n1267), .A2(n1013), .A3(G214), .ZN(n1265) );
XOR2_X1 U1005 ( .A(KEYINPUT52), .B(G237), .Z(n1267) );
XOR2_X1 U1006 ( .A(G902), .B(KEYINPUT6), .Z(n1257) );
XOR2_X1 U1007 ( .A(n1094), .B(KEYINPUT9), .Z(n1255) );
INV_X1 U1008 ( .A(G475), .ZN(n1094) );
XOR2_X1 U1009 ( .A(n1027), .B(KEYINPUT59), .Z(n1153) );
XNOR2_X1 U1010 ( .A(n1268), .B(G478), .ZN(n1027) );
NAND2_X1 U1011 ( .A1(n1087), .A2(n1211), .ZN(n1268) );
INV_X1 U1012 ( .A(G902), .ZN(n1211) );
XOR2_X1 U1013 ( .A(n1269), .B(n1270), .Z(n1087) );
XNOR2_X1 U1014 ( .A(n1233), .B(n1271), .ZN(n1270) );
XOR2_X1 U1015 ( .A(n1272), .B(n1273), .Z(n1271) );
NOR2_X1 U1016 ( .A1(KEYINPUT25), .A2(G143), .ZN(n1273) );
NAND2_X1 U1017 ( .A1(n1194), .A2(G217), .ZN(n1272) );
AND2_X1 U1018 ( .A1(G234), .A2(n1013), .ZN(n1194) );
INV_X1 U1019 ( .A(G953), .ZN(n1013) );
XOR2_X1 U1020 ( .A(G134), .B(KEYINPUT13), .Z(n1233) );
XOR2_X1 U1021 ( .A(n1274), .B(n1275), .Z(n1269) );
NOR2_X1 U1022 ( .A1(KEYINPUT41), .A2(n1276), .ZN(n1275) );
XOR2_X1 U1023 ( .A(n975), .B(n1277), .Z(n1276) );
NAND2_X1 U1024 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
OR2_X1 U1025 ( .A1(n1175), .A2(G116), .ZN(n1279) );
XOR2_X1 U1026 ( .A(n1280), .B(KEYINPUT26), .Z(n1278) );
NAND2_X1 U1027 ( .A1(G116), .A2(n1175), .ZN(n1280) );
INV_X1 U1028 ( .A(G122), .ZN(n1175) );
INV_X1 U1029 ( .A(G107), .ZN(n975) );
XOR2_X1 U1030 ( .A(n1205), .B(KEYINPUT19), .Z(n1274) );
INV_X1 U1031 ( .A(G128), .ZN(n1205) );
INV_X1 U1032 ( .A(G110), .ZN(n1185) );
endmodule


