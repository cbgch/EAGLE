//Key = 0000101111100010011001011000011010000101101001010111000000010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
n1431, n1432;

XNOR2_X1 U787 ( .A(G107), .B(n1091), .ZN(G9) );
NAND2_X1 U788 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U789 ( .A(KEYINPUT54), .B(n1094), .ZN(n1093) );
NOR2_X1 U790 ( .A1(n1095), .A2(n1096), .ZN(G75) );
NOR4_X1 U791 ( .A1(n1097), .A2(n1098), .A3(G953), .A4(n1099), .ZN(n1096) );
NOR3_X1 U792 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1098) );
INV_X1 U793 ( .A(n1103), .ZN(n1102) );
NOR2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1101) );
NOR2_X1 U795 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
INV_X1 U796 ( .A(n1108), .ZN(n1107) );
NOR2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
NOR2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U799 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
AND2_X1 U800 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NOR3_X1 U801 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1109) );
NOR3_X1 U802 ( .A1(n1119), .A2(n1112), .A3(n1094), .ZN(n1104) );
INV_X1 U803 ( .A(n1120), .ZN(n1112) );
NAND3_X1 U804 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1097) );
NAND2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
NAND2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND3_X1 U807 ( .A1(n1108), .A2(n1128), .A3(n1129), .ZN(n1127) );
NAND2_X1 U808 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NAND2_X1 U809 ( .A1(n1120), .A2(n1132), .ZN(n1131) );
NAND2_X1 U810 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U811 ( .A1(n1103), .A2(n1135), .ZN(n1130) );
XOR2_X1 U812 ( .A(n1136), .B(KEYINPUT27), .Z(n1126) );
NAND4_X1 U813 ( .A1(n1129), .A2(n1137), .A3(n1103), .A4(n1120), .ZN(n1136) );
INV_X1 U814 ( .A(n1100), .ZN(n1129) );
NOR3_X1 U815 ( .A1(n1099), .A2(G953), .A3(G952), .ZN(n1095) );
AND3_X1 U816 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1099) );
NOR3_X1 U817 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1140) );
AND2_X1 U818 ( .A1(n1134), .A2(KEYINPUT36), .ZN(n1143) );
INV_X1 U819 ( .A(n1144), .ZN(n1134) );
NOR2_X1 U820 ( .A1(KEYINPUT36), .A2(n1103), .ZN(n1142) );
XNOR2_X1 U821 ( .A(n1145), .B(n1146), .ZN(n1141) );
XNOR2_X1 U822 ( .A(G478), .B(KEYINPUT34), .ZN(n1146) );
XOR2_X1 U823 ( .A(KEYINPUT28), .B(n1147), .Z(n1139) );
NOR3_X1 U824 ( .A1(n1148), .A2(n1116), .A3(n1149), .ZN(n1147) );
XOR2_X1 U825 ( .A(n1115), .B(KEYINPUT10), .Z(n1149) );
NAND3_X1 U826 ( .A1(n1150), .A2(n1151), .A3(n1117), .ZN(n1148) );
XOR2_X1 U827 ( .A(n1152), .B(n1153), .Z(G72) );
XOR2_X1 U828 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U829 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U830 ( .A(n1158), .B(n1159), .Z(n1157) );
XNOR2_X1 U831 ( .A(n1160), .B(n1161), .ZN(n1159) );
XNOR2_X1 U832 ( .A(KEYINPUT7), .B(n1162), .ZN(n1161) );
INV_X1 U833 ( .A(G131), .ZN(n1160) );
XOR2_X1 U834 ( .A(n1163), .B(n1164), .Z(n1158) );
XOR2_X1 U835 ( .A(n1165), .B(G125), .Z(n1163) );
NAND2_X1 U836 ( .A1(KEYINPUT8), .A2(n1166), .ZN(n1165) );
NOR2_X1 U837 ( .A1(G900), .A2(n1167), .ZN(n1156) );
NOR3_X1 U838 ( .A1(n1168), .A2(KEYINPUT33), .A3(n1169), .ZN(n1154) );
AND2_X1 U839 ( .A1(G227), .A2(G900), .ZN(n1169) );
INV_X1 U840 ( .A(n1170), .ZN(n1168) );
NOR3_X1 U841 ( .A1(n1123), .A2(KEYINPUT60), .A3(G953), .ZN(n1152) );
XOR2_X1 U842 ( .A(n1171), .B(n1172), .Z(G69) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U845 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
XNOR2_X1 U846 ( .A(n1175), .B(KEYINPUT5), .ZN(n1178) );
AND2_X1 U847 ( .A1(n1179), .A2(n1180), .ZN(n1175) );
XOR2_X1 U848 ( .A(n1181), .B(n1182), .Z(n1179) );
NOR2_X1 U849 ( .A1(KEYINPUT11), .A2(n1183), .ZN(n1182) );
XOR2_X1 U850 ( .A(n1184), .B(n1185), .Z(n1183) );
XNOR2_X1 U851 ( .A(n1186), .B(KEYINPUT53), .ZN(n1184) );
XOR2_X1 U852 ( .A(n1176), .B(KEYINPUT50), .Z(n1177) );
NAND3_X1 U853 ( .A1(n1187), .A2(n1188), .A3(n1167), .ZN(n1176) );
OR2_X1 U854 ( .A1(n1189), .A2(KEYINPUT23), .ZN(n1188) );
NAND2_X1 U855 ( .A1(KEYINPUT23), .A2(n1121), .ZN(n1187) );
NAND2_X1 U856 ( .A1(n1170), .A2(n1190), .ZN(n1171) );
NAND2_X1 U857 ( .A1(G898), .A2(G224), .ZN(n1190) );
XOR2_X1 U858 ( .A(G953), .B(KEYINPUT35), .Z(n1170) );
NOR2_X1 U859 ( .A1(n1191), .A2(n1192), .ZN(G66) );
XOR2_X1 U860 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U861 ( .A1(KEYINPUT46), .A2(n1195), .ZN(n1194) );
OR2_X1 U862 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
NOR2_X1 U863 ( .A1(n1191), .A2(n1198), .ZN(G63) );
NOR3_X1 U864 ( .A1(n1145), .A2(n1199), .A3(n1200), .ZN(n1198) );
NOR3_X1 U865 ( .A1(n1201), .A2(n1202), .A3(n1196), .ZN(n1200) );
NOR2_X1 U866 ( .A1(n1203), .A2(n1204), .ZN(n1199) );
NOR2_X1 U867 ( .A1(n1205), .A2(n1202), .ZN(n1204) );
AND2_X1 U868 ( .A1(n1206), .A2(n1123), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1191), .A2(n1207), .ZN(G60) );
XOR2_X1 U870 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U871 ( .A1(n1210), .A2(n1196), .ZN(n1209) );
INV_X1 U872 ( .A(G475), .ZN(n1210) );
XOR2_X1 U873 ( .A(G104), .B(n1211), .Z(G6) );
NOR2_X1 U874 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NOR3_X1 U875 ( .A1(n1191), .A2(n1214), .A3(n1215), .ZN(G57) );
NOR2_X1 U876 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
INV_X1 U877 ( .A(n1218), .ZN(n1217) );
NOR2_X1 U878 ( .A1(n1219), .A2(n1220), .ZN(n1216) );
NOR3_X1 U879 ( .A1(n1221), .A2(KEYINPUT55), .A3(n1222), .ZN(n1220) );
AND2_X1 U880 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
INV_X1 U881 ( .A(KEYINPUT47), .ZN(n1221) );
NOR2_X1 U882 ( .A1(n1223), .A2(n1218), .ZN(n1214) );
XOR2_X1 U883 ( .A(n1224), .B(n1225), .Z(n1218) );
XNOR2_X1 U884 ( .A(n1226), .B(n1227), .ZN(n1224) );
NOR2_X1 U885 ( .A1(n1228), .A2(n1196), .ZN(n1227) );
NOR2_X1 U886 ( .A1(KEYINPUT55), .A2(n1222), .ZN(n1223) );
XNOR2_X1 U887 ( .A(n1229), .B(n1230), .ZN(n1222) );
NAND2_X1 U888 ( .A1(KEYINPUT29), .A2(n1231), .ZN(n1229) );
NOR2_X1 U889 ( .A1(n1232), .A2(n1233), .ZN(G54) );
XOR2_X1 U890 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U891 ( .A(n1236), .B(n1237), .Z(n1235) );
XNOR2_X1 U892 ( .A(n1238), .B(n1239), .ZN(n1236) );
NOR3_X1 U893 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
NOR2_X1 U894 ( .A1(G110), .A2(n1243), .ZN(n1242) );
NOR2_X1 U895 ( .A1(KEYINPUT22), .A2(n1244), .ZN(n1243) );
XNOR2_X1 U896 ( .A(KEYINPUT12), .B(n1162), .ZN(n1244) );
NOR3_X1 U897 ( .A1(n1245), .A2(KEYINPUT22), .A3(G140), .ZN(n1241) );
AND2_X1 U898 ( .A1(G140), .A2(KEYINPUT22), .ZN(n1240) );
XOR2_X1 U899 ( .A(n1246), .B(n1247), .Z(n1234) );
NOR2_X1 U900 ( .A1(n1248), .A2(n1196), .ZN(n1247) );
XOR2_X1 U901 ( .A(n1249), .B(KEYINPUT61), .Z(n1246) );
NOR2_X1 U902 ( .A1(n1250), .A2(n1251), .ZN(n1232) );
XNOR2_X1 U903 ( .A(KEYINPUT49), .B(n1167), .ZN(n1251) );
XOR2_X1 U904 ( .A(KEYINPUT56), .B(G952), .Z(n1250) );
NOR2_X1 U905 ( .A1(n1191), .A2(n1252), .ZN(G51) );
NOR2_X1 U906 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U907 ( .A(n1255), .B(n1256), .Z(n1254) );
NOR2_X1 U908 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NOR2_X1 U909 ( .A1(n1259), .A2(n1196), .ZN(n1255) );
NAND2_X1 U910 ( .A1(G902), .A2(n1260), .ZN(n1196) );
NAND2_X1 U911 ( .A1(n1123), .A2(n1206), .ZN(n1260) );
XOR2_X1 U912 ( .A(n1121), .B(KEYINPUT19), .Z(n1206) );
AND4_X1 U913 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1121) );
AND4_X1 U914 ( .A1(n1189), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1264) );
NAND2_X1 U915 ( .A1(n1092), .A2(n1268), .ZN(n1263) );
NAND2_X1 U916 ( .A1(n1213), .A2(n1094), .ZN(n1268) );
INV_X1 U917 ( .A(n1269), .ZN(n1094) );
INV_X1 U918 ( .A(n1137), .ZN(n1213) );
INV_X1 U919 ( .A(n1212), .ZN(n1092) );
NAND2_X1 U920 ( .A1(n1103), .A2(n1270), .ZN(n1212) );
AND4_X1 U921 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1123) );
NOR4_X1 U922 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1274) );
INV_X1 U923 ( .A(n1279), .ZN(n1277) );
NOR2_X1 U924 ( .A1(n1280), .A2(n1281), .ZN(n1273) );
INV_X1 U925 ( .A(n1282), .ZN(n1281) );
AND2_X1 U926 ( .A1(n1258), .A2(n1257), .ZN(n1253) );
XOR2_X1 U927 ( .A(n1283), .B(n1284), .Z(n1257) );
INV_X1 U928 ( .A(KEYINPUT39), .ZN(n1258) );
AND2_X1 U929 ( .A1(n1285), .A2(G953), .ZN(n1191) );
XNOR2_X1 U930 ( .A(KEYINPUT56), .B(G952), .ZN(n1285) );
XNOR2_X1 U931 ( .A(G146), .B(n1271), .ZN(G48) );
NAND3_X1 U932 ( .A1(n1137), .A2(n1114), .A3(n1286), .ZN(n1271) );
XNOR2_X1 U933 ( .A(G143), .B(n1272), .ZN(G45) );
NAND4_X1 U934 ( .A1(n1287), .A2(n1114), .A3(n1288), .A4(n1289), .ZN(n1272) );
XNOR2_X1 U935 ( .A(G140), .B(n1282), .ZN(G42) );
NAND3_X1 U936 ( .A1(n1290), .A2(n1135), .A3(n1124), .ZN(n1282) );
XOR2_X1 U937 ( .A(G137), .B(n1280), .Z(G39) );
AND3_X1 U938 ( .A1(n1124), .A2(n1286), .A3(n1108), .ZN(n1280) );
XOR2_X1 U939 ( .A(G134), .B(n1278), .Z(G36) );
AND3_X1 U940 ( .A1(n1287), .A2(n1269), .A3(n1124), .ZN(n1278) );
XNOR2_X1 U941 ( .A(G131), .B(n1279), .ZN(G33) );
NAND3_X1 U942 ( .A1(n1287), .A2(n1137), .A3(n1124), .ZN(n1279) );
INV_X1 U943 ( .A(n1119), .ZN(n1124) );
NAND2_X1 U944 ( .A1(n1115), .A2(n1291), .ZN(n1119) );
AND3_X1 U945 ( .A1(n1135), .A2(n1292), .A3(n1293), .ZN(n1287) );
XOR2_X1 U946 ( .A(G128), .B(n1276), .Z(G30) );
AND3_X1 U947 ( .A1(n1269), .A2(n1114), .A3(n1286), .ZN(n1276) );
AND4_X1 U948 ( .A1(n1135), .A2(n1294), .A3(n1292), .A4(n1295), .ZN(n1286) );
XNOR2_X1 U949 ( .A(G101), .B(n1261), .ZN(G3) );
NAND3_X1 U950 ( .A1(n1293), .A2(n1270), .A3(n1108), .ZN(n1261) );
XOR2_X1 U951 ( .A(G125), .B(n1275), .Z(G27) );
AND3_X1 U952 ( .A1(n1114), .A2(n1120), .A3(n1290), .ZN(n1275) );
AND3_X1 U953 ( .A1(n1144), .A2(n1292), .A3(n1137), .ZN(n1290) );
NAND2_X1 U954 ( .A1(n1100), .A2(n1296), .ZN(n1292) );
NAND4_X1 U955 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1298), .ZN(n1296) );
INV_X1 U956 ( .A(G900), .ZN(n1298) );
XNOR2_X1 U957 ( .A(G122), .B(n1262), .ZN(G24) );
NAND4_X1 U958 ( .A1(n1299), .A2(n1103), .A3(n1288), .A4(n1289), .ZN(n1262) );
NOR2_X1 U959 ( .A1(n1295), .A2(n1294), .ZN(n1103) );
XNOR2_X1 U960 ( .A(n1267), .B(n1300), .ZN(G21) );
NOR2_X1 U961 ( .A1(KEYINPUT2), .A2(n1301), .ZN(n1300) );
NAND4_X1 U962 ( .A1(n1299), .A2(n1108), .A3(n1294), .A4(n1295), .ZN(n1267) );
XNOR2_X1 U963 ( .A(G116), .B(n1266), .ZN(G18) );
NAND3_X1 U964 ( .A1(n1293), .A2(n1269), .A3(n1299), .ZN(n1266) );
NOR2_X1 U965 ( .A1(n1289), .A2(n1302), .ZN(n1269) );
INV_X1 U966 ( .A(n1288), .ZN(n1302) );
XNOR2_X1 U967 ( .A(G113), .B(n1189), .ZN(G15) );
NAND3_X1 U968 ( .A1(n1293), .A2(n1137), .A3(n1299), .ZN(n1189) );
AND3_X1 U969 ( .A1(n1120), .A2(n1303), .A3(n1114), .ZN(n1299) );
NOR2_X1 U970 ( .A1(n1288), .A2(n1138), .ZN(n1137) );
INV_X1 U971 ( .A(n1289), .ZN(n1138) );
INV_X1 U972 ( .A(n1133), .ZN(n1293) );
NAND2_X1 U973 ( .A1(n1304), .A2(n1294), .ZN(n1133) );
XNOR2_X1 U974 ( .A(G110), .B(n1265), .ZN(G12) );
NAND3_X1 U975 ( .A1(n1144), .A2(n1270), .A3(n1108), .ZN(n1265) );
NOR2_X1 U976 ( .A1(n1288), .A2(n1289), .ZN(n1108) );
XOR2_X1 U977 ( .A(G475), .B(n1305), .Z(n1289) );
NOR2_X1 U978 ( .A1(n1208), .A2(G902), .ZN(n1305) );
AND2_X1 U979 ( .A1(n1306), .A2(n1307), .ZN(n1208) );
NAND2_X1 U980 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XOR2_X1 U981 ( .A(n1310), .B(KEYINPUT3), .Z(n1306) );
OR2_X1 U982 ( .A1(n1309), .A2(n1308), .ZN(n1310) );
XOR2_X1 U983 ( .A(n1311), .B(n1312), .Z(n1308) );
XNOR2_X1 U984 ( .A(G113), .B(G122), .ZN(n1311) );
NAND3_X1 U985 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1309) );
NAND2_X1 U986 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
INV_X1 U987 ( .A(KEYINPUT30), .ZN(n1317) );
NAND3_X1 U988 ( .A1(KEYINPUT30), .A2(n1318), .A3(n1319), .ZN(n1314) );
OR2_X1 U989 ( .A1(n1319), .A2(n1318), .ZN(n1313) );
NOR2_X1 U990 ( .A1(KEYINPUT63), .A2(n1316), .ZN(n1318) );
XNOR2_X1 U991 ( .A(n1320), .B(n1321), .ZN(n1316) );
NOR2_X1 U992 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NOR2_X1 U993 ( .A1(G125), .A2(n1324), .ZN(n1323) );
XNOR2_X1 U994 ( .A(KEYINPUT48), .B(n1162), .ZN(n1324) );
NAND2_X1 U995 ( .A1(n1325), .A2(n1326), .ZN(n1319) );
NAND2_X1 U996 ( .A1(G131), .A2(n1327), .ZN(n1326) );
XOR2_X1 U997 ( .A(KEYINPUT32), .B(n1328), .Z(n1325) );
NOR2_X1 U998 ( .A1(G131), .A2(n1327), .ZN(n1328) );
XOR2_X1 U999 ( .A(n1329), .B(n1330), .Z(n1327) );
NAND2_X1 U1000 ( .A1(KEYINPUT37), .A2(n1331), .ZN(n1330) );
NAND3_X1 U1001 ( .A1(n1332), .A2(n1167), .A3(G214), .ZN(n1329) );
XOR2_X1 U1002 ( .A(n1145), .B(n1333), .Z(n1288) );
NOR2_X1 U1003 ( .A1(KEYINPUT0), .A2(n1202), .ZN(n1333) );
INV_X1 U1004 ( .A(G478), .ZN(n1202) );
NOR2_X1 U1005 ( .A1(n1203), .A2(G902), .ZN(n1145) );
INV_X1 U1006 ( .A(n1201), .ZN(n1203) );
NAND2_X1 U1007 ( .A1(n1334), .A2(n1335), .ZN(n1201) );
NAND2_X1 U1008 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1009 ( .A(n1338), .B(n1339), .Z(n1334) );
NOR2_X1 U1010 ( .A1(n1197), .A2(n1340), .ZN(n1339) );
OR2_X1 U1011 ( .A1(n1337), .A2(n1336), .ZN(n1338) );
XNOR2_X1 U1012 ( .A(n1341), .B(n1342), .ZN(n1336) );
XNOR2_X1 U1013 ( .A(G107), .B(n1343), .ZN(n1342) );
NAND2_X1 U1014 ( .A1(n1344), .A2(KEYINPUT24), .ZN(n1343) );
XNOR2_X1 U1015 ( .A(G134), .B(n1345), .ZN(n1344) );
XNOR2_X1 U1016 ( .A(G116), .B(G122), .ZN(n1341) );
INV_X1 U1017 ( .A(KEYINPUT42), .ZN(n1337) );
AND3_X1 U1018 ( .A1(n1135), .A2(n1303), .A3(n1114), .ZN(n1270) );
NOR2_X1 U1019 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
INV_X1 U1020 ( .A(n1291), .ZN(n1116) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1346), .ZN(n1291) );
XNOR2_X1 U1022 ( .A(n1347), .B(n1259), .ZN(n1115) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1346), .ZN(n1259) );
NAND2_X1 U1024 ( .A1(n1332), .A2(n1348), .ZN(n1346) );
NAND2_X1 U1025 ( .A1(n1349), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1026 ( .A(n1283), .B(n1350), .Z(n1349) );
NOR2_X1 U1027 ( .A1(KEYINPUT58), .A2(n1284), .ZN(n1350) );
NAND2_X1 U1028 ( .A1(G224), .A2(n1167), .ZN(n1284) );
XOR2_X1 U1029 ( .A(n1351), .B(n1352), .Z(n1283) );
XOR2_X1 U1030 ( .A(n1353), .B(n1185), .Z(n1352) );
XNOR2_X1 U1031 ( .A(n1354), .B(n1312), .ZN(n1185) );
XNOR2_X1 U1032 ( .A(n1355), .B(n1231), .ZN(n1354) );
NAND2_X1 U1033 ( .A1(KEYINPUT51), .A2(n1356), .ZN(n1355) );
XNOR2_X1 U1034 ( .A(n1357), .B(n1181), .ZN(n1351) );
NAND2_X1 U1035 ( .A1(n1358), .A2(n1359), .ZN(n1181) );
NAND2_X1 U1036 ( .A1(G110), .A2(n1360), .ZN(n1359) );
NAND2_X1 U1037 ( .A1(KEYINPUT4), .A2(n1361), .ZN(n1360) );
NAND2_X1 U1038 ( .A1(G122), .A2(n1362), .ZN(n1361) );
NAND2_X1 U1039 ( .A1(n1363), .A2(n1364), .ZN(n1358) );
INV_X1 U1040 ( .A(G122), .ZN(n1364) );
NAND2_X1 U1041 ( .A1(n1362), .A2(n1365), .ZN(n1363) );
NAND2_X1 U1042 ( .A1(KEYINPUT4), .A2(n1245), .ZN(n1365) );
INV_X1 U1043 ( .A(G110), .ZN(n1245) );
INV_X1 U1044 ( .A(KEYINPUT38), .ZN(n1362) );
XOR2_X1 U1045 ( .A(n1366), .B(G125), .Z(n1357) );
NAND2_X1 U1046 ( .A1(KEYINPUT17), .A2(n1186), .ZN(n1366) );
XOR2_X1 U1047 ( .A(n1226), .B(n1367), .Z(n1186) );
XOR2_X1 U1048 ( .A(KEYINPUT59), .B(KEYINPUT31), .Z(n1367) );
NAND2_X1 U1049 ( .A1(n1100), .A2(n1368), .ZN(n1303) );
NAND3_X1 U1050 ( .A1(G902), .A2(n1297), .A3(n1369), .ZN(n1368) );
INV_X1 U1051 ( .A(n1180), .ZN(n1369) );
NAND2_X1 U1052 ( .A1(n1370), .A2(G953), .ZN(n1180) );
XNOR2_X1 U1053 ( .A(G898), .B(KEYINPUT26), .ZN(n1370) );
NAND3_X1 U1054 ( .A1(n1297), .A2(n1167), .A3(n1371), .ZN(n1100) );
XNOR2_X1 U1055 ( .A(G952), .B(KEYINPUT6), .ZN(n1371) );
NAND2_X1 U1056 ( .A1(G237), .A2(G234), .ZN(n1297) );
NAND2_X1 U1057 ( .A1(n1372), .A2(n1373), .ZN(n1135) );
NAND3_X1 U1058 ( .A1(n1117), .A2(n1118), .A3(n1374), .ZN(n1373) );
INV_X1 U1059 ( .A(KEYINPUT25), .ZN(n1374) );
NAND2_X1 U1060 ( .A1(KEYINPUT25), .A2(n1120), .ZN(n1372) );
NOR2_X1 U1061 ( .A1(n1118), .A2(n1375), .ZN(n1120) );
INV_X1 U1062 ( .A(n1117), .ZN(n1375) );
NAND2_X1 U1063 ( .A1(G221), .A2(n1376), .ZN(n1117) );
NAND2_X1 U1064 ( .A1(G234), .A2(n1348), .ZN(n1376) );
NAND3_X1 U1065 ( .A1(n1377), .A2(n1378), .A3(n1151), .ZN(n1118) );
NAND2_X1 U1066 ( .A1(n1379), .A2(n1248), .ZN(n1151) );
NAND2_X1 U1067 ( .A1(KEYINPUT13), .A2(n1248), .ZN(n1378) );
OR2_X1 U1068 ( .A1(n1150), .A2(KEYINPUT13), .ZN(n1377) );
OR2_X1 U1069 ( .A1(n1248), .A2(n1379), .ZN(n1150) );
AND2_X1 U1070 ( .A1(n1380), .A2(n1348), .ZN(n1379) );
XNOR2_X1 U1071 ( .A(n1381), .B(n1382), .ZN(n1380) );
INV_X1 U1072 ( .A(n1238), .ZN(n1382) );
XOR2_X1 U1073 ( .A(n1164), .B(n1383), .Z(n1238) );
XOR2_X1 U1074 ( .A(G146), .B(n1345), .Z(n1164) );
XOR2_X1 U1075 ( .A(G128), .B(G143), .Z(n1345) );
XNOR2_X1 U1076 ( .A(n1384), .B(n1385), .ZN(n1381) );
NOR2_X1 U1077 ( .A1(KEYINPUT1), .A2(n1237), .ZN(n1385) );
XNOR2_X1 U1078 ( .A(n1386), .B(n1312), .ZN(n1237) );
XOR2_X1 U1079 ( .A(G104), .B(KEYINPUT44), .Z(n1312) );
XNOR2_X1 U1080 ( .A(n1387), .B(n1388), .ZN(n1386) );
NAND2_X1 U1081 ( .A1(KEYINPUT62), .A2(n1356), .ZN(n1388) );
INV_X1 U1082 ( .A(G107), .ZN(n1356) );
NAND2_X1 U1083 ( .A1(KEYINPUT40), .A2(n1231), .ZN(n1387) );
NOR2_X1 U1084 ( .A1(KEYINPUT15), .A2(n1389), .ZN(n1384) );
XOR2_X1 U1085 ( .A(n1249), .B(n1390), .Z(n1389) );
XNOR2_X1 U1086 ( .A(n1162), .B(G110), .ZN(n1390) );
NAND2_X1 U1087 ( .A1(G227), .A2(n1167), .ZN(n1249) );
INV_X1 U1088 ( .A(G469), .ZN(n1248) );
NOR2_X1 U1089 ( .A1(n1294), .A2(n1304), .ZN(n1144) );
INV_X1 U1090 ( .A(n1295), .ZN(n1304) );
NAND3_X1 U1091 ( .A1(n1391), .A2(n1392), .A3(n1393), .ZN(n1295) );
NAND2_X1 U1092 ( .A1(G902), .A2(G217), .ZN(n1393) );
OR3_X1 U1093 ( .A1(n1195), .A2(G902), .A3(n1394), .ZN(n1392) );
NAND2_X1 U1094 ( .A1(n1394), .A2(n1195), .ZN(n1391) );
XOR2_X1 U1095 ( .A(n1395), .B(n1396), .Z(n1195) );
XOR2_X1 U1096 ( .A(n1397), .B(n1398), .Z(n1396) );
XOR2_X1 U1097 ( .A(n1399), .B(n1400), .Z(n1398) );
NOR2_X1 U1098 ( .A1(G110), .A2(KEYINPUT43), .ZN(n1400) );
NAND2_X1 U1099 ( .A1(n1401), .A2(n1402), .ZN(n1399) );
NAND2_X1 U1100 ( .A1(n1403), .A2(n1162), .ZN(n1402) );
INV_X1 U1101 ( .A(G140), .ZN(n1162) );
NAND2_X1 U1102 ( .A1(G125), .A2(n1404), .ZN(n1403) );
NAND2_X1 U1103 ( .A1(n1322), .A2(n1404), .ZN(n1401) );
INV_X1 U1104 ( .A(KEYINPUT52), .ZN(n1404) );
AND2_X1 U1105 ( .A1(G140), .A2(G125), .ZN(n1322) );
NAND2_X1 U1106 ( .A1(KEYINPUT9), .A2(n1320), .ZN(n1397) );
XOR2_X1 U1107 ( .A(n1405), .B(n1406), .Z(n1395) );
NOR2_X1 U1108 ( .A1(n1407), .A2(n1408), .ZN(n1406) );
XOR2_X1 U1109 ( .A(n1409), .B(KEYINPUT14), .Z(n1408) );
NAND3_X1 U1110 ( .A1(n1410), .A2(n1411), .A3(G221), .ZN(n1409) );
NOR2_X1 U1111 ( .A1(n1412), .A2(n1411), .ZN(n1407) );
XOR2_X1 U1112 ( .A(G137), .B(KEYINPUT16), .Z(n1411) );
AND2_X1 U1113 ( .A1(n1410), .A2(G221), .ZN(n1412) );
INV_X1 U1114 ( .A(n1340), .ZN(n1410) );
NAND2_X1 U1115 ( .A1(G234), .A2(n1167), .ZN(n1340) );
XNOR2_X1 U1116 ( .A(G119), .B(G128), .ZN(n1405) );
NOR2_X1 U1117 ( .A1(n1197), .A2(G234), .ZN(n1394) );
INV_X1 U1118 ( .A(G217), .ZN(n1197) );
XOR2_X1 U1119 ( .A(n1413), .B(n1228), .Z(n1294) );
INV_X1 U1120 ( .A(G472), .ZN(n1228) );
NAND2_X1 U1121 ( .A1(n1414), .A2(n1348), .ZN(n1413) );
INV_X1 U1122 ( .A(G902), .ZN(n1348) );
XOR2_X1 U1123 ( .A(n1415), .B(n1416), .Z(n1414) );
XNOR2_X1 U1124 ( .A(n1417), .B(n1231), .ZN(n1416) );
INV_X1 U1125 ( .A(G101), .ZN(n1231) );
NAND2_X1 U1126 ( .A1(n1418), .A2(n1419), .ZN(n1417) );
NAND2_X1 U1127 ( .A1(n1225), .A2(n1420), .ZN(n1419) );
NAND2_X1 U1128 ( .A1(KEYINPUT45), .A2(n1421), .ZN(n1420) );
NAND2_X1 U1129 ( .A1(KEYINPUT18), .A2(n1422), .ZN(n1421) );
INV_X1 U1130 ( .A(n1226), .ZN(n1422) );
INV_X1 U1131 ( .A(n1423), .ZN(n1225) );
NAND2_X1 U1132 ( .A1(n1226), .A2(n1424), .ZN(n1418) );
NAND2_X1 U1133 ( .A1(KEYINPUT18), .A2(n1425), .ZN(n1424) );
NAND2_X1 U1134 ( .A1(KEYINPUT45), .A2(n1423), .ZN(n1425) );
XOR2_X1 U1135 ( .A(n1353), .B(n1383), .Z(n1423) );
XNOR2_X1 U1136 ( .A(n1426), .B(n1166), .ZN(n1383) );
XOR2_X1 U1137 ( .A(G134), .B(G137), .Z(n1166) );
XNOR2_X1 U1138 ( .A(G131), .B(KEYINPUT57), .ZN(n1426) );
XOR2_X1 U1139 ( .A(G128), .B(n1427), .Z(n1353) );
NOR2_X1 U1140 ( .A1(n1428), .A2(n1429), .ZN(n1427) );
XOR2_X1 U1141 ( .A(KEYINPUT20), .B(n1430), .Z(n1429) );
NOR2_X1 U1142 ( .A1(n1331), .A2(n1431), .ZN(n1430) );
XNOR2_X1 U1143 ( .A(KEYINPUT41), .B(n1320), .ZN(n1431) );
INV_X1 U1144 ( .A(G143), .ZN(n1331) );
NOR2_X1 U1145 ( .A1(G143), .A2(n1320), .ZN(n1428) );
INV_X1 U1146 ( .A(G146), .ZN(n1320) );
XOR2_X1 U1147 ( .A(G113), .B(n1432), .Z(n1226) );
XNOR2_X1 U1148 ( .A(n1301), .B(G116), .ZN(n1432) );
INV_X1 U1149 ( .A(G119), .ZN(n1301) );
NAND2_X1 U1150 ( .A1(KEYINPUT21), .A2(n1230), .ZN(n1415) );
NAND3_X1 U1151 ( .A1(n1332), .A2(n1167), .A3(G210), .ZN(n1230) );
INV_X1 U1152 ( .A(G953), .ZN(n1167) );
INV_X1 U1153 ( .A(G237), .ZN(n1332) );
endmodule


