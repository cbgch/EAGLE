//Key = 1111000111001010101100001110000011100000001011011000001010110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330;

XNOR2_X1 U734 ( .A(n1019), .B(n1020), .ZN(G9) );
NOR2_X1 U735 ( .A1(KEYINPUT50), .A2(n1021), .ZN(n1020) );
NOR2_X1 U736 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U737 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
NAND3_X1 U738 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1024) );
NAND2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND3_X1 U741 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NAND2_X1 U742 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NAND2_X1 U743 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U745 ( .A1(n1044), .A2(n1045), .ZN(n1038) );
NAND2_X1 U746 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U748 ( .A1(n1040), .A2(n1050), .A3(n1044), .ZN(n1033) );
NAND2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U750 ( .A1(n1035), .A2(n1053), .ZN(n1052) );
NAND2_X1 U751 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND4_X1 U752 ( .A1(n1056), .A2(KEYINPUT47), .A3(G221), .A4(n1057), .ZN(n1055) );
NAND2_X1 U753 ( .A1(n1037), .A2(n1058), .ZN(n1051) );
NAND3_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NAND2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
OR2_X1 U756 ( .A1(n1064), .A2(KEYINPUT47), .ZN(n1059) );
INV_X1 U757 ( .A(n1065), .ZN(n1031) );
NOR3_X1 U758 ( .A1(n1066), .A2(G953), .A3(n1067), .ZN(n1022) );
INV_X1 U759 ( .A(n1028), .ZN(n1067) );
NAND4_X1 U760 ( .A1(n1068), .A2(n1035), .A3(n1037), .A4(n1069), .ZN(n1028) );
NOR3_X1 U761 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
XOR2_X1 U762 ( .A(n1073), .B(KEYINPUT61), .Z(n1071) );
NAND2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U764 ( .A(n1026), .B(KEYINPUT25), .Z(n1066) );
INV_X1 U765 ( .A(G952), .ZN(n1026) );
XOR2_X1 U766 ( .A(n1076), .B(n1077), .Z(G72) );
XOR2_X1 U767 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U768 ( .A1(n1080), .A2(n1029), .ZN(n1079) );
AND2_X1 U769 ( .A1(G227), .A2(G900), .ZN(n1080) );
NAND3_X1 U770 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1078) );
NAND2_X1 U771 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U772 ( .A(KEYINPUT6), .B(G953), .Z(n1084) );
NAND2_X1 U773 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
XOR2_X1 U774 ( .A(n1088), .B(KEYINPUT41), .Z(n1087) );
XNOR2_X1 U775 ( .A(KEYINPUT5), .B(n1089), .ZN(n1086) );
NAND2_X1 U776 ( .A1(n1090), .A2(n1091), .ZN(n1081) );
XOR2_X1 U777 ( .A(KEYINPUT5), .B(n1089), .Z(n1091) );
XOR2_X1 U778 ( .A(n1088), .B(KEYINPUT56), .Z(n1090) );
XOR2_X1 U779 ( .A(n1092), .B(n1093), .Z(n1088) );
XOR2_X1 U780 ( .A(n1094), .B(G137), .Z(n1092) );
NAND2_X1 U781 ( .A1(n1029), .A2(n1025), .ZN(n1076) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(G69) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1029), .ZN(n1096) );
XOR2_X1 U784 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U785 ( .A1(n1100), .A2(G953), .ZN(n1095) );
NAND2_X1 U786 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1103), .ZN(n1102) );
NAND2_X1 U788 ( .A1(G224), .A2(n1104), .ZN(n1101) );
NAND2_X1 U789 ( .A1(G898), .A2(n1099), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1105), .A2(n1106), .ZN(n1099) );
NAND2_X1 U791 ( .A1(G953), .A2(n1107), .ZN(n1106) );
XNOR2_X1 U792 ( .A(n1108), .B(n1109), .ZN(n1105) );
XOR2_X1 U793 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U794 ( .A1(KEYINPUT48), .A2(n1112), .ZN(n1110) );
XOR2_X1 U795 ( .A(KEYINPUT26), .B(n1113), .Z(n1112) );
NOR2_X1 U796 ( .A1(n1114), .A2(n1115), .ZN(G66) );
XNOR2_X1 U797 ( .A(n1116), .B(n1117), .ZN(n1115) );
NOR2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U799 ( .A1(n1114), .A2(n1120), .ZN(G63) );
XOR2_X1 U800 ( .A(n1121), .B(n1122), .Z(n1120) );
AND2_X1 U801 ( .A1(G478), .A2(n1123), .ZN(n1121) );
NOR2_X1 U802 ( .A1(n1114), .A2(n1124), .ZN(G60) );
XOR2_X1 U803 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U804 ( .A1(KEYINPUT60), .A2(n1127), .ZN(n1126) );
NAND2_X1 U805 ( .A1(n1123), .A2(G475), .ZN(n1125) );
XNOR2_X1 U806 ( .A(G104), .B(n1128), .ZN(G6) );
NAND2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U808 ( .A1(n1114), .A2(n1131), .ZN(G57) );
XOR2_X1 U809 ( .A(n1132), .B(n1133), .Z(n1131) );
XOR2_X1 U810 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U812 ( .A(n1138), .B(KEYINPUT44), .Z(n1137) );
NAND2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
XOR2_X1 U815 ( .A(n1141), .B(KEYINPUT21), .Z(n1140) );
NAND2_X1 U816 ( .A1(KEYINPUT34), .A2(n1142), .ZN(n1134) );
XOR2_X1 U817 ( .A(n1143), .B(n1144), .Z(n1132) );
AND2_X1 U818 ( .A1(G472), .A2(n1123), .ZN(n1144) );
INV_X1 U819 ( .A(n1119), .ZN(n1123) );
NAND2_X1 U820 ( .A1(KEYINPUT14), .A2(n1145), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1114), .A2(n1146), .ZN(G54) );
XOR2_X1 U822 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U823 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR3_X1 U824 ( .A1(n1119), .A2(KEYINPUT22), .A3(n1151), .ZN(n1149) );
XOR2_X1 U825 ( .A(n1152), .B(n1153), .Z(n1147) );
NOR3_X1 U826 ( .A1(n1154), .A2(KEYINPUT10), .A3(n1155), .ZN(n1153) );
AND2_X1 U827 ( .A1(n1156), .A2(G140), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1114), .A2(n1157), .ZN(G51) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U830 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U831 ( .A1(KEYINPUT16), .A2(n1162), .ZN(n1160) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1158) );
NOR2_X1 U833 ( .A1(n1165), .A2(n1119), .ZN(n1164) );
NAND2_X1 U834 ( .A1(G902), .A2(n1166), .ZN(n1119) );
NAND2_X1 U835 ( .A1(n1167), .A2(n1098), .ZN(n1166) );
INV_X1 U836 ( .A(n1027), .ZN(n1098) );
NAND4_X1 U837 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1027) );
AND4_X1 U838 ( .A1(n1019), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1171) );
NAND2_X1 U839 ( .A1(n1175), .A2(n1130), .ZN(n1019) );
AND2_X1 U840 ( .A1(n1176), .A2(n1040), .ZN(n1130) );
NAND2_X1 U841 ( .A1(n1177), .A2(n1178), .ZN(n1170) );
NAND2_X1 U842 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XNOR2_X1 U843 ( .A(KEYINPUT24), .B(n1181), .ZN(n1180) );
XOR2_X1 U844 ( .A(n1182), .B(KEYINPUT38), .Z(n1179) );
NAND4_X1 U845 ( .A1(n1129), .A2(n1040), .A3(n1183), .A4(n1184), .ZN(n1168) );
NAND2_X1 U846 ( .A1(KEYINPUT7), .A2(n1185), .ZN(n1184) );
NAND2_X1 U847 ( .A1(n1186), .A2(n1187), .ZN(n1183) );
INV_X1 U848 ( .A(KEYINPUT7), .ZN(n1187) );
NAND3_X1 U849 ( .A1(n1054), .A2(n1188), .A3(n1189), .ZN(n1186) );
XOR2_X1 U850 ( .A(n1025), .B(KEYINPUT54), .Z(n1167) );
NAND4_X1 U851 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1025) );
NOR4_X1 U852 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NOR2_X1 U853 ( .A1(n1198), .A2(n1042), .ZN(n1197) );
NOR2_X1 U854 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
AND3_X1 U855 ( .A1(n1043), .A2(n1200), .A3(KEYINPUT28), .ZN(n1195) );
INV_X1 U856 ( .A(n1201), .ZN(n1200) );
NOR2_X1 U857 ( .A1(n1202), .A2(n1043), .ZN(n1194) );
NOR3_X1 U858 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
AND3_X1 U859 ( .A1(KEYINPUT13), .A2(n1064), .A3(n1206), .ZN(n1205) );
NOR2_X1 U860 ( .A1(KEYINPUT13), .A2(n1207), .ZN(n1204) );
NOR2_X1 U861 ( .A1(KEYINPUT28), .A2(n1201), .ZN(n1203) );
NOR2_X1 U862 ( .A1(n1029), .A2(G952), .ZN(n1114) );
XOR2_X1 U863 ( .A(G146), .B(n1208), .Z(G48) );
NOR3_X1 U864 ( .A1(n1201), .A2(KEYINPUT53), .A3(n1042), .ZN(n1208) );
XOR2_X1 U865 ( .A(G143), .B(n1196), .Z(G45) );
AND2_X1 U866 ( .A1(n1209), .A2(n1206), .ZN(n1196) );
XNOR2_X1 U867 ( .A(G140), .B(n1192), .ZN(G42) );
NAND4_X1 U868 ( .A1(n1210), .A2(n1129), .A3(n1048), .A4(n1035), .ZN(n1192) );
XOR2_X1 U869 ( .A(n1211), .B(n1190), .Z(G39) );
NAND4_X1 U870 ( .A1(n1044), .A2(n1210), .A3(n1035), .A4(n1070), .ZN(n1190) );
NAND2_X1 U871 ( .A1(n1212), .A2(n1213), .ZN(G36) );
NAND4_X1 U872 ( .A1(n1199), .A2(n1175), .A3(n1214), .A4(n1215), .ZN(n1213) );
NAND2_X1 U873 ( .A1(G134), .A2(n1216), .ZN(n1215) );
NAND2_X1 U874 ( .A1(KEYINPUT51), .A2(n1217), .ZN(n1214) );
INV_X1 U875 ( .A(G134), .ZN(n1217) );
NAND3_X1 U876 ( .A1(n1218), .A2(n1216), .A3(G134), .ZN(n1212) );
INV_X1 U877 ( .A(KEYINPUT46), .ZN(n1216) );
OR3_X1 U878 ( .A1(n1043), .A2(KEYINPUT51), .A3(n1207), .ZN(n1218) );
XOR2_X1 U879 ( .A(n1219), .B(n1220), .Z(G33) );
XNOR2_X1 U880 ( .A(G131), .B(KEYINPUT30), .ZN(n1220) );
NAND2_X1 U881 ( .A1(n1199), .A2(n1129), .ZN(n1219) );
INV_X1 U882 ( .A(n1207), .ZN(n1199) );
NAND2_X1 U883 ( .A1(n1206), .A2(n1035), .ZN(n1207) );
INV_X1 U884 ( .A(n1064), .ZN(n1035) );
NAND2_X1 U885 ( .A1(n1063), .A2(n1221), .ZN(n1064) );
NOR3_X1 U886 ( .A1(n1054), .A2(n1222), .A3(n1046), .ZN(n1206) );
XOR2_X1 U887 ( .A(G128), .B(n1223), .Z(G30) );
NOR2_X1 U888 ( .A1(n1043), .A2(n1201), .ZN(n1223) );
NAND3_X1 U889 ( .A1(n1177), .A2(n1070), .A3(n1210), .ZN(n1201) );
NOR3_X1 U890 ( .A1(n1224), .A2(n1222), .A3(n1054), .ZN(n1210) );
XNOR2_X1 U891 ( .A(G101), .B(n1169), .ZN(G3) );
NAND3_X1 U892 ( .A1(n1044), .A2(n1176), .A3(n1225), .ZN(n1169) );
XNOR2_X1 U893 ( .A(G125), .B(n1191), .ZN(G27) );
NAND4_X1 U894 ( .A1(n1048), .A2(n1037), .A3(n1129), .A4(n1226), .ZN(n1191) );
NOR3_X1 U895 ( .A1(n1060), .A2(n1222), .A3(n1224), .ZN(n1226) );
AND2_X1 U896 ( .A1(n1227), .A2(n1228), .ZN(n1222) );
NAND4_X1 U897 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1085), .ZN(n1228) );
INV_X1 U898 ( .A(G900), .ZN(n1085) );
XOR2_X1 U899 ( .A(n1065), .B(KEYINPUT35), .Z(n1227) );
XOR2_X1 U900 ( .A(n1230), .B(n1174), .Z(G24) );
NAND3_X1 U901 ( .A1(n1209), .A2(n1040), .A3(n1231), .ZN(n1174) );
NOR2_X1 U902 ( .A1(n1070), .A2(n1049), .ZN(n1040) );
AND3_X1 U903 ( .A1(n1232), .A2(n1233), .A3(n1177), .ZN(n1209) );
XOR2_X1 U904 ( .A(G119), .B(n1234), .Z(G21) );
NOR2_X1 U905 ( .A1(n1060), .A2(n1181), .ZN(n1234) );
NAND4_X1 U906 ( .A1(n1231), .A2(n1044), .A3(n1049), .A4(n1070), .ZN(n1181) );
XOR2_X1 U907 ( .A(G116), .B(n1235), .Z(G18) );
NOR2_X1 U908 ( .A1(n1060), .A2(n1182), .ZN(n1235) );
NAND3_X1 U909 ( .A1(n1225), .A2(n1175), .A3(n1231), .ZN(n1182) );
INV_X1 U910 ( .A(n1043), .ZN(n1175) );
NAND2_X1 U911 ( .A1(n1236), .A2(n1232), .ZN(n1043) );
XOR2_X1 U912 ( .A(n1233), .B(KEYINPUT58), .Z(n1236) );
INV_X1 U913 ( .A(n1177), .ZN(n1060) );
XNOR2_X1 U914 ( .A(G113), .B(n1173), .ZN(G15) );
NAND4_X1 U915 ( .A1(n1231), .A2(n1225), .A3(n1129), .A4(n1189), .ZN(n1173) );
INV_X1 U916 ( .A(n1042), .ZN(n1129) );
NAND2_X1 U917 ( .A1(n1068), .A2(n1233), .ZN(n1042) );
INV_X1 U918 ( .A(n1046), .ZN(n1225) );
NAND2_X1 U919 ( .A1(n1224), .A2(n1070), .ZN(n1046) );
INV_X1 U920 ( .A(n1048), .ZN(n1070) );
AND2_X1 U921 ( .A1(n1037), .A2(n1188), .ZN(n1231) );
AND2_X1 U922 ( .A1(n1056), .A2(n1237), .ZN(n1037) );
XOR2_X1 U923 ( .A(G110), .B(n1238), .Z(G12) );
NOR2_X1 U924 ( .A1(KEYINPUT63), .A2(n1172), .ZN(n1238) );
NAND4_X1 U925 ( .A1(n1044), .A2(n1176), .A3(n1048), .A4(n1049), .ZN(n1172) );
INV_X1 U926 ( .A(n1224), .ZN(n1049) );
XNOR2_X1 U927 ( .A(n1072), .B(KEYINPUT11), .ZN(n1224) );
XOR2_X1 U928 ( .A(n1239), .B(n1118), .Z(n1072) );
NAND2_X1 U929 ( .A1(G217), .A2(n1057), .ZN(n1118) );
NAND2_X1 U930 ( .A1(n1116), .A2(n1240), .ZN(n1239) );
XNOR2_X1 U931 ( .A(n1241), .B(n1089), .ZN(n1116) );
XOR2_X1 U932 ( .A(n1242), .B(n1243), .Z(n1241) );
XOR2_X1 U933 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U934 ( .A(G137), .B(G128), .Z(n1245) );
XOR2_X1 U935 ( .A(KEYINPUT33), .B(KEYINPUT0), .Z(n1244) );
XOR2_X1 U936 ( .A(n1246), .B(n1247), .Z(n1242) );
XOR2_X1 U937 ( .A(n1248), .B(n1249), .Z(n1247) );
NOR2_X1 U938 ( .A1(KEYINPUT39), .A2(n1250), .ZN(n1248) );
XOR2_X1 U939 ( .A(n1156), .B(n1251), .Z(n1246) );
AND2_X1 U940 ( .A1(n1252), .A2(G221), .ZN(n1251) );
XOR2_X1 U941 ( .A(n1253), .B(G472), .Z(n1048) );
NAND2_X1 U942 ( .A1(n1254), .A2(n1240), .ZN(n1253) );
XOR2_X1 U943 ( .A(n1145), .B(n1255), .Z(n1254) );
XOR2_X1 U944 ( .A(KEYINPUT57), .B(n1256), .Z(n1255) );
NOR2_X1 U945 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U946 ( .A(n1259), .B(KEYINPUT9), .Z(n1258) );
NAND2_X1 U947 ( .A1(n1142), .A2(n1260), .ZN(n1259) );
NOR2_X1 U948 ( .A1(n1142), .A2(n1260), .ZN(n1257) );
XNOR2_X1 U949 ( .A(n1141), .B(n1139), .ZN(n1260) );
AND2_X1 U950 ( .A1(n1261), .A2(n1262), .ZN(n1142) );
NAND2_X1 U951 ( .A1(G116), .A2(n1263), .ZN(n1262) );
NAND2_X1 U952 ( .A1(n1264), .A2(n1265), .ZN(n1261) );
XNOR2_X1 U953 ( .A(KEYINPUT31), .B(n1263), .ZN(n1264) );
XNOR2_X1 U954 ( .A(n1266), .B(G101), .ZN(n1145) );
NAND2_X1 U955 ( .A1(G210), .A2(n1267), .ZN(n1266) );
INV_X1 U956 ( .A(n1185), .ZN(n1176) );
NAND3_X1 U957 ( .A1(n1189), .A2(n1188), .A3(n1268), .ZN(n1185) );
INV_X1 U958 ( .A(n1054), .ZN(n1268) );
NAND2_X1 U959 ( .A1(n1269), .A2(n1237), .ZN(n1054) );
NAND2_X1 U960 ( .A1(G221), .A2(n1057), .ZN(n1237) );
NAND2_X1 U961 ( .A1(n1270), .A2(n1240), .ZN(n1057) );
XNOR2_X1 U962 ( .A(G234), .B(KEYINPUT32), .ZN(n1270) );
XNOR2_X1 U963 ( .A(KEYINPUT20), .B(n1056), .ZN(n1269) );
XNOR2_X1 U964 ( .A(n1271), .B(n1151), .ZN(n1056) );
INV_X1 U965 ( .A(G469), .ZN(n1151) );
NAND2_X1 U966 ( .A1(n1272), .A2(n1240), .ZN(n1271) );
XOR2_X1 U967 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U968 ( .A(KEYINPUT45), .B(n1152), .ZN(n1274) );
NAND2_X1 U969 ( .A1(G227), .A2(n1029), .ZN(n1152) );
XNOR2_X1 U970 ( .A(n1150), .B(n1275), .ZN(n1273) );
NOR2_X1 U971 ( .A1(n1276), .A2(n1155), .ZN(n1275) );
NOR2_X1 U972 ( .A1(n1156), .A2(G140), .ZN(n1155) );
NOR2_X1 U973 ( .A1(G110), .A2(n1277), .ZN(n1276) );
XOR2_X1 U974 ( .A(KEYINPUT42), .B(G140), .Z(n1277) );
XNOR2_X1 U975 ( .A(n1278), .B(n1279), .ZN(n1150) );
XNOR2_X1 U976 ( .A(n1280), .B(n1281), .ZN(n1279) );
XOR2_X1 U977 ( .A(n1141), .B(n1093), .Z(n1278) );
XNOR2_X1 U978 ( .A(n1282), .B(n1283), .ZN(n1093) );
NOR2_X1 U979 ( .A1(G128), .A2(KEYINPUT29), .ZN(n1283) );
NAND2_X1 U980 ( .A1(n1284), .A2(n1285), .ZN(n1141) );
NAND2_X1 U981 ( .A1(n1286), .A2(n1211), .ZN(n1285) );
INV_X1 U982 ( .A(G137), .ZN(n1211) );
XOR2_X1 U983 ( .A(KEYINPUT1), .B(n1287), .Z(n1286) );
NAND2_X1 U984 ( .A1(n1287), .A2(G137), .ZN(n1284) );
INV_X1 U985 ( .A(n1094), .ZN(n1287) );
XNOR2_X1 U986 ( .A(G131), .B(n1288), .ZN(n1094) );
XOR2_X1 U987 ( .A(KEYINPUT62), .B(G134), .Z(n1288) );
NAND2_X1 U988 ( .A1(n1065), .A2(n1289), .ZN(n1188) );
NAND4_X1 U989 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1107), .ZN(n1289) );
INV_X1 U990 ( .A(G898), .ZN(n1107) );
NAND3_X1 U991 ( .A1(n1229), .A2(n1029), .A3(G952), .ZN(n1065) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n1229) );
XOR2_X1 U993 ( .A(n1177), .B(KEYINPUT17), .Z(n1189) );
NOR2_X1 U994 ( .A1(n1063), .A2(n1062), .ZN(n1177) );
INV_X1 U995 ( .A(n1221), .ZN(n1062) );
NAND2_X1 U996 ( .A1(G214), .A2(n1290), .ZN(n1221) );
XNOR2_X1 U997 ( .A(n1291), .B(n1165), .ZN(n1063) );
NAND2_X1 U998 ( .A1(G210), .A2(n1290), .ZN(n1165) );
NAND2_X1 U999 ( .A1(n1240), .A2(n1292), .ZN(n1290) );
INV_X1 U1000 ( .A(G237), .ZN(n1292) );
NAND2_X1 U1001 ( .A1(n1293), .A2(n1240), .ZN(n1291) );
INV_X1 U1002 ( .A(G902), .ZN(n1240) );
XOR2_X1 U1003 ( .A(n1161), .B(n1294), .Z(n1293) );
XOR2_X1 U1004 ( .A(n1163), .B(n1162), .Z(n1294) );
XNOR2_X1 U1005 ( .A(G125), .B(n1139), .ZN(n1162) );
XNOR2_X1 U1006 ( .A(n1295), .B(n1282), .ZN(n1139) );
XOR2_X1 U1007 ( .A(G143), .B(n1250), .Z(n1282) );
INV_X1 U1008 ( .A(G146), .ZN(n1250) );
XNOR2_X1 U1009 ( .A(G128), .B(KEYINPUT55), .ZN(n1295) );
NOR2_X1 U1010 ( .A1(n1103), .A2(G953), .ZN(n1163) );
INV_X1 U1011 ( .A(G224), .ZN(n1103) );
XOR2_X1 U1012 ( .A(n1296), .B(n1297), .Z(n1161) );
INV_X1 U1013 ( .A(n1111), .ZN(n1297) );
XOR2_X1 U1014 ( .A(n1156), .B(n1298), .Z(n1111) );
XOR2_X1 U1015 ( .A(KEYINPUT2), .B(G122), .Z(n1298) );
INV_X1 U1016 ( .A(G110), .ZN(n1156) );
NAND2_X1 U1017 ( .A1(n1299), .A2(n1300), .ZN(n1296) );
OR2_X1 U1018 ( .A1(n1113), .A2(n1108), .ZN(n1300) );
XOR2_X1 U1019 ( .A(n1301), .B(KEYINPUT15), .Z(n1299) );
NAND2_X1 U1020 ( .A1(n1108), .A2(n1113), .ZN(n1301) );
XNOR2_X1 U1021 ( .A(n1302), .B(n1280), .ZN(n1113) );
XOR2_X1 U1022 ( .A(G101), .B(G107), .Z(n1280) );
NAND2_X1 U1023 ( .A1(KEYINPUT3), .A2(n1281), .ZN(n1302) );
XNOR2_X1 U1024 ( .A(G104), .B(KEYINPUT23), .ZN(n1281) );
XNOR2_X1 U1025 ( .A(n1303), .B(n1304), .ZN(n1108) );
XOR2_X1 U1026 ( .A(KEYINPUT8), .B(KEYINPUT40), .Z(n1304) );
XOR2_X1 U1027 ( .A(n1263), .B(G116), .Z(n1303) );
XNOR2_X1 U1028 ( .A(G113), .B(n1249), .ZN(n1263) );
XOR2_X1 U1029 ( .A(G119), .B(KEYINPUT49), .Z(n1249) );
NOR2_X1 U1030 ( .A1(n1232), .A2(n1233), .ZN(n1044) );
NAND2_X1 U1031 ( .A1(n1305), .A2(n1075), .ZN(n1233) );
OR3_X1 U1032 ( .A1(G475), .A2(G902), .A3(n1127), .ZN(n1075) );
XOR2_X1 U1033 ( .A(n1074), .B(KEYINPUT37), .Z(n1305) );
NAND2_X1 U1034 ( .A1(G475), .A2(n1306), .ZN(n1074) );
OR2_X1 U1035 ( .A1(n1127), .A2(G902), .ZN(n1306) );
XOR2_X1 U1036 ( .A(n1307), .B(n1308), .Z(n1127) );
XOR2_X1 U1037 ( .A(G104), .B(n1309), .Z(n1308) );
XOR2_X1 U1038 ( .A(KEYINPUT36), .B(G146), .Z(n1309) );
XNOR2_X1 U1039 ( .A(n1089), .B(n1310), .ZN(n1307) );
XOR2_X1 U1040 ( .A(n1311), .B(n1312), .Z(n1310) );
NAND2_X1 U1041 ( .A1(n1313), .A2(KEYINPUT59), .ZN(n1312) );
XOR2_X1 U1042 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1043 ( .A(G143), .B(G131), .Z(n1315) );
NAND3_X1 U1044 ( .A1(G214), .A2(n1267), .A3(KEYINPUT19), .ZN(n1314) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1267) );
NAND2_X1 U1046 ( .A1(n1316), .A2(n1317), .ZN(n1311) );
OR2_X1 U1047 ( .A1(n1230), .A2(G113), .ZN(n1317) );
XOR2_X1 U1048 ( .A(n1318), .B(KEYINPUT52), .Z(n1316) );
NAND2_X1 U1049 ( .A1(G113), .A2(n1230), .ZN(n1318) );
INV_X1 U1050 ( .A(G122), .ZN(n1230) );
XOR2_X1 U1051 ( .A(G125), .B(G140), .Z(n1089) );
INV_X1 U1052 ( .A(n1068), .ZN(n1232) );
XOR2_X1 U1053 ( .A(n1319), .B(G478), .Z(n1068) );
OR2_X1 U1054 ( .A1(n1122), .A2(G902), .ZN(n1319) );
XNOR2_X1 U1055 ( .A(n1320), .B(n1321), .ZN(n1122) );
NOR2_X1 U1056 ( .A1(KEYINPUT43), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1057 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1058 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1059 ( .A(n1265), .B(G122), .Z(n1326) );
INV_X1 U1060 ( .A(G116), .ZN(n1265) );
NAND2_X1 U1061 ( .A1(n1327), .A2(KEYINPUT18), .ZN(n1325) );
XOR2_X1 U1062 ( .A(n1021), .B(KEYINPUT12), .Z(n1327) );
INV_X1 U1063 ( .A(G107), .ZN(n1021) );
XOR2_X1 U1064 ( .A(n1328), .B(n1329), .Z(n1323) );
XOR2_X1 U1065 ( .A(G134), .B(G128), .Z(n1329) );
XOR2_X1 U1066 ( .A(KEYINPUT27), .B(G143), .Z(n1328) );
NAND2_X1 U1067 ( .A1(G217), .A2(n1252), .ZN(n1320) );
AND2_X1 U1068 ( .A1(n1330), .A2(n1029), .ZN(n1252) );
INV_X1 U1069 ( .A(G953), .ZN(n1029) );
XOR2_X1 U1070 ( .A(KEYINPUT4), .B(G234), .Z(n1330) );
endmodule


