//Key = 0110100011011100110011101111100010010101010101110000001010110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391;

XNOR2_X1 U771 ( .A(G107), .B(n1066), .ZN(G9) );
NAND3_X1 U772 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
XOR2_X1 U773 ( .A(n1070), .B(KEYINPUT47), .Z(n1069) );
INV_X1 U774 ( .A(n1071), .ZN(n1068) );
NOR2_X1 U775 ( .A1(n1072), .A2(n1073), .ZN(G75) );
NOR4_X1 U776 ( .A1(G953), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1073) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR2_X1 U778 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR3_X1 U779 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
AND2_X1 U781 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR3_X1 U782 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1084) );
NOR3_X1 U783 ( .A1(n1091), .A2(n1092), .A3(n1067), .ZN(n1090) );
NOR2_X1 U784 ( .A1(n1087), .A2(n1093), .ZN(n1089) );
NOR4_X1 U785 ( .A1(n1094), .A2(n1088), .A3(n1095), .A4(n1091), .ZN(n1079) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NOR2_X1 U787 ( .A1(n1098), .A2(n1081), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1083), .ZN(n1096) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U792 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR3_X1 U793 ( .A1(n1074), .A2(G953), .A3(G952), .ZN(n1072) );
AND4_X1 U794 ( .A1(n1108), .A2(n1109), .A3(n1093), .A4(n1110), .ZN(n1074) );
NOR3_X1 U795 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1110) );
XOR2_X1 U796 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U797 ( .A(n1116), .B(KEYINPUT19), .Z(n1111) );
NAND4_X1 U798 ( .A1(n1117), .A2(n1118), .A3(n1102), .A4(n1107), .ZN(n1116) );
XNOR2_X1 U799 ( .A(n1119), .B(n1120), .ZN(n1118) );
NOR2_X1 U800 ( .A1(G469), .A2(KEYINPUT40), .ZN(n1120) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(n1117) );
XOR2_X1 U802 ( .A(KEYINPUT18), .B(n1123), .Z(n1122) );
XOR2_X1 U803 ( .A(KEYINPUT24), .B(n1124), .Z(n1109) );
XOR2_X1 U804 ( .A(n1125), .B(n1126), .Z(G72) );
NOR2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U806 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
NAND2_X1 U807 ( .A1(n1131), .A2(n1132), .ZN(n1125) );
NAND2_X1 U808 ( .A1(n1133), .A2(n1128), .ZN(n1132) );
XNOR2_X1 U809 ( .A(n1134), .B(n1135), .ZN(n1133) );
NAND3_X1 U810 ( .A1(n1134), .A2(n1136), .A3(G953), .ZN(n1131) );
XOR2_X1 U811 ( .A(KEYINPUT34), .B(G900), .Z(n1136) );
AND2_X1 U812 ( .A1(KEYINPUT9), .A2(n1137), .ZN(n1134) );
XOR2_X1 U813 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U814 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U815 ( .A1(KEYINPUT0), .A2(n1142), .ZN(n1141) );
XOR2_X1 U816 ( .A(G131), .B(n1143), .Z(n1138) );
XOR2_X1 U817 ( .A(G137), .B(G134), .Z(n1143) );
XOR2_X1 U818 ( .A(n1144), .B(n1145), .Z(G69) );
XOR2_X1 U819 ( .A(n1146), .B(n1147), .Z(n1145) );
OR2_X1 U820 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U821 ( .A1(n1128), .A2(n1150), .ZN(n1146) );
NOR3_X1 U822 ( .A1(n1128), .A2(KEYINPUT36), .A3(n1151), .ZN(n1144) );
AND2_X1 U823 ( .A1(G224), .A2(G898), .ZN(n1151) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(G66) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U826 ( .A1(n1156), .A2(n1157), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1152), .A2(n1158), .ZN(G63) );
XOR2_X1 U828 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U829 ( .A1(n1156), .A2(G478), .ZN(n1159) );
NOR2_X1 U830 ( .A1(n1152), .A2(n1161), .ZN(G60) );
XOR2_X1 U831 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U832 ( .A1(n1156), .A2(G475), .ZN(n1162) );
XNOR2_X1 U833 ( .A(n1164), .B(n1165), .ZN(G6) );
NAND2_X1 U834 ( .A1(KEYINPUT63), .A2(G104), .ZN(n1165) );
NOR2_X1 U835 ( .A1(n1152), .A2(n1166), .ZN(G57) );
XOR2_X1 U836 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U838 ( .A(n1171), .B(n1172), .Z(n1167) );
NOR2_X1 U839 ( .A1(KEYINPUT23), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U840 ( .A(n1174), .B(n1175), .ZN(n1173) );
NAND2_X1 U841 ( .A1(KEYINPUT41), .A2(n1176), .ZN(n1174) );
NAND2_X1 U842 ( .A1(n1156), .A2(G472), .ZN(n1171) );
NOR2_X1 U843 ( .A1(n1152), .A2(n1177), .ZN(G54) );
XOR2_X1 U844 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1179) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND2_X1 U847 ( .A1(n1156), .A2(G469), .ZN(n1180) );
XOR2_X1 U848 ( .A(n1184), .B(n1185), .Z(n1178) );
XOR2_X1 U849 ( .A(n1186), .B(n1187), .Z(n1184) );
NOR2_X1 U850 ( .A1(n1152), .A2(n1188), .ZN(G51) );
NOR2_X1 U851 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U852 ( .A(KEYINPUT57), .B(n1191), .Z(n1190) );
AND2_X1 U853 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U854 ( .A1(n1192), .A2(n1193), .ZN(n1189) );
NAND2_X1 U855 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U856 ( .A1(n1196), .A2(n1148), .ZN(n1195) );
XOR2_X1 U857 ( .A(KEYINPUT58), .B(n1197), .Z(n1194) );
NOR2_X1 U858 ( .A1(n1148), .A2(n1196), .ZN(n1197) );
XNOR2_X1 U859 ( .A(n1198), .B(G125), .ZN(n1196) );
NAND3_X1 U860 ( .A1(G210), .A2(n1199), .A3(n1156), .ZN(n1192) );
AND2_X1 U861 ( .A1(G902), .A2(n1076), .ZN(n1156) );
NAND2_X1 U862 ( .A1(n1135), .A2(n1200), .ZN(n1076) );
INV_X1 U863 ( .A(n1150), .ZN(n1200) );
NAND3_X1 U864 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1150) );
NOR3_X1 U865 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
INV_X1 U866 ( .A(n1207), .ZN(n1206) );
NOR3_X1 U867 ( .A1(n1071), .A2(n1208), .A3(n1209), .ZN(n1204) );
NOR2_X1 U868 ( .A1(n1105), .A2(n1210), .ZN(n1209) );
NOR2_X1 U869 ( .A1(KEYINPUT11), .A2(n1211), .ZN(n1210) );
NOR2_X1 U870 ( .A1(n1067), .A2(n1070), .ZN(n1208) );
NAND2_X1 U871 ( .A1(n1100), .A2(n1212), .ZN(n1202) );
NAND3_X1 U872 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1212) );
XNOR2_X1 U873 ( .A(KEYINPUT46), .B(n1216), .ZN(n1215) );
NAND3_X1 U874 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1214) );
NAND2_X1 U875 ( .A1(n1220), .A2(n1221), .ZN(n1217) );
NAND2_X1 U876 ( .A1(n1087), .A2(n1222), .ZN(n1221) );
NAND2_X1 U877 ( .A1(n1092), .A2(n1086), .ZN(n1220) );
XNOR2_X1 U878 ( .A(KEYINPUT4), .B(n1223), .ZN(n1213) );
NAND2_X1 U879 ( .A1(KEYINPUT11), .A2(n1164), .ZN(n1201) );
NOR3_X1 U880 ( .A1(n1071), .A2(n1070), .A3(n1211), .ZN(n1164) );
NAND2_X1 U881 ( .A1(n1100), .A2(n1224), .ZN(n1071) );
AND2_X1 U882 ( .A1(n1225), .A2(n1226), .ZN(n1135) );
AND4_X1 U883 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1226) );
AND4_X1 U884 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1225) );
OR3_X1 U885 ( .A1(n1083), .A2(n1235), .A3(n1236), .ZN(n1234) );
NOR2_X1 U886 ( .A1(n1128), .A2(G952), .ZN(n1152) );
XOR2_X1 U887 ( .A(n1237), .B(n1233), .Z(G48) );
NAND2_X1 U888 ( .A1(n1238), .A2(n1092), .ZN(n1233) );
XOR2_X1 U889 ( .A(n1239), .B(n1232), .Z(G45) );
OR4_X1 U890 ( .A1(n1236), .A2(n1240), .A3(n1108), .A4(n1241), .ZN(n1232) );
XOR2_X1 U891 ( .A(n1242), .B(n1231), .Z(G42) );
NAND4_X1 U892 ( .A1(n1243), .A2(n1092), .A3(n1244), .A4(n1245), .ZN(n1231) );
INV_X1 U893 ( .A(n1211), .ZN(n1092) );
XOR2_X1 U894 ( .A(n1246), .B(n1230), .Z(G39) );
NAND4_X1 U895 ( .A1(n1087), .A2(n1222), .A3(n1244), .A4(n1245), .ZN(n1230) );
INV_X1 U896 ( .A(n1083), .ZN(n1244) );
INV_X1 U897 ( .A(n1095), .ZN(n1087) );
XOR2_X1 U898 ( .A(G134), .B(n1247), .Z(G36) );
NOR3_X1 U899 ( .A1(n1236), .A2(n1248), .A3(n1235), .ZN(n1247) );
XOR2_X1 U900 ( .A(n1083), .B(KEYINPUT48), .Z(n1248) );
XNOR2_X1 U901 ( .A(n1249), .B(n1227), .ZN(G33) );
OR3_X1 U902 ( .A1(n1083), .A2(n1236), .A3(n1211), .ZN(n1227) );
NAND2_X1 U903 ( .A1(n1086), .A2(n1245), .ZN(n1236) );
NAND2_X1 U904 ( .A1(n1250), .A2(n1102), .ZN(n1083) );
XOR2_X1 U905 ( .A(n1251), .B(KEYINPUT27), .Z(n1249) );
XOR2_X1 U906 ( .A(n1252), .B(n1229), .Z(G30) );
NAND2_X1 U907 ( .A1(n1238), .A2(n1067), .ZN(n1229) );
INV_X1 U908 ( .A(n1235), .ZN(n1067) );
AND3_X1 U909 ( .A1(n1245), .A2(n1100), .A3(n1222), .ZN(n1238) );
AND2_X1 U910 ( .A1(n1105), .A2(n1253), .ZN(n1245) );
XOR2_X1 U911 ( .A(n1176), .B(n1207), .Z(G3) );
NAND4_X1 U912 ( .A1(n1254), .A2(n1086), .A3(n1105), .A4(n1100), .ZN(n1207) );
NAND2_X1 U913 ( .A1(n1255), .A2(n1256), .ZN(G27) );
NAND2_X1 U914 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XOR2_X1 U915 ( .A(n1259), .B(KEYINPUT33), .Z(n1255) );
OR2_X1 U916 ( .A1(n1258), .A2(n1257), .ZN(n1259) );
INV_X1 U917 ( .A(n1228), .ZN(n1257) );
NAND3_X1 U918 ( .A1(n1243), .A2(n1253), .A3(n1260), .ZN(n1228) );
NAND2_X1 U919 ( .A1(n1078), .A2(n1261), .ZN(n1253) );
NAND4_X1 U920 ( .A1(G953), .A2(G902), .A3(n1262), .A4(n1130), .ZN(n1261) );
INV_X1 U921 ( .A(G900), .ZN(n1130) );
XOR2_X1 U922 ( .A(G125), .B(KEYINPUT21), .Z(n1258) );
XOR2_X1 U923 ( .A(G122), .B(n1263), .Z(G24) );
NOR2_X1 U924 ( .A1(n1240), .A2(n1216), .ZN(n1263) );
NAND4_X1 U925 ( .A1(n1219), .A2(n1224), .A3(n1264), .A4(n1265), .ZN(n1216) );
NOR3_X1 U926 ( .A1(n1088), .A2(n1266), .A3(n1091), .ZN(n1224) );
XNOR2_X1 U927 ( .A(G119), .B(n1267), .ZN(G21) );
NAND3_X1 U928 ( .A1(KEYINPUT54), .A2(n1100), .A3(n1268), .ZN(n1267) );
XOR2_X1 U929 ( .A(n1269), .B(KEYINPUT56), .Z(n1268) );
NAND3_X1 U930 ( .A1(n1254), .A2(n1219), .A3(n1270), .ZN(n1269) );
XNOR2_X1 U931 ( .A(n1222), .B(KEYINPUT35), .ZN(n1270) );
AND2_X1 U932 ( .A1(n1271), .A2(n1091), .ZN(n1222) );
INV_X1 U933 ( .A(n1093), .ZN(n1091) );
XNOR2_X1 U934 ( .A(KEYINPUT43), .B(n1088), .ZN(n1271) );
INV_X1 U935 ( .A(n1240), .ZN(n1100) );
XOR2_X1 U936 ( .A(n1272), .B(n1205), .Z(G18) );
AND3_X1 U937 ( .A1(n1219), .A2(n1086), .A3(n1273), .ZN(n1205) );
NOR3_X1 U938 ( .A1(n1235), .A2(n1266), .A3(n1240), .ZN(n1273) );
NAND2_X1 U939 ( .A1(n1108), .A2(n1265), .ZN(n1235) );
INV_X1 U940 ( .A(n1241), .ZN(n1265) );
NAND2_X1 U941 ( .A1(KEYINPUT39), .A2(n1274), .ZN(n1272) );
XNOR2_X1 U942 ( .A(G113), .B(n1275), .ZN(G15) );
NAND3_X1 U943 ( .A1(n1260), .A2(n1086), .A3(n1276), .ZN(n1275) );
XOR2_X1 U944 ( .A(n1218), .B(KEYINPUT10), .Z(n1276) );
AND2_X1 U945 ( .A1(n1088), .A2(n1093), .ZN(n1086) );
NOR3_X1 U946 ( .A1(n1211), .A2(n1240), .A3(n1081), .ZN(n1260) );
INV_X1 U947 ( .A(n1219), .ZN(n1081) );
NOR2_X1 U948 ( .A1(n1106), .A2(n1277), .ZN(n1219) );
INV_X1 U949 ( .A(n1107), .ZN(n1277) );
NAND2_X1 U950 ( .A1(n1241), .A2(n1264), .ZN(n1211) );
INV_X1 U951 ( .A(n1108), .ZN(n1264) );
XOR2_X1 U952 ( .A(n1278), .B(n1279), .Z(G12) );
NOR2_X1 U953 ( .A1(KEYINPUT53), .A2(n1182), .ZN(n1279) );
NOR2_X1 U954 ( .A1(n1280), .A2(n1240), .ZN(n1278) );
NAND2_X1 U955 ( .A1(n1101), .A2(n1102), .ZN(n1240) );
NAND2_X1 U956 ( .A1(G214), .A2(n1199), .ZN(n1102) );
INV_X1 U957 ( .A(n1250), .ZN(n1101) );
XNOR2_X1 U958 ( .A(n1121), .B(n1281), .ZN(n1250) );
NOR2_X1 U959 ( .A1(n1123), .A2(KEYINPUT29), .ZN(n1281) );
AND2_X1 U960 ( .A1(n1282), .A2(n1199), .ZN(n1123) );
NAND2_X1 U961 ( .A1(n1283), .A2(n1284), .ZN(n1199) );
INV_X1 U962 ( .A(G237), .ZN(n1284) );
XOR2_X1 U963 ( .A(KEYINPUT7), .B(G210), .Z(n1282) );
NAND2_X1 U964 ( .A1(n1285), .A2(n1286), .ZN(n1121) );
XOR2_X1 U965 ( .A(n1198), .B(n1287), .Z(n1285) );
XNOR2_X1 U966 ( .A(n1148), .B(n1288), .ZN(n1287) );
NOR2_X1 U967 ( .A1(G125), .A2(KEYINPUT51), .ZN(n1288) );
XNOR2_X1 U968 ( .A(n1289), .B(n1290), .ZN(n1148) );
XOR2_X1 U969 ( .A(n1182), .B(n1291), .Z(n1290) );
NAND2_X1 U970 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U971 ( .A1(n1294), .A2(n1176), .ZN(n1293) );
NAND2_X1 U972 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U973 ( .A1(KEYINPUT44), .A2(KEYINPUT37), .ZN(n1296) );
NAND3_X1 U974 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1292) );
INV_X1 U975 ( .A(KEYINPUT44), .ZN(n1299) );
NAND2_X1 U976 ( .A1(KEYINPUT37), .A2(n1300), .ZN(n1298) );
NAND2_X1 U977 ( .A1(G101), .A2(n1295), .ZN(n1300) );
NAND2_X1 U978 ( .A1(n1295), .A2(n1301), .ZN(n1297) );
INV_X1 U979 ( .A(KEYINPUT37), .ZN(n1301) );
XOR2_X1 U980 ( .A(n1302), .B(n1303), .Z(n1289) );
NOR2_X1 U981 ( .A1(G122), .A2(KEYINPUT6), .ZN(n1303) );
XNOR2_X1 U982 ( .A(n1304), .B(n1305), .ZN(n1198) );
AND2_X1 U983 ( .A1(n1128), .A2(G224), .ZN(n1305) );
XOR2_X1 U984 ( .A(n1223), .B(KEYINPUT14), .Z(n1280) );
NAND3_X1 U985 ( .A1(n1243), .A2(n1105), .A3(n1254), .ZN(n1223) );
NOR2_X1 U986 ( .A1(n1095), .A2(n1266), .ZN(n1254) );
INV_X1 U987 ( .A(n1218), .ZN(n1266) );
NAND2_X1 U988 ( .A1(n1078), .A2(n1306), .ZN(n1218) );
NAND3_X1 U989 ( .A1(G902), .A2(n1262), .A3(n1149), .ZN(n1306) );
NOR2_X1 U990 ( .A1(n1128), .A2(G898), .ZN(n1149) );
NAND3_X1 U991 ( .A1(n1262), .A2(n1128), .A3(G952), .ZN(n1078) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n1262) );
NAND2_X1 U993 ( .A1(n1241), .A2(n1108), .ZN(n1095) );
XOR2_X1 U994 ( .A(n1307), .B(G475), .Z(n1108) );
NAND2_X1 U995 ( .A1(n1163), .A2(n1286), .ZN(n1307) );
XOR2_X1 U996 ( .A(n1308), .B(n1309), .Z(n1163) );
XOR2_X1 U997 ( .A(G113), .B(n1310), .Z(n1309) );
XOR2_X1 U998 ( .A(G146), .B(G122), .Z(n1310) );
XOR2_X1 U999 ( .A(n1311), .B(n1140), .Z(n1308) );
AND2_X1 U1000 ( .A1(n1312), .A2(n1313), .ZN(n1140) );
NAND2_X1 U1001 ( .A1(G125), .A2(n1242), .ZN(n1313) );
XOR2_X1 U1002 ( .A(n1314), .B(G104), .Z(n1311) );
NAND3_X1 U1003 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1314) );
OR2_X1 U1004 ( .A1(n1251), .A2(n1318), .ZN(n1317) );
NAND3_X1 U1005 ( .A1(n1318), .A2(n1251), .A3(KEYINPUT1), .ZN(n1316) );
INV_X1 U1006 ( .A(G131), .ZN(n1251) );
NOR2_X1 U1007 ( .A1(KEYINPUT42), .A2(n1319), .ZN(n1318) );
NAND2_X1 U1008 ( .A1(n1319), .A2(n1320), .ZN(n1315) );
INV_X1 U1009 ( .A(KEYINPUT1), .ZN(n1320) );
XOR2_X1 U1010 ( .A(n1321), .B(n1239), .Z(n1319) );
INV_X1 U1011 ( .A(G143), .ZN(n1239) );
NAND2_X1 U1012 ( .A1(G214), .A2(n1322), .ZN(n1321) );
NOR2_X1 U1013 ( .A1(n1112), .A2(n1124), .ZN(n1241) );
NOR2_X1 U1014 ( .A1(n1323), .A2(n1324), .ZN(n1124) );
AND2_X1 U1015 ( .A1(n1323), .A2(n1324), .ZN(n1112) );
XOR2_X1 U1016 ( .A(G478), .B(KEYINPUT50), .Z(n1324) );
NAND2_X1 U1017 ( .A1(n1160), .A2(n1286), .ZN(n1323) );
XOR2_X1 U1018 ( .A(n1325), .B(n1326), .Z(n1160) );
XOR2_X1 U1019 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1020 ( .A(G107), .B(n1329), .ZN(n1328) );
NOR2_X1 U1021 ( .A1(G116), .A2(KEYINPUT49), .ZN(n1329) );
NAND2_X1 U1022 ( .A1(G217), .A2(n1330), .ZN(n1327) );
XOR2_X1 U1023 ( .A(n1331), .B(n1332), .Z(n1325) );
XOR2_X1 U1024 ( .A(G143), .B(G134), .Z(n1332) );
XOR2_X1 U1025 ( .A(G122), .B(n1252), .Z(n1331) );
INV_X1 U1026 ( .A(G128), .ZN(n1252) );
INV_X1 U1027 ( .A(n1070), .ZN(n1105) );
NAND2_X1 U1028 ( .A1(n1106), .A2(n1107), .ZN(n1070) );
NAND2_X1 U1029 ( .A1(G221), .A2(n1333), .ZN(n1107) );
XNOR2_X1 U1030 ( .A(n1119), .B(G469), .ZN(n1106) );
NAND2_X1 U1031 ( .A1(n1334), .A2(n1286), .ZN(n1119) );
XOR2_X1 U1032 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U1033 ( .A(n1186), .B(n1337), .Z(n1336) );
NOR2_X1 U1034 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NOR3_X1 U1035 ( .A1(KEYINPUT38), .A2(n1340), .A3(n1341), .ZN(n1339) );
NOR2_X1 U1036 ( .A1(G110), .A2(n1342), .ZN(n1341) );
NOR2_X1 U1037 ( .A1(KEYINPUT30), .A2(n1185), .ZN(n1342) );
INV_X1 U1038 ( .A(n1343), .ZN(n1185) );
NOR2_X1 U1039 ( .A1(KEYINPUT30), .A2(n1182), .ZN(n1340) );
NOR2_X1 U1040 ( .A1(n1344), .A2(n1343), .ZN(n1338) );
XOR2_X1 U1041 ( .A(n1242), .B(KEYINPUT16), .Z(n1343) );
NOR2_X1 U1042 ( .A1(n1345), .A2(G110), .ZN(n1344) );
NOR2_X1 U1043 ( .A1(KEYINPUT30), .A2(n1346), .ZN(n1345) );
INV_X1 U1044 ( .A(KEYINPUT38), .ZN(n1346) );
XNOR2_X1 U1045 ( .A(n1142), .B(n1347), .ZN(n1186) );
XNOR2_X1 U1046 ( .A(n1348), .B(G128), .ZN(n1142) );
NAND2_X1 U1047 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1048 ( .A1(G143), .A2(n1237), .ZN(n1350) );
XOR2_X1 U1049 ( .A(KEYINPUT25), .B(n1351), .Z(n1349) );
NOR2_X1 U1050 ( .A1(G143), .A2(n1237), .ZN(n1351) );
XOR2_X1 U1051 ( .A(n1352), .B(n1353), .Z(n1335) );
NOR2_X1 U1052 ( .A1(KEYINPUT62), .A2(n1187), .ZN(n1353) );
XOR2_X1 U1053 ( .A(G101), .B(n1295), .Z(n1187) );
XOR2_X1 U1054 ( .A(G104), .B(G107), .Z(n1295) );
XNOR2_X1 U1055 ( .A(n1183), .B(KEYINPUT20), .ZN(n1352) );
NOR2_X1 U1056 ( .A1(n1129), .A2(G953), .ZN(n1183) );
INV_X1 U1057 ( .A(G227), .ZN(n1129) );
NOR2_X1 U1058 ( .A1(n1088), .A2(n1093), .ZN(n1243) );
XOR2_X1 U1059 ( .A(n1354), .B(n1157), .Z(n1093) );
AND2_X1 U1060 ( .A1(G217), .A2(n1333), .ZN(n1157) );
NAND2_X1 U1061 ( .A1(n1283), .A2(G234), .ZN(n1333) );
XNOR2_X1 U1062 ( .A(G902), .B(KEYINPUT55), .ZN(n1283) );
NAND2_X1 U1063 ( .A1(n1155), .A2(n1286), .ZN(n1354) );
XNOR2_X1 U1064 ( .A(n1355), .B(n1356), .ZN(n1155) );
XOR2_X1 U1065 ( .A(n1357), .B(n1358), .Z(n1356) );
NAND2_X1 U1066 ( .A1(G221), .A2(n1330), .ZN(n1358) );
AND2_X1 U1067 ( .A1(G234), .A2(n1128), .ZN(n1330) );
INV_X1 U1068 ( .A(G953), .ZN(n1128) );
NAND2_X1 U1069 ( .A1(n1359), .A2(n1360), .ZN(n1357) );
NAND2_X1 U1070 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
XOR2_X1 U1071 ( .A(KEYINPUT22), .B(n1363), .Z(n1359) );
NOR2_X1 U1072 ( .A1(n1362), .A2(n1361), .ZN(n1363) );
XOR2_X1 U1073 ( .A(KEYINPUT31), .B(n1237), .Z(n1361) );
AND2_X1 U1074 ( .A1(n1364), .A2(n1365), .ZN(n1362) );
NAND2_X1 U1075 ( .A1(n1366), .A2(n1242), .ZN(n1365) );
XNOR2_X1 U1076 ( .A(G125), .B(KEYINPUT12), .ZN(n1366) );
XOR2_X1 U1077 ( .A(n1312), .B(KEYINPUT3), .Z(n1364) );
OR2_X1 U1078 ( .A1(n1242), .A2(G125), .ZN(n1312) );
INV_X1 U1079 ( .A(G140), .ZN(n1242) );
XOR2_X1 U1080 ( .A(n1367), .B(n1368), .Z(n1355) );
NOR2_X1 U1081 ( .A1(KEYINPUT60), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1082 ( .A(n1182), .B(n1370), .Z(n1369) );
XOR2_X1 U1083 ( .A(G128), .B(G119), .Z(n1370) );
INV_X1 U1084 ( .A(G110), .ZN(n1182) );
XOR2_X1 U1085 ( .A(n1246), .B(KEYINPUT15), .Z(n1367) );
XNOR2_X1 U1086 ( .A(n1371), .B(n1114), .ZN(n1088) );
NAND2_X1 U1087 ( .A1(n1286), .A2(n1372), .ZN(n1114) );
NAND2_X1 U1088 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NAND3_X1 U1089 ( .A1(n1375), .A2(n1376), .A3(n1377), .ZN(n1374) );
XOR2_X1 U1090 ( .A(n1378), .B(n1379), .Z(n1375) );
XOR2_X1 U1091 ( .A(n1380), .B(KEYINPUT52), .Z(n1373) );
NAND2_X1 U1092 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
NAND2_X1 U1093 ( .A1(n1377), .A2(n1376), .ZN(n1382) );
NAND2_X1 U1094 ( .A1(n1175), .A2(n1176), .ZN(n1376) );
XNOR2_X1 U1095 ( .A(n1383), .B(KEYINPUT59), .ZN(n1377) );
OR2_X1 U1096 ( .A1(n1175), .A2(n1176), .ZN(n1383) );
INV_X1 U1097 ( .A(G101), .ZN(n1176) );
NAND2_X1 U1098 ( .A1(G210), .A2(n1322), .ZN(n1175) );
NOR2_X1 U1099 ( .A1(G953), .A2(G237), .ZN(n1322) );
XOR2_X1 U1100 ( .A(n1378), .B(n1169), .Z(n1381) );
INV_X1 U1101 ( .A(n1379), .ZN(n1169) );
XOR2_X1 U1102 ( .A(n1302), .B(KEYINPUT28), .Z(n1379) );
XOR2_X1 U1103 ( .A(n1384), .B(n1385), .Z(n1302) );
XOR2_X1 U1104 ( .A(KEYINPUT45), .B(G119), .Z(n1385) );
XOR2_X1 U1105 ( .A(G113), .B(n1274), .Z(n1384) );
INV_X1 U1106 ( .A(G116), .ZN(n1274) );
NAND2_X1 U1107 ( .A1(KEYINPUT61), .A2(n1170), .ZN(n1378) );
XNOR2_X1 U1108 ( .A(n1386), .B(n1304), .ZN(n1170) );
XNOR2_X1 U1109 ( .A(n1387), .B(n1388), .ZN(n1304) );
XOR2_X1 U1110 ( .A(G143), .B(G128), .Z(n1388) );
NAND2_X1 U1111 ( .A1(KEYINPUT32), .A2(n1237), .ZN(n1387) );
INV_X1 U1112 ( .A(G146), .ZN(n1237) );
XNOR2_X1 U1113 ( .A(n1347), .B(KEYINPUT5), .ZN(n1386) );
XNOR2_X1 U1114 ( .A(n1389), .B(G131), .ZN(n1347) );
NAND2_X1 U1115 ( .A1(KEYINPUT2), .A2(n1390), .ZN(n1389) );
XOR2_X1 U1116 ( .A(n1246), .B(n1391), .Z(n1390) );
NAND2_X1 U1117 ( .A1(KEYINPUT17), .A2(G134), .ZN(n1391) );
INV_X1 U1118 ( .A(G137), .ZN(n1246) );
XOR2_X1 U1119 ( .A(G902), .B(KEYINPUT8), .Z(n1286) );
NAND2_X1 U1120 ( .A1(KEYINPUT13), .A2(n1115), .ZN(n1371) );
XOR2_X1 U1121 ( .A(G472), .B(KEYINPUT26), .Z(n1115) );
endmodule


