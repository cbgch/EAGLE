//Key = 0100001010110010011001010100111111001111101101110111111011001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318;

XNOR2_X1 U718 ( .A(G107), .B(n995), .ZN(G9) );
NOR2_X1 U719 ( .A1(n996), .A2(n997), .ZN(G75) );
NOR3_X1 U720 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
NOR2_X1 U721 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U722 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U723 ( .A1(KEYINPUT60), .A2(n1005), .ZN(n1004) );
NOR4_X1 U724 ( .A1(n1006), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n1005) );
INV_X1 U725 ( .A(n1010), .ZN(n1006) );
NOR2_X1 U726 ( .A1(n1011), .A2(n1009), .ZN(n1003) );
NOR2_X1 U727 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U728 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
INV_X1 U729 ( .A(n1016), .ZN(n1015) );
NOR2_X1 U730 ( .A1(n1017), .A2(n1018), .ZN(n1014) );
NOR2_X1 U731 ( .A1(n1019), .A2(n1008), .ZN(n1018) );
NOR2_X1 U732 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
AND2_X1 U733 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U734 ( .A1(n1024), .A2(n1007), .ZN(n1017) );
NOR2_X1 U735 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR3_X1 U736 ( .A1(n1008), .A2(n1027), .A3(n1007), .ZN(n1012) );
INV_X1 U737 ( .A(n1028), .ZN(n1007) );
NOR2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
AND2_X1 U739 ( .A1(n1010), .A2(KEYINPUT60), .ZN(n1030) );
NOR2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NAND3_X1 U741 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n998) );
NAND4_X1 U742 ( .A1(n1028), .A2(n1036), .A3(n1016), .A4(n1037), .ZN(n1035) );
NOR2_X1 U743 ( .A1(n1008), .A2(n1009), .ZN(n1037) );
INV_X1 U744 ( .A(n1038), .ZN(n1008) );
NAND2_X1 U745 ( .A1(n1039), .A2(n1040), .ZN(n1036) );
NAND2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
INV_X1 U747 ( .A(n1043), .ZN(n1039) );
NOR3_X1 U748 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n996) );
INV_X1 U749 ( .A(n1033), .ZN(n1044) );
NAND4_X1 U750 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1033) );
NOR4_X1 U751 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
XOR2_X1 U752 ( .A(n1053), .B(n1054), .Z(n1052) );
XNOR2_X1 U753 ( .A(G472), .B(KEYINPUT3), .ZN(n1054) );
XNOR2_X1 U754 ( .A(G475), .B(n1055), .ZN(n1051) );
NAND2_X1 U755 ( .A1(KEYINPUT49), .A2(n1056), .ZN(n1055) );
XNOR2_X1 U756 ( .A(n1057), .B(n1058), .ZN(n1049) );
NAND2_X1 U757 ( .A1(KEYINPUT43), .A2(n1059), .ZN(n1057) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1041), .ZN(n1047) );
XNOR2_X1 U759 ( .A(n1061), .B(n1062), .ZN(n1046) );
NAND2_X1 U760 ( .A1(KEYINPUT31), .A2(n1063), .ZN(n1062) );
XOR2_X1 U761 ( .A(n1064), .B(n1065), .Z(n1045) );
NOR2_X1 U762 ( .A1(n1066), .A2(KEYINPUT55), .ZN(n1065) );
XOR2_X1 U763 ( .A(n1067), .B(n1068), .Z(G72) );
NOR2_X1 U764 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XNOR2_X1 U765 ( .A(G953), .B(KEYINPUT16), .ZN(n1070) );
AND2_X1 U766 ( .A1(G227), .A2(G900), .ZN(n1069) );
NAND2_X1 U767 ( .A1(n1071), .A2(n1072), .ZN(n1067) );
NAND2_X1 U768 ( .A1(n1073), .A2(n1034), .ZN(n1072) );
XOR2_X1 U769 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
XNOR2_X1 U771 ( .A(n1078), .B(KEYINPUT18), .ZN(n1076) );
NAND3_X1 U772 ( .A1(G900), .A2(n1075), .A3(G953), .ZN(n1071) );
XNOR2_X1 U773 ( .A(n1079), .B(n1080), .ZN(n1075) );
XNOR2_X1 U774 ( .A(n1081), .B(n1082), .ZN(n1080) );
NOR2_X1 U775 ( .A1(KEYINPUT48), .A2(n1083), .ZN(n1082) );
XOR2_X1 U776 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U777 ( .A(n1086), .B(G134), .ZN(n1085) );
INV_X1 U778 ( .A(G137), .ZN(n1086) );
XNOR2_X1 U779 ( .A(n1087), .B(n1088), .ZN(n1084) );
NAND2_X1 U780 ( .A1(KEYINPUT50), .A2(G140), .ZN(n1081) );
XNOR2_X1 U781 ( .A(G125), .B(KEYINPUT53), .ZN(n1079) );
XOR2_X1 U782 ( .A(n1089), .B(n1090), .Z(G69) );
XOR2_X1 U783 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U784 ( .A1(n1093), .A2(n1034), .ZN(n1092) );
AND2_X1 U785 ( .A1(G224), .A2(G898), .ZN(n1093) );
NAND2_X1 U786 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
NAND2_X1 U787 ( .A1(G953), .A2(n1096), .ZN(n1095) );
XOR2_X1 U788 ( .A(n1097), .B(n1098), .Z(n1094) );
XOR2_X1 U789 ( .A(KEYINPUT40), .B(G110), .Z(n1098) );
XOR2_X1 U790 ( .A(n1099), .B(n1100), .Z(n1097) );
NAND2_X1 U791 ( .A1(n1034), .A2(n1101), .ZN(n1089) );
NAND2_X1 U792 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(G66) );
NOR3_X1 U794 ( .A1(n1061), .A2(n1106), .A3(n1107), .ZN(n1105) );
NOR3_X1 U795 ( .A1(n1108), .A2(n1063), .A3(n1109), .ZN(n1107) );
NOR2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1106) );
NOR2_X1 U797 ( .A1(n1112), .A2(n1063), .ZN(n1110) );
NOR2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(G63) );
XOR2_X1 U799 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND3_X1 U800 ( .A1(n1117), .A2(G478), .A3(KEYINPUT57), .ZN(n1115) );
NOR2_X1 U801 ( .A1(n1118), .A2(n1034), .ZN(n1113) );
XNOR2_X1 U802 ( .A(G952), .B(KEYINPUT21), .ZN(n1118) );
NOR2_X1 U803 ( .A1(n1104), .A2(n1119), .ZN(G60) );
NOR3_X1 U804 ( .A1(n1056), .A2(n1120), .A3(n1121), .ZN(n1119) );
AND2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR3_X1 U806 ( .A1(n1123), .A2(n1124), .A3(n1122), .ZN(n1120) );
NAND2_X1 U807 ( .A1(G475), .A2(n1125), .ZN(n1122) );
XNOR2_X1 U808 ( .A(KEYINPUT14), .B(n1000), .ZN(n1125) );
XNOR2_X1 U809 ( .A(G104), .B(n1126), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1104), .A2(n1127), .ZN(G57) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U812 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U813 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U814 ( .A1(n1134), .A2(n1109), .ZN(n1133) );
AND2_X1 U815 ( .A1(n1135), .A2(KEYINPUT17), .ZN(n1132) );
NOR2_X1 U816 ( .A1(KEYINPUT17), .A2(n1135), .ZN(n1130) );
XNOR2_X1 U817 ( .A(n1136), .B(n1137), .ZN(n1135) );
NAND4_X1 U818 ( .A1(KEYINPUT62), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1136) );
NAND2_X1 U819 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U820 ( .A(KEYINPUT1), .ZN(n1142) );
NAND2_X1 U821 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
XNOR2_X1 U822 ( .A(KEYINPUT56), .B(n1145), .ZN(n1143) );
NAND2_X1 U823 ( .A1(KEYINPUT1), .A2(n1146), .ZN(n1139) );
NAND2_X1 U824 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
OR2_X1 U825 ( .A1(n1145), .A2(KEYINPUT56), .ZN(n1148) );
NAND3_X1 U826 ( .A1(n1144), .A2(n1145), .A3(KEYINPUT56), .ZN(n1147) );
NAND2_X1 U827 ( .A1(n1149), .A2(n1150), .ZN(n1138) );
NAND2_X1 U828 ( .A1(n1151), .A2(n1152), .ZN(n1128) );
NAND2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U830 ( .A(KEYINPUT33), .B(n1155), .Z(n1151) );
NOR2_X1 U831 ( .A1(n1153), .A2(n1154), .ZN(n1155) );
NOR2_X1 U832 ( .A1(n1156), .A2(n1157), .ZN(G54) );
XOR2_X1 U833 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U834 ( .A(KEYINPUT63), .B(n1160), .Z(n1159) );
NOR2_X1 U835 ( .A1(n1058), .A2(n1109), .ZN(n1160) );
NOR2_X1 U836 ( .A1(G952), .A2(n1161), .ZN(n1156) );
XNOR2_X1 U837 ( .A(KEYINPUT46), .B(n1034), .ZN(n1161) );
NOR2_X1 U838 ( .A1(n1104), .A2(n1162), .ZN(G51) );
XOR2_X1 U839 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U840 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U841 ( .A1(n1167), .A2(n1109), .ZN(n1166) );
INV_X1 U842 ( .A(n1117), .ZN(n1109) );
NOR2_X1 U843 ( .A1(n1124), .A2(n1112), .ZN(n1117) );
INV_X1 U844 ( .A(n1000), .ZN(n1112) );
NAND4_X1 U845 ( .A1(n1168), .A2(n1078), .A3(n1102), .A4(n1077), .ZN(n1000) );
AND4_X1 U846 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1077) );
NAND3_X1 U847 ( .A1(n1173), .A2(n1174), .A3(n1038), .ZN(n1169) );
AND4_X1 U848 ( .A1(n1175), .A2(n1176), .A3(n1126), .A4(n1177), .ZN(n1102) );
AND4_X1 U849 ( .A1(n995), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1177) );
NAND3_X1 U850 ( .A1(n1028), .A2(n1181), .A3(n1025), .ZN(n995) );
NAND3_X1 U851 ( .A1(n1028), .A2(n1181), .A3(n1026), .ZN(n1126) );
AND4_X1 U852 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1078) );
NAND3_X1 U853 ( .A1(n1186), .A2(n1025), .A3(n1173), .ZN(n1182) );
XOR2_X1 U854 ( .A(n1103), .B(KEYINPUT13), .Z(n1168) );
XNOR2_X1 U855 ( .A(n1187), .B(n1188), .ZN(n1163) );
NOR2_X1 U856 ( .A1(KEYINPUT24), .A2(n1189), .ZN(n1188) );
NOR2_X1 U857 ( .A1(n1034), .A2(G952), .ZN(n1104) );
XNOR2_X1 U858 ( .A(G146), .B(n1170), .ZN(G48) );
NAND3_X1 U859 ( .A1(n1026), .A2(n1043), .A3(n1174), .ZN(n1170) );
XNOR2_X1 U860 ( .A(n1171), .B(n1190), .ZN(G45) );
NOR2_X1 U861 ( .A1(KEYINPUT34), .A2(n1191), .ZN(n1190) );
INV_X1 U862 ( .A(G143), .ZN(n1191) );
NAND4_X1 U863 ( .A1(n1186), .A2(n1043), .A3(n1050), .A4(n1192), .ZN(n1171) );
XNOR2_X1 U864 ( .A(G140), .B(n1172), .ZN(G42) );
NAND3_X1 U865 ( .A1(n1193), .A2(n1010), .A3(n1173), .ZN(n1172) );
XNOR2_X1 U866 ( .A(G137), .B(n1194), .ZN(G39) );
NAND3_X1 U867 ( .A1(n1038), .A2(n1174), .A3(n1195), .ZN(n1194) );
XNOR2_X1 U868 ( .A(n1173), .B(KEYINPUT52), .ZN(n1195) );
XOR2_X1 U869 ( .A(G134), .B(n1196), .Z(G36) );
NOR4_X1 U870 ( .A1(KEYINPUT59), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1196) );
XNOR2_X1 U871 ( .A(KEYINPUT10), .B(n1002), .ZN(n1199) );
INV_X1 U872 ( .A(n1173), .ZN(n1002) );
INV_X1 U873 ( .A(n1025), .ZN(n1197) );
XOR2_X1 U874 ( .A(n1183), .B(n1200), .Z(G33) );
XNOR2_X1 U875 ( .A(G131), .B(KEYINPUT15), .ZN(n1200) );
NAND3_X1 U876 ( .A1(n1186), .A2(n1026), .A3(n1173), .ZN(n1183) );
NOR2_X1 U877 ( .A1(n1201), .A2(n1041), .ZN(n1173) );
INV_X1 U878 ( .A(n1198), .ZN(n1186) );
NAND3_X1 U879 ( .A1(n1010), .A2(n1202), .A3(n1021), .ZN(n1198) );
XNOR2_X1 U880 ( .A(G128), .B(n1184), .ZN(G30) );
NAND3_X1 U881 ( .A1(n1025), .A2(n1043), .A3(n1174), .ZN(n1184) );
AND4_X1 U882 ( .A1(n1203), .A2(n1010), .A3(n1022), .A4(n1202), .ZN(n1174) );
XNOR2_X1 U883 ( .A(G101), .B(n1175), .ZN(G3) );
NAND3_X1 U884 ( .A1(n1021), .A2(n1181), .A3(n1038), .ZN(n1175) );
XNOR2_X1 U885 ( .A(G125), .B(n1185), .ZN(G27) );
NAND3_X1 U886 ( .A1(n1193), .A2(n1043), .A3(n1016), .ZN(n1185) );
AND4_X1 U887 ( .A1(n1026), .A2(n1023), .A3(n1022), .A4(n1202), .ZN(n1193) );
NAND2_X1 U888 ( .A1(n1009), .A2(n1204), .ZN(n1202) );
NAND4_X1 U889 ( .A1(G902), .A2(G953), .A3(n1205), .A4(n1206), .ZN(n1204) );
INV_X1 U890 ( .A(G900), .ZN(n1206) );
XNOR2_X1 U891 ( .A(G122), .B(n1176), .ZN(G24) );
NAND4_X1 U892 ( .A1(n1207), .A2(n1028), .A3(n1050), .A4(n1192), .ZN(n1176) );
NOR2_X1 U893 ( .A1(n1022), .A2(n1203), .ZN(n1028) );
XNOR2_X1 U894 ( .A(G119), .B(n1180), .ZN(G21) );
NAND4_X1 U895 ( .A1(n1038), .A2(n1207), .A3(n1203), .A4(n1022), .ZN(n1180) );
INV_X1 U896 ( .A(n1023), .ZN(n1203) );
XNOR2_X1 U897 ( .A(G116), .B(n1208), .ZN(G18) );
NAND2_X1 U898 ( .A1(KEYINPUT32), .A2(n1209), .ZN(n1208) );
INV_X1 U899 ( .A(n1179), .ZN(n1209) );
NAND3_X1 U900 ( .A1(n1021), .A2(n1025), .A3(n1207), .ZN(n1179) );
NOR2_X1 U901 ( .A1(n1192), .A2(n1210), .ZN(n1025) );
NAND2_X1 U902 ( .A1(n1211), .A2(n1212), .ZN(G15) );
OR2_X1 U903 ( .A1(n1178), .A2(G113), .ZN(n1212) );
XOR2_X1 U904 ( .A(n1213), .B(KEYINPUT5), .Z(n1211) );
NAND2_X1 U905 ( .A1(G113), .A2(n1178), .ZN(n1213) );
NAND3_X1 U906 ( .A1(n1021), .A2(n1026), .A3(n1207), .ZN(n1178) );
AND2_X1 U907 ( .A1(n1016), .A2(n1214), .ZN(n1207) );
NOR2_X1 U908 ( .A1(n1031), .A2(n1060), .ZN(n1016) );
XNOR2_X1 U909 ( .A(n1215), .B(KEYINPUT22), .ZN(n1031) );
AND2_X1 U910 ( .A1(n1210), .A2(n1192), .ZN(n1026) );
INV_X1 U911 ( .A(n1050), .ZN(n1210) );
NOR2_X1 U912 ( .A1(n1023), .A2(n1022), .ZN(n1021) );
XOR2_X1 U913 ( .A(n1103), .B(n1216), .Z(G12) );
NOR2_X1 U914 ( .A1(G110), .A2(KEYINPUT44), .ZN(n1216) );
NAND4_X1 U915 ( .A1(n1038), .A2(n1181), .A3(n1023), .A4(n1022), .ZN(n1103) );
XNOR2_X1 U916 ( .A(n1061), .B(n1063), .ZN(n1022) );
NAND2_X1 U917 ( .A1(G217), .A2(n1217), .ZN(n1063) );
NOR2_X1 U918 ( .A1(n1111), .A2(G902), .ZN(n1061) );
INV_X1 U919 ( .A(n1108), .ZN(n1111) );
XNOR2_X1 U920 ( .A(n1218), .B(n1219), .ZN(n1108) );
XNOR2_X1 U921 ( .A(n1220), .B(n1221), .ZN(n1219) );
NAND2_X1 U922 ( .A1(KEYINPUT54), .A2(G125), .ZN(n1220) );
XOR2_X1 U923 ( .A(n1222), .B(n1223), .Z(n1218) );
XNOR2_X1 U924 ( .A(n1224), .B(n1225), .ZN(n1223) );
NOR2_X1 U925 ( .A1(KEYINPUT4), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U926 ( .A(G119), .B(G128), .ZN(n1226) );
NAND2_X1 U927 ( .A1(n1227), .A2(n1228), .ZN(n1222) );
XOR2_X1 U928 ( .A(KEYINPUT6), .B(KEYINPUT20), .Z(n1228) );
XNOR2_X1 U929 ( .A(G137), .B(n1229), .ZN(n1227) );
NAND2_X1 U930 ( .A1(G221), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U931 ( .A(n1231), .B(n1232), .ZN(n1023) );
XNOR2_X1 U932 ( .A(KEYINPUT19), .B(n1053), .ZN(n1232) );
NAND2_X1 U933 ( .A1(n1233), .A2(n1124), .ZN(n1053) );
XOR2_X1 U934 ( .A(n1234), .B(n1235), .Z(n1233) );
XNOR2_X1 U935 ( .A(n1236), .B(n1144), .ZN(n1235) );
NAND2_X1 U936 ( .A1(KEYINPUT29), .A2(n1237), .ZN(n1236) );
XOR2_X1 U937 ( .A(n1153), .B(n1238), .Z(n1237) );
NAND2_X1 U938 ( .A1(KEYINPUT47), .A2(n1154), .ZN(n1238) );
NAND3_X1 U939 ( .A1(n1239), .A2(n1034), .A3(G210), .ZN(n1153) );
XNOR2_X1 U940 ( .A(n1137), .B(n1150), .ZN(n1234) );
XNOR2_X1 U941 ( .A(n1240), .B(n1241), .ZN(n1137) );
NOR2_X1 U942 ( .A1(KEYINPUT12), .A2(G116), .ZN(n1241) );
XNOR2_X1 U943 ( .A(G113), .B(G119), .ZN(n1240) );
NAND2_X1 U944 ( .A1(KEYINPUT28), .A2(n1134), .ZN(n1231) );
INV_X1 U945 ( .A(G472), .ZN(n1134) );
AND2_X1 U946 ( .A1(n1010), .A2(n1214), .ZN(n1181) );
AND2_X1 U947 ( .A1(n1043), .A2(n1242), .ZN(n1214) );
NAND2_X1 U948 ( .A1(n1009), .A2(n1243), .ZN(n1242) );
NAND4_X1 U949 ( .A1(G902), .A2(G953), .A3(n1205), .A4(n1096), .ZN(n1243) );
INV_X1 U950 ( .A(G898), .ZN(n1096) );
NAND3_X1 U951 ( .A1(n1205), .A2(n1034), .A3(G952), .ZN(n1009) );
NAND2_X1 U952 ( .A1(G237), .A2(n1244), .ZN(n1205) );
NOR2_X1 U953 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
AND2_X1 U954 ( .A1(G214), .A2(n1245), .ZN(n1041) );
INV_X1 U955 ( .A(n1201), .ZN(n1042) );
NAND2_X1 U956 ( .A1(n1246), .A2(n1247), .ZN(n1201) );
OR2_X1 U957 ( .A1(n1248), .A2(n1064), .ZN(n1247) );
XOR2_X1 U958 ( .A(n1249), .B(KEYINPUT9), .Z(n1246) );
NAND2_X1 U959 ( .A1(n1064), .A2(n1248), .ZN(n1249) );
XOR2_X1 U960 ( .A(n1066), .B(KEYINPUT11), .Z(n1248) );
INV_X1 U961 ( .A(n1167), .ZN(n1066) );
NAND2_X1 U962 ( .A1(G210), .A2(n1245), .ZN(n1167) );
NAND2_X1 U963 ( .A1(n1239), .A2(n1124), .ZN(n1245) );
AND3_X1 U964 ( .A1(n1250), .A2(n1124), .A3(n1251), .ZN(n1064) );
XOR2_X1 U965 ( .A(KEYINPUT51), .B(n1252), .Z(n1251) );
NOR2_X1 U966 ( .A1(n1165), .A2(n1253), .ZN(n1252) );
NAND2_X1 U967 ( .A1(n1165), .A2(n1253), .ZN(n1250) );
XNOR2_X1 U968 ( .A(n1254), .B(n1189), .ZN(n1253) );
NAND2_X1 U969 ( .A1(G224), .A2(n1034), .ZN(n1189) );
NAND2_X1 U970 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NAND3_X1 U971 ( .A1(n1257), .A2(n1149), .A3(n1258), .ZN(n1256) );
INV_X1 U972 ( .A(KEYINPUT37), .ZN(n1258) );
NAND2_X1 U973 ( .A1(n1187), .A2(KEYINPUT37), .ZN(n1255) );
XOR2_X1 U974 ( .A(n1257), .B(n1149), .Z(n1187) );
INV_X1 U975 ( .A(n1144), .ZN(n1149) );
XOR2_X1 U976 ( .A(G128), .B(n1259), .Z(n1144) );
NOR2_X1 U977 ( .A1(KEYINPUT26), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U978 ( .A(G143), .B(G146), .ZN(n1260) );
XNOR2_X1 U979 ( .A(G125), .B(KEYINPUT38), .ZN(n1257) );
AND2_X1 U980 ( .A1(n1261), .A2(n1262), .ZN(n1165) );
NAND2_X1 U981 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XNOR2_X1 U982 ( .A(n1265), .B(G110), .ZN(n1264) );
INV_X1 U983 ( .A(n1266), .ZN(n1263) );
XOR2_X1 U984 ( .A(n1267), .B(KEYINPUT7), .Z(n1261) );
NAND2_X1 U985 ( .A1(n1268), .A2(n1266), .ZN(n1267) );
XNOR2_X1 U986 ( .A(n1099), .B(n1269), .ZN(n1266) );
XNOR2_X1 U987 ( .A(KEYINPUT30), .B(n1270), .ZN(n1269) );
INV_X1 U988 ( .A(G113), .ZN(n1270) );
XOR2_X1 U989 ( .A(n1271), .B(n1272), .Z(n1099) );
XOR2_X1 U990 ( .A(n1273), .B(n1274), .Z(n1271) );
NOR2_X1 U991 ( .A1(G101), .A2(KEYINPUT41), .ZN(n1274) );
NAND3_X1 U992 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1273) );
NAND2_X1 U993 ( .A1(KEYINPUT0), .A2(G116), .ZN(n1277) );
NAND3_X1 U994 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1276) );
INV_X1 U995 ( .A(KEYINPUT0), .ZN(n1279) );
OR2_X1 U996 ( .A1(n1280), .A2(n1278), .ZN(n1275) );
NOR2_X1 U997 ( .A1(G116), .A2(KEYINPUT61), .ZN(n1278) );
INV_X1 U998 ( .A(G119), .ZN(n1280) );
XNOR2_X1 U999 ( .A(G110), .B(G122), .ZN(n1268) );
NOR2_X1 U1000 ( .A1(n1215), .A2(n1060), .ZN(n1010) );
INV_X1 U1001 ( .A(n1032), .ZN(n1060) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1217), .ZN(n1032) );
NAND2_X1 U1003 ( .A1(n1244), .A2(n1124), .ZN(n1217) );
XOR2_X1 U1004 ( .A(G234), .B(KEYINPUT2), .Z(n1244) );
NAND2_X1 U1005 ( .A1(n1281), .A2(n1282), .ZN(n1215) );
NAND2_X1 U1006 ( .A1(n1283), .A2(n1058), .ZN(n1282) );
INV_X1 U1007 ( .A(G469), .ZN(n1058) );
XNOR2_X1 U1008 ( .A(KEYINPUT25), .B(n1059), .ZN(n1283) );
INV_X1 U1009 ( .A(n1284), .ZN(n1059) );
NAND2_X1 U1010 ( .A1(n1285), .A2(G469), .ZN(n1281) );
XNOR2_X1 U1011 ( .A(n1284), .B(KEYINPUT39), .ZN(n1285) );
NOR2_X1 U1012 ( .A1(n1286), .A2(n1158), .ZN(n1284) );
XNOR2_X1 U1013 ( .A(n1287), .B(n1288), .ZN(n1158) );
XNOR2_X1 U1014 ( .A(n1272), .B(n1289), .ZN(n1288) );
XNOR2_X1 U1015 ( .A(n1290), .B(n1154), .ZN(n1289) );
INV_X1 U1016 ( .A(G101), .ZN(n1154) );
NAND2_X1 U1017 ( .A1(G227), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U1018 ( .A(KEYINPUT45), .B(n1034), .ZN(n1291) );
XNOR2_X1 U1019 ( .A(G104), .B(n1292), .ZN(n1272) );
XOR2_X1 U1020 ( .A(n1293), .B(n1221), .Z(n1287) );
XOR2_X1 U1021 ( .A(G110), .B(G140), .Z(n1221) );
XNOR2_X1 U1022 ( .A(n1087), .B(n1145), .ZN(n1293) );
INV_X1 U1023 ( .A(n1150), .ZN(n1145) );
XNOR2_X1 U1024 ( .A(n1294), .B(n1295), .ZN(n1150) );
NOR2_X1 U1025 ( .A1(G137), .A2(KEYINPUT27), .ZN(n1295) );
XNOR2_X1 U1026 ( .A(G131), .B(G134), .ZN(n1294) );
XNOR2_X1 U1027 ( .A(G146), .B(n1296), .ZN(n1087) );
XNOR2_X1 U1028 ( .A(n1124), .B(KEYINPUT58), .ZN(n1286) );
NOR2_X1 U1029 ( .A1(n1050), .A2(n1192), .ZN(n1038) );
XOR2_X1 U1030 ( .A(n1056), .B(G475), .Z(n1192) );
AND2_X1 U1031 ( .A1(n1123), .A2(n1124), .ZN(n1056) );
XNOR2_X1 U1032 ( .A(n1297), .B(n1298), .ZN(n1123) );
XNOR2_X1 U1033 ( .A(n1299), .B(n1100), .ZN(n1298) );
XNOR2_X1 U1034 ( .A(G113), .B(n1265), .ZN(n1100) );
NAND2_X1 U1035 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U1036 ( .A1(n1302), .A2(n1088), .ZN(n1301) );
XOR2_X1 U1037 ( .A(n1303), .B(KEYINPUT35), .Z(n1300) );
OR2_X1 U1038 ( .A1(n1088), .A2(n1302), .ZN(n1303) );
XOR2_X1 U1039 ( .A(G143), .B(n1304), .Z(n1302) );
AND3_X1 U1040 ( .A1(G214), .A2(n1034), .A3(n1239), .ZN(n1304) );
INV_X1 U1041 ( .A(G237), .ZN(n1239) );
INV_X1 U1042 ( .A(G131), .ZN(n1088) );
XNOR2_X1 U1043 ( .A(n1305), .B(n1306), .ZN(n1297) );
INV_X1 U1044 ( .A(G104), .ZN(n1306) );
NAND2_X1 U1045 ( .A1(KEYINPUT23), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1046 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1047 ( .A(G140), .B(G125), .Z(n1309) );
XNOR2_X1 U1048 ( .A(KEYINPUT8), .B(n1224), .ZN(n1308) );
INV_X1 U1049 ( .A(G146), .ZN(n1224) );
XNOR2_X1 U1050 ( .A(n1310), .B(G478), .ZN(n1050) );
NAND2_X1 U1051 ( .A1(n1116), .A2(n1124), .ZN(n1310) );
INV_X1 U1052 ( .A(G902), .ZN(n1124) );
XOR2_X1 U1053 ( .A(n1311), .B(n1312), .Z(n1116) );
AND2_X1 U1054 ( .A1(n1230), .A2(G217), .ZN(n1312) );
AND2_X1 U1055 ( .A1(G234), .A2(n1034), .ZN(n1230) );
INV_X1 U1056 ( .A(G953), .ZN(n1034) );
NAND2_X1 U1057 ( .A1(n1313), .A2(KEYINPUT42), .ZN(n1311) );
XOR2_X1 U1058 ( .A(n1314), .B(n1315), .Z(n1313) );
XNOR2_X1 U1059 ( .A(G134), .B(n1292), .ZN(n1315) );
INV_X1 U1060 ( .A(G107), .ZN(n1292) );
XOR2_X1 U1061 ( .A(n1316), .B(n1296), .Z(n1314) );
XNOR2_X1 U1062 ( .A(n1317), .B(G143), .ZN(n1296) );
INV_X1 U1063 ( .A(G128), .ZN(n1317) );
NAND2_X1 U1064 ( .A1(KEYINPUT36), .A2(n1318), .ZN(n1316) );
XNOR2_X1 U1065 ( .A(n1265), .B(G116), .ZN(n1318) );
INV_X1 U1066 ( .A(G122), .ZN(n1265) );
endmodule


