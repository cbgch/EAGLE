//Key = 1001000001010111100001010001000001000100101110100110000001100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;

XOR2_X1 U715 ( .A(G107), .B(n998), .Z(G9) );
NAND4_X1 U716 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(G75) );
NAND4_X1 U717 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1001) );
NOR3_X1 U718 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NOR2_X1 U719 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND3_X1 U720 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1007) );
NOR3_X1 U721 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1005) );
XNOR2_X1 U722 ( .A(G469), .B(n1018), .ZN(n1017) );
NOR2_X1 U723 ( .A1(n1019), .A2(KEYINPUT41), .ZN(n1018) );
NOR2_X1 U724 ( .A1(n1020), .A2(n1021), .ZN(n1016) );
XOR2_X1 U725 ( .A(n1022), .B(n1023), .Z(n1015) );
XOR2_X1 U726 ( .A(KEYINPUT39), .B(n1024), .Z(n1023) );
NOR2_X1 U727 ( .A1(KEYINPUT17), .A2(n1025), .ZN(n1024) );
XNOR2_X1 U728 ( .A(KEYINPUT58), .B(n1026), .ZN(n1004) );
NAND2_X1 U729 ( .A1(n1027), .A2(n1028), .ZN(n1000) );
NAND2_X1 U730 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND4_X1 U731 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NAND2_X1 U732 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U733 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
OR2_X1 U734 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U735 ( .A1(n1041), .A2(n1042), .ZN(n1033) );
NAND2_X1 U736 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
XNOR2_X1 U737 ( .A(n1037), .B(KEYINPUT50), .ZN(n1043) );
NAND2_X1 U738 ( .A1(n1044), .A2(n1045), .ZN(n1029) );
NAND2_X1 U739 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND3_X1 U740 ( .A1(n1032), .A2(n1048), .A3(n1035), .ZN(n1047) );
NAND2_X1 U741 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U742 ( .A1(n1031), .A2(n1051), .ZN(n1050) );
NAND2_X1 U743 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U744 ( .A1(n1008), .A2(n1054), .ZN(n1053) );
NAND2_X1 U745 ( .A1(n1037), .A2(n1055), .ZN(n1049) );
NAND2_X1 U746 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U747 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND3_X1 U748 ( .A1(n1060), .A2(n1031), .A3(n1037), .ZN(n1046) );
INV_X1 U749 ( .A(n1061), .ZN(n1027) );
XOR2_X1 U750 ( .A(n1062), .B(n1063), .Z(G72) );
NOR2_X1 U751 ( .A1(n1064), .A2(n1002), .ZN(n1063) );
AND2_X1 U752 ( .A1(G227), .A2(G900), .ZN(n1064) );
NAND2_X1 U753 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
NAND2_X1 U754 ( .A1(n1067), .A2(n1002), .ZN(n1066) );
XOR2_X1 U755 ( .A(n1068), .B(n1069), .Z(n1067) );
NAND2_X1 U756 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
XOR2_X1 U757 ( .A(n1072), .B(KEYINPUT30), .Z(n1070) );
NAND3_X1 U758 ( .A1(G900), .A2(n1069), .A3(G953), .ZN(n1065) );
XNOR2_X1 U759 ( .A(n1073), .B(n1074), .ZN(n1069) );
XOR2_X1 U760 ( .A(n1075), .B(n1076), .Z(n1074) );
NAND3_X1 U761 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
OR2_X1 U762 ( .A1(n1080), .A2(KEYINPUT40), .ZN(n1079) );
NAND3_X1 U763 ( .A1(KEYINPUT40), .A2(n1080), .A3(G140), .ZN(n1078) );
NAND2_X1 U764 ( .A1(n1081), .A2(n1082), .ZN(n1077) );
NAND2_X1 U765 ( .A1(KEYINPUT40), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U766 ( .A(KEYINPUT61), .B(n1080), .ZN(n1083) );
INV_X1 U767 ( .A(G125), .ZN(n1080) );
NAND2_X1 U768 ( .A1(n1084), .A2(n1085), .ZN(n1075) );
OR2_X1 U769 ( .A1(n1086), .A2(G131), .ZN(n1085) );
XOR2_X1 U770 ( .A(n1087), .B(KEYINPUT48), .Z(n1084) );
NAND2_X1 U771 ( .A1(G131), .A2(n1086), .ZN(n1087) );
XOR2_X1 U772 ( .A(n1088), .B(n1089), .Z(G69) );
XOR2_X1 U773 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U774 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U775 ( .A1(G953), .A2(n1094), .ZN(n1093) );
XNOR2_X1 U776 ( .A(n1095), .B(n1096), .ZN(n1092) );
XNOR2_X1 U777 ( .A(n1097), .B(n1098), .ZN(n1096) );
NAND2_X1 U778 ( .A1(KEYINPUT37), .A2(n1099), .ZN(n1097) );
NAND2_X1 U779 ( .A1(G953), .A2(n1100), .ZN(n1090) );
NAND2_X1 U780 ( .A1(n1101), .A2(G898), .ZN(n1100) );
XNOR2_X1 U781 ( .A(G224), .B(KEYINPUT49), .ZN(n1101) );
NOR2_X1 U782 ( .A1(n1102), .A2(G953), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1103), .A2(n1104), .ZN(G66) );
XOR2_X1 U784 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR3_X1 U785 ( .A1(n1107), .A2(KEYINPUT26), .A3(n1011), .ZN(n1105) );
NOR2_X1 U786 ( .A1(n1103), .A2(n1108), .ZN(G63) );
XOR2_X1 U787 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U788 ( .A1(n1111), .A2(KEYINPUT10), .ZN(n1109) );
NOR2_X1 U789 ( .A1(n1021), .A2(n1107), .ZN(n1111) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1112), .ZN(G60) );
XOR2_X1 U791 ( .A(n1113), .B(n1114), .Z(n1112) );
AND2_X1 U792 ( .A1(G475), .A2(n1115), .ZN(n1113) );
XOR2_X1 U793 ( .A(n1116), .B(n1117), .Z(G6) );
NOR2_X1 U794 ( .A1(KEYINPUT29), .A2(n1118), .ZN(n1117) );
NOR2_X1 U795 ( .A1(n1103), .A2(n1119), .ZN(G57) );
XOR2_X1 U796 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U797 ( .A1(KEYINPUT19), .A2(n1122), .ZN(n1121) );
XNOR2_X1 U798 ( .A(G101), .B(n1123), .ZN(n1120) );
NOR2_X1 U799 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U800 ( .A(KEYINPUT52), .B(n1126), .Z(n1125) );
AND2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U802 ( .A1(n1128), .A2(n1127), .ZN(n1124) );
NAND2_X1 U803 ( .A1(n1115), .A2(G472), .ZN(n1127) );
XOR2_X1 U804 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR3_X1 U805 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(G54) );
AND3_X1 U806 ( .A1(KEYINPUT38), .A2(G953), .A3(G952), .ZN(n1133) );
NOR2_X1 U807 ( .A1(KEYINPUT38), .A2(n1134), .ZN(n1132) );
INV_X1 U808 ( .A(n1103), .ZN(n1134) );
XOR2_X1 U809 ( .A(n1135), .B(n1136), .Z(n1131) );
XOR2_X1 U810 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U811 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U812 ( .A1(KEYINPUT31), .A2(n1141), .ZN(n1140) );
NOR3_X1 U813 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1139) );
AND2_X1 U814 ( .A1(n1145), .A2(KEYINPUT56), .ZN(n1144) );
NOR3_X1 U815 ( .A1(KEYINPUT56), .A2(n1145), .A3(n1146), .ZN(n1143) );
INV_X1 U816 ( .A(n1147), .ZN(n1145) );
NOR2_X1 U817 ( .A1(n1148), .A2(n1107), .ZN(n1137) );
INV_X1 U818 ( .A(n1115), .ZN(n1107) );
XNOR2_X1 U819 ( .A(n1073), .B(n1149), .ZN(n1135) );
NOR2_X1 U820 ( .A1(n1103), .A2(n1150), .ZN(G51) );
NOR2_X1 U821 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U822 ( .A(KEYINPUT22), .B(n1153), .Z(n1152) );
NOR2_X1 U823 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
AND2_X1 U824 ( .A1(n1155), .A2(n1154), .ZN(n1151) );
XOR2_X1 U825 ( .A(n1156), .B(n1157), .Z(n1154) );
XNOR2_X1 U826 ( .A(n1158), .B(n1159), .ZN(n1157) );
XNOR2_X1 U827 ( .A(n1160), .B(KEYINPUT23), .ZN(n1156) );
NAND2_X1 U828 ( .A1(n1115), .A2(n1025), .ZN(n1155) );
NOR2_X1 U829 ( .A1(n1161), .A2(n999), .ZN(n1115) );
AND3_X1 U830 ( .A1(n1102), .A2(n1072), .A3(n1071), .ZN(n999) );
AND4_X1 U831 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1071) );
NOR4_X1 U832 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
INV_X1 U833 ( .A(n1170), .ZN(n1167) );
NAND2_X1 U834 ( .A1(n1171), .A2(n1172), .ZN(n1164) );
AND4_X1 U835 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1102) );
NOR4_X1 U836 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
AND2_X1 U837 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U838 ( .A1(n998), .A2(n1116), .ZN(n1175) );
AND3_X1 U839 ( .A1(n1183), .A2(n1184), .A3(n1039), .ZN(n1116) );
AND3_X1 U840 ( .A1(n1040), .A2(n1184), .A3(n1183), .ZN(n998) );
NOR4_X1 U841 ( .A1(n1056), .A2(n1052), .A3(n1042), .A4(n1185), .ZN(n1183) );
NOR2_X1 U842 ( .A1(n1002), .A2(G952), .ZN(n1103) );
XNOR2_X1 U843 ( .A(G146), .B(n1186), .ZN(G48) );
NAND2_X1 U844 ( .A1(n1172), .A2(n1187), .ZN(n1186) );
XOR2_X1 U845 ( .A(KEYINPUT25), .B(n1171), .Z(n1187) );
AND2_X1 U846 ( .A1(n1039), .A2(n1188), .ZN(n1171) );
XNOR2_X1 U847 ( .A(G143), .B(n1163), .ZN(G45) );
NAND3_X1 U848 ( .A1(n1060), .A2(n1189), .A3(n1190), .ZN(n1163) );
NOR3_X1 U849 ( .A1(n1056), .A2(n1191), .A3(n1026), .ZN(n1190) );
INV_X1 U850 ( .A(n1172), .ZN(n1056) );
XNOR2_X1 U851 ( .A(n1082), .B(n1169), .ZN(G42) );
AND4_X1 U852 ( .A1(n1032), .A2(n1042), .A3(n1189), .A4(n1192), .ZN(n1169) );
NOR2_X1 U853 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XNOR2_X1 U854 ( .A(n1195), .B(n1168), .ZN(G39) );
AND3_X1 U855 ( .A1(n1031), .A2(n1188), .A3(n1044), .ZN(n1168) );
XOR2_X1 U856 ( .A(n1196), .B(G134), .Z(G36) );
NAND2_X1 U857 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
OR2_X1 U858 ( .A1(n1162), .A2(KEYINPUT35), .ZN(n1198) );
NAND3_X1 U859 ( .A1(n1031), .A2(n1189), .A3(n1181), .ZN(n1162) );
NAND4_X1 U860 ( .A1(n1199), .A2(n1181), .A3(n1200), .A4(KEYINPUT35), .ZN(n1197) );
NOR2_X1 U861 ( .A1(n1052), .A2(n1193), .ZN(n1200) );
XNOR2_X1 U862 ( .A(G131), .B(n1170), .ZN(G33) );
NAND4_X1 U863 ( .A1(n1060), .A2(n1039), .A3(n1031), .A4(n1189), .ZN(n1170) );
INV_X1 U864 ( .A(n1193), .ZN(n1031) );
NAND2_X1 U865 ( .A1(n1059), .A2(n1014), .ZN(n1193) );
XNOR2_X1 U866 ( .A(n1201), .B(KEYINPUT20), .ZN(n1059) );
XOR2_X1 U867 ( .A(G128), .B(n1166), .Z(G30) );
AND3_X1 U868 ( .A1(n1040), .A2(n1172), .A3(n1188), .ZN(n1166) );
AND3_X1 U869 ( .A1(n1185), .A2(n1042), .A3(n1189), .ZN(n1188) );
NOR2_X1 U870 ( .A1(n1052), .A2(n1199), .ZN(n1189) );
INV_X1 U871 ( .A(n1202), .ZN(n1052) );
XOR2_X1 U872 ( .A(G101), .B(n1179), .Z(G3) );
AND2_X1 U873 ( .A1(n1203), .A2(n1060), .ZN(n1179) );
XNOR2_X1 U874 ( .A(G125), .B(n1072), .ZN(G27) );
NAND4_X1 U875 ( .A1(n1039), .A2(n1172), .A3(n1037), .A4(n1204), .ZN(n1072) );
NOR3_X1 U876 ( .A1(n1185), .A2(n1035), .A3(n1199), .ZN(n1204) );
AND2_X1 U877 ( .A1(n1061), .A2(n1205), .ZN(n1199) );
NAND4_X1 U878 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1207), .ZN(n1205) );
INV_X1 U879 ( .A(G900), .ZN(n1207) );
XOR2_X1 U880 ( .A(G122), .B(n1178), .Z(G24) );
AND3_X1 U881 ( .A1(n1182), .A2(n1035), .A3(n1208), .ZN(n1178) );
NOR3_X1 U882 ( .A1(n1026), .A2(n1185), .A3(n1191), .ZN(n1208) );
INV_X1 U883 ( .A(n1209), .ZN(n1026) );
INV_X1 U884 ( .A(n1042), .ZN(n1035) );
XNOR2_X1 U885 ( .A(G119), .B(n1173), .ZN(G21) );
NAND4_X1 U886 ( .A1(n1182), .A2(n1044), .A3(n1185), .A4(n1042), .ZN(n1173) );
INV_X1 U887 ( .A(n1032), .ZN(n1185) );
XOR2_X1 U888 ( .A(n1210), .B(n1211), .Z(G18) );
XNOR2_X1 U889 ( .A(G116), .B(KEYINPUT5), .ZN(n1211) );
NAND4_X1 U890 ( .A1(n1212), .A2(n1037), .A3(n1213), .A4(n1181), .ZN(n1210) );
AND2_X1 U891 ( .A1(n1060), .A2(n1040), .ZN(n1181) );
NOR2_X1 U892 ( .A1(n1209), .A2(n1191), .ZN(n1040) );
XOR2_X1 U893 ( .A(n1214), .B(KEYINPUT3), .Z(n1191) );
NOR2_X1 U894 ( .A1(KEYINPUT7), .A2(n1215), .ZN(n1213) );
INV_X1 U895 ( .A(n1184), .ZN(n1215) );
XNOR2_X1 U896 ( .A(n1172), .B(KEYINPUT44), .ZN(n1212) );
XNOR2_X1 U897 ( .A(G113), .B(n1174), .ZN(G15) );
NAND3_X1 U898 ( .A1(n1060), .A2(n1039), .A3(n1182), .ZN(n1174) );
AND3_X1 U899 ( .A1(n1172), .A2(n1184), .A3(n1037), .ZN(n1182) );
NOR2_X1 U900 ( .A1(n1216), .A2(n1008), .ZN(n1037) );
INV_X1 U901 ( .A(n1054), .ZN(n1216) );
INV_X1 U902 ( .A(n1194), .ZN(n1039) );
NAND2_X1 U903 ( .A1(n1217), .A2(n1209), .ZN(n1194) );
XOR2_X1 U904 ( .A(n1214), .B(KEYINPUT14), .Z(n1217) );
NOR2_X1 U905 ( .A1(n1032), .A2(n1042), .ZN(n1060) );
NAND3_X1 U906 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(G12) );
NAND2_X1 U907 ( .A1(KEYINPUT60), .A2(n1221), .ZN(n1220) );
NAND3_X1 U908 ( .A1(G110), .A2(n1222), .A3(n1223), .ZN(n1219) );
NAND2_X1 U909 ( .A1(n1177), .A2(n1224), .ZN(n1218) );
NAND2_X1 U910 ( .A1(n1225), .A2(n1222), .ZN(n1224) );
INV_X1 U911 ( .A(KEYINPUT60), .ZN(n1222) );
XNOR2_X1 U912 ( .A(KEYINPUT28), .B(n1221), .ZN(n1225) );
INV_X1 U913 ( .A(G110), .ZN(n1221) );
INV_X1 U914 ( .A(n1223), .ZN(n1177) );
NAND3_X1 U915 ( .A1(n1032), .A2(n1042), .A3(n1203), .ZN(n1223) );
AND4_X1 U916 ( .A1(n1044), .A2(n1172), .A3(n1202), .A4(n1184), .ZN(n1203) );
NAND2_X1 U917 ( .A1(n1061), .A2(n1226), .ZN(n1184) );
NAND4_X1 U918 ( .A1(G953), .A2(G902), .A3(n1206), .A4(n1094), .ZN(n1226) );
INV_X1 U919 ( .A(G898), .ZN(n1094) );
NAND3_X1 U920 ( .A1(n1206), .A2(n1002), .A3(G952), .ZN(n1061) );
NAND2_X1 U921 ( .A1(G237), .A2(G234), .ZN(n1206) );
NOR2_X1 U922 ( .A1(n1054), .A2(n1008), .ZN(n1202) );
AND2_X1 U923 ( .A1(G221), .A2(n1227), .ZN(n1008) );
XOR2_X1 U924 ( .A(n1019), .B(n1148), .Z(n1054) );
INV_X1 U925 ( .A(G469), .ZN(n1148) );
AND2_X1 U926 ( .A1(n1228), .A2(n1161), .ZN(n1019) );
NAND2_X1 U927 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NAND2_X1 U928 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XNOR2_X1 U929 ( .A(n1147), .B(n1233), .ZN(n1232) );
XOR2_X1 U930 ( .A(n1234), .B(n1149), .Z(n1231) );
XOR2_X1 U931 ( .A(n1235), .B(KEYINPUT53), .Z(n1229) );
NAND3_X1 U932 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1235) );
XNOR2_X1 U933 ( .A(n1149), .B(n1234), .ZN(n1238) );
XOR2_X1 U934 ( .A(n1141), .B(n1239), .Z(n1234) );
NOR2_X1 U935 ( .A1(KEYINPUT62), .A2(n1073), .ZN(n1239) );
XOR2_X1 U936 ( .A(G128), .B(n1240), .Z(n1073) );
NOR2_X1 U937 ( .A1(KEYINPUT4), .A2(n1241), .ZN(n1240) );
XNOR2_X1 U938 ( .A(G146), .B(n1242), .ZN(n1241) );
NOR2_X1 U939 ( .A1(G143), .A2(KEYINPUT32), .ZN(n1242) );
INV_X1 U940 ( .A(n1142), .ZN(n1237) );
NOR2_X1 U941 ( .A1(n1147), .A2(n1233), .ZN(n1142) );
NAND2_X1 U942 ( .A1(n1233), .A2(n1147), .ZN(n1236) );
NAND2_X1 U943 ( .A1(G227), .A2(n1002), .ZN(n1147) );
NOR2_X1 U944 ( .A1(n1243), .A2(n1058), .ZN(n1172) );
INV_X1 U945 ( .A(n1014), .ZN(n1058) );
NAND2_X1 U946 ( .A1(G214), .A2(n1244), .ZN(n1014) );
INV_X1 U947 ( .A(n1201), .ZN(n1243) );
XNOR2_X1 U948 ( .A(n1022), .B(n1025), .ZN(n1201) );
AND2_X1 U949 ( .A1(G210), .A2(n1244), .ZN(n1025) );
NAND2_X1 U950 ( .A1(n1245), .A2(n1161), .ZN(n1244) );
INV_X1 U951 ( .A(G237), .ZN(n1245) );
NAND2_X1 U952 ( .A1(n1246), .A2(n1161), .ZN(n1022) );
XOR2_X1 U953 ( .A(n1158), .B(n1247), .Z(n1246) );
NOR2_X1 U954 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XOR2_X1 U955 ( .A(n1250), .B(KEYINPUT9), .Z(n1249) );
NAND2_X1 U956 ( .A1(n1251), .A2(n1159), .ZN(n1250) );
NOR2_X1 U957 ( .A1(n1251), .A2(n1159), .ZN(n1248) );
XNOR2_X1 U958 ( .A(n1252), .B(n1253), .ZN(n1159) );
XNOR2_X1 U959 ( .A(KEYINPUT34), .B(n1160), .ZN(n1251) );
AND2_X1 U960 ( .A1(G224), .A2(n1002), .ZN(n1160) );
XNOR2_X1 U961 ( .A(n1099), .B(n1254), .ZN(n1158) );
NOR2_X1 U962 ( .A1(KEYINPUT47), .A2(n1255), .ZN(n1254) );
NOR2_X1 U963 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U964 ( .A(KEYINPUT8), .B(n1258), .Z(n1257) );
NOR2_X1 U965 ( .A1(n1259), .A2(n1098), .ZN(n1258) );
XNOR2_X1 U966 ( .A(n1260), .B(KEYINPUT63), .ZN(n1259) );
INV_X1 U967 ( .A(n1095), .ZN(n1260) );
NOR2_X1 U968 ( .A1(n1261), .A2(n1262), .ZN(n1256) );
XNOR2_X1 U969 ( .A(KEYINPUT63), .B(n1095), .ZN(n1262) );
XNOR2_X1 U970 ( .A(n1263), .B(G113), .ZN(n1095) );
INV_X1 U971 ( .A(n1098), .ZN(n1261) );
XNOR2_X1 U972 ( .A(n1141), .B(KEYINPUT21), .ZN(n1098) );
XNOR2_X1 U973 ( .A(G101), .B(n1264), .ZN(n1141) );
XNOR2_X1 U974 ( .A(G107), .B(n1118), .ZN(n1264) );
XOR2_X1 U975 ( .A(G110), .B(n1265), .Z(n1099) );
NOR2_X1 U976 ( .A1(G122), .A2(KEYINPUT1), .ZN(n1265) );
NOR2_X1 U977 ( .A1(n1209), .A2(n1214), .ZN(n1044) );
NAND3_X1 U978 ( .A1(n1266), .A2(n1267), .A3(n1013), .ZN(n1214) );
NAND2_X1 U979 ( .A1(n1020), .A2(n1021), .ZN(n1013) );
INV_X1 U980 ( .A(G478), .ZN(n1021) );
INV_X1 U981 ( .A(n1268), .ZN(n1020) );
OR2_X1 U982 ( .A1(G478), .A2(KEYINPUT0), .ZN(n1267) );
NAND3_X1 U983 ( .A1(G478), .A2(n1268), .A3(KEYINPUT0), .ZN(n1266) );
NAND2_X1 U984 ( .A1(n1110), .A2(n1161), .ZN(n1268) );
XNOR2_X1 U985 ( .A(n1269), .B(n1270), .ZN(n1110) );
XOR2_X1 U986 ( .A(n1271), .B(n1272), .Z(n1270) );
XNOR2_X1 U987 ( .A(G134), .B(G122), .ZN(n1272) );
NAND3_X1 U988 ( .A1(G217), .A2(n1002), .A3(n1273), .ZN(n1271) );
XNOR2_X1 U989 ( .A(n1253), .B(n1274), .ZN(n1269) );
XOR2_X1 U990 ( .A(n1275), .B(n1276), .Z(n1274) );
NOR2_X1 U991 ( .A1(G107), .A2(KEYINPUT54), .ZN(n1275) );
XNOR2_X1 U992 ( .A(n1277), .B(G475), .ZN(n1209) );
OR2_X1 U993 ( .A1(n1114), .A2(G902), .ZN(n1277) );
XNOR2_X1 U994 ( .A(n1278), .B(n1279), .ZN(n1114) );
XOR2_X1 U995 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U996 ( .A(n1282), .B(n1118), .ZN(n1281) );
INV_X1 U997 ( .A(G104), .ZN(n1118) );
NAND2_X1 U998 ( .A1(n1283), .A2(G214), .ZN(n1282) );
XNOR2_X1 U999 ( .A(G122), .B(G140), .ZN(n1280) );
XOR2_X1 U1000 ( .A(n1284), .B(n1285), .Z(n1278) );
XOR2_X1 U1001 ( .A(n1286), .B(n1287), .Z(n1285) );
NOR2_X1 U1002 ( .A1(KEYINPUT36), .A2(n1288), .ZN(n1286) );
XOR2_X1 U1003 ( .A(n1289), .B(n1290), .Z(n1284) );
NOR2_X1 U1004 ( .A1(G113), .A2(KEYINPUT24), .ZN(n1290) );
NAND2_X1 U1005 ( .A1(KEYINPUT42), .A2(n1291), .ZN(n1289) );
INV_X1 U1006 ( .A(G131), .ZN(n1291) );
NAND3_X1 U1007 ( .A1(n1292), .A2(n1293), .A3(n1012), .ZN(n1042) );
NAND2_X1 U1008 ( .A1(n1010), .A2(n1011), .ZN(n1012) );
NAND2_X1 U1009 ( .A1(KEYINPUT12), .A2(n1011), .ZN(n1293) );
OR3_X1 U1010 ( .A1(n1010), .A2(KEYINPUT12), .A3(n1011), .ZN(n1292) );
NAND2_X1 U1011 ( .A1(G217), .A2(n1227), .ZN(n1011) );
NAND2_X1 U1012 ( .A1(G234), .A2(n1161), .ZN(n1227) );
NOR2_X1 U1013 ( .A1(n1106), .A2(G902), .ZN(n1010) );
XNOR2_X1 U1014 ( .A(n1294), .B(n1295), .ZN(n1106) );
AND3_X1 U1015 ( .A1(n1273), .A2(n1002), .A3(G221), .ZN(n1295) );
INV_X1 U1016 ( .A(G953), .ZN(n1002) );
XNOR2_X1 U1017 ( .A(G234), .B(KEYINPUT13), .ZN(n1273) );
XNOR2_X1 U1018 ( .A(n1296), .B(n1297), .ZN(n1294) );
NOR2_X1 U1019 ( .A1(KEYINPUT55), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U1020 ( .A(G137), .B(KEYINPUT57), .ZN(n1298) );
NOR2_X1 U1021 ( .A1(KEYINPUT6), .A2(n1299), .ZN(n1296) );
XOR2_X1 U1022 ( .A(n1300), .B(n1301), .Z(n1299) );
XNOR2_X1 U1023 ( .A(n1287), .B(n1146), .ZN(n1301) );
INV_X1 U1024 ( .A(n1233), .ZN(n1146) );
XNOR2_X1 U1025 ( .A(G110), .B(n1082), .ZN(n1233) );
INV_X1 U1026 ( .A(G140), .ZN(n1082) );
XNOR2_X1 U1027 ( .A(n1252), .B(KEYINPUT27), .ZN(n1287) );
XNOR2_X1 U1028 ( .A(G125), .B(G146), .ZN(n1252) );
XOR2_X1 U1029 ( .A(n1302), .B(KEYINPUT45), .Z(n1300) );
NAND2_X1 U1030 ( .A1(n1303), .A2(KEYINPUT43), .ZN(n1302) );
XNOR2_X1 U1031 ( .A(G119), .B(G128), .ZN(n1303) );
XNOR2_X1 U1032 ( .A(n1003), .B(KEYINPUT11), .ZN(n1032) );
XOR2_X1 U1033 ( .A(n1304), .B(G472), .Z(n1003) );
NAND2_X1 U1034 ( .A1(n1305), .A2(n1161), .ZN(n1304) );
INV_X1 U1035 ( .A(G902), .ZN(n1161) );
XOR2_X1 U1036 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1037 ( .A(n1122), .B(n1308), .Z(n1307) );
NOR2_X1 U1038 ( .A1(KEYINPUT2), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1039 ( .A(n1130), .B(n1310), .ZN(n1309) );
NOR2_X1 U1040 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NOR2_X1 U1041 ( .A1(KEYINPUT46), .A2(n1129), .ZN(n1312) );
NOR2_X1 U1042 ( .A1(KEYINPUT18), .A2(n1313), .ZN(n1311) );
INV_X1 U1043 ( .A(n1129), .ZN(n1313) );
XNOR2_X1 U1044 ( .A(n1314), .B(n1263), .ZN(n1129) );
XOR2_X1 U1045 ( .A(G119), .B(n1276), .Z(n1263) );
XOR2_X1 U1046 ( .A(G116), .B(KEYINPUT15), .Z(n1276) );
NAND2_X1 U1047 ( .A1(KEYINPUT33), .A2(G113), .ZN(n1314) );
XNOR2_X1 U1048 ( .A(n1315), .B(n1149), .ZN(n1130) );
XNOR2_X1 U1049 ( .A(n1316), .B(n1086), .ZN(n1149) );
XNOR2_X1 U1050 ( .A(G134), .B(n1195), .ZN(n1086) );
INV_X1 U1051 ( .A(G137), .ZN(n1195) );
XNOR2_X1 U1052 ( .A(G131), .B(KEYINPUT51), .ZN(n1316) );
XNOR2_X1 U1053 ( .A(G146), .B(n1253), .ZN(n1315) );
XNOR2_X1 U1054 ( .A(G128), .B(n1288), .ZN(n1253) );
INV_X1 U1055 ( .A(G143), .ZN(n1288) );
NAND2_X1 U1056 ( .A1(n1317), .A2(n1283), .ZN(n1122) );
NOR2_X1 U1057 ( .A1(G953), .A2(G237), .ZN(n1283) );
XNOR2_X1 U1058 ( .A(G210), .B(KEYINPUT16), .ZN(n1317) );
XNOR2_X1 U1059 ( .A(G101), .B(KEYINPUT59), .ZN(n1306) );
endmodule


