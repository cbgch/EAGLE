//Key = 0101101111110001000000000001110111010011011011000100101110100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
n1385, n1386, n1387;

XOR2_X1 U774 ( .A(G107), .B(n1065), .Z(G9) );
NOR2_X1 U775 ( .A1(n1066), .A2(n1067), .ZN(G75) );
NOR3_X1 U776 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NAND3_X1 U777 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1068) );
NAND2_X1 U778 ( .A1(n1074), .A2(n1075), .ZN(n1071) );
NAND2_X1 U779 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND3_X1 U780 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
NAND2_X1 U781 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
NAND2_X1 U782 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
OR2_X1 U783 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U784 ( .A1(n1087), .A2(n1088), .ZN(n1081) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND3_X1 U786 ( .A1(n1083), .A2(n1091), .A3(n1087), .ZN(n1076) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U788 ( .A1(n1078), .A2(n1094), .ZN(n1093) );
NAND2_X1 U789 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U790 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U791 ( .A(n1099), .B(KEYINPUT7), .Z(n1097) );
INV_X1 U792 ( .A(n1100), .ZN(n1095) );
NAND2_X1 U793 ( .A1(n1080), .A2(n1101), .ZN(n1092) );
NAND2_X1 U794 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U795 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
INV_X1 U796 ( .A(n1106), .ZN(n1074) );
AND3_X1 U797 ( .A1(n1073), .A2(n1072), .A3(n1107), .ZN(n1066) );
XOR2_X1 U798 ( .A(G952), .B(KEYINPUT28), .Z(n1107) );
NAND4_X1 U799 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1072) );
NOR4_X1 U800 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1111) );
XOR2_X1 U801 ( .A(n1116), .B(KEYINPUT15), .Z(n1114) );
XOR2_X1 U802 ( .A(KEYINPUT51), .B(n1117), .Z(n1113) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XNOR2_X1 U805 ( .A(n1122), .B(KEYINPUT17), .ZN(n1121) );
NOR2_X1 U806 ( .A1(n1123), .A2(n1122), .ZN(n1118) );
XNOR2_X1 U807 ( .A(n1124), .B(KEYINPUT25), .ZN(n1122) );
XNOR2_X1 U808 ( .A(n1125), .B(KEYINPUT62), .ZN(n1112) );
NOR3_X1 U809 ( .A1(n1098), .A2(n1126), .A3(n1127), .ZN(n1110) );
XOR2_X1 U810 ( .A(n1128), .B(n1129), .Z(n1108) );
NOR2_X1 U811 ( .A1(n1130), .A2(KEYINPUT20), .ZN(n1129) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(G72) );
XOR2_X1 U813 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR3_X1 U814 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1134) );
NOR2_X1 U815 ( .A1(G900), .A2(n1138), .ZN(n1137) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
XOR2_X1 U817 ( .A(n1141), .B(KEYINPUT42), .Z(n1135) );
NAND2_X1 U818 ( .A1(n1139), .A2(n1140), .ZN(n1141) );
XOR2_X1 U819 ( .A(G125), .B(G140), .Z(n1140) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1139) );
NAND2_X1 U821 ( .A1(KEYINPUT56), .A2(n1144), .ZN(n1142) );
XOR2_X1 U822 ( .A(n1145), .B(n1146), .Z(n1144) );
XNOR2_X1 U823 ( .A(n1147), .B(n1148), .ZN(n1146) );
NOR2_X1 U824 ( .A1(G131), .A2(KEYINPUT0), .ZN(n1148) );
NAND2_X1 U825 ( .A1(KEYINPUT32), .A2(n1149), .ZN(n1147) );
NOR2_X1 U826 ( .A1(G953), .A2(n1150), .ZN(n1133) );
NOR3_X1 U827 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
XOR2_X1 U828 ( .A(n1154), .B(KEYINPUT3), .Z(n1152) );
XNOR2_X1 U829 ( .A(KEYINPUT57), .B(n1155), .ZN(n1151) );
NOR2_X1 U830 ( .A1(n1156), .A2(n1138), .ZN(n1131) );
AND2_X1 U831 ( .A1(G227), .A2(G900), .ZN(n1156) );
XOR2_X1 U832 ( .A(n1157), .B(n1158), .Z(G69) );
NOR2_X1 U833 ( .A1(n1159), .A2(n1138), .ZN(n1158) );
AND2_X1 U834 ( .A1(G224), .A2(G898), .ZN(n1159) );
NAND2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NAND2_X1 U836 ( .A1(n1162), .A2(n1138), .ZN(n1161) );
XNOR2_X1 U837 ( .A(n1163), .B(n1164), .ZN(n1162) );
NOR3_X1 U838 ( .A1(n1165), .A2(n1065), .A3(n1166), .ZN(n1163) );
XOR2_X1 U839 ( .A(n1167), .B(KEYINPUT47), .Z(n1166) );
INV_X1 U840 ( .A(n1168), .ZN(n1065) );
NAND3_X1 U841 ( .A1(G898), .A2(n1164), .A3(G953), .ZN(n1160) );
NAND2_X1 U842 ( .A1(n1169), .A2(n1170), .ZN(n1164) );
NAND2_X1 U843 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
INV_X1 U844 ( .A(KEYINPUT31), .ZN(n1172) );
XOR2_X1 U845 ( .A(n1173), .B(n1174), .Z(n1171) );
NAND2_X1 U846 ( .A1(KEYINPUT31), .A2(n1175), .ZN(n1169) );
XOR2_X1 U847 ( .A(n1176), .B(n1177), .Z(n1175) );
INV_X1 U848 ( .A(n1173), .ZN(n1177) );
XOR2_X1 U849 ( .A(n1178), .B(n1179), .Z(n1173) );
XOR2_X1 U850 ( .A(KEYINPUT24), .B(G122), .Z(n1179) );
NOR2_X1 U851 ( .A1(n1180), .A2(n1181), .ZN(G66) );
XNOR2_X1 U852 ( .A(n1182), .B(n1183), .ZN(n1181) );
NOR2_X1 U853 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U854 ( .A1(n1180), .A2(n1186), .ZN(G63) );
XOR2_X1 U855 ( .A(n1187), .B(n1188), .Z(n1186) );
AND2_X1 U856 ( .A1(G478), .A2(n1189), .ZN(n1187) );
NOR3_X1 U857 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(G60) );
AND2_X1 U858 ( .A1(KEYINPUT52), .A2(n1180), .ZN(n1192) );
NOR3_X1 U859 ( .A1(KEYINPUT52), .A2(n1138), .A3(n1069), .ZN(n1191) );
INV_X1 U860 ( .A(G952), .ZN(n1069) );
XOR2_X1 U861 ( .A(n1193), .B(n1194), .Z(n1190) );
NOR2_X1 U862 ( .A1(n1195), .A2(n1185), .ZN(n1194) );
XOR2_X1 U863 ( .A(n1124), .B(KEYINPUT61), .Z(n1195) );
XOR2_X1 U864 ( .A(n1196), .B(n1197), .Z(G6) );
NAND2_X1 U865 ( .A1(KEYINPUT55), .A2(G104), .ZN(n1197) );
NOR2_X1 U866 ( .A1(n1180), .A2(n1198), .ZN(G57) );
XOR2_X1 U867 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U868 ( .A(n1201), .B(n1202), .Z(n1200) );
NOR2_X1 U869 ( .A1(G101), .A2(KEYINPUT50), .ZN(n1201) );
XOR2_X1 U870 ( .A(n1203), .B(n1204), .Z(n1199) );
NOR3_X1 U871 ( .A1(n1185), .A2(KEYINPUT37), .A3(n1205), .ZN(n1204) );
INV_X1 U872 ( .A(G472), .ZN(n1205) );
NOR2_X1 U873 ( .A1(n1180), .A2(n1206), .ZN(G54) );
XOR2_X1 U874 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U875 ( .A(n1209), .B(n1210), .Z(n1208) );
XOR2_X1 U876 ( .A(n1143), .B(n1211), .Z(n1207) );
XOR2_X1 U877 ( .A(n1212), .B(n1213), .Z(n1211) );
NAND2_X1 U878 ( .A1(n1189), .A2(G469), .ZN(n1213) );
INV_X1 U879 ( .A(n1185), .ZN(n1189) );
NAND3_X1 U880 ( .A1(n1214), .A2(n1215), .A3(KEYINPUT58), .ZN(n1212) );
NAND2_X1 U881 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
XOR2_X1 U882 ( .A(n1218), .B(n1219), .Z(n1216) );
OR3_X1 U883 ( .A1(n1218), .A2(n1219), .A3(n1217), .ZN(n1214) );
INV_X1 U884 ( .A(KEYINPUT30), .ZN(n1217) );
XOR2_X1 U885 ( .A(n1178), .B(n1220), .Z(n1219) );
NOR2_X1 U886 ( .A1(n1180), .A2(n1221), .ZN(G51) );
XOR2_X1 U887 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U888 ( .A1(n1224), .A2(n1185), .ZN(n1223) );
NAND2_X1 U889 ( .A1(G902), .A2(n1070), .ZN(n1185) );
NAND4_X1 U890 ( .A1(n1154), .A2(n1168), .A3(n1155), .A4(n1225), .ZN(n1070) );
NOR3_X1 U891 ( .A1(n1167), .A2(n1165), .A3(n1153), .ZN(n1225) );
NAND4_X1 U892 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1153) );
AND3_X1 U893 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1229) );
NAND2_X1 U894 ( .A1(n1078), .A2(n1233), .ZN(n1228) );
XOR2_X1 U895 ( .A(KEYINPUT36), .B(n1234), .Z(n1233) );
NOR2_X1 U896 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND3_X1 U897 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1226) );
XOR2_X1 U898 ( .A(KEYINPUT60), .B(n1085), .Z(n1238) );
NAND3_X1 U899 ( .A1(n1196), .A2(n1240), .A3(n1241), .ZN(n1165) );
NAND3_X1 U900 ( .A1(n1087), .A2(n1242), .A3(n1239), .ZN(n1241) );
NAND3_X1 U901 ( .A1(n1083), .A2(n1242), .A3(n1085), .ZN(n1196) );
NAND4_X1 U902 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1167) );
OR2_X1 U903 ( .A1(n1247), .A2(n1102), .ZN(n1243) );
OR2_X1 U904 ( .A1(n1248), .A2(n1249), .ZN(n1155) );
XOR2_X1 U905 ( .A(KEYINPUT33), .B(n1250), .Z(n1249) );
NAND3_X1 U906 ( .A1(n1083), .A2(n1242), .A3(n1086), .ZN(n1168) );
NOR2_X1 U907 ( .A1(n1251), .A2(n1252), .ZN(n1222) );
XOR2_X1 U908 ( .A(n1253), .B(KEYINPUT44), .Z(n1252) );
NAND2_X1 U909 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NOR2_X1 U910 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
XOR2_X1 U911 ( .A(G125), .B(n1256), .Z(n1255) );
XOR2_X1 U912 ( .A(n1257), .B(n1258), .Z(n1254) );
XNOR2_X1 U913 ( .A(G122), .B(KEYINPUT26), .ZN(n1257) );
NOR2_X1 U914 ( .A1(n1138), .A2(G952), .ZN(n1180) );
XOR2_X1 U915 ( .A(n1227), .B(n1259), .Z(G48) );
NAND2_X1 U916 ( .A1(KEYINPUT29), .A2(G146), .ZN(n1259) );
NAND3_X1 U917 ( .A1(n1085), .A2(n1260), .A3(n1261), .ZN(n1227) );
XOR2_X1 U918 ( .A(G143), .B(n1262), .Z(G45) );
NOR2_X1 U919 ( .A1(n1263), .A2(n1248), .ZN(n1262) );
NAND4_X1 U920 ( .A1(n1100), .A2(n1264), .A3(n1260), .A4(n1265), .ZN(n1248) );
NOR2_X1 U921 ( .A1(n1090), .A2(n1266), .ZN(n1265) );
NAND3_X1 U922 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(G42) );
NAND2_X1 U923 ( .A1(G140), .A2(n1270), .ZN(n1269) );
NAND2_X1 U924 ( .A1(n1271), .A2(n1272), .ZN(n1268) );
INV_X1 U925 ( .A(KEYINPUT54), .ZN(n1272) );
NAND2_X1 U926 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
XOR2_X1 U927 ( .A(KEYINPUT4), .B(G140), .Z(n1274) );
NAND2_X1 U928 ( .A1(KEYINPUT54), .A2(n1275), .ZN(n1267) );
NAND2_X1 U929 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND3_X1 U930 ( .A1(KEYINPUT4), .A2(n1273), .A3(n1220), .ZN(n1277) );
INV_X1 U931 ( .A(n1270), .ZN(n1273) );
NAND3_X1 U932 ( .A1(n1237), .A2(n1085), .A3(n1239), .ZN(n1270) );
OR2_X1 U933 ( .A1(n1220), .A2(KEYINPUT4), .ZN(n1276) );
XNOR2_X1 U934 ( .A(G137), .B(n1278), .ZN(G39) );
NAND4_X1 U935 ( .A1(n1279), .A2(n1078), .A3(n1280), .A4(n1250), .ZN(n1278) );
XOR2_X1 U936 ( .A(KEYINPUT46), .B(n1100), .Z(n1280) );
XOR2_X1 U937 ( .A(n1149), .B(n1230), .Z(G36) );
NAND3_X1 U938 ( .A1(n1281), .A2(n1086), .A3(n1237), .ZN(n1230) );
INV_X1 U939 ( .A(G134), .ZN(n1149) );
XOR2_X1 U940 ( .A(n1282), .B(G131), .Z(G33) );
NAND2_X1 U941 ( .A1(KEYINPUT41), .A2(n1231), .ZN(n1282) );
NAND3_X1 U942 ( .A1(n1085), .A2(n1281), .A3(n1237), .ZN(n1231) );
AND3_X1 U943 ( .A1(n1100), .A2(n1250), .A3(n1078), .ZN(n1237) );
AND2_X1 U944 ( .A1(n1105), .A2(n1109), .ZN(n1078) );
XNOR2_X1 U945 ( .A(G128), .B(n1154), .ZN(G30) );
NAND3_X1 U946 ( .A1(n1086), .A2(n1260), .A3(n1261), .ZN(n1154) );
INV_X1 U947 ( .A(n1236), .ZN(n1261) );
NAND4_X1 U948 ( .A1(n1100), .A2(n1115), .A3(n1125), .A4(n1250), .ZN(n1236) );
XNOR2_X1 U949 ( .A(n1240), .B(n1283), .ZN(G3) );
NOR2_X1 U950 ( .A1(KEYINPUT5), .A2(n1284), .ZN(n1283) );
NAND3_X1 U951 ( .A1(n1087), .A2(n1242), .A3(n1281), .ZN(n1240) );
INV_X1 U952 ( .A(n1285), .ZN(n1242) );
XOR2_X1 U953 ( .A(n1232), .B(n1286), .Z(G27) );
NAND2_X1 U954 ( .A1(KEYINPUT10), .A2(G125), .ZN(n1286) );
NAND4_X1 U955 ( .A1(n1239), .A2(n1085), .A3(n1287), .A4(n1080), .ZN(n1232) );
NOR2_X1 U956 ( .A1(n1263), .A2(n1102), .ZN(n1287) );
INV_X1 U957 ( .A(n1260), .ZN(n1102) );
INV_X1 U958 ( .A(n1250), .ZN(n1263) );
NAND2_X1 U959 ( .A1(n1106), .A2(n1288), .ZN(n1250) );
NAND4_X1 U960 ( .A1(G953), .A2(G902), .A3(n1289), .A4(n1290), .ZN(n1288) );
INV_X1 U961 ( .A(G900), .ZN(n1290) );
XNOR2_X1 U962 ( .A(G122), .B(n1245), .ZN(G24) );
NAND4_X1 U963 ( .A1(n1291), .A2(n1292), .A3(n1083), .A4(n1264), .ZN(n1245) );
NOR2_X1 U964 ( .A1(n1125), .A2(n1115), .ZN(n1083) );
XNOR2_X1 U965 ( .A(G119), .B(n1293), .ZN(G21) );
NAND2_X1 U966 ( .A1(n1294), .A2(n1260), .ZN(n1293) );
XOR2_X1 U967 ( .A(n1247), .B(KEYINPUT11), .Z(n1294) );
NAND3_X1 U968 ( .A1(n1080), .A2(n1295), .A3(n1279), .ZN(n1247) );
AND3_X1 U969 ( .A1(n1115), .A2(n1125), .A3(n1087), .ZN(n1279) );
INV_X1 U970 ( .A(n1235), .ZN(n1087) );
INV_X1 U971 ( .A(n1296), .ZN(n1115) );
XNOR2_X1 U972 ( .A(G116), .B(n1246), .ZN(G18) );
NAND3_X1 U973 ( .A1(n1292), .A2(n1086), .A3(n1281), .ZN(n1246) );
NOR2_X1 U974 ( .A1(n1291), .A2(n1116), .ZN(n1086) );
XOR2_X1 U975 ( .A(G113), .B(n1297), .Z(G15) );
NOR2_X1 U976 ( .A1(KEYINPUT2), .A2(n1244), .ZN(n1297) );
NAND3_X1 U977 ( .A1(n1281), .A2(n1292), .A3(n1085), .ZN(n1244) );
NOR2_X1 U978 ( .A1(n1266), .A2(n1264), .ZN(n1085) );
INV_X1 U979 ( .A(n1116), .ZN(n1264) );
AND3_X1 U980 ( .A1(n1260), .A2(n1295), .A3(n1080), .ZN(n1292) );
NOR2_X1 U981 ( .A1(n1099), .A2(n1098), .ZN(n1080) );
INV_X1 U982 ( .A(n1298), .ZN(n1099) );
INV_X1 U983 ( .A(n1090), .ZN(n1281) );
NAND2_X1 U984 ( .A1(n1296), .A2(n1125), .ZN(n1090) );
XOR2_X1 U985 ( .A(G110), .B(n1299), .Z(G12) );
NOR4_X1 U986 ( .A1(KEYINPUT18), .A2(n1285), .A3(n1235), .A4(n1089), .ZN(n1299) );
INV_X1 U987 ( .A(n1239), .ZN(n1089) );
NOR2_X1 U988 ( .A1(n1125), .A2(n1296), .ZN(n1239) );
XNOR2_X1 U989 ( .A(n1300), .B(n1184), .ZN(n1296) );
NAND2_X1 U990 ( .A1(G217), .A2(n1301), .ZN(n1184) );
NAND2_X1 U991 ( .A1(n1182), .A2(n1302), .ZN(n1300) );
XNOR2_X1 U992 ( .A(n1303), .B(n1304), .ZN(n1182) );
XOR2_X1 U993 ( .A(n1305), .B(n1306), .Z(n1303) );
XOR2_X1 U994 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U995 ( .A(G125), .B(G119), .Z(n1308) );
XOR2_X1 U996 ( .A(KEYINPUT38), .B(KEYINPUT21), .Z(n1307) );
XOR2_X1 U997 ( .A(n1309), .B(n1310), .Z(n1305) );
XNOR2_X1 U998 ( .A(n1311), .B(n1312), .ZN(n1310) );
NOR2_X1 U999 ( .A1(KEYINPUT16), .A2(n1220), .ZN(n1312) );
NAND2_X1 U1000 ( .A1(KEYINPUT6), .A2(n1145), .ZN(n1311) );
INV_X1 U1001 ( .A(n1313), .ZN(n1145) );
XOR2_X1 U1002 ( .A(n1314), .B(n1315), .Z(n1309) );
AND3_X1 U1003 ( .A1(G221), .A2(n1138), .A3(G234), .ZN(n1315) );
NAND2_X1 U1004 ( .A1(KEYINPUT35), .A2(n1178), .ZN(n1314) );
XNOR2_X1 U1005 ( .A(n1316), .B(G472), .ZN(n1125) );
NAND2_X1 U1006 ( .A1(n1317), .A2(n1302), .ZN(n1316) );
XNOR2_X1 U1007 ( .A(n1202), .B(n1318), .ZN(n1317) );
XOR2_X1 U1008 ( .A(n1284), .B(n1203), .Z(n1318) );
NAND2_X1 U1009 ( .A1(G210), .A2(n1319), .ZN(n1203) );
XNOR2_X1 U1010 ( .A(n1320), .B(n1321), .ZN(n1202) );
XOR2_X1 U1011 ( .A(G113), .B(n1143), .Z(n1321) );
XOR2_X1 U1012 ( .A(n1209), .B(n1322), .Z(n1320) );
NAND2_X1 U1013 ( .A1(n1116), .A2(n1266), .ZN(n1235) );
INV_X1 U1014 ( .A(n1291), .ZN(n1266) );
XOR2_X1 U1015 ( .A(n1323), .B(n1123), .Z(n1291) );
INV_X1 U1016 ( .A(n1120), .ZN(n1123) );
NAND2_X1 U1017 ( .A1(n1324), .A2(n1302), .ZN(n1120) );
INV_X1 U1018 ( .A(n1193), .ZN(n1324) );
XOR2_X1 U1019 ( .A(n1325), .B(n1326), .Z(n1193) );
XOR2_X1 U1020 ( .A(n1327), .B(n1328), .Z(n1326) );
XOR2_X1 U1021 ( .A(G140), .B(G113), .Z(n1328) );
XOR2_X1 U1022 ( .A(G146), .B(G143), .Z(n1327) );
XOR2_X1 U1023 ( .A(n1329), .B(n1330), .Z(n1325) );
XOR2_X1 U1024 ( .A(n1331), .B(n1332), .Z(n1330) );
NOR2_X1 U1025 ( .A1(KEYINPUT40), .A2(n1333), .ZN(n1331) );
INV_X1 U1026 ( .A(G131), .ZN(n1333) );
XOR2_X1 U1027 ( .A(n1334), .B(G104), .Z(n1329) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1319), .ZN(n1334) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1319) );
NAND2_X1 U1030 ( .A1(KEYINPUT49), .A2(n1124), .ZN(n1323) );
INV_X1 U1031 ( .A(G475), .ZN(n1124) );
XNOR2_X1 U1032 ( .A(G478), .B(n1335), .ZN(n1116) );
NOR2_X1 U1033 ( .A1(G902), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1034 ( .A(KEYINPUT22), .B(n1188), .Z(n1336) );
XNOR2_X1 U1035 ( .A(n1337), .B(n1338), .ZN(n1188) );
NOR3_X1 U1036 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(n1338) );
NOR2_X1 U1037 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NOR2_X1 U1038 ( .A1(KEYINPUT19), .A2(n1344), .ZN(n1342) );
XNOR2_X1 U1039 ( .A(KEYINPUT39), .B(n1345), .ZN(n1344) );
NOR3_X1 U1040 ( .A1(n1346), .A2(KEYINPUT19), .A3(n1345), .ZN(n1340) );
INV_X1 U1041 ( .A(n1343), .ZN(n1346) );
XNOR2_X1 U1042 ( .A(G128), .B(n1347), .ZN(n1343) );
XOR2_X1 U1043 ( .A(G143), .B(G134), .Z(n1347) );
AND2_X1 U1044 ( .A1(n1345), .A2(KEYINPUT19), .ZN(n1339) );
XNOR2_X1 U1045 ( .A(G107), .B(n1348), .ZN(n1345) );
XOR2_X1 U1046 ( .A(G122), .B(G116), .Z(n1348) );
NAND4_X1 U1047 ( .A1(KEYINPUT45), .A2(G234), .A3(G217), .A4(n1138), .ZN(n1337) );
NAND3_X1 U1048 ( .A1(n1100), .A2(n1295), .A3(n1260), .ZN(n1285) );
NOR2_X1 U1049 ( .A1(n1105), .A2(n1104), .ZN(n1260) );
INV_X1 U1050 ( .A(n1109), .ZN(n1104) );
NAND2_X1 U1051 ( .A1(G214), .A2(n1349), .ZN(n1109) );
XOR2_X1 U1052 ( .A(n1130), .B(n1350), .Z(n1105) );
NOR2_X1 U1053 ( .A1(n1128), .A2(KEYINPUT53), .ZN(n1350) );
INV_X1 U1054 ( .A(n1224), .ZN(n1128) );
NAND2_X1 U1055 ( .A1(G210), .A2(n1349), .ZN(n1224) );
NAND2_X1 U1056 ( .A1(n1351), .A2(n1302), .ZN(n1349) );
INV_X1 U1057 ( .A(G237), .ZN(n1351) );
AND2_X1 U1058 ( .A1(n1352), .A2(n1302), .ZN(n1130) );
XOR2_X1 U1059 ( .A(n1258), .B(n1353), .Z(n1352) );
XOR2_X1 U1060 ( .A(n1256), .B(n1332), .Z(n1353) );
XOR2_X1 U1061 ( .A(G122), .B(G125), .Z(n1332) );
XNOR2_X1 U1062 ( .A(n1354), .B(n1143), .ZN(n1256) );
NAND2_X1 U1063 ( .A1(G224), .A2(n1138), .ZN(n1354) );
XOR2_X1 U1064 ( .A(n1176), .B(n1178), .Z(n1258) );
INV_X1 U1065 ( .A(G110), .ZN(n1178) );
NAND2_X1 U1066 ( .A1(n1355), .A2(n1356), .ZN(n1176) );
NAND2_X1 U1067 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
INV_X1 U1068 ( .A(n1174), .ZN(n1355) );
NOR2_X1 U1069 ( .A1(n1358), .A2(n1357), .ZN(n1174) );
XNOR2_X1 U1070 ( .A(G101), .B(n1359), .ZN(n1357) );
NOR2_X1 U1071 ( .A1(KEYINPUT13), .A2(n1360), .ZN(n1359) );
XOR2_X1 U1072 ( .A(G104), .B(n1361), .Z(n1360) );
NOR2_X1 U1073 ( .A1(G107), .A2(KEYINPUT12), .ZN(n1361) );
NAND2_X1 U1074 ( .A1(n1362), .A2(n1363), .ZN(n1358) );
NAND2_X1 U1075 ( .A1(n1364), .A2(n1365), .ZN(n1363) );
INV_X1 U1076 ( .A(G113), .ZN(n1365) );
NAND2_X1 U1077 ( .A1(n1366), .A2(n1367), .ZN(n1364) );
NAND2_X1 U1078 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
NAND2_X1 U1079 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1080 ( .A1(n1322), .A2(n1370), .ZN(n1366) );
XOR2_X1 U1081 ( .A(KEYINPUT48), .B(KEYINPUT1), .Z(n1370) );
INV_X1 U1082 ( .A(n1368), .ZN(n1322) );
NAND3_X1 U1083 ( .A1(n1368), .A2(n1371), .A3(G113), .ZN(n1362) );
INV_X1 U1084 ( .A(KEYINPUT63), .ZN(n1371) );
XOR2_X1 U1085 ( .A(G116), .B(G119), .Z(n1368) );
NAND2_X1 U1086 ( .A1(n1106), .A2(n1372), .ZN(n1295) );
NAND4_X1 U1087 ( .A1(G953), .A2(G902), .A3(n1289), .A4(n1373), .ZN(n1372) );
INV_X1 U1088 ( .A(G898), .ZN(n1373) );
NAND3_X1 U1089 ( .A1(n1073), .A2(n1289), .A3(G952), .ZN(n1106) );
NAND2_X1 U1090 ( .A1(G237), .A2(G234), .ZN(n1289) );
XOR2_X1 U1091 ( .A(n1138), .B(KEYINPUT59), .Z(n1073) );
NOR2_X1 U1092 ( .A1(n1298), .A2(n1098), .ZN(n1100) );
AND2_X1 U1093 ( .A1(G221), .A2(n1301), .ZN(n1098) );
NAND2_X1 U1094 ( .A1(G234), .A2(n1302), .ZN(n1301) );
INV_X1 U1095 ( .A(G902), .ZN(n1302) );
NOR2_X1 U1096 ( .A1(n1374), .A2(n1127), .ZN(n1298) );
NOR3_X1 U1097 ( .A1(G469), .A2(G902), .A3(n1375), .ZN(n1127) );
XNOR2_X1 U1098 ( .A(KEYINPUT8), .B(n1126), .ZN(n1374) );
AND2_X1 U1099 ( .A1(G469), .A2(n1376), .ZN(n1126) );
OR2_X1 U1100 ( .A1(n1375), .A2(G902), .ZN(n1376) );
XOR2_X1 U1101 ( .A(n1377), .B(n1378), .Z(n1375) );
XNOR2_X1 U1102 ( .A(n1209), .B(n1379), .ZN(n1378) );
XNOR2_X1 U1103 ( .A(n1143), .B(n1380), .ZN(n1379) );
NOR2_X1 U1104 ( .A1(KEYINPUT23), .A2(n1210), .ZN(n1380) );
XNOR2_X1 U1105 ( .A(n1381), .B(n1382), .ZN(n1210) );
XOR2_X1 U1106 ( .A(KEYINPUT34), .B(G107), .Z(n1382) );
XOR2_X1 U1107 ( .A(n1284), .B(G104), .Z(n1381) );
INV_X1 U1108 ( .A(G101), .ZN(n1284) );
XOR2_X1 U1109 ( .A(G143), .B(n1304), .Z(n1143) );
XOR2_X1 U1110 ( .A(G128), .B(G146), .Z(n1304) );
XNOR2_X1 U1111 ( .A(n1383), .B(n1384), .ZN(n1209) );
XOR2_X1 U1112 ( .A(G134), .B(G131), .Z(n1384) );
NAND2_X1 U1113 ( .A1(KEYINPUT9), .A2(n1313), .ZN(n1383) );
XNOR2_X1 U1114 ( .A(G137), .B(KEYINPUT14), .ZN(n1313) );
XOR2_X1 U1115 ( .A(n1385), .B(n1386), .Z(n1377) );
XNOR2_X1 U1116 ( .A(n1387), .B(n1218), .ZN(n1386) );
NAND2_X1 U1117 ( .A1(G227), .A2(n1138), .ZN(n1218) );
INV_X1 U1118 ( .A(G953), .ZN(n1138) );
NOR2_X1 U1119 ( .A1(G110), .A2(KEYINPUT43), .ZN(n1387) );
XOR2_X1 U1120 ( .A(n1220), .B(KEYINPUT27), .Z(n1385) );
INV_X1 U1121 ( .A(G140), .ZN(n1220) );
endmodule


