//Key = 0000011101001001111101111000011110101100100100101100001101000011


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
n2292, n2293, n2294;

OR2_X1 U1287 ( .A1(n2294), .A2(n1723), .ZN(U280) );
OR2_X1 U1288 ( .A1(n1753), .A2(STATO_REG_0__SCAN_IN), .ZN(n1722) );
INV_X2 U1289 ( .A(n1722), .ZN(n1723) );
INV_X2 U1290 ( .A(U280), .ZN(n1724) );
INV_X1 U1291 ( .A(n1725), .ZN(U375) );
NAND2_X1 U1292 ( .A1(n1726), .A2(n1727), .ZN(U344) );
NAND2_X1 U1293 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1728), .ZN(n1727) );
NAND2_X1 U1294 ( .A1(DATA_IN_7_), .A2(n1729), .ZN(n1726) );
NAND2_X1 U1295 ( .A1(n1730), .A2(n1731), .ZN(U343) );
NAND2_X1 U1296 ( .A1(n1732), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1731) );
XOR2_X1 U1297 ( .A(n1728), .B(KEYINPUT42), .Z(n1732) );
NAND2_X1 U1298 ( .A1(DATA_IN_6_), .A2(n1729), .ZN(n1730) );
NAND2_X1 U1299 ( .A1(n1733), .A2(n1734), .ZN(U342) );
NAND2_X1 U1300 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1728), .ZN(n1734) );
NAND2_X1 U1301 ( .A1(DATA_IN_5_), .A2(n1729), .ZN(n1733) );
NAND2_X1 U1302 ( .A1(n1735), .A2(n1736), .ZN(U341) );
NAND2_X1 U1303 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1728), .ZN(n1736) );
NAND2_X1 U1304 ( .A1(DATA_IN_4_), .A2(n1729), .ZN(n1735) );
NAND2_X1 U1305 ( .A1(n1737), .A2(n1738), .ZN(U340) );
NAND2_X1 U1306 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1728), .ZN(n1738) );
NAND2_X1 U1307 ( .A1(DATA_IN_3_), .A2(n1729), .ZN(n1737) );
NAND2_X1 U1308 ( .A1(n1739), .A2(n1740), .ZN(U339) );
NAND2_X1 U1309 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1728), .ZN(n1740) );
NAND2_X1 U1310 ( .A1(DATA_IN_2_), .A2(n1729), .ZN(n1739) );
NAND2_X1 U1311 ( .A1(n1741), .A2(n1742), .ZN(U338) );
NAND2_X1 U1312 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1728), .ZN(n1742) );
NAND2_X1 U1313 ( .A1(DATA_IN_1_), .A2(n1729), .ZN(n1741) );
NAND2_X1 U1314 ( .A1(n1743), .A2(n1744), .ZN(U337) );
NAND2_X1 U1315 ( .A1(n1745), .A2(n1728), .ZN(n1744) );
NAND2_X1 U1316 ( .A1(n1725), .A2(n1746), .ZN(n1728) );
NAND2_X1 U1317 ( .A1(n1747), .A2(n1748), .ZN(n1746) );
XOR2_X1 U1318 ( .A(n1749), .B(KEYINPUT30), .Z(n1745) );
NAND2_X1 U1319 ( .A1(DATA_IN_0_), .A2(n1729), .ZN(n1743) );
NAND2_X1 U1320 ( .A1(n1748), .A2(n1750), .ZN(n1729) );
NAND2_X1 U1321 ( .A1(n1751), .A2(n1752), .ZN(n1750) );
XOR2_X1 U1322 ( .A(n1753), .B(KEYINPUT40), .Z(n1751) );
NAND2_X1 U1323 ( .A1(n1754), .A2(n1755), .ZN(U336) );
NAND2_X1 U1324 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1756), .ZN(n1755) );
NAND2_X1 U1325 ( .A1(n1757), .A2(DATA_IN_7_), .ZN(n1754) );
NAND2_X1 U1326 ( .A1(n1758), .A2(n1759), .ZN(U335) );
NAND2_X1 U1327 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1756), .ZN(n1759) );
NAND2_X1 U1328 ( .A1(n1757), .A2(DATA_IN_6_), .ZN(n1758) );
NAND2_X1 U1329 ( .A1(n1760), .A2(n1761), .ZN(U334) );
NAND2_X1 U1330 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1756), .ZN(n1761) );
NAND2_X1 U1331 ( .A1(n1757), .A2(DATA_IN_5_), .ZN(n1760) );
NAND2_X1 U1332 ( .A1(n1762), .A2(n1763), .ZN(U333) );
NAND2_X1 U1333 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1756), .ZN(n1763) );
NAND2_X1 U1334 ( .A1(n1757), .A2(DATA_IN_4_), .ZN(n1762) );
NAND2_X1 U1335 ( .A1(n1764), .A2(n1765), .ZN(U332) );
NAND2_X1 U1336 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1756), .ZN(n1765) );
NAND2_X1 U1337 ( .A1(n1757), .A2(DATA_IN_3_), .ZN(n1764) );
NAND2_X1 U1338 ( .A1(n1766), .A2(n1767), .ZN(U331) );
NAND2_X1 U1339 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1756), .ZN(n1767) );
NAND2_X1 U1340 ( .A1(n1757), .A2(DATA_IN_2_), .ZN(n1766) );
NAND2_X1 U1341 ( .A1(n1768), .A2(n1769), .ZN(U330) );
NAND2_X1 U1342 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1756), .ZN(n1769) );
NAND2_X1 U1343 ( .A1(n1757), .A2(DATA_IN_1_), .ZN(n1768) );
NAND2_X1 U1344 ( .A1(n1770), .A2(n1771), .ZN(U329) );
NAND2_X1 U1345 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1756), .ZN(n1771) );
NAND2_X1 U1346 ( .A1(n1757), .A2(DATA_IN_0_), .ZN(n1770) );
INV_X1 U1347 ( .A(n1756), .ZN(n1757) );
NAND2_X1 U1348 ( .A1(n1725), .A2(n1772), .ZN(n1756) );
NAND2_X1 U1349 ( .A1(n1773), .A2(n1748), .ZN(n1772) );
NAND2_X1 U1350 ( .A1(n1747), .A2(n1774), .ZN(n1773) );
NAND2_X1 U1351 ( .A1(n1775), .A2(n1776), .ZN(n1774) );
NAND3_X1 U1352 ( .A1(n1777), .A2(n1778), .A3(n1779), .ZN(n1776) );
NAND2_X1 U1353 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1780), .ZN(n1779) );
NAND3_X1 U1354 ( .A1(n1781), .A2(n1782), .A3(n1783), .ZN(n1778) );
NAND2_X1 U1355 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1784), .ZN(n1783) );
NAND3_X1 U1356 ( .A1(n1785), .A2(n1786), .A3(n1787), .ZN(n1782) );
NAND2_X1 U1357 ( .A1(DATA_IN_5_), .A2(n1788), .ZN(n1787) );
NAND3_X1 U1358 ( .A1(n1789), .A2(n1790), .A3(n1791), .ZN(n1786) );
XOR2_X1 U1359 ( .A(KEYINPUT62), .B(n1792), .Z(n1791) );
NOR2_X1 U1360 ( .A1(DATA_IN_3_), .A2(n1793), .ZN(n1792) );
NAND3_X1 U1361 ( .A1(n1794), .A2(n1795), .A3(n1796), .ZN(n1790) );
NAND2_X1 U1362 ( .A1(DATA_IN_3_), .A2(n1793), .ZN(n1796) );
NAND3_X1 U1363 ( .A1(n1797), .A2(n1798), .A3(n1799), .ZN(n1795) );
NAND2_X1 U1364 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1800), .ZN(n1799) );
NAND3_X1 U1365 ( .A1(n1801), .A2(n1802), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1798) );
XOR2_X1 U1366 ( .A(KEYINPUT17), .B(n1803), .Z(n1801) );
NOR2_X1 U1367 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1804), .ZN(n1803) );
NAND2_X1 U1368 ( .A1(n1805), .A2(n1804), .ZN(n1797) );
XOR2_X1 U1369 ( .A(RMIN_REG_1__SCAN_IN), .B(KEYINPUT33), .Z(n1805) );
NAND2_X1 U1370 ( .A1(DATA_IN_2_), .A2(n1806), .ZN(n1794) );
NAND2_X1 U1371 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1807), .ZN(n1789) );
NAND2_X1 U1372 ( .A1(DATA_IN_4_), .A2(n1808), .ZN(n1785) );
NAND2_X1 U1373 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1809), .ZN(n1781) );
OR2_X1 U1374 ( .A1(n1784), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1777) );
NAND2_X1 U1375 ( .A1(DATA_IN_7_), .A2(n1810), .ZN(n1775) );
INV_X1 U1376 ( .A(n1752), .ZN(n1747) );
NAND2_X1 U1377 ( .A1(n1811), .A2(n1812), .ZN(n1752) );
NAND2_X1 U1378 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1780), .ZN(n1812) );
NAND3_X1 U1379 ( .A1(n1813), .A2(n1814), .A3(n1815), .ZN(n1811) );
NAND2_X1 U1380 ( .A1(DATA_IN_7_), .A2(n1816), .ZN(n1815) );
NAND3_X1 U1381 ( .A1(n1817), .A2(n1818), .A3(n1819), .ZN(n1814) );
NAND2_X1 U1382 ( .A1(DATA_IN_6_), .A2(n1820), .ZN(n1819) );
NAND3_X1 U1383 ( .A1(n1821), .A2(n1822), .A3(n1823), .ZN(n1818) );
NAND2_X1 U1384 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1809), .ZN(n1823) );
NAND3_X1 U1385 ( .A1(n1824), .A2(n1825), .A3(n1826), .ZN(n1822) );
NAND2_X1 U1386 ( .A1(DATA_IN_4_), .A2(n1827), .ZN(n1826) );
NAND3_X1 U1387 ( .A1(n1828), .A2(n1829), .A3(n1830), .ZN(n1825) );
NAND2_X1 U1388 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1831), .ZN(n1830) );
NAND3_X1 U1389 ( .A1(n1832), .A2(n1833), .A3(n1834), .ZN(n1829) );
XOR2_X1 U1390 ( .A(n1835), .B(KEYINPUT52), .Z(n1834) );
NAND2_X1 U1391 ( .A1(DATA_IN_2_), .A2(n1836), .ZN(n1835) );
NAND3_X1 U1392 ( .A1(n1837), .A2(n1749), .A3(DATA_IN_0_), .ZN(n1833) );
NAND2_X1 U1393 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1804), .ZN(n1837) );
NAND2_X1 U1394 ( .A1(DATA_IN_1_), .A2(n1838), .ZN(n1832) );
NAND2_X1 U1395 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1800), .ZN(n1828) );
NAND2_X1 U1396 ( .A1(DATA_IN_3_), .A2(n1839), .ZN(n1824) );
NAND2_X1 U1397 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1807), .ZN(n1821) );
NAND2_X1 U1398 ( .A1(n1840), .A2(n1841), .ZN(n1817) );
INV_X1 U1399 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1841) );
XOR2_X1 U1400 ( .A(n1809), .B(KEYINPUT24), .Z(n1840) );
NAND2_X1 U1401 ( .A1(n1842), .A2(RMAX_REG_6__SCAN_IN), .ZN(n1813) );
XOR2_X1 U1402 ( .A(n1784), .B(KEYINPUT0), .Z(n1842) );
NAND2_X1 U1403 ( .A1(n1843), .A2(n1844), .ZN(U328) );
NAND2_X1 U1404 ( .A1(n1845), .A2(DATA_IN_7_), .ZN(n1844) );
NAND2_X1 U1405 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1846), .ZN(n1843) );
NAND2_X1 U1406 ( .A1(n1847), .A2(n1848), .ZN(U327) );
NAND2_X1 U1407 ( .A1(n1845), .A2(DATA_IN_6_), .ZN(n1848) );
NAND2_X1 U1408 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1846), .ZN(n1847) );
NAND2_X1 U1409 ( .A1(n1849), .A2(n1850), .ZN(U326) );
NAND2_X1 U1410 ( .A1(n1845), .A2(DATA_IN_5_), .ZN(n1850) );
NAND2_X1 U1411 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1846), .ZN(n1849) );
NAND2_X1 U1412 ( .A1(n1851), .A2(n1852), .ZN(U325) );
NAND2_X1 U1413 ( .A1(n1845), .A2(DATA_IN_4_), .ZN(n1852) );
NAND2_X1 U1414 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1846), .ZN(n1851) );
NAND2_X1 U1415 ( .A1(n1853), .A2(n1854), .ZN(U324) );
NAND2_X1 U1416 ( .A1(n1845), .A2(DATA_IN_3_), .ZN(n1854) );
NAND2_X1 U1417 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1846), .ZN(n1853) );
NAND2_X1 U1418 ( .A1(n1855), .A2(n1856), .ZN(U323) );
NAND2_X1 U1419 ( .A1(n1857), .A2(n1845), .ZN(n1856) );
XOR2_X1 U1420 ( .A(n1800), .B(KEYINPUT34), .Z(n1857) );
NAND2_X1 U1421 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1846), .ZN(n1855) );
NAND2_X1 U1422 ( .A1(n1858), .A2(n1859), .ZN(U322) );
NAND2_X1 U1423 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1846), .ZN(n1859) );
XOR2_X1 U1424 ( .A(KEYINPUT46), .B(n1860), .Z(n1858) );
NOR2_X1 U1425 ( .A1(n1804), .A2(n1861), .ZN(n1860) );
NAND2_X1 U1426 ( .A1(n1862), .A2(n1863), .ZN(U321) );
NAND2_X1 U1427 ( .A1(n1845), .A2(DATA_IN_0_), .ZN(n1863) );
INV_X1 U1428 ( .A(n1861), .ZN(n1845) );
NAND2_X1 U1429 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1864), .ZN(n1861) );
NAND2_X1 U1430 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1846), .ZN(n1862) );
NAND2_X1 U1431 ( .A1(n1725), .A2(n1864), .ZN(n1846) );
NAND2_X1 U1432 ( .A1(n1865), .A2(n1748), .ZN(n1864) );
NAND2_X1 U1433 ( .A1(n1748), .A2(n1753), .ZN(n1725) );
NAND2_X1 U1434 ( .A1(n1866), .A2(n1867), .ZN(U320) );
NAND2_X1 U1435 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1724), .ZN(n1867) );
NAND2_X1 U1436 ( .A1(n1723), .A2(DATA_IN_7_), .ZN(n1866) );
NAND2_X1 U1437 ( .A1(n1868), .A2(n1869), .ZN(U319) );
NAND2_X1 U1438 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1724), .ZN(n1869) );
NAND2_X1 U1439 ( .A1(n1723), .A2(DATA_IN_6_), .ZN(n1868) );
NAND2_X1 U1440 ( .A1(n1870), .A2(n1871), .ZN(U318) );
NAND2_X1 U1441 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1724), .ZN(n1871) );
NAND2_X1 U1442 ( .A1(n1723), .A2(DATA_IN_5_), .ZN(n1870) );
NAND2_X1 U1443 ( .A1(n1872), .A2(n1873), .ZN(U317) );
NAND2_X1 U1444 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1724), .ZN(n1873) );
NAND2_X1 U1445 ( .A1(n1723), .A2(DATA_IN_4_), .ZN(n1872) );
NAND2_X1 U1446 ( .A1(n1874), .A2(n1875), .ZN(U316) );
NAND2_X1 U1447 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1724), .ZN(n1875) );
NAND2_X1 U1448 ( .A1(n1723), .A2(DATA_IN_3_), .ZN(n1874) );
NAND2_X1 U1449 ( .A1(n1876), .A2(n1877), .ZN(U315) );
NAND2_X1 U1450 ( .A1(n1878), .A2(n1724), .ZN(n1877) );
XNOR2_X1 U1451 ( .A(REG1_REG_2__SCAN_IN), .B(KEYINPUT12), .ZN(n1878) );
NAND2_X1 U1452 ( .A1(n1723), .A2(DATA_IN_2_), .ZN(n1876) );
NAND2_X1 U1453 ( .A1(n1879), .A2(n1880), .ZN(U314) );
NAND2_X1 U1454 ( .A1(n1723), .A2(DATA_IN_1_), .ZN(n1880) );
XOR2_X1 U1455 ( .A(n1881), .B(KEYINPUT41), .Z(n1879) );
NAND2_X1 U1456 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1724), .ZN(n1881) );
NAND2_X1 U1457 ( .A1(n1882), .A2(n1883), .ZN(U313) );
NAND2_X1 U1458 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1724), .ZN(n1883) );
NAND2_X1 U1459 ( .A1(n1723), .A2(DATA_IN_0_), .ZN(n1882) );
NAND2_X1 U1460 ( .A1(n1884), .A2(n1885), .ZN(U312) );
NAND2_X1 U1461 ( .A1(n1886), .A2(REG2_REG_7__SCAN_IN), .ZN(n1885) );
XOR2_X1 U1462 ( .A(U280), .B(KEYINPUT5), .Z(n1886) );
NAND2_X1 U1463 ( .A1(n1723), .A2(REG1_REG_7__SCAN_IN), .ZN(n1884) );
NAND2_X1 U1464 ( .A1(n1887), .A2(n1888), .ZN(U311) );
NAND2_X1 U1465 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1724), .ZN(n1888) );
NAND2_X1 U1466 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1723), .ZN(n1887) );
NAND2_X1 U1467 ( .A1(n1889), .A2(n1890), .ZN(U310) );
NAND2_X1 U1468 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1724), .ZN(n1890) );
XOR2_X1 U1469 ( .A(n1891), .B(KEYINPUT4), .Z(n1889) );
NAND2_X1 U1470 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1723), .ZN(n1891) );
NAND2_X1 U1471 ( .A1(n1892), .A2(n1893), .ZN(U309) );
NAND2_X1 U1472 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1724), .ZN(n1893) );
NAND2_X1 U1473 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1723), .ZN(n1892) );
NAND2_X1 U1474 ( .A1(n1894), .A2(n1895), .ZN(U308) );
NAND2_X1 U1475 ( .A1(n1896), .A2(n1724), .ZN(n1895) );
XOR2_X1 U1476 ( .A(REG2_REG_3__SCAN_IN), .B(KEYINPUT45), .Z(n1896) );
NAND2_X1 U1477 ( .A1(n1723), .A2(n1897), .ZN(n1894) );
XOR2_X1 U1478 ( .A(REG1_REG_3__SCAN_IN), .B(KEYINPUT61), .Z(n1897) );
NAND2_X1 U1479 ( .A1(n1898), .A2(n1899), .ZN(U307) );
NAND2_X1 U1480 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1724), .ZN(n1899) );
XOR2_X1 U1481 ( .A(n1900), .B(KEYINPUT56), .Z(n1898) );
NAND2_X1 U1482 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1723), .ZN(n1900) );
NAND2_X1 U1483 ( .A1(n1901), .A2(n1902), .ZN(U306) );
NAND2_X1 U1484 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1724), .ZN(n1902) );
NAND2_X1 U1485 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1723), .ZN(n1901) );
NAND2_X1 U1486 ( .A1(n1903), .A2(n1904), .ZN(U305) );
NAND2_X1 U1487 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1724), .ZN(n1904) );
NAND2_X1 U1488 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1723), .ZN(n1903) );
NAND2_X1 U1489 ( .A1(n1905), .A2(n1906), .ZN(U304) );
NAND2_X1 U1490 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1724), .ZN(n1906) );
NAND2_X1 U1491 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1723), .ZN(n1905) );
NAND2_X1 U1492 ( .A1(n1907), .A2(n1908), .ZN(U303) );
NAND2_X1 U1493 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1724), .ZN(n1908) );
NAND2_X1 U1494 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1723), .ZN(n1907) );
NAND2_X1 U1495 ( .A1(n1909), .A2(n1910), .ZN(U302) );
NAND2_X1 U1496 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1724), .ZN(n1910) );
XOR2_X1 U1497 ( .A(n1911), .B(KEYINPUT11), .Z(n1909) );
NAND2_X1 U1498 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1723), .ZN(n1911) );
NAND2_X1 U1499 ( .A1(n1912), .A2(n1913), .ZN(U301) );
NAND2_X1 U1500 ( .A1(n1914), .A2(n1724), .ZN(n1913) );
XNOR2_X1 U1501 ( .A(REG3_REG_4__SCAN_IN), .B(KEYINPUT43), .ZN(n1914) );
NAND2_X1 U1502 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1723), .ZN(n1912) );
NAND2_X1 U1503 ( .A1(n1915), .A2(n1916), .ZN(U300) );
NAND2_X1 U1504 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1724), .ZN(n1916) );
XOR2_X1 U1505 ( .A(KEYINPUT37), .B(n1917), .Z(n1915) );
AND2_X1 U1506 ( .A1(n1723), .A2(REG2_REG_3__SCAN_IN), .ZN(n1917) );
NAND2_X1 U1507 ( .A1(n1918), .A2(n1919), .ZN(U299) );
NAND2_X1 U1508 ( .A1(n1723), .A2(n1920), .ZN(n1919) );
XOR2_X1 U1509 ( .A(REG2_REG_2__SCAN_IN), .B(KEYINPUT20), .Z(n1920) );
NAND2_X1 U1510 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1724), .ZN(n1918) );
NAND2_X1 U1511 ( .A1(n1921), .A2(n1922), .ZN(U298) );
NAND2_X1 U1512 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1724), .ZN(n1922) );
NAND2_X1 U1513 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1723), .ZN(n1921) );
NAND2_X1 U1514 ( .A1(n1923), .A2(n1924), .ZN(U297) );
NAND2_X1 U1515 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1724), .ZN(n1924) );
NAND2_X1 U1516 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1723), .ZN(n1923) );
NAND2_X1 U1517 ( .A1(n1925), .A2(n1926), .ZN(U296) );
NAND2_X1 U1518 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1724), .ZN(n1926) );
NAND2_X1 U1519 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1723), .ZN(n1925) );
NAND2_X1 U1520 ( .A1(n1927), .A2(n1928), .ZN(U295) );
NAND2_X1 U1521 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1724), .ZN(n1928) );
NAND2_X1 U1522 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1723), .ZN(n1927) );
NAND2_X1 U1523 ( .A1(n1929), .A2(n1930), .ZN(U294) );
NAND2_X1 U1524 ( .A1(n1931), .A2(n1724), .ZN(n1930) );
XOR2_X1 U1525 ( .A(n1932), .B(KEYINPUT48), .Z(n1931) );
NAND2_X1 U1526 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1723), .ZN(n1929) );
NAND2_X1 U1527 ( .A1(n1933), .A2(n1934), .ZN(U293) );
NAND2_X1 U1528 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1724), .ZN(n1934) );
NAND2_X1 U1529 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1723), .ZN(n1933) );
NAND2_X1 U1530 ( .A1(n1935), .A2(n1936), .ZN(U292) );
NAND2_X1 U1531 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1724), .ZN(n1936) );
NAND2_X1 U1532 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1723), .ZN(n1935) );
NAND2_X1 U1533 ( .A1(n1937), .A2(n1938), .ZN(U291) );
NAND2_X1 U1534 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1724), .ZN(n1938) );
NAND2_X1 U1535 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1723), .ZN(n1937) );
NAND2_X1 U1536 ( .A1(n1939), .A2(n1940), .ZN(U290) );
NAND2_X1 U1537 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1724), .ZN(n1940) );
NAND2_X1 U1538 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1723), .ZN(n1939) );
NAND2_X1 U1539 ( .A1(n1941), .A2(n1942), .ZN(U289) );
NAND2_X1 U1540 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1724), .ZN(n1942) );
NAND2_X1 U1541 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1723), .ZN(n1941) );
NAND4_X1 U1542 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .ZN(U288));
NAND2_X1 U1543 ( .A1(n1947), .A2(REG4_REG_7__SCAN_IN), .ZN(n1946) );
NOR2_X1 U1544 ( .A1(n1948), .A2(n1949), .ZN(n1945) );
AND2_X1 U1545 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1950), .ZN(n1949) );
AND4_X1 U1546 ( .A1(n1951), .A2(n1952), .A3(n1953), .A4(KEYINPUT8), .ZN(n1948) );
NAND2_X1 U1547 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1724), .ZN(n1944) );
NAND2_X1 U1548 ( .A1(n1954), .A2(n1955), .ZN(U287) );
NAND2_X1 U1549 ( .A1(n1947), .A2(REG4_REG_6__SCAN_IN), .ZN(n1955) );
XOR2_X1 U1550 ( .A(n1956), .B(KEYINPUT31), .Z(n1954) );
NAND3_X1 U1551 ( .A1(n1943), .A2(n1957), .A3(n1958), .ZN(n1956) );
NOR3_X1 U1552 ( .A1(n1959), .A2(n1960), .A3(n1961), .ZN(n1958) );
NOR3_X1 U1553 ( .A1(n1962), .A2(n1963), .A3(n1964), .ZN(n1961) );
NOR3_X1 U1554 ( .A1(n1965), .A2(n1966), .A3(n1967), .ZN(n1960) );
AND2_X1 U1555 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1950), .ZN(n1959) );
NAND2_X1 U1556 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1724), .ZN(n1957) );
AND2_X1 U1557 ( .A1(n1968), .A2(n1969), .ZN(n1943) );
NAND3_X1 U1558 ( .A1(n1952), .A2(n1965), .A3(n1966), .ZN(n1969) );
NOR3_X1 U1559 ( .A1(n1970), .A2(KEYINPUT8), .A3(n1971), .ZN(n1966) );
NAND3_X1 U1560 ( .A1(n1963), .A2(n1962), .A3(n1972), .ZN(n1968) );
NAND2_X1 U1561 ( .A1(n1973), .A2(n1974), .ZN(n1962) );
XOR2_X1 U1562 ( .A(n1975), .B(KEYINPUT9), .Z(n1973) );
INV_X1 U1563 ( .A(n1976), .ZN(n1963) );
NAND4_X1 U1564 ( .A1(n1977), .A2(n1978), .A3(n1979), .A4(n1980), .ZN(U286));
NOR3_X1 U1565 ( .A1(n1981), .A2(n1982), .A3(n1983), .ZN(n1980) );
NOR2_X1 U1566 ( .A1(n1984), .A2(n1964), .ZN(n1983) );
XOR2_X1 U1567 ( .A(n1985), .B(n1986), .Z(n1984) );
NAND2_X1 U1568 ( .A1(KEYINPUT9), .A2(n1974), .ZN(n1985) );
NAND2_X1 U1569 ( .A1(n1987), .A2(n1976), .ZN(n1974) );
NAND3_X1 U1570 ( .A1(n1988), .A2(n1951), .A3(n1989), .ZN(n1976) );
NAND2_X1 U1571 ( .A1(n1970), .A2(n1990), .ZN(n1987) );
NAND2_X1 U1572 ( .A1(n1989), .A2(n1988), .ZN(n1990) );
NOR3_X1 U1573 ( .A1(n1967), .A2(n1953), .A3(n1991), .ZN(n1982) );
NOR2_X1 U1574 ( .A1(n1992), .A2(n1993), .ZN(n1991) );
INV_X1 U1575 ( .A(n1965), .ZN(n1953) );
NAND2_X1 U1576 ( .A1(n1992), .A2(n1993), .ZN(n1965) );
XOR2_X1 U1577 ( .A(n1970), .B(n1994), .Z(n1993) );
INV_X1 U1578 ( .A(n1951), .ZN(n1970) );
NOR2_X1 U1579 ( .A1(n1951), .A2(n1995), .ZN(n1981) );
NAND2_X1 U1580 ( .A1(n1996), .A2(n1997), .ZN(n1951) );
NAND4_X1 U1581 ( .A1(n1998), .A2(n1999), .A3(n2000), .A4(n2001), .ZN(n1997));
NAND2_X1 U1582 ( .A1(n2002), .A2(n2003), .ZN(n2001) );
XOR2_X1 U1583 ( .A(REG4_REG_6__SCAN_IN), .B(DATA_IN_6_), .Z(n2002) );
NAND2_X1 U1584 ( .A1(n2004), .A2(RESTART), .ZN(n2000) );
XOR2_X1 U1585 ( .A(RMIN_REG_6__SCAN_IN), .B(RMAX_REG_6__SCAN_IN), .Z(n2004));
NAND2_X1 U1586 ( .A1(n2005), .A2(n2006), .ZN(n1999) );
NAND2_X1 U1587 ( .A1(n2007), .A2(n2008), .ZN(n2006) );
XOR2_X1 U1588 ( .A(KEYINPUT39), .B(n2009), .Z(n2008) );
NAND2_X1 U1589 ( .A1(n2010), .A2(n2011), .ZN(n1998) );
NAND4_X1 U1590 ( .A1(n2012), .A2(n2013), .A3(n2014), .A4(n2015), .ZN(n1996));
NAND2_X1 U1591 ( .A1(n2016), .A2(n2003), .ZN(n2015) );
XOR2_X1 U1592 ( .A(REG4_REG_6__SCAN_IN), .B(n1784), .Z(n2016) );
NAND2_X1 U1593 ( .A1(n2017), .A2(RESTART), .ZN(n2014) );
XOR2_X1 U1594 ( .A(n1820), .B(RMIN_REG_6__SCAN_IN), .Z(n2017) );
NAND2_X1 U1595 ( .A1(n2009), .A2(n2018), .ZN(n2013) );
NAND2_X1 U1596 ( .A1(n2005), .A2(n2010), .ZN(n2018) );
NAND2_X1 U1597 ( .A1(n2007), .A2(n2019), .ZN(n2012) );
NAND2_X1 U1598 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1724), .ZN(n1979) );
NAND2_X1 U1599 ( .A1(n1950), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1978) );
NAND2_X1 U1600 ( .A1(n1947), .A2(REG4_REG_5__SCAN_IN), .ZN(n1977) );
NAND4_X1 U1601 ( .A1(n2020), .A2(n2021), .A3(n2022), .A4(n2023), .ZN(U285));
NOR3_X1 U1602 ( .A1(n2024), .A2(n2025), .A3(n2026), .ZN(n2023) );
NOR3_X1 U1603 ( .A1(n1964), .A2(n1986), .A3(n2027), .ZN(n2026) );
NOR2_X1 U1604 ( .A1(n2028), .A2(n2029), .ZN(n2027) );
INV_X1 U1605 ( .A(n1975), .ZN(n1986) );
NAND2_X1 U1606 ( .A1(n2028), .A2(n2029), .ZN(n1975) );
XOR2_X1 U1607 ( .A(n2030), .B(n1989), .Z(n2029) );
INV_X1 U1608 ( .A(n2031), .ZN(n1989) );
NOR3_X1 U1609 ( .A1(n1967), .A2(n1992), .A3(n2032), .ZN(n2025) );
NOR2_X1 U1610 ( .A1(n2033), .A2(n2034), .ZN(n2032) );
NOR3_X1 U1611 ( .A1(n2035), .A2(n2036), .A3(n2037), .ZN(n1992) );
INV_X1 U1612 ( .A(n2034), .ZN(n2035) );
NAND2_X1 U1613 ( .A1(n1971), .A2(n2038), .ZN(n2034) );
NAND2_X1 U1614 ( .A1(n2030), .A2(n2039), .ZN(n2038) );
INV_X1 U1615 ( .A(n1994), .ZN(n1971) );
NOR2_X1 U1616 ( .A1(n2039), .A2(n2030), .ZN(n1994) );
NOR2_X1 U1617 ( .A1(n2040), .A2(n1995), .ZN(n2024) );
XOR2_X1 U1618 ( .A(KEYINPUT60), .B(n1988), .Z(n2040) );
INV_X1 U1619 ( .A(n2030), .ZN(n1988) );
NAND2_X1 U1620 ( .A1(n2041), .A2(n2042), .ZN(n2030) );
NAND2_X1 U1621 ( .A1(n2043), .A2(n2010), .ZN(n2042) );
XOR2_X1 U1622 ( .A(n2044), .B(n2009), .Z(n2043) );
XNOR2_X1 U1623 ( .A(KEYINPUT27), .B(n2045), .ZN(n2044) );
NOR2_X1 U1624 ( .A1(KEYINPUT47), .A2(n2005), .ZN(n2045) );
INV_X1 U1625 ( .A(n2019), .ZN(n2005) );
NAND2_X1 U1626 ( .A1(n2046), .A2(n2007), .ZN(n2041) );
INV_X1 U1627 ( .A(n2010), .ZN(n2007) );
NAND3_X1 U1628 ( .A1(n2047), .A2(n2048), .A3(n2049), .ZN(n2010) );
NAND2_X1 U1629 ( .A1(KEYINPUT50), .A2(n1788), .ZN(n2049) );
NAND3_X1 U1630 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n2050), .A3(RESTART), .ZN(n2048) );
NAND2_X1 U1631 ( .A1(n2051), .A2(n2003), .ZN(n2047) );
NAND2_X1 U1632 ( .A1(n1932), .A2(n2050), .ZN(n2051) );
INV_X1 U1633 ( .A(KEYINPUT50), .ZN(n2050) );
XOR2_X1 U1634 ( .A(n2019), .B(n2009), .Z(n2046) );
INV_X1 U1635 ( .A(n2011), .ZN(n2009) );
NAND3_X1 U1636 ( .A1(n2052), .A2(n2053), .A3(n2054), .ZN(n2011) );
OR2_X1 U1637 ( .A1(KEYINPUT22), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2054) );
NAND3_X1 U1638 ( .A1(KEYINPUT22), .A2(RMAX_REG_5__SCAN_IN), .A3(RESTART),
.ZN(n2053) );
NAND2_X1 U1639 ( .A1(n2055), .A2(n2003), .ZN(n2052) );
NAND2_X1 U1640 ( .A1(KEYINPUT22), .A2(n1809), .ZN(n2055) );
NAND2_X1 U1641 ( .A1(n2056), .A2(n2057), .ZN(n2019) );
NAND2_X1 U1642 ( .A1(n2058), .A2(n2059), .ZN(n2057) );
NAND2_X1 U1643 ( .A1(n2060), .A2(n2061), .ZN(n2059) );
XNOR2_X1 U1644 ( .A(KEYINPUT28), .B(n2062), .ZN(n2060) );
NAND2_X1 U1645 ( .A1(n2062), .A2(n2063), .ZN(n2056) );
NAND2_X1 U1646 ( .A1(n1947), .A2(REG4_REG_4__SCAN_IN), .ZN(n2022) );
NAND2_X1 U1647 ( .A1(n2064), .A2(DATA_OUT_REG_4__SCAN_IN), .ZN(n2021) );
XOR2_X1 U1648 ( .A(U280), .B(KEYINPUT21), .Z(n2064) );
NAND2_X1 U1649 ( .A1(n1950), .A2(RLAST_REG_4__SCAN_IN), .ZN(n2020) );
NAND4_X1 U1650 ( .A1(n2065), .A2(n2066), .A3(n2067), .A4(n2068), .ZN(U284));
NOR3_X1 U1651 ( .A1(n2069), .A2(n2070), .A3(n2071), .ZN(n2068) );
NOR3_X1 U1652 ( .A1(n1967), .A2(n2072), .A3(n2033), .ZN(n2071) );
NOR2_X1 U1653 ( .A1(n2036), .A2(n2037), .ZN(n2033) );
XOR2_X1 U1654 ( .A(n2073), .B(KEYINPUT15), .Z(n2037) );
INV_X1 U1655 ( .A(n2074), .ZN(n2036) );
NOR2_X1 U1656 ( .A1(n2073), .A2(n2074), .ZN(n2072) );
NAND2_X1 U1657 ( .A1(n2039), .A2(n2075), .ZN(n2074) );
OR2_X1 U1658 ( .A1(n2076), .A2(n2077), .ZN(n2039) );
NOR3_X1 U1659 ( .A1(n1964), .A2(n2028), .A3(n2078), .ZN(n2070) );
NOR2_X1 U1660 ( .A1(n2079), .A2(n2080), .ZN(n2078) );
AND2_X1 U1661 ( .A1(n2079), .A2(n2080), .ZN(n2028) );
NAND2_X1 U1662 ( .A1(n2031), .A2(n2075), .ZN(n2080) );
NAND2_X1 U1663 ( .A1(n2077), .A2(n2076), .ZN(n2075) );
INV_X1 U1664 ( .A(n2081), .ZN(n2077) );
NAND3_X1 U1665 ( .A1(n2082), .A2(n2083), .A3(n2081), .ZN(n2031) );
XOR2_X1 U1666 ( .A(KEYINPUT25), .B(n2084), .Z(n2083) );
NOR2_X1 U1667 ( .A1(n2081), .A2(n1995), .ZN(n2069) );
XNOR2_X1 U1668 ( .A(n2085), .B(n2058), .ZN(n2081) );
NAND2_X1 U1669 ( .A1(n2086), .A2(n2087), .ZN(n2058) );
NAND2_X1 U1670 ( .A1(RESTART), .A2(n1808), .ZN(n2087) );
OR2_X1 U1671 ( .A1(REG4_REG_4__SCAN_IN), .A2(RESTART), .ZN(n2086) );
XOR2_X1 U1672 ( .A(n2061), .B(n2062), .Z(n2085) );
NAND2_X1 U1673 ( .A1(n2088), .A2(n2089), .ZN(n2062) );
NAND2_X1 U1674 ( .A1(RESTART), .A2(n1827), .ZN(n2089) );
NAND2_X1 U1675 ( .A1(n1807), .A2(n2003), .ZN(n2088) );
INV_X1 U1676 ( .A(n2063), .ZN(n2061) );
NAND2_X1 U1677 ( .A1(n2090), .A2(n2091), .ZN(n2063) );
NAND2_X1 U1678 ( .A1(n2092), .A2(n2093), .ZN(n2091) );
NAND2_X1 U1679 ( .A1(n2094), .A2(n2095), .ZN(n2093) );
XOR2_X1 U1680 ( .A(n2096), .B(KEYINPUT54), .Z(n2095) );
NAND2_X1 U1681 ( .A1(n2096), .A2(n2097), .ZN(n2090) );
NAND2_X1 U1682 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1724), .ZN(n2067) );
NAND2_X1 U1683 ( .A1(n1950), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2066) );
NAND2_X1 U1684 ( .A1(n1947), .A2(REG4_REG_3__SCAN_IN), .ZN(n2065) );
NAND4_X1 U1685 ( .A1(n2098), .A2(n2099), .A3(n2100), .A4(n2101), .ZN(U283));
NOR3_X1 U1686 ( .A1(n2102), .A2(n2103), .A3(n2104), .ZN(n2101) );
NOR3_X1 U1687 ( .A1(n1964), .A2(n2079), .A3(n2105), .ZN(n2104) );
NOR3_X1 U1688 ( .A1(n2106), .A2(n2107), .A3(n2108), .ZN(n2105) );
AND3_X1 U1689 ( .A1(KEYINPUT35), .A2(n2109), .A3(n2110), .ZN(n2108) );
NOR2_X1 U1690 ( .A1(KEYINPUT35), .A2(n2111), .ZN(n2107) );
AND2_X1 U1691 ( .A1(n2112), .A2(n2113), .ZN(n2079) );
NAND3_X1 U1692 ( .A1(n2076), .A2(n2114), .A3(n2115), .ZN(n2113) );
NAND2_X1 U1693 ( .A1(KEYINPUT2), .A2(n2084), .ZN(n2115) );
INV_X1 U1694 ( .A(n2106), .ZN(n2114) );
NOR3_X1 U1695 ( .A1(n2084), .A2(KEYINPUT2), .A3(n2082), .ZN(n2106) );
NAND2_X1 U1696 ( .A1(n2084), .A2(n2082), .ZN(n2076) );
NOR3_X1 U1697 ( .A1(n1967), .A2(n2073), .A3(n2116), .ZN(n2103) );
XOR2_X1 U1698 ( .A(n2117), .B(KEYINPUT29), .Z(n2116) );
NAND3_X1 U1699 ( .A1(n2118), .A2(n2119), .A3(n2120), .ZN(n2117) );
NAND2_X1 U1700 ( .A1(n2121), .A2(n2122), .ZN(n2120) );
OR2_X1 U1701 ( .A1(n2111), .A2(KEYINPUT3), .ZN(n2119) );
NAND3_X1 U1702 ( .A1(n2123), .A2(n2124), .A3(KEYINPUT3), .ZN(n2118) );
AND2_X1 U1703 ( .A1(n2112), .A2(n2125), .ZN(n2073) );
XOR2_X1 U1704 ( .A(n2122), .B(n2082), .Z(n2125) );
INV_X1 U1705 ( .A(n2111), .ZN(n2112) );
NAND2_X1 U1706 ( .A1(n2124), .A2(n2109), .ZN(n2111) );
NOR2_X1 U1707 ( .A1(n2082), .A2(n1995), .ZN(n2102) );
INV_X1 U1708 ( .A(n2121), .ZN(n2082) );
NAND2_X1 U1709 ( .A1(n2126), .A2(n2127), .ZN(n2121) );
NAND2_X1 U1710 ( .A1(n2128), .A2(n2097), .ZN(n2127) );
NAND2_X1 U1711 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
NAND2_X1 U1712 ( .A1(n2131), .A2(n2092), .ZN(n2130) );
XOR2_X1 U1713 ( .A(KEYINPUT36), .B(n2132), .Z(n2129) );
NOR2_X1 U1714 ( .A1(n2133), .A2(n2092), .ZN(n2132) );
NAND2_X1 U1715 ( .A1(n2134), .A2(n2094), .ZN(n2126) );
INV_X1 U1716 ( .A(n2097), .ZN(n2094) );
NAND2_X1 U1717 ( .A1(n2135), .A2(n2136), .ZN(n2097) );
NAND2_X1 U1718 ( .A1(n2137), .A2(n2138), .ZN(n2136) );
NAND2_X1 U1719 ( .A1(n2139), .A2(n2140), .ZN(n2137) );
XOR2_X1 U1720 ( .A(n2141), .B(KEYINPUT23), .Z(n2140) );
NAND2_X1 U1721 ( .A1(n2141), .A2(n2142), .ZN(n2135) );
NAND2_X1 U1722 ( .A1(n2143), .A2(n2144), .ZN(n2134) );
NAND2_X1 U1723 ( .A1(n2145), .A2(n2133), .ZN(n2144) );
XOR2_X1 U1724 ( .A(n2131), .B(KEYINPUT14), .Z(n2133) );
INV_X1 U1725 ( .A(n2096), .ZN(n2131) );
INV_X1 U1726 ( .A(n2092), .ZN(n2145) );
NAND2_X1 U1727 ( .A1(n2092), .A2(n2096), .ZN(n2143) );
NAND2_X1 U1728 ( .A1(n2146), .A2(n2147), .ZN(n2096) );
NAND2_X1 U1729 ( .A1(RESTART), .A2(n1839), .ZN(n2147) );
NAND2_X1 U1730 ( .A1(n1831), .A2(n2003), .ZN(n2146) );
NAND2_X1 U1731 ( .A1(n2148), .A2(n2149), .ZN(n2092) );
NAND2_X1 U1732 ( .A1(RESTART), .A2(n1793), .ZN(n2149) );
OR2_X1 U1733 ( .A1(REG4_REG_3__SCAN_IN), .A2(RESTART), .ZN(n2148) );
XOR2_X1 U1734 ( .A(n2150), .B(KEYINPUT26), .Z(n2100) );
NAND2_X1 U1735 ( .A1(n1947), .A2(REG4_REG_2__SCAN_IN), .ZN(n2150) );
NAND2_X1 U1736 ( .A1(n1950), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2099) );
NAND2_X1 U1737 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1724), .ZN(n2098) );
NAND4_X1 U1738 ( .A1(n2151), .A2(n2152), .A3(n2153), .A4(n2154), .ZN(U282));
NOR3_X1 U1739 ( .A1(n2155), .A2(n2156), .A3(n2157), .ZN(n2154) );
NOR2_X1 U1740 ( .A1(n2158), .A2(n1964), .ZN(n2157) );
XOR2_X1 U1741 ( .A(n2159), .B(n2123), .Z(n2158) );
INV_X1 U1742 ( .A(n2109), .ZN(n2123) );
NAND2_X1 U1743 ( .A1(KEYINPUT6), .A2(n2110), .ZN(n2159) );
INV_X1 U1744 ( .A(n2124), .ZN(n2110) );
NOR2_X1 U1745 ( .A1(n1967), .A2(n2160), .ZN(n2156) );
XOR2_X1 U1746 ( .A(n2161), .B(n2162), .Z(n2160) );
XOR2_X1 U1747 ( .A(n2124), .B(KEYINPUT10), .Z(n2162) );
NAND2_X1 U1748 ( .A1(n2122), .A2(n2163), .ZN(n2124) );
NAND2_X1 U1749 ( .A1(n2164), .A2(n2165), .ZN(n2163) );
INV_X1 U1750 ( .A(n2084), .ZN(n2122) );
NOR2_X1 U1751 ( .A1(n2165), .A2(n2164), .ZN(n2084) );
NAND2_X1 U1752 ( .A1(KEYINPUT16), .A2(n2109), .ZN(n2161) );
NOR2_X1 U1753 ( .A1(n2166), .A2(n1995), .ZN(n2155) );
INV_X1 U1754 ( .A(n2164), .ZN(n2166) );
XOR2_X1 U1755 ( .A(n2167), .B(n2139), .Z(n2164) );
INV_X1 U1756 ( .A(n2142), .ZN(n2139) );
NAND2_X1 U1757 ( .A1(n2168), .A2(n2169), .ZN(n2142) );
NAND2_X1 U1758 ( .A1(RESTART), .A2(n1836), .ZN(n2169) );
NAND2_X1 U1759 ( .A1(n1800), .A2(n2003), .ZN(n2168) );
NAND2_X1 U1760 ( .A1(n2170), .A2(n2171), .ZN(n2167) );
NAND2_X1 U1761 ( .A1(n2172), .A2(n2138), .ZN(n2171) );
INV_X1 U1762 ( .A(n2173), .ZN(n2138) );
NAND2_X1 U1763 ( .A1(KEYINPUT63), .A2(n2141), .ZN(n2172) );
NAND3_X1 U1764 ( .A1(KEYINPUT7), .A2(n2141), .A3(n2173), .ZN(n2170) );
NOR2_X1 U1765 ( .A1(n2174), .A2(n2175), .ZN(n2173) );
AND2_X1 U1766 ( .A1(n2176), .A2(n2177), .ZN(n2175) );
NAND2_X1 U1767 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
XOR2_X1 U1768 ( .A(n2180), .B(KEYINPUT19), .Z(n2178) );
NAND2_X1 U1769 ( .A1(n2181), .A2(n2182), .ZN(n2141) );
NAND2_X1 U1770 ( .A1(RESTART), .A2(n1806), .ZN(n2182) );
NAND2_X1 U1771 ( .A1(n2183), .A2(n2003), .ZN(n2181) );
NAND2_X1 U1772 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1724), .ZN(n2153) );
NAND2_X1 U1773 ( .A1(n1950), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2152) );
NAND2_X1 U1774 ( .A1(n1947), .A2(REG4_REG_1__SCAN_IN), .ZN(n2151) );
NAND3_X1 U1775 ( .A1(n2184), .A2(n2185), .A3(n2186), .ZN(U281) );
NOR3_X1 U1776 ( .A1(n2187), .A2(n2188), .A3(n2189), .ZN(n2186) );
AND2_X1 U1777 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1950), .ZN(n2189) );
AND3_X1 U1778 ( .A1(n1865), .A2(n2003), .A3(n2190), .ZN(n1950) );
NOR2_X1 U1779 ( .A1(n2191), .A2(n2109), .ZN(n2188) );
NAND2_X1 U1780 ( .A1(n2165), .A2(n2192), .ZN(n2109) );
NAND3_X1 U1781 ( .A1(n2193), .A2(n2194), .A3(n2195), .ZN(n2192) );
NAND2_X1 U1782 ( .A1(n2196), .A2(n2197), .ZN(n2165) );
NAND2_X1 U1783 ( .A1(n2195), .A2(n2193), .ZN(n2197) );
NAND2_X1 U1784 ( .A1(n2198), .A2(n2199), .ZN(n2193) );
NAND2_X1 U1785 ( .A1(n2200), .A2(n2201), .ZN(n2195) );
NAND2_X1 U1786 ( .A1(RESTART), .A2(n2202), .ZN(n2201) );
NAND2_X1 U1787 ( .A1(n1749), .A2(n2203), .ZN(n2202) );
NAND2_X1 U1788 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n2199), .ZN(n2203) );
INV_X1 U1789 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1749) );
NAND2_X1 U1790 ( .A1(n2204), .A2(n2003), .ZN(n2200) );
NAND2_X1 U1791 ( .A1(n1802), .A2(n2205), .ZN(n2204) );
NAND2_X1 U1792 ( .A1(REG4_REG_0__SCAN_IN), .A2(n2199), .ZN(n2205) );
INV_X1 U1793 ( .A(KEYINPUT53), .ZN(n2199) );
INV_X1 U1794 ( .A(DATA_IN_0_), .ZN(n1802) );
NOR2_X1 U1795 ( .A1(n1952), .A2(n1972), .ZN(n2191) );
INV_X1 U1796 ( .A(n1964), .ZN(n1972) );
NAND3_X1 U1797 ( .A1(n2190), .A2(RESTART), .A3(n2206), .ZN(n1964) );
INV_X1 U1798 ( .A(n1967), .ZN(n1952) );
NAND4_X1 U1799 ( .A1(ENABLE), .A2(n2190), .A3(n2207), .A4(n2208), .ZN(n1967));
NOR2_X1 U1800 ( .A1(RESTART), .A2(AVERAGE), .ZN(n2207) );
NOR2_X1 U1801 ( .A1(n2196), .A2(n1995), .ZN(n2187) );
NAND3_X1 U1802 ( .A1(n2209), .A2(n2210), .A3(n2190), .ZN(n1995) );
NAND2_X1 U1803 ( .A1(n2211), .A2(n2003), .ZN(n2210) );
OR4_X1 U1804 ( .A1(n2208), .A2(n1865), .A3(n2212), .A4(AVERAGE), .ZN(n2211));
NOR2_X1 U1805 ( .A1(n2213), .A2(KEYINPUT18), .ZN(n2212) );
INV_X1 U1806 ( .A(n2206), .ZN(n2213) );
INV_X1 U1807 ( .A(ENABLE), .ZN(n1865) );
NAND3_X1 U1808 ( .A1(n2214), .A2(n2215), .A3(n2216), .ZN(n2208) );
OR2_X1 U1809 ( .A1(n1780), .A2(n2217), .ZN(n2216) );
NAND2_X1 U1810 ( .A1(KEYINPUT38), .A2(n2218), .ZN(n2215) );
NAND2_X1 U1811 ( .A1(REG4_REG_7__SCAN_IN), .A2(DATA_IN_7_), .ZN(n2218) );
NAND2_X1 U1812 ( .A1(REG4_REG_7__SCAN_IN), .A2(n2219), .ZN(n2214) );
NAND2_X1 U1813 ( .A1(n2217), .A2(n2220), .ZN(n2219) );
OR2_X1 U1814 ( .A1(n1780), .A2(KEYINPUT38), .ZN(n2220) );
INV_X1 U1815 ( .A(DATA_IN_7_), .ZN(n1780) );
XOR2_X1 U1816 ( .A(n2221), .B(KEYINPUT58), .Z(n2217) );
NAND2_X1 U1817 ( .A1(n2222), .A2(n2223), .ZN(n2221) );
NAND2_X1 U1818 ( .A1(REG4_REG_6__SCAN_IN), .A2(n2224), .ZN(n2223) );
NAND2_X1 U1819 ( .A1(n2225), .A2(n2226), .ZN(n2224) );
XOR2_X1 U1820 ( .A(KEYINPUT55), .B(DATA_IN_6_), .Z(n2225) );
OR2_X1 U1821 ( .A1(n2226), .A2(n1784), .ZN(n2222) );
INV_X1 U1822 ( .A(DATA_IN_6_), .ZN(n1784) );
NAND2_X1 U1823 ( .A1(n2227), .A2(n2228), .ZN(n2226) );
NAND3_X1 U1824 ( .A1(n2229), .A2(n2230), .A3(n2231), .ZN(n2228) );
NAND2_X1 U1825 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2231) );
NAND3_X1 U1826 ( .A1(n2232), .A2(n2233), .A3(n2234), .ZN(n2230) );
NAND2_X1 U1827 ( .A1(n2235), .A2(n1807), .ZN(n2234) );
INV_X1 U1828 ( .A(DATA_IN_4_), .ZN(n1807) );
XOR2_X1 U1829 ( .A(REG4_REG_4__SCAN_IN), .B(KEYINPUT57), .Z(n2235) );
NAND3_X1 U1830 ( .A1(n2236), .A2(n2237), .A3(n2238), .ZN(n2233) );
NAND2_X1 U1831 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2238) );
NAND3_X1 U1832 ( .A1(n2239), .A2(n2240), .A3(n2241), .ZN(n2237) );
NAND2_X1 U1833 ( .A1(n1800), .A2(n2183), .ZN(n2241) );
INV_X1 U1834 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2183) );
INV_X1 U1835 ( .A(DATA_IN_2_), .ZN(n1800) );
NAND2_X1 U1836 ( .A1(n2242), .A2(n2243), .ZN(n2240) );
INV_X1 U1837 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2243) );
OR2_X1 U1838 ( .A1(n2244), .A2(n1804), .ZN(n2242) );
NAND2_X1 U1839 ( .A1(n2244), .A2(n1804), .ZN(n2239) );
NAND2_X1 U1840 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2236) );
NAND2_X1 U1841 ( .A1(n2245), .A2(n1831), .ZN(n2232) );
INV_X1 U1842 ( .A(DATA_IN_3_), .ZN(n1831) );
XNOR2_X1 U1843 ( .A(REG4_REG_3__SCAN_IN), .B(KEYINPUT59), .ZN(n2245) );
NAND2_X1 U1844 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2229) );
NAND2_X1 U1845 ( .A1(n1932), .A2(n1809), .ZN(n2227) );
INV_X1 U1846 ( .A(DATA_IN_5_), .ZN(n1809) );
INV_X1 U1847 ( .A(REG4_REG_5__SCAN_IN), .ZN(n1932) );
NAND3_X1 U1848 ( .A1(KEYINPUT18), .A2(n2206), .A3(RESTART), .ZN(n2209) );
XOR2_X1 U1849 ( .A(n2246), .B(KEYINPUT49), .Z(n2206) );
NAND2_X1 U1850 ( .A1(n2247), .A2(n2248), .ZN(n2246) );
NAND2_X1 U1851 ( .A1(n2249), .A2(n1810), .ZN(n2248) );
INV_X1 U1852 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1810) );
OR2_X1 U1853 ( .A1(n2250), .A2(n1816), .ZN(n2249) );
NAND2_X1 U1854 ( .A1(n2250), .A2(n1816), .ZN(n2247) );
INV_X1 U1855 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1816) );
NAND2_X1 U1856 ( .A1(n2251), .A2(n2252), .ZN(n2250) );
NAND2_X1 U1857 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n2253), .ZN(n2252) );
NAND2_X1 U1858 ( .A1(n1820), .A2(n2254), .ZN(n2253) );
OR2_X1 U1859 ( .A1(n2254), .A2(n1820), .ZN(n2251) );
INV_X1 U1860 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1820) );
NAND2_X1 U1861 ( .A1(n2255), .A2(n2256), .ZN(n2254) );
NAND2_X1 U1862 ( .A1(n2257), .A2(n1788), .ZN(n2256) );
INV_X1 U1863 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1788) );
NAND2_X1 U1864 ( .A1(n2258), .A2(n2259), .ZN(n2257) );
XOR2_X1 U1865 ( .A(RMAX_REG_5__SCAN_IN), .B(KEYINPUT51), .Z(n2258) );
OR2_X1 U1866 ( .A1(n2259), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2255) );
NAND2_X1 U1867 ( .A1(n2260), .A2(n2261), .ZN(n2259) );
NAND2_X1 U1868 ( .A1(n2262), .A2(RMIN_REG_4__SCAN_IN), .ZN(n2261) );
XOR2_X1 U1869 ( .A(n1827), .B(KEYINPUT32), .Z(n2262) );
NAND3_X1 U1870 ( .A1(n2263), .A2(n2264), .A3(n2265), .ZN(n2260) );
NAND2_X1 U1871 ( .A1(n1827), .A2(n1808), .ZN(n2265) );
INV_X1 U1872 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1808) );
INV_X1 U1873 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1827) );
NAND3_X1 U1874 ( .A1(n2266), .A2(n2267), .A3(n2268), .ZN(n2264) );
NAND2_X1 U1875 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2268) );
NAND3_X1 U1876 ( .A1(n2269), .A2(n2270), .A3(n2271), .ZN(n2267) );
NAND2_X1 U1877 ( .A1(n1836), .A2(n1806), .ZN(n2271) );
INV_X1 U1878 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1806) );
INV_X1 U1879 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1836) );
NAND2_X1 U1880 ( .A1(n2272), .A2(n2273), .ZN(n2270) );
INV_X1 U1881 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n2273) );
OR2_X1 U1882 ( .A1(n2274), .A2(n1838), .ZN(n2272) );
NAND2_X1 U1883 ( .A1(n2274), .A2(n1838), .ZN(n2269) );
NAND2_X1 U1884 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n2275), .ZN(n2266) );
XOR2_X1 U1885 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT13), .Z(n2275) );
NAND2_X1 U1886 ( .A1(n1839), .A2(n1793), .ZN(n2263) );
INV_X1 U1887 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1793) );
INV_X1 U1888 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1839) );
INV_X1 U1889 ( .A(n2194), .ZN(n2196) );
NAND4_X1 U1890 ( .A1(n2276), .A2(n2277), .A3(n2278), .A4(n2279), .ZN(n2194));
NAND3_X1 U1891 ( .A1(n2280), .A2(n2281), .A3(n2282), .ZN(n2279) );
OR2_X1 U1892 ( .A1(n2282), .A2(n2280), .ZN(n2278) );
NOR2_X1 U1893 ( .A1(n2180), .A2(n2198), .ZN(n2280) );
NAND2_X1 U1894 ( .A1(n2174), .A2(n2283), .ZN(n2277) );
NAND2_X1 U1895 ( .A1(n2176), .A2(n2284), .ZN(n2283) );
AND2_X1 U1896 ( .A1(n2281), .A2(n2180), .ZN(n2174) );
INV_X1 U1897 ( .A(n2179), .ZN(n2281) );
NAND2_X1 U1898 ( .A1(n2179), .A2(n2285), .ZN(n2276) );
NAND2_X1 U1899 ( .A1(n2286), .A2(n2282), .ZN(n2285) );
INV_X1 U1900 ( .A(KEYINPUT1), .ZN(n2282) );
XOR2_X1 U1901 ( .A(n2287), .B(n2198), .Z(n2286) );
INV_X1 U1902 ( .A(n2176), .ZN(n2198) );
NAND2_X1 U1903 ( .A1(n2288), .A2(n2289), .ZN(n2176) );
NAND2_X1 U1904 ( .A1(n2244), .A2(n2003), .ZN(n2289) );
NAND2_X1 U1905 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2244) );
NAND2_X1 U1906 ( .A1(RESTART), .A2(n2274), .ZN(n2288) );
NAND2_X1 U1907 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2274) );
NAND2_X1 U1908 ( .A1(n2180), .A2(n2284), .ZN(n2287) );
INV_X1 U1909 ( .A(KEYINPUT44), .ZN(n2284) );
NAND2_X1 U1910 ( .A1(n2290), .A2(n2291), .ZN(n2180) );
NAND2_X1 U1911 ( .A1(RESTART), .A2(n1838), .ZN(n2291) );
INV_X1 U1912 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1838) );
NAND2_X1 U1913 ( .A1(n1804), .A2(n2003), .ZN(n2290) );
INV_X1 U1914 ( .A(DATA_IN_1_), .ZN(n1804) );
NAND2_X1 U1915 ( .A1(n2292), .A2(n2293), .ZN(n2179) );
NAND2_X1 U1916 ( .A1(REG4_REG_1__SCAN_IN), .A2(n2003), .ZN(n2293) );
NAND2_X1 U1917 ( .A1(RMIN_REG_1__SCAN_IN), .A2(RESTART), .ZN(n2292) );
NAND2_X1 U1918 ( .A1(n1947), .A2(REG4_REG_0__SCAN_IN), .ZN(n2185) );
AND4_X1 U1919 ( .A1(AVERAGE), .A2(ENABLE), .A3(n2190), .A4(n2003), .ZN(n1947) );
INV_X1 U1920 ( .A(RESTART), .ZN(n2003) );
NOR2_X1 U1921 ( .A1(n1753), .A2(n1724), .ZN(n2190) );
NAND2_X1 U1922 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1724), .ZN(n2184) );
INV_X1 U1923 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1753) );
NOR2_X1 U1924 ( .A1(n1748), .A2(STATO_REG_1__SCAN_IN), .ZN(n2294) );
INV_X1 U1925 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1748) );
endmodule


