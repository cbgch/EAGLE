//Key = 1110100001100001001100000101011101010101101001011111011000000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287;

XNOR2_X1 U724 ( .A(G107), .B(n984), .ZN(G9) );
NOR2_X1 U725 ( .A1(n985), .A2(n986), .ZN(G75) );
NOR4_X1 U726 ( .A1(n987), .A2(n988), .A3(n989), .A4(n990), .ZN(n986) );
NAND3_X1 U727 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n987) );
NAND2_X1 U728 ( .A1(n994), .A2(n995), .ZN(n993) );
NAND2_X1 U729 ( .A1(n996), .A2(n997), .ZN(n994) );
NAND3_X1 U730 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
NAND2_X1 U731 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NAND2_X1 U732 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U733 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U734 ( .A1(n1007), .A2(n1008), .ZN(n1001) );
NAND2_X1 U735 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U736 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
INV_X1 U737 ( .A(n1013), .ZN(n1009) );
NAND3_X1 U738 ( .A1(n1007), .A2(n1014), .A3(n1003), .ZN(n996) );
NAND3_X1 U739 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND2_X1 U740 ( .A1(n1000), .A2(n1018), .ZN(n1017) );
NAND2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
XNOR2_X1 U742 ( .A(n1000), .B(KEYINPUT10), .ZN(n1019) );
NAND2_X1 U743 ( .A1(n998), .A2(n1021), .ZN(n1015) );
NAND3_X1 U744 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1021) );
OR2_X1 U745 ( .A1(n1025), .A2(KEYINPUT61), .ZN(n1023) );
NAND3_X1 U746 ( .A1(n1026), .A2(n1027), .A3(KEYINPUT61), .ZN(n1022) );
NOR3_X1 U747 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n985) );
INV_X1 U748 ( .A(n991), .ZN(n1028) );
NAND4_X1 U749 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n991) );
NOR4_X1 U750 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
XOR2_X1 U751 ( .A(KEYINPUT16), .B(n1037), .Z(n1036) );
NOR2_X1 U752 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XNOR2_X1 U753 ( .A(n1040), .B(KEYINPUT36), .ZN(n1038) );
XOR2_X1 U754 ( .A(G472), .B(n1041), .Z(n1035) );
NOR2_X1 U755 ( .A1(KEYINPUT34), .A2(n1042), .ZN(n1041) );
INV_X1 U756 ( .A(n1007), .ZN(n1033) );
NOR3_X1 U757 ( .A1(n1026), .A2(n1043), .A3(n1011), .ZN(n1031) );
NAND2_X1 U758 ( .A1(n1044), .A2(n1045), .ZN(n1030) );
XOR2_X1 U759 ( .A(KEYINPUT7), .B(n1046), .Z(n1044) );
NAND2_X1 U760 ( .A1(n1039), .A2(n1047), .ZN(n1029) );
XOR2_X1 U761 ( .A(KEYINPUT11), .B(G469), .Z(n1039) );
XOR2_X1 U762 ( .A(n1048), .B(n1049), .Z(G72) );
XOR2_X1 U763 ( .A(n1050), .B(n1051), .Z(n1049) );
NOR2_X1 U764 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U765 ( .A(n1054), .B(n1055), .Z(n1053) );
XNOR2_X1 U766 ( .A(n1056), .B(n1057), .ZN(n1055) );
XNOR2_X1 U767 ( .A(KEYINPUT6), .B(n1058), .ZN(n1057) );
XNOR2_X1 U768 ( .A(n1059), .B(n1060), .ZN(n1054) );
NOR2_X1 U769 ( .A1(G953), .A2(n1061), .ZN(n1050) );
NOR2_X1 U770 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
XNOR2_X1 U771 ( .A(KEYINPUT18), .B(n990), .ZN(n1063) );
NOR2_X1 U772 ( .A1(n1064), .A2(n992), .ZN(n1048) );
AND2_X1 U773 ( .A1(G227), .A2(G900), .ZN(n1064) );
NAND2_X1 U774 ( .A1(n1065), .A2(n1066), .ZN(G69) );
NAND2_X1 U775 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U776 ( .A(KEYINPUT4), .B(n1069), .Z(n1065) );
NOR2_X1 U777 ( .A1(n1067), .A2(n1068), .ZN(n1069) );
NAND2_X1 U778 ( .A1(G953), .A2(n1070), .ZN(n1068) );
NAND2_X1 U779 ( .A1(G898), .A2(G224), .ZN(n1070) );
NAND2_X1 U780 ( .A1(n1071), .A2(n1072), .ZN(n1067) );
NAND2_X1 U781 ( .A1(n1073), .A2(n992), .ZN(n1072) );
XOR2_X1 U782 ( .A(n988), .B(n1074), .Z(n1073) );
NAND3_X1 U783 ( .A1(G898), .A2(n1074), .A3(G953), .ZN(n1071) );
XNOR2_X1 U784 ( .A(n1075), .B(n1076), .ZN(n1074) );
XOR2_X1 U785 ( .A(KEYINPUT62), .B(KEYINPUT2), .Z(n1076) );
NOR2_X1 U786 ( .A1(n1077), .A2(n1078), .ZN(G66) );
XOR2_X1 U787 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U788 ( .A1(n1081), .A2(KEYINPUT32), .ZN(n1079) );
NOR2_X1 U789 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR2_X1 U790 ( .A1(n1077), .A2(n1084), .ZN(G63) );
XOR2_X1 U791 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U792 ( .A1(n1087), .A2(G478), .ZN(n1085) );
NOR2_X1 U793 ( .A1(n1077), .A2(n1088), .ZN(G60) );
XOR2_X1 U794 ( .A(n1089), .B(n1090), .Z(n1088) );
NAND2_X1 U795 ( .A1(n1087), .A2(G475), .ZN(n1089) );
XNOR2_X1 U796 ( .A(G104), .B(n1091), .ZN(G6) );
NOR2_X1 U797 ( .A1(n1077), .A2(n1092), .ZN(G57) );
XOR2_X1 U798 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U799 ( .A1(n1095), .A2(KEYINPUT63), .ZN(n1093) );
XOR2_X1 U800 ( .A(n1096), .B(n1097), .Z(n1095) );
XOR2_X1 U801 ( .A(n1098), .B(n1099), .Z(n1096) );
NOR2_X1 U802 ( .A1(KEYINPUT5), .A2(n1100), .ZN(n1099) );
XOR2_X1 U803 ( .A(n1101), .B(n1102), .Z(n1100) );
XNOR2_X1 U804 ( .A(KEYINPUT50), .B(n1056), .ZN(n1102) );
NAND2_X1 U805 ( .A1(n1087), .A2(G472), .ZN(n1098) );
NOR2_X1 U806 ( .A1(n1077), .A2(n1103), .ZN(G54) );
XOR2_X1 U807 ( .A(n1104), .B(n1105), .Z(n1103) );
XNOR2_X1 U808 ( .A(n1106), .B(n1107), .ZN(n1105) );
NAND2_X1 U809 ( .A1(n1087), .A2(G469), .ZN(n1106) );
INV_X1 U810 ( .A(n1083), .ZN(n1087) );
XOR2_X1 U811 ( .A(n1108), .B(n1109), .Z(n1104) );
XNOR2_X1 U812 ( .A(KEYINPUT42), .B(n1110), .ZN(n1109) );
NOR2_X1 U813 ( .A1(KEYINPUT12), .A2(n1111), .ZN(n1110) );
XNOR2_X1 U814 ( .A(n1112), .B(n1113), .ZN(n1111) );
NAND2_X1 U815 ( .A1(KEYINPUT49), .A2(n1056), .ZN(n1108) );
NOR2_X1 U816 ( .A1(n1077), .A2(n1114), .ZN(G51) );
XOR2_X1 U817 ( .A(n1075), .B(n1115), .Z(n1114) );
XOR2_X1 U818 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U819 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U820 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U821 ( .A1(n1122), .A2(KEYINPUT13), .ZN(n1120) );
NOR2_X1 U822 ( .A1(KEYINPUT59), .A2(n1123), .ZN(n1122) );
NOR2_X1 U823 ( .A1(n1124), .A2(n1125), .ZN(n1118) );
NOR2_X1 U824 ( .A1(n1126), .A2(KEYINPUT59), .ZN(n1125) );
NOR2_X1 U825 ( .A1(KEYINPUT13), .A2(n1127), .ZN(n1126) );
INV_X1 U826 ( .A(n1121), .ZN(n1127) );
XNOR2_X1 U827 ( .A(n1101), .B(n1060), .ZN(n1121) );
OR2_X1 U828 ( .A1(n1083), .A2(n1045), .ZN(n1116) );
NAND2_X1 U829 ( .A1(G902), .A2(n1128), .ZN(n1083) );
OR3_X1 U830 ( .A1(n990), .A2(n989), .A3(n988), .ZN(n1128) );
NAND4_X1 U831 ( .A1(n1091), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n988) );
AND3_X1 U832 ( .A1(n1132), .A2(n984), .A3(n1133), .ZN(n1131) );
NAND3_X1 U833 ( .A1(n998), .A2(n1134), .A3(n1135), .ZN(n984) );
NAND2_X1 U834 ( .A1(n1136), .A2(n1137), .ZN(n1130) );
NAND2_X1 U835 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U836 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U837 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U838 ( .A1(n1144), .A2(n1007), .ZN(n1143) );
NAND2_X1 U839 ( .A1(n1018), .A2(n1135), .ZN(n1142) );
XNOR2_X1 U840 ( .A(KEYINPUT30), .B(n1145), .ZN(n1138) );
NAND3_X1 U841 ( .A1(n998), .A2(n1134), .A3(n1146), .ZN(n1091) );
XOR2_X1 U842 ( .A(n1062), .B(KEYINPUT21), .Z(n989) );
NAND4_X1 U843 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1062) );
NAND3_X1 U844 ( .A1(n1135), .A2(n1151), .A3(n1152), .ZN(n1148) );
XNOR2_X1 U845 ( .A(KEYINPUT22), .B(n1153), .ZN(n1151) );
NAND2_X1 U846 ( .A1(n1154), .A2(n1000), .ZN(n1147) );
XOR2_X1 U847 ( .A(n1155), .B(KEYINPUT37), .Z(n1154) );
NAND4_X1 U848 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n990) );
NOR2_X1 U849 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND3_X1 U850 ( .A1(n1020), .A2(n1146), .A3(n1152), .ZN(n1158) );
NAND4_X1 U851 ( .A1(n1018), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1157) );
INV_X1 U852 ( .A(KEYINPUT45), .ZN(n1164) );
NAND2_X1 U853 ( .A1(n1165), .A2(KEYINPUT45), .ZN(n1156) );
NOR2_X1 U854 ( .A1(n992), .A2(G952), .ZN(n1077) );
XOR2_X1 U855 ( .A(G146), .B(n1161), .Z(G48) );
AND3_X1 U856 ( .A1(n1144), .A2(n1146), .A3(n1163), .ZN(n1161) );
XOR2_X1 U857 ( .A(G143), .B(n1165), .Z(G45) );
AND3_X1 U858 ( .A1(n1166), .A2(n1018), .A3(n1163), .ZN(n1165) );
XNOR2_X1 U859 ( .A(n1058), .B(n1167), .ZN(G42) );
NOR4_X1 U860 ( .A1(KEYINPUT14), .A2(n1005), .A3(n1168), .A4(n1169), .ZN(n1167) );
INV_X1 U861 ( .A(n1020), .ZN(n1168) );
XOR2_X1 U862 ( .A(G137), .B(n1160), .Z(G39) );
AND3_X1 U863 ( .A1(n1144), .A2(n1007), .A3(n1152), .ZN(n1160) );
INV_X1 U864 ( .A(n1169), .ZN(n1152) );
XOR2_X1 U865 ( .A(G134), .B(n1170), .Z(G36) );
NOR3_X1 U866 ( .A1(n1169), .A2(n1006), .A3(n1153), .ZN(n1170) );
NAND2_X1 U867 ( .A1(n1171), .A2(n1000), .ZN(n1169) );
INV_X1 U868 ( .A(n1025), .ZN(n1000) );
XOR2_X1 U869 ( .A(G131), .B(n1172), .Z(G33) );
NOR2_X1 U870 ( .A1(n1155), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U871 ( .A(KEYINPUT19), .B(n1025), .ZN(n1173) );
NAND2_X1 U872 ( .A1(n1027), .A2(n1174), .ZN(n1025) );
NAND3_X1 U873 ( .A1(n1018), .A2(n1146), .A3(n1171), .ZN(n1155) );
XNOR2_X1 U874 ( .A(G128), .B(n1149), .ZN(G30) );
NAND3_X1 U875 ( .A1(n1144), .A2(n1135), .A3(n1163), .ZN(n1149) );
AND2_X1 U876 ( .A1(n1171), .A2(n1136), .ZN(n1163) );
AND2_X1 U877 ( .A1(n1013), .A2(n1175), .ZN(n1171) );
XNOR2_X1 U878 ( .A(G101), .B(n1129), .ZN(G3) );
NAND3_X1 U879 ( .A1(n1007), .A2(n1134), .A3(n1018), .ZN(n1129) );
AND3_X1 U880 ( .A1(n1013), .A2(n1176), .A3(n1136), .ZN(n1134) );
XNOR2_X1 U881 ( .A(G125), .B(n1150), .ZN(G27) );
NAND3_X1 U882 ( .A1(n1020), .A2(n1146), .A3(n1177), .ZN(n1150) );
AND3_X1 U883 ( .A1(n1003), .A2(n1175), .A3(n1136), .ZN(n1177) );
NAND2_X1 U884 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
NAND3_X1 U885 ( .A1(G902), .A2(n995), .A3(n1052), .ZN(n1179) );
NOR2_X1 U886 ( .A1(n992), .A2(G900), .ZN(n1052) );
XNOR2_X1 U887 ( .A(G122), .B(n1132), .ZN(G24) );
NAND4_X1 U888 ( .A1(n1166), .A2(n1140), .A3(n998), .A4(n1136), .ZN(n1132) );
NOR2_X1 U889 ( .A1(n1180), .A2(n1181), .ZN(n998) );
INV_X1 U890 ( .A(n1162), .ZN(n1166) );
NAND2_X1 U891 ( .A1(n1182), .A2(n1183), .ZN(n1162) );
XNOR2_X1 U892 ( .A(G119), .B(n1184), .ZN(G21) );
NAND4_X1 U893 ( .A1(n1185), .A2(n1144), .A3(n1140), .A4(n1007), .ZN(n1184) );
AND2_X1 U894 ( .A1(n1181), .A2(n1180), .ZN(n1144) );
XNOR2_X1 U895 ( .A(n1136), .B(KEYINPUT27), .ZN(n1185) );
XNOR2_X1 U896 ( .A(G116), .B(n1186), .ZN(G18) );
NAND4_X1 U897 ( .A1(n1018), .A2(n1140), .A3(n1187), .A4(n1188), .ZN(n1186) );
XNOR2_X1 U898 ( .A(KEYINPUT56), .B(n1006), .ZN(n1188) );
INV_X1 U899 ( .A(n1135), .ZN(n1006) );
NOR2_X1 U900 ( .A1(n1183), .A2(n1189), .ZN(n1135) );
XNOR2_X1 U901 ( .A(KEYINPUT24), .B(n1024), .ZN(n1187) );
XNOR2_X1 U902 ( .A(G113), .B(n1133), .ZN(G15) );
NAND4_X1 U903 ( .A1(n1018), .A2(n1146), .A3(n1140), .A4(n1136), .ZN(n1133) );
AND2_X1 U904 ( .A1(n1003), .A2(n1176), .ZN(n1140) );
NOR2_X1 U905 ( .A1(n1190), .A2(n1011), .ZN(n1003) );
INV_X1 U906 ( .A(n1005), .ZN(n1146) );
NAND2_X1 U907 ( .A1(n1189), .A2(n1183), .ZN(n1005) );
INV_X1 U908 ( .A(n1182), .ZN(n1189) );
INV_X1 U909 ( .A(n1153), .ZN(n1018) );
NAND2_X1 U910 ( .A1(n1191), .A2(n1180), .ZN(n1153) );
XNOR2_X1 U911 ( .A(n1192), .B(n1193), .ZN(G12) );
NOR2_X1 U912 ( .A1(n1024), .A2(n1145), .ZN(n1193) );
NAND4_X1 U913 ( .A1(n1020), .A2(n1007), .A3(n1013), .A4(n1176), .ZN(n1145) );
NAND2_X1 U914 ( .A1(n1178), .A2(n1194), .ZN(n1176) );
NAND4_X1 U915 ( .A1(G953), .A2(G902), .A3(n995), .A4(n1195), .ZN(n1194) );
INV_X1 U916 ( .A(G898), .ZN(n1195) );
NAND3_X1 U917 ( .A1(n995), .A2(n992), .A3(G952), .ZN(n1178) );
NAND2_X1 U918 ( .A1(n1196), .A2(G237), .ZN(n995) );
XNOR2_X1 U919 ( .A(G234), .B(KEYINPUT25), .ZN(n1196) );
NOR2_X1 U920 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
AND2_X1 U921 ( .A1(G221), .A2(n1197), .ZN(n1011) );
INV_X1 U922 ( .A(n1190), .ZN(n1012) );
XNOR2_X1 U923 ( .A(n1198), .B(G469), .ZN(n1190) );
NAND2_X1 U924 ( .A1(KEYINPUT48), .A2(n1040), .ZN(n1198) );
INV_X1 U925 ( .A(n1047), .ZN(n1040) );
NAND2_X1 U926 ( .A1(n1199), .A2(n1200), .ZN(n1047) );
XOR2_X1 U927 ( .A(n1201), .B(n1202), .Z(n1199) );
XOR2_X1 U928 ( .A(n1203), .B(n1113), .Z(n1202) );
AND2_X1 U929 ( .A1(G227), .A2(n992), .ZN(n1113) );
NAND2_X1 U930 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NAND2_X1 U931 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
INV_X1 U932 ( .A(n1107), .ZN(n1206) );
XOR2_X1 U933 ( .A(n1208), .B(KEYINPUT55), .Z(n1204) );
NAND2_X1 U934 ( .A1(n1056), .A2(n1107), .ZN(n1208) );
XNOR2_X1 U935 ( .A(n1209), .B(n1210), .ZN(n1107) );
XNOR2_X1 U936 ( .A(n1211), .B(n1212), .ZN(n1209) );
INV_X1 U937 ( .A(n1059), .ZN(n1212) );
XOR2_X1 U938 ( .A(G143), .B(n1213), .Z(n1059) );
NAND2_X1 U939 ( .A1(KEYINPUT29), .A2(n1214), .ZN(n1211) );
NAND2_X1 U940 ( .A1(KEYINPUT53), .A2(n1112), .ZN(n1201) );
XOR2_X1 U941 ( .A(G110), .B(n1215), .Z(n1112) );
XNOR2_X1 U942 ( .A(KEYINPUT44), .B(n1058), .ZN(n1215) );
NOR2_X1 U943 ( .A1(n1182), .A2(n1183), .ZN(n1007) );
XNOR2_X1 U944 ( .A(n1216), .B(G475), .ZN(n1183) );
NAND2_X1 U945 ( .A1(n1090), .A2(n1200), .ZN(n1216) );
XNOR2_X1 U946 ( .A(n1217), .B(n1218), .ZN(n1090) );
XOR2_X1 U947 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U948 ( .A(KEYINPUT0), .B(G131), .Z(n1220) );
NOR2_X1 U949 ( .A1(KEYINPUT8), .A2(n1221), .ZN(n1219) );
XNOR2_X1 U950 ( .A(G143), .B(n1222), .ZN(n1221) );
NAND2_X1 U951 ( .A1(G214), .A2(n1223), .ZN(n1222) );
XOR2_X1 U952 ( .A(n1224), .B(n1225), .Z(n1217) );
XNOR2_X1 U953 ( .A(n1226), .B(n1227), .ZN(n1225) );
NOR2_X1 U954 ( .A1(KEYINPUT26), .A2(n1058), .ZN(n1227) );
INV_X1 U955 ( .A(G140), .ZN(n1058) );
NAND2_X1 U956 ( .A1(KEYINPUT9), .A2(n1228), .ZN(n1226) );
XOR2_X1 U957 ( .A(n1229), .B(n1230), .Z(n1228) );
XNOR2_X1 U958 ( .A(n1231), .B(KEYINPUT43), .ZN(n1230) );
NAND2_X1 U959 ( .A1(KEYINPUT40), .A2(n1214), .ZN(n1231) );
XNOR2_X1 U960 ( .A(n1232), .B(G478), .ZN(n1182) );
NAND2_X1 U961 ( .A1(n1086), .A2(n1233), .ZN(n1232) );
XNOR2_X1 U962 ( .A(KEYINPUT33), .B(n1200), .ZN(n1233) );
XOR2_X1 U963 ( .A(n1234), .B(n1235), .Z(n1086) );
XNOR2_X1 U964 ( .A(G134), .B(n1236), .ZN(n1235) );
NAND2_X1 U965 ( .A1(KEYINPUT1), .A2(n1237), .ZN(n1236) );
XOR2_X1 U966 ( .A(G128), .B(n1238), .Z(n1237) );
XOR2_X1 U967 ( .A(KEYINPUT60), .B(G143), .Z(n1238) );
XOR2_X1 U968 ( .A(n1239), .B(n1240), .Z(n1234) );
NOR2_X1 U969 ( .A1(n1241), .A2(KEYINPUT46), .ZN(n1240) );
NOR2_X1 U970 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U971 ( .A(KEYINPUT28), .B(n1244), .Z(n1243) );
NOR2_X1 U972 ( .A1(G107), .A2(n1245), .ZN(n1244) );
XNOR2_X1 U973 ( .A(n1246), .B(KEYINPUT52), .ZN(n1245) );
NOR2_X1 U974 ( .A1(n1246), .A2(n1247), .ZN(n1242) );
XNOR2_X1 U975 ( .A(n1248), .B(G122), .ZN(n1246) );
NAND2_X1 U976 ( .A1(KEYINPUT47), .A2(n1249), .ZN(n1248) );
NAND2_X1 U977 ( .A1(G217), .A2(n1250), .ZN(n1239) );
NOR2_X1 U978 ( .A1(n1180), .A2(n1191), .ZN(n1020) );
INV_X1 U979 ( .A(n1181), .ZN(n1191) );
XOR2_X1 U980 ( .A(n1034), .B(KEYINPUT23), .Z(n1181) );
XOR2_X1 U981 ( .A(n1251), .B(n1082), .Z(n1034) );
NAND2_X1 U982 ( .A1(G217), .A2(n1197), .ZN(n1082) );
NAND2_X1 U983 ( .A1(G234), .A2(n1200), .ZN(n1197) );
NAND2_X1 U984 ( .A1(n1080), .A2(n1200), .ZN(n1251) );
XNOR2_X1 U985 ( .A(n1252), .B(n1253), .ZN(n1080) );
XOR2_X1 U986 ( .A(n1254), .B(n1255), .Z(n1253) );
XNOR2_X1 U987 ( .A(G140), .B(n1256), .ZN(n1255) );
NOR2_X1 U988 ( .A1(KEYINPUT58), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U989 ( .A(n1258), .B(n1259), .ZN(n1257) );
NAND2_X1 U990 ( .A1(G221), .A2(n1250), .ZN(n1258) );
AND2_X1 U991 ( .A1(G234), .A2(n992), .ZN(n1250) );
NAND2_X1 U992 ( .A1(KEYINPUT31), .A2(G128), .ZN(n1254) );
XOR2_X1 U993 ( .A(n1224), .B(n1260), .Z(n1252) );
XNOR2_X1 U994 ( .A(G146), .B(n1060), .ZN(n1224) );
NAND2_X1 U995 ( .A1(n1261), .A2(n1262), .ZN(n1180) );
OR2_X1 U996 ( .A1(n1042), .A2(G472), .ZN(n1262) );
XOR2_X1 U997 ( .A(n1263), .B(KEYINPUT38), .Z(n1261) );
NAND2_X1 U998 ( .A1(G472), .A2(n1042), .ZN(n1263) );
NAND2_X1 U999 ( .A1(n1264), .A2(n1200), .ZN(n1042) );
XOR2_X1 U1000 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U1001 ( .A(n1267), .B(n1056), .ZN(n1266) );
INV_X1 U1002 ( .A(n1207), .ZN(n1056) );
XOR2_X1 U1003 ( .A(n1268), .B(n1269), .Z(n1207) );
INV_X1 U1004 ( .A(n1259), .ZN(n1269) );
XOR2_X1 U1005 ( .A(G137), .B(KEYINPUT17), .Z(n1259) );
XNOR2_X1 U1006 ( .A(G131), .B(G134), .ZN(n1268) );
NOR2_X1 U1007 ( .A1(KEYINPUT3), .A2(n1101), .ZN(n1267) );
XOR2_X1 U1008 ( .A(n1094), .B(n1097), .Z(n1265) );
XNOR2_X1 U1009 ( .A(n1270), .B(n1271), .ZN(n1097) );
NOR2_X1 U1010 ( .A1(KEYINPUT20), .A2(G116), .ZN(n1271) );
XNOR2_X1 U1011 ( .A(G113), .B(G119), .ZN(n1270) );
XOR2_X1 U1012 ( .A(n1272), .B(G101), .Z(n1094) );
NAND2_X1 U1013 ( .A1(G210), .A2(n1223), .ZN(n1272) );
NOR2_X1 U1014 ( .A1(G953), .A2(G237), .ZN(n1223) );
INV_X1 U1015 ( .A(n1136), .ZN(n1024) );
NOR2_X1 U1016 ( .A1(n1026), .A2(n1027), .ZN(n1136) );
NOR2_X1 U1017 ( .A1(n1273), .A2(n1043), .ZN(n1027) );
NOR2_X1 U1018 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
AND2_X1 U1019 ( .A1(n1046), .A2(n1045), .ZN(n1273) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1274), .ZN(n1045) );
AND2_X1 U1021 ( .A1(n1275), .A2(n1200), .ZN(n1046) );
XOR2_X1 U1022 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U1023 ( .A(n1075), .B(n1101), .Z(n1277) );
NAND2_X1 U1024 ( .A1(n1278), .A2(n1279), .ZN(n1101) );
OR2_X1 U1025 ( .A1(n1213), .A2(G143), .ZN(n1279) );
NAND2_X1 U1026 ( .A1(G143), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U1027 ( .A(n1213), .B(KEYINPUT51), .ZN(n1280) );
XOR2_X1 U1028 ( .A(G146), .B(G128), .Z(n1213) );
XOR2_X1 U1029 ( .A(n1281), .B(n1282), .Z(n1075) );
XOR2_X1 U1030 ( .A(n1283), .B(n1284), .Z(n1282) );
XNOR2_X1 U1031 ( .A(n1249), .B(n1210), .ZN(n1284) );
XNOR2_X1 U1032 ( .A(G101), .B(n1247), .ZN(n1210) );
INV_X1 U1033 ( .A(G107), .ZN(n1247) );
INV_X1 U1034 ( .A(G116), .ZN(n1249) );
XOR2_X1 U1035 ( .A(KEYINPUT57), .B(KEYINPUT41), .Z(n1283) );
XNOR2_X1 U1036 ( .A(n1229), .B(n1285), .ZN(n1281) );
XOR2_X1 U1037 ( .A(n1214), .B(n1260), .Z(n1285) );
XNOR2_X1 U1038 ( .A(n1192), .B(G119), .ZN(n1260) );
XOR2_X1 U1039 ( .A(G104), .B(KEYINPUT15), .Z(n1214) );
XOR2_X1 U1040 ( .A(G113), .B(G122), .Z(n1229) );
XNOR2_X1 U1041 ( .A(n1124), .B(n1286), .ZN(n1276) );
NAND2_X1 U1042 ( .A1(KEYINPUT54), .A2(n1060), .ZN(n1286) );
XOR2_X1 U1043 ( .A(G125), .B(KEYINPUT39), .Z(n1060) );
INV_X1 U1044 ( .A(n1123), .ZN(n1124) );
NAND2_X1 U1045 ( .A1(G224), .A2(n992), .ZN(n1123) );
INV_X1 U1046 ( .A(G953), .ZN(n992) );
INV_X1 U1047 ( .A(n1174), .ZN(n1026) );
NAND2_X1 U1048 ( .A1(G214), .A2(n1274), .ZN(n1174) );
NAND2_X1 U1049 ( .A1(n1287), .A2(n1200), .ZN(n1274) );
INV_X1 U1050 ( .A(G902), .ZN(n1200) );
XOR2_X1 U1051 ( .A(KEYINPUT35), .B(G237), .Z(n1287) );
INV_X1 U1052 ( .A(G110), .ZN(n1192) );
endmodule


