//Key = 0001101111110111011101001110110011100100011111011110110101010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318;

XOR2_X1 U736 ( .A(G107), .B(n1004), .Z(G9) );
NOR2_X1 U737 ( .A1(KEYINPUT1), .A2(n1005), .ZN(n1004) );
NOR2_X1 U738 ( .A1(n1006), .A2(n1007), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1008), .A2(n1009), .A3(G953), .A4(n1010), .ZN(n1007) );
NOR3_X1 U740 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1009) );
INV_X1 U741 ( .A(n1014), .ZN(n1013) );
NAND3_X1 U742 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1011) );
NAND2_X1 U743 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
NAND2_X1 U744 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND3_X1 U745 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1018) );
OR2_X1 U746 ( .A1(n1025), .A2(n1020), .ZN(n1023) );
NAND3_X1 U747 ( .A1(n1026), .A2(n1027), .A3(n1025), .ZN(n1022) );
NAND2_X1 U748 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND3_X1 U749 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1008) );
NAND4_X1 U750 ( .A1(n1020), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NAND2_X1 U751 ( .A1(n1036), .A2(n1012), .ZN(n1035) );
NAND2_X1 U752 ( .A1(KEYINPUT54), .A2(n1037), .ZN(n1036) );
NAND3_X1 U753 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1034) );
INV_X1 U754 ( .A(n1012), .ZN(n1040) );
NAND3_X1 U755 ( .A1(n1041), .A2(n1042), .A3(n1014), .ZN(n1039) );
OR2_X1 U756 ( .A1(n1016), .A2(n1017), .ZN(n1042) );
OR3_X1 U757 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1041) );
NAND2_X1 U758 ( .A1(n1037), .A2(n1046), .ZN(n1038) );
INV_X1 U759 ( .A(KEYINPUT54), .ZN(n1046) );
NOR3_X1 U760 ( .A1(n1010), .A2(G953), .A3(G952), .ZN(n1006) );
AND4_X1 U761 ( .A1(n1025), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1010) );
NOR3_X1 U762 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1049) );
XOR2_X1 U763 ( .A(n1053), .B(n1054), .Z(n1052) );
XNOR2_X1 U764 ( .A(KEYINPUT55), .B(n1055), .ZN(n1054) );
NOR2_X1 U765 ( .A1(G469), .A2(KEYINPUT56), .ZN(n1053) );
NAND4_X1 U766 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1050) );
NAND2_X1 U767 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U768 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NAND2_X1 U769 ( .A1(KEYINPUT37), .A2(n1064), .ZN(n1063) );
NAND2_X1 U770 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
NAND2_X1 U771 ( .A1(KEYINPUT37), .A2(n1067), .ZN(n1065) );
INV_X1 U772 ( .A(KEYINPUT2), .ZN(n1067) );
OR3_X1 U773 ( .A1(n1064), .A2(KEYINPUT2), .A3(n1061), .ZN(n1058) );
INV_X1 U774 ( .A(n1066), .ZN(n1064) );
NAND3_X1 U775 ( .A1(G472), .A2(n1068), .A3(n1069), .ZN(n1057) );
INV_X1 U776 ( .A(KEYINPUT39), .ZN(n1069) );
NAND2_X1 U777 ( .A1(KEYINPUT39), .A2(n1070), .ZN(n1056) );
NOR3_X1 U778 ( .A1(n1028), .A2(n1071), .A3(n1045), .ZN(n1048) );
NAND2_X1 U779 ( .A1(n1072), .A2(n1073), .ZN(n1047) );
NAND2_X1 U780 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND2_X1 U781 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U782 ( .A(KEYINPUT19), .B(G475), .Z(n1076) );
NAND2_X1 U783 ( .A1(n1078), .A2(n1070), .ZN(n1074) );
XOR2_X1 U784 ( .A(n1079), .B(n1080), .Z(G72) );
XOR2_X1 U785 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U786 ( .A1(KEYINPUT18), .A2(n1083), .ZN(n1082) );
NAND2_X1 U787 ( .A1(G953), .A2(n1084), .ZN(n1083) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1084) );
NAND2_X1 U789 ( .A1(n1085), .A2(n1086), .ZN(n1081) );
NAND2_X1 U790 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
XOR2_X1 U791 ( .A(n1089), .B(n1090), .Z(n1085) );
XOR2_X1 U792 ( .A(n1091), .B(KEYINPUT35), .Z(n1089) );
NAND2_X1 U793 ( .A1(n1092), .A2(n1093), .ZN(n1079) );
XOR2_X1 U794 ( .A(n1094), .B(n1095), .Z(G69) );
XOR2_X1 U795 ( .A(n1096), .B(n1097), .Z(n1095) );
NOR2_X1 U796 ( .A1(n1098), .A2(n1092), .ZN(n1097) );
NOR2_X1 U797 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U798 ( .A1(n1101), .A2(n1102), .ZN(n1096) );
NAND2_X1 U799 ( .A1(n1087), .A2(n1100), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1092), .A2(n1103), .ZN(n1094) );
NOR2_X1 U801 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U802 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U803 ( .A(n1108), .B(KEYINPUT6), .Z(n1107) );
NAND2_X1 U804 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U805 ( .A1(KEYINPUT41), .A2(n1111), .ZN(n1106) );
NOR2_X1 U806 ( .A1(n1104), .A2(n1112), .ZN(G63) );
XOR2_X1 U807 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U808 ( .A(KEYINPUT14), .B(n1115), .Z(n1114) );
AND2_X1 U809 ( .A1(G478), .A2(n1109), .ZN(n1115) );
NOR2_X1 U810 ( .A1(n1104), .A2(n1116), .ZN(G60) );
XOR2_X1 U811 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U812 ( .A1(n1119), .A2(KEYINPUT58), .ZN(n1118) );
NAND2_X1 U813 ( .A1(n1109), .A2(G475), .ZN(n1117) );
XOR2_X1 U814 ( .A(G104), .B(n1120), .Z(G6) );
NOR2_X1 U815 ( .A1(n1104), .A2(n1121), .ZN(G57) );
XOR2_X1 U816 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U817 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U818 ( .A1(n1070), .A2(n1126), .ZN(n1125) );
INV_X1 U819 ( .A(G472), .ZN(n1070) );
XOR2_X1 U820 ( .A(n1127), .B(KEYINPUT4), .Z(n1122) );
NAND2_X1 U821 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U822 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U823 ( .A(KEYINPUT61), .B(n1132), .Z(n1130) );
XOR2_X1 U824 ( .A(KEYINPUT32), .B(n1133), .Z(n1128) );
NOR2_X1 U825 ( .A1(n1134), .A2(n1132), .ZN(n1133) );
XOR2_X1 U826 ( .A(n1135), .B(n1136), .Z(n1132) );
XNOR2_X1 U827 ( .A(n1131), .B(KEYINPUT29), .ZN(n1134) );
NOR2_X1 U828 ( .A1(n1104), .A2(n1137), .ZN(G54) );
XOR2_X1 U829 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U830 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U831 ( .A1(n1142), .A2(KEYINPUT10), .ZN(n1140) );
XOR2_X1 U832 ( .A(n1091), .B(n1143), .Z(n1142) );
XNOR2_X1 U833 ( .A(n1144), .B(n1145), .ZN(n1138) );
AND2_X1 U834 ( .A1(G469), .A2(n1109), .ZN(n1145) );
INV_X1 U835 ( .A(n1126), .ZN(n1109) );
NOR2_X1 U836 ( .A1(n1104), .A2(n1146), .ZN(G51) );
NOR2_X1 U837 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U838 ( .A(KEYINPUT27), .B(n1149), .Z(n1148) );
AND2_X1 U839 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U840 ( .A1(n1151), .A2(n1150), .ZN(n1147) );
XNOR2_X1 U841 ( .A(n1152), .B(n1153), .ZN(n1150) );
NAND2_X1 U842 ( .A1(KEYINPUT45), .A2(n1154), .ZN(n1152) );
NOR2_X1 U843 ( .A1(n1126), .A2(n1066), .ZN(n1151) );
NAND2_X1 U844 ( .A1(G902), .A2(n1155), .ZN(n1126) );
NAND2_X1 U845 ( .A1(n1032), .A2(n1030), .ZN(n1155) );
INV_X1 U846 ( .A(n1093), .ZN(n1030) );
NAND4_X1 U847 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1093) );
AND4_X1 U848 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1159) );
AND2_X1 U849 ( .A1(n1164), .A2(n1165), .ZN(n1158) );
NAND3_X1 U850 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1156) );
XNOR2_X1 U851 ( .A(n1169), .B(KEYINPUT5), .ZN(n1168) );
INV_X1 U852 ( .A(n1170), .ZN(n1167) );
XNOR2_X1 U853 ( .A(n1171), .B(KEYINPUT13), .ZN(n1166) );
INV_X1 U854 ( .A(n1103), .ZN(n1032) );
NAND4_X1 U855 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1103) );
NOR4_X1 U856 ( .A1(n1120), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1175) );
NOR2_X1 U857 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
INV_X1 U858 ( .A(n1181), .ZN(n1177) );
INV_X1 U859 ( .A(n1005), .ZN(n1176) );
NAND2_X1 U860 ( .A1(n1043), .A2(n1182), .ZN(n1005) );
AND2_X1 U861 ( .A1(n1044), .A2(n1182), .ZN(n1120) );
AND4_X1 U862 ( .A1(n1183), .A2(n1033), .A3(n1171), .A4(n1184), .ZN(n1182) );
NOR2_X1 U863 ( .A1(n1185), .A2(n1186), .ZN(n1174) );
NOR2_X1 U864 ( .A1(n1092), .A2(G952), .ZN(n1104) );
XOR2_X1 U865 ( .A(G146), .B(n1187), .Z(G48) );
NOR2_X1 U866 ( .A1(KEYINPUT0), .A2(n1157), .ZN(n1187) );
NAND3_X1 U867 ( .A1(n1044), .A2(n1171), .A3(n1188), .ZN(n1157) );
XOR2_X1 U868 ( .A(G143), .B(n1189), .Z(G45) );
NOR4_X1 U869 ( .A1(KEYINPUT38), .A2(n1169), .A3(n1027), .A4(n1170), .ZN(n1189) );
NAND4_X1 U870 ( .A1(n1021), .A2(n1183), .A3(n1051), .A4(n1190), .ZN(n1170) );
INV_X1 U871 ( .A(n1171), .ZN(n1027) );
XNOR2_X1 U872 ( .A(G140), .B(n1165), .ZN(G42) );
NAND2_X1 U873 ( .A1(n1191), .A2(n1192), .ZN(n1165) );
XNOR2_X1 U874 ( .A(G137), .B(n1160), .ZN(G39) );
NAND3_X1 U875 ( .A1(n1020), .A2(n1017), .A3(n1188), .ZN(n1160) );
XNOR2_X1 U876 ( .A(G134), .B(n1164), .ZN(G36) );
NAND3_X1 U877 ( .A1(n1021), .A2(n1043), .A3(n1191), .ZN(n1164) );
XOR2_X1 U878 ( .A(n1193), .B(G131), .Z(G33) );
NAND2_X1 U879 ( .A1(KEYINPUT52), .A2(n1163), .ZN(n1193) );
NAND3_X1 U880 ( .A1(n1044), .A2(n1021), .A3(n1191), .ZN(n1163) );
AND3_X1 U881 ( .A1(n1183), .A2(n1194), .A3(n1020), .ZN(n1191) );
NOR2_X1 U882 ( .A1(n1195), .A2(n1028), .ZN(n1020) );
XOR2_X1 U883 ( .A(n1162), .B(n1196), .Z(G30) );
XOR2_X1 U884 ( .A(KEYINPUT7), .B(G128), .Z(n1196) );
NAND3_X1 U885 ( .A1(n1043), .A2(n1171), .A3(n1188), .ZN(n1162) );
AND4_X1 U886 ( .A1(n1183), .A2(n1197), .A3(n1194), .A4(n1198), .ZN(n1188) );
XOR2_X1 U887 ( .A(G101), .B(n1199), .Z(G3) );
NOR2_X1 U888 ( .A1(n1179), .A2(n1200), .ZN(n1199) );
XNOR2_X1 U889 ( .A(KEYINPUT43), .B(n1180), .ZN(n1200) );
INV_X1 U890 ( .A(n1021), .ZN(n1180) );
XNOR2_X1 U891 ( .A(G125), .B(n1161), .ZN(G27) );
NAND4_X1 U892 ( .A1(n1014), .A2(n1192), .A3(n1201), .A4(n1171), .ZN(n1161) );
NOR2_X1 U893 ( .A1(n1045), .A2(n1169), .ZN(n1201) );
INV_X1 U894 ( .A(n1194), .ZN(n1169) );
NAND2_X1 U895 ( .A1(n1012), .A2(n1202), .ZN(n1194) );
NAND2_X1 U896 ( .A1(n1203), .A2(n1088), .ZN(n1202) );
INV_X1 U897 ( .A(G900), .ZN(n1088) );
NOR3_X1 U898 ( .A1(n1198), .A2(n1025), .A3(n1204), .ZN(n1192) );
NAND2_X1 U899 ( .A1(n1205), .A2(n1206), .ZN(G24) );
NAND2_X1 U900 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U901 ( .A(KEYINPUT34), .B(n1209), .Z(n1205) );
NOR2_X1 U902 ( .A1(n1207), .A2(n1208), .ZN(n1209) );
INV_X1 U903 ( .A(n1172), .ZN(n1207) );
NAND4_X1 U904 ( .A1(n1210), .A2(n1033), .A3(n1051), .A4(n1190), .ZN(n1172) );
NOR2_X1 U905 ( .A1(n1198), .A2(n1197), .ZN(n1033) );
XNOR2_X1 U906 ( .A(G119), .B(n1211), .ZN(G21) );
NAND2_X1 U907 ( .A1(KEYINPUT28), .A2(n1212), .ZN(n1211) );
INV_X1 U908 ( .A(n1173), .ZN(n1212) );
NAND4_X1 U909 ( .A1(n1210), .A2(n1017), .A3(n1197), .A4(n1198), .ZN(n1173) );
NAND2_X1 U910 ( .A1(n1213), .A2(n1214), .ZN(G18) );
NAND2_X1 U911 ( .A1(G116), .A2(n1181), .ZN(n1214) );
XOR2_X1 U912 ( .A(KEYINPUT44), .B(n1215), .Z(n1213) );
NOR2_X1 U913 ( .A1(G116), .A2(n1181), .ZN(n1215) );
NAND3_X1 U914 ( .A1(n1021), .A2(n1043), .A3(n1210), .ZN(n1181) );
NOR2_X1 U915 ( .A1(n1190), .A2(n1216), .ZN(n1043) );
XNOR2_X1 U916 ( .A(n1217), .B(n1186), .ZN(G15) );
AND3_X1 U917 ( .A1(n1210), .A2(n1021), .A3(n1044), .ZN(n1186) );
INV_X1 U918 ( .A(n1204), .ZN(n1044) );
NAND2_X1 U919 ( .A1(n1216), .A2(n1190), .ZN(n1204) );
INV_X1 U920 ( .A(n1051), .ZN(n1216) );
NOR2_X1 U921 ( .A1(n1197), .A2(n1024), .ZN(n1021) );
INV_X1 U922 ( .A(n1198), .ZN(n1024) );
AND4_X1 U923 ( .A1(n1014), .A2(n1171), .A3(n1184), .A4(n1016), .ZN(n1210) );
NAND2_X1 U924 ( .A1(n1218), .A2(n1219), .ZN(G12) );
NAND3_X1 U925 ( .A1(n1185), .A2(KEYINPUT3), .A3(n1220), .ZN(n1219) );
INV_X1 U926 ( .A(n1221), .ZN(n1220) );
NAND2_X1 U927 ( .A1(n1221), .A2(n1222), .ZN(n1218) );
NAND2_X1 U928 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NAND2_X1 U929 ( .A1(n1185), .A2(n1225), .ZN(n1224) );
NAND2_X1 U930 ( .A1(KEYINPUT3), .A2(n1226), .ZN(n1225) );
NAND2_X1 U931 ( .A1(n1226), .A2(n1227), .ZN(n1223) );
INV_X1 U932 ( .A(n1185), .ZN(n1227) );
NOR3_X1 U933 ( .A1(n1198), .A2(n1025), .A3(n1179), .ZN(n1185) );
NAND3_X1 U934 ( .A1(n1171), .A2(n1184), .A3(n1037), .ZN(n1179) );
AND2_X1 U935 ( .A1(n1017), .A2(n1183), .ZN(n1037) );
NOR2_X1 U936 ( .A1(n1014), .A2(n1045), .ZN(n1183) );
INV_X1 U937 ( .A(n1016), .ZN(n1045) );
NAND2_X1 U938 ( .A1(G221), .A2(n1228), .ZN(n1016) );
XOR2_X1 U939 ( .A(n1055), .B(G469), .Z(n1014) );
NAND2_X1 U940 ( .A1(n1229), .A2(n1073), .ZN(n1055) );
XOR2_X1 U941 ( .A(n1141), .B(n1230), .Z(n1229) );
XNOR2_X1 U942 ( .A(n1091), .B(n1231), .ZN(n1230) );
INV_X1 U943 ( .A(n1232), .ZN(n1231) );
XOR2_X1 U944 ( .A(n1233), .B(n1234), .Z(n1091) );
XOR2_X1 U945 ( .A(n1235), .B(n1236), .Z(n1234) );
XOR2_X1 U946 ( .A(KEYINPUT26), .B(KEYINPUT22), .Z(n1236) );
NOR2_X1 U947 ( .A1(G128), .A2(KEYINPUT46), .ZN(n1235) );
XOR2_X1 U948 ( .A(n1136), .B(n1237), .Z(n1233) );
XOR2_X1 U949 ( .A(n1238), .B(n1239), .Z(n1141) );
XOR2_X1 U950 ( .A(KEYINPUT53), .B(G140), .Z(n1239) );
NAND2_X1 U951 ( .A1(G227), .A2(n1092), .ZN(n1238) );
NOR2_X1 U952 ( .A1(n1051), .A2(n1190), .ZN(n1017) );
NAND2_X1 U953 ( .A1(n1240), .A2(n1241), .ZN(n1190) );
OR3_X1 U954 ( .A1(G475), .A2(G902), .A3(n1119), .ZN(n1241) );
INV_X1 U955 ( .A(n1077), .ZN(n1119) );
XOR2_X1 U956 ( .A(KEYINPUT50), .B(n1071), .Z(n1240) );
AND2_X1 U957 ( .A1(G475), .A2(n1242), .ZN(n1071) );
NAND2_X1 U958 ( .A1(n1073), .A2(n1077), .ZN(n1242) );
NAND2_X1 U959 ( .A1(n1243), .A2(n1244), .ZN(n1077) );
NAND2_X1 U960 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U961 ( .A(KEYINPUT47), .B(n1247), .Z(n1243) );
NOR2_X1 U962 ( .A1(n1246), .A2(n1245), .ZN(n1247) );
XOR2_X1 U963 ( .A(n1248), .B(n1249), .Z(n1245) );
XOR2_X1 U964 ( .A(n1250), .B(n1251), .Z(n1249) );
NOR2_X1 U965 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U966 ( .A(G214), .ZN(n1253) );
XNOR2_X1 U967 ( .A(G131), .B(G143), .ZN(n1250) );
NAND2_X1 U968 ( .A1(n1254), .A2(KEYINPUT11), .ZN(n1248) );
XNOR2_X1 U969 ( .A(G146), .B(n1090), .ZN(n1254) );
XOR2_X1 U970 ( .A(G125), .B(G140), .Z(n1090) );
XNOR2_X1 U971 ( .A(n1255), .B(G104), .ZN(n1246) );
NAND2_X1 U972 ( .A1(KEYINPUT8), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U973 ( .A(n1257), .B(G478), .ZN(n1051) );
NAND2_X1 U974 ( .A1(n1258), .A2(n1073), .ZN(n1257) );
XOR2_X1 U975 ( .A(KEYINPUT23), .B(n1113), .Z(n1258) );
XNOR2_X1 U976 ( .A(n1259), .B(n1260), .ZN(n1113) );
XNOR2_X1 U977 ( .A(n1261), .B(n1262), .ZN(n1260) );
NAND3_X1 U978 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1261) );
OR2_X1 U979 ( .A1(n1208), .A2(G116), .ZN(n1265) );
NAND2_X1 U980 ( .A1(n1266), .A2(n1267), .ZN(n1264) );
INV_X1 U981 ( .A(KEYINPUT49), .ZN(n1267) );
NAND2_X1 U982 ( .A1(n1268), .A2(n1208), .ZN(n1266) );
XNOR2_X1 U983 ( .A(KEYINPUT21), .B(G116), .ZN(n1268) );
NAND2_X1 U984 ( .A1(KEYINPUT49), .A2(n1269), .ZN(n1263) );
NAND2_X1 U985 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
OR2_X1 U986 ( .A1(G116), .A2(KEYINPUT21), .ZN(n1271) );
NAND3_X1 U987 ( .A1(G116), .A2(n1208), .A3(KEYINPUT21), .ZN(n1270) );
INV_X1 U988 ( .A(G122), .ZN(n1208) );
XOR2_X1 U989 ( .A(n1272), .B(n1273), .Z(n1259) );
NOR2_X1 U990 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U991 ( .A(n1276), .B(KEYINPUT62), .Z(n1275) );
NAND2_X1 U992 ( .A1(G134), .A2(n1277), .ZN(n1276) );
NOR2_X1 U993 ( .A1(G134), .A2(n1277), .ZN(n1274) );
XOR2_X1 U994 ( .A(G143), .B(G128), .Z(n1277) );
NAND3_X1 U995 ( .A1(KEYINPUT15), .A2(n1278), .A3(n1279), .ZN(n1272) );
XNOR2_X1 U996 ( .A(G217), .B(KEYINPUT17), .ZN(n1279) );
NAND2_X1 U997 ( .A1(n1012), .A2(n1280), .ZN(n1184) );
NAND2_X1 U998 ( .A1(n1203), .A2(n1100), .ZN(n1280) );
INV_X1 U999 ( .A(G898), .ZN(n1100) );
AND3_X1 U1000 ( .A1(n1087), .A2(n1281), .A3(G902), .ZN(n1203) );
XNOR2_X1 U1001 ( .A(G953), .B(KEYINPUT48), .ZN(n1087) );
NAND3_X1 U1002 ( .A1(n1281), .A2(n1092), .A3(G952), .ZN(n1012) );
NAND2_X1 U1003 ( .A1(G234), .A2(G237), .ZN(n1281) );
NOR2_X1 U1004 ( .A1(n1029), .A2(n1028), .ZN(n1171) );
AND2_X1 U1005 ( .A1(G214), .A2(n1282), .ZN(n1028) );
INV_X1 U1006 ( .A(n1195), .ZN(n1029) );
XOR2_X1 U1007 ( .A(n1061), .B(n1066), .Z(n1195) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1282), .ZN(n1066) );
NAND2_X1 U1009 ( .A1(n1283), .A2(n1073), .ZN(n1282) );
NAND2_X1 U1010 ( .A1(n1284), .A2(n1073), .ZN(n1061) );
XNOR2_X1 U1011 ( .A(n1153), .B(n1154), .ZN(n1284) );
XNOR2_X1 U1012 ( .A(n1285), .B(n1286), .ZN(n1153) );
XOR2_X1 U1013 ( .A(KEYINPUT20), .B(G125), .Z(n1286) );
XNOR2_X1 U1014 ( .A(n1101), .B(n1287), .ZN(n1285) );
NOR2_X1 U1015 ( .A1(G953), .A2(n1099), .ZN(n1287) );
INV_X1 U1016 ( .A(G224), .ZN(n1099) );
XOR2_X1 U1017 ( .A(n1288), .B(n1289), .Z(n1101) );
XNOR2_X1 U1018 ( .A(n1232), .B(n1256), .ZN(n1288) );
XNOR2_X1 U1019 ( .A(n1217), .B(G122), .ZN(n1256) );
INV_X1 U1020 ( .A(G113), .ZN(n1217) );
XOR2_X1 U1021 ( .A(G110), .B(n1143), .Z(n1232) );
XNOR2_X1 U1022 ( .A(n1290), .B(n1262), .ZN(n1143) );
XOR2_X1 U1023 ( .A(G107), .B(KEYINPUT25), .Z(n1262) );
XNOR2_X1 U1024 ( .A(G101), .B(G104), .ZN(n1290) );
INV_X1 U1025 ( .A(n1197), .ZN(n1025) );
XNOR2_X1 U1026 ( .A(n1291), .B(n1110), .ZN(n1197) );
AND2_X1 U1027 ( .A1(G217), .A2(n1228), .ZN(n1110) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1073), .ZN(n1228) );
NAND2_X1 U1029 ( .A1(n1111), .A2(n1073), .ZN(n1291) );
XNOR2_X1 U1030 ( .A(n1292), .B(n1293), .ZN(n1111) );
XOR2_X1 U1031 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1032 ( .A(G125), .B(n1144), .ZN(n1295) );
INV_X1 U1033 ( .A(G110), .ZN(n1144) );
XOR2_X1 U1034 ( .A(G146), .B(G137), .Z(n1294) );
XOR2_X1 U1035 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U1036 ( .A(n1298), .B(n1299), .Z(n1297) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1278), .ZN(n1299) );
AND2_X1 U1038 ( .A1(G234), .A2(n1092), .ZN(n1278) );
NAND2_X1 U1039 ( .A1(n1300), .A2(KEYINPUT24), .ZN(n1298) );
XOR2_X1 U1040 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U1041 ( .A(G128), .B(KEYINPUT57), .ZN(n1301) );
NAND2_X1 U1042 ( .A1(KEYINPUT59), .A2(G140), .ZN(n1296) );
NAND2_X1 U1043 ( .A1(n1303), .A2(n1304), .ZN(n1198) );
NAND2_X1 U1044 ( .A1(G472), .A2(n1068), .ZN(n1304) );
XOR2_X1 U1045 ( .A(KEYINPUT42), .B(n1305), .Z(n1303) );
NOR2_X1 U1046 ( .A1(G472), .A2(n1068), .ZN(n1305) );
NAND2_X1 U1047 ( .A1(n1073), .A2(n1078), .ZN(n1068) );
NAND2_X1 U1048 ( .A1(n1306), .A2(n1307), .ZN(n1078) );
NAND2_X1 U1049 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XOR2_X1 U1050 ( .A(KEYINPUT63), .B(n1310), .Z(n1306) );
NOR2_X1 U1051 ( .A1(n1308), .A2(n1309), .ZN(n1310) );
XNOR2_X1 U1052 ( .A(n1311), .B(n1131), .ZN(n1309) );
XOR2_X1 U1053 ( .A(G113), .B(n1312), .Z(n1131) );
NOR2_X1 U1054 ( .A1(KEYINPUT16), .A2(n1289), .ZN(n1312) );
XNOR2_X1 U1055 ( .A(G116), .B(n1302), .ZN(n1289) );
XOR2_X1 U1056 ( .A(G119), .B(KEYINPUT51), .Z(n1302) );
NAND2_X1 U1057 ( .A1(n1313), .A2(KEYINPUT9), .ZN(n1311) );
XOR2_X1 U1058 ( .A(n1135), .B(n1314), .Z(n1313) );
NOR2_X1 U1059 ( .A1(KEYINPUT30), .A2(n1136), .ZN(n1314) );
XNOR2_X1 U1060 ( .A(G131), .B(n1315), .ZN(n1136) );
XOR2_X1 U1061 ( .A(G137), .B(G134), .Z(n1315) );
XNOR2_X1 U1062 ( .A(n1154), .B(KEYINPUT40), .ZN(n1135) );
XOR2_X1 U1063 ( .A(G128), .B(n1237), .Z(n1154) );
XOR2_X1 U1064 ( .A(G143), .B(G146), .Z(n1237) );
XNOR2_X1 U1065 ( .A(n1124), .B(KEYINPUT31), .ZN(n1308) );
XNOR2_X1 U1066 ( .A(G101), .B(n1316), .ZN(n1124) );
NOR2_X1 U1067 ( .A1(n1252), .A2(n1317), .ZN(n1316) );
INV_X1 U1068 ( .A(G210), .ZN(n1317) );
NAND2_X1 U1069 ( .A1(n1318), .A2(n1092), .ZN(n1252) );
INV_X1 U1070 ( .A(G953), .ZN(n1092) );
XNOR2_X1 U1071 ( .A(KEYINPUT33), .B(n1283), .ZN(n1318) );
INV_X1 U1072 ( .A(G237), .ZN(n1283) );
INV_X1 U1073 ( .A(G902), .ZN(n1073) );
XNOR2_X1 U1074 ( .A(KEYINPUT60), .B(KEYINPUT36), .ZN(n1226) );
XOR2_X1 U1075 ( .A(G110), .B(KEYINPUT12), .Z(n1221) );
endmodule


