//Key = 1100100010100101000001110000010101000011111011111100001001011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;

NAND2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(G9) );
NAND2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XNOR2_X1 U796 ( .A(KEYINPUT28), .B(n1115), .ZN(n1113) );
NAND2_X1 U797 ( .A1(n1116), .A2(G107), .ZN(n1111) );
XNOR2_X1 U798 ( .A(KEYINPUT0), .B(n1115), .ZN(n1116) );
NOR2_X1 U799 ( .A1(n1117), .A2(n1118), .ZN(G75) );
NOR4_X1 U800 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
XOR2_X1 U802 ( .A(KEYINPUT22), .B(n1125), .Z(n1124) );
NAND4_X1 U803 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1119) );
NAND3_X1 U804 ( .A1(n1130), .A2(n1125), .A3(n1131), .ZN(n1127) );
AND3_X1 U805 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1125) );
NAND2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U808 ( .A1(n1134), .A2(n1139), .ZN(n1138) );
NAND2_X1 U809 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NAND2_X1 U810 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XNOR2_X1 U811 ( .A(KEYINPUT24), .B(n1144), .ZN(n1143) );
NAND2_X1 U812 ( .A1(n1132), .A2(n1145), .ZN(n1140) );
OR2_X1 U813 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U814 ( .A1(n1133), .A2(n1148), .ZN(n1137) );
NAND2_X1 U815 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND3_X1 U816 ( .A1(n1151), .A2(n1152), .A3(n1134), .ZN(n1150) );
NOR2_X1 U817 ( .A1(n1153), .A2(n1154), .ZN(n1134) );
INV_X1 U818 ( .A(n1155), .ZN(n1154) );
NAND2_X1 U819 ( .A1(n1132), .A2(n1156), .ZN(n1149) );
NAND2_X1 U820 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U821 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U822 ( .A(KEYINPUT63), .B(n1153), .ZN(n1160) );
NAND2_X1 U823 ( .A1(n1161), .A2(n1162), .ZN(n1157) );
XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n1153), .ZN(n1162) );
AND3_X1 U825 ( .A1(n1128), .A2(n1129), .A3(n1163), .ZN(n1117) );
NAND4_X1 U826 ( .A1(n1151), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1128) );
NOR4_X1 U827 ( .A1(n1131), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1166) );
XOR2_X1 U828 ( .A(n1170), .B(KEYINPUT21), .Z(n1169) );
XOR2_X1 U829 ( .A(n1171), .B(n1172), .Z(n1168) );
XOR2_X1 U830 ( .A(KEYINPUT60), .B(G472), .Z(n1172) );
AND2_X1 U831 ( .A1(n1173), .A2(n1174), .ZN(n1167) );
NOR3_X1 U832 ( .A1(n1144), .A2(n1175), .A3(n1176), .ZN(n1165) );
NOR2_X1 U833 ( .A1(KEYINPUT19), .A2(n1177), .ZN(n1176) );
NOR2_X1 U834 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
AND2_X1 U835 ( .A1(n1174), .A2(KEYINPUT3), .ZN(n1179) );
NOR3_X1 U836 ( .A1(KEYINPUT3), .A2(n1174), .A3(n1173), .ZN(n1178) );
INV_X1 U837 ( .A(n1180), .ZN(n1174) );
NOR2_X1 U838 ( .A1(n1181), .A2(n1182), .ZN(n1175) );
INV_X1 U839 ( .A(KEYINPUT19), .ZN(n1182) );
NOR2_X1 U840 ( .A1(n1173), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U841 ( .A(KEYINPUT3), .B(n1180), .ZN(n1183) );
XOR2_X1 U842 ( .A(n1184), .B(n1185), .Z(G72) );
NOR2_X1 U843 ( .A1(n1186), .A2(n1129), .ZN(n1185) );
NOR2_X1 U844 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U845 ( .A1(n1189), .A2(n1190), .ZN(n1184) );
NAND2_X1 U846 ( .A1(n1191), .A2(n1129), .ZN(n1190) );
XOR2_X1 U847 ( .A(n1122), .B(n1192), .Z(n1191) );
NAND3_X1 U848 ( .A1(G900), .A2(n1192), .A3(G953), .ZN(n1189) );
XOR2_X1 U849 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U850 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U851 ( .A(G140), .B(KEYINPUT10), .ZN(n1196) );
NAND2_X1 U852 ( .A1(KEYINPUT39), .A2(n1197), .ZN(n1195) );
XOR2_X1 U853 ( .A(n1198), .B(n1199), .Z(n1193) );
XNOR2_X1 U854 ( .A(n1200), .B(n1201), .ZN(n1198) );
NAND2_X1 U855 ( .A1(KEYINPUT13), .A2(n1202), .ZN(n1201) );
NAND2_X1 U856 ( .A1(n1203), .A2(KEYINPUT48), .ZN(n1200) );
XNOR2_X1 U857 ( .A(G125), .B(KEYINPUT40), .ZN(n1203) );
NAND2_X1 U858 ( .A1(n1204), .A2(n1205), .ZN(G69) );
NAND2_X1 U859 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U860 ( .A1(G953), .A2(n1208), .ZN(n1206) );
NAND2_X1 U861 ( .A1(G898), .A2(G224), .ZN(n1208) );
NAND2_X1 U862 ( .A1(n1209), .A2(n1210), .ZN(n1204) );
NAND2_X1 U863 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
OR2_X1 U864 ( .A1(n1129), .A2(G224), .ZN(n1212) );
INV_X1 U865 ( .A(n1207), .ZN(n1209) );
NAND3_X1 U866 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1207) );
NAND3_X1 U867 ( .A1(n1120), .A2(n1129), .A3(n1216), .ZN(n1215) );
NAND2_X1 U868 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U869 ( .A1(KEYINPUT42), .A2(n1219), .ZN(n1218) );
NAND2_X1 U870 ( .A1(KEYINPUT18), .A2(n1219), .ZN(n1214) );
NAND3_X1 U871 ( .A1(n1220), .A2(n1217), .A3(n1221), .ZN(n1213) );
INV_X1 U872 ( .A(n1219), .ZN(n1221) );
NAND3_X1 U873 ( .A1(n1222), .A2(n1223), .A3(n1211), .ZN(n1219) );
INV_X1 U874 ( .A(n1224), .ZN(n1211) );
NAND2_X1 U875 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
XOR2_X1 U876 ( .A(KEYINPUT55), .B(n1227), .Z(n1225) );
NAND2_X1 U877 ( .A1(n1228), .A2(n1229), .ZN(n1222) );
XNOR2_X1 U878 ( .A(n1227), .B(KEYINPUT50), .ZN(n1229) );
INV_X1 U879 ( .A(KEYINPUT18), .ZN(n1217) );
NAND2_X1 U880 ( .A1(KEYINPUT42), .A2(n1120), .ZN(n1220) );
NOR2_X1 U881 ( .A1(n1230), .A2(n1231), .ZN(G66) );
NOR2_X1 U882 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
XOR2_X1 U883 ( .A(KEYINPUT6), .B(n1234), .Z(n1233) );
NOR2_X1 U884 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
AND2_X1 U885 ( .A1(n1236), .A2(n1235), .ZN(n1232) );
NAND2_X1 U886 ( .A1(n1237), .A2(G217), .ZN(n1236) );
NOR2_X1 U887 ( .A1(n1230), .A2(n1238), .ZN(G63) );
XOR2_X1 U888 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U889 ( .A1(n1237), .A2(G478), .ZN(n1239) );
NOR2_X1 U890 ( .A1(n1230), .A2(n1241), .ZN(G60) );
XOR2_X1 U891 ( .A(n1242), .B(n1243), .Z(n1241) );
NAND2_X1 U892 ( .A1(n1237), .A2(G475), .ZN(n1242) );
XNOR2_X1 U893 ( .A(n1244), .B(n1245), .ZN(G6) );
NAND2_X1 U894 ( .A1(KEYINPUT1), .A2(n1246), .ZN(n1245) );
XOR2_X1 U895 ( .A(KEYINPUT34), .B(G104), .Z(n1246) );
NOR2_X1 U896 ( .A1(n1247), .A2(n1248), .ZN(G57) );
XOR2_X1 U897 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U898 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U899 ( .A(n1253), .B(n1254), .Z(n1252) );
NAND2_X1 U900 ( .A1(KEYINPUT45), .A2(n1255), .ZN(n1253) );
XOR2_X1 U901 ( .A(n1256), .B(n1257), .Z(n1249) );
XOR2_X1 U902 ( .A(n1258), .B(KEYINPUT46), .Z(n1257) );
NAND2_X1 U903 ( .A1(n1237), .A2(G472), .ZN(n1256) );
NOR2_X1 U904 ( .A1(n1259), .A2(n1260), .ZN(n1247) );
XNOR2_X1 U905 ( .A(KEYINPUT4), .B(n1129), .ZN(n1260) );
XNOR2_X1 U906 ( .A(G952), .B(KEYINPUT38), .ZN(n1259) );
NOR2_X1 U907 ( .A1(n1230), .A2(n1261), .ZN(G54) );
XOR2_X1 U908 ( .A(n1262), .B(n1263), .Z(n1261) );
XNOR2_X1 U909 ( .A(n1264), .B(n1265), .ZN(n1263) );
NAND2_X1 U910 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U911 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
INV_X1 U912 ( .A(n1270), .ZN(n1269) );
NAND2_X1 U913 ( .A1(n1270), .A2(n1271), .ZN(n1266) );
XNOR2_X1 U914 ( .A(n1268), .B(KEYINPUT5), .ZN(n1271) );
XOR2_X1 U915 ( .A(n1272), .B(n1273), .Z(n1262) );
NAND2_X1 U916 ( .A1(n1237), .A2(G469), .ZN(n1272) );
INV_X1 U917 ( .A(n1274), .ZN(n1237) );
NOR2_X1 U918 ( .A1(n1230), .A2(n1275), .ZN(G51) );
XOR2_X1 U919 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U920 ( .A(n1278), .B(n1279), .ZN(n1277) );
NOR2_X1 U921 ( .A1(KEYINPUT11), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U922 ( .A(n1281), .B(n1282), .ZN(n1276) );
NOR2_X1 U923 ( .A1(KEYINPUT53), .A2(n1283), .ZN(n1282) );
NOR2_X1 U924 ( .A1(KEYINPUT51), .A2(n1284), .ZN(n1281) );
NOR2_X1 U925 ( .A1(n1180), .A2(n1274), .ZN(n1284) );
NAND2_X1 U926 ( .A1(G902), .A2(n1285), .ZN(n1274) );
OR2_X1 U927 ( .A1(n1120), .A2(n1122), .ZN(n1285) );
NAND4_X1 U928 ( .A1(n1286), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n1122) );
AND3_X1 U929 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1289) );
NAND2_X1 U930 ( .A1(n1293), .A2(n1294), .ZN(n1288) );
NAND3_X1 U931 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
NAND4_X1 U932 ( .A1(n1146), .A2(n1132), .A3(n1161), .A4(n1298), .ZN(n1295) );
NAND4_X1 U933 ( .A1(n1299), .A2(n1115), .A3(n1300), .A4(n1301), .ZN(n1120) );
NOR4_X1 U934 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1244), .ZN(n1301) );
AND3_X1 U935 ( .A1(n1305), .A2(n1155), .A3(n1146), .ZN(n1244) );
NAND2_X1 U936 ( .A1(n1306), .A2(n1307), .ZN(n1300) );
NAND2_X1 U937 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND2_X1 U938 ( .A1(n1133), .A2(n1310), .ZN(n1309) );
NAND2_X1 U939 ( .A1(n1159), .A2(n1147), .ZN(n1308) );
NAND3_X1 U940 ( .A1(n1147), .A2(n1155), .A3(n1305), .ZN(n1115) );
AND2_X1 U941 ( .A1(n1311), .A2(n1163), .ZN(n1230) );
INV_X1 U942 ( .A(G952), .ZN(n1163) );
XNOR2_X1 U943 ( .A(KEYINPUT4), .B(G953), .ZN(n1311) );
XNOR2_X1 U944 ( .A(G146), .B(n1286), .ZN(G48) );
NAND4_X1 U945 ( .A1(n1312), .A2(n1146), .A3(n1293), .A4(n1310), .ZN(n1286) );
XNOR2_X1 U946 ( .A(n1313), .B(n1314), .ZN(G45) );
NOR2_X1 U947 ( .A1(n1297), .A2(n1315), .ZN(n1314) );
XNOR2_X1 U948 ( .A(KEYINPUT54), .B(n1123), .ZN(n1315) );
NAND4_X1 U949 ( .A1(n1312), .A2(n1159), .A3(n1316), .A4(n1317), .ZN(n1297) );
XNOR2_X1 U950 ( .A(G140), .B(n1287), .ZN(G42) );
NAND3_X1 U951 ( .A1(n1146), .A2(n1161), .A3(n1318), .ZN(n1287) );
XNOR2_X1 U952 ( .A(G137), .B(n1290), .ZN(G39) );
NAND3_X1 U953 ( .A1(n1133), .A2(n1310), .A3(n1318), .ZN(n1290) );
XOR2_X1 U954 ( .A(n1292), .B(n1319), .Z(G36) );
NOR2_X1 U955 ( .A1(G134), .A2(KEYINPUT35), .ZN(n1319) );
NAND3_X1 U956 ( .A1(n1159), .A2(n1147), .A3(n1318), .ZN(n1292) );
XNOR2_X1 U957 ( .A(G131), .B(n1291), .ZN(G33) );
NAND3_X1 U958 ( .A1(n1146), .A2(n1159), .A3(n1318), .ZN(n1291) );
AND2_X1 U959 ( .A1(n1312), .A2(n1135), .ZN(n1318) );
NOR2_X1 U960 ( .A1(n1320), .A2(n1131), .ZN(n1135) );
NAND3_X1 U961 ( .A1(n1321), .A2(n1322), .A3(n1323), .ZN(G30) );
OR2_X1 U962 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND3_X1 U963 ( .A1(n1325), .A2(n1324), .A3(G128), .ZN(n1322) );
NAND2_X1 U964 ( .A1(n1326), .A2(n1327), .ZN(n1321) );
NAND2_X1 U965 ( .A1(n1328), .A2(n1324), .ZN(n1326) );
INV_X1 U966 ( .A(KEYINPUT30), .ZN(n1324) );
XNOR2_X1 U967 ( .A(KEYINPUT62), .B(n1325), .ZN(n1328) );
NAND2_X1 U968 ( .A1(n1293), .A2(n1329), .ZN(n1325) );
XNOR2_X1 U969 ( .A(KEYINPUT37), .B(n1296), .ZN(n1329) );
NAND3_X1 U970 ( .A1(n1147), .A2(n1310), .A3(n1312), .ZN(n1296) );
AND2_X1 U971 ( .A1(n1142), .A2(n1298), .ZN(n1312) );
XNOR2_X1 U972 ( .A(n1255), .B(n1304), .ZN(G3) );
AND3_X1 U973 ( .A1(n1133), .A2(n1305), .A3(n1159), .ZN(n1304) );
INV_X1 U974 ( .A(n1330), .ZN(n1159) );
XNOR2_X1 U975 ( .A(G125), .B(n1331), .ZN(G27) );
NAND4_X1 U976 ( .A1(n1332), .A2(n1132), .A3(n1333), .A4(n1161), .ZN(n1331) );
AND2_X1 U977 ( .A1(n1298), .A2(n1293), .ZN(n1333) );
NAND2_X1 U978 ( .A1(n1153), .A2(n1334), .ZN(n1298) );
NAND4_X1 U979 ( .A1(G902), .A2(G953), .A3(n1335), .A4(n1188), .ZN(n1334) );
INV_X1 U980 ( .A(G900), .ZN(n1188) );
XNOR2_X1 U981 ( .A(n1146), .B(KEYINPUT31), .ZN(n1332) );
INV_X1 U982 ( .A(n1336), .ZN(n1146) );
XOR2_X1 U983 ( .A(n1299), .B(n1337), .Z(G24) );
NOR2_X1 U984 ( .A1(G122), .A2(KEYINPUT2), .ZN(n1337) );
NAND4_X1 U985 ( .A1(n1306), .A2(n1155), .A3(n1316), .A4(n1317), .ZN(n1299) );
NOR2_X1 U986 ( .A1(n1338), .A2(n1339), .ZN(n1155) );
INV_X1 U987 ( .A(n1340), .ZN(n1306) );
XNOR2_X1 U988 ( .A(n1341), .B(n1342), .ZN(G21) );
NOR4_X1 U989 ( .A1(KEYINPUT7), .A2(n1343), .A3(n1144), .A4(n1340), .ZN(n1342) );
INV_X1 U990 ( .A(n1133), .ZN(n1144) );
INV_X1 U991 ( .A(n1310), .ZN(n1343) );
NAND2_X1 U992 ( .A1(n1344), .A2(n1345), .ZN(n1310) );
NAND3_X1 U993 ( .A1(n1339), .A2(n1338), .A3(n1346), .ZN(n1345) );
NAND2_X1 U994 ( .A1(KEYINPUT26), .A2(n1161), .ZN(n1344) );
XOR2_X1 U995 ( .A(G116), .B(n1347), .Z(G18) );
NOR3_X1 U996 ( .A1(n1348), .A2(n1349), .A3(n1330), .ZN(n1347) );
NAND3_X1 U997 ( .A1(n1350), .A2(n1351), .A3(n1147), .ZN(n1348) );
NOR2_X1 U998 ( .A1(n1317), .A2(n1352), .ZN(n1147) );
XNOR2_X1 U999 ( .A(KEYINPUT27), .B(n1123), .ZN(n1350) );
INV_X1 U1000 ( .A(n1293), .ZN(n1123) );
XOR2_X1 U1001 ( .A(n1303), .B(n1353), .Z(G15) );
XOR2_X1 U1002 ( .A(KEYINPUT56), .B(G113), .Z(n1353) );
NOR3_X1 U1003 ( .A1(n1340), .A2(n1330), .A3(n1336), .ZN(n1303) );
NAND2_X1 U1004 ( .A1(n1352), .A2(n1317), .ZN(n1336) );
INV_X1 U1005 ( .A(n1316), .ZN(n1352) );
NAND2_X1 U1006 ( .A1(n1354), .A2(n1164), .ZN(n1330) );
XNOR2_X1 U1007 ( .A(n1338), .B(n1346), .ZN(n1354) );
INV_X1 U1008 ( .A(KEYINPUT26), .ZN(n1346) );
NAND3_X1 U1009 ( .A1(n1293), .A2(n1351), .A3(n1132), .ZN(n1340) );
INV_X1 U1010 ( .A(n1349), .ZN(n1132) );
NAND2_X1 U1011 ( .A1(n1151), .A2(n1170), .ZN(n1349) );
XOR2_X1 U1012 ( .A(G110), .B(n1302), .Z(G12) );
AND3_X1 U1013 ( .A1(n1133), .A2(n1305), .A3(n1161), .ZN(n1302) );
NOR2_X1 U1014 ( .A1(n1338), .A2(n1164), .ZN(n1161) );
INV_X1 U1015 ( .A(n1339), .ZN(n1164) );
NAND3_X1 U1016 ( .A1(n1355), .A2(n1356), .A3(n1357), .ZN(n1339) );
NAND2_X1 U1017 ( .A1(G217), .A2(G902), .ZN(n1357) );
NAND3_X1 U1018 ( .A1(n1235), .A2(n1358), .A3(n1359), .ZN(n1356) );
OR2_X1 U1019 ( .A1(n1359), .A2(n1235), .ZN(n1355) );
XNOR2_X1 U1020 ( .A(n1197), .B(n1360), .ZN(n1235) );
XOR2_X1 U1021 ( .A(n1361), .B(n1362), .Z(n1360) );
NOR2_X1 U1022 ( .A1(KEYINPUT58), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1023 ( .A(n1364), .B(n1365), .Z(n1363) );
XNOR2_X1 U1024 ( .A(n1327), .B(G119), .ZN(n1365) );
XOR2_X1 U1025 ( .A(n1366), .B(G110), .Z(n1364) );
NAND3_X1 U1026 ( .A1(n1367), .A2(n1368), .A3(n1369), .ZN(n1366) );
NAND2_X1 U1027 ( .A1(n1370), .A2(n1371), .ZN(n1368) );
INV_X1 U1028 ( .A(KEYINPUT8), .ZN(n1371) );
XNOR2_X1 U1029 ( .A(n1372), .B(n1373), .ZN(n1370) );
NOR2_X1 U1030 ( .A1(G140), .A2(n1374), .ZN(n1373) );
NAND2_X1 U1031 ( .A1(KEYINPUT8), .A2(n1375), .ZN(n1367) );
NOR3_X1 U1032 ( .A1(n1376), .A2(G953), .A3(n1377), .ZN(n1361) );
XNOR2_X1 U1033 ( .A(G234), .B(KEYINPUT20), .ZN(n1377) );
INV_X1 U1034 ( .A(G221), .ZN(n1376) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1378), .ZN(n1359) );
INV_X1 U1036 ( .A(G234), .ZN(n1378) );
NAND2_X1 U1037 ( .A1(n1379), .A2(n1380), .ZN(n1338) );
NAND2_X1 U1038 ( .A1(G472), .A2(n1171), .ZN(n1380) );
XOR2_X1 U1039 ( .A(KEYINPUT15), .B(n1381), .Z(n1379) );
NOR2_X1 U1040 ( .A1(G472), .A2(n1171), .ZN(n1381) );
NAND2_X1 U1041 ( .A1(n1382), .A2(n1358), .ZN(n1171) );
XOR2_X1 U1042 ( .A(n1383), .B(n1384), .Z(n1382) );
XOR2_X1 U1043 ( .A(n1385), .B(n1254), .Z(n1384) );
XOR2_X1 U1044 ( .A(G113), .B(n1386), .Z(n1254) );
NOR2_X1 U1045 ( .A1(KEYINPUT25), .A2(n1387), .ZN(n1386) );
XNOR2_X1 U1046 ( .A(n1388), .B(n1389), .ZN(n1387) );
NOR2_X1 U1047 ( .A1(KEYINPUT36), .A2(n1341), .ZN(n1389) );
XOR2_X1 U1048 ( .A(n1258), .B(n1390), .Z(n1385) );
NOR2_X1 U1049 ( .A1(KEYINPUT17), .A2(n1251), .ZN(n1390) );
XNOR2_X1 U1050 ( .A(n1391), .B(n1392), .ZN(n1251) );
NAND2_X1 U1051 ( .A1(n1393), .A2(G210), .ZN(n1258) );
XNOR2_X1 U1052 ( .A(n1394), .B(n1255), .ZN(n1383) );
XNOR2_X1 U1053 ( .A(KEYINPUT32), .B(KEYINPUT29), .ZN(n1394) );
AND3_X1 U1054 ( .A1(n1142), .A2(n1351), .A3(n1293), .ZN(n1305) );
NOR2_X1 U1055 ( .A1(n1130), .A2(n1131), .ZN(n1293) );
AND2_X1 U1056 ( .A1(G214), .A2(n1395), .ZN(n1131) );
INV_X1 U1057 ( .A(n1320), .ZN(n1130) );
XOR2_X1 U1058 ( .A(n1173), .B(n1180), .Z(n1320) );
NAND2_X1 U1059 ( .A1(G210), .A2(n1395), .ZN(n1180) );
NAND2_X1 U1060 ( .A1(n1358), .A2(n1396), .ZN(n1395) );
INV_X1 U1061 ( .A(G237), .ZN(n1396) );
NAND2_X1 U1062 ( .A1(n1397), .A2(n1358), .ZN(n1173) );
XNOR2_X1 U1063 ( .A(n1398), .B(n1283), .ZN(n1397) );
XNOR2_X1 U1064 ( .A(n1227), .B(n1228), .ZN(n1283) );
INV_X1 U1065 ( .A(n1226), .ZN(n1228) );
XOR2_X1 U1066 ( .A(G110), .B(n1399), .Z(n1226) );
XNOR2_X1 U1067 ( .A(n1400), .B(n1401), .ZN(n1227) );
XNOR2_X1 U1068 ( .A(n1341), .B(G113), .ZN(n1401) );
INV_X1 U1069 ( .A(G119), .ZN(n1341) );
XNOR2_X1 U1070 ( .A(n1402), .B(n1403), .ZN(n1400) );
NAND2_X1 U1071 ( .A1(n1404), .A2(n1405), .ZN(n1402) );
NAND2_X1 U1072 ( .A1(G101), .A2(n1406), .ZN(n1405) );
XOR2_X1 U1073 ( .A(KEYINPUT44), .B(n1407), .Z(n1404) );
NOR2_X1 U1074 ( .A1(G101), .A2(n1406), .ZN(n1407) );
XNOR2_X1 U1075 ( .A(n1114), .B(G104), .ZN(n1406) );
NAND2_X1 U1076 ( .A1(n1408), .A2(KEYINPUT47), .ZN(n1398) );
XNOR2_X1 U1077 ( .A(n1280), .B(n1409), .ZN(n1408) );
INV_X1 U1078 ( .A(n1278), .ZN(n1409) );
XOR2_X1 U1079 ( .A(G125), .B(n1392), .Z(n1278) );
AND2_X1 U1080 ( .A1(n1410), .A2(n1411), .ZN(n1392) );
NAND2_X1 U1081 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
NAND2_X1 U1082 ( .A1(n1414), .A2(n1415), .ZN(n1413) );
XNOR2_X1 U1083 ( .A(KEYINPUT16), .B(n1327), .ZN(n1412) );
XOR2_X1 U1084 ( .A(KEYINPUT41), .B(n1416), .Z(n1410) );
AND3_X1 U1085 ( .A1(n1414), .A2(n1327), .A3(n1415), .ZN(n1416) );
NAND2_X1 U1086 ( .A1(n1417), .A2(n1372), .ZN(n1415) );
XNOR2_X1 U1087 ( .A(KEYINPUT52), .B(n1313), .ZN(n1417) );
NAND2_X1 U1088 ( .A1(G224), .A2(n1129), .ZN(n1280) );
NAND2_X1 U1089 ( .A1(n1153), .A2(n1418), .ZN(n1351) );
NAND3_X1 U1090 ( .A1(n1224), .A2(n1335), .A3(G902), .ZN(n1418) );
NOR2_X1 U1091 ( .A1(n1129), .A2(G898), .ZN(n1224) );
NAND3_X1 U1092 ( .A1(n1335), .A2(n1129), .A3(n1419), .ZN(n1153) );
XNOR2_X1 U1093 ( .A(G952), .B(KEYINPUT57), .ZN(n1419) );
NAND2_X1 U1094 ( .A1(G237), .A2(G234), .ZN(n1335) );
NOR2_X1 U1095 ( .A1(n1151), .A2(n1152), .ZN(n1142) );
INV_X1 U1096 ( .A(n1170), .ZN(n1152) );
NAND2_X1 U1097 ( .A1(G221), .A2(n1420), .ZN(n1170) );
NAND2_X1 U1098 ( .A1(G234), .A2(n1358), .ZN(n1420) );
XOR2_X1 U1099 ( .A(n1421), .B(G469), .Z(n1151) );
NAND2_X1 U1100 ( .A1(n1422), .A2(n1358), .ZN(n1421) );
XOR2_X1 U1101 ( .A(n1423), .B(n1424), .Z(n1422) );
XOR2_X1 U1102 ( .A(n1273), .B(n1425), .Z(n1424) );
XOR2_X1 U1103 ( .A(KEYINPUT9), .B(KEYINPUT43), .Z(n1425) );
NOR2_X1 U1104 ( .A1(n1187), .A2(G953), .ZN(n1273) );
INV_X1 U1105 ( .A(G227), .ZN(n1187) );
XOR2_X1 U1106 ( .A(n1426), .B(n1427), .Z(n1423) );
NOR2_X1 U1107 ( .A1(n1428), .A2(n1429), .ZN(n1427) );
NOR3_X1 U1108 ( .A1(KEYINPUT49), .A2(G110), .A3(n1430), .ZN(n1429) );
NOR2_X1 U1109 ( .A1(n1264), .A2(n1431), .ZN(n1428) );
INV_X1 U1110 ( .A(KEYINPUT49), .ZN(n1431) );
XNOR2_X1 U1111 ( .A(G110), .B(n1430), .ZN(n1264) );
XNOR2_X1 U1112 ( .A(n1268), .B(n1270), .ZN(n1426) );
XNOR2_X1 U1113 ( .A(n1432), .B(n1433), .ZN(n1270) );
XNOR2_X1 U1114 ( .A(G104), .B(n1255), .ZN(n1433) );
INV_X1 U1115 ( .A(G101), .ZN(n1255) );
NAND2_X1 U1116 ( .A1(KEYINPUT33), .A2(n1114), .ZN(n1432) );
INV_X1 U1117 ( .A(G107), .ZN(n1114) );
XNOR2_X1 U1118 ( .A(n1202), .B(n1391), .ZN(n1268) );
XOR2_X1 U1119 ( .A(n1199), .B(n1197), .Z(n1391) );
XOR2_X1 U1120 ( .A(G137), .B(KEYINPUT59), .Z(n1197) );
XOR2_X1 U1121 ( .A(G131), .B(G134), .Z(n1199) );
NAND3_X1 U1122 ( .A1(n1434), .A2(n1435), .A3(n1436), .ZN(n1202) );
OR2_X1 U1123 ( .A1(n1414), .A2(G128), .ZN(n1436) );
NAND2_X1 U1124 ( .A1(G146), .A2(n1313), .ZN(n1414) );
NAND3_X1 U1125 ( .A1(G128), .A2(G143), .A3(G146), .ZN(n1435) );
NAND2_X1 U1126 ( .A1(n1437), .A2(n1372), .ZN(n1434) );
XNOR2_X1 U1127 ( .A(n1313), .B(G128), .ZN(n1437) );
NOR2_X1 U1128 ( .A1(n1316), .A2(n1317), .ZN(n1133) );
XNOR2_X1 U1129 ( .A(n1438), .B(G475), .ZN(n1317) );
NAND2_X1 U1130 ( .A1(n1243), .A2(n1358), .ZN(n1438) );
XOR2_X1 U1131 ( .A(n1439), .B(n1440), .Z(n1243) );
XOR2_X1 U1132 ( .A(G104), .B(n1441), .Z(n1440) );
XNOR2_X1 U1133 ( .A(n1313), .B(G131), .ZN(n1441) );
XOR2_X1 U1134 ( .A(n1442), .B(n1443), .Z(n1439) );
AND2_X1 U1135 ( .A1(G214), .A2(n1393), .ZN(n1443) );
NOR2_X1 U1136 ( .A1(G953), .A2(G237), .ZN(n1393) );
XOR2_X1 U1137 ( .A(n1444), .B(n1445), .Z(n1442) );
NOR2_X1 U1138 ( .A1(n1446), .A2(n1447), .ZN(n1445) );
XOR2_X1 U1139 ( .A(KEYINPUT12), .B(n1448), .Z(n1447) );
NOR2_X1 U1140 ( .A1(G113), .A2(n1399), .ZN(n1448) );
AND2_X1 U1141 ( .A1(n1399), .A2(G113), .ZN(n1446) );
INV_X1 U1142 ( .A(G122), .ZN(n1399) );
NAND2_X1 U1143 ( .A1(n1449), .A2(n1369), .ZN(n1444) );
NAND3_X1 U1144 ( .A1(G146), .A2(n1374), .A3(G140), .ZN(n1369) );
INV_X1 U1145 ( .A(G125), .ZN(n1374) );
INV_X1 U1146 ( .A(n1375), .ZN(n1449) );
NAND2_X1 U1147 ( .A1(n1450), .A2(n1451), .ZN(n1375) );
NAND2_X1 U1148 ( .A1(n1452), .A2(n1372), .ZN(n1451) );
INV_X1 U1149 ( .A(G146), .ZN(n1372) );
XNOR2_X1 U1150 ( .A(G125), .B(G140), .ZN(n1452) );
NAND3_X1 U1151 ( .A1(G125), .A2(n1430), .A3(G146), .ZN(n1450) );
INV_X1 U1152 ( .A(G140), .ZN(n1430) );
XNOR2_X1 U1153 ( .A(n1453), .B(G478), .ZN(n1316) );
NAND2_X1 U1154 ( .A1(n1240), .A2(n1358), .ZN(n1453) );
INV_X1 U1155 ( .A(G902), .ZN(n1358) );
XOR2_X1 U1156 ( .A(n1454), .B(n1455), .Z(n1240) );
XOR2_X1 U1157 ( .A(n1456), .B(n1457), .Z(n1455) );
XNOR2_X1 U1158 ( .A(G134), .B(n1327), .ZN(n1457) );
INV_X1 U1159 ( .A(G128), .ZN(n1327) );
XNOR2_X1 U1160 ( .A(KEYINPUT23), .B(n1313), .ZN(n1456) );
INV_X1 U1161 ( .A(G143), .ZN(n1313) );
XOR2_X1 U1162 ( .A(n1458), .B(n1459), .Z(n1454) );
XNOR2_X1 U1163 ( .A(n1460), .B(n1403), .ZN(n1459) );
INV_X1 U1164 ( .A(n1388), .ZN(n1403) );
XOR2_X1 U1165 ( .A(G116), .B(KEYINPUT14), .Z(n1388) );
AND3_X1 U1166 ( .A1(G217), .A2(n1129), .A3(G234), .ZN(n1460) );
INV_X1 U1167 ( .A(G953), .ZN(n1129) );
XNOR2_X1 U1168 ( .A(G122), .B(G107), .ZN(n1458) );
endmodule


