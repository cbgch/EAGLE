//Key = 0000110011100101010000010000001100000010110000011101101110101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;

XOR2_X1 U781 ( .A(G107), .B(n1072), .Z(G9) );
NOR2_X1 U782 ( .A1(n1073), .A2(n1074), .ZN(G75) );
NOR4_X1 U783 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
INV_X1 U784 ( .A(n1079), .ZN(n1077) );
NOR2_X1 U785 ( .A1(n1080), .A2(n1081), .ZN(n1076) );
NOR2_X1 U786 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR4_X1 U787 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1083) );
NOR2_X1 U788 ( .A1(n1088), .A2(n1089), .ZN(n1085) );
NOR2_X1 U789 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NOR3_X1 U790 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
XNOR2_X1 U791 ( .A(KEYINPUT61), .B(n1095), .ZN(n1094) );
NOR2_X1 U792 ( .A1(n1096), .A2(n1097), .ZN(n1090) );
NOR2_X1 U793 ( .A1(n1098), .A2(n1099), .ZN(n1084) );
NOR2_X1 U794 ( .A1(n1092), .A2(n1100), .ZN(n1099) );
NOR4_X1 U795 ( .A1(n1092), .A2(n1101), .A3(n1100), .A4(n1088), .ZN(n1082) );
NOR3_X1 U796 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NOR2_X1 U797 ( .A1(n1105), .A2(n1086), .ZN(n1104) );
INV_X1 U798 ( .A(n1106), .ZN(n1086) );
NOR3_X1 U799 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1105) );
NOR3_X1 U800 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
INV_X1 U801 ( .A(KEYINPUT15), .ZN(n1110) );
NOR2_X1 U802 ( .A1(KEYINPUT15), .A2(n1087), .ZN(n1108) );
NOR2_X1 U803 ( .A1(n1113), .A2(n1114), .ZN(n1103) );
XNOR2_X1 U804 ( .A(KEYINPUT47), .B(n1087), .ZN(n1114) );
AND2_X1 U805 ( .A1(n1115), .A2(n1116), .ZN(n1102) );
NOR3_X1 U806 ( .A1(n1078), .A2(G952), .A3(n1075), .ZN(n1073) );
AND4_X1 U807 ( .A1(n1117), .A2(n1097), .A3(n1118), .A4(n1119), .ZN(n1075) );
NOR4_X1 U808 ( .A1(n1120), .A2(n1121), .A3(n1087), .A4(n1122), .ZN(n1119) );
AND2_X1 U809 ( .A1(n1123), .A2(G469), .ZN(n1121) );
NOR3_X1 U810 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1120) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
AND3_X1 U812 ( .A1(n1128), .A2(n1127), .A3(KEYINPUT23), .ZN(n1125) );
NOR2_X1 U813 ( .A1(n1129), .A2(KEYINPUT46), .ZN(n1127) );
NOR2_X1 U814 ( .A1(KEYINPUT23), .A2(n1130), .ZN(n1124) );
NOR3_X1 U815 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1118) );
INV_X1 U816 ( .A(n1134), .ZN(n1131) );
NAND2_X1 U817 ( .A1(n1135), .A2(n1136), .ZN(n1117) );
NAND2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U819 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U820 ( .A1(KEYINPUT48), .A2(G472), .ZN(n1140) );
NAND2_X1 U821 ( .A1(n1141), .A2(n1142), .ZN(n1135) );
NAND2_X1 U822 ( .A1(KEYINPUT48), .A2(n1143), .ZN(n1141) );
NAND2_X1 U823 ( .A1(n1144), .A2(n1139), .ZN(n1143) );
INV_X1 U824 ( .A(KEYINPUT36), .ZN(n1139) );
XOR2_X1 U825 ( .A(n1145), .B(n1146), .Z(G72) );
NOR3_X1 U826 ( .A1(n1147), .A2(KEYINPUT50), .A3(n1148), .ZN(n1146) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
INV_X1 U828 ( .A(G900), .ZN(n1150) );
XNOR2_X1 U829 ( .A(G227), .B(KEYINPUT24), .ZN(n1149) );
NAND2_X1 U830 ( .A1(n1151), .A2(n1152), .ZN(n1145) );
NAND2_X1 U831 ( .A1(n1153), .A2(n1147), .ZN(n1152) );
XOR2_X1 U832 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND3_X1 U833 ( .A1(n1155), .A2(n1156), .A3(G953), .ZN(n1151) );
NOR2_X1 U834 ( .A1(KEYINPUT3), .A2(n1157), .ZN(n1155) );
NOR3_X1 U835 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1157) );
NOR2_X1 U836 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
AND3_X1 U837 ( .A1(n1162), .A2(n1161), .A3(KEYINPUT51), .ZN(n1159) );
AND2_X1 U838 ( .A1(KEYINPUT9), .A2(n1163), .ZN(n1161) );
NAND2_X1 U839 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NAND2_X1 U840 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U841 ( .A(KEYINPUT41), .B(n1168), .Z(n1164) );
NOR2_X1 U842 ( .A1(n1166), .A2(n1167), .ZN(n1168) );
XOR2_X1 U843 ( .A(G131), .B(n1169), .Z(n1167) );
NOR2_X1 U844 ( .A1(KEYINPUT51), .A2(n1163), .ZN(n1158) );
XNOR2_X1 U845 ( .A(G140), .B(G125), .ZN(n1163) );
XOR2_X1 U846 ( .A(n1170), .B(n1171), .Z(G69) );
NOR2_X1 U847 ( .A1(KEYINPUT11), .A2(n1172), .ZN(n1171) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U849 ( .A1(n1147), .A2(n1175), .ZN(n1174) );
NAND2_X1 U850 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
NAND2_X1 U851 ( .A1(G953), .A2(n1178), .ZN(n1177) );
XOR2_X1 U852 ( .A(n1179), .B(n1180), .Z(n1176) );
NOR2_X1 U853 ( .A1(KEYINPUT7), .A2(n1181), .ZN(n1179) );
XOR2_X1 U854 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U855 ( .A(n1184), .B(KEYINPUT31), .ZN(n1182) );
NAND2_X1 U856 ( .A1(n1185), .A2(G953), .ZN(n1170) );
XOR2_X1 U857 ( .A(n1186), .B(KEYINPUT18), .Z(n1185) );
NAND2_X1 U858 ( .A1(G898), .A2(G224), .ZN(n1186) );
NOR2_X1 U859 ( .A1(n1187), .A2(n1188), .ZN(G66) );
NOR3_X1 U860 ( .A1(n1129), .A2(n1189), .A3(n1190), .ZN(n1188) );
NOR3_X1 U861 ( .A1(n1191), .A2(n1128), .A3(n1192), .ZN(n1190) );
INV_X1 U862 ( .A(n1193), .ZN(n1191) );
NOR2_X1 U863 ( .A1(n1194), .A2(n1193), .ZN(n1189) );
NOR2_X1 U864 ( .A1(n1079), .A2(n1128), .ZN(n1194) );
NOR2_X1 U865 ( .A1(n1187), .A2(n1195), .ZN(G63) );
XOR2_X1 U866 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U867 ( .A1(n1198), .A2(n1192), .ZN(n1197) );
NAND2_X1 U868 ( .A1(KEYINPUT58), .A2(n1199), .ZN(n1196) );
NOR2_X1 U869 ( .A1(n1187), .A2(n1200), .ZN(G60) );
XOR2_X1 U870 ( .A(n1201), .B(n1202), .Z(n1200) );
AND2_X1 U871 ( .A1(G475), .A2(n1203), .ZN(n1201) );
XOR2_X1 U872 ( .A(G104), .B(n1204), .Z(G6) );
NOR2_X1 U873 ( .A1(n1187), .A2(n1205), .ZN(G57) );
XOR2_X1 U874 ( .A(n1206), .B(n1207), .Z(n1205) );
XNOR2_X1 U875 ( .A(n1208), .B(n1209), .ZN(n1207) );
XNOR2_X1 U876 ( .A(n1210), .B(n1211), .ZN(n1209) );
XOR2_X1 U877 ( .A(n1212), .B(n1213), .Z(n1206) );
XOR2_X1 U878 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U879 ( .A1(n1142), .A2(n1192), .ZN(n1215) );
INV_X1 U880 ( .A(n1203), .ZN(n1192) );
INV_X1 U881 ( .A(G472), .ZN(n1142) );
NAND2_X1 U882 ( .A1(KEYINPUT55), .A2(n1216), .ZN(n1212) );
NOR2_X1 U883 ( .A1(n1187), .A2(n1217), .ZN(G54) );
XOR2_X1 U884 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U885 ( .A(n1220), .B(n1221), .Z(n1219) );
NOR2_X1 U886 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
XOR2_X1 U887 ( .A(KEYINPUT44), .B(KEYINPUT16), .Z(n1223) );
NOR2_X1 U888 ( .A1(KEYINPUT35), .A2(n1224), .ZN(n1220) );
XOR2_X1 U889 ( .A(n1225), .B(n1226), .Z(n1218) );
NOR2_X1 U890 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NOR2_X1 U891 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NOR2_X1 U892 ( .A1(n1231), .A2(n1232), .ZN(n1229) );
INV_X1 U893 ( .A(KEYINPUT5), .ZN(n1232) );
NOR2_X1 U894 ( .A1(KEYINPUT57), .A2(n1166), .ZN(n1231) );
INV_X1 U895 ( .A(n1233), .ZN(n1166) );
NOR2_X1 U896 ( .A1(n1234), .A2(n1233), .ZN(n1227) );
XOR2_X1 U897 ( .A(G128), .B(n1235), .Z(n1233) );
NOR2_X1 U898 ( .A1(n1236), .A2(KEYINPUT57), .ZN(n1234) );
AND2_X1 U899 ( .A1(n1230), .A2(KEYINPUT5), .ZN(n1236) );
XNOR2_X1 U900 ( .A(G101), .B(n1237), .ZN(n1230) );
NAND2_X1 U901 ( .A1(n1203), .A2(G469), .ZN(n1225) );
NOR2_X1 U902 ( .A1(n1187), .A2(n1238), .ZN(G51) );
XOR2_X1 U903 ( .A(n1239), .B(n1240), .Z(n1238) );
XNOR2_X1 U904 ( .A(n1241), .B(n1242), .ZN(n1240) );
NAND2_X1 U905 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
NAND2_X1 U906 ( .A1(G125), .A2(n1245), .ZN(n1244) );
XOR2_X1 U907 ( .A(KEYINPUT38), .B(n1246), .Z(n1243) );
NOR2_X1 U908 ( .A1(G125), .A2(n1245), .ZN(n1246) );
XOR2_X1 U909 ( .A(n1247), .B(n1248), .Z(n1239) );
NAND2_X1 U910 ( .A1(n1203), .A2(n1249), .ZN(n1247) );
NOR2_X1 U911 ( .A1(n1250), .A2(n1079), .ZN(n1203) );
NOR2_X1 U912 ( .A1(n1175), .A2(n1154), .ZN(n1079) );
NAND4_X1 U913 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1154) );
NOR4_X1 U914 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1254) );
NOR4_X1 U915 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1258) );
INV_X1 U916 ( .A(n1263), .ZN(n1257) );
NOR2_X1 U917 ( .A1(n1264), .A2(n1265), .ZN(n1253) );
NOR2_X1 U918 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND4_X1 U919 ( .A1(n1268), .A2(n1093), .A3(n1269), .A4(n1113), .ZN(n1267) );
INV_X1 U920 ( .A(KEYINPUT45), .ZN(n1266) );
NOR2_X1 U921 ( .A1(KEYINPUT45), .A2(n1270), .ZN(n1264) );
NAND2_X1 U922 ( .A1(n1271), .A2(n1115), .ZN(n1252) );
XOR2_X1 U923 ( .A(n1272), .B(KEYINPUT8), .Z(n1271) );
NAND2_X1 U924 ( .A1(n1273), .A2(n1274), .ZN(n1251) );
NAND2_X1 U925 ( .A1(n1275), .A2(n1095), .ZN(n1274) );
XNOR2_X1 U926 ( .A(n1093), .B(KEYINPUT63), .ZN(n1275) );
NAND2_X1 U927 ( .A1(n1276), .A2(n1277), .ZN(n1175) );
NOR4_X1 U928 ( .A1(n1278), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1277) );
NOR4_X1 U929 ( .A1(n1282), .A2(n1283), .A3(n1204), .A4(n1072), .ZN(n1276) );
AND3_X1 U930 ( .A1(n1284), .A2(n1106), .A3(n1285), .ZN(n1072) );
AND3_X1 U931 ( .A1(n1285), .A2(n1106), .A3(n1093), .ZN(n1204) );
NOR2_X1 U932 ( .A1(n1147), .A2(G952), .ZN(n1187) );
XOR2_X1 U933 ( .A(G146), .B(n1286), .Z(G48) );
NOR2_X1 U934 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U935 ( .A(G143), .B(n1289), .ZN(G45) );
NAND4_X1 U936 ( .A1(n1290), .A2(n1291), .A3(n1122), .A4(n1292), .ZN(n1289) );
XNOR2_X1 U937 ( .A(KEYINPUT53), .B(n1261), .ZN(n1291) );
XNOR2_X1 U938 ( .A(n1293), .B(n1256), .ZN(G42) );
NOR4_X1 U939 ( .A1(n1294), .A2(n1287), .A3(n1113), .A4(n1087), .ZN(n1256) );
INV_X1 U940 ( .A(n1093), .ZN(n1287) );
NAND2_X1 U941 ( .A1(n1295), .A2(n1296), .ZN(G39) );
OR2_X1 U942 ( .A1(n1263), .A2(G137), .ZN(n1296) );
XOR2_X1 U943 ( .A(n1297), .B(KEYINPUT62), .Z(n1295) );
NAND2_X1 U944 ( .A1(G137), .A2(n1263), .ZN(n1297) );
NAND4_X1 U945 ( .A1(n1298), .A2(n1299), .A3(n1115), .A4(n1300), .ZN(n1263) );
NOR2_X1 U946 ( .A1(n1100), .A2(n1294), .ZN(n1300) );
INV_X1 U947 ( .A(n1096), .ZN(n1100) );
INV_X1 U948 ( .A(n1087), .ZN(n1115) );
XOR2_X1 U949 ( .A(G134), .B(n1255), .Z(G36) );
NOR3_X1 U950 ( .A1(n1087), .A2(n1095), .A3(n1262), .ZN(n1255) );
INV_X1 U951 ( .A(n1284), .ZN(n1095) );
XOR2_X1 U952 ( .A(G131), .B(n1301), .Z(G33) );
NOR2_X1 U953 ( .A1(n1087), .A2(n1272), .ZN(n1301) );
NAND2_X1 U954 ( .A1(n1290), .A2(n1093), .ZN(n1272) );
INV_X1 U955 ( .A(n1262), .ZN(n1290) );
NAND2_X1 U956 ( .A1(n1302), .A2(n1116), .ZN(n1262) );
NAND2_X1 U957 ( .A1(n1303), .A2(n1112), .ZN(n1087) );
INV_X1 U958 ( .A(n1111), .ZN(n1303) );
XNOR2_X1 U959 ( .A(G128), .B(n1304), .ZN(G30) );
NAND3_X1 U960 ( .A1(n1273), .A2(n1284), .A3(KEYINPUT17), .ZN(n1304) );
INV_X1 U961 ( .A(n1288), .ZN(n1273) );
NAND4_X1 U962 ( .A1(n1302), .A2(n1107), .A3(n1298), .A4(n1299), .ZN(n1288) );
INV_X1 U963 ( .A(n1261), .ZN(n1107) );
INV_X1 U964 ( .A(n1294), .ZN(n1302) );
NAND3_X1 U965 ( .A1(n1097), .A2(n1088), .A3(n1269), .ZN(n1294) );
XNOR2_X1 U966 ( .A(n1216), .B(n1283), .ZN(G3) );
AND3_X1 U967 ( .A1(n1096), .A2(n1285), .A3(n1116), .ZN(n1283) );
XNOR2_X1 U968 ( .A(G125), .B(n1270), .ZN(G27) );
NAND4_X1 U969 ( .A1(n1268), .A2(n1093), .A3(n1305), .A4(n1269), .ZN(n1270) );
NAND2_X1 U970 ( .A1(n1081), .A2(n1306), .ZN(n1269) );
NAND4_X1 U971 ( .A1(n1307), .A2(G953), .A3(G902), .A4(n1308), .ZN(n1306) );
INV_X1 U972 ( .A(n1156), .ZN(n1307) );
XOR2_X1 U973 ( .A(G900), .B(KEYINPUT28), .Z(n1156) );
XOR2_X1 U974 ( .A(G122), .B(n1282), .Z(G24) );
AND4_X1 U975 ( .A1(n1309), .A2(n1106), .A3(n1122), .A4(n1292), .ZN(n1282) );
NOR2_X1 U976 ( .A1(n1299), .A2(n1298), .ZN(n1106) );
XOR2_X1 U977 ( .A(G119), .B(n1281), .Z(G21) );
AND4_X1 U978 ( .A1(n1309), .A2(n1096), .A3(n1298), .A4(n1299), .ZN(n1281) );
NAND2_X1 U979 ( .A1(n1310), .A2(n1311), .ZN(G18) );
NAND2_X1 U980 ( .A1(n1280), .A2(n1312), .ZN(n1311) );
XOR2_X1 U981 ( .A(KEYINPUT52), .B(n1313), .Z(n1310) );
NOR2_X1 U982 ( .A1(n1280), .A2(n1312), .ZN(n1313) );
AND3_X1 U983 ( .A1(n1116), .A2(n1284), .A3(n1309), .ZN(n1280) );
AND2_X1 U984 ( .A1(n1268), .A2(n1314), .ZN(n1309) );
NOR3_X1 U985 ( .A1(n1261), .A2(n1092), .A3(n1088), .ZN(n1268) );
INV_X1 U986 ( .A(n1098), .ZN(n1088) );
NOR2_X1 U987 ( .A1(n1122), .A2(n1259), .ZN(n1284) );
INV_X1 U988 ( .A(n1292), .ZN(n1259) );
XNOR2_X1 U989 ( .A(n1279), .B(n1315), .ZN(G15) );
XNOR2_X1 U990 ( .A(G113), .B(KEYINPUT25), .ZN(n1315) );
AND4_X1 U991 ( .A1(n1116), .A2(n1093), .A3(n1098), .A4(n1316), .ZN(n1279) );
NOR3_X1 U992 ( .A1(n1317), .A2(n1092), .A3(n1318), .ZN(n1316) );
NOR2_X1 U993 ( .A1(n1292), .A2(n1260), .ZN(n1093) );
INV_X1 U994 ( .A(n1122), .ZN(n1260) );
NOR2_X1 U995 ( .A1(n1298), .A2(n1319), .ZN(n1116) );
XOR2_X1 U996 ( .A(G110), .B(n1278), .Z(G12) );
AND3_X1 U997 ( .A1(n1305), .A2(n1285), .A3(n1096), .ZN(n1278) );
NOR2_X1 U998 ( .A1(n1292), .A2(n1122), .ZN(n1096) );
XNOR2_X1 U999 ( .A(n1320), .B(G475), .ZN(n1122) );
OR2_X1 U1000 ( .A1(n1202), .A2(G902), .ZN(n1320) );
XNOR2_X1 U1001 ( .A(n1321), .B(n1322), .ZN(n1202) );
XOR2_X1 U1002 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1003 ( .A(n1325), .B(G113), .Z(n1324) );
NAND2_X1 U1004 ( .A1(n1326), .A2(G214), .ZN(n1325) );
XNOR2_X1 U1005 ( .A(G146), .B(G140), .ZN(n1323) );
XNOR2_X1 U1006 ( .A(n1327), .B(n1328), .ZN(n1321) );
INV_X1 U1007 ( .A(n1329), .ZN(n1328) );
XOR2_X1 U1008 ( .A(n1330), .B(n1331), .Z(n1327) );
NAND2_X1 U1009 ( .A1(KEYINPUT49), .A2(n1332), .ZN(n1330) );
NAND2_X1 U1010 ( .A1(n1333), .A2(n1134), .ZN(n1292) );
NAND2_X1 U1011 ( .A1(G478), .A2(n1334), .ZN(n1134) );
NAND2_X1 U1012 ( .A1(n1250), .A2(n1199), .ZN(n1334) );
XNOR2_X1 U1013 ( .A(n1132), .B(KEYINPUT37), .ZN(n1333) );
AND3_X1 U1014 ( .A1(n1198), .A2(n1250), .A3(n1199), .ZN(n1132) );
NAND2_X1 U1015 ( .A1(n1335), .A2(n1336), .ZN(n1199) );
NAND3_X1 U1016 ( .A1(n1337), .A2(n1338), .A3(G217), .ZN(n1336) );
NAND2_X1 U1017 ( .A1(n1339), .A2(n1340), .ZN(n1335) );
NAND2_X1 U1018 ( .A1(G217), .A2(n1338), .ZN(n1340) );
INV_X1 U1019 ( .A(n1341), .ZN(n1338) );
XOR2_X1 U1020 ( .A(n1337), .B(KEYINPUT40), .Z(n1339) );
XOR2_X1 U1021 ( .A(n1342), .B(n1343), .Z(n1337) );
XOR2_X1 U1022 ( .A(n1331), .B(n1344), .Z(n1343) );
XOR2_X1 U1023 ( .A(G122), .B(G143), .Z(n1331) );
XNOR2_X1 U1024 ( .A(G134), .B(G116), .ZN(n1342) );
INV_X1 U1025 ( .A(G478), .ZN(n1198) );
NOR4_X1 U1026 ( .A1(n1317), .A2(n1318), .A3(n1092), .A4(n1098), .ZN(n1285) );
NOR2_X1 U1027 ( .A1(n1345), .A2(n1133), .ZN(n1098) );
NOR2_X1 U1028 ( .A1(n1123), .A2(G469), .ZN(n1133) );
AND2_X1 U1029 ( .A1(n1346), .A2(n1123), .ZN(n1345) );
NAND2_X1 U1030 ( .A1(n1347), .A2(n1250), .ZN(n1123) );
XOR2_X1 U1031 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1032 ( .A(n1350), .B(n1235), .Z(n1349) );
XNOR2_X1 U1033 ( .A(n1351), .B(n1352), .ZN(n1235) );
NOR2_X1 U1034 ( .A1(G146), .A2(KEYINPUT14), .ZN(n1352) );
XNOR2_X1 U1035 ( .A(G143), .B(KEYINPUT1), .ZN(n1351) );
XNOR2_X1 U1036 ( .A(n1329), .B(n1344), .ZN(n1350) );
XOR2_X1 U1037 ( .A(G107), .B(G128), .Z(n1344) );
XOR2_X1 U1038 ( .A(G104), .B(G131), .Z(n1329) );
XOR2_X1 U1039 ( .A(n1353), .B(n1354), .Z(n1348) );
NOR2_X1 U1040 ( .A1(KEYINPUT59), .A2(n1222), .ZN(n1354) );
XNOR2_X1 U1041 ( .A(n1355), .B(n1356), .ZN(n1222) );
XNOR2_X1 U1042 ( .A(n1293), .B(G110), .ZN(n1356) );
NAND2_X1 U1043 ( .A1(G227), .A2(n1147), .ZN(n1355) );
XNOR2_X1 U1044 ( .A(n1357), .B(n1216), .ZN(n1353) );
XNOR2_X1 U1045 ( .A(G469), .B(KEYINPUT30), .ZN(n1346) );
INV_X1 U1046 ( .A(n1097), .ZN(n1092) );
NAND2_X1 U1047 ( .A1(n1358), .A2(G221), .ZN(n1097) );
XOR2_X1 U1048 ( .A(n1359), .B(KEYINPUT19), .Z(n1358) );
INV_X1 U1049 ( .A(n1314), .ZN(n1318) );
NAND2_X1 U1050 ( .A1(n1081), .A2(n1360), .ZN(n1314) );
NAND4_X1 U1051 ( .A1(G953), .A2(G902), .A3(n1308), .A4(n1178), .ZN(n1360) );
INV_X1 U1052 ( .A(G898), .ZN(n1178) );
NAND3_X1 U1053 ( .A1(n1361), .A2(n1308), .A3(G952), .ZN(n1081) );
NAND2_X1 U1054 ( .A1(G237), .A2(n1362), .ZN(n1308) );
XOR2_X1 U1055 ( .A(KEYINPUT0), .B(G234), .Z(n1362) );
INV_X1 U1056 ( .A(n1078), .ZN(n1361) );
XOR2_X1 U1057 ( .A(G953), .B(KEYINPUT42), .Z(n1078) );
XOR2_X1 U1058 ( .A(n1261), .B(KEYINPUT22), .Z(n1317) );
NAND2_X1 U1059 ( .A1(n1111), .A2(n1112), .ZN(n1261) );
NAND2_X1 U1060 ( .A1(G214), .A2(n1363), .ZN(n1112) );
XNOR2_X1 U1061 ( .A(n1364), .B(n1249), .ZN(n1111) );
AND2_X1 U1062 ( .A1(G210), .A2(n1363), .ZN(n1249) );
NAND2_X1 U1063 ( .A1(n1365), .A2(n1250), .ZN(n1363) );
XNOR2_X1 U1064 ( .A(G237), .B(KEYINPUT27), .ZN(n1365) );
NAND2_X1 U1065 ( .A1(n1366), .A2(n1250), .ZN(n1364) );
XOR2_X1 U1066 ( .A(n1367), .B(n1368), .Z(n1366) );
XNOR2_X1 U1067 ( .A(n1369), .B(n1208), .ZN(n1368) );
NOR2_X1 U1068 ( .A1(KEYINPUT20), .A2(n1242), .ZN(n1369) );
XOR2_X1 U1069 ( .A(n1370), .B(n1180), .Z(n1242) );
XOR2_X1 U1070 ( .A(G122), .B(G110), .Z(n1180) );
XNOR2_X1 U1071 ( .A(KEYINPUT6), .B(n1371), .ZN(n1370) );
NOR2_X1 U1072 ( .A1(KEYINPUT21), .A2(n1372), .ZN(n1371) );
XNOR2_X1 U1073 ( .A(n1373), .B(n1183), .ZN(n1372) );
XOR2_X1 U1074 ( .A(n1374), .B(n1216), .Z(n1183) );
NAND2_X1 U1075 ( .A1(KEYINPUT54), .A2(n1237), .ZN(n1374) );
XOR2_X1 U1076 ( .A(G104), .B(G107), .Z(n1237) );
NAND2_X1 U1077 ( .A1(KEYINPUT13), .A2(n1210), .ZN(n1373) );
XNOR2_X1 U1078 ( .A(G125), .B(n1248), .ZN(n1367) );
AND2_X1 U1079 ( .A1(G224), .A2(n1147), .ZN(n1248) );
INV_X1 U1080 ( .A(n1113), .ZN(n1305) );
NAND2_X1 U1081 ( .A1(n1319), .A2(n1298), .ZN(n1113) );
NAND3_X1 U1082 ( .A1(n1375), .A2(n1376), .A3(n1377), .ZN(n1298) );
NAND2_X1 U1083 ( .A1(n1129), .A2(n1128), .ZN(n1377) );
NAND2_X1 U1084 ( .A1(KEYINPUT2), .A2(n1378), .ZN(n1376) );
NAND2_X1 U1085 ( .A1(n1379), .A2(n1130), .ZN(n1378) );
INV_X1 U1086 ( .A(n1129), .ZN(n1130) );
XNOR2_X1 U1087 ( .A(KEYINPUT34), .B(n1128), .ZN(n1379) );
NAND2_X1 U1088 ( .A1(n1380), .A2(n1381), .ZN(n1375) );
INV_X1 U1089 ( .A(KEYINPUT2), .ZN(n1381) );
NAND2_X1 U1090 ( .A1(n1382), .A2(n1383), .ZN(n1380) );
NAND2_X1 U1091 ( .A1(KEYINPUT34), .A2(n1128), .ZN(n1383) );
OR3_X1 U1092 ( .A1(n1129), .A2(KEYINPUT34), .A3(n1128), .ZN(n1382) );
NAND2_X1 U1093 ( .A1(G217), .A2(n1359), .ZN(n1128) );
NAND2_X1 U1094 ( .A1(G234), .A2(n1250), .ZN(n1359) );
NOR2_X1 U1095 ( .A1(n1193), .A2(G902), .ZN(n1129) );
XNOR2_X1 U1096 ( .A(n1384), .B(n1385), .ZN(n1193) );
XOR2_X1 U1097 ( .A(n1386), .B(n1387), .Z(n1385) );
XNOR2_X1 U1098 ( .A(n1388), .B(G119), .ZN(n1387) );
INV_X1 U1099 ( .A(G128), .ZN(n1388) );
XOR2_X1 U1100 ( .A(G146), .B(G137), .Z(n1386) );
XOR2_X1 U1101 ( .A(n1389), .B(n1390), .Z(n1384) );
XOR2_X1 U1102 ( .A(G110), .B(n1391), .Z(n1390) );
NOR3_X1 U1103 ( .A1(n1341), .A2(KEYINPUT26), .A3(n1392), .ZN(n1391) );
INV_X1 U1104 ( .A(G221), .ZN(n1392) );
NAND2_X1 U1105 ( .A1(G234), .A2(n1147), .ZN(n1341) );
INV_X1 U1106 ( .A(G953), .ZN(n1147) );
NAND2_X1 U1107 ( .A1(n1393), .A2(n1394), .ZN(n1389) );
NAND2_X1 U1108 ( .A1(n1395), .A2(n1332), .ZN(n1394) );
XOR2_X1 U1109 ( .A(KEYINPUT10), .B(n1396), .Z(n1393) );
NOR2_X1 U1110 ( .A1(n1332), .A2(n1395), .ZN(n1396) );
XNOR2_X1 U1111 ( .A(KEYINPUT32), .B(n1293), .ZN(n1395) );
INV_X1 U1112 ( .A(G140), .ZN(n1293) );
INV_X1 U1113 ( .A(G125), .ZN(n1332) );
INV_X1 U1114 ( .A(n1299), .ZN(n1319) );
NAND2_X1 U1115 ( .A1(n1397), .A2(n1398), .ZN(n1299) );
OR2_X1 U1116 ( .A1(n1399), .A2(G472), .ZN(n1398) );
XOR2_X1 U1117 ( .A(n1400), .B(KEYINPUT43), .Z(n1397) );
NAND2_X1 U1118 ( .A1(G472), .A2(n1399), .ZN(n1400) );
XOR2_X1 U1119 ( .A(n1137), .B(KEYINPUT60), .Z(n1399) );
INV_X1 U1120 ( .A(n1144), .ZN(n1137) );
NAND2_X1 U1121 ( .A1(n1401), .A2(n1250), .ZN(n1144) );
INV_X1 U1122 ( .A(G902), .ZN(n1250) );
XOR2_X1 U1123 ( .A(n1214), .B(n1402), .Z(n1401) );
XNOR2_X1 U1124 ( .A(n1216), .B(n1403), .ZN(n1402) );
NOR2_X1 U1125 ( .A1(KEYINPUT12), .A2(n1404), .ZN(n1403) );
XNOR2_X1 U1126 ( .A(n1405), .B(n1224), .ZN(n1404) );
INV_X1 U1127 ( .A(n1211), .ZN(n1224) );
XNOR2_X1 U1128 ( .A(n1357), .B(G131), .ZN(n1211) );
NAND2_X1 U1129 ( .A1(KEYINPUT56), .A2(n1169), .ZN(n1357) );
XOR2_X1 U1130 ( .A(G134), .B(n1406), .Z(n1169) );
XOR2_X1 U1131 ( .A(KEYINPUT33), .B(G137), .Z(n1406) );
XNOR2_X1 U1132 ( .A(n1407), .B(n1210), .ZN(n1405) );
INV_X1 U1133 ( .A(n1184), .ZN(n1210) );
XOR2_X1 U1134 ( .A(G113), .B(n1408), .Z(n1184) );
XNOR2_X1 U1135 ( .A(G119), .B(n1312), .ZN(n1408) );
INV_X1 U1136 ( .A(G116), .ZN(n1312) );
NAND2_X1 U1137 ( .A1(KEYINPUT4), .A2(n1208), .ZN(n1407) );
INV_X1 U1138 ( .A(n1245), .ZN(n1208) );
XOR2_X1 U1139 ( .A(G128), .B(n1409), .Z(n1245) );
NOR2_X1 U1140 ( .A1(KEYINPUT39), .A2(n1410), .ZN(n1409) );
XNOR2_X1 U1141 ( .A(G146), .B(n1411), .ZN(n1410) );
NOR2_X1 U1142 ( .A1(G143), .A2(KEYINPUT29), .ZN(n1411) );
INV_X1 U1143 ( .A(G101), .ZN(n1216) );
AND2_X1 U1144 ( .A1(n1326), .A2(G210), .ZN(n1214) );
NOR2_X1 U1145 ( .A1(G953), .A2(G237), .ZN(n1326) );
endmodule


