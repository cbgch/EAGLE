//Key = 1111100111001111000011001111100111100110111001100000001010000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
n1375, n1376, n1377, n1378, n1379;

XOR2_X1 U759 ( .A(n1035), .B(n1036), .Z(G9) );
NOR2_X1 U760 ( .A1(n1037), .A2(n1038), .ZN(G75) );
NOR4_X1 U761 ( .A1(G953), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1038) );
NOR2_X1 U762 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U763 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U764 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U765 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U766 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U767 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U768 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR3_X1 U769 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1048) );
NOR2_X1 U770 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U771 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
XOR2_X1 U772 ( .A(KEYINPUT8), .B(n1062), .Z(n1061) );
NOR3_X1 U773 ( .A1(n1051), .A2(n1063), .A3(n1057), .ZN(n1044) );
INV_X1 U774 ( .A(n1064), .ZN(n1057) );
NOR2_X1 U775 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR3_X1 U776 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NOR3_X1 U777 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
AND2_X1 U778 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
INV_X1 U779 ( .A(n1075), .ZN(n1070) );
NOR2_X1 U780 ( .A1(n1076), .A2(n1075), .ZN(n1068) );
NOR2_X1 U781 ( .A1(n1077), .A2(n1047), .ZN(n1065) );
INV_X1 U782 ( .A(n1076), .ZN(n1047) );
NOR3_X1 U783 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n1037) );
AND4_X1 U784 ( .A1(n1078), .A2(n1075), .A3(n1079), .A4(n1080), .ZN(n1039) );
NOR3_X1 U785 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1080) );
XNOR2_X1 U786 ( .A(KEYINPUT35), .B(n1084), .ZN(n1083) );
XNOR2_X1 U787 ( .A(G478), .B(n1085), .ZN(n1082) );
NAND2_X1 U788 ( .A1(KEYINPUT34), .A2(n1086), .ZN(n1085) );
INV_X1 U789 ( .A(n1087), .ZN(n1086) );
NAND3_X1 U790 ( .A1(n1088), .A2(n1089), .A3(n1074), .ZN(n1081) );
XOR2_X1 U791 ( .A(n1090), .B(n1091), .Z(n1089) );
XOR2_X1 U792 ( .A(n1092), .B(KEYINPUT3), .Z(n1091) );
XOR2_X1 U793 ( .A(G469), .B(n1093), .Z(n1088) );
NOR2_X1 U794 ( .A1(n1094), .A2(KEYINPUT36), .ZN(n1093) );
INV_X1 U795 ( .A(n1095), .ZN(n1094) );
NOR3_X1 U796 ( .A1(n1096), .A2(n1062), .A3(n1097), .ZN(n1079) );
INV_X1 U797 ( .A(n1098), .ZN(n1096) );
XOR2_X1 U798 ( .A(n1099), .B(n1100), .Z(G72) );
XOR2_X1 U799 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U800 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U801 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U802 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U803 ( .A(n1109), .B(n1110), .Z(n1105) );
NOR3_X1 U804 ( .A1(KEYINPUT57), .A2(n1111), .A3(n1112), .ZN(n1110) );
NOR2_X1 U805 ( .A1(KEYINPUT55), .A2(n1113), .ZN(n1112) );
XOR2_X1 U806 ( .A(n1114), .B(G137), .Z(n1113) );
NOR2_X1 U807 ( .A1(n1115), .A2(n1116), .ZN(n1111) );
INV_X1 U808 ( .A(KEYINPUT55), .ZN(n1116) );
NOR2_X1 U809 ( .A1(G137), .A2(n1114), .ZN(n1115) );
XOR2_X1 U810 ( .A(n1117), .B(n1118), .Z(n1109) );
NOR2_X1 U811 ( .A1(n1119), .A2(n1120), .ZN(n1103) );
XOR2_X1 U812 ( .A(KEYINPUT51), .B(G900), .Z(n1120) );
NAND2_X1 U813 ( .A1(n1119), .A2(n1121), .ZN(n1101) );
NAND2_X1 U814 ( .A1(G953), .A2(n1122), .ZN(n1099) );
NAND2_X1 U815 ( .A1(G900), .A2(G227), .ZN(n1122) );
NAND2_X1 U816 ( .A1(n1123), .A2(n1124), .ZN(G69) );
NAND2_X1 U817 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U818 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NAND3_X1 U819 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
NAND2_X1 U820 ( .A1(G953), .A2(n1132), .ZN(n1130) );
NAND3_X1 U821 ( .A1(n1133), .A2(n1127), .A3(n1134), .ZN(n1123) );
NAND2_X1 U822 ( .A1(n1131), .A2(n1129), .ZN(n1134) );
INV_X1 U823 ( .A(n1135), .ZN(n1129) );
NAND3_X1 U824 ( .A1(n1135), .A2(n1119), .A3(n1136), .ZN(n1127) );
XOR2_X1 U825 ( .A(KEYINPUT27), .B(n1131), .Z(n1136) );
AND2_X1 U826 ( .A1(n1137), .A2(n1138), .ZN(n1131) );
NAND2_X1 U827 ( .A1(G953), .A2(n1139), .ZN(n1138) );
XOR2_X1 U828 ( .A(n1140), .B(n1141), .Z(n1137) );
NAND2_X1 U829 ( .A1(KEYINPUT45), .A2(n1142), .ZN(n1140) );
INV_X1 U830 ( .A(n1143), .ZN(n1142) );
NAND2_X1 U831 ( .A1(n1144), .A2(n1126), .ZN(n1133) );
INV_X1 U832 ( .A(KEYINPUT5), .ZN(n1126) );
NAND2_X1 U833 ( .A1(G953), .A2(n1145), .ZN(n1144) );
NAND2_X1 U834 ( .A1(G898), .A2(G224), .ZN(n1145) );
NOR2_X1 U835 ( .A1(n1146), .A2(n1147), .ZN(G66) );
XOR2_X1 U836 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U837 ( .A1(n1150), .A2(n1151), .ZN(n1148) );
NOR2_X1 U838 ( .A1(n1146), .A2(n1152), .ZN(G63) );
XOR2_X1 U839 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U840 ( .A1(n1150), .A2(G478), .ZN(n1153) );
NOR2_X1 U841 ( .A1(n1146), .A2(n1155), .ZN(G60) );
XOR2_X1 U842 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U843 ( .A1(n1150), .A2(G475), .ZN(n1156) );
XOR2_X1 U844 ( .A(n1158), .B(n1159), .Z(G6) );
NOR2_X1 U845 ( .A1(n1146), .A2(n1160), .ZN(G57) );
XOR2_X1 U846 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U847 ( .A(n1163), .B(KEYINPUT39), .ZN(n1162) );
NAND2_X1 U848 ( .A1(n1164), .A2(KEYINPUT12), .ZN(n1163) );
XNOR2_X1 U849 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U850 ( .A1(n1150), .A2(G472), .ZN(n1165) );
NOR2_X1 U851 ( .A1(n1146), .A2(n1167), .ZN(G54) );
XOR2_X1 U852 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U853 ( .A1(n1170), .A2(n1150), .ZN(n1169) );
INV_X1 U854 ( .A(n1171), .ZN(n1150) );
XOR2_X1 U855 ( .A(n1172), .B(KEYINPUT13), .Z(n1170) );
NAND2_X1 U856 ( .A1(n1173), .A2(n1174), .ZN(n1168) );
NAND2_X1 U857 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U858 ( .A(KEYINPUT14), .B(n1177), .Z(n1173) );
NOR2_X1 U859 ( .A1(n1176), .A2(n1175), .ZN(n1177) );
XNOR2_X1 U860 ( .A(n1178), .B(n1179), .ZN(n1175) );
NAND2_X1 U861 ( .A1(KEYINPUT62), .A2(n1180), .ZN(n1178) );
NOR2_X1 U862 ( .A1(n1181), .A2(n1182), .ZN(G51) );
XNOR2_X1 U863 ( .A(n1146), .B(KEYINPUT28), .ZN(n1182) );
NOR2_X1 U864 ( .A1(n1119), .A2(G952), .ZN(n1146) );
XOR2_X1 U865 ( .A(n1183), .B(n1184), .Z(n1181) );
NOR2_X1 U866 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U867 ( .A(KEYINPUT47), .B(n1187), .Z(n1186) );
XOR2_X1 U868 ( .A(n1188), .B(n1189), .Z(n1183) );
NOR3_X1 U869 ( .A1(n1171), .A2(KEYINPUT53), .A3(n1092), .ZN(n1189) );
NAND2_X1 U870 ( .A1(G902), .A2(n1041), .ZN(n1171) );
OR2_X1 U871 ( .A1(n1135), .A2(n1121), .ZN(n1041) );
NAND4_X1 U872 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1121) );
AND4_X1 U873 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
NAND2_X1 U874 ( .A1(KEYINPUT0), .A2(n1198), .ZN(n1192) );
NAND2_X1 U875 ( .A1(n1059), .A2(n1199), .ZN(n1191) );
XOR2_X1 U876 ( .A(KEYINPUT48), .B(n1200), .Z(n1199) );
NAND2_X1 U877 ( .A1(n1201), .A2(n1202), .ZN(n1190) );
NAND3_X1 U878 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
NAND2_X1 U879 ( .A1(KEYINPUT18), .A2(n1206), .ZN(n1205) );
NAND4_X1 U880 ( .A1(n1207), .A2(n1208), .A3(n1077), .A4(n1209), .ZN(n1204) );
INV_X1 U881 ( .A(KEYINPUT0), .ZN(n1209) );
NAND2_X1 U882 ( .A1(n1210), .A2(n1211), .ZN(n1203) );
NAND2_X1 U883 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
OR2_X1 U884 ( .A1(n1054), .A2(KEYINPUT18), .ZN(n1213) );
INV_X1 U885 ( .A(n1214), .ZN(n1054) );
NAND2_X1 U886 ( .A1(n1215), .A2(n1216), .ZN(n1135) );
NOR4_X1 U887 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
INV_X1 U888 ( .A(n1221), .ZN(n1220) );
AND4_X1 U889 ( .A1(n1222), .A2(n1036), .A3(n1159), .A4(n1223), .ZN(n1215) );
NAND3_X1 U890 ( .A1(n1053), .A2(n1224), .A3(n1071), .ZN(n1223) );
INV_X1 U891 ( .A(n1225), .ZN(n1224) );
NAND2_X1 U892 ( .A1(n1226), .A2(n1227), .ZN(n1159) );
NAND2_X1 U893 ( .A1(n1214), .A2(n1227), .ZN(n1036) );
AND2_X1 U894 ( .A1(n1228), .A2(n1076), .ZN(n1227) );
XOR2_X1 U895 ( .A(n1229), .B(n1230), .Z(G48) );
NAND2_X1 U896 ( .A1(n1200), .A2(n1059), .ZN(n1230) );
AND2_X1 U897 ( .A1(n1231), .A2(n1226), .ZN(n1200) );
XNOR2_X1 U898 ( .A(G143), .B(n1197), .ZN(G45) );
NAND4_X1 U899 ( .A1(n1210), .A2(n1059), .A3(n1232), .A4(n1233), .ZN(n1197) );
XOR2_X1 U900 ( .A(n1117), .B(n1234), .Z(G42) );
NOR2_X1 U901 ( .A1(n1235), .A2(KEYINPUT43), .ZN(n1234) );
INV_X1 U902 ( .A(n1196), .ZN(n1235) );
NAND4_X1 U903 ( .A1(n1201), .A2(n1236), .A3(n1226), .A4(n1237), .ZN(n1196) );
INV_X1 U904 ( .A(n1212), .ZN(n1226) );
XOR2_X1 U905 ( .A(G137), .B(n1198), .Z(G39) );
AND3_X1 U906 ( .A1(n1231), .A2(n1064), .A3(n1201), .ZN(n1198) );
INV_X1 U907 ( .A(n1051), .ZN(n1201) );
XOR2_X1 U908 ( .A(n1114), .B(n1238), .Z(G36) );
OR2_X1 U909 ( .A1(n1206), .A2(n1051), .ZN(n1238) );
NAND2_X1 U910 ( .A1(n1210), .A2(n1214), .ZN(n1206) );
INV_X1 U911 ( .A(n1239), .ZN(n1210) );
XOR2_X1 U912 ( .A(G131), .B(n1240), .Z(G33) );
NOR4_X1 U913 ( .A1(KEYINPUT60), .A2(n1212), .A3(n1051), .A4(n1239), .ZN(n1240) );
NAND3_X1 U914 ( .A1(n1237), .A2(n1208), .A3(n1071), .ZN(n1239) );
NAND2_X1 U915 ( .A1(n1241), .A2(n1242), .ZN(n1051) );
XOR2_X1 U916 ( .A(n1243), .B(KEYINPUT49), .Z(n1241) );
XOR2_X1 U917 ( .A(n1195), .B(n1244), .Z(G30) );
NOR2_X1 U918 ( .A1(G128), .A2(KEYINPUT10), .ZN(n1244) );
NAND3_X1 U919 ( .A1(n1214), .A2(n1059), .A3(n1231), .ZN(n1195) );
AND4_X1 U920 ( .A1(n1237), .A2(n1245), .A3(n1208), .A4(n1073), .ZN(n1231) );
INV_X1 U921 ( .A(n1077), .ZN(n1237) );
XOR2_X1 U922 ( .A(n1246), .B(n1222), .Z(G3) );
NAND3_X1 U923 ( .A1(n1064), .A2(n1228), .A3(n1071), .ZN(n1222) );
XNOR2_X1 U924 ( .A(G125), .B(n1194), .ZN(G27) );
NAND3_X1 U925 ( .A1(n1053), .A2(n1059), .A3(n1236), .ZN(n1194) );
AND3_X1 U926 ( .A1(n1208), .A2(n1073), .A3(n1074), .ZN(n1236) );
NAND2_X1 U927 ( .A1(n1043), .A2(n1247), .ZN(n1208) );
NAND4_X1 U928 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1249), .ZN(n1247) );
INV_X1 U929 ( .A(G900), .ZN(n1249) );
XOR2_X1 U930 ( .A(n1250), .B(n1221), .Z(G24) );
NAND4_X1 U931 ( .A1(n1251), .A2(n1076), .A3(n1232), .A4(n1233), .ZN(n1221) );
NOR2_X1 U932 ( .A1(n1073), .A2(n1245), .ZN(n1076) );
XOR2_X1 U933 ( .A(G119), .B(n1219), .Z(G21) );
AND2_X1 U934 ( .A1(n1207), .A2(n1251), .ZN(n1219) );
AND3_X1 U935 ( .A1(n1245), .A2(n1073), .A3(n1064), .ZN(n1207) );
INV_X1 U936 ( .A(n1074), .ZN(n1245) );
XNOR2_X1 U937 ( .A(n1218), .B(n1252), .ZN(G18) );
NAND2_X1 U938 ( .A1(KEYINPUT41), .A2(G116), .ZN(n1252) );
AND3_X1 U939 ( .A1(n1251), .A2(n1214), .A3(n1071), .ZN(n1218) );
NOR2_X1 U940 ( .A1(n1253), .A2(n1254), .ZN(n1214) );
NOR2_X1 U941 ( .A1(n1055), .A2(n1225), .ZN(n1251) );
NAND3_X1 U942 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(G15) );
NAND2_X1 U943 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND2_X1 U944 ( .A1(KEYINPUT23), .A2(n1260), .ZN(n1256) );
NAND2_X1 U945 ( .A1(n1261), .A2(G113), .ZN(n1260) );
XNOR2_X1 U946 ( .A(n1258), .B(KEYINPUT63), .ZN(n1261) );
NAND2_X1 U947 ( .A1(n1262), .A2(n1263), .ZN(n1255) );
INV_X1 U948 ( .A(KEYINPUT23), .ZN(n1263) );
NAND2_X1 U949 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
OR3_X1 U950 ( .A1(n1259), .A2(n1258), .A3(KEYINPUT63), .ZN(n1265) );
NAND2_X1 U951 ( .A1(KEYINPUT63), .A2(n1258), .ZN(n1264) );
AND4_X1 U952 ( .A1(n1266), .A2(n1053), .A3(n1071), .A4(n1267), .ZN(n1258) );
NOR2_X1 U953 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U954 ( .A1(n1212), .A2(n1055), .ZN(n1053) );
NAND2_X1 U955 ( .A1(n1268), .A2(n1075), .ZN(n1055) );
NAND2_X1 U956 ( .A1(n1233), .A2(n1254), .ZN(n1212) );
INV_X1 U957 ( .A(n1232), .ZN(n1254) );
XNOR2_X1 U958 ( .A(n1253), .B(KEYINPUT40), .ZN(n1233) );
XNOR2_X1 U959 ( .A(n1059), .B(KEYINPUT61), .ZN(n1266) );
XOR2_X1 U960 ( .A(n1217), .B(n1269), .Z(G12) );
NOR2_X1 U961 ( .A1(KEYINPUT11), .A2(n1270), .ZN(n1269) );
AND4_X1 U962 ( .A1(n1064), .A2(n1228), .A3(n1074), .A4(n1073), .ZN(n1217) );
NAND2_X1 U963 ( .A1(n1271), .A2(n1078), .ZN(n1073) );
NAND2_X1 U964 ( .A1(n1151), .A2(n1272), .ZN(n1078) );
NAND2_X1 U965 ( .A1(n1149), .A2(n1273), .ZN(n1272) );
INV_X1 U966 ( .A(n1274), .ZN(n1151) );
XNOR2_X1 U967 ( .A(n1097), .B(KEYINPUT44), .ZN(n1271) );
AND3_X1 U968 ( .A1(n1274), .A2(n1273), .A3(n1149), .ZN(n1097) );
XOR2_X1 U969 ( .A(n1275), .B(n1276), .Z(n1149) );
XOR2_X1 U970 ( .A(G137), .B(n1277), .Z(n1276) );
AND3_X1 U971 ( .A1(G221), .A2(n1119), .A3(G234), .ZN(n1277) );
NAND3_X1 U972 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1275) );
NAND2_X1 U973 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U974 ( .A1(KEYINPUT46), .A2(n1283), .ZN(n1282) );
XOR2_X1 U975 ( .A(KEYINPUT52), .B(n1284), .Z(n1283) );
NAND3_X1 U976 ( .A1(KEYINPUT46), .A2(n1285), .A3(n1284), .ZN(n1279) );
INV_X1 U977 ( .A(n1281), .ZN(n1285) );
XNOR2_X1 U978 ( .A(G125), .B(n1286), .ZN(n1281) );
XOR2_X1 U979 ( .A(G146), .B(G140), .Z(n1286) );
OR2_X1 U980 ( .A1(n1284), .A2(KEYINPUT46), .ZN(n1278) );
XNOR2_X1 U981 ( .A(n1287), .B(n1288), .ZN(n1284) );
XOR2_X1 U982 ( .A(G128), .B(G119), .Z(n1288) );
NAND2_X1 U983 ( .A1(KEYINPUT56), .A2(n1270), .ZN(n1287) );
INV_X1 U984 ( .A(G110), .ZN(n1270) );
NAND2_X1 U985 ( .A1(G217), .A2(n1289), .ZN(n1274) );
XOR2_X1 U986 ( .A(n1290), .B(G472), .Z(n1074) );
NAND3_X1 U987 ( .A1(n1291), .A2(n1292), .A3(n1273), .ZN(n1290) );
NAND2_X1 U988 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XOR2_X1 U989 ( .A(n1166), .B(n1161), .Z(n1293) );
OR3_X1 U990 ( .A1(n1166), .A2(n1161), .A3(n1294), .ZN(n1291) );
INV_X1 U991 ( .A(KEYINPUT6), .ZN(n1294) );
XNOR2_X1 U992 ( .A(n1295), .B(G101), .ZN(n1161) );
NAND2_X1 U993 ( .A1(G210), .A2(n1296), .ZN(n1295) );
XOR2_X1 U994 ( .A(n1297), .B(n1298), .Z(n1166) );
XOR2_X1 U995 ( .A(n1299), .B(n1300), .Z(n1297) );
NAND3_X1 U996 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1299) );
XOR2_X1 U997 ( .A(n1304), .B(KEYINPUT29), .Z(n1303) );
NAND2_X1 U998 ( .A1(G113), .A2(n1305), .ZN(n1304) );
XOR2_X1 U999 ( .A(G119), .B(G116), .Z(n1305) );
OR2_X1 U1000 ( .A1(n1306), .A2(G116), .ZN(n1302) );
NAND2_X1 U1001 ( .A1(n1307), .A2(G116), .ZN(n1301) );
INV_X1 U1002 ( .A(n1308), .ZN(n1307) );
NOR2_X1 U1003 ( .A1(n1225), .A2(n1077), .ZN(n1228) );
NAND2_X1 U1004 ( .A1(n1067), .A2(n1075), .ZN(n1077) );
NAND2_X1 U1005 ( .A1(G221), .A2(n1289), .ZN(n1075) );
NAND2_X1 U1006 ( .A1(G234), .A2(n1273), .ZN(n1289) );
INV_X1 U1007 ( .A(n1268), .ZN(n1067) );
XOR2_X1 U1008 ( .A(n1172), .B(n1309), .Z(n1268) );
NOR2_X1 U1009 ( .A1(KEYINPUT22), .A2(n1095), .ZN(n1309) );
NAND2_X1 U1010 ( .A1(n1310), .A2(n1273), .ZN(n1095) );
XOR2_X1 U1011 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U1012 ( .A(n1180), .B(n1313), .Z(n1312) );
NOR2_X1 U1013 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
AND2_X1 U1014 ( .A1(KEYINPUT42), .A2(n1316), .ZN(n1315) );
NOR2_X1 U1015 ( .A1(KEYINPUT38), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U1016 ( .A(n1176), .B(n1317), .ZN(n1316) );
XOR2_X1 U1017 ( .A(KEYINPUT58), .B(KEYINPUT15), .Z(n1317) );
XNOR2_X1 U1018 ( .A(n1318), .B(n1319), .ZN(n1176) );
XOR2_X1 U1019 ( .A(G101), .B(n1320), .Z(n1319) );
XOR2_X1 U1020 ( .A(G107), .B(G104), .Z(n1320) );
XOR2_X1 U1021 ( .A(n1321), .B(n1322), .Z(n1318) );
XNOR2_X1 U1022 ( .A(n1300), .B(n1118), .ZN(n1321) );
NOR2_X1 U1023 ( .A1(KEYINPUT16), .A2(G143), .ZN(n1118) );
XOR2_X1 U1024 ( .A(G137), .B(n1107), .Z(n1300) );
XOR2_X1 U1025 ( .A(G131), .B(G146), .Z(n1107) );
XOR2_X1 U1026 ( .A(G110), .B(G140), .Z(n1180) );
XNOR2_X1 U1027 ( .A(n1179), .B(KEYINPUT7), .ZN(n1311) );
AND2_X1 U1028 ( .A1(G227), .A2(n1119), .ZN(n1179) );
INV_X1 U1029 ( .A(G469), .ZN(n1172) );
NAND2_X1 U1030 ( .A1(n1059), .A2(n1267), .ZN(n1225) );
NAND2_X1 U1031 ( .A1(n1043), .A2(n1323), .ZN(n1267) );
NAND4_X1 U1032 ( .A1(G953), .A2(G902), .A3(n1248), .A4(n1139), .ZN(n1323) );
INV_X1 U1033 ( .A(G898), .ZN(n1139) );
NAND3_X1 U1034 ( .A1(n1248), .A2(n1119), .A3(n1324), .ZN(n1043) );
XNOR2_X1 U1035 ( .A(G952), .B(KEYINPUT2), .ZN(n1324) );
NAND2_X1 U1036 ( .A1(G237), .A2(G234), .ZN(n1248) );
NOR2_X1 U1037 ( .A1(n1242), .A2(n1062), .ZN(n1059) );
INV_X1 U1038 ( .A(n1243), .ZN(n1062) );
NAND2_X1 U1039 ( .A1(G214), .A2(n1325), .ZN(n1243) );
INV_X1 U1040 ( .A(n1060), .ZN(n1242) );
NAND2_X1 U1041 ( .A1(n1326), .A2(n1327), .ZN(n1060) );
NAND2_X1 U1042 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
XOR2_X1 U1043 ( .A(KEYINPUT26), .B(n1330), .Z(n1326) );
NOR2_X1 U1044 ( .A1(n1328), .A2(n1329), .ZN(n1330) );
XOR2_X1 U1045 ( .A(n1090), .B(KEYINPUT30), .Z(n1329) );
NAND2_X1 U1046 ( .A1(n1331), .A2(n1273), .ZN(n1090) );
XOR2_X1 U1047 ( .A(n1188), .B(n1332), .Z(n1331) );
OR2_X1 U1048 ( .A1(n1187), .A2(n1185), .ZN(n1332) );
AND2_X1 U1049 ( .A1(n1333), .A2(n1334), .ZN(n1185) );
NOR2_X1 U1050 ( .A1(n1334), .A2(n1333), .ZN(n1187) );
NOR2_X1 U1051 ( .A1(n1132), .A2(G953), .ZN(n1333) );
INV_X1 U1052 ( .A(G224), .ZN(n1132) );
XNOR2_X1 U1053 ( .A(n1335), .B(n1336), .ZN(n1334) );
XOR2_X1 U1054 ( .A(KEYINPUT31), .B(G146), .Z(n1336) );
XNOR2_X1 U1055 ( .A(G143), .B(n1108), .ZN(n1335) );
XOR2_X1 U1056 ( .A(G125), .B(G128), .Z(n1108) );
NAND2_X1 U1057 ( .A1(n1337), .A2(n1338), .ZN(n1188) );
NAND2_X1 U1058 ( .A1(n1143), .A2(n1141), .ZN(n1338) );
XOR2_X1 U1059 ( .A(KEYINPUT20), .B(n1339), .Z(n1337) );
NOR2_X1 U1060 ( .A1(n1143), .A2(n1141), .ZN(n1339) );
XNOR2_X1 U1061 ( .A(n1340), .B(n1341), .ZN(n1141) );
XOR2_X1 U1062 ( .A(n1342), .B(n1343), .Z(n1341) );
NAND2_X1 U1063 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
NAND2_X1 U1064 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
INV_X1 U1065 ( .A(n1348), .ZN(n1347) );
NAND2_X1 U1066 ( .A1(n1308), .A2(n1349), .ZN(n1346) );
NAND2_X1 U1067 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NAND2_X1 U1068 ( .A1(G119), .A2(n1259), .ZN(n1308) );
NAND2_X1 U1069 ( .A1(n1348), .A2(n1352), .ZN(n1344) );
NAND2_X1 U1070 ( .A1(n1353), .A2(n1306), .ZN(n1352) );
NAND2_X1 U1071 ( .A1(n1259), .A2(n1351), .ZN(n1306) );
INV_X1 U1072 ( .A(G119), .ZN(n1351) );
NAND2_X1 U1073 ( .A1(G119), .A2(n1350), .ZN(n1353) );
XOR2_X1 U1074 ( .A(n1259), .B(KEYINPUT9), .Z(n1350) );
INV_X1 U1075 ( .A(G113), .ZN(n1259) );
NOR2_X1 U1076 ( .A1(G116), .A2(KEYINPUT59), .ZN(n1348) );
NAND2_X1 U1077 ( .A1(n1354), .A2(KEYINPUT54), .ZN(n1342) );
XOR2_X1 U1078 ( .A(n1035), .B(n1355), .Z(n1354) );
NOR2_X1 U1079 ( .A1(KEYINPUT50), .A2(n1158), .ZN(n1355) );
INV_X1 U1080 ( .A(G104), .ZN(n1158) );
INV_X1 U1081 ( .A(G107), .ZN(n1035) );
XOR2_X1 U1082 ( .A(n1246), .B(KEYINPUT19), .Z(n1340) );
INV_X1 U1083 ( .A(G101), .ZN(n1246) );
XOR2_X1 U1084 ( .A(n1356), .B(G110), .Z(n1143) );
NAND2_X1 U1085 ( .A1(KEYINPUT1), .A2(n1250), .ZN(n1356) );
INV_X1 U1086 ( .A(n1092), .ZN(n1328) );
NAND2_X1 U1087 ( .A1(G210), .A2(n1325), .ZN(n1092) );
NAND2_X1 U1088 ( .A1(n1273), .A2(n1357), .ZN(n1325) );
INV_X1 U1089 ( .A(G237), .ZN(n1357) );
NOR2_X1 U1090 ( .A1(n1253), .A2(n1232), .ZN(n1064) );
XOR2_X1 U1091 ( .A(n1358), .B(G478), .Z(n1232) );
NAND2_X1 U1092 ( .A1(KEYINPUT33), .A2(n1087), .ZN(n1358) );
NAND2_X1 U1093 ( .A1(n1154), .A2(n1273), .ZN(n1087) );
XOR2_X1 U1094 ( .A(n1359), .B(n1360), .Z(n1154) );
XOR2_X1 U1095 ( .A(G116), .B(n1361), .Z(n1360) );
XOR2_X1 U1096 ( .A(KEYINPUT4), .B(G122), .Z(n1361) );
XNOR2_X1 U1097 ( .A(n1298), .B(n1362), .ZN(n1359) );
XOR2_X1 U1098 ( .A(G107), .B(n1363), .Z(n1362) );
AND3_X1 U1099 ( .A1(G234), .A2(n1119), .A3(G217), .ZN(n1363) );
INV_X1 U1100 ( .A(G953), .ZN(n1119) );
XOR2_X1 U1101 ( .A(G143), .B(n1322), .Z(n1298) );
XNOR2_X1 U1102 ( .A(G128), .B(n1114), .ZN(n1322) );
INV_X1 U1103 ( .A(G134), .ZN(n1114) );
NAND2_X1 U1104 ( .A1(n1098), .A2(n1084), .ZN(n1253) );
NAND3_X1 U1105 ( .A1(n1364), .A2(n1273), .A3(n1157), .ZN(n1084) );
XOR2_X1 U1106 ( .A(KEYINPUT32), .B(G475), .Z(n1364) );
NAND2_X1 U1107 ( .A1(n1365), .A2(n1366), .ZN(n1098) );
NAND2_X1 U1108 ( .A1(n1157), .A2(n1273), .ZN(n1366) );
INV_X1 U1109 ( .A(G902), .ZN(n1273) );
XOR2_X1 U1110 ( .A(n1367), .B(n1368), .Z(n1157) );
XOR2_X1 U1111 ( .A(G104), .B(n1369), .Z(n1368) );
NOR2_X1 U1112 ( .A1(KEYINPUT17), .A2(n1370), .ZN(n1369) );
XOR2_X1 U1113 ( .A(n1371), .B(n1372), .Z(n1370) );
XNOR2_X1 U1114 ( .A(n1373), .B(n1374), .ZN(n1372) );
NAND2_X1 U1115 ( .A1(KEYINPUT37), .A2(n1229), .ZN(n1374) );
INV_X1 U1116 ( .A(G146), .ZN(n1229) );
NAND2_X1 U1117 ( .A1(KEYINPUT24), .A2(n1375), .ZN(n1373) );
XOR2_X1 U1118 ( .A(n1376), .B(n1377), .Z(n1375) );
XNOR2_X1 U1119 ( .A(G131), .B(G143), .ZN(n1377) );
NAND2_X1 U1120 ( .A1(G214), .A2(n1296), .ZN(n1376) );
NOR2_X1 U1121 ( .A1(G953), .A2(G237), .ZN(n1296) );
XOR2_X1 U1122 ( .A(n1378), .B(G125), .Z(n1371) );
NAND2_X1 U1123 ( .A1(n1379), .A2(n1117), .ZN(n1378) );
INV_X1 U1124 ( .A(G140), .ZN(n1117) );
XNOR2_X1 U1125 ( .A(KEYINPUT25), .B(KEYINPUT21), .ZN(n1379) );
XOR2_X1 U1126 ( .A(n1250), .B(G113), .Z(n1367) );
INV_X1 U1127 ( .A(G122), .ZN(n1250) );
XNOR2_X1 U1128 ( .A(G475), .B(KEYINPUT32), .ZN(n1365) );
endmodule


