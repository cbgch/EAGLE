//Key = 0110111010010010110101100101110110111010101010110101000000011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;

XNOR2_X1 U725 ( .A(G107), .B(n999), .ZN(G9) );
NOR2_X1 U726 ( .A1(n1000), .A2(n1001), .ZN(G75) );
NOR4_X1 U727 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1001) );
XOR2_X1 U728 ( .A(n1006), .B(KEYINPUT35), .Z(n1004) );
NAND3_X1 U729 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
XOR2_X1 U730 ( .A(KEYINPUT37), .B(n1010), .Z(n1008) );
NOR2_X1 U731 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
XOR2_X1 U732 ( .A(KEYINPUT23), .B(n1013), .Z(n1012) );
NAND4_X1 U733 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1002) );
NAND4_X1 U734 ( .A1(n1018), .A2(n1019), .A3(n1007), .A4(n1020), .ZN(n1015) );
NAND2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U737 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U738 ( .A1(n1027), .A2(n1028), .ZN(n1021) );
NAND3_X1 U739 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
OR3_X1 U740 ( .A1(n1032), .A2(n1033), .A3(KEYINPUT63), .ZN(n1030) );
NAND2_X1 U741 ( .A1(KEYINPUT63), .A2(n1023), .ZN(n1029) );
NAND2_X1 U742 ( .A1(n1009), .A2(n1034), .ZN(n1014) );
NAND2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U744 ( .A1(n1019), .A2(n1037), .ZN(n1036) );
NAND2_X1 U745 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U747 ( .A1(n1007), .A2(n1042), .ZN(n1035) );
AND3_X1 U748 ( .A1(n1027), .A2(n1023), .A3(n1018), .ZN(n1009) );
INV_X1 U749 ( .A(n1043), .ZN(n1018) );
NOR3_X1 U750 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n1000) );
INV_X1 U751 ( .A(n1016), .ZN(n1044) );
NAND4_X1 U752 ( .A1(n1019), .A2(n1045), .A3(n1023), .A4(n1046), .ZN(n1016) );
NOR2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
XOR2_X1 U754 ( .A(n1049), .B(n1050), .Z(n1048) );
XNOR2_X1 U755 ( .A(G472), .B(KEYINPUT55), .ZN(n1050) );
XNOR2_X1 U756 ( .A(KEYINPUT40), .B(n1051), .ZN(n1045) );
XOR2_X1 U757 ( .A(n1052), .B(n1053), .Z(G72) );
XOR2_X1 U758 ( .A(n1054), .B(n1055), .Z(n1053) );
NAND2_X1 U759 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
INV_X1 U760 ( .A(n1058), .ZN(n1057) );
XOR2_X1 U761 ( .A(n1059), .B(n1060), .Z(n1056) );
XOR2_X1 U762 ( .A(n1061), .B(n1062), .Z(n1060) );
NAND3_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NAND2_X1 U764 ( .A1(KEYINPUT57), .A2(n1066), .ZN(n1065) );
NAND3_X1 U765 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1064) );
INV_X1 U766 ( .A(KEYINPUT57), .ZN(n1068) );
OR2_X1 U767 ( .A1(n1069), .A2(n1067), .ZN(n1063) );
NOR2_X1 U768 ( .A1(KEYINPUT53), .A2(n1066), .ZN(n1067) );
XNOR2_X1 U769 ( .A(G134), .B(G137), .ZN(n1066) );
NAND2_X1 U770 ( .A1(n1005), .A2(n1017), .ZN(n1054) );
NOR2_X1 U771 ( .A1(n1070), .A2(n1017), .ZN(n1052) );
AND2_X1 U772 ( .A1(G227), .A2(G900), .ZN(n1070) );
XOR2_X1 U773 ( .A(n1071), .B(n1072), .Z(G69) );
NOR2_X1 U774 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XOR2_X1 U775 ( .A(n1075), .B(KEYINPUT38), .Z(n1074) );
NAND3_X1 U776 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
INV_X1 U777 ( .A(n1079), .ZN(n1078) );
NAND2_X1 U778 ( .A1(n1080), .A2(n1017), .ZN(n1077) );
XOR2_X1 U779 ( .A(KEYINPUT52), .B(n1003), .Z(n1080) );
XOR2_X1 U780 ( .A(n1081), .B(n1082), .Z(n1076) );
NOR3_X1 U781 ( .A1(n1083), .A2(G953), .A3(n1084), .ZN(n1073) );
NOR2_X1 U782 ( .A1(n1085), .A2(n1079), .ZN(n1084) );
XOR2_X1 U783 ( .A(n1086), .B(KEYINPUT7), .Z(n1079) );
XNOR2_X1 U784 ( .A(n1081), .B(n1082), .ZN(n1085) );
XNOR2_X1 U785 ( .A(n1087), .B(n1088), .ZN(n1082) );
NOR2_X1 U786 ( .A1(KEYINPUT54), .A2(n1089), .ZN(n1088) );
NAND2_X1 U787 ( .A1(KEYINPUT17), .A2(n1090), .ZN(n1087) );
XNOR2_X1 U788 ( .A(KEYINPUT52), .B(n1003), .ZN(n1083) );
NAND2_X1 U789 ( .A1(G953), .A2(n1091), .ZN(n1071) );
NAND2_X1 U790 ( .A1(G898), .A2(G224), .ZN(n1091) );
NOR2_X1 U791 ( .A1(n1092), .A2(n1093), .ZN(G66) );
XOR2_X1 U792 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NOR2_X1 U794 ( .A1(n1092), .A2(n1098), .ZN(G63) );
XOR2_X1 U795 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U796 ( .A1(n1101), .A2(n1097), .ZN(n1099) );
NOR2_X1 U797 ( .A1(n1092), .A2(n1102), .ZN(G60) );
XNOR2_X1 U798 ( .A(n1103), .B(n1104), .ZN(n1102) );
NOR2_X1 U799 ( .A1(n1097), .A2(n1105), .ZN(n1104) );
XOR2_X1 U800 ( .A(KEYINPUT4), .B(G475), .Z(n1105) );
XNOR2_X1 U801 ( .A(G104), .B(n1106), .ZN(G6) );
NOR2_X1 U802 ( .A1(n1092), .A2(n1107), .ZN(G57) );
XOR2_X1 U803 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U804 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U805 ( .A1(n1112), .A2(n1097), .ZN(n1111) );
INV_X1 U806 ( .A(G472), .ZN(n1112) );
NOR2_X1 U807 ( .A1(KEYINPUT41), .A2(n1113), .ZN(n1110) );
XOR2_X1 U808 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U809 ( .A1(KEYINPUT60), .A2(n1116), .ZN(n1114) );
XOR2_X1 U810 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U811 ( .A1(KEYINPUT27), .A2(n1119), .ZN(n1117) );
NOR2_X1 U812 ( .A1(n1120), .A2(n1121), .ZN(n1108) );
XOR2_X1 U813 ( .A(KEYINPUT43), .B(n1122), .Z(n1121) );
NOR2_X1 U814 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U815 ( .A1(G101), .A2(n1125), .ZN(n1120) );
NOR2_X1 U816 ( .A1(n1092), .A2(n1126), .ZN(G54) );
XOR2_X1 U817 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U818 ( .A1(n1129), .A2(KEYINPUT26), .ZN(n1128) );
NOR2_X1 U819 ( .A1(n1130), .A2(n1097), .ZN(n1129) );
NAND2_X1 U820 ( .A1(n1131), .A2(n1132), .ZN(n1127) );
NAND2_X1 U821 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U822 ( .A(n1135), .B(KEYINPUT24), .Z(n1131) );
OR2_X1 U823 ( .A1(n1134), .A2(n1133), .ZN(n1135) );
XNOR2_X1 U824 ( .A(n1136), .B(n1059), .ZN(n1133) );
XNOR2_X1 U825 ( .A(n1137), .B(n1138), .ZN(n1136) );
NAND2_X1 U826 ( .A1(KEYINPUT34), .A2(n1139), .ZN(n1138) );
NAND2_X1 U827 ( .A1(KEYINPUT19), .A2(n1140), .ZN(n1137) );
XNOR2_X1 U828 ( .A(n1141), .B(n1142), .ZN(n1134) );
XNOR2_X1 U829 ( .A(KEYINPUT28), .B(n1143), .ZN(n1142) );
XNOR2_X1 U830 ( .A(n1144), .B(n1145), .ZN(n1141) );
NOR2_X1 U831 ( .A1(KEYINPUT18), .A2(n1146), .ZN(n1145) );
NOR2_X1 U832 ( .A1(KEYINPUT39), .A2(n1147), .ZN(n1144) );
INV_X1 U833 ( .A(n1148), .ZN(n1147) );
NOR2_X1 U834 ( .A1(n1092), .A2(n1149), .ZN(G51) );
XOR2_X1 U835 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U836 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U837 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U838 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XOR2_X1 U839 ( .A(n1158), .B(KEYINPUT58), .Z(n1154) );
OR2_X1 U840 ( .A1(n1157), .A2(n1156), .ZN(n1158) );
XOR2_X1 U841 ( .A(n1159), .B(n1160), .Z(n1157) );
NAND2_X1 U842 ( .A1(KEYINPUT44), .A2(n1118), .ZN(n1159) );
XOR2_X1 U843 ( .A(KEYINPUT47), .B(n1161), .Z(n1150) );
NOR2_X1 U844 ( .A1(n1162), .A2(n1097), .ZN(n1161) );
NAND2_X1 U845 ( .A1(n1163), .A2(n1164), .ZN(n1097) );
OR2_X1 U846 ( .A1(n1003), .A2(n1005), .ZN(n1164) );
NAND4_X1 U847 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1005) );
AND4_X1 U848 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1168) );
NOR2_X1 U849 ( .A1(n1173), .A2(n1174), .ZN(n1167) );
NOR3_X1 U850 ( .A1(n1175), .A2(n1051), .A3(n1176), .ZN(n1174) );
NAND3_X1 U851 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1175) );
NAND2_X1 U852 ( .A1(KEYINPUT5), .A2(n1180), .ZN(n1178) );
NAND2_X1 U853 ( .A1(n1181), .A2(n1182), .ZN(n1177) );
INV_X1 U854 ( .A(KEYINPUT5), .ZN(n1182) );
NAND3_X1 U855 ( .A1(n1019), .A2(n1183), .A3(n1184), .ZN(n1181) );
NAND2_X1 U856 ( .A1(n1185), .A2(n1186), .ZN(n1166) );
NAND2_X1 U857 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND3_X1 U858 ( .A1(n1189), .A2(n1031), .A3(KEYINPUT0), .ZN(n1188) );
NAND2_X1 U859 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
NAND2_X1 U860 ( .A1(n1192), .A2(n1193), .ZN(n1165) );
INV_X1 U861 ( .A(KEYINPUT0), .ZN(n1193) );
NAND4_X1 U862 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1003) );
AND4_X1 U863 ( .A1(n1106), .A2(n999), .A3(n1198), .A4(n1199), .ZN(n1197) );
NAND3_X1 U864 ( .A1(n1191), .A2(n1007), .A3(n1200), .ZN(n999) );
NAND3_X1 U865 ( .A1(n1200), .A2(n1007), .A3(n1179), .ZN(n1106) );
NOR2_X1 U866 ( .A1(n1201), .A2(n1202), .ZN(n1196) );
NOR2_X1 U867 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
XOR2_X1 U868 ( .A(n1205), .B(KEYINPUT56), .Z(n1203) );
INV_X1 U869 ( .A(n1206), .ZN(n1201) );
XNOR2_X1 U870 ( .A(KEYINPUT61), .B(n1207), .ZN(n1163) );
NOR2_X1 U871 ( .A1(n1017), .A2(G952), .ZN(n1092) );
XNOR2_X1 U872 ( .A(G146), .B(n1171), .ZN(G48) );
NAND2_X1 U873 ( .A1(n1208), .A2(n1179), .ZN(n1171) );
XOR2_X1 U874 ( .A(G143), .B(n1192), .Z(G45) );
AND3_X1 U875 ( .A1(n1185), .A2(n1183), .A3(n1189), .ZN(n1192) );
AND4_X1 U876 ( .A1(n1042), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1189) );
XNOR2_X1 U877 ( .A(G140), .B(n1212), .ZN(G42) );
NAND4_X1 U878 ( .A1(n1190), .A2(n1179), .A3(n1040), .A4(n1041), .ZN(n1212) );
XNOR2_X1 U879 ( .A(n1213), .B(n1173), .ZN(G39) );
AND3_X1 U880 ( .A1(n1176), .A2(n1214), .A3(n1190), .ZN(n1173) );
XNOR2_X1 U881 ( .A(n1215), .B(n1216), .ZN(G36) );
NOR3_X1 U882 ( .A1(n1217), .A2(n1026), .A3(n1180), .ZN(n1216) );
INV_X1 U883 ( .A(n1191), .ZN(n1026) );
XNOR2_X1 U884 ( .A(KEYINPUT59), .B(n1038), .ZN(n1217) );
INV_X1 U885 ( .A(n1185), .ZN(n1038) );
XNOR2_X1 U886 ( .A(G131), .B(n1172), .ZN(G33) );
NAND3_X1 U887 ( .A1(n1185), .A2(n1179), .A3(n1190), .ZN(n1172) );
INV_X1 U888 ( .A(n1180), .ZN(n1190) );
NAND3_X1 U889 ( .A1(n1183), .A2(n1211), .A3(n1019), .ZN(n1180) );
NOR2_X1 U890 ( .A1(n1013), .A2(n1218), .ZN(n1019) );
INV_X1 U891 ( .A(n1011), .ZN(n1218) );
XNOR2_X1 U892 ( .A(G128), .B(n1170), .ZN(G30) );
NAND2_X1 U893 ( .A1(n1208), .A2(n1191), .ZN(n1170) );
AND3_X1 U894 ( .A1(n1176), .A2(n1183), .A3(n1219), .ZN(n1208) );
XNOR2_X1 U895 ( .A(G101), .B(n1206), .ZN(G3) );
NAND3_X1 U896 ( .A1(n1027), .A2(n1200), .A3(n1185), .ZN(n1206) );
XNOR2_X1 U897 ( .A(G125), .B(n1169), .ZN(G27) );
NAND4_X1 U898 ( .A1(n1219), .A2(n1179), .A3(n1023), .A4(n1040), .ZN(n1169) );
NOR3_X1 U899 ( .A1(n1051), .A2(n1184), .A3(n1204), .ZN(n1219) );
INV_X1 U900 ( .A(n1211), .ZN(n1184) );
NAND2_X1 U901 ( .A1(n1043), .A2(n1220), .ZN(n1211) );
NAND3_X1 U902 ( .A1(G902), .A2(n1221), .A3(n1058), .ZN(n1220) );
NOR2_X1 U903 ( .A1(n1017), .A2(G900), .ZN(n1058) );
XNOR2_X1 U904 ( .A(G122), .B(n1194), .ZN(G24) );
NAND4_X1 U905 ( .A1(n1222), .A2(n1007), .A3(n1209), .A4(n1210), .ZN(n1194) );
NOR2_X1 U906 ( .A1(n1041), .A2(n1176), .ZN(n1007) );
XOR2_X1 U907 ( .A(n1223), .B(n1224), .Z(G21) );
XOR2_X1 U908 ( .A(KEYINPUT12), .B(G119), .Z(n1224) );
NOR2_X1 U909 ( .A1(n1204), .A2(n1205), .ZN(n1223) );
NAND4_X1 U910 ( .A1(n1176), .A2(n1214), .A3(n1023), .A4(n1225), .ZN(n1205) );
INV_X1 U911 ( .A(n1040), .ZN(n1176) );
XNOR2_X1 U912 ( .A(G116), .B(n1195), .ZN(G18) );
NAND3_X1 U913 ( .A1(n1222), .A2(n1191), .A3(n1185), .ZN(n1195) );
NOR2_X1 U914 ( .A1(n1210), .A2(n1226), .ZN(n1191) );
XNOR2_X1 U915 ( .A(G113), .B(n1199), .ZN(G15) );
NAND3_X1 U916 ( .A1(n1222), .A2(n1179), .A3(n1185), .ZN(n1199) );
NOR2_X1 U917 ( .A1(n1040), .A2(n1041), .ZN(n1185) );
INV_X1 U918 ( .A(n1025), .ZN(n1179) );
NAND2_X1 U919 ( .A1(n1226), .A2(n1210), .ZN(n1025) );
INV_X1 U920 ( .A(n1209), .ZN(n1226) );
AND3_X1 U921 ( .A1(n1042), .A2(n1225), .A3(n1023), .ZN(n1222) );
NOR2_X1 U922 ( .A1(n1033), .A2(n1227), .ZN(n1023) );
INV_X1 U923 ( .A(n1032), .ZN(n1227) );
XNOR2_X1 U924 ( .A(G110), .B(n1198), .ZN(G12) );
NAND3_X1 U925 ( .A1(n1200), .A2(n1040), .A3(n1214), .ZN(n1198) );
NOR2_X1 U926 ( .A1(n1047), .A2(n1051), .ZN(n1214) );
INV_X1 U927 ( .A(n1041), .ZN(n1051) );
XOR2_X1 U928 ( .A(n1228), .B(n1096), .Z(n1041) );
NAND2_X1 U929 ( .A1(G217), .A2(n1229), .ZN(n1096) );
OR2_X1 U930 ( .A1(n1095), .A2(G902), .ZN(n1228) );
XNOR2_X1 U931 ( .A(n1230), .B(n1231), .ZN(n1095) );
XNOR2_X1 U932 ( .A(n1232), .B(n1233), .ZN(n1231) );
NOR3_X1 U933 ( .A1(n1234), .A2(KEYINPUT9), .A3(n1235), .ZN(n1233) );
NOR2_X1 U934 ( .A1(G146), .A2(n1236), .ZN(n1235) );
XOR2_X1 U935 ( .A(n1237), .B(KEYINPUT21), .Z(n1234) );
NAND2_X1 U936 ( .A1(G146), .A2(n1236), .ZN(n1237) );
XNOR2_X1 U937 ( .A(n1062), .B(KEYINPUT50), .ZN(n1236) );
XNOR2_X1 U938 ( .A(G140), .B(G125), .ZN(n1062) );
NAND2_X1 U939 ( .A1(KEYINPUT11), .A2(n1238), .ZN(n1232) );
XNOR2_X1 U940 ( .A(G137), .B(n1239), .ZN(n1238) );
NAND2_X1 U941 ( .A1(n1240), .A2(G221), .ZN(n1239) );
XOR2_X1 U942 ( .A(n1241), .B(n1242), .Z(n1230) );
NOR2_X1 U943 ( .A1(KEYINPUT13), .A2(G128), .ZN(n1242) );
XNOR2_X1 U944 ( .A(G119), .B(G110), .ZN(n1241) );
INV_X1 U945 ( .A(n1027), .ZN(n1047) );
NOR2_X1 U946 ( .A1(n1209), .A2(n1210), .ZN(n1027) );
XNOR2_X1 U947 ( .A(n1243), .B(G475), .ZN(n1210) );
NAND2_X1 U948 ( .A1(n1103), .A2(n1207), .ZN(n1243) );
XNOR2_X1 U949 ( .A(n1244), .B(n1245), .ZN(n1103) );
XNOR2_X1 U950 ( .A(n1246), .B(n1247), .ZN(n1245) );
XOR2_X1 U951 ( .A(n1248), .B(n1249), .Z(n1247) );
AND2_X1 U952 ( .A1(G214), .A2(n1250), .ZN(n1249) );
NAND2_X1 U953 ( .A1(n1251), .A2(KEYINPUT8), .ZN(n1248) );
XNOR2_X1 U954 ( .A(n1252), .B(n1143), .ZN(n1251) );
NAND2_X1 U955 ( .A1(KEYINPUT36), .A2(n1160), .ZN(n1252) );
XOR2_X1 U956 ( .A(n1253), .B(n1254), .Z(n1244) );
XNOR2_X1 U957 ( .A(n1069), .B(G122), .ZN(n1254) );
INV_X1 U958 ( .A(G131), .ZN(n1069) );
XNOR2_X1 U959 ( .A(G104), .B(G113), .ZN(n1253) );
XOR2_X1 U960 ( .A(n1255), .B(n1101), .Z(n1209) );
INV_X1 U961 ( .A(G478), .ZN(n1101) );
OR2_X1 U962 ( .A1(n1100), .A2(G902), .ZN(n1255) );
XNOR2_X1 U963 ( .A(n1256), .B(n1257), .ZN(n1100) );
XOR2_X1 U964 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U965 ( .A(G128), .B(G122), .Z(n1259) );
XOR2_X1 U966 ( .A(KEYINPUT14), .B(G143), .Z(n1258) );
XOR2_X1 U967 ( .A(n1260), .B(n1261), .Z(n1256) );
XOR2_X1 U968 ( .A(n1262), .B(n1263), .Z(n1261) );
NAND2_X1 U969 ( .A1(KEYINPUT22), .A2(n1215), .ZN(n1263) );
INV_X1 U970 ( .A(G134), .ZN(n1215) );
NAND2_X1 U971 ( .A1(G217), .A2(n1240), .ZN(n1262) );
AND2_X1 U972 ( .A1(G234), .A2(n1017), .ZN(n1240) );
XOR2_X1 U973 ( .A(n1264), .B(G107), .Z(n1260) );
NAND2_X1 U974 ( .A1(KEYINPUT31), .A2(n1265), .ZN(n1264) );
INV_X1 U975 ( .A(G116), .ZN(n1265) );
XOR2_X1 U976 ( .A(G472), .B(n1266), .Z(n1040) );
NOR2_X1 U977 ( .A1(KEYINPUT30), .A2(n1267), .ZN(n1266) );
XNOR2_X1 U978 ( .A(KEYINPUT10), .B(n1049), .ZN(n1267) );
NAND2_X1 U979 ( .A1(n1268), .A2(n1269), .ZN(n1049) );
XNOR2_X1 U980 ( .A(KEYINPUT51), .B(n1207), .ZN(n1269) );
XOR2_X1 U981 ( .A(n1270), .B(n1271), .Z(n1268) );
XOR2_X1 U982 ( .A(n1118), .B(n1272), .Z(n1271) );
NAND2_X1 U983 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U984 ( .A1(n1275), .A2(n1119), .ZN(n1274) );
XNOR2_X1 U985 ( .A(KEYINPUT1), .B(n1124), .ZN(n1275) );
NAND2_X1 U986 ( .A1(n1276), .A2(n1139), .ZN(n1273) );
XNOR2_X1 U987 ( .A(n1125), .B(KEYINPUT32), .ZN(n1276) );
INV_X1 U988 ( .A(n1124), .ZN(n1125) );
NAND2_X1 U989 ( .A1(n1250), .A2(G210), .ZN(n1124) );
NOR2_X1 U990 ( .A1(G953), .A2(G237), .ZN(n1250) );
XOR2_X1 U991 ( .A(n1277), .B(n1278), .Z(n1270) );
XNOR2_X1 U992 ( .A(G101), .B(KEYINPUT45), .ZN(n1278) );
NAND2_X1 U993 ( .A1(n1279), .A2(n1115), .ZN(n1277) );
XNOR2_X1 U994 ( .A(G113), .B(n1280), .ZN(n1115) );
XNOR2_X1 U995 ( .A(KEYINPUT6), .B(KEYINPUT2), .ZN(n1279) );
AND3_X1 U996 ( .A1(n1183), .A2(n1225), .A3(n1042), .ZN(n1200) );
INV_X1 U997 ( .A(n1204), .ZN(n1042) );
NAND2_X1 U998 ( .A1(n1013), .A2(n1011), .ZN(n1204) );
NAND2_X1 U999 ( .A1(G214), .A2(n1281), .ZN(n1011) );
XOR2_X1 U1000 ( .A(n1282), .B(n1162), .Z(n1013) );
NAND2_X1 U1001 ( .A1(G210), .A2(n1281), .ZN(n1162) );
NAND2_X1 U1002 ( .A1(n1283), .A2(n1207), .ZN(n1281) );
INV_X1 U1003 ( .A(G237), .ZN(n1283) );
NAND2_X1 U1004 ( .A1(n1284), .A2(n1207), .ZN(n1282) );
XOR2_X1 U1005 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U1006 ( .A(n1152), .B(n1156), .Z(n1286) );
AND2_X1 U1007 ( .A1(G224), .A2(n1017), .ZN(n1156) );
NAND2_X1 U1008 ( .A1(n1287), .A2(n1288), .ZN(n1152) );
NAND2_X1 U1009 ( .A1(n1289), .A2(n1090), .ZN(n1288) );
XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n1290), .Z(n1287) );
NOR2_X1 U1011 ( .A1(n1090), .A2(n1289), .ZN(n1290) );
XNOR2_X1 U1012 ( .A(n1081), .B(n1089), .ZN(n1289) );
XNOR2_X1 U1013 ( .A(n1291), .B(n1292), .ZN(n1089) );
NOR2_X1 U1014 ( .A1(KEYINPUT48), .A2(n1280), .ZN(n1292) );
XNOR2_X1 U1015 ( .A(G116), .B(G119), .ZN(n1280) );
INV_X1 U1016 ( .A(G113), .ZN(n1291) );
XNOR2_X1 U1017 ( .A(n1293), .B(n1294), .ZN(n1081) );
NAND2_X1 U1018 ( .A1(KEYINPUT29), .A2(n1123), .ZN(n1293) );
INV_X1 U1019 ( .A(G101), .ZN(n1123) );
XNOR2_X1 U1020 ( .A(G110), .B(G122), .ZN(n1090) );
NAND2_X1 U1021 ( .A1(n1295), .A2(n1296), .ZN(n1285) );
NAND2_X1 U1022 ( .A1(n1297), .A2(n1160), .ZN(n1296) );
INV_X1 U1023 ( .A(G125), .ZN(n1160) );
NAND2_X1 U1024 ( .A1(n1118), .A2(n1298), .ZN(n1297) );
OR2_X1 U1025 ( .A1(n1299), .A2(KEYINPUT42), .ZN(n1298) );
NAND3_X1 U1026 ( .A1(n1300), .A2(n1301), .A3(KEYINPUT42), .ZN(n1295) );
NAND2_X1 U1027 ( .A1(KEYINPUT25), .A2(n1302), .ZN(n1301) );
NAND2_X1 U1028 ( .A1(G125), .A2(n1118), .ZN(n1302) );
NAND2_X1 U1029 ( .A1(n1118), .A2(n1299), .ZN(n1300) );
INV_X1 U1030 ( .A(KEYINPUT25), .ZN(n1299) );
XNOR2_X1 U1031 ( .A(G128), .B(n1246), .ZN(n1118) );
NAND2_X1 U1032 ( .A1(n1043), .A2(n1303), .ZN(n1225) );
NAND3_X1 U1033 ( .A1(n1086), .A2(n1221), .A3(G902), .ZN(n1303) );
AND2_X1 U1034 ( .A1(n1304), .A2(G953), .ZN(n1086) );
XNOR2_X1 U1035 ( .A(G898), .B(KEYINPUT33), .ZN(n1304) );
NAND3_X1 U1036 ( .A1(n1221), .A2(n1017), .A3(G952), .ZN(n1043) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1221) );
INV_X1 U1038 ( .A(n1031), .ZN(n1183) );
NAND2_X1 U1039 ( .A1(n1033), .A2(n1032), .ZN(n1031) );
NAND2_X1 U1040 ( .A1(G221), .A2(n1229), .ZN(n1032) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1207), .ZN(n1229) );
XOR2_X1 U1042 ( .A(n1305), .B(n1130), .Z(n1033) );
INV_X1 U1043 ( .A(G469), .ZN(n1130) );
NAND2_X1 U1044 ( .A1(n1306), .A2(n1207), .ZN(n1305) );
INV_X1 U1045 ( .A(G902), .ZN(n1207) );
XOR2_X1 U1046 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1047 ( .A(n1309), .B(n1310), .ZN(n1308) );
NOR2_X1 U1048 ( .A1(KEYINPUT20), .A2(n1148), .ZN(n1310) );
NAND2_X1 U1049 ( .A1(G227), .A2(n1017), .ZN(n1148) );
INV_X1 U1050 ( .A(G953), .ZN(n1017) );
NAND2_X1 U1051 ( .A1(KEYINPUT46), .A2(n1311), .ZN(n1309) );
XNOR2_X1 U1052 ( .A(n1059), .B(n1312), .ZN(n1311) );
XNOR2_X1 U1053 ( .A(n1140), .B(n1119), .ZN(n1312) );
INV_X1 U1054 ( .A(n1139), .ZN(n1119) );
XNOR2_X1 U1055 ( .A(n1313), .B(n1314), .ZN(n1139) );
NOR2_X1 U1056 ( .A1(KEYINPUT62), .A2(n1213), .ZN(n1314) );
INV_X1 U1057 ( .A(G137), .ZN(n1213) );
XNOR2_X1 U1058 ( .A(G131), .B(G134), .ZN(n1313) );
XNOR2_X1 U1059 ( .A(G101), .B(n1294), .ZN(n1140) );
XNOR2_X1 U1060 ( .A(n1315), .B(G107), .ZN(n1294) );
INV_X1 U1061 ( .A(G104), .ZN(n1315) );
XNOR2_X1 U1062 ( .A(n1316), .B(n1246), .ZN(n1059) );
XOR2_X1 U1063 ( .A(G143), .B(G146), .Z(n1246) );
XNOR2_X1 U1064 ( .A(KEYINPUT16), .B(n1317), .ZN(n1316) );
NOR2_X1 U1065 ( .A1(G128), .A2(KEYINPUT15), .ZN(n1317) );
XNOR2_X1 U1066 ( .A(n1146), .B(n1318), .ZN(n1307) );
XNOR2_X1 U1067 ( .A(KEYINPUT3), .B(n1143), .ZN(n1318) );
INV_X1 U1068 ( .A(G140), .ZN(n1143) );
INV_X1 U1069 ( .A(G110), .ZN(n1146) );
endmodule


