//Key = 1101101000000110100111011010100110000001111101101100000001111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377;

XOR2_X1 U744 ( .A(G107), .B(n1036), .Z(G9) );
NOR2_X1 U745 ( .A1(KEYINPUT37), .A2(n1037), .ZN(n1036) );
NOR2_X1 U746 ( .A1(n1038), .A2(n1039), .ZN(G75) );
NOR4_X1 U747 ( .A1(G953), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1039) );
NOR3_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1041) );
XOR2_X1 U749 ( .A(n1046), .B(KEYINPUT20), .Z(n1045) );
NOR2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1044) );
NOR3_X1 U751 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NOR2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U753 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U754 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U757 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U758 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR3_X1 U759 ( .A1(n1066), .A2(n1054), .A3(n1067), .ZN(n1058) );
AND3_X1 U760 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1054) );
NAND2_X1 U761 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND2_X1 U762 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U763 ( .A1(n1075), .A2(n1066), .ZN(n1074) );
INV_X1 U764 ( .A(n1076), .ZN(n1073) );
NAND2_X1 U765 ( .A1(n1077), .A2(n1078), .ZN(n1068) );
NAND2_X1 U766 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U767 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
INV_X1 U768 ( .A(KEYINPUT61), .ZN(n1066) );
NOR4_X1 U769 ( .A1(n1083), .A2(n1055), .A3(n1057), .A4(n1061), .ZN(n1047) );
NOR2_X1 U770 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
INV_X1 U771 ( .A(KEYINPUT19), .ZN(n1043) );
NOR3_X1 U772 ( .A1(n1040), .A2(G953), .A3(G952), .ZN(n1038) );
AND4_X1 U773 ( .A1(n1086), .A2(n1070), .A3(n1087), .A4(n1088), .ZN(n1040) );
NOR4_X1 U774 ( .A1(n1082), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1088) );
NOR2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
INV_X1 U776 ( .A(G478), .ZN(n1093) );
NOR2_X1 U777 ( .A1(G902), .A2(n1094), .ZN(n1092) );
NOR2_X1 U778 ( .A1(n1095), .A2(n1096), .ZN(n1087) );
XOR2_X1 U779 ( .A(n1097), .B(G472), .Z(n1086) );
XOR2_X1 U780 ( .A(n1098), .B(n1099), .Z(G72) );
NOR2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
AND2_X1 U782 ( .A1(G227), .A2(G900), .ZN(n1100) );
NAND2_X1 U783 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
NAND3_X1 U784 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
NAND2_X1 U785 ( .A1(G953), .A2(n1107), .ZN(n1105) );
OR2_X1 U786 ( .A1(n1106), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U787 ( .A(n1108), .B(n1109), .ZN(n1104) );
NOR2_X1 U788 ( .A1(KEYINPUT12), .A2(n1110), .ZN(n1109) );
XOR2_X1 U789 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U790 ( .A(n1113), .B(n1114), .Z(n1112) );
XNOR2_X1 U791 ( .A(KEYINPUT29), .B(n1115), .ZN(n1114) );
XNOR2_X1 U792 ( .A(n1116), .B(n1117), .ZN(n1111) );
NAND3_X1 U793 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1108) );
INV_X1 U794 ( .A(n1121), .ZN(n1120) );
OR2_X1 U795 ( .A1(G140), .A2(KEYINPUT48), .ZN(n1119) );
NAND2_X1 U796 ( .A1(n1122), .A2(KEYINPUT48), .ZN(n1118) );
NAND2_X1 U797 ( .A1(n1101), .A2(n1123), .ZN(n1106) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U799 ( .A(n1126), .B(n1127), .Z(G69) );
NOR2_X1 U800 ( .A1(n1128), .A2(n1101), .ZN(n1127) );
NOR2_X1 U801 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U802 ( .A1(n1131), .A2(n1132), .ZN(n1126) );
NAND2_X1 U803 ( .A1(n1133), .A2(n1101), .ZN(n1132) );
XNOR2_X1 U804 ( .A(n1134), .B(n1135), .ZN(n1133) );
NAND3_X1 U805 ( .A1(G898), .A2(n1135), .A3(G953), .ZN(n1131) );
NOR2_X1 U806 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XNOR2_X1 U807 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U808 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NOR2_X1 U809 ( .A1(n1136), .A2(n1142), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1143), .B(n1094), .ZN(n1142) );
NAND3_X1 U811 ( .A1(n1144), .A2(n1042), .A3(G478), .ZN(n1143) );
XNOR2_X1 U812 ( .A(KEYINPUT34), .B(n1145), .ZN(n1144) );
NOR2_X1 U813 ( .A1(n1136), .A2(n1146), .ZN(G60) );
XOR2_X1 U814 ( .A(n1147), .B(n1148), .Z(n1146) );
NOR2_X1 U815 ( .A1(KEYINPUT35), .A2(n1149), .ZN(n1148) );
XOR2_X1 U816 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U817 ( .A1(n1152), .A2(G475), .ZN(n1147) );
XNOR2_X1 U818 ( .A(G104), .B(n1153), .ZN(G6) );
NOR2_X1 U819 ( .A1(n1136), .A2(n1154), .ZN(G57) );
NOR2_X1 U820 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
XOR2_X1 U821 ( .A(KEYINPUT30), .B(n1157), .Z(n1156) );
NOR2_X1 U822 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U823 ( .A(KEYINPUT54), .B(n1160), .Z(n1159) );
NOR2_X1 U824 ( .A1(n1161), .A2(n1162), .ZN(n1155) );
INV_X1 U825 ( .A(n1158), .ZN(n1162) );
XOR2_X1 U826 ( .A(n1163), .B(n1164), .Z(n1158) );
XOR2_X1 U827 ( .A(n1165), .B(n1166), .Z(n1163) );
AND2_X1 U828 ( .A1(G472), .A2(n1152), .ZN(n1166) );
NAND2_X1 U829 ( .A1(KEYINPUT21), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U830 ( .A(KEYINPUT54), .B(n1160), .ZN(n1161) );
NOR2_X1 U831 ( .A1(n1136), .A2(n1168), .ZN(G54) );
XOR2_X1 U832 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U833 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U834 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U835 ( .A(n1175), .B(KEYINPUT58), .Z(n1174) );
INV_X1 U836 ( .A(G110), .ZN(n1173) );
NOR2_X1 U837 ( .A1(G110), .A2(n1176), .ZN(n1171) );
XNOR2_X1 U838 ( .A(KEYINPUT14), .B(n1175), .ZN(n1176) );
XNOR2_X1 U839 ( .A(n1177), .B(n1178), .ZN(n1169) );
AND2_X1 U840 ( .A1(G469), .A2(n1152), .ZN(n1178) );
INV_X1 U841 ( .A(n1141), .ZN(n1152) );
NOR2_X1 U842 ( .A1(n1136), .A2(n1179), .ZN(G51) );
XOR2_X1 U843 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U844 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U845 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U846 ( .A1(n1186), .A2(n1187), .ZN(n1184) );
NOR2_X1 U847 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
INV_X1 U848 ( .A(n1190), .ZN(n1188) );
NOR2_X1 U849 ( .A1(n1191), .A2(n1190), .ZN(n1186) );
XOR2_X1 U850 ( .A(KEYINPUT60), .B(n1189), .Z(n1191) );
NOR2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1182) );
XNOR2_X1 U852 ( .A(n1194), .B(n1189), .ZN(n1193) );
XOR2_X1 U853 ( .A(n1135), .B(KEYINPUT39), .Z(n1189) );
NAND2_X1 U854 ( .A1(n1190), .A2(KEYINPUT60), .ZN(n1194) );
XOR2_X1 U855 ( .A(n1195), .B(n1196), .Z(n1190) );
INV_X1 U856 ( .A(n1185), .ZN(n1192) );
NAND2_X1 U857 ( .A1(n1197), .A2(n1198), .ZN(n1185) );
XOR2_X1 U858 ( .A(KEYINPUT5), .B(KEYINPUT46), .Z(n1198) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1141), .ZN(n1180) );
NAND2_X1 U860 ( .A1(G902), .A2(n1042), .ZN(n1141) );
NAND3_X1 U861 ( .A1(n1124), .A2(n1200), .A3(n1134), .ZN(n1042) );
AND4_X1 U862 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1134) );
AND4_X1 U863 ( .A1(n1037), .A2(n1205), .A3(n1206), .A4(n1153), .ZN(n1204) );
NAND3_X1 U864 ( .A1(n1207), .A2(n1208), .A3(n1075), .ZN(n1153) );
NAND3_X1 U865 ( .A1(n1207), .A2(n1208), .A3(n1076), .ZN(n1037) );
NOR2_X1 U866 ( .A1(n1209), .A2(n1210), .ZN(n1203) );
NOR2_X1 U867 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U868 ( .A1(n1084), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U869 ( .A(n1085), .B(KEYINPUT6), .ZN(n1213) );
NOR4_X1 U870 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1209) );
XNOR2_X1 U871 ( .A(KEYINPUT49), .B(n1057), .ZN(n1217) );
NAND2_X1 U872 ( .A1(n1218), .A2(n1219), .ZN(n1202) );
INV_X1 U873 ( .A(KEYINPUT53), .ZN(n1219) );
NAND3_X1 U874 ( .A1(n1063), .A2(n1220), .A3(KEYINPUT53), .ZN(n1201) );
XOR2_X1 U875 ( .A(KEYINPUT44), .B(n1125), .Z(n1200) );
AND4_X1 U876 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1125) );
NOR2_X1 U877 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
AND4_X1 U878 ( .A1(KEYINPUT33), .A2(n1227), .A3(n1076), .A4(n1228), .ZN(n1226) );
AND3_X1 U879 ( .A1(n1229), .A2(n1230), .A3(n1208), .ZN(n1227) );
NOR2_X1 U880 ( .A1(KEYINPUT33), .A2(n1231), .ZN(n1225) );
AND4_X1 U881 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1124) );
NOR2_X1 U882 ( .A1(n1101), .A2(G952), .ZN(n1136) );
XNOR2_X1 U883 ( .A(G146), .B(n1232), .ZN(G48) );
NAND4_X1 U884 ( .A1(n1236), .A2(n1228), .A3(n1075), .A4(n1237), .ZN(n1232) );
XOR2_X1 U885 ( .A(n1233), .B(n1238), .Z(G45) );
XNOR2_X1 U886 ( .A(G143), .B(KEYINPUT47), .ZN(n1238) );
NAND3_X1 U887 ( .A1(n1236), .A2(n1084), .A3(n1239), .ZN(n1233) );
NOR3_X1 U888 ( .A1(n1079), .A2(n1214), .A3(n1215), .ZN(n1239) );
XNOR2_X1 U889 ( .A(G140), .B(n1234), .ZN(G42) );
NAND3_X1 U890 ( .A1(n1085), .A2(n1075), .A3(n1240), .ZN(n1234) );
XNOR2_X1 U891 ( .A(G137), .B(n1235), .ZN(G39) );
NAND3_X1 U892 ( .A1(n1228), .A2(n1077), .A3(n1240), .ZN(n1235) );
XNOR2_X1 U893 ( .A(G134), .B(n1222), .ZN(G36) );
NAND3_X1 U894 ( .A1(n1084), .A2(n1076), .A3(n1240), .ZN(n1222) );
XNOR2_X1 U895 ( .A(G131), .B(n1223), .ZN(G33) );
NAND3_X1 U896 ( .A1(n1075), .A2(n1084), .A3(n1240), .ZN(n1223) );
AND3_X1 U897 ( .A1(n1237), .A2(n1229), .A3(n1070), .ZN(n1240) );
INV_X1 U898 ( .A(n1055), .ZN(n1070) );
NAND2_X1 U899 ( .A1(n1241), .A2(n1065), .ZN(n1055) );
INV_X1 U900 ( .A(n1064), .ZN(n1241) );
INV_X1 U901 ( .A(n1079), .ZN(n1237) );
XNOR2_X1 U902 ( .A(G128), .B(n1231), .ZN(G30) );
NAND4_X1 U903 ( .A1(n1236), .A2(n1228), .A3(n1076), .A4(n1208), .ZN(n1231) );
XNOR2_X1 U904 ( .A(G101), .B(n1242), .ZN(G3) );
NAND2_X1 U905 ( .A1(n1243), .A2(n1084), .ZN(n1242) );
XNOR2_X1 U906 ( .A(G125), .B(n1224), .ZN(G27) );
NAND4_X1 U907 ( .A1(n1236), .A2(n1085), .A3(n1075), .A4(n1071), .ZN(n1224) );
AND2_X1 U908 ( .A1(n1063), .A2(n1229), .ZN(n1236) );
NAND2_X1 U909 ( .A1(n1244), .A2(n1245), .ZN(n1229) );
NAND2_X1 U910 ( .A1(n1246), .A2(n1107), .ZN(n1245) );
INV_X1 U911 ( .A(G900), .ZN(n1107) );
XNOR2_X1 U912 ( .A(G122), .B(n1247), .ZN(G24) );
NAND3_X1 U913 ( .A1(n1071), .A2(n1207), .A3(n1248), .ZN(n1247) );
NOR3_X1 U914 ( .A1(n1215), .A2(KEYINPUT51), .A3(n1214), .ZN(n1248) );
INV_X1 U915 ( .A(n1216), .ZN(n1207) );
NAND4_X1 U916 ( .A1(n1063), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1216) );
XNOR2_X1 U917 ( .A(G119), .B(n1206), .ZN(G21) );
NAND3_X1 U918 ( .A1(n1252), .A2(n1071), .A3(n1228), .ZN(n1206) );
NOR2_X1 U919 ( .A1(n1250), .A2(n1249), .ZN(n1228) );
XOR2_X1 U920 ( .A(n1253), .B(n1218), .Z(G18) );
NOR2_X1 U921 ( .A1(n1220), .A2(n1230), .ZN(n1218) );
NAND2_X1 U922 ( .A1(n1254), .A2(n1076), .ZN(n1220) );
NOR2_X1 U923 ( .A1(n1091), .A2(n1214), .ZN(n1076) );
NAND2_X1 U924 ( .A1(KEYINPUT16), .A2(n1255), .ZN(n1253) );
NAND2_X1 U925 ( .A1(n1256), .A2(n1257), .ZN(G15) );
OR2_X1 U926 ( .A1(n1205), .A2(G113), .ZN(n1257) );
XOR2_X1 U927 ( .A(n1258), .B(KEYINPUT56), .Z(n1256) );
NAND2_X1 U928 ( .A1(G113), .A2(n1205), .ZN(n1258) );
NAND3_X1 U929 ( .A1(n1254), .A2(n1063), .A3(n1075), .ZN(n1205) );
INV_X1 U930 ( .A(n1067), .ZN(n1075) );
NAND2_X1 U931 ( .A1(n1214), .A2(n1091), .ZN(n1067) );
AND3_X1 U932 ( .A1(n1084), .A2(n1251), .A3(n1071), .ZN(n1254) );
INV_X1 U933 ( .A(n1057), .ZN(n1071) );
NAND2_X1 U934 ( .A1(n1081), .A2(n1259), .ZN(n1057) );
INV_X1 U935 ( .A(n1095), .ZN(n1081) );
NOR2_X1 U936 ( .A1(n1249), .A2(n1051), .ZN(n1084) );
INV_X1 U937 ( .A(n1250), .ZN(n1051) );
XNOR2_X1 U938 ( .A(G110), .B(n1260), .ZN(G12) );
NAND2_X1 U939 ( .A1(n1243), .A2(n1085), .ZN(n1260) );
NOR2_X1 U940 ( .A1(n1250), .A2(n1049), .ZN(n1085) );
INV_X1 U941 ( .A(n1249), .ZN(n1049) );
XNOR2_X1 U942 ( .A(n1097), .B(n1261), .ZN(n1249) );
NOR2_X1 U943 ( .A1(G472), .A2(KEYINPUT22), .ZN(n1261) );
NAND2_X1 U944 ( .A1(n1262), .A2(n1145), .ZN(n1097) );
XOR2_X1 U945 ( .A(n1164), .B(n1263), .Z(n1262) );
XOR2_X1 U946 ( .A(n1160), .B(n1167), .Z(n1263) );
XNOR2_X1 U947 ( .A(n1195), .B(n1264), .ZN(n1167) );
XOR2_X1 U948 ( .A(n1265), .B(n1266), .Z(n1160) );
INV_X1 U949 ( .A(G101), .ZN(n1266) );
NAND3_X1 U950 ( .A1(n1267), .A2(n1101), .A3(G210), .ZN(n1265) );
NAND2_X1 U951 ( .A1(n1268), .A2(n1269), .ZN(n1164) );
NAND2_X1 U952 ( .A1(G119), .A2(n1270), .ZN(n1269) );
NAND2_X1 U953 ( .A1(n1271), .A2(n1272), .ZN(n1268) );
XNOR2_X1 U954 ( .A(n1273), .B(KEYINPUT3), .ZN(n1271) );
XOR2_X1 U955 ( .A(n1096), .B(KEYINPUT45), .Z(n1250) );
XOR2_X1 U956 ( .A(n1274), .B(n1140), .Z(n1096) );
NAND2_X1 U957 ( .A1(G217), .A2(n1275), .ZN(n1140) );
NAND2_X1 U958 ( .A1(n1276), .A2(n1139), .ZN(n1274) );
XOR2_X1 U959 ( .A(n1277), .B(n1278), .Z(n1139) );
XOR2_X1 U960 ( .A(n1279), .B(n1280), .Z(n1278) );
NAND2_X1 U961 ( .A1(KEYINPUT4), .A2(n1281), .ZN(n1280) );
XNOR2_X1 U962 ( .A(n1282), .B(G119), .ZN(n1281) );
NAND3_X1 U963 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1279) );
NAND2_X1 U964 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U965 ( .A1(n1288), .A2(n1289), .ZN(n1284) );
INV_X1 U966 ( .A(KEYINPUT1), .ZN(n1289) );
NAND2_X1 U967 ( .A1(n1290), .A2(n1291), .ZN(n1288) );
XNOR2_X1 U968 ( .A(KEYINPUT38), .B(n1287), .ZN(n1291) );
NAND2_X1 U969 ( .A1(KEYINPUT1), .A2(n1292), .ZN(n1283) );
NAND2_X1 U970 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
OR3_X1 U971 ( .A1(n1286), .A2(n1287), .A3(KEYINPUT38), .ZN(n1294) );
INV_X1 U972 ( .A(n1290), .ZN(n1286) );
NOR2_X1 U973 ( .A1(n1121), .A2(n1122), .ZN(n1290) );
NAND2_X1 U974 ( .A1(KEYINPUT38), .A2(n1287), .ZN(n1293) );
XNOR2_X1 U975 ( .A(G110), .B(n1295), .ZN(n1277) );
NOR2_X1 U976 ( .A1(KEYINPUT52), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U977 ( .A(G137), .B(n1297), .ZN(n1296) );
NAND2_X1 U978 ( .A1(G221), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U979 ( .A(G902), .B(KEYINPUT15), .ZN(n1276) );
INV_X1 U980 ( .A(n1212), .ZN(n1243) );
NAND2_X1 U981 ( .A1(n1252), .A2(n1208), .ZN(n1212) );
XNOR2_X1 U982 ( .A(n1079), .B(KEYINPUT62), .ZN(n1208) );
NAND2_X1 U983 ( .A1(n1259), .A2(n1095), .ZN(n1079) );
XNOR2_X1 U984 ( .A(n1299), .B(G469), .ZN(n1095) );
NAND2_X1 U985 ( .A1(n1300), .A2(n1145), .ZN(n1299) );
XOR2_X1 U986 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U987 ( .A(G110), .B(n1303), .ZN(n1302) );
XNOR2_X1 U988 ( .A(KEYINPUT25), .B(KEYINPUT18), .ZN(n1303) );
XNOR2_X1 U989 ( .A(n1304), .B(n1305), .ZN(n1301) );
INV_X1 U990 ( .A(n1177), .ZN(n1305) );
XNOR2_X1 U991 ( .A(n1306), .B(n1307), .ZN(n1177) );
XNOR2_X1 U992 ( .A(n1264), .B(n1117), .ZN(n1307) );
XNOR2_X1 U993 ( .A(n1308), .B(n1309), .ZN(n1117) );
NOR2_X1 U994 ( .A1(G128), .A2(KEYINPUT27), .ZN(n1309) );
XOR2_X1 U995 ( .A(n1310), .B(n1113), .Z(n1264) );
NAND2_X1 U996 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND2_X1 U997 ( .A1(n1313), .A2(n1115), .ZN(n1312) );
INV_X1 U998 ( .A(G137), .ZN(n1115) );
INV_X1 U999 ( .A(n1116), .ZN(n1313) );
XOR2_X1 U1000 ( .A(n1314), .B(KEYINPUT36), .Z(n1311) );
NAND2_X1 U1001 ( .A1(G137), .A2(n1116), .ZN(n1314) );
XOR2_X1 U1002 ( .A(G134), .B(KEYINPUT42), .Z(n1116) );
XNOR2_X1 U1003 ( .A(n1315), .B(n1316), .ZN(n1306) );
NAND2_X1 U1004 ( .A1(n1317), .A2(n1318), .ZN(n1315) );
OR2_X1 U1005 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XOR2_X1 U1006 ( .A(n1321), .B(KEYINPUT8), .Z(n1317) );
NAND2_X1 U1007 ( .A1(n1319), .A2(n1320), .ZN(n1321) );
NAND2_X1 U1008 ( .A1(KEYINPUT24), .A2(n1322), .ZN(n1304) );
XNOR2_X1 U1009 ( .A(KEYINPUT10), .B(n1175), .ZN(n1322) );
NAND2_X1 U1010 ( .A1(G227), .A2(n1101), .ZN(n1175) );
XOR2_X1 U1011 ( .A(KEYINPUT23), .B(n1082), .Z(n1259) );
AND2_X1 U1012 ( .A1(G221), .A2(n1275), .ZN(n1082) );
NAND2_X1 U1013 ( .A1(G234), .A2(n1145), .ZN(n1275) );
AND3_X1 U1014 ( .A1(n1063), .A2(n1251), .A3(n1077), .ZN(n1252) );
INV_X1 U1015 ( .A(n1061), .ZN(n1077) );
NAND2_X1 U1016 ( .A1(n1214), .A2(n1215), .ZN(n1061) );
INV_X1 U1017 ( .A(n1091), .ZN(n1215) );
XNOR2_X1 U1018 ( .A(n1323), .B(G475), .ZN(n1091) );
NAND2_X1 U1019 ( .A1(n1324), .A2(n1145), .ZN(n1323) );
XNOR2_X1 U1020 ( .A(n1151), .B(n1150), .ZN(n1324) );
XOR2_X1 U1021 ( .A(n1325), .B(n1326), .Z(n1150) );
XOR2_X1 U1022 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR3_X1 U1023 ( .A1(n1329), .A2(G953), .A3(n1330), .ZN(n1328) );
INV_X1 U1024 ( .A(G214), .ZN(n1330) );
XNOR2_X1 U1025 ( .A(KEYINPUT55), .B(n1267), .ZN(n1329) );
NOR2_X1 U1026 ( .A1(G113), .A2(KEYINPUT2), .ZN(n1327) );
XOR2_X1 U1027 ( .A(n1331), .B(G122), .Z(n1325) );
NAND3_X1 U1028 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1331) );
INV_X1 U1029 ( .A(n1122), .ZN(n1334) );
NOR2_X1 U1030 ( .A1(n1316), .A2(n1335), .ZN(n1122) );
INV_X1 U1031 ( .A(G140), .ZN(n1316) );
NAND2_X1 U1032 ( .A1(n1121), .A2(KEYINPUT26), .ZN(n1333) );
NOR2_X1 U1033 ( .A1(n1196), .A2(G140), .ZN(n1121) );
INV_X1 U1034 ( .A(n1335), .ZN(n1196) );
OR2_X1 U1035 ( .A1(n1335), .A2(KEYINPUT26), .ZN(n1332) );
XNOR2_X1 U1036 ( .A(n1308), .B(n1336), .ZN(n1151) );
XOR2_X1 U1037 ( .A(n1337), .B(n1113), .Z(n1336) );
XOR2_X1 U1038 ( .A(G131), .B(KEYINPUT59), .Z(n1113) );
XNOR2_X1 U1039 ( .A(G143), .B(G146), .ZN(n1308) );
NOR2_X1 U1040 ( .A1(n1338), .A2(n1089), .ZN(n1214) );
NOR3_X1 U1041 ( .A1(G478), .A2(G902), .A3(n1094), .ZN(n1089) );
AND2_X1 U1042 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
OR2_X1 U1043 ( .A1(n1094), .A2(G902), .ZN(n1340) );
XOR2_X1 U1044 ( .A(n1341), .B(n1342), .Z(n1094) );
XOR2_X1 U1045 ( .A(n1343), .B(n1344), .Z(n1342) );
NAND2_X1 U1046 ( .A1(G217), .A2(n1298), .ZN(n1344) );
AND2_X1 U1047 ( .A1(G234), .A2(n1101), .ZN(n1298) );
NAND2_X1 U1048 ( .A1(n1345), .A2(n1346), .ZN(n1343) );
NAND2_X1 U1049 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
XOR2_X1 U1050 ( .A(n1349), .B(KEYINPUT11), .Z(n1345) );
OR2_X1 U1051 ( .A1(n1348), .A2(n1347), .ZN(n1349) );
XNOR2_X1 U1052 ( .A(n1350), .B(G122), .ZN(n1347) );
NAND2_X1 U1053 ( .A1(KEYINPUT43), .A2(n1255), .ZN(n1350) );
XNOR2_X1 U1054 ( .A(G128), .B(n1351), .ZN(n1341) );
XNOR2_X1 U1055 ( .A(n1352), .B(G134), .ZN(n1351) );
INV_X1 U1056 ( .A(G143), .ZN(n1352) );
XNOR2_X1 U1057 ( .A(G478), .B(KEYINPUT32), .ZN(n1339) );
NAND2_X1 U1058 ( .A1(n1244), .A2(n1353), .ZN(n1251) );
NAND2_X1 U1059 ( .A1(n1246), .A2(n1130), .ZN(n1353) );
INV_X1 U1060 ( .A(G898), .ZN(n1130) );
AND3_X1 U1061 ( .A1(G902), .A2(n1046), .A3(G953), .ZN(n1246) );
NAND3_X1 U1062 ( .A1(n1046), .A2(n1101), .A3(n1354), .ZN(n1244) );
XNOR2_X1 U1063 ( .A(G952), .B(KEYINPUT19), .ZN(n1354) );
INV_X1 U1064 ( .A(G953), .ZN(n1101) );
NAND2_X1 U1065 ( .A1(G237), .A2(G234), .ZN(n1046) );
INV_X1 U1066 ( .A(n1230), .ZN(n1063) );
NAND2_X1 U1067 ( .A1(n1064), .A2(n1065), .ZN(n1230) );
NAND2_X1 U1068 ( .A1(G214), .A2(n1355), .ZN(n1065) );
XOR2_X1 U1069 ( .A(n1356), .B(n1199), .Z(n1064) );
NAND2_X1 U1070 ( .A1(G210), .A2(n1355), .ZN(n1199) );
NAND2_X1 U1071 ( .A1(n1145), .A2(n1267), .ZN(n1355) );
INV_X1 U1072 ( .A(G237), .ZN(n1267) );
NAND2_X1 U1073 ( .A1(n1357), .A2(n1145), .ZN(n1356) );
INV_X1 U1074 ( .A(G902), .ZN(n1145) );
XOR2_X1 U1075 ( .A(n1358), .B(KEYINPUT40), .Z(n1357) );
NAND2_X1 U1076 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
NAND2_X1 U1077 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
XOR2_X1 U1078 ( .A(KEYINPUT57), .B(n1363), .Z(n1359) );
NOR2_X1 U1079 ( .A1(n1361), .A2(n1362), .ZN(n1363) );
XNOR2_X1 U1080 ( .A(n1364), .B(n1335), .ZN(n1362) );
XOR2_X1 U1081 ( .A(G125), .B(KEYINPUT63), .Z(n1335) );
XOR2_X1 U1082 ( .A(n1365), .B(n1197), .Z(n1364) );
NOR2_X1 U1083 ( .A1(n1129), .A2(G953), .ZN(n1197) );
INV_X1 U1084 ( .A(G224), .ZN(n1129) );
NAND2_X1 U1085 ( .A1(KEYINPUT31), .A2(n1195), .ZN(n1365) );
XOR2_X1 U1086 ( .A(n1366), .B(n1367), .Z(n1195) );
NOR2_X1 U1087 ( .A1(KEYINPUT17), .A2(n1282), .ZN(n1367) );
INV_X1 U1088 ( .A(G128), .ZN(n1282) );
NAND2_X1 U1089 ( .A1(n1368), .A2(n1369), .ZN(n1366) );
NAND2_X1 U1090 ( .A1(n1370), .A2(n1287), .ZN(n1369) );
INV_X1 U1091 ( .A(G146), .ZN(n1287) );
XNOR2_X1 U1092 ( .A(G143), .B(KEYINPUT7), .ZN(n1370) );
NAND2_X1 U1093 ( .A1(n1371), .A2(G146), .ZN(n1368) );
XNOR2_X1 U1094 ( .A(G143), .B(KEYINPUT28), .ZN(n1371) );
INV_X1 U1095 ( .A(n1135), .ZN(n1361) );
XNOR2_X1 U1096 ( .A(n1372), .B(n1373), .ZN(n1135) );
XOR2_X1 U1097 ( .A(n1374), .B(n1375), .Z(n1373) );
XNOR2_X1 U1098 ( .A(n1272), .B(G110), .ZN(n1375) );
INV_X1 U1099 ( .A(G119), .ZN(n1272) );
XOR2_X1 U1100 ( .A(KEYINPUT50), .B(G122), .Z(n1374) );
XNOR2_X1 U1101 ( .A(n1376), .B(n1270), .ZN(n1372) );
INV_X1 U1102 ( .A(n1273), .ZN(n1270) );
XOR2_X1 U1103 ( .A(G113), .B(n1377), .Z(n1273) );
XNOR2_X1 U1104 ( .A(KEYINPUT13), .B(n1255), .ZN(n1377) );
INV_X1 U1105 ( .A(G116), .ZN(n1255) );
XNOR2_X1 U1106 ( .A(n1320), .B(n1319), .ZN(n1376) );
XOR2_X1 U1107 ( .A(n1348), .B(n1337), .Z(n1319) );
XOR2_X1 U1108 ( .A(G104), .B(KEYINPUT9), .Z(n1337) );
XOR2_X1 U1109 ( .A(G107), .B(KEYINPUT41), .Z(n1348) );
XOR2_X1 U1110 ( .A(G101), .B(KEYINPUT0), .Z(n1320) );
endmodule


