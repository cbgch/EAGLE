//Key = 0111001001111010000100000000010001011100111000100011010011101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322;

XNOR2_X1 U731 ( .A(G107), .B(n1015), .ZN(G9) );
NOR2_X1 U732 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
XOR2_X1 U736 ( .A(KEYINPUT31), .B(n1026), .Z(n1025) );
NOR3_X1 U737 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
NOR2_X1 U738 ( .A1(n1030), .A2(n1028), .ZN(n1024) );
NAND3_X1 U739 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1028) );
NAND3_X1 U740 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1018) );
NAND4_X1 U741 ( .A1(n1037), .A2(n1033), .A3(n1038), .A4(n1027), .ZN(n1036) );
NAND2_X1 U742 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND3_X1 U743 ( .A1(n1041), .A2(n1042), .A3(n1032), .ZN(n1040) );
OR2_X1 U744 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U745 ( .A1(n1031), .A2(n1045), .ZN(n1039) );
NAND3_X1 U746 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NAND2_X1 U747 ( .A1(n1049), .A2(n1041), .ZN(n1048) );
NAND2_X1 U748 ( .A1(n1032), .A2(n1050), .ZN(n1046) );
NAND2_X1 U749 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
XNOR2_X1 U751 ( .A(KEYINPUT45), .B(n1055), .ZN(n1053) );
INV_X1 U752 ( .A(n1056), .ZN(n1033) );
NOR3_X1 U753 ( .A1(n1057), .A2(G953), .A3(n1058), .ZN(n1016) );
INV_X1 U754 ( .A(n1034), .ZN(n1058) );
NAND4_X1 U755 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1034) );
NOR3_X1 U756 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
XOR2_X1 U757 ( .A(KEYINPUT8), .B(n1066), .Z(n1065) );
XNOR2_X1 U758 ( .A(G469), .B(n1067), .ZN(n1064) );
NAND3_X1 U759 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1063) );
XNOR2_X1 U760 ( .A(n1071), .B(G472), .ZN(n1070) );
XNOR2_X1 U761 ( .A(KEYINPUT40), .B(n1072), .ZN(n1069) );
NOR3_X1 U762 ( .A1(n1073), .A2(n1054), .A3(n1074), .ZN(n1061) );
AND2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND2_X1 U764 ( .A1(G475), .A2(n1077), .ZN(n1060) );
XOR2_X1 U765 ( .A(KEYINPUT46), .B(n1078), .Z(n1059) );
NOR2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1078) );
XNOR2_X1 U767 ( .A(n1079), .B(KEYINPUT23), .ZN(n1076) );
XNOR2_X1 U768 ( .A(KEYINPUT38), .B(n1021), .ZN(n1057) );
INV_X1 U769 ( .A(G952), .ZN(n1021) );
XOR2_X1 U770 ( .A(n1080), .B(n1081), .Z(G72) );
XOR2_X1 U771 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XOR2_X1 U773 ( .A(n1086), .B(n1087), .Z(n1085) );
XNOR2_X1 U774 ( .A(n1088), .B(n1089), .ZN(n1087) );
NAND2_X1 U775 ( .A1(KEYINPUT53), .A2(G140), .ZN(n1089) );
NAND2_X1 U776 ( .A1(n1090), .A2(KEYINPUT12), .ZN(n1088) );
XNOR2_X1 U777 ( .A(n1091), .B(n1092), .ZN(n1090) );
XOR2_X1 U778 ( .A(n1093), .B(KEYINPUT27), .Z(n1091) );
XNOR2_X1 U779 ( .A(G125), .B(KEYINPUT37), .ZN(n1086) );
NOR2_X1 U780 ( .A1(G900), .A2(n1035), .ZN(n1084) );
NAND3_X1 U781 ( .A1(KEYINPUT50), .A2(n1094), .A3(n1095), .ZN(n1082) );
XNOR2_X1 U782 ( .A(n1096), .B(n1035), .ZN(n1095) );
XNOR2_X1 U783 ( .A(KEYINPUT60), .B(KEYINPUT33), .ZN(n1096) );
NAND2_X1 U784 ( .A1(G953), .A2(n1097), .ZN(n1080) );
NAND2_X1 U785 ( .A1(G900), .A2(G227), .ZN(n1097) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(G69) );
XOR2_X1 U787 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U788 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U789 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XNOR2_X1 U790 ( .A(KEYINPUT63), .B(n1106), .ZN(n1105) );
XNOR2_X1 U791 ( .A(KEYINPUT14), .B(n1035), .ZN(n1102) );
NAND2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(n1100) );
NAND2_X1 U793 ( .A1(n1109), .A2(G953), .ZN(n1108) );
XNOR2_X1 U794 ( .A(G898), .B(KEYINPUT17), .ZN(n1109) );
XNOR2_X1 U795 ( .A(n1110), .B(n1111), .ZN(n1107) );
NOR2_X1 U796 ( .A1(n1112), .A2(n1035), .ZN(n1098) );
NOR2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XOR2_X1 U799 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1121), .ZN(G63) );
XNOR2_X1 U802 ( .A(n1122), .B(n1123), .ZN(n1121) );
AND2_X1 U803 ( .A1(G478), .A2(n1124), .ZN(n1122) );
NOR2_X1 U804 ( .A1(n1115), .A2(n1125), .ZN(G60) );
XOR2_X1 U805 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U806 ( .A1(KEYINPUT3), .A2(n1128), .ZN(n1126) );
NAND2_X1 U807 ( .A1(n1124), .A2(G475), .ZN(n1128) );
XNOR2_X1 U808 ( .A(G104), .B(n1129), .ZN(G6) );
NOR2_X1 U809 ( .A1(n1115), .A2(n1130), .ZN(G57) );
XOR2_X1 U810 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U811 ( .A(KEYINPUT18), .B(n1133), .Z(n1132) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1120), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1135), .A2(n1136), .ZN(G54) );
XNOR2_X1 U814 ( .A(n1115), .B(KEYINPUT11), .ZN(n1136) );
XOR2_X1 U815 ( .A(n1137), .B(n1138), .Z(n1135) );
XOR2_X1 U816 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U817 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NAND2_X1 U818 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U819 ( .A1(n1092), .A2(n1145), .ZN(n1144) );
NAND2_X1 U820 ( .A1(KEYINPUT54), .A2(KEYINPUT35), .ZN(n1145) );
NAND3_X1 U821 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1141) );
INV_X1 U822 ( .A(KEYINPUT54), .ZN(n1148) );
NAND2_X1 U823 ( .A1(KEYINPUT35), .A2(n1149), .ZN(n1147) );
NAND2_X1 U824 ( .A1(n1150), .A2(n1092), .ZN(n1149) );
OR2_X1 U825 ( .A1(n1151), .A2(KEYINPUT35), .ZN(n1146) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1137) );
AND2_X1 U827 ( .A1(G469), .A2(n1124), .ZN(n1153) );
INV_X1 U828 ( .A(n1120), .ZN(n1124) );
NAND2_X1 U829 ( .A1(n1154), .A2(n1155), .ZN(n1152) );
NAND2_X1 U830 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR2_X1 U831 ( .A1(n1115), .A2(n1158), .ZN(G51) );
XOR2_X1 U832 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR3_X1 U833 ( .A1(n1120), .A2(KEYINPUT47), .A3(n1075), .ZN(n1160) );
NAND2_X1 U834 ( .A1(G902), .A2(n1019), .ZN(n1120) );
NAND3_X1 U835 ( .A1(n1104), .A2(n1106), .A3(n1161), .ZN(n1019) );
INV_X1 U836 ( .A(n1094), .ZN(n1161) );
NAND4_X1 U837 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1094) );
NOR4_X1 U838 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
NAND2_X1 U839 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
NAND2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XNOR2_X1 U842 ( .A(n1176), .B(KEYINPUT10), .ZN(n1174) );
NAND4_X1 U843 ( .A1(n1049), .A2(n1177), .A3(n1178), .A4(n1043), .ZN(n1162) );
XNOR2_X1 U844 ( .A(n1023), .B(KEYINPUT4), .ZN(n1178) );
INV_X1 U845 ( .A(n1041), .ZN(n1023) );
AND4_X1 U846 ( .A1(n1179), .A2(n1129), .A3(n1180), .A4(n1181), .ZN(n1104) );
NOR4_X1 U847 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181) );
INV_X1 U848 ( .A(n1015), .ZN(n1185) );
NAND3_X1 U849 ( .A1(n1043), .A2(n1032), .A3(n1186), .ZN(n1015) );
NAND2_X1 U850 ( .A1(n1187), .A2(n1170), .ZN(n1180) );
NAND3_X1 U851 ( .A1(n1186), .A2(n1032), .A3(n1044), .ZN(n1129) );
NAND3_X1 U852 ( .A1(n1031), .A2(n1186), .A3(n1049), .ZN(n1179) );
NAND3_X1 U853 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1159) );
NAND2_X1 U854 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
INV_X1 U855 ( .A(KEYINPUT51), .ZN(n1192) );
NAND3_X1 U856 ( .A1(KEYINPUT51), .A2(n1193), .A3(n1194), .ZN(n1189) );
OR2_X1 U857 ( .A1(n1194), .A2(n1193), .ZN(n1188) );
NOR2_X1 U858 ( .A1(KEYINPUT5), .A2(n1191), .ZN(n1193) );
XNOR2_X1 U859 ( .A(n1195), .B(n1196), .ZN(n1191) );
NAND2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
NAND2_X1 U861 ( .A1(n1151), .A2(n1199), .ZN(n1198) );
XOR2_X1 U862 ( .A(n1200), .B(KEYINPUT39), .Z(n1197) );
NAND2_X1 U863 ( .A1(n1092), .A2(G125), .ZN(n1200) );
NOR2_X1 U864 ( .A1(n1035), .A2(G952), .ZN(n1115) );
XOR2_X1 U865 ( .A(n1201), .B(n1202), .Z(G48) );
AND3_X1 U866 ( .A1(n1175), .A2(n1170), .A3(n1176), .ZN(n1202) );
NOR2_X1 U867 ( .A1(KEYINPUT44), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U868 ( .A(n1163), .B(n1204), .ZN(G45) );
NOR2_X1 U869 ( .A1(KEYINPUT21), .A2(n1205), .ZN(n1204) );
NAND4_X1 U870 ( .A1(n1049), .A2(n1177), .A3(n1206), .A4(n1170), .ZN(n1163) );
NOR2_X1 U871 ( .A1(n1207), .A2(n1072), .ZN(n1206) );
XNOR2_X1 U872 ( .A(G140), .B(n1208), .ZN(G42) );
NAND2_X1 U873 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U874 ( .A1(KEYINPUT55), .A2(n1169), .ZN(n1210) );
OR2_X1 U875 ( .A1(KEYINPUT52), .A2(n1169), .ZN(n1209) );
NOR2_X1 U876 ( .A1(n1047), .A2(n1211), .ZN(n1169) );
NAND3_X1 U877 ( .A1(n1041), .A2(n1212), .A3(n1213), .ZN(n1047) );
XOR2_X1 U878 ( .A(G137), .B(n1168), .Z(G39) );
AND4_X1 U879 ( .A1(n1177), .A2(n1176), .A3(n1031), .A4(n1041), .ZN(n1168) );
XNOR2_X1 U880 ( .A(G134), .B(n1214), .ZN(G36) );
NAND4_X1 U881 ( .A1(n1215), .A2(n1049), .A3(n1177), .A4(n1043), .ZN(n1214) );
XNOR2_X1 U882 ( .A(KEYINPUT19), .B(n1041), .ZN(n1215) );
XOR2_X1 U883 ( .A(n1167), .B(n1216), .Z(G33) );
NOR2_X1 U884 ( .A1(KEYINPUT24), .A2(n1217), .ZN(n1216) );
INV_X1 U885 ( .A(G131), .ZN(n1217) );
AND3_X1 U886 ( .A1(n1175), .A2(n1041), .A3(n1049), .ZN(n1167) );
NAND2_X1 U887 ( .A1(n1218), .A2(n1219), .ZN(n1041) );
OR3_X1 U888 ( .A1(n1055), .A2(n1054), .A3(KEYINPUT45), .ZN(n1219) );
NAND2_X1 U889 ( .A1(KEYINPUT45), .A2(n1170), .ZN(n1218) );
INV_X1 U890 ( .A(n1211), .ZN(n1175) );
NAND2_X1 U891 ( .A1(n1044), .A2(n1177), .ZN(n1211) );
XOR2_X1 U892 ( .A(G128), .B(n1166), .Z(G30) );
AND4_X1 U893 ( .A1(n1177), .A2(n1176), .A3(n1043), .A4(n1170), .ZN(n1166) );
AND2_X1 U894 ( .A1(n1220), .A2(n1221), .ZN(n1177) );
XOR2_X1 U895 ( .A(n1222), .B(n1223), .Z(G3) );
NOR2_X1 U896 ( .A1(KEYINPUT13), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U897 ( .A(G101), .B(KEYINPUT1), .ZN(n1224) );
NAND4_X1 U898 ( .A1(n1049), .A2(n1031), .A3(n1225), .A4(n1170), .ZN(n1222) );
NOR2_X1 U899 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XNOR2_X1 U900 ( .A(n1220), .B(KEYINPUT59), .ZN(n1227) );
XOR2_X1 U901 ( .A(n1228), .B(n1229), .Z(G27) );
NAND2_X1 U902 ( .A1(KEYINPUT29), .A2(G125), .ZN(n1229) );
NAND2_X1 U903 ( .A1(n1170), .A2(n1230), .ZN(n1228) );
XNOR2_X1 U904 ( .A(KEYINPUT16), .B(n1172), .ZN(n1230) );
NAND4_X1 U905 ( .A1(n1231), .A2(n1213), .A3(n1212), .A4(n1221), .ZN(n1172) );
NAND2_X1 U906 ( .A1(n1056), .A2(n1232), .ZN(n1221) );
NAND4_X1 U907 ( .A1(G953), .A2(G902), .A3(n1233), .A4(n1234), .ZN(n1232) );
INV_X1 U908 ( .A(G900), .ZN(n1234) );
XNOR2_X1 U909 ( .A(G122), .B(n1235), .ZN(G24) );
NAND2_X1 U910 ( .A1(KEYINPUT58), .A2(n1184), .ZN(n1235) );
AND4_X1 U911 ( .A1(n1236), .A2(n1032), .A3(n1237), .A4(n1238), .ZN(n1184) );
NOR2_X1 U912 ( .A1(n1239), .A2(n1212), .ZN(n1032) );
XOR2_X1 U913 ( .A(G119), .B(n1183), .Z(G21) );
AND3_X1 U914 ( .A1(n1176), .A2(n1031), .A3(n1236), .ZN(n1183) );
NOR2_X1 U915 ( .A1(n1068), .A2(n1213), .ZN(n1176) );
INV_X1 U916 ( .A(n1212), .ZN(n1068) );
XNOR2_X1 U917 ( .A(n1240), .B(n1182), .ZN(G18) );
AND3_X1 U918 ( .A1(n1049), .A2(n1043), .A3(n1236), .ZN(n1182) );
NOR4_X1 U919 ( .A1(n1029), .A2(n1051), .A3(n1074), .A4(n1226), .ZN(n1236) );
NOR2_X1 U920 ( .A1(n1238), .A2(n1072), .ZN(n1043) );
INV_X1 U921 ( .A(n1237), .ZN(n1072) );
XNOR2_X1 U922 ( .A(G113), .B(n1241), .ZN(G15) );
NAND2_X1 U923 ( .A1(n1170), .A2(n1242), .ZN(n1241) );
XOR2_X1 U924 ( .A(KEYINPUT26), .B(n1187), .Z(n1242) );
AND3_X1 U925 ( .A1(n1049), .A2(n1243), .A3(n1231), .ZN(n1187) );
AND3_X1 U926 ( .A1(n1044), .A2(n1027), .A3(n1037), .ZN(n1231) );
NOR2_X1 U927 ( .A1(n1237), .A2(n1207), .ZN(n1044) );
NOR2_X1 U928 ( .A1(n1212), .A2(n1213), .ZN(n1049) );
XOR2_X1 U929 ( .A(G110), .B(n1244), .Z(G12) );
NOR2_X1 U930 ( .A1(KEYINPUT30), .A2(n1106), .ZN(n1244) );
NAND4_X1 U931 ( .A1(n1031), .A2(n1186), .A3(n1213), .A4(n1212), .ZN(n1106) );
XOR2_X1 U932 ( .A(n1245), .B(n1119), .Z(n1212) );
NAND2_X1 U933 ( .A1(G217), .A2(n1246), .ZN(n1119) );
OR2_X1 U934 ( .A1(n1118), .A2(G902), .ZN(n1245) );
XNOR2_X1 U935 ( .A(n1247), .B(n1248), .ZN(n1118) );
XOR2_X1 U936 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U937 ( .A(n1251), .B(n1252), .Z(n1250) );
AND3_X1 U938 ( .A1(G221), .A2(n1035), .A3(G234), .ZN(n1251) );
XOR2_X1 U939 ( .A(n1253), .B(n1254), .Z(n1247) );
NOR2_X1 U940 ( .A1(G137), .A2(KEYINPUT0), .ZN(n1254) );
XNOR2_X1 U941 ( .A(G119), .B(n1255), .ZN(n1253) );
NOR2_X1 U942 ( .A1(KEYINPUT61), .A2(n1256), .ZN(n1255) );
INV_X1 U943 ( .A(n1239), .ZN(n1213) );
NAND3_X1 U944 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1239) );
NAND2_X1 U945 ( .A1(G472), .A2(n1260), .ZN(n1259) );
OR3_X1 U946 ( .A1(n1260), .A2(G472), .A3(KEYINPUT22), .ZN(n1258) );
NOR2_X1 U947 ( .A1(n1071), .A2(KEYINPUT43), .ZN(n1260) );
NAND2_X1 U948 ( .A1(KEYINPUT22), .A2(n1261), .ZN(n1257) );
NAND2_X1 U949 ( .A1(n1071), .A2(n1134), .ZN(n1261) );
INV_X1 U950 ( .A(G472), .ZN(n1134) );
NOR2_X1 U951 ( .A1(n1131), .A2(G902), .ZN(n1071) );
XNOR2_X1 U952 ( .A(n1262), .B(n1263), .ZN(n1131) );
XOR2_X1 U953 ( .A(G101), .B(n1264), .Z(n1263) );
NOR2_X1 U954 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XOR2_X1 U955 ( .A(n1267), .B(KEYINPUT2), .Z(n1266) );
NAND2_X1 U956 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NOR2_X1 U957 ( .A1(n1269), .A2(n1268), .ZN(n1265) );
XNOR2_X1 U958 ( .A(n1270), .B(G119), .ZN(n1268) );
NAND2_X1 U959 ( .A1(KEYINPUT42), .A2(n1240), .ZN(n1270) );
INV_X1 U960 ( .A(G113), .ZN(n1269) );
XNOR2_X1 U961 ( .A(n1271), .B(n1272), .ZN(n1262) );
AND2_X1 U962 ( .A1(G210), .A2(n1273), .ZN(n1272) );
NOR3_X1 U963 ( .A1(n1030), .A2(n1226), .A3(n1051), .ZN(n1186) );
INV_X1 U964 ( .A(n1170), .ZN(n1051) );
NOR2_X1 U965 ( .A1(n1274), .A2(n1054), .ZN(n1170) );
AND2_X1 U966 ( .A1(G214), .A2(n1275), .ZN(n1054) );
INV_X1 U967 ( .A(n1055), .ZN(n1274) );
XOR2_X1 U968 ( .A(n1079), .B(n1075), .Z(n1055) );
NAND2_X1 U969 ( .A1(G210), .A2(n1275), .ZN(n1075) );
NAND2_X1 U970 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
INV_X1 U971 ( .A(G237), .ZN(n1277) );
XOR2_X1 U972 ( .A(KEYINPUT49), .B(n1278), .Z(n1276) );
NAND2_X1 U973 ( .A1(n1279), .A2(n1280), .ZN(n1079) );
XOR2_X1 U974 ( .A(n1281), .B(n1282), .Z(n1279) );
XNOR2_X1 U975 ( .A(n1199), .B(n1196), .ZN(n1282) );
NOR2_X1 U976 ( .A1(n1113), .A2(G953), .ZN(n1196) );
INV_X1 U977 ( .A(G224), .ZN(n1113) );
INV_X1 U978 ( .A(G125), .ZN(n1199) );
XNOR2_X1 U979 ( .A(n1194), .B(n1283), .ZN(n1281) );
NOR2_X1 U980 ( .A1(KEYINPUT34), .A2(n1151), .ZN(n1283) );
XOR2_X1 U981 ( .A(n1284), .B(n1285), .Z(n1194) );
INV_X1 U982 ( .A(n1110), .ZN(n1285) );
XNOR2_X1 U983 ( .A(n1286), .B(n1287), .ZN(n1110) );
XNOR2_X1 U984 ( .A(n1240), .B(n1288), .ZN(n1287) );
XOR2_X1 U985 ( .A(KEYINPUT9), .B(G119), .Z(n1288) );
XNOR2_X1 U986 ( .A(n1143), .B(G113), .ZN(n1286) );
NAND2_X1 U987 ( .A1(KEYINPUT36), .A2(n1111), .ZN(n1284) );
XNOR2_X1 U988 ( .A(G122), .B(n1252), .ZN(n1111) );
INV_X1 U989 ( .A(n1243), .ZN(n1226) );
NAND2_X1 U990 ( .A1(n1056), .A2(n1289), .ZN(n1243) );
NAND4_X1 U991 ( .A1(G953), .A2(G902), .A3(n1233), .A4(n1114), .ZN(n1289) );
INV_X1 U992 ( .A(G898), .ZN(n1114) );
NAND3_X1 U993 ( .A1(n1233), .A2(n1035), .A3(G952), .ZN(n1056) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1233) );
INV_X1 U995 ( .A(n1220), .ZN(n1030) );
NOR2_X1 U996 ( .A1(n1037), .A2(n1074), .ZN(n1220) );
INV_X1 U997 ( .A(n1027), .ZN(n1074) );
NAND2_X1 U998 ( .A1(G221), .A2(n1246), .ZN(n1027) );
NAND2_X1 U999 ( .A1(G234), .A2(n1278), .ZN(n1246) );
XNOR2_X1 U1000 ( .A(n1280), .B(KEYINPUT62), .ZN(n1278) );
INV_X1 U1001 ( .A(n1029), .ZN(n1037) );
XOR2_X1 U1002 ( .A(n1290), .B(n1067), .Z(n1029) );
NAND2_X1 U1003 ( .A1(n1291), .A2(n1280), .ZN(n1067) );
XOR2_X1 U1004 ( .A(n1292), .B(n1293), .Z(n1291) );
NAND2_X1 U1005 ( .A1(KEYINPUT56), .A2(n1294), .ZN(n1293) );
XNOR2_X1 U1006 ( .A(n1271), .B(n1150), .ZN(n1294) );
INV_X1 U1007 ( .A(n1143), .ZN(n1150) );
XOR2_X1 U1008 ( .A(G101), .B(n1295), .Z(n1143) );
XNOR2_X1 U1009 ( .A(n1296), .B(G104), .ZN(n1295) );
INV_X1 U1010 ( .A(G107), .ZN(n1296) );
XOR2_X1 U1011 ( .A(n1140), .B(n1092), .Z(n1271) );
INV_X1 U1012 ( .A(n1151), .ZN(n1092) );
XOR2_X1 U1013 ( .A(G143), .B(n1249), .Z(n1151) );
XNOR2_X1 U1014 ( .A(G128), .B(n1203), .ZN(n1249) );
INV_X1 U1015 ( .A(G146), .ZN(n1203) );
XOR2_X1 U1016 ( .A(n1093), .B(KEYINPUT57), .Z(n1140) );
XNOR2_X1 U1017 ( .A(G131), .B(n1297), .ZN(n1093) );
XOR2_X1 U1018 ( .A(G137), .B(G134), .Z(n1297) );
NAND3_X1 U1019 ( .A1(n1298), .A2(n1299), .A3(n1154), .ZN(n1292) );
OR2_X1 U1020 ( .A1(n1157), .A2(n1156), .ZN(n1154) );
OR2_X1 U1021 ( .A1(n1157), .A2(KEYINPUT6), .ZN(n1299) );
NAND3_X1 U1022 ( .A1(n1156), .A2(n1157), .A3(KEYINPUT6), .ZN(n1298) );
NAND2_X1 U1023 ( .A1(G227), .A2(n1035), .ZN(n1157) );
XNOR2_X1 U1024 ( .A(n1300), .B(n1252), .ZN(n1156) );
XOR2_X1 U1025 ( .A(G110), .B(KEYINPUT32), .Z(n1252) );
XNOR2_X1 U1026 ( .A(G140), .B(KEYINPUT25), .ZN(n1300) );
NAND2_X1 U1027 ( .A1(KEYINPUT41), .A2(G469), .ZN(n1290) );
NOR2_X1 U1028 ( .A1(n1237), .A2(n1238), .ZN(n1031) );
INV_X1 U1029 ( .A(n1207), .ZN(n1238) );
NOR2_X1 U1030 ( .A1(n1066), .A2(n1301), .ZN(n1207) );
AND2_X1 U1031 ( .A1(G475), .A2(n1077), .ZN(n1301) );
NOR2_X1 U1032 ( .A1(n1077), .A2(G475), .ZN(n1066) );
OR2_X1 U1033 ( .A1(n1127), .A2(G902), .ZN(n1077) );
XNOR2_X1 U1034 ( .A(n1302), .B(n1303), .ZN(n1127) );
XNOR2_X1 U1035 ( .A(n1304), .B(n1256), .ZN(n1303) );
XNOR2_X1 U1036 ( .A(G140), .B(G125), .ZN(n1256) );
NOR2_X1 U1037 ( .A1(KEYINPUT15), .A2(n1305), .ZN(n1304) );
XOR2_X1 U1038 ( .A(G122), .B(n1306), .Z(n1305) );
NOR2_X1 U1039 ( .A1(G113), .A2(KEYINPUT48), .ZN(n1306) );
XOR2_X1 U1040 ( .A(n1307), .B(n1308), .Z(n1302) );
NOR2_X1 U1041 ( .A1(KEYINPUT28), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1042 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1043 ( .A(G131), .B(G143), .ZN(n1311) );
NAND3_X1 U1044 ( .A1(n1273), .A2(G214), .A3(n1312), .ZN(n1310) );
XNOR2_X1 U1045 ( .A(KEYINPUT7), .B(KEYINPUT20), .ZN(n1312) );
NOR2_X1 U1046 ( .A1(G953), .A2(G237), .ZN(n1273) );
XNOR2_X1 U1047 ( .A(G104), .B(G146), .ZN(n1307) );
XNOR2_X1 U1048 ( .A(n1313), .B(G478), .ZN(n1237) );
NAND2_X1 U1049 ( .A1(n1123), .A2(n1280), .ZN(n1313) );
INV_X1 U1050 ( .A(G902), .ZN(n1280) );
NAND2_X1 U1051 ( .A1(n1314), .A2(n1315), .ZN(n1123) );
NAND2_X1 U1052 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND3_X1 U1053 ( .A1(G234), .A2(n1035), .A3(G217), .ZN(n1317) );
NAND4_X1 U1054 ( .A1(G234), .A2(n1035), .A3(G217), .A4(n1318), .ZN(n1314) );
INV_X1 U1055 ( .A(n1316), .ZN(n1318) );
XNOR2_X1 U1056 ( .A(n1319), .B(n1320), .ZN(n1316) );
XOR2_X1 U1057 ( .A(G128), .B(n1321), .Z(n1320) );
XNOR2_X1 U1058 ( .A(n1205), .B(G134), .ZN(n1321) );
INV_X1 U1059 ( .A(G143), .ZN(n1205) );
XNOR2_X1 U1060 ( .A(G107), .B(n1322), .ZN(n1319) );
XNOR2_X1 U1061 ( .A(G122), .B(n1240), .ZN(n1322) );
INV_X1 U1062 ( .A(G116), .ZN(n1240) );
INV_X1 U1063 ( .A(G953), .ZN(n1035) );
endmodule


