//Key = 1111011100100010011110111001011100011011111111011110100011000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278;

XNOR2_X1 U713 ( .A(G107), .B(n975), .ZN(G9) );
NAND2_X1 U714 ( .A1(n976), .A2(n977), .ZN(n975) );
XOR2_X1 U715 ( .A(n978), .B(KEYINPUT39), .Z(n976) );
NOR2_X1 U716 ( .A1(n979), .A2(n980), .ZN(G75) );
NOR4_X1 U717 ( .A1(n981), .A2(n982), .A3(n983), .A4(n984), .ZN(n980) );
XNOR2_X1 U718 ( .A(G952), .B(KEYINPUT4), .ZN(n983) );
NAND3_X1 U719 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n981) );
NAND2_X1 U720 ( .A1(n988), .A2(n989), .ZN(n987) );
NAND2_X1 U721 ( .A1(n990), .A2(n991), .ZN(n989) );
NAND3_X1 U722 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND2_X1 U723 ( .A1(n995), .A2(n996), .ZN(n993) );
NAND2_X1 U724 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U725 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U726 ( .A1(n1001), .A2(n1002), .ZN(n995) );
NAND2_X1 U727 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U728 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND3_X1 U729 ( .A1(n997), .A2(n1007), .A3(n1001), .ZN(n990) );
NAND3_X1 U730 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NAND2_X1 U731 ( .A1(n1011), .A2(n992), .ZN(n1010) );
NAND3_X1 U732 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1009) );
XNOR2_X1 U733 ( .A(n992), .B(KEYINPUT48), .ZN(n1014) );
NAND2_X1 U734 ( .A1(n994), .A2(n1015), .ZN(n1008) );
OR2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
INV_X1 U736 ( .A(n1018), .ZN(n988) );
NOR3_X1 U737 ( .A1(n1019), .A2(G953), .A3(G952), .ZN(n979) );
XNOR2_X1 U738 ( .A(KEYINPUT11), .B(n985), .ZN(n1019) );
NAND2_X1 U739 ( .A1(n1020), .A2(n1021), .ZN(n985) );
NOR4_X1 U740 ( .A1(n1005), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n1021) );
NOR2_X1 U741 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U742 ( .A1(G902), .A2(n1027), .ZN(n1025) );
NOR4_X1 U743 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1020) );
XOR2_X1 U744 ( .A(n1032), .B(n1033), .Z(G72) );
XOR2_X1 U745 ( .A(n1034), .B(n1035), .Z(n1033) );
NOR2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
XOR2_X1 U747 ( .A(n1038), .B(n1039), .Z(n1037) );
XOR2_X1 U748 ( .A(n1040), .B(n1041), .Z(n1039) );
XNOR2_X1 U749 ( .A(KEYINPUT31), .B(n1042), .ZN(n1038) );
NOR2_X1 U750 ( .A1(KEYINPUT21), .A2(n1043), .ZN(n1042) );
XOR2_X1 U751 ( .A(n1044), .B(n1045), .Z(n1043) );
NAND2_X1 U752 ( .A1(KEYINPUT41), .A2(n1046), .ZN(n1045) );
INV_X1 U753 ( .A(G131), .ZN(n1046) );
NAND3_X1 U754 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1044) );
NAND2_X1 U755 ( .A1(KEYINPUT16), .A2(n1050), .ZN(n1049) );
NAND3_X1 U756 ( .A1(G137), .A2(n1051), .A3(n1052), .ZN(n1048) );
NAND2_X1 U757 ( .A1(G134), .A2(n1053), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1054), .A2(n1051), .ZN(n1053) );
INV_X1 U759 ( .A(KEYINPUT16), .ZN(n1051) );
XOR2_X1 U760 ( .A(n1050), .B(KEYINPUT49), .Z(n1054) );
NOR2_X1 U761 ( .A1(G900), .A2(n986), .ZN(n1036) );
NOR2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1034) );
INV_X1 U763 ( .A(n1057), .ZN(n1056) );
AND2_X1 U764 ( .A1(G227), .A2(G900), .ZN(n1055) );
NOR3_X1 U765 ( .A1(n1058), .A2(KEYINPUT8), .A3(G953), .ZN(n1032) );
INV_X1 U766 ( .A(n982), .ZN(n1058) );
XOR2_X1 U767 ( .A(n1059), .B(n1060), .Z(G69) );
NAND2_X1 U768 ( .A1(n1057), .A2(n1061), .ZN(n1060) );
NAND2_X1 U769 ( .A1(n1062), .A2(G898), .ZN(n1061) );
XNOR2_X1 U770 ( .A(G224), .B(KEYINPUT5), .ZN(n1062) );
XOR2_X1 U771 ( .A(n986), .B(KEYINPUT56), .Z(n1057) );
NAND3_X1 U772 ( .A1(n1063), .A2(n1064), .A3(KEYINPUT1), .ZN(n1059) );
NAND2_X1 U773 ( .A1(G953), .A2(n1065), .ZN(n1064) );
XNOR2_X1 U774 ( .A(n984), .B(n1066), .ZN(n1063) );
NOR2_X1 U775 ( .A1(n1067), .A2(n1068), .ZN(G66) );
XOR2_X1 U776 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR2_X1 U777 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U778 ( .A1(KEYINPUT6), .A2(n1073), .ZN(n1069) );
NOR2_X1 U779 ( .A1(n1067), .A2(n1074), .ZN(G63) );
NOR2_X1 U780 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XOR2_X1 U781 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U782 ( .A1(n1079), .A2(n1072), .ZN(n1078) );
INV_X1 U783 ( .A(G478), .ZN(n1079) );
NOR2_X1 U784 ( .A1(KEYINPUT61), .A2(n1080), .ZN(n1077) );
AND2_X1 U785 ( .A1(n1080), .A2(KEYINPUT61), .ZN(n1075) );
NOR2_X1 U786 ( .A1(n1067), .A2(n1081), .ZN(G60) );
NOR2_X1 U787 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U788 ( .A(KEYINPUT33), .B(n1084), .Z(n1083) );
AND2_X1 U789 ( .A1(n1027), .A2(n1085), .ZN(n1084) );
NOR2_X1 U790 ( .A1(n1085), .A2(n1027), .ZN(n1082) );
NOR2_X1 U791 ( .A1(n1072), .A2(n1026), .ZN(n1085) );
INV_X1 U792 ( .A(G475), .ZN(n1026) );
XNOR2_X1 U793 ( .A(G104), .B(n1086), .ZN(G6) );
NOR2_X1 U794 ( .A1(n1067), .A2(n1087), .ZN(G57) );
XOR2_X1 U795 ( .A(n1088), .B(n1089), .Z(n1087) );
XOR2_X1 U796 ( .A(n1040), .B(n1090), .Z(n1089) );
XOR2_X1 U797 ( .A(n1091), .B(n1092), .Z(n1088) );
XOR2_X1 U798 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U799 ( .A1(KEYINPUT9), .A2(n1095), .ZN(n1094) );
NOR2_X1 U800 ( .A1(n1096), .A2(n1072), .ZN(n1093) );
INV_X1 U801 ( .A(G472), .ZN(n1096) );
NOR2_X1 U802 ( .A1(n1067), .A2(n1097), .ZN(G54) );
NOR2_X1 U803 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U804 ( .A(n1100), .B(KEYINPUT45), .Z(n1099) );
NAND2_X1 U805 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U806 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
XNOR2_X1 U807 ( .A(n1103), .B(n1104), .ZN(n1102) );
XOR2_X1 U808 ( .A(n1105), .B(n1040), .Z(n1103) );
NAND2_X1 U809 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND3_X1 U810 ( .A1(G227), .A2(n986), .A3(n1108), .ZN(n1107) );
XOR2_X1 U811 ( .A(n1109), .B(KEYINPUT53), .Z(n1108) );
NOR2_X1 U812 ( .A1(n1072), .A2(n1110), .ZN(n1101) );
NOR2_X1 U813 ( .A1(n1067), .A2(n1111), .ZN(G51) );
XOR2_X1 U814 ( .A(n1112), .B(n1113), .Z(n1111) );
NOR4_X1 U815 ( .A1(KEYINPUT59), .A2(n1114), .A3(n1072), .A4(n1115), .ZN(n1113) );
XOR2_X1 U816 ( .A(KEYINPUT7), .B(G210), .Z(n1115) );
NAND2_X1 U817 ( .A1(n1116), .A2(n1117), .ZN(n1072) );
OR2_X1 U818 ( .A1(n982), .A2(n984), .ZN(n1117) );
NAND2_X1 U819 ( .A1(n1118), .A2(n1119), .ZN(n984) );
AND4_X1 U820 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1119) );
AND4_X1 U821 ( .A1(n1124), .A2(n1125), .A3(n1086), .A4(n1126), .ZN(n1118) );
OR2_X1 U822 ( .A1(n978), .A2(n1003), .ZN(n1126) );
NAND4_X1 U823 ( .A1(n1127), .A2(n1011), .A3(n992), .A4(n1128), .ZN(n978) );
NAND3_X1 U824 ( .A1(n1129), .A2(n992), .A3(n1130), .ZN(n1086) );
NAND4_X1 U825 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n982) );
NOR4_X1 U826 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1134) );
INV_X1 U827 ( .A(n1139), .ZN(n1138) );
NOR2_X1 U828 ( .A1(n1140), .A2(n1141), .ZN(n1133) );
NOR3_X1 U829 ( .A1(n1142), .A2(n1000), .A3(n1003), .ZN(n1141) );
NOR2_X1 U830 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
XOR2_X1 U831 ( .A(n1145), .B(KEYINPUT55), .Z(n1143) );
NAND2_X1 U832 ( .A1(n1146), .A2(n1129), .ZN(n1145) );
XOR2_X1 U833 ( .A(KEYINPUT54), .B(G902), .Z(n1116) );
NAND3_X1 U834 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1112) );
NAND2_X1 U835 ( .A1(KEYINPUT37), .A2(n1150), .ZN(n1149) );
OR3_X1 U836 ( .A1(n1151), .A2(KEYINPUT37), .A3(n1066), .ZN(n1148) );
NAND2_X1 U837 ( .A1(n1066), .A2(n1151), .ZN(n1147) );
NAND2_X1 U838 ( .A1(KEYINPUT19), .A2(n1152), .ZN(n1151) );
INV_X1 U839 ( .A(n1150), .ZN(n1152) );
XOR2_X1 U840 ( .A(n1153), .B(n1040), .Z(n1150) );
XOR2_X1 U841 ( .A(n1154), .B(n1155), .Z(n1153) );
NOR2_X1 U842 ( .A1(KEYINPUT28), .A2(n1156), .ZN(n1155) );
NOR2_X1 U843 ( .A1(n986), .A2(G952), .ZN(n1067) );
XOR2_X1 U844 ( .A(G146), .B(n1137), .Z(G48) );
NOR3_X1 U845 ( .A1(n1142), .A2(n1003), .A3(n999), .ZN(n1137) );
XNOR2_X1 U846 ( .A(G143), .B(n1131), .ZN(G45) );
NAND4_X1 U847 ( .A1(n1146), .A2(n977), .A3(n1028), .A4(n1157), .ZN(n1131) );
XOR2_X1 U848 ( .A(G140), .B(n1136), .Z(G42) );
AND4_X1 U849 ( .A1(n1129), .A2(n1017), .A3(n997), .A4(n1158), .ZN(n1136) );
XOR2_X1 U850 ( .A(G137), .B(n1135), .Z(G39) );
NOR3_X1 U851 ( .A1(n1144), .A2(n1142), .A3(n1159), .ZN(n1135) );
INV_X1 U852 ( .A(n1001), .ZN(n1159) );
XOR2_X1 U853 ( .A(n1052), .B(n1132), .Z(G36) );
NAND3_X1 U854 ( .A1(n997), .A2(n1127), .A3(n1146), .ZN(n1132) );
AND2_X1 U855 ( .A1(n1016), .A2(n1158), .ZN(n1146) );
NAND2_X1 U856 ( .A1(n1160), .A2(n1161), .ZN(G33) );
NAND2_X1 U857 ( .A1(G131), .A2(n1162), .ZN(n1161) );
XOR2_X1 U858 ( .A(KEYINPUT44), .B(n1163), .Z(n1160) );
NOR2_X1 U859 ( .A1(G131), .A2(n1162), .ZN(n1163) );
NAND4_X1 U860 ( .A1(n1164), .A2(n1129), .A3(n997), .A4(n1158), .ZN(n1162) );
INV_X1 U861 ( .A(n1144), .ZN(n997) );
NAND2_X1 U862 ( .A1(n1165), .A2(n1006), .ZN(n1144) );
XOR2_X1 U863 ( .A(n1031), .B(KEYINPUT24), .Z(n1006) );
XNOR2_X1 U864 ( .A(n1016), .B(KEYINPUT23), .ZN(n1164) );
XOR2_X1 U865 ( .A(G128), .B(n1166), .Z(G30) );
NOR3_X1 U866 ( .A1(n1167), .A2(n1000), .A3(n1142), .ZN(n1166) );
NAND3_X1 U867 ( .A1(n1168), .A2(n1169), .A3(n1158), .ZN(n1142) );
AND2_X1 U868 ( .A1(n1011), .A2(n1170), .ZN(n1158) );
INV_X1 U869 ( .A(n1127), .ZN(n1000) );
XOR2_X1 U870 ( .A(KEYINPUT47), .B(n977), .Z(n1167) );
XOR2_X1 U871 ( .A(n1171), .B(n1172), .Z(G3) );
NAND2_X1 U872 ( .A1(KEYINPUT35), .A2(n1173), .ZN(n1172) );
INV_X1 U873 ( .A(n1122), .ZN(n1173) );
NAND3_X1 U874 ( .A1(n1016), .A2(n1001), .A3(n1130), .ZN(n1122) );
XOR2_X1 U875 ( .A(n1154), .B(n1139), .Z(G27) );
NAND3_X1 U876 ( .A1(n1129), .A2(n1017), .A3(n1174), .ZN(n1139) );
AND3_X1 U877 ( .A1(n994), .A2(n1170), .A3(n977), .ZN(n1174) );
NAND2_X1 U878 ( .A1(n1018), .A2(n1175), .ZN(n1170) );
NAND4_X1 U879 ( .A1(G953), .A2(G902), .A3(n1176), .A4(n1177), .ZN(n1175) );
INV_X1 U880 ( .A(G900), .ZN(n1177) );
NAND2_X1 U881 ( .A1(n1178), .A2(n1179), .ZN(G24) );
OR2_X1 U882 ( .A1(n1121), .A2(G122), .ZN(n1179) );
XOR2_X1 U883 ( .A(n1180), .B(KEYINPUT26), .Z(n1178) );
NAND2_X1 U884 ( .A1(G122), .A2(n1121), .ZN(n1180) );
NAND4_X1 U885 ( .A1(n1181), .A2(n992), .A3(n1028), .A4(n1157), .ZN(n1121) );
AND2_X1 U886 ( .A1(n1182), .A2(n1183), .ZN(n992) );
XOR2_X1 U887 ( .A(n1168), .B(KEYINPUT3), .Z(n1182) );
XNOR2_X1 U888 ( .A(G119), .B(n1120), .ZN(G21) );
NAND4_X1 U889 ( .A1(n1181), .A2(n1001), .A3(n1168), .A4(n1169), .ZN(n1120) );
XOR2_X1 U890 ( .A(n1184), .B(n1125), .Z(G18) );
NAND3_X1 U891 ( .A1(n1016), .A2(n1127), .A3(n1181), .ZN(n1125) );
NOR2_X1 U892 ( .A1(n1185), .A2(n1186), .ZN(n1127) );
XNOR2_X1 U893 ( .A(G113), .B(n1124), .ZN(G15) );
NAND3_X1 U894 ( .A1(n1016), .A2(n1129), .A3(n1181), .ZN(n1124) );
AND3_X1 U895 ( .A1(n977), .A2(n1128), .A3(n994), .ZN(n1181) );
INV_X1 U896 ( .A(n1030), .ZN(n994) );
NAND2_X1 U897 ( .A1(n1012), .A2(n1187), .ZN(n1030) );
INV_X1 U898 ( .A(n999), .ZN(n1129) );
NAND2_X1 U899 ( .A1(n1157), .A2(n1186), .ZN(n999) );
INV_X1 U900 ( .A(n1028), .ZN(n1186) );
XNOR2_X1 U901 ( .A(n1185), .B(KEYINPUT10), .ZN(n1157) );
AND2_X1 U902 ( .A1(n1183), .A2(n1168), .ZN(n1016) );
XNOR2_X1 U903 ( .A(G110), .B(n1123), .ZN(G12) );
NAND3_X1 U904 ( .A1(n1017), .A2(n1001), .A3(n1130), .ZN(n1123) );
AND3_X1 U905 ( .A1(n1011), .A2(n1128), .A3(n977), .ZN(n1130) );
INV_X1 U906 ( .A(n1003), .ZN(n977) );
NAND2_X1 U907 ( .A1(n1165), .A2(n1031), .ZN(n1003) );
XNOR2_X1 U908 ( .A(n1188), .B(n1189), .ZN(n1031) );
NOR2_X1 U909 ( .A1(n1114), .A2(n1190), .ZN(n1189) );
INV_X1 U910 ( .A(G210), .ZN(n1190) );
NAND2_X1 U911 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
XOR2_X1 U912 ( .A(n1193), .B(n1194), .Z(n1191) );
XOR2_X1 U913 ( .A(n1156), .B(n1195), .Z(n1194) );
XNOR2_X1 U914 ( .A(KEYINPUT52), .B(KEYINPUT0), .ZN(n1195) );
NAND2_X1 U915 ( .A1(G224), .A2(n986), .ZN(n1156) );
XNOR2_X1 U916 ( .A(n1066), .B(n1196), .ZN(n1193) );
XOR2_X1 U917 ( .A(n1197), .B(n1040), .Z(n1196) );
NOR2_X1 U918 ( .A1(KEYINPUT63), .A2(n1154), .ZN(n1197) );
INV_X1 U919 ( .A(G125), .ZN(n1154) );
XNOR2_X1 U920 ( .A(n1198), .B(n1199), .ZN(n1066) );
XOR2_X1 U921 ( .A(G101), .B(n1200), .Z(n1199) );
XOR2_X1 U922 ( .A(G113), .B(G110), .Z(n1200) );
XOR2_X1 U923 ( .A(n1201), .B(n1202), .Z(n1198) );
XOR2_X1 U924 ( .A(n1203), .B(n1204), .Z(n1201) );
NOR2_X1 U925 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U926 ( .A(KEYINPUT36), .B(KEYINPUT17), .Z(n1206) );
NAND2_X1 U927 ( .A1(KEYINPUT2), .A2(n1207), .ZN(n1203) );
XOR2_X1 U928 ( .A(KEYINPUT22), .B(n1005), .Z(n1165) );
NOR2_X1 U929 ( .A1(n1208), .A2(n1114), .ZN(n1005) );
NOR2_X1 U930 ( .A1(G902), .A2(G237), .ZN(n1114) );
INV_X1 U931 ( .A(G214), .ZN(n1208) );
NAND2_X1 U932 ( .A1(n1018), .A2(n1209), .ZN(n1128) );
NAND4_X1 U933 ( .A1(G953), .A2(G902), .A3(n1176), .A4(n1065), .ZN(n1209) );
INV_X1 U934 ( .A(G898), .ZN(n1065) );
NAND3_X1 U935 ( .A1(n1176), .A2(n986), .A3(G952), .ZN(n1018) );
NAND2_X1 U936 ( .A1(G237), .A2(G234), .ZN(n1176) );
NOR2_X1 U937 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
INV_X1 U938 ( .A(n1187), .ZN(n1013) );
NAND2_X1 U939 ( .A1(G221), .A2(n1210), .ZN(n1187) );
XNOR2_X1 U940 ( .A(n1211), .B(n1110), .ZN(n1012) );
INV_X1 U941 ( .A(G469), .ZN(n1110) );
NAND2_X1 U942 ( .A1(n1192), .A2(n1212), .ZN(n1211) );
NAND2_X1 U943 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND3_X1 U944 ( .A1(n1215), .A2(n1106), .A3(n1216), .ZN(n1214) );
XNOR2_X1 U945 ( .A(n1217), .B(n1104), .ZN(n1216) );
XOR2_X1 U946 ( .A(n1218), .B(KEYINPUT34), .Z(n1213) );
NAND2_X1 U947 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND2_X1 U948 ( .A1(n1215), .A2(n1106), .ZN(n1220) );
NAND2_X1 U949 ( .A1(n1221), .A2(n1222), .ZN(n1106) );
NAND2_X1 U950 ( .A1(G227), .A2(n986), .ZN(n1222) );
NAND2_X1 U951 ( .A1(n1109), .A2(G227), .ZN(n1215) );
INV_X1 U952 ( .A(n1221), .ZN(n1109) );
XOR2_X1 U953 ( .A(G140), .B(G110), .Z(n1221) );
XOR2_X1 U954 ( .A(n1217), .B(n1104), .Z(n1219) );
XOR2_X1 U955 ( .A(n1207), .B(n1090), .Z(n1104) );
XOR2_X1 U956 ( .A(G101), .B(n1223), .Z(n1090) );
XOR2_X1 U957 ( .A(G104), .B(n1224), .Z(n1207) );
NOR2_X1 U958 ( .A1(KEYINPUT58), .A2(n1040), .ZN(n1217) );
NOR2_X1 U959 ( .A1(n1185), .A2(n1028), .ZN(n1001) );
XOR2_X1 U960 ( .A(n1225), .B(n1226), .Z(n1028) );
XOR2_X1 U961 ( .A(KEYINPUT14), .B(G478), .Z(n1226) );
NAND2_X1 U962 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
INV_X1 U963 ( .A(n1080), .ZN(n1228) );
XOR2_X1 U964 ( .A(n1229), .B(n1230), .Z(n1080) );
XOR2_X1 U965 ( .A(n1224), .B(n1202), .Z(n1230) );
XOR2_X1 U966 ( .A(G107), .B(KEYINPUT25), .Z(n1224) );
XOR2_X1 U967 ( .A(n1231), .B(n1232), .Z(n1229) );
NOR2_X1 U968 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
INV_X1 U969 ( .A(G217), .ZN(n1234) );
XNOR2_X1 U970 ( .A(n1235), .B(n1236), .ZN(n1231) );
NAND2_X1 U971 ( .A1(KEYINPUT18), .A2(n1184), .ZN(n1236) );
NAND2_X1 U972 ( .A1(KEYINPUT42), .A2(n1237), .ZN(n1235) );
XNOR2_X1 U973 ( .A(n1238), .B(n1239), .ZN(n1237) );
NAND2_X1 U974 ( .A1(KEYINPUT50), .A2(n1052), .ZN(n1238) );
INV_X1 U975 ( .A(G134), .ZN(n1052) );
XOR2_X1 U976 ( .A(n1192), .B(KEYINPUT60), .Z(n1227) );
NAND2_X1 U977 ( .A1(n1240), .A2(n1241), .ZN(n1185) );
NAND2_X1 U978 ( .A1(G475), .A2(n1242), .ZN(n1241) );
NAND3_X1 U979 ( .A1(n1243), .A2(n1192), .A3(KEYINPUT38), .ZN(n1242) );
NAND2_X1 U980 ( .A1(n1022), .A2(KEYINPUT38), .ZN(n1240) );
NOR3_X1 U981 ( .A1(G475), .A2(G902), .A3(n1027), .ZN(n1022) );
INV_X1 U982 ( .A(n1243), .ZN(n1027) );
XOR2_X1 U983 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U984 ( .A(n1246), .B(n1247), .Z(n1245) );
XOR2_X1 U985 ( .A(G113), .B(G104), .Z(n1247) );
XOR2_X1 U986 ( .A(G143), .B(G131), .Z(n1246) );
XOR2_X1 U987 ( .A(n1248), .B(n1249), .Z(n1244) );
XOR2_X1 U988 ( .A(n1041), .B(n1202), .Z(n1249) );
XOR2_X1 U989 ( .A(G122), .B(KEYINPUT15), .Z(n1202) );
XNOR2_X1 U990 ( .A(n1250), .B(n1251), .ZN(n1248) );
NAND2_X1 U991 ( .A1(n1252), .A2(G214), .ZN(n1250) );
NOR2_X1 U992 ( .A1(n1253), .A2(n1168), .ZN(n1017) );
XOR2_X1 U993 ( .A(n1024), .B(KEYINPUT12), .Z(n1168) );
XOR2_X1 U994 ( .A(n1254), .B(n1255), .Z(n1024) );
XOR2_X1 U995 ( .A(KEYINPUT57), .B(G472), .Z(n1255) );
NAND2_X1 U996 ( .A1(n1256), .A2(n1192), .ZN(n1254) );
XNOR2_X1 U997 ( .A(n1095), .B(n1257), .ZN(n1256) );
XOR2_X1 U998 ( .A(n1171), .B(n1258), .Z(n1257) );
NAND2_X1 U999 ( .A1(n1259), .A2(KEYINPUT29), .ZN(n1258) );
XOR2_X1 U1000 ( .A(n1260), .B(n1223), .Z(n1259) );
XNOR2_X1 U1001 ( .A(n1261), .B(n1262), .ZN(n1223) );
XOR2_X1 U1002 ( .A(G137), .B(n1263), .Z(n1262) );
NOR2_X1 U1003 ( .A1(G134), .A2(KEYINPUT46), .ZN(n1263) );
NAND2_X1 U1004 ( .A1(KEYINPUT43), .A2(G131), .ZN(n1261) );
XOR2_X1 U1005 ( .A(n1264), .B(n1091), .Z(n1260) );
XNOR2_X1 U1006 ( .A(n1265), .B(n1266), .ZN(n1091) );
XOR2_X1 U1007 ( .A(KEYINPUT27), .B(KEYINPUT13), .Z(n1266) );
XOR2_X1 U1008 ( .A(G113), .B(n1205), .Z(n1265) );
XOR2_X1 U1009 ( .A(n1184), .B(G119), .Z(n1205) );
INV_X1 U1010 ( .A(G116), .ZN(n1184) );
NAND2_X1 U1011 ( .A1(KEYINPUT20), .A2(n1040), .ZN(n1264) );
XNOR2_X1 U1012 ( .A(n1251), .B(n1239), .ZN(n1040) );
XOR2_X1 U1013 ( .A(G128), .B(G143), .Z(n1239) );
INV_X1 U1014 ( .A(G101), .ZN(n1171) );
NAND2_X1 U1015 ( .A1(n1252), .A2(G210), .ZN(n1095) );
NOR2_X1 U1016 ( .A1(G953), .A2(G237), .ZN(n1252) );
INV_X1 U1017 ( .A(n1169), .ZN(n1253) );
XOR2_X1 U1018 ( .A(n1029), .B(KEYINPUT51), .Z(n1169) );
INV_X1 U1019 ( .A(n1183), .ZN(n1029) );
XNOR2_X1 U1020 ( .A(n1267), .B(n1071), .ZN(n1183) );
NAND2_X1 U1021 ( .A1(G217), .A2(n1210), .ZN(n1071) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1192), .ZN(n1210) );
NAND2_X1 U1023 ( .A1(n1073), .A2(n1192), .ZN(n1267) );
INV_X1 U1024 ( .A(G902), .ZN(n1192) );
XOR2_X1 U1025 ( .A(n1268), .B(n1269), .Z(n1073) );
XOR2_X1 U1026 ( .A(n1270), .B(n1271), .Z(n1269) );
INV_X1 U1027 ( .A(n1041), .ZN(n1271) );
XOR2_X1 U1028 ( .A(G140), .B(G125), .Z(n1041) );
NAND2_X1 U1029 ( .A1(n1272), .A2(KEYINPUT40), .ZN(n1270) );
XOR2_X1 U1030 ( .A(n1273), .B(n1274), .Z(n1272) );
XOR2_X1 U1031 ( .A(KEYINPUT30), .B(G128), .Z(n1274) );
XNOR2_X1 U1032 ( .A(G119), .B(G110), .ZN(n1273) );
XOR2_X1 U1033 ( .A(n1275), .B(n1276), .Z(n1268) );
NOR2_X1 U1034 ( .A1(n1233), .A2(n1277), .ZN(n1276) );
INV_X1 U1035 ( .A(G221), .ZN(n1277) );
NAND2_X1 U1036 ( .A1(G234), .A2(n986), .ZN(n1233) );
INV_X1 U1037 ( .A(G953), .ZN(n986) );
XOR2_X1 U1038 ( .A(n1050), .B(n1278), .Z(n1275) );
NOR2_X1 U1039 ( .A1(KEYINPUT32), .A2(n1251), .ZN(n1278) );
XNOR2_X1 U1040 ( .A(G146), .B(KEYINPUT62), .ZN(n1251) );
INV_X1 U1041 ( .A(G137), .ZN(n1050) );
endmodule


