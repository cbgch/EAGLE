//Key = 1010111000010101101110011001000110010001100011000111111110011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296;

XNOR2_X1 U735 ( .A(n998), .B(n999), .ZN(G9) );
NOR2_X1 U736 ( .A1(KEYINPUT8), .A2(n1000), .ZN(n999) );
INV_X1 U737 ( .A(G107), .ZN(n1000) );
NAND3_X1 U738 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(G75) );
NAND2_X1 U739 ( .A1(G952), .A2(n1004), .ZN(n1003) );
NAND3_X1 U740 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
NAND2_X1 U741 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NAND2_X1 U742 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND4_X1 U743 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
NOR2_X1 U744 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U745 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
OR2_X1 U746 ( .A1(n1020), .A2(n1021), .ZN(n1013) );
OR3_X1 U747 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1012) );
NAND4_X1 U748 ( .A1(n1025), .A2(n1020), .A3(n1021), .A4(n1026), .ZN(n1010) );
NAND2_X1 U749 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XOR2_X1 U750 ( .A(KEYINPUT28), .B(n1029), .Z(n1028) );
NOR2_X1 U751 ( .A1(n1030), .A2(n1031), .ZN(n1025) );
NOR3_X1 U752 ( .A1(n1017), .A2(n1032), .A3(n1033), .ZN(n1031) );
INV_X1 U753 ( .A(n1034), .ZN(n1017) );
NOR2_X1 U754 ( .A1(n1034), .A2(n1014), .ZN(n1030) );
INV_X1 U755 ( .A(n1035), .ZN(n1008) );
NAND2_X1 U756 ( .A1(KEYINPUT7), .A2(n1036), .ZN(n1005) );
NAND2_X1 U757 ( .A1(n1037), .A2(n1038), .ZN(n1001) );
NAND2_X1 U758 ( .A1(KEYINPUT7), .A2(G952), .ZN(n1038) );
INV_X1 U759 ( .A(n1036), .ZN(n1037) );
NAND4_X1 U760 ( .A1(n1034), .A2(n1020), .A3(n1039), .A4(n1040), .ZN(n1036) );
NOR3_X1 U761 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
XNOR2_X1 U762 ( .A(n1044), .B(n1045), .ZN(n1039) );
XOR2_X1 U763 ( .A(n1046), .B(n1047), .Z(G72) );
NOR3_X1 U764 ( .A1(n1048), .A2(KEYINPUT47), .A3(n1049), .ZN(n1047) );
NOR2_X1 U765 ( .A1(G900), .A2(n1050), .ZN(n1049) );
XNOR2_X1 U766 ( .A(G953), .B(KEYINPUT14), .ZN(n1050) );
XOR2_X1 U767 ( .A(n1051), .B(n1052), .Z(n1048) );
XOR2_X1 U768 ( .A(n1053), .B(n1054), .Z(n1052) );
XOR2_X1 U769 ( .A(n1055), .B(n1056), .Z(n1051) );
XOR2_X1 U770 ( .A(KEYINPUT4), .B(KEYINPUT16), .Z(n1056) );
NAND2_X1 U771 ( .A1(n1057), .A2(n1058), .ZN(n1046) );
NAND2_X1 U772 ( .A1(n1059), .A2(n1002), .ZN(n1058) );
NAND2_X1 U773 ( .A1(G953), .A2(n1060), .ZN(n1057) );
NAND2_X1 U774 ( .A1(G227), .A2(n1061), .ZN(n1060) );
XNOR2_X1 U775 ( .A(KEYINPUT38), .B(n1062), .ZN(n1061) );
XOR2_X1 U776 ( .A(n1063), .B(n1064), .Z(G69) );
XOR2_X1 U777 ( .A(n1065), .B(n1066), .Z(n1064) );
OR2_X1 U778 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U779 ( .A1(n1069), .A2(n1002), .ZN(n1065) );
NOR3_X1 U780 ( .A1(n1002), .A2(KEYINPUT34), .A3(n1070), .ZN(n1063) );
AND2_X1 U781 ( .A1(G224), .A2(G898), .ZN(n1070) );
NOR2_X1 U782 ( .A1(n1071), .A2(n1072), .ZN(G66) );
XOR2_X1 U783 ( .A(n1073), .B(n1074), .Z(n1072) );
NAND2_X1 U784 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR2_X1 U785 ( .A1(n1071), .A2(n1077), .ZN(G63) );
XOR2_X1 U786 ( .A(n1078), .B(n1079), .Z(n1077) );
NAND2_X1 U787 ( .A1(n1075), .A2(G478), .ZN(n1079) );
NOR2_X1 U788 ( .A1(n1080), .A2(n1081), .ZN(G60) );
XOR2_X1 U789 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U790 ( .A1(KEYINPUT25), .A2(n1084), .ZN(n1083) );
NOR3_X1 U791 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1082) );
NOR2_X1 U792 ( .A1(KEYINPUT27), .A2(n1088), .ZN(n1087) );
AND2_X1 U793 ( .A1(G902), .A2(n1007), .ZN(n1088) );
NOR2_X1 U794 ( .A1(n1075), .A2(n1089), .ZN(n1086) );
INV_X1 U795 ( .A(KEYINPUT27), .ZN(n1089) );
NOR2_X1 U796 ( .A1(n1090), .A2(n1091), .ZN(n1080) );
XOR2_X1 U797 ( .A(KEYINPUT58), .B(n1092), .Z(n1090) );
XNOR2_X1 U798 ( .A(G104), .B(n1093), .ZN(G6) );
NOR2_X1 U799 ( .A1(n1071), .A2(n1094), .ZN(G57) );
XOR2_X1 U800 ( .A(n1095), .B(n1096), .Z(n1094) );
XOR2_X1 U801 ( .A(n1097), .B(n1098), .Z(n1096) );
XNOR2_X1 U802 ( .A(KEYINPUT35), .B(KEYINPUT29), .ZN(n1098) );
XOR2_X1 U803 ( .A(n1099), .B(n1100), .Z(n1095) );
XOR2_X1 U804 ( .A(n1101), .B(n1102), .Z(n1099) );
NAND2_X1 U805 ( .A1(n1075), .A2(G472), .ZN(n1101) );
NOR2_X1 U806 ( .A1(n1071), .A2(n1103), .ZN(G54) );
XOR2_X1 U807 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U808 ( .A1(KEYINPUT43), .A2(n1106), .ZN(n1105) );
XOR2_X1 U809 ( .A(n1107), .B(n1108), .Z(n1106) );
XNOR2_X1 U810 ( .A(n1109), .B(n1110), .ZN(n1108) );
XNOR2_X1 U811 ( .A(n1111), .B(n1112), .ZN(n1107) );
XNOR2_X1 U812 ( .A(G140), .B(n1113), .ZN(n1112) );
NAND2_X1 U813 ( .A1(n1075), .A2(G469), .ZN(n1104) );
NOR2_X1 U814 ( .A1(n1071), .A2(n1114), .ZN(G51) );
XOR2_X1 U815 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U816 ( .A1(n1075), .A2(n1117), .ZN(n1116) );
NOR2_X1 U817 ( .A1(n1118), .A2(n1007), .ZN(n1075) );
NOR2_X1 U818 ( .A1(n1069), .A2(n1059), .ZN(n1007) );
NAND2_X1 U819 ( .A1(n1119), .A2(n1120), .ZN(n1059) );
AND4_X1 U820 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
NOR4_X1 U821 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1119) );
NOR3_X1 U822 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
INV_X1 U823 ( .A(n1132), .ZN(n1127) );
NAND4_X1 U824 ( .A1(n1133), .A2(n1093), .A3(n1134), .A4(n1135), .ZN(n1069) );
NOR4_X1 U825 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1135) );
NOR3_X1 U826 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1134) );
NOR2_X1 U827 ( .A1(n1143), .A2(n998), .ZN(n1142) );
NAND3_X1 U828 ( .A1(n1033), .A2(n1144), .A3(n1021), .ZN(n998) );
INV_X1 U829 ( .A(KEYINPUT13), .ZN(n1143) );
NOR4_X1 U830 ( .A1(KEYINPUT13), .A2(n1145), .A3(n1146), .A4(n1130), .ZN(n1141) );
NAND2_X1 U831 ( .A1(n1147), .A2(n1021), .ZN(n1145) );
NOR2_X1 U832 ( .A1(n1147), .A2(n1148), .ZN(n1140) );
NAND3_X1 U833 ( .A1(n1021), .A2(n1144), .A3(n1032), .ZN(n1093) );
NAND2_X1 U834 ( .A1(n1149), .A2(n1150), .ZN(n1133) );
XNOR2_X1 U835 ( .A(KEYINPUT26), .B(n1131), .ZN(n1150) );
NAND2_X1 U836 ( .A1(n1151), .A2(KEYINPUT49), .ZN(n1115) );
XOR2_X1 U837 ( .A(n1067), .B(n1152), .Z(n1151) );
NOR2_X1 U838 ( .A1(KEYINPUT37), .A2(n1153), .ZN(n1152) );
XOR2_X1 U839 ( .A(n1154), .B(n1155), .Z(n1153) );
XNOR2_X1 U840 ( .A(n1156), .B(n1157), .ZN(n1155) );
NOR2_X1 U841 ( .A1(G125), .A2(KEYINPUT46), .ZN(n1157) );
NOR2_X1 U842 ( .A1(n1091), .A2(n1092), .ZN(n1071) );
XOR2_X1 U843 ( .A(G952), .B(KEYINPUT10), .Z(n1092) );
XNOR2_X1 U844 ( .A(KEYINPUT19), .B(n1002), .ZN(n1091) );
XNOR2_X1 U845 ( .A(G146), .B(n1124), .ZN(G48) );
NAND2_X1 U846 ( .A1(n1158), .A2(n1032), .ZN(n1124) );
XNOR2_X1 U847 ( .A(n1159), .B(n1160), .ZN(G45) );
NOR2_X1 U848 ( .A1(KEYINPUT41), .A2(n1132), .ZN(n1160) );
NAND4_X1 U849 ( .A1(n1042), .A2(n1161), .A3(n1041), .A4(n1162), .ZN(n1132) );
NOR2_X1 U850 ( .A1(n1146), .A2(n1131), .ZN(n1162) );
XOR2_X1 U851 ( .A(G140), .B(n1126), .Z(G42) );
AND3_X1 U852 ( .A1(n1032), .A2(n1022), .A3(n1163), .ZN(n1126) );
XOR2_X1 U853 ( .A(G137), .B(n1125), .Z(G39) );
AND2_X1 U854 ( .A1(n1163), .A2(n1164), .ZN(n1125) );
XNOR2_X1 U855 ( .A(G134), .B(n1165), .ZN(G36) );
NAND4_X1 U856 ( .A1(KEYINPUT20), .A2(n1163), .A3(n1023), .A4(n1033), .ZN(n1165) );
XNOR2_X1 U857 ( .A(G131), .B(n1123), .ZN(G33) );
NAND3_X1 U858 ( .A1(n1032), .A2(n1023), .A3(n1163), .ZN(n1123) );
INV_X1 U859 ( .A(n1129), .ZN(n1163) );
NAND4_X1 U860 ( .A1(n1020), .A2(n1029), .A3(n1161), .A4(n1166), .ZN(n1129) );
INV_X1 U861 ( .A(n1024), .ZN(n1020) );
NAND2_X1 U862 ( .A1(n1018), .A2(n1019), .ZN(n1024) );
INV_X1 U863 ( .A(n1167), .ZN(n1018) );
XNOR2_X1 U864 ( .A(G128), .B(n1122), .ZN(G30) );
NAND2_X1 U865 ( .A1(n1158), .A2(n1033), .ZN(n1122) );
NOR4_X1 U866 ( .A1(n1168), .A2(n1146), .A3(n1169), .A4(n1170), .ZN(n1158) );
INV_X1 U867 ( .A(n1161), .ZN(n1170) );
XOR2_X1 U868 ( .A(G101), .B(n1171), .Z(G3) );
NOR2_X1 U869 ( .A1(n1172), .A2(n1131), .ZN(n1171) );
INV_X1 U870 ( .A(n1023), .ZN(n1131) );
XNOR2_X1 U871 ( .A(G125), .B(n1121), .ZN(G27) );
NAND4_X1 U872 ( .A1(n1032), .A2(n1173), .A3(n1022), .A4(n1161), .ZN(n1121) );
NAND2_X1 U873 ( .A1(n1035), .A2(n1174), .ZN(n1161) );
NAND4_X1 U874 ( .A1(G902), .A2(G953), .A3(n1175), .A4(n1062), .ZN(n1174) );
INV_X1 U875 ( .A(G900), .ZN(n1062) );
XOR2_X1 U876 ( .A(G122), .B(n1176), .Z(G24) );
NOR2_X1 U877 ( .A1(n1148), .A2(n1177), .ZN(n1176) );
XNOR2_X1 U878 ( .A(KEYINPUT17), .B(n1178), .ZN(n1177) );
NAND4_X1 U879 ( .A1(n1173), .A2(n1021), .A3(n1041), .A4(n1042), .ZN(n1148) );
NOR2_X1 U880 ( .A1(n1043), .A2(n1179), .ZN(n1021) );
XOR2_X1 U881 ( .A(G119), .B(n1139), .Z(G21) );
AND3_X1 U882 ( .A1(n1173), .A2(n1178), .A3(n1164), .ZN(n1139) );
AND3_X1 U883 ( .A1(n1014), .A2(n1043), .A3(n1179), .ZN(n1164) );
XOR2_X1 U884 ( .A(G116), .B(n1138), .Z(G18) );
AND2_X1 U885 ( .A1(n1180), .A2(n1033), .ZN(n1138) );
INV_X1 U886 ( .A(n1130), .ZN(n1033) );
NAND2_X1 U887 ( .A1(n1181), .A2(n1041), .ZN(n1130) );
XOR2_X1 U888 ( .A(G113), .B(n1137), .Z(G15) );
AND2_X1 U889 ( .A1(n1032), .A2(n1180), .ZN(n1137) );
AND3_X1 U890 ( .A1(n1173), .A2(n1178), .A3(n1023), .ZN(n1180) );
NOR2_X1 U891 ( .A1(n1168), .A2(n1043), .ZN(n1023) );
AND3_X1 U892 ( .A1(n1167), .A2(n1019), .A3(n1034), .ZN(n1173) );
NOR2_X1 U893 ( .A1(n1029), .A2(n1027), .ZN(n1034) );
INV_X1 U894 ( .A(n1166), .ZN(n1027) );
AND2_X1 U895 ( .A1(n1182), .A2(n1042), .ZN(n1032) );
XNOR2_X1 U896 ( .A(n1113), .B(n1136), .ZN(G12) );
AND2_X1 U897 ( .A1(n1149), .A2(n1022), .ZN(n1136) );
NOR2_X1 U898 ( .A1(n1169), .A2(n1179), .ZN(n1022) );
INV_X1 U899 ( .A(n1168), .ZN(n1179) );
NAND3_X1 U900 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1168) );
OR2_X1 U901 ( .A1(n1044), .A2(n1186), .ZN(n1185) );
NAND3_X1 U902 ( .A1(n1186), .A2(n1044), .A3(KEYINPUT32), .ZN(n1184) );
NAND2_X1 U903 ( .A1(n1187), .A2(n1118), .ZN(n1044) );
XOR2_X1 U904 ( .A(n1188), .B(n1189), .Z(n1187) );
XOR2_X1 U905 ( .A(n1097), .B(G101), .Z(n1189) );
NAND3_X1 U906 ( .A1(n1190), .A2(n1002), .A3(G210), .ZN(n1097) );
NAND2_X1 U907 ( .A1(KEYINPUT45), .A2(n1191), .ZN(n1188) );
XNOR2_X1 U908 ( .A(n1100), .B(n1192), .ZN(n1191) );
XNOR2_X1 U909 ( .A(n1193), .B(n1194), .ZN(n1100) );
XNOR2_X1 U910 ( .A(n1195), .B(KEYINPUT61), .ZN(n1194) );
NAND2_X1 U911 ( .A1(KEYINPUT0), .A2(n1196), .ZN(n1195) );
XOR2_X1 U912 ( .A(KEYINPUT3), .B(G116), .Z(n1196) );
XOR2_X1 U913 ( .A(n1154), .B(n1053), .Z(n1193) );
AND2_X1 U914 ( .A1(n1197), .A2(n1045), .ZN(n1186) );
XNOR2_X1 U915 ( .A(KEYINPUT60), .B(KEYINPUT51), .ZN(n1197) );
OR2_X1 U916 ( .A1(n1045), .A2(KEYINPUT32), .ZN(n1183) );
INV_X1 U917 ( .A(G472), .ZN(n1045) );
INV_X1 U918 ( .A(n1043), .ZN(n1169) );
XNOR2_X1 U919 ( .A(n1198), .B(n1076), .ZN(n1043) );
AND2_X1 U920 ( .A1(G217), .A2(n1199), .ZN(n1076) );
NAND2_X1 U921 ( .A1(n1074), .A2(n1118), .ZN(n1198) );
XNOR2_X1 U922 ( .A(n1200), .B(n1201), .ZN(n1074) );
XOR2_X1 U923 ( .A(n1202), .B(n1203), .Z(n1201) );
XNOR2_X1 U924 ( .A(n1204), .B(n1205), .ZN(n1203) );
NOR2_X1 U925 ( .A1(G146), .A2(KEYINPUT12), .ZN(n1205) );
NAND4_X1 U926 ( .A1(KEYINPUT2), .A2(G221), .A3(G234), .A4(n1002), .ZN(n1204) );
XOR2_X1 U927 ( .A(n1206), .B(n1207), .Z(n1200) );
XNOR2_X1 U928 ( .A(G137), .B(n1208), .ZN(n1207) );
XNOR2_X1 U929 ( .A(G119), .B(n1209), .ZN(n1206) );
NOR2_X1 U930 ( .A1(KEYINPUT33), .A2(n1113), .ZN(n1209) );
INV_X1 U931 ( .A(n1172), .ZN(n1149) );
NAND2_X1 U932 ( .A1(n1014), .A2(n1144), .ZN(n1172) );
NOR2_X1 U933 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
INV_X1 U934 ( .A(n1178), .ZN(n1147) );
NAND2_X1 U935 ( .A1(n1035), .A2(n1210), .ZN(n1178) );
NAND3_X1 U936 ( .A1(n1068), .A2(n1175), .A3(G902), .ZN(n1210) );
NOR2_X1 U937 ( .A1(n1002), .A2(G898), .ZN(n1068) );
NAND3_X1 U938 ( .A1(n1175), .A2(n1002), .A3(G952), .ZN(n1035) );
NAND2_X1 U939 ( .A1(G237), .A2(n1211), .ZN(n1175) );
NAND4_X1 U940 ( .A1(n1167), .A2(n1029), .A3(n1019), .A4(n1166), .ZN(n1146) );
NAND2_X1 U941 ( .A1(G221), .A2(n1199), .ZN(n1166) );
NAND2_X1 U942 ( .A1(n1211), .A2(n1118), .ZN(n1199) );
XNOR2_X1 U943 ( .A(G234), .B(KEYINPUT52), .ZN(n1211) );
NAND2_X1 U944 ( .A1(G214), .A2(n1212), .ZN(n1019) );
XNOR2_X1 U945 ( .A(n1213), .B(G469), .ZN(n1029) );
NAND2_X1 U946 ( .A1(n1214), .A2(n1118), .ZN(n1213) );
XOR2_X1 U947 ( .A(n1215), .B(n1216), .Z(n1214) );
XOR2_X1 U948 ( .A(n1217), .B(n1110), .Z(n1216) );
XNOR2_X1 U949 ( .A(n1218), .B(n1053), .ZN(n1110) );
XNOR2_X1 U950 ( .A(n1219), .B(n1220), .ZN(n1053) );
XNOR2_X1 U951 ( .A(G131), .B(G137), .ZN(n1219) );
NAND2_X1 U952 ( .A1(G227), .A2(n1002), .ZN(n1218) );
NOR2_X1 U953 ( .A1(G110), .A2(KEYINPUT22), .ZN(n1217) );
XOR2_X1 U954 ( .A(n1221), .B(n1222), .Z(n1215) );
XOR2_X1 U955 ( .A(KEYINPUT48), .B(G140), .Z(n1222) );
NOR2_X1 U956 ( .A1(KEYINPUT30), .A2(n1223), .ZN(n1221) );
XNOR2_X1 U957 ( .A(n1224), .B(n1225), .ZN(n1223) );
INV_X1 U958 ( .A(n1111), .ZN(n1225) );
XNOR2_X1 U959 ( .A(n1226), .B(n1227), .ZN(n1111) );
NOR2_X1 U960 ( .A1(G101), .A2(KEYINPUT1), .ZN(n1227) );
NAND3_X1 U961 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(n1226) );
NAND2_X1 U962 ( .A1(G104), .A2(n1231), .ZN(n1230) );
NAND2_X1 U963 ( .A1(KEYINPUT63), .A2(n1232), .ZN(n1229) );
NAND2_X1 U964 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XNOR2_X1 U965 ( .A(KEYINPUT44), .B(n1235), .ZN(n1233) );
NAND2_X1 U966 ( .A1(n1236), .A2(n1237), .ZN(n1228) );
INV_X1 U967 ( .A(KEYINPUT63), .ZN(n1237) );
NAND2_X1 U968 ( .A1(n1238), .A2(n1239), .ZN(n1236) );
NAND3_X1 U969 ( .A1(KEYINPUT44), .A2(n1234), .A3(n1235), .ZN(n1239) );
INV_X1 U970 ( .A(G104), .ZN(n1234) );
OR2_X1 U971 ( .A1(n1235), .A2(KEYINPUT44), .ZN(n1238) );
NAND2_X1 U972 ( .A1(KEYINPUT55), .A2(n1109), .ZN(n1224) );
XOR2_X1 U973 ( .A(n1055), .B(KEYINPUT6), .Z(n1109) );
XNOR2_X1 U974 ( .A(G128), .B(n1240), .ZN(n1055) );
XNOR2_X1 U975 ( .A(n1241), .B(n1117), .ZN(n1167) );
AND2_X1 U976 ( .A1(G210), .A2(n1212), .ZN(n1117) );
NAND2_X1 U977 ( .A1(n1190), .A2(n1118), .ZN(n1212) );
NAND2_X1 U978 ( .A1(n1242), .A2(n1118), .ZN(n1241) );
XOR2_X1 U979 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U980 ( .A(n1067), .B(n1154), .Z(n1244) );
NAND2_X1 U981 ( .A1(n1245), .A2(n1246), .ZN(n1154) );
NAND2_X1 U982 ( .A1(G128), .A2(n1247), .ZN(n1246) );
NAND2_X1 U983 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U984 ( .A1(G143), .A2(n1250), .ZN(n1249) );
XOR2_X1 U985 ( .A(KEYINPUT39), .B(n1251), .Z(n1248) );
NOR2_X1 U986 ( .A1(G143), .A2(n1250), .ZN(n1251) );
NAND2_X1 U987 ( .A1(n1252), .A2(n1208), .ZN(n1245) );
INV_X1 U988 ( .A(G128), .ZN(n1208) );
NAND2_X1 U989 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NAND2_X1 U990 ( .A1(KEYINPUT39), .A2(n1255), .ZN(n1254) );
OR3_X1 U991 ( .A1(n1250), .A2(G143), .A3(KEYINPUT39), .ZN(n1253) );
XOR2_X1 U992 ( .A(n1256), .B(n1257), .Z(n1067) );
XOR2_X1 U993 ( .A(n1258), .B(n1259), .Z(n1257) );
XNOR2_X1 U994 ( .A(n1113), .B(G104), .ZN(n1259) );
XOR2_X1 U995 ( .A(KEYINPUT18), .B(G116), .Z(n1258) );
XNOR2_X1 U996 ( .A(n1102), .B(n1260), .ZN(n1256) );
XNOR2_X1 U997 ( .A(n1261), .B(n1235), .ZN(n1260) );
INV_X1 U998 ( .A(n1231), .ZN(n1235) );
NOR2_X1 U999 ( .A1(G122), .A2(KEYINPUT9), .ZN(n1261) );
XOR2_X1 U1000 ( .A(G101), .B(n1192), .Z(n1102) );
XOR2_X1 U1001 ( .A(G113), .B(G119), .Z(n1192) );
XNOR2_X1 U1002 ( .A(G125), .B(n1262), .ZN(n1243) );
NAND2_X1 U1003 ( .A1(KEYINPUT40), .A2(n1156), .ZN(n1262) );
NAND2_X1 U1004 ( .A1(G224), .A2(n1002), .ZN(n1156) );
AND2_X1 U1005 ( .A1(n1182), .A2(n1181), .ZN(n1014) );
XNOR2_X1 U1006 ( .A(n1042), .B(KEYINPUT57), .ZN(n1181) );
XNOR2_X1 U1007 ( .A(n1263), .B(n1264), .ZN(n1042) );
XNOR2_X1 U1008 ( .A(KEYINPUT21), .B(n1085), .ZN(n1264) );
INV_X1 U1009 ( .A(G475), .ZN(n1085) );
NAND2_X1 U1010 ( .A1(n1084), .A2(n1118), .ZN(n1263) );
XOR2_X1 U1011 ( .A(n1265), .B(n1266), .Z(n1084) );
XNOR2_X1 U1012 ( .A(G104), .B(n1267), .ZN(n1266) );
NAND2_X1 U1013 ( .A1(n1268), .A2(KEYINPUT15), .ZN(n1267) );
XOR2_X1 U1014 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U1015 ( .A(G131), .B(n1271), .ZN(n1270) );
XNOR2_X1 U1016 ( .A(KEYINPUT36), .B(KEYINPUT24), .ZN(n1271) );
XOR2_X1 U1017 ( .A(n1272), .B(n1202), .Z(n1269) );
XOR2_X1 U1018 ( .A(n1054), .B(KEYINPUT54), .Z(n1202) );
XOR2_X1 U1019 ( .A(G125), .B(G140), .Z(n1054) );
XNOR2_X1 U1020 ( .A(n1273), .B(n1255), .ZN(n1272) );
INV_X1 U1021 ( .A(n1240), .ZN(n1255) );
XNOR2_X1 U1022 ( .A(G143), .B(n1250), .ZN(n1240) );
INV_X1 U1023 ( .A(G146), .ZN(n1250) );
NAND4_X1 U1024 ( .A1(KEYINPUT23), .A2(G214), .A3(n1190), .A4(n1002), .ZN(n1273) );
INV_X1 U1025 ( .A(G237), .ZN(n1190) );
XNOR2_X1 U1026 ( .A(G113), .B(G122), .ZN(n1265) );
INV_X1 U1027 ( .A(n1041), .ZN(n1182) );
XOR2_X1 U1028 ( .A(G478), .B(n1274), .Z(n1041) );
AND2_X1 U1029 ( .A1(n1078), .A2(n1118), .ZN(n1274) );
INV_X1 U1030 ( .A(G902), .ZN(n1118) );
NAND2_X1 U1031 ( .A1(n1275), .A2(n1276), .ZN(n1078) );
NAND2_X1 U1032 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND3_X1 U1033 ( .A1(G234), .A2(n1002), .A3(G217), .ZN(n1278) );
INV_X1 U1034 ( .A(n1279), .ZN(n1277) );
XOR2_X1 U1035 ( .A(KEYINPUT53), .B(n1280), .Z(n1275) );
AND4_X1 U1036 ( .A1(n1002), .A2(G234), .A3(G217), .A4(n1279), .ZN(n1280) );
XNOR2_X1 U1037 ( .A(n1281), .B(n1282), .ZN(n1279) );
NOR2_X1 U1038 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
AND2_X1 U1039 ( .A1(n1285), .A2(n1220), .ZN(n1284) );
NOR2_X1 U1040 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
XNOR2_X1 U1041 ( .A(n1220), .B(KEYINPUT5), .ZN(n1286) );
XOR2_X1 U1042 ( .A(G134), .B(KEYINPUT56), .Z(n1220) );
AND2_X1 U1043 ( .A1(n1287), .A2(n1288), .ZN(n1285) );
NAND2_X1 U1044 ( .A1(G128), .A2(n1159), .ZN(n1288) );
XOR2_X1 U1045 ( .A(KEYINPUT31), .B(n1289), .Z(n1287) );
NOR2_X1 U1046 ( .A1(G128), .A2(n1159), .ZN(n1289) );
INV_X1 U1047 ( .A(G143), .ZN(n1159) );
NAND3_X1 U1048 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1281) );
NAND2_X1 U1049 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
OR3_X1 U1050 ( .A1(n1294), .A2(n1293), .A3(KEYINPUT62), .ZN(n1291) );
XOR2_X1 U1051 ( .A(n1231), .B(KEYINPUT50), .Z(n1293) );
XOR2_X1 U1052 ( .A(G107), .B(KEYINPUT59), .Z(n1231) );
OR2_X1 U1053 ( .A1(KEYINPUT42), .A2(n1295), .ZN(n1294) );
NAND2_X1 U1054 ( .A1(n1295), .A2(KEYINPUT62), .ZN(n1290) );
XOR2_X1 U1055 ( .A(G116), .B(n1296), .Z(n1295) );
XOR2_X1 U1056 ( .A(KEYINPUT11), .B(G122), .Z(n1296) );
INV_X1 U1057 ( .A(G953), .ZN(n1002) );
INV_X1 U1058 ( .A(G110), .ZN(n1113) );
endmodule


