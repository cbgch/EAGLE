//Key = 1110000101111011001001100010011011111110010011111110011010111001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402;

XNOR2_X1 U759 ( .A(G107), .B(n1072), .ZN(G9) );
NAND2_X1 U760 ( .A1(KEYINPUT47), .A2(n1073), .ZN(n1072) );
NOR2_X1 U761 ( .A1(n1074), .A2(n1075), .ZN(G75) );
NOR4_X1 U762 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075) );
XOR2_X1 U763 ( .A(KEYINPUT36), .B(n1080), .Z(n1077) );
NOR2_X1 U764 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR3_X1 U765 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NOR2_X1 U766 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U767 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U768 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U769 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
AND2_X1 U770 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
NOR3_X1 U771 ( .A1(n1096), .A2(n1093), .A3(n1097), .ZN(n1086) );
XOR2_X1 U772 ( .A(KEYINPUT48), .B(n1095), .Z(n1096) );
AND3_X1 U773 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1081) );
NAND3_X1 U774 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1076) );
NAND3_X1 U775 ( .A1(n1099), .A2(n1104), .A3(n1105), .ZN(n1103) );
INV_X1 U776 ( .A(n1083), .ZN(n1105) );
NAND2_X1 U777 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NAND3_X1 U778 ( .A1(n1108), .A2(n1109), .A3(n1095), .ZN(n1107) );
NAND2_X1 U779 ( .A1(n1110), .A2(n1111), .ZN(n1106) );
NAND2_X1 U780 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND3_X1 U781 ( .A1(n1114), .A2(n1095), .A3(n1115), .ZN(n1113) );
NAND3_X1 U782 ( .A1(n1108), .A2(n1116), .A3(n1117), .ZN(n1112) );
NAND3_X1 U783 ( .A1(n1110), .A2(n1118), .A3(n1098), .ZN(n1101) );
NOR3_X1 U784 ( .A1(n1119), .A2(n1093), .A3(n1083), .ZN(n1098) );
NOR3_X1 U785 ( .A1(n1078), .A2(G952), .A3(n1120), .ZN(n1074) );
INV_X1 U786 ( .A(n1102), .ZN(n1120) );
NAND4_X1 U787 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1102) );
NOR4_X1 U788 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1124) );
XOR2_X1 U789 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U790 ( .A(n1131), .B(n1132), .Z(n1127) );
NAND2_X1 U791 ( .A1(KEYINPUT2), .A2(n1133), .ZN(n1131) );
XOR2_X1 U792 ( .A(n1134), .B(n1135), .Z(n1126) );
XNOR2_X1 U793 ( .A(KEYINPUT45), .B(n1136), .ZN(n1135) );
NAND2_X1 U794 ( .A1(KEYINPUT30), .A2(G469), .ZN(n1134) );
XNOR2_X1 U795 ( .A(n1137), .B(KEYINPUT0), .ZN(n1125) );
NOR3_X1 U796 ( .A1(n1138), .A2(n1117), .A3(n1115), .ZN(n1123) );
NOR2_X1 U797 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
AND3_X1 U798 ( .A1(KEYINPUT63), .A2(n1141), .A3(n1142), .ZN(n1139) );
NAND2_X1 U799 ( .A1(n1141), .A2(n1143), .ZN(n1122) );
NAND2_X1 U800 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND3_X1 U801 ( .A1(n1142), .A2(n1140), .A3(KEYINPUT63), .ZN(n1145) );
NAND2_X1 U802 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
INV_X1 U803 ( .A(n1148), .ZN(n1147) );
NAND2_X1 U804 ( .A1(n1148), .A2(n1149), .ZN(n1121) );
NOR2_X1 U805 ( .A1(KEYINPUT27), .A2(n1150), .ZN(n1148) );
XOR2_X1 U806 ( .A(n1151), .B(KEYINPUT24), .Z(n1150) );
NAND3_X1 U807 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(G72) );
NAND2_X1 U808 ( .A1(KEYINPUT31), .A2(n1155), .ZN(n1154) );
OR3_X1 U809 ( .A1(n1155), .A2(KEYINPUT31), .A3(n1156), .ZN(n1153) );
NAND2_X1 U810 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
NAND2_X1 U811 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
INV_X1 U812 ( .A(KEYINPUT31), .ZN(n1159) );
XOR2_X1 U813 ( .A(n1155), .B(KEYINPUT54), .Z(n1158) );
NAND2_X1 U814 ( .A1(G953), .A2(n1160), .ZN(n1155) );
NAND2_X1 U815 ( .A1(G900), .A2(G227), .ZN(n1160) );
XNOR2_X1 U816 ( .A(n1161), .B(n1162), .ZN(n1156) );
NOR2_X1 U817 ( .A1(n1163), .A2(G953), .ZN(n1162) );
NAND3_X1 U818 ( .A1(n1164), .A2(n1165), .A3(KEYINPUT44), .ZN(n1161) );
NAND2_X1 U819 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U820 ( .A(KEYINPUT4), .B(G953), .Z(n1166) );
XOR2_X1 U821 ( .A(n1168), .B(n1169), .Z(n1164) );
XNOR2_X1 U822 ( .A(n1170), .B(n1171), .ZN(n1169) );
XOR2_X1 U823 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U824 ( .A1(KEYINPUT43), .A2(n1174), .ZN(n1172) );
XOR2_X1 U825 ( .A(G137), .B(n1175), .Z(n1168) );
XOR2_X1 U826 ( .A(KEYINPUT8), .B(G140), .Z(n1175) );
NAND2_X1 U827 ( .A1(n1176), .A2(n1177), .ZN(G69) );
NAND2_X1 U828 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
OR2_X1 U829 ( .A1(n1180), .A2(G224), .ZN(n1179) );
NAND3_X1 U830 ( .A1(n1181), .A2(n1182), .A3(G953), .ZN(n1176) );
NAND2_X1 U831 ( .A1(G898), .A2(G224), .ZN(n1182) );
XOR2_X1 U832 ( .A(KEYINPUT22), .B(n1178), .Z(n1181) );
XNOR2_X1 U833 ( .A(n1183), .B(n1184), .ZN(n1178) );
NOR2_X1 U834 ( .A1(n1185), .A2(G953), .ZN(n1184) );
NAND3_X1 U835 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1183) );
XOR2_X1 U836 ( .A(KEYINPUT12), .B(n1189), .Z(n1188) );
NOR2_X1 U837 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U838 ( .A1(n1191), .A2(n1190), .ZN(n1187) );
NAND2_X1 U839 ( .A1(n1192), .A2(n1193), .ZN(n1190) );
NAND3_X1 U840 ( .A1(n1194), .A2(n1195), .A3(n1196), .ZN(n1193) );
INV_X1 U841 ( .A(KEYINPUT56), .ZN(n1196) );
NAND2_X1 U842 ( .A1(n1197), .A2(KEYINPUT56), .ZN(n1192) );
XOR2_X1 U843 ( .A(KEYINPUT39), .B(n1198), .Z(n1191) );
NAND2_X1 U844 ( .A1(G953), .A2(n1199), .ZN(n1186) );
NOR2_X1 U845 ( .A1(n1200), .A2(n1201), .ZN(G66) );
NOR3_X1 U846 ( .A1(n1130), .A2(n1202), .A3(n1203), .ZN(n1201) );
NOR2_X1 U847 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
AND3_X1 U848 ( .A1(n1205), .A2(G902), .A3(n1204), .ZN(n1202) );
NOR3_X1 U849 ( .A1(KEYINPUT40), .A2(n1206), .A3(n1207), .ZN(n1204) );
INV_X1 U850 ( .A(G217), .ZN(n1207) );
NOR2_X1 U851 ( .A1(n1200), .A2(n1208), .ZN(G63) );
XNOR2_X1 U852 ( .A(n1142), .B(n1209), .ZN(n1208) );
NOR2_X1 U853 ( .A1(n1140), .A2(n1210), .ZN(n1209) );
INV_X1 U854 ( .A(G478), .ZN(n1140) );
NOR2_X1 U855 ( .A1(n1200), .A2(n1211), .ZN(G60) );
NOR3_X1 U856 ( .A1(n1132), .A2(n1212), .A3(n1213), .ZN(n1211) );
NOR3_X1 U857 ( .A1(n1214), .A2(n1210), .A3(n1133), .ZN(n1213) );
INV_X1 U858 ( .A(n1215), .ZN(n1214) );
NOR2_X1 U859 ( .A1(n1216), .A2(n1215), .ZN(n1212) );
NOR2_X1 U860 ( .A1(n1206), .A2(n1133), .ZN(n1216) );
INV_X1 U861 ( .A(n1079), .ZN(n1206) );
XOR2_X1 U862 ( .A(G104), .B(n1217), .Z(G6) );
NOR2_X1 U863 ( .A1(n1200), .A2(n1218), .ZN(G57) );
XOR2_X1 U864 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U865 ( .A1(KEYINPUT13), .A2(n1221), .ZN(n1220) );
XOR2_X1 U866 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR3_X1 U867 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1223) );
NOR3_X1 U868 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1226) );
AND3_X1 U869 ( .A1(n1227), .A2(n1230), .A3(n1228), .ZN(n1225) );
NOR2_X1 U870 ( .A1(n1230), .A2(n1231), .ZN(n1224) );
NAND3_X1 U871 ( .A1(G472), .A2(G902), .A3(n1232), .ZN(n1222) );
XOR2_X1 U872 ( .A(n1079), .B(KEYINPUT16), .Z(n1232) );
NAND3_X1 U873 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1219) );
NAND2_X1 U874 ( .A1(KEYINPUT20), .A2(n1236), .ZN(n1235) );
NAND3_X1 U875 ( .A1(n1237), .A2(n1238), .A3(G101), .ZN(n1234) );
NAND2_X1 U876 ( .A1(n1239), .A2(n1240), .ZN(n1233) );
NAND2_X1 U877 ( .A1(n1241), .A2(n1238), .ZN(n1239) );
INV_X1 U878 ( .A(KEYINPUT20), .ZN(n1238) );
XOR2_X1 U879 ( .A(n1236), .B(KEYINPUT60), .Z(n1241) );
NOR2_X1 U880 ( .A1(n1200), .A2(n1242), .ZN(G54) );
XOR2_X1 U881 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U882 ( .A(n1228), .B(n1245), .ZN(n1244) );
XOR2_X1 U883 ( .A(n1246), .B(n1247), .Z(n1243) );
NOR2_X1 U884 ( .A1(n1248), .A2(n1210), .ZN(n1247) );
INV_X1 U885 ( .A(G469), .ZN(n1248) );
NAND2_X1 U886 ( .A1(n1249), .A2(n1250), .ZN(n1246) );
NAND2_X1 U887 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U888 ( .A(n1253), .ZN(n1249) );
NOR2_X1 U889 ( .A1(n1200), .A2(n1254), .ZN(G51) );
NOR2_X1 U890 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U891 ( .A(KEYINPUT61), .B(n1257), .Z(n1256) );
NOR2_X1 U892 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U893 ( .A(KEYINPUT17), .B(n1260), .Z(n1259) );
AND2_X1 U894 ( .A1(n1258), .A2(n1260), .ZN(n1255) );
NOR2_X1 U895 ( .A1(n1210), .A2(n1151), .ZN(n1260) );
NAND2_X1 U896 ( .A1(G902), .A2(n1079), .ZN(n1210) );
NAND2_X1 U897 ( .A1(n1185), .A2(n1163), .ZN(n1079) );
AND4_X1 U898 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1163) );
NOR4_X1 U899 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1264) );
INV_X1 U900 ( .A(n1269), .ZN(n1268) );
AND2_X1 U901 ( .A1(n1270), .A2(n1271), .ZN(n1263) );
NAND4_X1 U902 ( .A1(n1272), .A2(n1273), .A3(n1274), .A4(n1275), .ZN(n1262) );
OR2_X1 U903 ( .A1(n1276), .A2(KEYINPUT25), .ZN(n1273) );
NAND2_X1 U904 ( .A1(KEYINPUT25), .A2(n1277), .ZN(n1272) );
NAND2_X1 U905 ( .A1(n1278), .A2(n1094), .ZN(n1277) );
INV_X1 U906 ( .A(n1279), .ZN(n1278) );
NAND2_X1 U907 ( .A1(n1280), .A2(n1095), .ZN(n1261) );
XOR2_X1 U908 ( .A(n1281), .B(KEYINPUT32), .Z(n1280) );
AND4_X1 U909 ( .A1(n1282), .A2(n1283), .A3(n1284), .A4(n1285), .ZN(n1185) );
NOR4_X1 U910 ( .A1(n1286), .A2(n1287), .A3(n1217), .A4(n1288), .ZN(n1285) );
AND3_X1 U911 ( .A1(n1289), .A2(n1099), .A3(n1290), .ZN(n1288) );
AND3_X1 U912 ( .A1(n1291), .A2(n1099), .A3(n1100), .ZN(n1217) );
NOR2_X1 U913 ( .A1(n1073), .A2(n1292), .ZN(n1284) );
AND3_X1 U914 ( .A1(n1109), .A2(n1099), .A3(n1291), .ZN(n1073) );
XNOR2_X1 U915 ( .A(n1293), .B(n1294), .ZN(n1258) );
XOR2_X1 U916 ( .A(n1229), .B(n1295), .Z(n1294) );
NOR2_X1 U917 ( .A1(n1180), .A2(G952), .ZN(n1200) );
XOR2_X1 U918 ( .A(n1296), .B(n1267), .Z(G48) );
AND4_X1 U919 ( .A1(n1276), .A2(n1274), .A3(n1100), .A4(n1297), .ZN(n1267) );
NAND2_X1 U920 ( .A1(KEYINPUT26), .A2(n1298), .ZN(n1296) );
INV_X1 U921 ( .A(G146), .ZN(n1298) );
XOR2_X1 U922 ( .A(n1299), .B(n1271), .Z(G45) );
NAND4_X1 U923 ( .A1(n1276), .A2(n1289), .A3(n1300), .A4(n1297), .ZN(n1271) );
XNOR2_X1 U924 ( .A(G140), .B(n1270), .ZN(G42) );
NAND4_X1 U925 ( .A1(n1276), .A2(n1095), .A3(n1100), .A4(n1118), .ZN(n1270) );
XOR2_X1 U926 ( .A(n1301), .B(n1302), .Z(G39) );
NOR2_X1 U927 ( .A1(n1266), .A2(KEYINPUT19), .ZN(n1302) );
AND4_X1 U928 ( .A1(n1276), .A2(n1095), .A3(n1274), .A4(n1110), .ZN(n1266) );
INV_X1 U929 ( .A(n1119), .ZN(n1095) );
NAND2_X1 U930 ( .A1(n1303), .A2(n1304), .ZN(G36) );
NAND2_X1 U931 ( .A1(n1265), .A2(n1305), .ZN(n1304) );
XOR2_X1 U932 ( .A(KEYINPUT1), .B(n1306), .Z(n1303) );
NOR2_X1 U933 ( .A1(n1265), .A2(n1305), .ZN(n1306) );
INV_X1 U934 ( .A(G134), .ZN(n1305) );
NOR4_X1 U935 ( .A1(n1307), .A2(n1119), .A3(n1097), .A4(n1308), .ZN(n1265) );
XOR2_X1 U936 ( .A(G131), .B(n1309), .Z(G33) );
NOR2_X1 U937 ( .A1(n1119), .A2(n1281), .ZN(n1309) );
NAND3_X1 U938 ( .A1(n1300), .A2(n1100), .A3(n1276), .ZN(n1281) );
NAND2_X1 U939 ( .A1(n1116), .A2(n1310), .ZN(n1119) );
XNOR2_X1 U940 ( .A(G128), .B(n1311), .ZN(G30) );
NAND4_X1 U941 ( .A1(KEYINPUT50), .A2(n1276), .A3(n1275), .A4(n1274), .ZN(n1311) );
NOR2_X1 U942 ( .A1(n1092), .A2(n1308), .ZN(n1275) );
INV_X1 U943 ( .A(n1297), .ZN(n1092) );
INV_X1 U944 ( .A(n1307), .ZN(n1276) );
NAND2_X1 U945 ( .A1(n1094), .A2(n1279), .ZN(n1307) );
XOR2_X1 U946 ( .A(G101), .B(n1287), .Z(G3) );
AND3_X1 U947 ( .A1(n1110), .A2(n1291), .A3(n1300), .ZN(n1287) );
XOR2_X1 U948 ( .A(n1174), .B(n1269), .Z(G27) );
NAND4_X1 U949 ( .A1(n1118), .A2(n1279), .A3(n1297), .A4(n1312), .ZN(n1269) );
AND2_X1 U950 ( .A1(n1108), .A2(n1100), .ZN(n1312) );
NAND2_X1 U951 ( .A1(n1083), .A2(n1313), .ZN(n1279) );
NAND4_X1 U952 ( .A1(G953), .A2(G902), .A3(n1314), .A4(n1167), .ZN(n1313) );
INV_X1 U953 ( .A(G900), .ZN(n1167) );
XOR2_X1 U954 ( .A(G122), .B(n1315), .Z(G24) );
NOR3_X1 U955 ( .A1(n1316), .A2(n1089), .A3(n1317), .ZN(n1315) );
INV_X1 U956 ( .A(n1099), .ZN(n1089) );
XOR2_X1 U957 ( .A(KEYINPUT53), .B(n1289), .Z(n1316) );
NOR2_X1 U958 ( .A1(n1318), .A2(n1319), .ZN(n1289) );
XOR2_X1 U959 ( .A(G119), .B(n1286), .Z(G21) );
AND3_X1 U960 ( .A1(n1290), .A2(n1110), .A3(n1274), .ZN(n1286) );
AND2_X1 U961 ( .A1(n1137), .A2(n1320), .ZN(n1274) );
XNOR2_X1 U962 ( .A(G116), .B(n1282), .ZN(G18) );
NAND3_X1 U963 ( .A1(n1290), .A2(n1109), .A3(n1300), .ZN(n1282) );
INV_X1 U964 ( .A(n1308), .ZN(n1109) );
NAND2_X1 U965 ( .A1(n1318), .A2(n1321), .ZN(n1308) );
XNOR2_X1 U966 ( .A(G113), .B(n1283), .ZN(G15) );
NAND3_X1 U967 ( .A1(n1290), .A2(n1100), .A3(n1300), .ZN(n1283) );
INV_X1 U968 ( .A(n1097), .ZN(n1300) );
NAND2_X1 U969 ( .A1(n1322), .A2(n1137), .ZN(n1097) );
NOR2_X1 U970 ( .A1(n1318), .A2(n1321), .ZN(n1100) );
INV_X1 U971 ( .A(n1319), .ZN(n1321) );
INV_X1 U972 ( .A(n1317), .ZN(n1290) );
NAND2_X1 U973 ( .A1(n1108), .A2(n1323), .ZN(n1317) );
INV_X1 U974 ( .A(n1093), .ZN(n1108) );
NAND2_X1 U975 ( .A1(n1114), .A2(n1324), .ZN(n1093) );
XOR2_X1 U976 ( .A(G110), .B(n1292), .Z(G12) );
AND3_X1 U977 ( .A1(n1291), .A2(n1118), .A3(n1110), .ZN(n1292) );
INV_X1 U978 ( .A(n1085), .ZN(n1110) );
NAND2_X1 U979 ( .A1(n1319), .A2(n1318), .ZN(n1085) );
XNOR2_X1 U980 ( .A(n1325), .B(n1326), .ZN(n1318) );
XOR2_X1 U981 ( .A(KEYINPUT62), .B(n1132), .Z(n1326) );
NOR2_X1 U982 ( .A1(n1215), .A2(G902), .ZN(n1132) );
XNOR2_X1 U983 ( .A(n1327), .B(n1328), .ZN(n1215) );
XOR2_X1 U984 ( .A(G122), .B(G113), .Z(n1328) );
XOR2_X1 U985 ( .A(n1329), .B(G104), .Z(n1327) );
NAND2_X1 U986 ( .A1(KEYINPUT18), .A2(n1330), .ZN(n1329) );
XOR2_X1 U987 ( .A(n1331), .B(n1332), .Z(n1330) );
XOR2_X1 U988 ( .A(n1333), .B(n1334), .Z(n1332) );
AND2_X1 U989 ( .A1(G214), .A2(n1335), .ZN(n1334) );
NAND2_X1 U990 ( .A1(KEYINPUT46), .A2(n1336), .ZN(n1333) );
XOR2_X1 U991 ( .A(n1337), .B(n1338), .Z(n1336) );
NOR2_X1 U992 ( .A1(G146), .A2(KEYINPUT23), .ZN(n1337) );
XOR2_X1 U993 ( .A(G131), .B(n1299), .Z(n1331) );
NAND2_X1 U994 ( .A1(KEYINPUT29), .A2(n1133), .ZN(n1325) );
INV_X1 U995 ( .A(G475), .ZN(n1133) );
XOR2_X1 U996 ( .A(n1339), .B(G478), .Z(n1319) );
NAND2_X1 U997 ( .A1(n1141), .A2(n1142), .ZN(n1339) );
NAND2_X1 U998 ( .A1(n1340), .A2(n1341), .ZN(n1142) );
NAND2_X1 U999 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1000 ( .A(n1344), .B(KEYINPUT5), .Z(n1340) );
OR2_X1 U1001 ( .A1(n1343), .A2(n1342), .ZN(n1344) );
AND3_X1 U1002 ( .A1(G234), .A2(n1180), .A3(G217), .ZN(n1342) );
XNOR2_X1 U1003 ( .A(n1345), .B(n1346), .ZN(n1343) );
XOR2_X1 U1004 ( .A(G128), .B(n1347), .Z(n1346) );
XOR2_X1 U1005 ( .A(G143), .B(G134), .Z(n1347) );
XOR2_X1 U1006 ( .A(n1348), .B(n1349), .Z(n1345) );
NOR2_X1 U1007 ( .A1(G107), .A2(KEYINPUT6), .ZN(n1349) );
XOR2_X1 U1008 ( .A(n1350), .B(G116), .Z(n1348) );
NAND2_X1 U1009 ( .A1(KEYINPUT9), .A2(G122), .ZN(n1350) );
NAND2_X1 U1010 ( .A1(n1351), .A2(n1352), .ZN(n1118) );
OR3_X1 U1011 ( .A1(n1322), .A2(n1137), .A3(KEYINPUT55), .ZN(n1352) );
NAND2_X1 U1012 ( .A1(KEYINPUT55), .A2(n1099), .ZN(n1351) );
NOR2_X1 U1013 ( .A1(n1320), .A2(n1137), .ZN(n1099) );
XNOR2_X1 U1014 ( .A(n1353), .B(G472), .ZN(n1137) );
NAND2_X1 U1015 ( .A1(n1354), .A2(n1141), .ZN(n1353) );
XOR2_X1 U1016 ( .A(n1355), .B(n1356), .Z(n1354) );
XOR2_X1 U1017 ( .A(n1231), .B(n1237), .Z(n1356) );
INV_X1 U1018 ( .A(n1236), .ZN(n1237) );
NAND2_X1 U1019 ( .A1(n1335), .A2(G210), .ZN(n1236) );
NOR2_X1 U1020 ( .A1(G953), .A2(G237), .ZN(n1335) );
XNOR2_X1 U1021 ( .A(n1228), .B(n1227), .ZN(n1231) );
XNOR2_X1 U1022 ( .A(n1357), .B(n1358), .ZN(n1227) );
NAND2_X1 U1023 ( .A1(KEYINPUT38), .A2(G113), .ZN(n1357) );
XOR2_X1 U1024 ( .A(n1359), .B(n1360), .Z(n1355) );
XOR2_X1 U1025 ( .A(KEYINPUT42), .B(G101), .Z(n1360) );
NAND2_X1 U1026 ( .A1(KEYINPUT49), .A2(n1229), .ZN(n1359) );
INV_X1 U1027 ( .A(n1322), .ZN(n1320) );
XOR2_X1 U1028 ( .A(n1361), .B(n1130), .Z(n1322) );
NOR2_X1 U1029 ( .A1(n1205), .A2(G902), .ZN(n1130) );
XOR2_X1 U1030 ( .A(n1362), .B(n1363), .Z(n1205) );
XOR2_X1 U1031 ( .A(G110), .B(n1364), .Z(n1363) );
XOR2_X1 U1032 ( .A(G137), .B(G119), .Z(n1364) );
XOR2_X1 U1033 ( .A(n1365), .B(n1338), .Z(n1362) );
XOR2_X1 U1034 ( .A(G125), .B(G140), .Z(n1338) );
XOR2_X1 U1035 ( .A(n1366), .B(n1367), .Z(n1365) );
NAND3_X1 U1036 ( .A1(G234), .A2(n1180), .A3(G221), .ZN(n1366) );
NAND2_X1 U1037 ( .A1(KEYINPUT7), .A2(n1129), .ZN(n1361) );
AND2_X1 U1038 ( .A1(G217), .A2(n1368), .ZN(n1129) );
AND2_X1 U1039 ( .A1(n1323), .A2(n1094), .ZN(n1291) );
NOR2_X1 U1040 ( .A1(n1114), .A2(n1115), .ZN(n1094) );
INV_X1 U1041 ( .A(n1324), .ZN(n1115) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1368), .ZN(n1324) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1141), .ZN(n1368) );
XOR2_X1 U1044 ( .A(n1136), .B(G469), .Z(n1114) );
NAND2_X1 U1045 ( .A1(n1369), .A2(n1141), .ZN(n1136) );
XOR2_X1 U1046 ( .A(n1370), .B(n1371), .Z(n1369) );
NOR2_X1 U1047 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
NOR3_X1 U1048 ( .A1(KEYINPUT21), .A2(n1374), .A3(n1170), .ZN(n1373) );
NOR2_X1 U1049 ( .A1(n1245), .A2(n1375), .ZN(n1372) );
INV_X1 U1050 ( .A(KEYINPUT21), .ZN(n1375) );
XNOR2_X1 U1051 ( .A(n1374), .B(n1170), .ZN(n1245) );
XOR2_X1 U1052 ( .A(n1229), .B(KEYINPUT15), .Z(n1170) );
XNOR2_X1 U1053 ( .A(n1376), .B(n1377), .ZN(n1374) );
XOR2_X1 U1054 ( .A(KEYINPUT52), .B(G107), .Z(n1377) );
XOR2_X1 U1055 ( .A(G104), .B(n1240), .Z(n1376) );
INV_X1 U1056 ( .A(G101), .ZN(n1240) );
XNOR2_X1 U1057 ( .A(n1228), .B(n1378), .ZN(n1370) );
NOR3_X1 U1058 ( .A1(n1253), .A2(n1379), .A3(n1380), .ZN(n1378) );
AND3_X1 U1059 ( .A1(KEYINPUT33), .A2(n1252), .A3(n1251), .ZN(n1380) );
NOR2_X1 U1060 ( .A1(KEYINPUT33), .A2(n1251), .ZN(n1379) );
NOR2_X1 U1061 ( .A1(n1252), .A2(n1251), .ZN(n1253) );
XOR2_X1 U1062 ( .A(G110), .B(G140), .Z(n1251) );
NAND2_X1 U1063 ( .A1(G227), .A2(n1180), .ZN(n1252) );
XNOR2_X1 U1064 ( .A(n1381), .B(KEYINPUT58), .ZN(n1228) );
NAND2_X1 U1065 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
NAND2_X1 U1066 ( .A1(n1384), .A2(n1301), .ZN(n1383) );
INV_X1 U1067 ( .A(G137), .ZN(n1301) );
XOR2_X1 U1068 ( .A(KEYINPUT11), .B(n1173), .Z(n1384) );
NAND2_X1 U1069 ( .A1(n1173), .A2(G137), .ZN(n1382) );
XOR2_X1 U1070 ( .A(G131), .B(n1385), .Z(n1173) );
XOR2_X1 U1071 ( .A(KEYINPUT57), .B(G134), .Z(n1385) );
AND2_X1 U1072 ( .A1(n1297), .A2(n1386), .ZN(n1323) );
NAND2_X1 U1073 ( .A1(n1083), .A2(n1387), .ZN(n1386) );
NAND4_X1 U1074 ( .A1(G953), .A2(G902), .A3(n1314), .A4(n1199), .ZN(n1387) );
INV_X1 U1075 ( .A(G898), .ZN(n1199) );
NAND3_X1 U1076 ( .A1(n1388), .A2(n1314), .A3(G952), .ZN(n1083) );
NAND2_X1 U1077 ( .A1(G237), .A2(G234), .ZN(n1314) );
INV_X1 U1078 ( .A(n1078), .ZN(n1388) );
XOR2_X1 U1079 ( .A(n1180), .B(KEYINPUT10), .Z(n1078) );
NOR2_X1 U1080 ( .A1(n1116), .A2(n1117), .ZN(n1297) );
INV_X1 U1081 ( .A(n1310), .ZN(n1117) );
NAND2_X1 U1082 ( .A1(G214), .A2(n1389), .ZN(n1310) );
XOR2_X1 U1083 ( .A(n1390), .B(n1151), .Z(n1116) );
NAND2_X1 U1084 ( .A1(G210), .A2(n1389), .ZN(n1151) );
NAND2_X1 U1085 ( .A1(n1391), .A2(n1141), .ZN(n1389) );
INV_X1 U1086 ( .A(G237), .ZN(n1391) );
NAND2_X1 U1087 ( .A1(KEYINPUT41), .A2(n1149), .ZN(n1390) );
NAND2_X1 U1088 ( .A1(n1146), .A2(n1141), .ZN(n1149) );
INV_X1 U1089 ( .A(G902), .ZN(n1141) );
XNOR2_X1 U1090 ( .A(n1392), .B(n1393), .ZN(n1146) );
XOR2_X1 U1091 ( .A(KEYINPUT28), .B(n1394), .Z(n1393) );
NOR2_X1 U1092 ( .A1(KEYINPUT51), .A2(n1230), .ZN(n1394) );
INV_X1 U1093 ( .A(n1229), .ZN(n1230) );
XOR2_X1 U1094 ( .A(n1299), .B(n1367), .Z(n1229) );
XOR2_X1 U1095 ( .A(G128), .B(G146), .Z(n1367) );
INV_X1 U1096 ( .A(G143), .ZN(n1299) );
XNOR2_X1 U1097 ( .A(n1293), .B(n1295), .ZN(n1392) );
XNOR2_X1 U1098 ( .A(n1395), .B(n1174), .ZN(n1295) );
INV_X1 U1099 ( .A(G125), .ZN(n1174) );
NAND2_X1 U1100 ( .A1(n1396), .A2(n1180), .ZN(n1395) );
INV_X1 U1101 ( .A(G953), .ZN(n1180) );
XNOR2_X1 U1102 ( .A(G224), .B(KEYINPUT59), .ZN(n1396) );
XNOR2_X1 U1103 ( .A(n1197), .B(n1198), .ZN(n1293) );
XOR2_X1 U1104 ( .A(G110), .B(n1397), .Z(n1198) );
XOR2_X1 U1105 ( .A(KEYINPUT35), .B(G122), .Z(n1397) );
XOR2_X1 U1106 ( .A(n1195), .B(n1194), .Z(n1197) );
XNOR2_X1 U1107 ( .A(n1398), .B(n1399), .ZN(n1194) );
XOR2_X1 U1108 ( .A(KEYINPUT3), .B(G104), .Z(n1399) );
XOR2_X1 U1109 ( .A(n1400), .B(G101), .Z(n1398) );
NAND2_X1 U1110 ( .A1(KEYINPUT34), .A2(G107), .ZN(n1400) );
XNOR2_X1 U1111 ( .A(n1401), .B(n1402), .ZN(n1195) );
XOR2_X1 U1112 ( .A(KEYINPUT37), .B(KEYINPUT14), .Z(n1402) );
XNOR2_X1 U1113 ( .A(G113), .B(n1358), .ZN(n1401) );
XOR2_X1 U1114 ( .A(G116), .B(G119), .Z(n1358) );
endmodule


