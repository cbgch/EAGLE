//Key = 1111110010100001000101110001011100111110100111110001101001001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312;

XNOR2_X1 U720 ( .A(n998), .B(n999), .ZN(G9) );
NOR2_X1 U721 ( .A1(n1000), .A2(n1001), .ZN(G75) );
NOR4_X1 U722 ( .A1(n1002), .A2(n1003), .A3(G953), .A4(n1004), .ZN(n1001) );
NOR2_X1 U723 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NOR2_X1 U724 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR2_X1 U725 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NOR2_X1 U726 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NOR4_X1 U727 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NOR3_X1 U728 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1014) );
NOR2_X1 U729 ( .A1(n1020), .A2(n1021), .ZN(n1013) );
NOR3_X1 U730 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1011) );
XOR2_X1 U731 ( .A(n1016), .B(KEYINPUT50), .Z(n1024) );
NOR3_X1 U732 ( .A1(n1025), .A2(n1026), .A3(n1023), .ZN(n1007) );
NOR3_X1 U733 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
NOR2_X1 U734 ( .A1(n1030), .A2(n1010), .ZN(n1029) );
NOR2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR3_X1 U736 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1031) );
INV_X1 U737 ( .A(n1036), .ZN(n1035) );
NOR2_X1 U738 ( .A1(n1037), .A2(n1038), .ZN(n1028) );
XOR2_X1 U739 ( .A(n1016), .B(KEYINPUT16), .Z(n1037) );
NOR2_X1 U740 ( .A1(n1039), .A2(n1016), .ZN(n1027) );
NAND2_X1 U741 ( .A1(n1040), .A2(n1041), .ZN(n1002) );
NOR3_X1 U742 ( .A1(n1004), .A2(G953), .A3(G952), .ZN(n1000) );
AND4_X1 U743 ( .A1(n1042), .A2(n1033), .A3(n1043), .A4(n1044), .ZN(n1004) );
NOR4_X1 U744 ( .A1(n1045), .A2(n1046), .A3(n1010), .A4(n1047), .ZN(n1044) );
XOR2_X1 U745 ( .A(n1048), .B(KEYINPUT8), .Z(n1045) );
NOR3_X1 U746 ( .A1(n1034), .A2(n1049), .A3(n1017), .ZN(n1043) );
INV_X1 U747 ( .A(n1021), .ZN(n1017) );
INV_X1 U748 ( .A(n1050), .ZN(n1034) );
NAND2_X1 U749 ( .A1(G469), .A2(n1051), .ZN(n1042) );
XOR2_X1 U750 ( .A(n1052), .B(n1053), .Z(G72) );
XOR2_X1 U751 ( .A(n1054), .B(n1055), .Z(n1053) );
NAND2_X1 U752 ( .A1(G953), .A2(n1056), .ZN(n1055) );
NAND2_X1 U753 ( .A1(G900), .A2(G227), .ZN(n1056) );
NAND2_X1 U754 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
NAND2_X1 U755 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U756 ( .A(n1061), .B(n1062), .Z(n1057) );
XOR2_X1 U757 ( .A(n1063), .B(n1064), .Z(n1062) );
XNOR2_X1 U758 ( .A(n1065), .B(n1066), .ZN(n1064) );
XNOR2_X1 U759 ( .A(G134), .B(n1067), .ZN(n1061) );
XNOR2_X1 U760 ( .A(KEYINPUT12), .B(n1068), .ZN(n1067) );
NOR2_X1 U761 ( .A1(n1041), .A2(G953), .ZN(n1052) );
NAND2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(G69) );
NAND3_X1 U763 ( .A1(G953), .A2(n1071), .A3(n1072), .ZN(n1070) );
XNOR2_X1 U764 ( .A(n1073), .B(KEYINPUT24), .ZN(n1072) );
XOR2_X1 U765 ( .A(n1074), .B(KEYINPUT49), .Z(n1069) );
NAND2_X1 U766 ( .A1(n1073), .A2(n1075), .ZN(n1074) );
NAND2_X1 U767 ( .A1(G953), .A2(n1071), .ZN(n1075) );
NAND2_X1 U768 ( .A1(G898), .A2(G224), .ZN(n1071) );
XNOR2_X1 U769 ( .A(n1076), .B(n1077), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1040), .A2(G953), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
XOR2_X1 U772 ( .A(KEYINPUT4), .B(n1080), .Z(n1079) );
NOR2_X1 U773 ( .A1(G898), .A2(n1081), .ZN(n1080) );
XOR2_X1 U774 ( .A(n1082), .B(KEYINPUT23), .Z(n1078) );
NOR2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(G66) );
XOR2_X1 U776 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U778 ( .A1(n1083), .A2(n1089), .ZN(G63) );
XOR2_X1 U779 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR2_X1 U780 ( .A1(KEYINPUT25), .A2(n1092), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1093), .A2(n1087), .ZN(n1090) );
XNOR2_X1 U782 ( .A(G478), .B(KEYINPUT47), .ZN(n1093) );
NOR2_X1 U783 ( .A1(n1083), .A2(n1094), .ZN(G60) );
NOR3_X1 U784 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
AND2_X1 U785 ( .A1(n1098), .A2(KEYINPUT61), .ZN(n1097) );
NOR3_X1 U786 ( .A1(KEYINPUT61), .A2(n1099), .A3(n1098), .ZN(n1096) );
NOR3_X1 U787 ( .A1(n1100), .A2(KEYINPUT41), .A3(n1101), .ZN(n1099) );
NOR3_X1 U788 ( .A1(n1100), .A2(n1102), .A3(n1101), .ZN(n1095) );
INV_X1 U789 ( .A(G475), .ZN(n1101) );
NOR2_X1 U790 ( .A1(n1103), .A2(KEYINPUT61), .ZN(n1102) );
NOR2_X1 U791 ( .A1(KEYINPUT41), .A2(n1104), .ZN(n1103) );
INV_X1 U792 ( .A(n1098), .ZN(n1104) );
NAND2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(G6) );
NAND2_X1 U794 ( .A1(G104), .A2(n1107), .ZN(n1106) );
XOR2_X1 U795 ( .A(KEYINPUT40), .B(n1108), .Z(n1105) );
NOR2_X1 U796 ( .A1(G104), .A2(n1107), .ZN(n1108) );
INV_X1 U797 ( .A(n1109), .ZN(n1107) );
NOR2_X1 U798 ( .A1(n1083), .A2(n1110), .ZN(G57) );
XOR2_X1 U799 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U800 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(n1111) );
NAND2_X1 U802 ( .A1(n1087), .A2(G472), .ZN(n1115) );
NOR2_X1 U803 ( .A1(n1083), .A2(n1117), .ZN(G54) );
XOR2_X1 U804 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U805 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U806 ( .A(n1122), .B(n1063), .Z(n1120) );
NAND2_X1 U807 ( .A1(KEYINPUT30), .A2(n1123), .ZN(n1122) );
XOR2_X1 U808 ( .A(n1124), .B(n1125), .Z(n1118) );
XNOR2_X1 U809 ( .A(G140), .B(n1126), .ZN(n1125) );
XOR2_X1 U810 ( .A(n1127), .B(n1128), .Z(n1124) );
NAND2_X1 U811 ( .A1(n1087), .A2(G469), .ZN(n1127) );
NOR2_X1 U812 ( .A1(n1083), .A2(n1129), .ZN(G51) );
XOR2_X1 U813 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U814 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U815 ( .A1(KEYINPUT36), .A2(n1134), .ZN(n1133) );
NAND2_X1 U816 ( .A1(n1087), .A2(G210), .ZN(n1132) );
INV_X1 U817 ( .A(n1100), .ZN(n1087) );
NAND2_X1 U818 ( .A1(G902), .A2(n1135), .ZN(n1100) );
NAND2_X1 U819 ( .A1(n1136), .A2(n1041), .ZN(n1135) );
AND4_X1 U820 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1041) );
NOR4_X1 U821 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
AND2_X1 U822 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
XNOR2_X1 U823 ( .A(n1040), .B(KEYINPUT2), .ZN(n1136) );
AND4_X1 U824 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1040) );
NOR4_X1 U825 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n999), .ZN(n1150) );
NOR3_X1 U826 ( .A1(n1154), .A2(n1023), .A3(n1038), .ZN(n999) );
INV_X1 U827 ( .A(n1155), .ZN(n1038) );
NOR2_X1 U828 ( .A1(n1109), .A2(n1156), .ZN(n1149) );
NOR3_X1 U829 ( .A1(n1157), .A2(n1158), .A3(n1154), .ZN(n1156) );
XNOR2_X1 U830 ( .A(KEYINPUT60), .B(n1010), .ZN(n1157) );
NOR3_X1 U831 ( .A1(n1154), .A2(n1023), .A3(n1039), .ZN(n1109) );
INV_X1 U832 ( .A(n1020), .ZN(n1023) );
XNOR2_X1 U833 ( .A(n1159), .B(n1160), .ZN(n1130) );
NOR2_X1 U834 ( .A1(n1161), .A2(G952), .ZN(n1083) );
XOR2_X1 U835 ( .A(n1144), .B(n1162), .Z(G48) );
NOR2_X1 U836 ( .A1(KEYINPUT17), .A2(n1163), .ZN(n1162) );
AND3_X1 U837 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1144) );
XOR2_X1 U838 ( .A(n1143), .B(n1167), .Z(G45) );
NOR2_X1 U839 ( .A1(KEYINPUT18), .A2(n1168), .ZN(n1167) );
AND3_X1 U840 ( .A1(n1169), .A2(n1018), .A3(n1166), .ZN(n1143) );
XNOR2_X1 U841 ( .A(G140), .B(n1146), .ZN(G42) );
NAND3_X1 U842 ( .A1(n1164), .A2(n1019), .A3(n1170), .ZN(n1146) );
XNOR2_X1 U843 ( .A(n1142), .B(n1171), .ZN(G39) );
XNOR2_X1 U844 ( .A(G137), .B(KEYINPUT55), .ZN(n1171) );
AND4_X1 U845 ( .A1(n1172), .A2(n1170), .A3(n1173), .A4(n1047), .ZN(n1142) );
XNOR2_X1 U846 ( .A(G134), .B(n1145), .ZN(G36) );
NAND3_X1 U847 ( .A1(n1018), .A2(n1155), .A3(n1170), .ZN(n1145) );
XNOR2_X1 U848 ( .A(G131), .B(n1137), .ZN(G33) );
NAND3_X1 U849 ( .A1(n1164), .A2(n1018), .A3(n1170), .ZN(n1137) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1016), .ZN(n1170) );
NAND3_X1 U851 ( .A1(n1033), .A2(n1050), .A3(n1036), .ZN(n1016) );
INV_X1 U852 ( .A(n1166), .ZN(n1174) );
NOR2_X1 U853 ( .A1(n1022), .A2(n1175), .ZN(n1166) );
INV_X1 U854 ( .A(n1176), .ZN(n1175) );
XNOR2_X1 U855 ( .A(G128), .B(n1138), .ZN(G30) );
NAND4_X1 U856 ( .A1(n1165), .A2(n1155), .A3(n1177), .A4(n1176), .ZN(n1138) );
XNOR2_X1 U857 ( .A(G101), .B(n1147), .ZN(G3) );
NAND2_X1 U858 ( .A1(n1178), .A2(n1018), .ZN(n1147) );
XOR2_X1 U859 ( .A(n1141), .B(n1179), .Z(G27) );
NOR2_X1 U860 ( .A1(KEYINPUT42), .A2(n1134), .ZN(n1179) );
AND4_X1 U861 ( .A1(n1032), .A2(n1176), .A3(n1019), .A4(n1180), .ZN(n1141) );
NOR2_X1 U862 ( .A1(n1025), .A2(n1039), .ZN(n1180) );
NAND2_X1 U863 ( .A1(n1006), .A2(n1181), .ZN(n1176) );
NAND4_X1 U864 ( .A1(G902), .A2(n1059), .A3(n1182), .A4(n1060), .ZN(n1181) );
INV_X1 U865 ( .A(G900), .ZN(n1060) );
XOR2_X1 U866 ( .A(G122), .B(n1153), .Z(G24) );
AND3_X1 U867 ( .A1(n1183), .A2(n1020), .A3(n1169), .ZN(n1153) );
AND3_X1 U868 ( .A1(n1184), .A2(n1185), .A3(n1032), .ZN(n1169) );
NAND2_X1 U869 ( .A1(n1186), .A2(n1187), .ZN(n1020) );
OR3_X1 U870 ( .A1(n1046), .A2(n1047), .A3(KEYINPUT48), .ZN(n1187) );
NAND2_X1 U871 ( .A1(KEYINPUT48), .A2(n1019), .ZN(n1186) );
XNOR2_X1 U872 ( .A(G119), .B(n1188), .ZN(G21) );
NAND2_X1 U873 ( .A1(KEYINPUT19), .A2(n1152), .ZN(n1188) );
AND3_X1 U874 ( .A1(n1183), .A2(n1173), .A3(n1165), .ZN(n1152) );
AND3_X1 U875 ( .A1(n1032), .A2(n1047), .A3(n1172), .ZN(n1165) );
XNOR2_X1 U876 ( .A(n1046), .B(KEYINPUT37), .ZN(n1172) );
XOR2_X1 U877 ( .A(G116), .B(n1151), .Z(G18) );
AND4_X1 U878 ( .A1(n1183), .A2(n1018), .A3(n1155), .A4(n1032), .ZN(n1151) );
NOR2_X1 U879 ( .A1(n1184), .A2(n1189), .ZN(n1155) );
XNOR2_X1 U880 ( .A(G113), .B(n1148), .ZN(G15) );
NAND4_X1 U881 ( .A1(n1164), .A2(n1183), .A3(n1190), .A4(n1018), .ZN(n1148) );
NOR2_X1 U882 ( .A1(n1047), .A2(n1191), .ZN(n1018) );
NOR2_X1 U883 ( .A1(n1025), .A2(n1192), .ZN(n1183) );
INV_X1 U884 ( .A(n1193), .ZN(n1192) );
NAND2_X1 U885 ( .A1(n1194), .A2(n1021), .ZN(n1025) );
INV_X1 U886 ( .A(n1039), .ZN(n1164) );
NAND2_X1 U887 ( .A1(n1189), .A2(n1184), .ZN(n1039) );
INV_X1 U888 ( .A(n1185), .ZN(n1189) );
XNOR2_X1 U889 ( .A(G110), .B(n1195), .ZN(G12) );
NAND2_X1 U890 ( .A1(n1178), .A2(n1019), .ZN(n1195) );
INV_X1 U891 ( .A(n1158), .ZN(n1019) );
NAND2_X1 U892 ( .A1(n1191), .A2(n1047), .ZN(n1158) );
XNOR2_X1 U893 ( .A(n1196), .B(n1088), .ZN(n1047) );
AND2_X1 U894 ( .A1(G217), .A2(n1197), .ZN(n1088) );
NAND2_X1 U895 ( .A1(n1086), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U896 ( .A(n1199), .B(n1200), .ZN(n1086) );
XOR2_X1 U897 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U898 ( .A(n1203), .B(n1066), .Z(n1202) );
NAND2_X1 U899 ( .A1(KEYINPUT27), .A2(n1204), .ZN(n1203) );
XNOR2_X1 U900 ( .A(G137), .B(n1205), .ZN(n1204) );
NAND2_X1 U901 ( .A1(G221), .A2(n1206), .ZN(n1205) );
XNOR2_X1 U902 ( .A(n1207), .B(n1126), .ZN(n1201) );
NAND2_X1 U903 ( .A1(n1208), .A2(KEYINPUT57), .ZN(n1207) );
XNOR2_X1 U904 ( .A(G119), .B(KEYINPUT10), .ZN(n1208) );
XOR2_X1 U905 ( .A(n1209), .B(n1210), .Z(n1199) );
XNOR2_X1 U906 ( .A(n1163), .B(G128), .ZN(n1210) );
INV_X1 U907 ( .A(G146), .ZN(n1163) );
XNOR2_X1 U908 ( .A(KEYINPUT29), .B(KEYINPUT21), .ZN(n1209) );
INV_X1 U909 ( .A(n1046), .ZN(n1191) );
XNOR2_X1 U910 ( .A(n1211), .B(G472), .ZN(n1046) );
NAND2_X1 U911 ( .A1(n1212), .A2(n1198), .ZN(n1211) );
XOR2_X1 U912 ( .A(n1213), .B(n1214), .Z(n1212) );
XNOR2_X1 U913 ( .A(n1215), .B(n1113), .ZN(n1214) );
XNOR2_X1 U914 ( .A(n1216), .B(n1217), .ZN(n1113) );
NAND3_X1 U915 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1215) );
NAND2_X1 U916 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
OR3_X1 U917 ( .A1(n1222), .A2(n1221), .A3(n1116), .ZN(n1219) );
INV_X1 U918 ( .A(KEYINPUT46), .ZN(n1222) );
NAND2_X1 U919 ( .A1(n1116), .A2(n1223), .ZN(n1218) );
NAND2_X1 U920 ( .A1(n1224), .A2(KEYINPUT46), .ZN(n1223) );
XNOR2_X1 U921 ( .A(n1221), .B(KEYINPUT20), .ZN(n1224) );
XOR2_X1 U922 ( .A(n1225), .B(KEYINPUT28), .Z(n1221) );
AND3_X1 U923 ( .A1(n1226), .A2(n1161), .A3(G210), .ZN(n1116) );
NOR2_X1 U924 ( .A1(n1010), .A2(n1154), .ZN(n1178) );
NAND3_X1 U925 ( .A1(n1190), .A2(n1193), .A3(n1177), .ZN(n1154) );
XOR2_X1 U926 ( .A(n1022), .B(KEYINPUT38), .Z(n1177) );
NAND2_X1 U927 ( .A1(n1021), .A2(n1015), .ZN(n1022) );
INV_X1 U928 ( .A(n1194), .ZN(n1015) );
NOR2_X1 U929 ( .A1(n1227), .A2(n1049), .ZN(n1194) );
NOR2_X1 U930 ( .A1(n1051), .A2(G469), .ZN(n1049) );
AND2_X1 U931 ( .A1(n1228), .A2(n1051), .ZN(n1227) );
NAND2_X1 U932 ( .A1(n1229), .A2(n1198), .ZN(n1051) );
XOR2_X1 U933 ( .A(n1230), .B(n1231), .Z(n1229) );
NAND3_X1 U934 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
NAND2_X1 U935 ( .A1(KEYINPUT59), .A2(n1235), .ZN(n1234) );
NAND3_X1 U936 ( .A1(n1236), .A2(n1237), .A3(n1121), .ZN(n1233) );
INV_X1 U937 ( .A(KEYINPUT59), .ZN(n1237) );
OR2_X1 U938 ( .A1(n1121), .A2(n1236), .ZN(n1232) );
NOR2_X1 U939 ( .A1(KEYINPUT9), .A2(n1235), .ZN(n1236) );
XNOR2_X1 U940 ( .A(n1123), .B(n1063), .ZN(n1235) );
XNOR2_X1 U941 ( .A(n1238), .B(G128), .ZN(n1063) );
NAND2_X1 U942 ( .A1(KEYINPUT63), .A2(n1239), .ZN(n1238) );
XOR2_X1 U943 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U944 ( .A(KEYINPUT54), .B(n1168), .ZN(n1241) );
NOR2_X1 U945 ( .A1(G146), .A2(KEYINPUT39), .ZN(n1240) );
NAND2_X1 U946 ( .A1(n1242), .A2(n1243), .ZN(n1123) );
NAND2_X1 U947 ( .A1(n1244), .A2(n1225), .ZN(n1243) );
XOR2_X1 U948 ( .A(n1245), .B(KEYINPUT14), .Z(n1242) );
OR2_X1 U949 ( .A1(n1225), .A2(n1244), .ZN(n1245) );
XNOR2_X1 U950 ( .A(G104), .B(n998), .ZN(n1244) );
INV_X1 U951 ( .A(G107), .ZN(n998) );
XOR2_X1 U952 ( .A(n1217), .B(KEYINPUT1), .Z(n1121) );
XNOR2_X1 U953 ( .A(n1246), .B(n1247), .ZN(n1217) );
XNOR2_X1 U954 ( .A(KEYINPUT45), .B(n1065), .ZN(n1247) );
NAND2_X1 U955 ( .A1(n1248), .A2(KEYINPUT22), .ZN(n1246) );
XNOR2_X1 U956 ( .A(n1249), .B(n1068), .ZN(n1248) );
INV_X1 U957 ( .A(G137), .ZN(n1068) );
NAND2_X1 U958 ( .A1(KEYINPUT43), .A2(n1250), .ZN(n1249) );
NAND2_X1 U959 ( .A1(n1251), .A2(n1252), .ZN(n1230) );
NAND2_X1 U960 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U961 ( .A(n1255), .B(n1128), .Z(n1251) );
AND2_X1 U962 ( .A1(G227), .A2(n1161), .ZN(n1128) );
OR2_X1 U963 ( .A1(n1254), .A2(n1253), .ZN(n1255) );
XNOR2_X1 U964 ( .A(n1256), .B(G140), .ZN(n1253) );
NAND2_X1 U965 ( .A1(KEYINPUT15), .A2(n1126), .ZN(n1256) );
INV_X1 U966 ( .A(KEYINPUT35), .ZN(n1254) );
XOR2_X1 U967 ( .A(KEYINPUT11), .B(G469), .Z(n1228) );
NAND2_X1 U968 ( .A1(G221), .A2(n1197), .ZN(n1021) );
NAND2_X1 U969 ( .A1(G234), .A2(n1198), .ZN(n1197) );
NAND2_X1 U970 ( .A1(n1006), .A2(n1257), .ZN(n1193) );
NAND4_X1 U971 ( .A1(G902), .A2(n1258), .A3(n1182), .A4(n1259), .ZN(n1257) );
INV_X1 U972 ( .A(G898), .ZN(n1259) );
XNOR2_X1 U973 ( .A(KEYINPUT33), .B(n1081), .ZN(n1258) );
INV_X1 U974 ( .A(n1059), .ZN(n1081) );
XOR2_X1 U975 ( .A(G953), .B(KEYINPUT56), .Z(n1059) );
NAND3_X1 U976 ( .A1(n1182), .A2(n1161), .A3(G952), .ZN(n1006) );
NAND2_X1 U977 ( .A1(G237), .A2(G234), .ZN(n1182) );
XNOR2_X1 U978 ( .A(n1032), .B(KEYINPUT31), .ZN(n1190) );
AND2_X1 U979 ( .A1(n1033), .A2(n1260), .ZN(n1032) );
NAND2_X1 U980 ( .A1(n1036), .A2(n1050), .ZN(n1260) );
NAND3_X1 U981 ( .A1(n1261), .A2(n1198), .A3(n1262), .ZN(n1050) );
XNOR2_X1 U982 ( .A(n1048), .B(KEYINPUT44), .ZN(n1036) );
NAND2_X1 U983 ( .A1(n1263), .A2(n1264), .ZN(n1048) );
NAND2_X1 U984 ( .A1(n1262), .A2(n1198), .ZN(n1264) );
XOR2_X1 U985 ( .A(n1265), .B(n1266), .Z(n1262) );
XOR2_X1 U986 ( .A(n1267), .B(n1160), .Z(n1266) );
XNOR2_X1 U987 ( .A(n1216), .B(n1268), .ZN(n1160) );
AND2_X1 U988 ( .A1(n1161), .A2(G224), .ZN(n1268) );
XOR2_X1 U989 ( .A(n1269), .B(n1270), .Z(n1216) );
XOR2_X1 U990 ( .A(KEYINPUT54), .B(KEYINPUT13), .Z(n1270) );
XNOR2_X1 U991 ( .A(G146), .B(n1271), .ZN(n1269) );
NAND2_X1 U992 ( .A1(KEYINPUT3), .A2(n1159), .ZN(n1267) );
XNOR2_X1 U993 ( .A(n1082), .B(KEYINPUT0), .ZN(n1159) );
XOR2_X1 U994 ( .A(n1272), .B(n1273), .Z(n1082) );
XOR2_X1 U995 ( .A(G104), .B(n1274), .Z(n1273) );
XNOR2_X1 U996 ( .A(G122), .B(n1126), .ZN(n1274) );
INV_X1 U997 ( .A(G110), .ZN(n1126) );
XNOR2_X1 U998 ( .A(n1114), .B(n1275), .ZN(n1272) );
NOR2_X1 U999 ( .A1(G107), .A2(KEYINPUT7), .ZN(n1275) );
XNOR2_X1 U1000 ( .A(n1213), .B(n1276), .ZN(n1114) );
INV_X1 U1001 ( .A(n1225), .ZN(n1276) );
XOR2_X1 U1002 ( .A(G101), .B(KEYINPUT26), .Z(n1225) );
XOR2_X1 U1003 ( .A(G113), .B(n1277), .Z(n1213) );
XOR2_X1 U1004 ( .A(G119), .B(G116), .Z(n1277) );
XNOR2_X1 U1005 ( .A(n1278), .B(n1134), .ZN(n1265) );
XNOR2_X1 U1006 ( .A(KEYINPUT58), .B(KEYINPUT34), .ZN(n1278) );
INV_X1 U1007 ( .A(n1261), .ZN(n1263) );
NAND2_X1 U1008 ( .A1(G210), .A2(n1279), .ZN(n1261) );
XOR2_X1 U1009 ( .A(KEYINPUT62), .B(n1280), .Z(n1279) );
NOR2_X1 U1010 ( .A1(G237), .A2(G902), .ZN(n1280) );
NAND2_X1 U1011 ( .A1(G214), .A2(n1281), .ZN(n1033) );
NAND2_X1 U1012 ( .A1(n1226), .A2(n1198), .ZN(n1281) );
INV_X1 U1013 ( .A(n1173), .ZN(n1010) );
NOR2_X1 U1014 ( .A1(n1185), .A2(n1184), .ZN(n1173) );
XOR2_X1 U1015 ( .A(G475), .B(n1282), .Z(n1184) );
NOR2_X1 U1016 ( .A1(G902), .A2(n1098), .ZN(n1282) );
XNOR2_X1 U1017 ( .A(n1283), .B(n1284), .ZN(n1098) );
XNOR2_X1 U1018 ( .A(G104), .B(n1285), .ZN(n1284) );
NAND2_X1 U1019 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U1020 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U1021 ( .A1(KEYINPUT5), .A2(n1290), .ZN(n1289) );
NAND2_X1 U1022 ( .A1(KEYINPUT52), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U1023 ( .A(n1065), .B(n1292), .ZN(n1291) );
INV_X1 U1024 ( .A(G131), .ZN(n1065) );
XNOR2_X1 U1025 ( .A(n1293), .B(n1066), .ZN(n1288) );
NAND2_X1 U1026 ( .A1(n1294), .A2(n1295), .ZN(n1286) );
NAND2_X1 U1027 ( .A1(KEYINPUT52), .A2(n1296), .ZN(n1295) );
NAND2_X1 U1028 ( .A1(KEYINPUT5), .A2(n1297), .ZN(n1296) );
XOR2_X1 U1029 ( .A(n1293), .B(n1066), .Z(n1297) );
XNOR2_X1 U1030 ( .A(n1134), .B(G140), .ZN(n1066) );
INV_X1 U1031 ( .A(G125), .ZN(n1134) );
NOR2_X1 U1032 ( .A1(G146), .A2(KEYINPUT53), .ZN(n1293) );
XNOR2_X1 U1033 ( .A(G131), .B(n1292), .ZN(n1294) );
NOR3_X1 U1034 ( .A1(n1298), .A2(n1299), .A3(KEYINPUT32), .ZN(n1292) );
NOR2_X1 U1035 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
XNOR2_X1 U1036 ( .A(KEYINPUT51), .B(n1168), .ZN(n1301) );
INV_X1 U1037 ( .A(n1302), .ZN(n1300) );
NOR2_X1 U1038 ( .A1(G143), .A2(n1302), .ZN(n1298) );
NAND3_X1 U1039 ( .A1(n1226), .A2(n1161), .A3(G214), .ZN(n1302) );
INV_X1 U1040 ( .A(G237), .ZN(n1226) );
XNOR2_X1 U1041 ( .A(G113), .B(G122), .ZN(n1283) );
XNOR2_X1 U1042 ( .A(n1303), .B(G478), .ZN(n1185) );
NAND2_X1 U1043 ( .A1(n1304), .A2(n1198), .ZN(n1303) );
INV_X1 U1044 ( .A(G902), .ZN(n1198) );
XNOR2_X1 U1045 ( .A(n1092), .B(KEYINPUT6), .ZN(n1304) );
AND2_X1 U1046 ( .A1(n1305), .A2(n1306), .ZN(n1092) );
NAND2_X1 U1047 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1048 ( .A1(G217), .A2(n1206), .ZN(n1308) );
NAND3_X1 U1049 ( .A1(G217), .A2(n1206), .A3(n1309), .ZN(n1305) );
INV_X1 U1050 ( .A(n1307), .ZN(n1309) );
XNOR2_X1 U1051 ( .A(n1310), .B(n1311), .ZN(n1307) );
XOR2_X1 U1052 ( .A(G116), .B(n1312), .Z(n1311) );
XNOR2_X1 U1053 ( .A(n1250), .B(G122), .ZN(n1312) );
INV_X1 U1054 ( .A(G134), .ZN(n1250) );
XNOR2_X1 U1055 ( .A(G107), .B(n1271), .ZN(n1310) );
XNOR2_X1 U1056 ( .A(G128), .B(n1168), .ZN(n1271) );
INV_X1 U1057 ( .A(G143), .ZN(n1168) );
AND2_X1 U1058 ( .A1(G234), .A2(n1161), .ZN(n1206) );
INV_X1 U1059 ( .A(G953), .ZN(n1161) );
endmodule


