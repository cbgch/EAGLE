//Key = 1100111110111100001000100011001010100110100101001001101111010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328;

NAND2_X1 U738 ( .A1(n1017), .A2(n1018), .ZN(G9) );
NAND2_X1 U739 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
XOR2_X1 U740 ( .A(KEYINPUT37), .B(n1021), .Z(n1017) );
NOR2_X1 U741 ( .A1(n1019), .A2(n1020), .ZN(n1021) );
NOR2_X1 U742 ( .A1(n1022), .A2(n1023), .ZN(G75) );
XOR2_X1 U743 ( .A(n1024), .B(KEYINPUT18), .Z(n1023) );
OR3_X1 U744 ( .A1(G952), .A2(G953), .A3(n1025), .ZN(n1024) );
NOR4_X1 U745 ( .A1(n1026), .A2(n1027), .A3(G953), .A4(n1025), .ZN(n1022) );
AND4_X1 U746 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1025) );
NOR4_X1 U747 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
XOR2_X1 U748 ( .A(n1036), .B(n1037), .Z(n1034) );
XNOR2_X1 U749 ( .A(n1038), .B(KEYINPUT32), .ZN(n1037) );
NAND2_X1 U750 ( .A1(KEYINPUT10), .A2(n1039), .ZN(n1038) );
XNOR2_X1 U751 ( .A(n1040), .B(n1041), .ZN(n1033) );
NAND2_X1 U752 ( .A1(KEYINPUT0), .A2(n1042), .ZN(n1040) );
XNOR2_X1 U753 ( .A(n1043), .B(n1044), .ZN(n1030) );
NAND2_X1 U754 ( .A1(KEYINPUT43), .A2(n1045), .ZN(n1043) );
INV_X1 U755 ( .A(n1046), .ZN(n1045) );
XOR2_X1 U756 ( .A(n1047), .B(KEYINPUT16), .Z(n1028) );
NOR2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1027) );
NOR2_X1 U758 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR3_X1 U759 ( .A1(n1035), .A2(n1052), .A3(n1053), .ZN(n1051) );
NOR2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR3_X1 U762 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1056) );
NOR3_X1 U763 ( .A1(n1047), .A2(n1061), .A3(n1062), .ZN(n1060) );
INV_X1 U764 ( .A(n1063), .ZN(n1061) );
NOR2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U767 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR3_X1 U768 ( .A1(n1065), .A2(n1070), .A3(n1062), .ZN(n1054) );
NOR2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR4_X1 U770 ( .A1(n1073), .A2(n1062), .A3(n1057), .A4(n1065), .ZN(n1050) );
NOR2_X1 U771 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U772 ( .A1(n1076), .A2(G952), .A3(n1077), .ZN(n1026) );
XOR2_X1 U773 ( .A(n1078), .B(n1079), .Z(G72) );
XOR2_X1 U774 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XOR2_X1 U776 ( .A(n1084), .B(n1085), .Z(n1083) );
XOR2_X1 U777 ( .A(n1086), .B(n1087), .Z(n1085) );
XNOR2_X1 U778 ( .A(n1088), .B(KEYINPUT14), .ZN(n1084) );
NAND2_X1 U779 ( .A1(KEYINPUT51), .A2(n1089), .ZN(n1088) );
XNOR2_X1 U780 ( .A(n1090), .B(KEYINPUT45), .ZN(n1082) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1080) );
XNOR2_X1 U782 ( .A(G953), .B(n1093), .ZN(n1091) );
XNOR2_X1 U783 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n1093) );
NAND2_X1 U784 ( .A1(G953), .A2(n1094), .ZN(n1078) );
NAND2_X1 U785 ( .A1(G900), .A2(G227), .ZN(n1094) );
NAND2_X1 U786 ( .A1(n1095), .A2(n1096), .ZN(G69) );
NAND2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U788 ( .A(n1099), .B(n1077), .Z(n1097) );
NAND2_X1 U789 ( .A1(n1100), .A2(G953), .ZN(n1095) );
NAND2_X1 U790 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U791 ( .A1(n1099), .A2(n1103), .ZN(n1102) );
INV_X1 U792 ( .A(G224), .ZN(n1103) );
NAND2_X1 U793 ( .A1(G224), .A2(n1104), .ZN(n1101) );
NAND2_X1 U794 ( .A1(G898), .A2(n1099), .ZN(n1104) );
NAND2_X1 U795 ( .A1(n1105), .A2(n1106), .ZN(n1099) );
NAND2_X1 U796 ( .A1(G953), .A2(n1107), .ZN(n1106) );
XNOR2_X1 U797 ( .A(n1108), .B(n1109), .ZN(n1105) );
NOR2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(G66) );
XOR2_X1 U799 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U800 ( .A(KEYINPUT40), .B(n1114), .Z(n1113) );
NOR2_X1 U801 ( .A1(n1046), .A2(n1115), .ZN(n1114) );
NOR2_X1 U802 ( .A1(n1110), .A2(n1116), .ZN(G63) );
XOR2_X1 U803 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U804 ( .A1(n1119), .A2(n1115), .ZN(n1117) );
NOR2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(G60) );
XNOR2_X1 U806 ( .A(n1110), .B(KEYINPUT12), .ZN(n1121) );
XNOR2_X1 U807 ( .A(n1122), .B(n1123), .ZN(n1120) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1115), .ZN(n1123) );
XNOR2_X1 U809 ( .A(G104), .B(n1125), .ZN(G6) );
NOR2_X1 U810 ( .A1(n1110), .A2(n1126), .ZN(G57) );
XOR2_X1 U811 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U812 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U813 ( .A(G101), .B(n1131), .ZN(n1130) );
NOR2_X1 U814 ( .A1(KEYINPUT19), .A2(n1132), .ZN(n1129) );
XOR2_X1 U815 ( .A(n1133), .B(n1134), .Z(n1127) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1115), .ZN(n1134) );
NOR2_X1 U817 ( .A1(n1110), .A2(n1136), .ZN(G54) );
XOR2_X1 U818 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U819 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
OR2_X1 U820 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U821 ( .A(n1143), .B(KEYINPUT50), .Z(n1139) );
NAND2_X1 U822 ( .A1(n1142), .A2(n1141), .ZN(n1143) );
XNOR2_X1 U823 ( .A(n1144), .B(n1145), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1146), .B(n1087), .Z(n1142) );
NAND3_X1 U825 ( .A1(n1147), .A2(n1148), .A3(G469), .ZN(n1137) );
NAND2_X1 U826 ( .A1(n1115), .A2(n1149), .ZN(n1148) );
INV_X1 U827 ( .A(KEYINPUT33), .ZN(n1149) );
NAND2_X1 U828 ( .A1(KEYINPUT33), .A2(n1150), .ZN(n1147) );
NAND2_X1 U829 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U830 ( .A1(n1153), .A2(n1154), .ZN(G51) );
XNOR2_X1 U831 ( .A(n1110), .B(KEYINPUT5), .ZN(n1154) );
NOR2_X1 U832 ( .A1(n1098), .A2(G952), .ZN(n1110) );
XOR2_X1 U833 ( .A(n1155), .B(n1156), .Z(n1153) );
XOR2_X1 U834 ( .A(n1157), .B(n1158), .Z(n1155) );
NOR2_X1 U835 ( .A1(n1041), .A2(n1115), .ZN(n1158) );
NAND2_X1 U836 ( .A1(G902), .A2(n1152), .ZN(n1115) );
NAND2_X1 U837 ( .A1(n1077), .A2(n1076), .ZN(n1152) );
INV_X1 U838 ( .A(n1092), .ZN(n1076) );
NAND4_X1 U839 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1092) );
NOR4_X1 U840 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
NOR2_X1 U841 ( .A1(n1065), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U842 ( .A(KEYINPUT57), .B(n1168), .ZN(n1167) );
NOR4_X1 U843 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1164) );
INV_X1 U844 ( .A(KEYINPUT31), .ZN(n1170) );
NOR2_X1 U845 ( .A1(n1173), .A2(n1174), .ZN(n1163) );
NOR2_X1 U846 ( .A1(n1175), .A2(n1176), .ZN(n1173) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1172), .ZN(n1176) );
NOR2_X1 U848 ( .A1(n1178), .A2(n1072), .ZN(n1177) );
NOR2_X1 U849 ( .A1(KEYINPUT31), .A2(n1171), .ZN(n1178) );
NOR2_X1 U850 ( .A1(n1179), .A2(n1180), .ZN(n1175) );
AND4_X1 U851 ( .A1(n1181), .A2(n1125), .A3(n1182), .A4(n1183), .ZN(n1077) );
NOR4_X1 U852 ( .A1(n1019), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1183) );
INV_X1 U853 ( .A(n1187), .ZN(n1186) );
AND2_X1 U854 ( .A1(n1071), .A2(n1188), .ZN(n1019) );
NAND2_X1 U855 ( .A1(n1169), .A2(n1189), .ZN(n1182) );
NAND2_X1 U856 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND4_X1 U857 ( .A1(n1072), .A2(n1074), .A3(n1192), .A4(n1193), .ZN(n1191) );
XNOR2_X1 U858 ( .A(KEYINPUT22), .B(n1194), .ZN(n1190) );
NAND2_X1 U859 ( .A1(n1072), .A2(n1188), .ZN(n1125) );
AND3_X1 U860 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1188) );
NAND3_X1 U861 ( .A1(n1029), .A2(n1197), .A3(n1075), .ZN(n1181) );
NAND3_X1 U862 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(n1157) );
XNOR2_X1 U863 ( .A(n1201), .B(KEYINPUT3), .ZN(n1200) );
OR3_X1 U864 ( .A1(n1202), .A2(n1203), .A3(KEYINPUT52), .ZN(n1199) );
NAND2_X1 U865 ( .A1(n1204), .A2(KEYINPUT52), .ZN(n1198) );
XNOR2_X1 U866 ( .A(G146), .B(n1205), .ZN(G48) );
NAND2_X1 U867 ( .A1(n1169), .A2(n1206), .ZN(n1205) );
XOR2_X1 U868 ( .A(KEYINPUT17), .B(n1207), .Z(n1206) );
NOR2_X1 U869 ( .A1(n1208), .A2(n1172), .ZN(n1207) );
XNOR2_X1 U870 ( .A(n1209), .B(n1210), .ZN(G45) );
NOR3_X1 U871 ( .A1(n1211), .A2(n1174), .A3(n1180), .ZN(n1210) );
NAND4_X1 U872 ( .A1(n1074), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1180) );
XNOR2_X1 U873 ( .A(KEYINPUT4), .B(n1179), .ZN(n1211) );
XNOR2_X1 U874 ( .A(G140), .B(n1161), .ZN(G42) );
NAND2_X1 U875 ( .A1(n1215), .A2(n1075), .ZN(n1161) );
XNOR2_X1 U876 ( .A(G137), .B(n1159), .ZN(G39) );
OR3_X1 U877 ( .A1(n1065), .A2(n1057), .A3(n1172), .ZN(n1159) );
XNOR2_X1 U878 ( .A(n1216), .B(n1217), .ZN(G36) );
NOR2_X1 U879 ( .A1(n1065), .A2(n1168), .ZN(n1217) );
NAND4_X1 U880 ( .A1(n1074), .A2(n1071), .A3(n1067), .A4(n1214), .ZN(n1168) );
XNOR2_X1 U881 ( .A(G131), .B(n1218), .ZN(G33) );
NAND2_X1 U882 ( .A1(KEYINPUT34), .A2(n1166), .ZN(n1218) );
AND2_X1 U883 ( .A1(n1215), .A2(n1074), .ZN(n1166) );
NOR4_X1 U884 ( .A1(n1065), .A2(n1208), .A3(n1179), .A4(n1219), .ZN(n1215) );
INV_X1 U885 ( .A(n1214), .ZN(n1219) );
NAND2_X1 U886 ( .A1(n1063), .A2(n1047), .ZN(n1065) );
XNOR2_X1 U887 ( .A(n1220), .B(KEYINPUT39), .ZN(n1063) );
XNOR2_X1 U888 ( .A(n1221), .B(n1222), .ZN(G30) );
NOR3_X1 U889 ( .A1(n1172), .A2(n1174), .A3(n1171), .ZN(n1222) );
INV_X1 U890 ( .A(n1071), .ZN(n1171) );
NAND4_X1 U891 ( .A1(n1053), .A2(n1067), .A3(n1035), .A4(n1214), .ZN(n1172) );
XNOR2_X1 U892 ( .A(G101), .B(n1187), .ZN(G3) );
NAND3_X1 U893 ( .A1(n1029), .A2(n1197), .A3(n1074), .ZN(n1187) );
XNOR2_X1 U894 ( .A(G125), .B(n1160), .ZN(G27) );
NAND4_X1 U895 ( .A1(n1075), .A2(n1072), .A3(n1059), .A4(n1214), .ZN(n1160) );
NAND2_X1 U896 ( .A1(n1049), .A2(n1223), .ZN(n1214) );
NAND3_X1 U897 ( .A1(G902), .A2(n1224), .A3(n1090), .ZN(n1223) );
NOR2_X1 U898 ( .A1(n1098), .A2(G900), .ZN(n1090) );
XNOR2_X1 U899 ( .A(n1225), .B(n1185), .ZN(G24) );
AND4_X1 U900 ( .A1(n1212), .A2(n1213), .A3(n1196), .A4(n1226), .ZN(n1185) );
NOR2_X1 U901 ( .A1(n1227), .A2(n1035), .ZN(n1226) );
XNOR2_X1 U902 ( .A(n1228), .B(n1184), .ZN(G21) );
NOR4_X1 U903 ( .A1(n1057), .A2(n1227), .A3(n1196), .A4(n1195), .ZN(n1184) );
INV_X1 U904 ( .A(n1035), .ZN(n1195) );
NAND2_X1 U905 ( .A1(n1059), .A2(n1193), .ZN(n1227) );
XOR2_X1 U906 ( .A(G116), .B(n1229), .Z(G18) );
NOR2_X1 U907 ( .A1(n1174), .A2(n1194), .ZN(n1229) );
NAND4_X1 U908 ( .A1(n1074), .A2(n1192), .A3(n1071), .A4(n1193), .ZN(n1194) );
NOR2_X1 U909 ( .A1(n1213), .A2(n1230), .ZN(n1071) );
XNOR2_X1 U910 ( .A(G113), .B(n1231), .ZN(G15) );
NAND4_X1 U911 ( .A1(n1072), .A2(n1074), .A3(n1059), .A4(n1232), .ZN(n1231) );
XNOR2_X1 U912 ( .A(KEYINPUT13), .B(n1193), .ZN(n1232) );
NOR2_X1 U913 ( .A1(n1062), .A2(n1174), .ZN(n1059) );
INV_X1 U914 ( .A(n1192), .ZN(n1062) );
NOR2_X1 U915 ( .A1(n1068), .A2(n1032), .ZN(n1192) );
INV_X1 U916 ( .A(n1069), .ZN(n1032) );
AND2_X1 U917 ( .A1(n1233), .A2(n1035), .ZN(n1074) );
XNOR2_X1 U918 ( .A(KEYINPUT49), .B(n1053), .ZN(n1233) );
INV_X1 U919 ( .A(n1196), .ZN(n1053) );
INV_X1 U920 ( .A(n1208), .ZN(n1072) );
NAND2_X1 U921 ( .A1(n1230), .A2(n1213), .ZN(n1208) );
INV_X1 U922 ( .A(n1212), .ZN(n1230) );
XNOR2_X1 U923 ( .A(G110), .B(n1234), .ZN(G12) );
NAND3_X1 U924 ( .A1(n1197), .A2(n1235), .A3(n1075), .ZN(n1234) );
NOR2_X1 U925 ( .A1(n1196), .A2(n1035), .ZN(n1075) );
XOR2_X1 U926 ( .A(n1236), .B(n1135), .Z(n1035) );
INV_X1 U927 ( .A(G472), .ZN(n1135) );
NAND2_X1 U928 ( .A1(n1237), .A2(n1151), .ZN(n1236) );
XOR2_X1 U929 ( .A(n1133), .B(n1238), .Z(n1237) );
XOR2_X1 U930 ( .A(n1132), .B(n1239), .Z(n1238) );
NOR2_X1 U931 ( .A1(KEYINPUT28), .A2(n1240), .ZN(n1239) );
XOR2_X1 U932 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U933 ( .A(n1131), .B(KEYINPUT15), .Z(n1242) );
NAND2_X1 U934 ( .A1(G210), .A2(n1243), .ZN(n1131) );
NAND2_X1 U935 ( .A1(KEYINPUT38), .A2(n1244), .ZN(n1241) );
XOR2_X1 U936 ( .A(n1245), .B(n1246), .Z(n1132) );
XNOR2_X1 U937 ( .A(G116), .B(KEYINPUT61), .ZN(n1245) );
XNOR2_X1 U938 ( .A(n1247), .B(n1087), .ZN(n1133) );
XOR2_X1 U939 ( .A(n1248), .B(n1046), .Z(n1196) );
NAND2_X1 U940 ( .A1(G217), .A2(n1249), .ZN(n1046) );
XOR2_X1 U941 ( .A(n1044), .B(KEYINPUT62), .Z(n1248) );
NAND2_X1 U942 ( .A1(n1112), .A2(n1151), .ZN(n1044) );
XOR2_X1 U943 ( .A(n1250), .B(n1251), .Z(n1112) );
XOR2_X1 U944 ( .A(n1086), .B(n1252), .Z(n1251) );
NOR2_X1 U945 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
NOR2_X1 U946 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XNOR2_X1 U947 ( .A(G110), .B(KEYINPUT6), .ZN(n1256) );
INV_X1 U948 ( .A(n1257), .ZN(n1255) );
NOR2_X1 U949 ( .A1(n1257), .A2(n1258), .ZN(n1253) );
XNOR2_X1 U950 ( .A(KEYINPUT54), .B(n1145), .ZN(n1258) );
XNOR2_X1 U951 ( .A(G119), .B(n1221), .ZN(n1257) );
XOR2_X1 U952 ( .A(n1259), .B(n1260), .Z(n1250) );
XNOR2_X1 U953 ( .A(n1261), .B(G137), .ZN(n1260) );
NAND3_X1 U954 ( .A1(G234), .A2(n1098), .A3(G221), .ZN(n1259) );
XNOR2_X1 U955 ( .A(KEYINPUT25), .B(n1057), .ZN(n1235) );
INV_X1 U956 ( .A(n1029), .ZN(n1057) );
NOR2_X1 U957 ( .A1(n1212), .A2(n1213), .ZN(n1029) );
XOR2_X1 U958 ( .A(n1262), .B(n1124), .Z(n1213) );
INV_X1 U959 ( .A(G475), .ZN(n1124) );
NAND2_X1 U960 ( .A1(n1122), .A2(n1151), .ZN(n1262) );
XNOR2_X1 U961 ( .A(n1263), .B(n1264), .ZN(n1122) );
XOR2_X1 U962 ( .A(G104), .B(n1265), .Z(n1264) );
XNOR2_X1 U963 ( .A(n1225), .B(G113), .ZN(n1265) );
XOR2_X1 U964 ( .A(n1266), .B(n1267), .Z(n1263) );
NOR2_X1 U965 ( .A1(KEYINPUT21), .A2(n1268), .ZN(n1267) );
XOR2_X1 U966 ( .A(n1269), .B(n1270), .Z(n1268) );
XNOR2_X1 U967 ( .A(n1271), .B(n1209), .ZN(n1269) );
INV_X1 U968 ( .A(G143), .ZN(n1209) );
NAND2_X1 U969 ( .A1(G214), .A2(n1243), .ZN(n1271) );
NOR2_X1 U970 ( .A1(G953), .A2(G237), .ZN(n1243) );
NAND2_X1 U971 ( .A1(n1272), .A2(n1273), .ZN(n1266) );
NAND2_X1 U972 ( .A1(G146), .A2(n1086), .ZN(n1273) );
XOR2_X1 U973 ( .A(n1274), .B(KEYINPUT9), .Z(n1272) );
OR2_X1 U974 ( .A1(n1086), .A2(G146), .ZN(n1274) );
XOR2_X1 U975 ( .A(G125), .B(n1275), .Z(n1086) );
XOR2_X1 U976 ( .A(n1276), .B(n1119), .Z(n1212) );
INV_X1 U977 ( .A(G478), .ZN(n1119) );
OR2_X1 U978 ( .A1(n1118), .A2(G902), .ZN(n1276) );
XNOR2_X1 U979 ( .A(n1277), .B(n1278), .ZN(n1118) );
NOR2_X1 U980 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XOR2_X1 U981 ( .A(n1281), .B(KEYINPUT27), .Z(n1280) );
NAND2_X1 U982 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NOR2_X1 U983 ( .A1(n1282), .A2(n1284), .ZN(n1279) );
XOR2_X1 U984 ( .A(n1283), .B(KEYINPUT36), .Z(n1284) );
XNOR2_X1 U985 ( .A(G107), .B(n1285), .ZN(n1283) );
XNOR2_X1 U986 ( .A(n1225), .B(G116), .ZN(n1285) );
INV_X1 U987 ( .A(G122), .ZN(n1225) );
XOR2_X1 U988 ( .A(n1286), .B(n1287), .Z(n1282) );
NAND2_X1 U989 ( .A1(KEYINPUT30), .A2(n1216), .ZN(n1286) );
INV_X1 U990 ( .A(G134), .ZN(n1216) );
NAND4_X1 U991 ( .A1(G234), .A2(G217), .A3(n1288), .A4(n1098), .ZN(n1277) );
XOR2_X1 U992 ( .A(KEYINPUT7), .B(KEYINPUT42), .Z(n1288) );
AND3_X1 U993 ( .A1(n1169), .A2(n1193), .A3(n1067), .ZN(n1197) );
INV_X1 U994 ( .A(n1179), .ZN(n1067) );
NAND2_X1 U995 ( .A1(n1068), .A2(n1069), .ZN(n1179) );
NAND2_X1 U996 ( .A1(G221), .A2(n1249), .ZN(n1069) );
NAND2_X1 U997 ( .A1(n1289), .A2(n1151), .ZN(n1249) );
NAND2_X1 U998 ( .A1(n1290), .A2(n1291), .ZN(n1068) );
NAND2_X1 U999 ( .A1(n1039), .A2(n1036), .ZN(n1291) );
XOR2_X1 U1000 ( .A(KEYINPUT59), .B(n1292), .Z(n1290) );
NOR2_X1 U1001 ( .A1(n1039), .A2(n1036), .ZN(n1292) );
XNOR2_X1 U1002 ( .A(G469), .B(KEYINPUT60), .ZN(n1036) );
AND2_X1 U1003 ( .A1(n1293), .A2(n1151), .ZN(n1039) );
XOR2_X1 U1004 ( .A(n1294), .B(n1295), .Z(n1293) );
NOR2_X1 U1005 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U1006 ( .A(KEYINPUT24), .B(n1298), .Z(n1297) );
AND2_X1 U1007 ( .A1(n1299), .A2(n1146), .ZN(n1298) );
NOR2_X1 U1008 ( .A1(n1146), .A2(n1299), .ZN(n1296) );
XOR2_X1 U1009 ( .A(n1087), .B(KEYINPUT55), .Z(n1299) );
XNOR2_X1 U1010 ( .A(n1300), .B(n1270), .ZN(n1087) );
XOR2_X1 U1011 ( .A(G131), .B(KEYINPUT20), .Z(n1270) );
XNOR2_X1 U1012 ( .A(G134), .B(G137), .ZN(n1300) );
XNOR2_X1 U1013 ( .A(n1301), .B(n1089), .ZN(n1146) );
AND2_X1 U1014 ( .A1(n1302), .A2(n1303), .ZN(n1089) );
NAND2_X1 U1015 ( .A1(n1287), .A2(G146), .ZN(n1303) );
NAND2_X1 U1016 ( .A1(n1304), .A2(n1261), .ZN(n1302) );
INV_X1 U1017 ( .A(G146), .ZN(n1261) );
XNOR2_X1 U1018 ( .A(n1287), .B(KEYINPUT23), .ZN(n1304) );
XOR2_X1 U1019 ( .A(G128), .B(G143), .Z(n1287) );
XNOR2_X1 U1020 ( .A(n1305), .B(n1244), .ZN(n1301) );
INV_X1 U1021 ( .A(G101), .ZN(n1244) );
NAND2_X1 U1022 ( .A1(KEYINPUT1), .A2(n1306), .ZN(n1294) );
XNOR2_X1 U1023 ( .A(n1307), .B(n1308), .ZN(n1306) );
INV_X1 U1024 ( .A(n1144), .ZN(n1308) );
XNOR2_X1 U1025 ( .A(n1309), .B(n1275), .ZN(n1144) );
XOR2_X1 U1026 ( .A(G140), .B(KEYINPUT47), .Z(n1275) );
NAND2_X1 U1027 ( .A1(G227), .A2(n1098), .ZN(n1309) );
NOR2_X1 U1028 ( .A1(G110), .A2(KEYINPUT2), .ZN(n1307) );
NAND2_X1 U1029 ( .A1(n1049), .A2(n1310), .ZN(n1193) );
NAND4_X1 U1030 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1107), .ZN(n1310) );
INV_X1 U1031 ( .A(G898), .ZN(n1107) );
NAND3_X1 U1032 ( .A1(n1224), .A2(n1098), .A3(G952), .ZN(n1049) );
NAND2_X1 U1033 ( .A1(G237), .A2(n1289), .ZN(n1224) );
XNOR2_X1 U1034 ( .A(G234), .B(KEYINPUT26), .ZN(n1289) );
INV_X1 U1035 ( .A(n1174), .ZN(n1169) );
NAND2_X1 U1036 ( .A1(n1220), .A2(n1047), .ZN(n1174) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1311), .ZN(n1047) );
XNOR2_X1 U1038 ( .A(n1312), .B(n1041), .ZN(n1220) );
NAND2_X1 U1039 ( .A1(G210), .A2(n1311), .ZN(n1041) );
NAND2_X1 U1040 ( .A1(n1313), .A2(n1151), .ZN(n1311) );
INV_X1 U1041 ( .A(G237), .ZN(n1313) );
XOR2_X1 U1042 ( .A(n1042), .B(KEYINPUT56), .Z(n1312) );
NAND2_X1 U1043 ( .A1(n1314), .A2(n1151), .ZN(n1042) );
INV_X1 U1044 ( .A(G902), .ZN(n1151) );
XOR2_X1 U1045 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1046 ( .A(n1156), .B(n1317), .ZN(n1316) );
NOR2_X1 U1047 ( .A1(n1204), .A2(n1201), .ZN(n1317) );
AND2_X1 U1048 ( .A1(n1318), .A2(n1203), .ZN(n1201) );
NOR2_X1 U1049 ( .A1(n1203), .A2(n1318), .ZN(n1204) );
INV_X1 U1050 ( .A(n1202), .ZN(n1318) );
NAND2_X1 U1051 ( .A1(G224), .A2(n1098), .ZN(n1202) );
INV_X1 U1052 ( .A(G953), .ZN(n1098) );
XNOR2_X1 U1053 ( .A(G125), .B(n1247), .ZN(n1203) );
XNOR2_X1 U1054 ( .A(n1319), .B(n1320), .ZN(n1247) );
NOR2_X1 U1055 ( .A1(KEYINPUT63), .A2(n1221), .ZN(n1320) );
INV_X1 U1056 ( .A(G128), .ZN(n1221) );
XNOR2_X1 U1057 ( .A(G143), .B(G146), .ZN(n1319) );
XOR2_X1 U1058 ( .A(n1108), .B(n1321), .Z(n1156) );
NOR2_X1 U1059 ( .A1(KEYINPUT44), .A2(n1109), .ZN(n1321) );
XOR2_X1 U1060 ( .A(n1322), .B(n1323), .Z(n1109) );
XNOR2_X1 U1061 ( .A(n1324), .B(n1246), .ZN(n1323) );
XNOR2_X1 U1062 ( .A(G113), .B(n1228), .ZN(n1246) );
INV_X1 U1063 ( .A(G119), .ZN(n1228) );
NAND2_X1 U1064 ( .A1(n1325), .A2(KEYINPUT11), .ZN(n1324) );
XOR2_X1 U1065 ( .A(n1305), .B(KEYINPUT58), .Z(n1325) );
XNOR2_X1 U1066 ( .A(G104), .B(n1326), .ZN(n1305) );
XNOR2_X1 U1067 ( .A(KEYINPUT8), .B(n1020), .ZN(n1326) );
INV_X1 U1068 ( .A(G107), .ZN(n1020) );
XOR2_X1 U1069 ( .A(n1327), .B(n1328), .Z(n1322) );
NOR2_X1 U1070 ( .A1(KEYINPUT53), .A2(G116), .ZN(n1328) );
XNOR2_X1 U1071 ( .A(G101), .B(KEYINPUT35), .ZN(n1327) );
XNOR2_X1 U1072 ( .A(G122), .B(n1145), .ZN(n1108) );
INV_X1 U1073 ( .A(G110), .ZN(n1145) );
XNOR2_X1 U1074 ( .A(KEYINPUT41), .B(KEYINPUT29), .ZN(n1315) );
endmodule


