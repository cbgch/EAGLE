//Key = 0011001000010000010100001000111100010110111100101010010001100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
n1456, n1457;

XOR2_X1 U790 ( .A(n1096), .B(n1097), .Z(G9) );
NAND3_X1 U791 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(n1097) );
NAND2_X1 U792 ( .A1(KEYINPUT63), .A2(n1101), .ZN(n1099) );
NAND2_X1 U793 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
INV_X1 U794 ( .A(KEYINPUT63), .ZN(n1103) );
NAND3_X1 U795 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1102) );
INV_X1 U796 ( .A(n1107), .ZN(n1104) );
NOR2_X1 U797 ( .A1(n1108), .A2(n1109), .ZN(G75) );
NOR4_X1 U798 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1109) );
NOR3_X1 U799 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1112) );
NOR2_X1 U800 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U801 ( .A(KEYINPUT1), .B(n1119), .Z(n1118) );
NOR4_X1 U802 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1119) );
NOR2_X1 U803 ( .A1(n1124), .A2(n1123), .ZN(n1117) );
NOR2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U805 ( .A1(n1127), .A2(n1121), .ZN(n1126) );
INV_X1 U806 ( .A(n1128), .ZN(n1121) );
NOR2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
NOR2_X1 U808 ( .A1(n1122), .A2(n1131), .ZN(n1130) );
INV_X1 U809 ( .A(n1132), .ZN(n1122) );
NOR2_X1 U810 ( .A1(n1133), .A2(n1134), .ZN(n1129) );
INV_X1 U811 ( .A(n1106), .ZN(n1134) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NOR2_X1 U813 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1125) );
NAND3_X1 U815 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1110) );
NAND4_X1 U816 ( .A1(n1144), .A2(n1145), .A3(n1128), .A4(n1146), .ZN(n1143) );
NAND2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U818 ( .A1(n1115), .A2(n1149), .ZN(n1148) );
INV_X1 U819 ( .A(n1123), .ZN(n1144) );
NOR3_X1 U820 ( .A1(n1150), .A2(G953), .A3(G952), .ZN(n1108) );
INV_X1 U821 ( .A(n1141), .ZN(n1150) );
NAND4_X1 U822 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1141) );
NOR3_X1 U823 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1154) );
NAND3_X1 U824 ( .A1(n1158), .A2(n1159), .A3(n1149), .ZN(n1155) );
NAND2_X1 U825 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(n1158) );
XOR2_X1 U827 ( .A(KEYINPUT56), .B(n1164), .Z(n1162) );
NOR3_X1 U828 ( .A1(n1165), .A2(n1166), .A3(n1115), .ZN(n1153) );
NAND3_X1 U829 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1152) );
NAND2_X1 U830 ( .A1(G469), .A2(n1170), .ZN(n1169) );
OR2_X1 U831 ( .A1(n1171), .A2(KEYINPUT18), .ZN(n1170) );
OR4_X1 U832 ( .A1(G469), .A2(KEYINPUT18), .A3(n1171), .A4(KEYINPUT15), .ZN(n1168) );
NAND2_X1 U833 ( .A1(n1171), .A2(KEYINPUT15), .ZN(n1167) );
NAND2_X1 U834 ( .A1(n1172), .A2(n1173), .ZN(G72) );
NAND4_X1 U835 ( .A1(G953), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1173) );
XOR2_X1 U836 ( .A(n1177), .B(KEYINPUT16), .Z(n1172) );
NAND2_X1 U837 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U838 ( .A1(G953), .A2(n1174), .ZN(n1179) );
NAND2_X1 U839 ( .A1(G900), .A2(G227), .ZN(n1174) );
NAND2_X1 U840 ( .A1(n1175), .A2(n1176), .ZN(n1178) );
NAND3_X1 U841 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1176) );
XNOR2_X1 U842 ( .A(n1183), .B(n1184), .ZN(n1182) );
NAND2_X1 U843 ( .A1(n1185), .A2(n1186), .ZN(n1181) );
NAND2_X1 U844 ( .A1(G953), .A2(n1187), .ZN(n1180) );
NAND3_X1 U845 ( .A1(n1188), .A2(n1189), .A3(n1185), .ZN(n1175) );
NAND2_X1 U846 ( .A1(n1190), .A2(n1191), .ZN(n1185) );
NAND2_X1 U847 ( .A1(G953), .A2(n1186), .ZN(n1189) );
NAND2_X1 U848 ( .A1(n1192), .A2(n1142), .ZN(n1188) );
NAND2_X1 U849 ( .A1(n1193), .A2(n1186), .ZN(n1192) );
INV_X1 U850 ( .A(KEYINPUT23), .ZN(n1186) );
XOR2_X1 U851 ( .A(n1183), .B(n1184), .Z(n1193) );
NAND2_X1 U852 ( .A1(KEYINPUT41), .A2(n1194), .ZN(n1183) );
XOR2_X1 U853 ( .A(n1195), .B(n1196), .Z(n1194) );
NAND2_X1 U854 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND2_X1 U855 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U856 ( .A(KEYINPUT20), .B(n1201), .Z(n1200) );
XOR2_X1 U857 ( .A(n1202), .B(KEYINPUT54), .Z(n1199) );
NAND2_X1 U858 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
XNOR2_X1 U859 ( .A(KEYINPUT20), .B(n1201), .ZN(n1204) );
XOR2_X1 U860 ( .A(n1202), .B(KEYINPUT11), .Z(n1203) );
INV_X1 U861 ( .A(G131), .ZN(n1202) );
XOR2_X1 U862 ( .A(n1205), .B(n1206), .Z(G69) );
XOR2_X1 U863 ( .A(n1207), .B(n1208), .Z(n1206) );
NAND2_X1 U864 ( .A1(G953), .A2(n1209), .ZN(n1208) );
NAND2_X1 U865 ( .A1(G224), .A2(G898), .ZN(n1209) );
NAND3_X1 U866 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1207) );
NAND2_X1 U867 ( .A1(n1213), .A2(G953), .ZN(n1212) );
NAND2_X1 U868 ( .A1(n1214), .A2(n1215), .ZN(n1211) );
NAND2_X1 U869 ( .A1(n1216), .A2(n1217), .ZN(n1210) );
INV_X1 U870 ( .A(n1215), .ZN(n1217) );
XOR2_X1 U871 ( .A(n1214), .B(KEYINPUT19), .Z(n1216) );
NOR2_X1 U872 ( .A1(n1218), .A2(G953), .ZN(n1205) );
NOR2_X1 U873 ( .A1(n1219), .A2(n1220), .ZN(G66) );
NOR3_X1 U874 ( .A1(n1164), .A2(n1221), .A3(n1222), .ZN(n1220) );
NOR3_X1 U875 ( .A1(n1223), .A2(n1163), .A3(n1224), .ZN(n1222) );
NOR2_X1 U876 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
AND2_X1 U877 ( .A1(n1227), .A2(n1160), .ZN(n1225) );
NOR2_X1 U878 ( .A1(n1219), .A2(n1228), .ZN(G63) );
XNOR2_X1 U879 ( .A(n1229), .B(n1230), .ZN(n1228) );
NOR2_X1 U880 ( .A1(n1231), .A2(n1224), .ZN(n1230) );
INV_X1 U881 ( .A(G478), .ZN(n1231) );
NOR2_X1 U882 ( .A1(n1219), .A2(n1232), .ZN(G60) );
XNOR2_X1 U883 ( .A(n1233), .B(n1234), .ZN(n1232) );
NOR2_X1 U884 ( .A1(n1235), .A2(n1224), .ZN(n1234) );
INV_X1 U885 ( .A(G475), .ZN(n1235) );
XOR2_X1 U886 ( .A(n1236), .B(n1237), .Z(G6) );
OR2_X1 U887 ( .A1(n1101), .A2(n1238), .ZN(n1237) );
NOR2_X1 U888 ( .A1(n1219), .A2(n1239), .ZN(G57) );
XOR2_X1 U889 ( .A(n1240), .B(n1241), .Z(n1239) );
XOR2_X1 U890 ( .A(n1242), .B(n1243), .Z(n1241) );
NAND2_X1 U891 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NAND2_X1 U892 ( .A1(KEYINPUT30), .A2(n1246), .ZN(n1245) );
NAND3_X1 U893 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1244) );
INV_X1 U894 ( .A(KEYINPUT30), .ZN(n1249) );
XOR2_X1 U895 ( .A(n1250), .B(n1251), .Z(n1240) );
NOR2_X1 U896 ( .A1(n1252), .A2(KEYINPUT45), .ZN(n1250) );
NOR2_X1 U897 ( .A1(n1253), .A2(n1224), .ZN(n1252) );
INV_X1 U898 ( .A(G472), .ZN(n1253) );
NOR2_X1 U899 ( .A1(n1219), .A2(n1254), .ZN(G54) );
XOR2_X1 U900 ( .A(n1255), .B(n1256), .Z(n1254) );
NOR2_X1 U901 ( .A1(n1257), .A2(n1224), .ZN(n1256) );
INV_X1 U902 ( .A(G469), .ZN(n1257) );
NAND2_X1 U903 ( .A1(KEYINPUT46), .A2(n1258), .ZN(n1255) );
XOR2_X1 U904 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U905 ( .A(n1261), .B(n1262), .Z(n1260) );
NOR2_X1 U906 ( .A1(n1263), .A2(KEYINPUT7), .ZN(n1262) );
XOR2_X1 U907 ( .A(n1264), .B(n1265), .Z(n1259) );
NOR2_X1 U908 ( .A1(KEYINPUT12), .A2(n1266), .ZN(n1265) );
XOR2_X1 U909 ( .A(n1267), .B(KEYINPUT14), .Z(n1266) );
XOR2_X1 U910 ( .A(n1268), .B(KEYINPUT49), .Z(n1264) );
NOR2_X1 U911 ( .A1(n1219), .A2(n1269), .ZN(G51) );
XOR2_X1 U912 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U913 ( .A(n1272), .B(n1273), .ZN(n1271) );
NAND2_X1 U914 ( .A1(KEYINPUT24), .A2(n1274), .ZN(n1272) );
INV_X1 U915 ( .A(n1275), .ZN(n1274) );
XOR2_X1 U916 ( .A(n1276), .B(n1277), .Z(n1270) );
XOR2_X1 U917 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR2_X1 U918 ( .A1(n1280), .A2(n1224), .ZN(n1279) );
NAND2_X1 U919 ( .A1(G902), .A2(n1227), .ZN(n1224) );
NAND2_X1 U920 ( .A1(n1218), .A2(n1281), .ZN(n1227) );
XNOR2_X1 U921 ( .A(KEYINPUT9), .B(n1113), .ZN(n1281) );
NAND2_X1 U922 ( .A1(n1282), .A2(n1190), .ZN(n1113) );
AND4_X1 U923 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1190) );
NOR4_X1 U924 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1286) );
OR2_X1 U925 ( .A1(n1291), .A2(n1292), .ZN(n1285) );
NAND2_X1 U926 ( .A1(n1293), .A2(n1136), .ZN(n1283) );
INV_X1 U927 ( .A(n1294), .ZN(n1136) );
XOR2_X1 U928 ( .A(n1191), .B(KEYINPUT22), .Z(n1282) );
INV_X1 U929 ( .A(n1111), .ZN(n1218) );
NAND2_X1 U930 ( .A1(n1295), .A2(n1296), .ZN(n1111) );
AND4_X1 U931 ( .A1(n1297), .A2(n1298), .A3(n1299), .A4(n1300), .ZN(n1296) );
NOR4_X1 U932 ( .A1(n1301), .A2(n1302), .A3(n1303), .A4(n1304), .ZN(n1295) );
NOR2_X1 U933 ( .A1(n1139), .A2(n1101), .ZN(n1304) );
NAND2_X1 U934 ( .A1(n1305), .A2(n1106), .ZN(n1101) );
NOR2_X1 U935 ( .A1(n1306), .A2(n1100), .ZN(n1139) );
NOR3_X1 U936 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1303) );
INV_X1 U937 ( .A(n1100), .ZN(n1308) );
XOR2_X1 U938 ( .A(KEYINPUT3), .B(n1310), .Z(n1307) );
AND2_X1 U939 ( .A1(n1311), .A2(KEYINPUT28), .ZN(n1302) );
NOR2_X1 U940 ( .A1(KEYINPUT28), .A2(n1312), .ZN(n1301) );
NAND4_X1 U941 ( .A1(n1145), .A2(n1313), .A3(n1107), .A4(n1147), .ZN(n1312) );
INV_X1 U942 ( .A(n1140), .ZN(n1145) );
NAND2_X1 U943 ( .A1(n1132), .A2(n1106), .ZN(n1140) );
NAND2_X1 U944 ( .A1(KEYINPUT17), .A2(n1247), .ZN(n1276) );
NOR2_X1 U945 ( .A1(n1142), .A2(G952), .ZN(n1219) );
NAND2_X1 U946 ( .A1(n1314), .A2(n1315), .ZN(G48) );
NAND3_X1 U947 ( .A1(n1293), .A2(n1316), .A3(n1317), .ZN(n1315) );
XOR2_X1 U948 ( .A(n1318), .B(KEYINPUT52), .Z(n1314) );
NAND2_X1 U949 ( .A1(G146), .A2(n1319), .ZN(n1318) );
NAND2_X1 U950 ( .A1(n1317), .A2(n1293), .ZN(n1319) );
AND4_X1 U951 ( .A1(n1306), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1293) );
XOR2_X1 U952 ( .A(n1294), .B(KEYINPUT43), .Z(n1317) );
XOR2_X1 U953 ( .A(n1323), .B(n1290), .Z(G45) );
AND4_X1 U954 ( .A1(n1313), .A2(n1310), .A3(n1105), .A4(n1322), .ZN(n1290) );
NAND2_X1 U955 ( .A1(KEYINPUT50), .A2(n1324), .ZN(n1323) );
INV_X1 U956 ( .A(G143), .ZN(n1324) );
XOR2_X1 U957 ( .A(n1289), .B(n1325), .Z(G42) );
NOR2_X1 U958 ( .A1(KEYINPUT21), .A2(n1268), .ZN(n1325) );
INV_X1 U959 ( .A(G140), .ZN(n1268) );
NOR3_X1 U960 ( .A1(n1238), .A2(n1120), .A3(n1292), .ZN(n1289) );
XOR2_X1 U961 ( .A(G137), .B(n1288), .Z(G39) );
AND3_X1 U962 ( .A1(n1128), .A2(n1321), .A3(n1326), .ZN(n1288) );
XOR2_X1 U963 ( .A(n1327), .B(n1328), .Z(G36) );
XOR2_X1 U964 ( .A(KEYINPUT27), .B(G134), .Z(n1328) );
NOR3_X1 U965 ( .A1(n1291), .A2(KEYINPUT5), .A3(n1292), .ZN(n1327) );
XOR2_X1 U966 ( .A(G131), .B(n1287), .Z(G33) );
NOR3_X1 U967 ( .A1(n1238), .A2(n1131), .A3(n1292), .ZN(n1287) );
INV_X1 U968 ( .A(n1326), .ZN(n1292) );
NOR4_X1 U969 ( .A1(n1294), .A2(n1114), .A3(n1329), .A4(n1115), .ZN(n1326) );
XOR2_X1 U970 ( .A(n1149), .B(KEYINPUT42), .Z(n1114) );
NAND2_X1 U971 ( .A1(n1330), .A2(n1331), .ZN(G30) );
NAND2_X1 U972 ( .A1(G128), .A2(n1191), .ZN(n1331) );
XOR2_X1 U973 ( .A(n1332), .B(KEYINPUT26), .Z(n1330) );
OR2_X1 U974 ( .A1(n1191), .A2(G128), .ZN(n1332) );
NAND4_X1 U975 ( .A1(n1100), .A2(n1105), .A3(n1321), .A4(n1322), .ZN(n1191) );
XOR2_X1 U976 ( .A(n1333), .B(n1300), .Z(G3) );
NAND3_X1 U977 ( .A1(n1128), .A2(n1305), .A3(n1310), .ZN(n1300) );
XOR2_X1 U978 ( .A(n1278), .B(n1284), .Z(G27) );
NAND4_X1 U979 ( .A1(n1306), .A2(n1132), .A3(n1334), .A4(n1335), .ZN(n1284) );
NOR2_X1 U980 ( .A1(n1329), .A2(n1147), .ZN(n1334) );
INV_X1 U981 ( .A(n1322), .ZN(n1329) );
NAND2_X1 U982 ( .A1(n1123), .A2(n1336), .ZN(n1322) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1337), .A4(n1187), .ZN(n1336) );
INV_X1 U984 ( .A(G900), .ZN(n1187) );
NAND3_X1 U985 ( .A1(n1338), .A2(n1339), .A3(n1340), .ZN(G24) );
NAND2_X1 U986 ( .A1(G122), .A2(n1341), .ZN(n1340) );
NAND2_X1 U987 ( .A1(KEYINPUT44), .A2(n1342), .ZN(n1339) );
NAND2_X1 U988 ( .A1(n1311), .A2(n1343), .ZN(n1342) );
XOR2_X1 U989 ( .A(KEYINPUT40), .B(G122), .Z(n1343) );
NAND2_X1 U990 ( .A1(n1344), .A2(n1345), .ZN(n1338) );
INV_X1 U991 ( .A(KEYINPUT44), .ZN(n1345) );
NAND2_X1 U992 ( .A1(n1346), .A2(n1347), .ZN(n1344) );
OR2_X1 U993 ( .A1(n1348), .A2(KEYINPUT40), .ZN(n1347) );
NAND3_X1 U994 ( .A1(n1311), .A2(n1348), .A3(KEYINPUT40), .ZN(n1346) );
INV_X1 U995 ( .A(n1341), .ZN(n1311) );
NAND3_X1 U996 ( .A1(n1349), .A2(n1106), .A3(n1313), .ZN(n1341) );
AND2_X1 U997 ( .A1(n1157), .A2(n1350), .ZN(n1313) );
NOR2_X1 U998 ( .A1(n1351), .A2(n1352), .ZN(n1106) );
XNOR2_X1 U999 ( .A(G119), .B(n1299), .ZN(G21) );
NAND3_X1 U1000 ( .A1(n1128), .A2(n1321), .A3(n1349), .ZN(n1299) );
NAND2_X1 U1001 ( .A1(n1353), .A2(n1354), .ZN(n1321) );
OR2_X1 U1002 ( .A1(n1131), .A2(KEYINPUT62), .ZN(n1354) );
INV_X1 U1003 ( .A(n1310), .ZN(n1131) );
NAND3_X1 U1004 ( .A1(n1351), .A2(n1352), .A3(KEYINPUT62), .ZN(n1353) );
INV_X1 U1005 ( .A(n1355), .ZN(n1351) );
XOR2_X1 U1006 ( .A(n1356), .B(n1357), .Z(G18) );
XOR2_X1 U1007 ( .A(KEYINPUT0), .B(G116), .Z(n1357) );
NOR2_X1 U1008 ( .A1(n1309), .A2(n1291), .ZN(n1356) );
NAND2_X1 U1009 ( .A1(n1310), .A2(n1100), .ZN(n1291) );
NOR2_X1 U1010 ( .A1(n1157), .A2(n1358), .ZN(n1100) );
XNOR2_X1 U1011 ( .A(G113), .B(n1298), .ZN(G15) );
NAND3_X1 U1012 ( .A1(n1349), .A2(n1310), .A3(n1306), .ZN(n1298) );
INV_X1 U1013 ( .A(n1238), .ZN(n1306) );
NAND2_X1 U1014 ( .A1(n1358), .A2(n1157), .ZN(n1238) );
INV_X1 U1015 ( .A(n1350), .ZN(n1358) );
NOR2_X1 U1016 ( .A1(n1352), .A2(n1355), .ZN(n1310) );
INV_X1 U1017 ( .A(n1309), .ZN(n1349) );
NAND3_X1 U1018 ( .A1(n1320), .A2(n1107), .A3(n1132), .ZN(n1309) );
NOR2_X1 U1019 ( .A1(n1137), .A2(n1165), .ZN(n1132) );
INV_X1 U1020 ( .A(n1138), .ZN(n1165) );
XOR2_X1 U1021 ( .A(n1267), .B(n1297), .Z(G12) );
NAND3_X1 U1022 ( .A1(n1335), .A2(n1305), .A3(n1128), .ZN(n1297) );
NOR2_X1 U1023 ( .A1(n1350), .A2(n1157), .ZN(n1128) );
XNOR2_X1 U1024 ( .A(n1359), .B(G475), .ZN(n1157) );
NAND2_X1 U1025 ( .A1(n1233), .A2(n1360), .ZN(n1359) );
XNOR2_X1 U1026 ( .A(n1361), .B(n1362), .ZN(n1233) );
XOR2_X1 U1027 ( .A(G122), .B(G104), .Z(n1362) );
XOR2_X1 U1028 ( .A(n1363), .B(n1364), .Z(n1361) );
NOR2_X1 U1029 ( .A1(KEYINPUT59), .A2(n1365), .ZN(n1364) );
XOR2_X1 U1030 ( .A(n1366), .B(n1367), .Z(n1365) );
NAND2_X1 U1031 ( .A1(n1368), .A2(KEYINPUT2), .ZN(n1366) );
XNOR2_X1 U1032 ( .A(n1369), .B(n1370), .ZN(n1368) );
XOR2_X1 U1033 ( .A(n1371), .B(G131), .Z(n1369) );
NAND2_X1 U1034 ( .A1(G214), .A2(n1372), .ZN(n1371) );
NAND2_X1 U1035 ( .A1(n1373), .A2(n1151), .ZN(n1350) );
NAND2_X1 U1036 ( .A1(G478), .A2(n1374), .ZN(n1151) );
XNOR2_X1 U1037 ( .A(n1166), .B(KEYINPUT8), .ZN(n1373) );
NOR2_X1 U1038 ( .A1(n1374), .A2(G478), .ZN(n1166) );
NAND2_X1 U1039 ( .A1(n1229), .A2(n1360), .ZN(n1374) );
XNOR2_X1 U1040 ( .A(n1375), .B(n1376), .ZN(n1229) );
XOR2_X1 U1041 ( .A(G134), .B(n1377), .Z(n1376) );
NOR2_X1 U1042 ( .A1(KEYINPUT13), .A2(n1378), .ZN(n1377) );
XOR2_X1 U1043 ( .A(n1379), .B(n1380), .Z(n1378) );
XOR2_X1 U1044 ( .A(G116), .B(n1348), .Z(n1380) );
INV_X1 U1045 ( .A(G122), .ZN(n1348) );
NAND2_X1 U1046 ( .A1(KEYINPUT37), .A2(n1096), .ZN(n1379) );
XOR2_X1 U1047 ( .A(n1381), .B(n1382), .Z(n1375) );
NOR2_X1 U1048 ( .A1(n1383), .A2(n1384), .ZN(n1382) );
INV_X1 U1049 ( .A(G217), .ZN(n1384) );
NAND2_X1 U1050 ( .A1(n1385), .A2(KEYINPUT57), .ZN(n1381) );
XOR2_X1 U1051 ( .A(n1386), .B(n1387), .Z(n1385) );
NOR2_X1 U1052 ( .A1(KEYINPUT51), .A2(n1370), .ZN(n1387) );
AND2_X1 U1053 ( .A1(n1105), .A2(n1107), .ZN(n1305) );
NAND2_X1 U1054 ( .A1(n1123), .A2(n1388), .ZN(n1107) );
NAND4_X1 U1055 ( .A1(n1213), .A2(G953), .A3(G902), .A4(n1337), .ZN(n1388) );
XNOR2_X1 U1056 ( .A(G898), .B(KEYINPUT25), .ZN(n1213) );
NAND3_X1 U1057 ( .A1(n1337), .A2(n1142), .A3(G952), .ZN(n1123) );
NAND2_X1 U1058 ( .A1(G237), .A2(G234), .ZN(n1337) );
NOR2_X1 U1059 ( .A1(n1147), .A2(n1294), .ZN(n1105) );
NAND2_X1 U1060 ( .A1(n1137), .A2(n1138), .ZN(n1294) );
NAND2_X1 U1061 ( .A1(G221), .A2(n1389), .ZN(n1138) );
XOR2_X1 U1062 ( .A(n1171), .B(G469), .Z(n1137) );
AND2_X1 U1063 ( .A1(n1390), .A2(n1360), .ZN(n1171) );
XOR2_X1 U1064 ( .A(n1391), .B(n1392), .Z(n1390) );
XOR2_X1 U1065 ( .A(G140), .B(G110), .Z(n1392) );
XOR2_X1 U1066 ( .A(n1261), .B(n1263), .Z(n1391) );
AND2_X1 U1067 ( .A1(G227), .A2(n1142), .ZN(n1263) );
XOR2_X1 U1068 ( .A(n1393), .B(n1248), .Z(n1261) );
XOR2_X1 U1069 ( .A(n1195), .B(n1394), .Z(n1393) );
NOR3_X1 U1070 ( .A1(n1395), .A2(n1396), .A3(n1397), .ZN(n1394) );
NOR2_X1 U1071 ( .A1(n1096), .A2(n1398), .ZN(n1397) );
XOR2_X1 U1072 ( .A(G104), .B(G101), .Z(n1398) );
NOR3_X1 U1073 ( .A1(G107), .A2(G101), .A3(n1236), .ZN(n1396) );
NOR2_X1 U1074 ( .A1(n1333), .A2(n1399), .ZN(n1395) );
INV_X1 U1075 ( .A(G101), .ZN(n1333) );
NAND3_X1 U1076 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n1195) );
OR2_X1 U1077 ( .A1(n1403), .A2(KEYINPUT58), .ZN(n1402) );
NAND3_X1 U1078 ( .A1(KEYINPUT58), .A2(n1403), .A3(n1386), .ZN(n1401) );
INV_X1 U1079 ( .A(G128), .ZN(n1386) );
NAND2_X1 U1080 ( .A1(G128), .A2(n1404), .ZN(n1400) );
NAND2_X1 U1081 ( .A1(KEYINPUT58), .A2(n1405), .ZN(n1404) );
XOR2_X1 U1082 ( .A(KEYINPUT34), .B(n1403), .Z(n1405) );
INV_X1 U1083 ( .A(n1320), .ZN(n1147) );
NOR2_X1 U1084 ( .A1(n1149), .A2(n1115), .ZN(n1320) );
AND2_X1 U1085 ( .A1(G214), .A2(n1406), .ZN(n1115) );
XOR2_X1 U1086 ( .A(n1280), .B(n1407), .Z(n1149) );
NOR2_X1 U1087 ( .A1(G902), .A2(n1408), .ZN(n1407) );
XOR2_X1 U1088 ( .A(n1409), .B(n1410), .Z(n1408) );
NOR2_X1 U1089 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
XOR2_X1 U1090 ( .A(n1413), .B(KEYINPUT48), .Z(n1412) );
NAND2_X1 U1091 ( .A1(n1414), .A2(n1275), .ZN(n1413) );
NOR2_X1 U1092 ( .A1(n1275), .A2(n1414), .ZN(n1411) );
NAND2_X1 U1093 ( .A1(n1415), .A2(n1416), .ZN(n1414) );
OR2_X1 U1094 ( .A1(n1278), .A2(n1247), .ZN(n1416) );
XOR2_X1 U1095 ( .A(n1417), .B(KEYINPUT10), .Z(n1415) );
NAND2_X1 U1096 ( .A1(n1247), .A2(n1278), .ZN(n1417) );
NAND2_X1 U1097 ( .A1(G224), .A2(n1142), .ZN(n1275) );
NAND2_X1 U1098 ( .A1(KEYINPUT38), .A2(n1273), .ZN(n1409) );
XOR2_X1 U1099 ( .A(n1215), .B(n1214), .Z(n1273) );
XOR2_X1 U1100 ( .A(n1418), .B(n1419), .Z(n1214) );
XOR2_X1 U1101 ( .A(G122), .B(G110), .Z(n1419) );
NAND2_X1 U1102 ( .A1(n1420), .A2(n1421), .ZN(n1418) );
OR2_X1 U1103 ( .A1(n1422), .A2(n1251), .ZN(n1421) );
NAND3_X1 U1104 ( .A1(n1423), .A2(n1424), .A3(n1422), .ZN(n1420) );
INV_X1 U1105 ( .A(KEYINPUT6), .ZN(n1422) );
NAND2_X1 U1106 ( .A1(n1425), .A2(n1426), .ZN(n1215) );
NAND3_X1 U1107 ( .A1(n1399), .A2(n1427), .A3(G101), .ZN(n1426) );
XOR2_X1 U1108 ( .A(KEYINPUT29), .B(n1428), .Z(n1425) );
NOR2_X1 U1109 ( .A1(G101), .A2(n1429), .ZN(n1428) );
AND2_X1 U1110 ( .A1(n1399), .A2(n1427), .ZN(n1429) );
NAND2_X1 U1111 ( .A1(G107), .A2(n1430), .ZN(n1427) );
XOR2_X1 U1112 ( .A(KEYINPUT60), .B(G104), .Z(n1430) );
NAND2_X1 U1113 ( .A1(n1096), .A2(n1236), .ZN(n1399) );
INV_X1 U1114 ( .A(G104), .ZN(n1236) );
INV_X1 U1115 ( .A(G107), .ZN(n1096) );
NAND2_X1 U1116 ( .A1(G210), .A2(n1406), .ZN(n1280) );
NAND2_X1 U1117 ( .A1(n1431), .A2(n1360), .ZN(n1406) );
INV_X1 U1118 ( .A(G237), .ZN(n1431) );
INV_X1 U1119 ( .A(n1120), .ZN(n1335) );
NAND2_X1 U1120 ( .A1(n1355), .A2(n1432), .ZN(n1120) );
XNOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1352), .ZN(n1432) );
XNOR2_X1 U1122 ( .A(n1164), .B(n1433), .ZN(n1352) );
NOR2_X1 U1123 ( .A1(n1160), .A2(KEYINPUT32), .ZN(n1433) );
INV_X1 U1124 ( .A(n1163), .ZN(n1160) );
NAND2_X1 U1125 ( .A1(G217), .A2(n1389), .ZN(n1163) );
NAND2_X1 U1126 ( .A1(G234), .A2(n1360), .ZN(n1389) );
INV_X1 U1127 ( .A(n1161), .ZN(n1164) );
NAND2_X1 U1128 ( .A1(n1223), .A2(n1360), .ZN(n1161) );
INV_X1 U1129 ( .A(n1226), .ZN(n1223) );
XOR2_X1 U1130 ( .A(n1434), .B(n1435), .Z(n1226) );
XOR2_X1 U1131 ( .A(n1436), .B(n1367), .Z(n1435) );
XOR2_X1 U1132 ( .A(G146), .B(n1184), .Z(n1367) );
XNOR2_X1 U1133 ( .A(n1278), .B(G140), .ZN(n1184) );
INV_X1 U1134 ( .A(G125), .ZN(n1278) );
NOR2_X1 U1135 ( .A1(n1383), .A2(n1437), .ZN(n1436) );
INV_X1 U1136 ( .A(G221), .ZN(n1437) );
NAND2_X1 U1137 ( .A1(G234), .A2(n1142), .ZN(n1383) );
INV_X1 U1138 ( .A(G953), .ZN(n1142) );
XOR2_X1 U1139 ( .A(n1438), .B(n1439), .Z(n1434) );
XOR2_X1 U1140 ( .A(KEYINPUT31), .B(G137), .Z(n1439) );
NAND3_X1 U1141 ( .A1(n1440), .A2(n1441), .A3(n1442), .ZN(n1438) );
NAND2_X1 U1142 ( .A1(KEYINPUT39), .A2(n1443), .ZN(n1442) );
NAND3_X1 U1143 ( .A1(n1444), .A2(n1445), .A3(n1267), .ZN(n1441) );
INV_X1 U1144 ( .A(KEYINPUT39), .ZN(n1445) );
OR2_X1 U1145 ( .A1(n1267), .A2(n1444), .ZN(n1440) );
NOR2_X1 U1146 ( .A1(KEYINPUT4), .A2(n1443), .ZN(n1444) );
XOR2_X1 U1147 ( .A(G128), .B(n1446), .Z(n1443) );
XNOR2_X1 U1148 ( .A(n1156), .B(KEYINPUT47), .ZN(n1355) );
XNOR2_X1 U1149 ( .A(n1447), .B(G472), .ZN(n1156) );
NAND2_X1 U1150 ( .A1(n1448), .A2(n1360), .ZN(n1447) );
INV_X1 U1151 ( .A(G902), .ZN(n1360) );
XOR2_X1 U1152 ( .A(n1449), .B(n1450), .Z(n1448) );
INV_X1 U1153 ( .A(n1242), .ZN(n1450) );
XOR2_X1 U1154 ( .A(n1451), .B(G101), .Z(n1242) );
NAND2_X1 U1155 ( .A1(G210), .A2(n1372), .ZN(n1451) );
NOR2_X1 U1156 ( .A1(G953), .A2(G237), .ZN(n1372) );
NOR2_X1 U1157 ( .A1(KEYINPUT33), .A2(n1452), .ZN(n1449) );
XOR2_X1 U1158 ( .A(n1251), .B(n1246), .Z(n1452) );
XOR2_X1 U1159 ( .A(n1248), .B(n1247), .Z(n1246) );
XNOR2_X1 U1160 ( .A(n1453), .B(n1454), .ZN(n1247) );
NOR2_X1 U1161 ( .A1(n1455), .A2(n1456), .ZN(n1454) );
AND3_X1 U1162 ( .A1(KEYINPUT55), .A2(n1316), .A3(n1370), .ZN(n1456) );
NOR2_X1 U1163 ( .A1(KEYINPUT55), .A2(n1457), .ZN(n1455) );
INV_X1 U1164 ( .A(n1403), .ZN(n1457) );
XOR2_X1 U1165 ( .A(n1316), .B(n1370), .Z(n1403) );
XNOR2_X1 U1166 ( .A(G143), .B(KEYINPUT35), .ZN(n1370) );
INV_X1 U1167 ( .A(G146), .ZN(n1316) );
NAND2_X1 U1168 ( .A1(KEYINPUT61), .A2(G128), .ZN(n1453) );
XOR2_X1 U1169 ( .A(G131), .B(n1201), .Z(n1248) );
XOR2_X1 U1170 ( .A(G134), .B(G137), .Z(n1201) );
XNOR2_X1 U1171 ( .A(n1424), .B(n1423), .ZN(n1251) );
INV_X1 U1172 ( .A(n1363), .ZN(n1423) );
XNOR2_X1 U1173 ( .A(G113), .B(KEYINPUT36), .ZN(n1363) );
XNOR2_X1 U1174 ( .A(G116), .B(n1446), .ZN(n1424) );
XOR2_X1 U1175 ( .A(G119), .B(KEYINPUT53), .Z(n1446) );
INV_X1 U1176 ( .A(G110), .ZN(n1267) );
endmodule


