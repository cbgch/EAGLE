//Key = 0110100011101111101110011101100010010010111000101001111111011011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301;

XNOR2_X1 U728 ( .A(n1000), .B(n1001), .ZN(G9) );
NAND3_X1 U729 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(G75) );
NAND2_X1 U730 ( .A1(G952), .A2(n1005), .ZN(n1004) );
NAND3_X1 U731 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1005) );
NAND2_X1 U732 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NAND2_X1 U733 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NAND3_X1 U734 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NAND2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND2_X1 U736 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
XOR2_X1 U737 ( .A(KEYINPUT0), .B(n1020), .Z(n1019) );
NAND2_X1 U738 ( .A1(n1021), .A2(n1020), .ZN(n1016) );
NAND2_X1 U739 ( .A1(n1022), .A2(n1023), .ZN(n1011) );
NAND2_X1 U740 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NAND3_X1 U741 ( .A1(n1020), .A2(n1026), .A3(n1015), .ZN(n1025) );
XNOR2_X1 U742 ( .A(n1027), .B(n1028), .ZN(n1026) );
NAND2_X1 U743 ( .A1(n1013), .A2(n1029), .ZN(n1024) );
NAND3_X1 U744 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND2_X1 U745 ( .A1(n1015), .A2(n1033), .ZN(n1032) );
NAND2_X1 U746 ( .A1(n1020), .A2(n1034), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U748 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
XNOR2_X1 U749 ( .A(n1039), .B(KEYINPUT28), .ZN(n1037) );
INV_X1 U750 ( .A(n1040), .ZN(n1035) );
NAND2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(n1030) );
XOR2_X1 U752 ( .A(KEYINPUT49), .B(n1015), .Z(n1042) );
NAND4_X1 U753 ( .A1(n1043), .A2(n1013), .A3(n1044), .A4(n1045), .ZN(n1002) );
NOR4_X1 U754 ( .A1(n1039), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1045) );
XNOR2_X1 U755 ( .A(n1049), .B(n1050), .ZN(n1048) );
XNOR2_X1 U756 ( .A(n1051), .B(KEYINPUT41), .ZN(n1049) );
AND2_X1 U757 ( .A1(n1052), .A2(G217), .ZN(n1047) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1044) );
XOR2_X1 U759 ( .A(n1055), .B(n1056), .Z(G72) );
XOR2_X1 U760 ( .A(n1057), .B(n1058), .Z(n1056) );
NAND2_X1 U761 ( .A1(G953), .A2(n1059), .ZN(n1058) );
NAND2_X1 U762 ( .A1(G900), .A2(G227), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1060), .A2(n1061), .ZN(n1057) );
NAND2_X1 U764 ( .A1(G953), .A2(n1062), .ZN(n1061) );
XOR2_X1 U765 ( .A(n1063), .B(n1064), .Z(n1060) );
XOR2_X1 U766 ( .A(n1065), .B(n1066), .Z(n1064) );
XNOR2_X1 U767 ( .A(n1067), .B(KEYINPUT57), .ZN(n1063) );
NOR2_X1 U768 ( .A1(n1006), .A2(G953), .ZN(n1055) );
XOR2_X1 U769 ( .A(n1068), .B(n1069), .Z(G69) );
XOR2_X1 U770 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U771 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
INV_X1 U772 ( .A(n1074), .ZN(n1073) );
NAND2_X1 U773 ( .A1(G953), .A2(n1075), .ZN(n1070) );
NAND2_X1 U774 ( .A1(G898), .A2(G224), .ZN(n1075) );
NOR2_X1 U775 ( .A1(n1008), .A2(G953), .ZN(n1068) );
NOR2_X1 U776 ( .A1(n1076), .A2(n1077), .ZN(G66) );
NOR3_X1 U777 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
INV_X1 U780 ( .A(KEYINPUT32), .ZN(n1084) );
XOR2_X1 U781 ( .A(n1085), .B(KEYINPUT48), .Z(n1083) );
AND3_X1 U782 ( .A1(n1082), .A2(n1085), .A3(KEYINPUT32), .ZN(n1079) );
XNOR2_X1 U783 ( .A(n1086), .B(KEYINPUT1), .ZN(n1082) );
NOR2_X1 U784 ( .A1(KEYINPUT32), .A2(n1085), .ZN(n1078) );
NAND2_X1 U785 ( .A1(n1087), .A2(G217), .ZN(n1085) );
NOR2_X1 U786 ( .A1(n1076), .A2(n1088), .ZN(G63) );
XNOR2_X1 U787 ( .A(n1089), .B(n1090), .ZN(n1088) );
AND2_X1 U788 ( .A1(G478), .A2(n1087), .ZN(n1089) );
NOR2_X1 U789 ( .A1(n1076), .A2(n1091), .ZN(G60) );
XNOR2_X1 U790 ( .A(n1092), .B(n1093), .ZN(n1091) );
AND2_X1 U791 ( .A1(G475), .A2(n1087), .ZN(n1093) );
XOR2_X1 U792 ( .A(G104), .B(n1094), .Z(G6) );
NOR2_X1 U793 ( .A1(KEYINPUT43), .A2(n1095), .ZN(n1094) );
NOR2_X1 U794 ( .A1(n1076), .A2(n1096), .ZN(G57) );
XOR2_X1 U795 ( .A(KEYINPUT17), .B(n1097), .Z(n1096) );
NOR2_X1 U796 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U797 ( .A(KEYINPUT45), .B(n1100), .Z(n1099) );
NOR2_X1 U798 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
AND2_X1 U799 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
XNOR2_X1 U800 ( .A(n1103), .B(n1104), .ZN(n1102) );
XOR2_X1 U801 ( .A(KEYINPUT21), .B(n1105), .Z(n1104) );
NOR2_X1 U802 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U803 ( .A(n1108), .B(KEYINPUT27), .Z(n1107) );
NAND2_X1 U804 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U805 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
XNOR2_X1 U806 ( .A(n1067), .B(KEYINPUT60), .ZN(n1109) );
XOR2_X1 U807 ( .A(n1111), .B(n1112), .Z(n1103) );
AND2_X1 U808 ( .A1(G472), .A2(n1087), .ZN(n1112) );
NOR2_X1 U809 ( .A1(n1076), .A2(n1113), .ZN(G54) );
XOR2_X1 U810 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND3_X1 U811 ( .A1(n1087), .A2(G469), .A3(KEYINPUT18), .ZN(n1115) );
INV_X1 U812 ( .A(n1116), .ZN(n1087) );
NAND3_X1 U813 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1114) );
OR2_X1 U814 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U815 ( .A1(KEYINPUT58), .A2(n1122), .ZN(n1118) );
NAND2_X1 U816 ( .A1(n1123), .A2(n1121), .ZN(n1122) );
XNOR2_X1 U817 ( .A(n1120), .B(KEYINPUT38), .ZN(n1123) );
NAND2_X1 U818 ( .A1(n1124), .A2(n1125), .ZN(n1117) );
INV_X1 U819 ( .A(KEYINPUT58), .ZN(n1125) );
NAND2_X1 U820 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
OR2_X1 U821 ( .A1(n1120), .A2(KEYINPUT38), .ZN(n1127) );
NAND3_X1 U822 ( .A1(n1120), .A2(n1121), .A3(KEYINPUT38), .ZN(n1126) );
XNOR2_X1 U823 ( .A(G101), .B(n1128), .ZN(n1121) );
XOR2_X1 U824 ( .A(n1129), .B(n1130), .Z(n1120) );
NAND3_X1 U825 ( .A1(n1131), .A2(n1132), .A3(KEYINPUT13), .ZN(n1129) );
OR3_X1 U826 ( .A1(n1133), .A2(G110), .A3(KEYINPUT15), .ZN(n1132) );
NAND2_X1 U827 ( .A1(n1134), .A2(KEYINPUT15), .ZN(n1131) );
XOR2_X1 U828 ( .A(G110), .B(n1133), .Z(n1134) );
NOR3_X1 U829 ( .A1(n1135), .A2(n1076), .A3(n1136), .ZN(G51) );
NOR3_X1 U830 ( .A1(n1137), .A2(n1072), .A3(n1138), .ZN(n1136) );
XOR2_X1 U831 ( .A(n1139), .B(n1140), .Z(n1137) );
NOR2_X1 U832 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U833 ( .A(KEYINPUT46), .ZN(n1142) );
NOR2_X1 U834 ( .A1(n1003), .A2(G952), .ZN(n1076) );
NOR2_X1 U835 ( .A1(n1143), .A2(n1144), .ZN(n1135) );
XOR2_X1 U836 ( .A(n1139), .B(n1145), .Z(n1144) );
AND2_X1 U837 ( .A1(n1141), .A2(KEYINPUT46), .ZN(n1145) );
XNOR2_X1 U838 ( .A(n1146), .B(n1147), .ZN(n1141) );
NOR2_X1 U839 ( .A1(KEYINPUT6), .A2(n1148), .ZN(n1147) );
NOR2_X1 U840 ( .A1(n1116), .A2(n1050), .ZN(n1139) );
NAND2_X1 U841 ( .A1(G902), .A2(n1149), .ZN(n1116) );
NAND2_X1 U842 ( .A1(n1008), .A2(n1006), .ZN(n1149) );
AND2_X1 U843 ( .A1(n1150), .A2(n1151), .ZN(n1006) );
AND4_X1 U844 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1151) );
NAND3_X1 U845 ( .A1(n1156), .A2(n1040), .A3(n1157), .ZN(n1154) );
AND4_X1 U846 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1150) );
AND4_X1 U847 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1008) );
NOR4_X1 U848 ( .A1(n1166), .A2(n1001), .A3(n1167), .A4(n1168), .ZN(n1165) );
AND3_X1 U849 ( .A1(n1020), .A2(n1169), .A3(n1018), .ZN(n1001) );
AND2_X1 U850 ( .A1(n1170), .A2(n1095), .ZN(n1164) );
NAND3_X1 U851 ( .A1(n1020), .A2(n1169), .A3(n1021), .ZN(n1095) );
NOR2_X1 U852 ( .A1(n1072), .A2(n1138), .ZN(n1143) );
INV_X1 U853 ( .A(KEYINPUT59), .ZN(n1138) );
XNOR2_X1 U854 ( .A(G146), .B(n1171), .ZN(G48) );
NAND2_X1 U855 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U856 ( .A1(KEYINPUT22), .A2(n1174), .ZN(n1173) );
OR2_X1 U857 ( .A1(KEYINPUT61), .A2(n1174), .ZN(n1172) );
INV_X1 U858 ( .A(n1161), .ZN(n1174) );
NAND3_X1 U859 ( .A1(n1021), .A2(n1040), .A3(n1175), .ZN(n1161) );
XNOR2_X1 U860 ( .A(G143), .B(n1176), .ZN(G45) );
NAND3_X1 U861 ( .A1(n1156), .A2(n1177), .A3(n1178), .ZN(n1176) );
XNOR2_X1 U862 ( .A(n1040), .B(KEYINPUT4), .ZN(n1178) );
XOR2_X1 U863 ( .A(KEYINPUT5), .B(n1157), .Z(n1177) );
XNOR2_X1 U864 ( .A(G140), .B(n1160), .ZN(G42) );
NAND4_X1 U865 ( .A1(n1015), .A2(n1179), .A3(n1021), .A4(n1033), .ZN(n1160) );
NAND2_X1 U866 ( .A1(n1180), .A2(n1181), .ZN(G39) );
NAND2_X1 U867 ( .A1(G137), .A2(n1159), .ZN(n1181) );
XOR2_X1 U868 ( .A(n1182), .B(KEYINPUT30), .Z(n1180) );
OR2_X1 U869 ( .A1(n1159), .A2(G137), .ZN(n1182) );
NAND3_X1 U870 ( .A1(n1015), .A2(n1022), .A3(n1175), .ZN(n1159) );
XNOR2_X1 U871 ( .A(G134), .B(n1153), .ZN(G36) );
NAND3_X1 U872 ( .A1(n1156), .A2(n1018), .A3(n1015), .ZN(n1153) );
XNOR2_X1 U873 ( .A(G131), .B(n1152), .ZN(G33) );
NAND3_X1 U874 ( .A1(n1156), .A2(n1021), .A3(n1015), .ZN(n1152) );
NOR2_X1 U875 ( .A1(n1183), .A2(n1184), .ZN(n1015) );
AND2_X1 U876 ( .A1(n1179), .A2(n1041), .ZN(n1156) );
XNOR2_X1 U877 ( .A(G128), .B(n1158), .ZN(G30) );
NAND3_X1 U878 ( .A1(n1018), .A2(n1040), .A3(n1175), .ZN(n1158) );
AND3_X1 U879 ( .A1(n1185), .A2(n1186), .A3(n1179), .ZN(n1175) );
AND3_X1 U880 ( .A1(n1187), .A2(n1027), .A3(n1028), .ZN(n1179) );
OR2_X1 U881 ( .A1(n1188), .A2(n1041), .ZN(n1186) );
NAND2_X1 U882 ( .A1(n1189), .A2(n1188), .ZN(n1185) );
NAND2_X1 U883 ( .A1(n1053), .A2(n1190), .ZN(n1189) );
XOR2_X1 U884 ( .A(G101), .B(n1166), .Z(G3) );
AND3_X1 U885 ( .A1(n1041), .A2(n1169), .A3(n1022), .ZN(n1166) );
XNOR2_X1 U886 ( .A(n1191), .B(n1192), .ZN(G27) );
NAND2_X1 U887 ( .A1(KEYINPUT54), .A2(n1155), .ZN(n1191) );
NAND4_X1 U888 ( .A1(n1021), .A2(n1033), .A3(n1193), .A4(n1013), .ZN(n1155) );
AND2_X1 U889 ( .A1(n1187), .A2(n1040), .ZN(n1193) );
NAND2_X1 U890 ( .A1(n1194), .A2(n1195), .ZN(n1187) );
NAND4_X1 U891 ( .A1(G953), .A2(G902), .A3(n1010), .A4(n1062), .ZN(n1195) );
INV_X1 U892 ( .A(G900), .ZN(n1062) );
XNOR2_X1 U893 ( .A(G122), .B(n1170), .ZN(G24) );
NAND3_X1 U894 ( .A1(n1196), .A2(n1020), .A3(n1157), .ZN(n1170) );
NOR2_X1 U895 ( .A1(n1197), .A2(n1043), .ZN(n1157) );
NOR2_X1 U896 ( .A1(n1190), .A2(n1053), .ZN(n1020) );
XOR2_X1 U897 ( .A(n1162), .B(n1198), .Z(G21) );
XNOR2_X1 U898 ( .A(KEYINPUT35), .B(n1199), .ZN(n1198) );
NAND4_X1 U899 ( .A1(n1200), .A2(n1196), .A3(n1022), .A4(n1053), .ZN(n1162) );
XNOR2_X1 U900 ( .A(n1190), .B(n1188), .ZN(n1200) );
INV_X1 U901 ( .A(KEYINPUT31), .ZN(n1188) );
XNOR2_X1 U902 ( .A(G116), .B(n1163), .ZN(G18) );
NAND3_X1 U903 ( .A1(n1041), .A2(n1018), .A3(n1196), .ZN(n1163) );
NOR2_X1 U904 ( .A1(n1201), .A2(n1043), .ZN(n1018) );
INV_X1 U905 ( .A(n1202), .ZN(n1043) );
XNOR2_X1 U906 ( .A(G113), .B(n1203), .ZN(G15) );
NAND2_X1 U907 ( .A1(KEYINPUT24), .A2(n1168), .ZN(n1203) );
AND3_X1 U908 ( .A1(n1196), .A2(n1041), .A3(n1021), .ZN(n1168) );
NOR2_X1 U909 ( .A1(n1197), .A2(n1202), .ZN(n1021) );
NOR2_X1 U910 ( .A1(n1190), .A2(n1204), .ZN(n1041) );
AND2_X1 U911 ( .A1(n1013), .A2(n1205), .ZN(n1196) );
NOR2_X1 U912 ( .A1(n1028), .A2(n1206), .ZN(n1013) );
INV_X1 U913 ( .A(n1027), .ZN(n1206) );
XOR2_X1 U914 ( .A(G110), .B(n1167), .Z(G12) );
AND3_X1 U915 ( .A1(n1022), .A2(n1169), .A3(n1033), .ZN(n1167) );
AND2_X1 U916 ( .A1(n1204), .A2(n1190), .ZN(n1033) );
NAND2_X1 U917 ( .A1(n1207), .A2(n1208), .ZN(n1190) );
NAND2_X1 U918 ( .A1(G217), .A2(n1052), .ZN(n1208) );
NAND2_X1 U919 ( .A1(n1209), .A2(n1210), .ZN(n1052) );
OR2_X1 U920 ( .A1(n1086), .A2(G234), .ZN(n1210) );
XNOR2_X1 U921 ( .A(n1046), .B(KEYINPUT47), .ZN(n1207) );
AND3_X1 U922 ( .A1(n1086), .A2(n1209), .A3(n1211), .ZN(n1046) );
NAND2_X1 U923 ( .A1(G217), .A2(n1212), .ZN(n1211) );
NAND2_X1 U924 ( .A1(n1213), .A2(n1214), .ZN(n1086) );
NAND2_X1 U925 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XOR2_X1 U926 ( .A(n1217), .B(KEYINPUT39), .Z(n1213) );
OR2_X1 U927 ( .A1(n1216), .A2(n1215), .ZN(n1217) );
XOR2_X1 U928 ( .A(n1218), .B(n1219), .Z(n1215) );
XOR2_X1 U929 ( .A(n1220), .B(n1221), .Z(n1219) );
XNOR2_X1 U930 ( .A(n1222), .B(G128), .ZN(n1221) );
XOR2_X1 U931 ( .A(KEYINPUT8), .B(KEYINPUT52), .Z(n1220) );
XOR2_X1 U932 ( .A(n1223), .B(n1066), .Z(n1218) );
XNOR2_X1 U933 ( .A(n1224), .B(n1199), .ZN(n1223) );
NAND2_X1 U934 ( .A1(n1225), .A2(KEYINPUT19), .ZN(n1224) );
XNOR2_X1 U935 ( .A(G110), .B(KEYINPUT51), .ZN(n1225) );
XNOR2_X1 U936 ( .A(n1226), .B(G137), .ZN(n1216) );
NAND3_X1 U937 ( .A1(G221), .A2(n1227), .A3(KEYINPUT56), .ZN(n1226) );
INV_X1 U938 ( .A(n1053), .ZN(n1204) );
XNOR2_X1 U939 ( .A(n1228), .B(G472), .ZN(n1053) );
NAND2_X1 U940 ( .A1(n1229), .A2(n1209), .ZN(n1228) );
XOR2_X1 U941 ( .A(n1230), .B(n1231), .Z(n1229) );
XOR2_X1 U942 ( .A(KEYINPUT37), .B(n1232), .Z(n1231) );
XNOR2_X1 U943 ( .A(n1111), .B(n1101), .ZN(n1230) );
XOR2_X1 U944 ( .A(n1233), .B(G101), .Z(n1101) );
NAND2_X1 U945 ( .A1(G210), .A2(n1234), .ZN(n1233) );
NAND2_X1 U946 ( .A1(n1235), .A2(n1236), .ZN(n1111) );
NAND2_X1 U947 ( .A1(G119), .A2(n1237), .ZN(n1236) );
NAND2_X1 U948 ( .A1(n1238), .A2(n1199), .ZN(n1235) );
XNOR2_X1 U949 ( .A(KEYINPUT50), .B(n1237), .ZN(n1238) );
XNOR2_X1 U950 ( .A(G116), .B(n1239), .ZN(n1237) );
AND3_X1 U951 ( .A1(n1028), .A2(n1027), .A3(n1205), .ZN(n1169) );
AND2_X1 U952 ( .A1(n1040), .A2(n1240), .ZN(n1205) );
NAND2_X1 U953 ( .A1(n1194), .A2(n1241), .ZN(n1240) );
NAND3_X1 U954 ( .A1(G902), .A2(n1010), .A3(n1074), .ZN(n1241) );
NOR2_X1 U955 ( .A1(n1003), .A2(G898), .ZN(n1074) );
NAND3_X1 U956 ( .A1(n1242), .A2(n1003), .A3(G952), .ZN(n1194) );
XNOR2_X1 U957 ( .A(KEYINPUT63), .B(n1010), .ZN(n1242) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1010) );
NOR2_X1 U959 ( .A1(n1038), .A2(n1183), .ZN(n1040) );
XOR2_X1 U960 ( .A(n1039), .B(KEYINPUT11), .Z(n1183) );
AND2_X1 U961 ( .A1(G214), .A2(n1243), .ZN(n1039) );
INV_X1 U962 ( .A(n1184), .ZN(n1038) );
XOR2_X1 U963 ( .A(n1050), .B(n1244), .Z(n1184) );
NOR2_X1 U964 ( .A1(n1051), .A2(KEYINPUT44), .ZN(n1244) );
AND2_X1 U965 ( .A1(n1245), .A2(n1246), .ZN(n1051) );
XNOR2_X1 U966 ( .A(G902), .B(KEYINPUT3), .ZN(n1246) );
XOR2_X1 U967 ( .A(n1072), .B(n1247), .Z(n1245) );
NOR2_X1 U968 ( .A1(KEYINPUT7), .A2(n1248), .ZN(n1247) );
XNOR2_X1 U969 ( .A(n1249), .B(n1148), .ZN(n1248) );
NAND2_X1 U970 ( .A1(G224), .A2(n1003), .ZN(n1148) );
NAND2_X1 U971 ( .A1(KEYINPUT14), .A2(n1146), .ZN(n1249) );
XNOR2_X1 U972 ( .A(G125), .B(n1067), .ZN(n1146) );
XOR2_X1 U973 ( .A(n1250), .B(n1251), .Z(n1072) );
XOR2_X1 U974 ( .A(n1252), .B(n1253), .Z(n1251) );
XNOR2_X1 U975 ( .A(G104), .B(G122), .ZN(n1253) );
NAND2_X1 U976 ( .A1(KEYINPUT10), .A2(n1254), .ZN(n1252) );
XNOR2_X1 U977 ( .A(n1199), .B(G116), .ZN(n1254) );
INV_X1 U978 ( .A(G119), .ZN(n1199) );
XOR2_X1 U979 ( .A(n1255), .B(n1239), .Z(n1250) );
XNOR2_X1 U980 ( .A(n1256), .B(KEYINPUT12), .ZN(n1239) );
XOR2_X1 U981 ( .A(n1257), .B(n1258), .Z(n1255) );
NAND2_X1 U982 ( .A1(KEYINPUT23), .A2(n1000), .ZN(n1257) );
INV_X1 U983 ( .A(G107), .ZN(n1000) );
NAND2_X1 U984 ( .A1(G210), .A2(n1243), .ZN(n1050) );
NAND2_X1 U985 ( .A1(n1259), .A2(n1209), .ZN(n1243) );
XNOR2_X1 U986 ( .A(G237), .B(KEYINPUT29), .ZN(n1259) );
NAND2_X1 U987 ( .A1(G221), .A2(n1260), .ZN(n1027) );
NAND2_X1 U988 ( .A1(G234), .A2(n1209), .ZN(n1260) );
XNOR2_X1 U989 ( .A(n1261), .B(G469), .ZN(n1028) );
NAND2_X1 U990 ( .A1(n1262), .A2(n1209), .ZN(n1261) );
XOR2_X1 U991 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U992 ( .A(n1130), .B(n1265), .Z(n1264) );
XNOR2_X1 U993 ( .A(KEYINPUT9), .B(KEYINPUT40), .ZN(n1265) );
NAND2_X1 U994 ( .A1(G227), .A2(n1003), .ZN(n1130) );
INV_X1 U995 ( .A(G953), .ZN(n1003) );
XNOR2_X1 U996 ( .A(n1128), .B(n1266), .ZN(n1263) );
XOR2_X1 U997 ( .A(n1133), .B(n1258), .Z(n1266) );
XOR2_X1 U998 ( .A(G101), .B(G110), .Z(n1258) );
XOR2_X1 U999 ( .A(G140), .B(KEYINPUT55), .Z(n1133) );
XNOR2_X1 U1000 ( .A(n1267), .B(n1232), .ZN(n1128) );
XNOR2_X1 U1001 ( .A(n1110), .B(n1067), .ZN(n1232) );
XOR2_X1 U1002 ( .A(G146), .B(n1268), .Z(n1067) );
XOR2_X1 U1003 ( .A(n1269), .B(KEYINPUT2), .Z(n1110) );
NAND2_X1 U1004 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U1005 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
INV_X1 U1006 ( .A(KEYINPUT16), .ZN(n1273) );
NAND2_X1 U1007 ( .A1(G131), .A2(n1274), .ZN(n1272) );
NAND2_X1 U1008 ( .A1(KEYINPUT16), .A2(n1065), .ZN(n1270) );
XNOR2_X1 U1009 ( .A(G131), .B(n1274), .ZN(n1065) );
XOR2_X1 U1010 ( .A(G134), .B(G137), .Z(n1274) );
XNOR2_X1 U1011 ( .A(KEYINPUT57), .B(n1275), .ZN(n1267) );
NOR2_X1 U1012 ( .A1(KEYINPUT26), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U1013 ( .A(G104), .B(G107), .ZN(n1276) );
NOR2_X1 U1014 ( .A1(n1202), .A2(n1201), .ZN(n1022) );
INV_X1 U1015 ( .A(n1197), .ZN(n1201) );
XOR2_X1 U1016 ( .A(n1054), .B(KEYINPUT20), .Z(n1197) );
XNOR2_X1 U1017 ( .A(n1277), .B(G475), .ZN(n1054) );
NAND2_X1 U1018 ( .A1(n1092), .A2(n1209), .ZN(n1277) );
INV_X1 U1019 ( .A(G902), .ZN(n1209) );
XNOR2_X1 U1020 ( .A(n1278), .B(n1279), .ZN(n1092) );
XOR2_X1 U1021 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U1022 ( .A(n1282), .B(G104), .ZN(n1281) );
INV_X1 U1023 ( .A(G131), .ZN(n1282) );
XNOR2_X1 U1024 ( .A(n1222), .B(G143), .ZN(n1280) );
INV_X1 U1025 ( .A(G146), .ZN(n1222) );
XOR2_X1 U1026 ( .A(n1283), .B(n1284), .Z(n1278) );
XOR2_X1 U1027 ( .A(n1285), .B(n1286), .Z(n1284) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1234), .ZN(n1286) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1234) );
NAND3_X1 U1030 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1285) );
NAND2_X1 U1031 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
INV_X1 U1032 ( .A(KEYINPUT53), .ZN(n1291) );
NAND3_X1 U1033 ( .A1(KEYINPUT53), .A2(n1292), .A3(n1293), .ZN(n1288) );
OR2_X1 U1034 ( .A1(n1293), .A2(n1292), .ZN(n1287) );
NOR2_X1 U1035 ( .A1(KEYINPUT34), .A2(n1290), .ZN(n1292) );
XOR2_X1 U1036 ( .A(n1256), .B(KEYINPUT25), .Z(n1290) );
XNOR2_X1 U1037 ( .A(G113), .B(KEYINPUT36), .ZN(n1256) );
NAND2_X1 U1038 ( .A1(KEYINPUT62), .A2(n1066), .ZN(n1283) );
XNOR2_X1 U1039 ( .A(n1192), .B(G140), .ZN(n1066) );
INV_X1 U1040 ( .A(G125), .ZN(n1192) );
XNOR2_X1 U1041 ( .A(n1294), .B(G478), .ZN(n1202) );
NAND2_X1 U1042 ( .A1(n1295), .A2(n1090), .ZN(n1294) );
XOR2_X1 U1043 ( .A(n1296), .B(n1297), .Z(n1090) );
XOR2_X1 U1044 ( .A(n1298), .B(n1299), .Z(n1297) );
NAND2_X1 U1045 ( .A1(G217), .A2(n1227), .ZN(n1299) );
NOR2_X1 U1046 ( .A1(n1212), .A2(G953), .ZN(n1227) );
INV_X1 U1047 ( .A(G234), .ZN(n1212) );
NAND2_X1 U1048 ( .A1(n1300), .A2(KEYINPUT42), .ZN(n1298) );
XNOR2_X1 U1049 ( .A(G134), .B(n1268), .ZN(n1300) );
XOR2_X1 U1050 ( .A(G128), .B(G143), .Z(n1268) );
XNOR2_X1 U1051 ( .A(G107), .B(n1301), .ZN(n1296) );
XNOR2_X1 U1052 ( .A(n1293), .B(G116), .ZN(n1301) );
INV_X1 U1053 ( .A(G122), .ZN(n1293) );
XNOR2_X1 U1054 ( .A(G902), .B(KEYINPUT33), .ZN(n1295) );
endmodule


