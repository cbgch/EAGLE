//Key = 0000110000011000101010000000001101101011100111101000010010001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370;

XNOR2_X1 U750 ( .A(G107), .B(n1036), .ZN(G9) );
NAND4_X1 U751 ( .A1(KEYINPUT30), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1036) );
INV_X1 U752 ( .A(n1040), .ZN(n1038) );
NAND3_X1 U753 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(G75) );
NAND2_X1 U754 ( .A1(G952), .A2(n1044), .ZN(n1043) );
NAND4_X1 U755 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1044) );
NAND2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NAND3_X1 U758 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NAND2_X1 U759 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NAND3_X1 U760 ( .A1(n1037), .A2(n1058), .A3(n1059), .ZN(n1057) );
NAND2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U762 ( .A1(n1062), .A2(n1063), .ZN(n1056) );
NAND2_X1 U763 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U764 ( .A1(n1059), .A2(n1066), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U766 ( .A1(n1037), .A2(n1069), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND4_X1 U769 ( .A1(n1062), .A2(n1059), .A3(n1037), .A4(n1074), .ZN(n1051) );
NAND2_X1 U770 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U771 ( .A1(n1077), .A2(n1055), .ZN(n1075) );
NAND4_X1 U772 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1041) );
NOR4_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
XNOR2_X1 U774 ( .A(n1086), .B(n1087), .ZN(n1085) );
XOR2_X1 U775 ( .A(KEYINPUT51), .B(n1088), .Z(n1084) );
NOR2_X1 U776 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XNOR2_X1 U777 ( .A(n1091), .B(n1092), .ZN(n1083) );
NOR2_X1 U778 ( .A1(KEYINPUT0), .A2(n1093), .ZN(n1092) );
NOR3_X1 U779 ( .A1(n1094), .A2(n1095), .A3(n1077), .ZN(n1080) );
NOR2_X1 U780 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
XNOR2_X1 U781 ( .A(n1098), .B(KEYINPUT24), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1079) );
XOR2_X1 U783 ( .A(n1099), .B(n1100), .Z(G72) );
XOR2_X1 U784 ( .A(n1101), .B(n1102), .Z(n1100) );
NOR2_X1 U785 ( .A1(n1103), .A2(G953), .ZN(n1102) );
NOR3_X1 U786 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
INV_X1 U787 ( .A(n1107), .ZN(n1105) );
NAND3_X1 U788 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1104) );
NOR2_X1 U789 ( .A1(n1111), .A2(n1112), .ZN(n1101) );
XOR2_X1 U790 ( .A(KEYINPUT9), .B(n1113), .Z(n1112) );
NOR2_X1 U791 ( .A1(G900), .A2(n1042), .ZN(n1113) );
XOR2_X1 U792 ( .A(n1114), .B(n1115), .Z(n1111) );
NOR2_X1 U793 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
INV_X1 U794 ( .A(n1118), .ZN(n1117) );
NAND3_X1 U795 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1114) );
NAND2_X1 U796 ( .A1(KEYINPUT57), .A2(n1122), .ZN(n1121) );
NAND3_X1 U797 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1120) );
INV_X1 U798 ( .A(KEYINPUT57), .ZN(n1124) );
OR2_X1 U799 ( .A1(n1125), .A2(n1123), .ZN(n1119) );
AND2_X1 U800 ( .A1(KEYINPUT40), .A2(n1126), .ZN(n1123) );
XOR2_X1 U801 ( .A(n1127), .B(KEYINPUT34), .Z(n1125) );
NOR2_X1 U802 ( .A1(n1128), .A2(n1042), .ZN(n1099) );
AND2_X1 U803 ( .A1(G227), .A2(G900), .ZN(n1128) );
XOR2_X1 U804 ( .A(n1129), .B(n1130), .Z(G69) );
NOR2_X1 U805 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U806 ( .A1(G224), .A2(n1042), .ZN(n1131) );
NOR3_X1 U807 ( .A1(KEYINPUT23), .A2(n1133), .A3(n1134), .ZN(n1129) );
NOR3_X1 U808 ( .A1(n1135), .A2(G953), .A3(n1136), .ZN(n1134) );
NOR3_X1 U809 ( .A1(n1137), .A2(n1132), .A3(n1138), .ZN(n1133) );
NOR2_X1 U810 ( .A1(G953), .A2(n1136), .ZN(n1138) );
AND2_X1 U811 ( .A1(n1139), .A2(n1048), .ZN(n1136) );
XNOR2_X1 U812 ( .A(n1046), .B(KEYINPUT4), .ZN(n1139) );
INV_X1 U813 ( .A(n1135), .ZN(n1137) );
XOR2_X1 U814 ( .A(n1140), .B(n1141), .Z(n1135) );
NAND2_X1 U815 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
INV_X1 U817 ( .A(KEYINPUT25), .ZN(n1145) );
NAND3_X1 U818 ( .A1(n1146), .A2(n1147), .A3(KEYINPUT25), .ZN(n1142) );
NOR2_X1 U819 ( .A1(n1148), .A2(n1149), .ZN(G66) );
XNOR2_X1 U820 ( .A(n1150), .B(n1151), .ZN(n1149) );
NOR2_X1 U821 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XNOR2_X1 U822 ( .A(KEYINPUT31), .B(n1154), .ZN(n1153) );
NOR3_X1 U823 ( .A1(n1148), .A2(n1155), .A3(n1156), .ZN(G63) );
NOR2_X1 U824 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XNOR2_X1 U825 ( .A(n1159), .B(KEYINPUT53), .ZN(n1158) );
INV_X1 U826 ( .A(n1160), .ZN(n1157) );
NOR2_X1 U827 ( .A1(n1160), .A2(n1161), .ZN(n1155) );
XNOR2_X1 U828 ( .A(KEYINPUT43), .B(n1162), .ZN(n1161) );
INV_X1 U829 ( .A(n1159), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1152), .A2(n1086), .ZN(n1159) );
NOR2_X1 U831 ( .A1(n1148), .A2(n1163), .ZN(G60) );
XOR2_X1 U832 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U833 ( .A(n1166), .B(KEYINPUT14), .Z(n1164) );
NAND2_X1 U834 ( .A1(n1167), .A2(G475), .ZN(n1166) );
XNOR2_X1 U835 ( .A(G104), .B(n1168), .ZN(G6) );
NAND4_X1 U836 ( .A1(n1169), .A2(n1170), .A3(n1037), .A4(n1171), .ZN(n1168) );
XNOR2_X1 U837 ( .A(n1172), .B(KEYINPUT49), .ZN(n1169) );
NOR2_X1 U838 ( .A1(n1148), .A2(n1173), .ZN(G57) );
XNOR2_X1 U839 ( .A(n1174), .B(n1175), .ZN(n1173) );
NOR3_X1 U840 ( .A1(n1176), .A2(KEYINPUT61), .A3(n1177), .ZN(n1175) );
NOR3_X1 U841 ( .A1(n1178), .A2(n1093), .A3(n1152), .ZN(n1177) );
XOR2_X1 U842 ( .A(KEYINPUT45), .B(n1179), .Z(n1178) );
NOR2_X1 U843 ( .A1(n1180), .A2(n1179), .ZN(n1176) );
XNOR2_X1 U844 ( .A(n1181), .B(KEYINPUT38), .ZN(n1179) );
NOR2_X1 U845 ( .A1(n1093), .A2(n1152), .ZN(n1180) );
NOR2_X1 U846 ( .A1(n1148), .A2(n1182), .ZN(G54) );
XOR2_X1 U847 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U848 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U849 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
AND2_X1 U850 ( .A1(KEYINPUT10), .A2(n1189), .ZN(n1188) );
NOR2_X1 U851 ( .A1(KEYINPUT59), .A2(n1189), .ZN(n1187) );
NAND2_X1 U852 ( .A1(n1167), .A2(G469), .ZN(n1189) );
NAND2_X1 U853 ( .A1(KEYINPUT18), .A2(n1190), .ZN(n1185) );
XOR2_X1 U854 ( .A(n1191), .B(n1192), .Z(n1183) );
NOR2_X1 U855 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U856 ( .A1(G110), .A2(n1195), .ZN(n1193) );
NAND2_X1 U857 ( .A1(n1196), .A2(n1197), .ZN(n1191) );
NOR2_X1 U858 ( .A1(n1148), .A2(n1198), .ZN(G51) );
XOR2_X1 U859 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U860 ( .A(n1201), .B(n1202), .Z(n1199) );
NOR2_X1 U861 ( .A1(KEYINPUT15), .A2(n1203), .ZN(n1202) );
NAND2_X1 U862 ( .A1(n1167), .A2(n1204), .ZN(n1201) );
INV_X1 U863 ( .A(n1152), .ZN(n1167) );
NAND2_X1 U864 ( .A1(G902), .A2(n1205), .ZN(n1152) );
NAND3_X1 U865 ( .A1(n1206), .A2(n1048), .A3(n1046), .ZN(n1205) );
AND4_X1 U866 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1046) );
NAND2_X1 U867 ( .A1(n1211), .A2(n1212), .ZN(n1207) );
XOR2_X1 U868 ( .A(n1213), .B(KEYINPUT36), .Z(n1211) );
NAND3_X1 U869 ( .A1(n1214), .A2(n1215), .A3(n1171), .ZN(n1048) );
NAND3_X1 U870 ( .A1(n1216), .A2(n1217), .A3(n1039), .ZN(n1215) );
NAND2_X1 U871 ( .A1(n1037), .A2(n1218), .ZN(n1217) );
NAND2_X1 U872 ( .A1(n1060), .A2(n1219), .ZN(n1218) );
OR2_X1 U873 ( .A1(n1061), .A2(KEYINPUT27), .ZN(n1219) );
INV_X1 U874 ( .A(n1170), .ZN(n1060) );
NAND2_X1 U875 ( .A1(n1062), .A2(n1220), .ZN(n1216) );
NAND2_X1 U876 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
OR2_X1 U877 ( .A1(n1067), .A2(KEYINPUT41), .ZN(n1222) );
XNOR2_X1 U878 ( .A(n1223), .B(KEYINPUT6), .ZN(n1221) );
NAND3_X1 U879 ( .A1(n1224), .A2(n1225), .A3(n1172), .ZN(n1214) );
INV_X1 U880 ( .A(n1039), .ZN(n1172) );
NAND3_X1 U881 ( .A1(n1037), .A2(n1226), .A3(KEYINPUT27), .ZN(n1225) );
NAND3_X1 U882 ( .A1(n1227), .A2(n1062), .A3(KEYINPUT41), .ZN(n1224) );
XOR2_X1 U883 ( .A(KEYINPUT54), .B(n1045), .Z(n1206) );
NOR2_X1 U884 ( .A1(n1228), .A2(n1106), .ZN(n1045) );
NAND4_X1 U885 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1106) );
NAND4_X1 U886 ( .A1(n1233), .A2(n1170), .A3(n1234), .A4(n1235), .ZN(n1229) );
XNOR2_X1 U887 ( .A(KEYINPUT3), .B(n1070), .ZN(n1235) );
XNOR2_X1 U888 ( .A(n1236), .B(KEYINPUT12), .ZN(n1228) );
NAND4_X1 U889 ( .A1(n1237), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1236) );
NAND4_X1 U890 ( .A1(n1233), .A2(n1226), .A3(n1212), .A4(n1238), .ZN(n1107) );
XNOR2_X1 U891 ( .A(KEYINPUT58), .B(n1076), .ZN(n1238) );
XOR2_X1 U892 ( .A(n1110), .B(KEYINPUT50), .Z(n1237) );
NAND2_X1 U893 ( .A1(n1239), .A2(n1240), .ZN(n1110) );
NOR2_X1 U894 ( .A1(n1042), .A2(G952), .ZN(n1148) );
NAND2_X1 U895 ( .A1(n1241), .A2(n1242), .ZN(G48) );
NAND2_X1 U896 ( .A1(G146), .A2(n1243), .ZN(n1242) );
XOR2_X1 U897 ( .A(n1244), .B(KEYINPUT7), .Z(n1241) );
OR2_X1 U898 ( .A1(n1243), .A2(G146), .ZN(n1244) );
NAND3_X1 U899 ( .A1(n1170), .A2(n1171), .A3(n1233), .ZN(n1243) );
INV_X1 U900 ( .A(n1245), .ZN(n1233) );
XOR2_X1 U901 ( .A(n1246), .B(G143), .Z(G45) );
NAND2_X1 U902 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
OR2_X1 U903 ( .A1(n1230), .A2(KEYINPUT55), .ZN(n1248) );
NAND3_X1 U904 ( .A1(n1249), .A2(n1171), .A3(n1223), .ZN(n1230) );
NAND4_X1 U905 ( .A1(n1171), .A2(n1068), .A3(n1249), .A4(KEYINPUT55), .ZN(n1247) );
AND3_X1 U906 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1249) );
XNOR2_X1 U907 ( .A(G140), .B(n1231), .ZN(G42) );
NAND3_X1 U908 ( .A1(n1227), .A2(n1240), .A3(n1170), .ZN(n1231) );
XNOR2_X1 U909 ( .A(G137), .B(n1232), .ZN(G39) );
NAND4_X1 U910 ( .A1(n1062), .A2(n1240), .A3(n1253), .A4(n1254), .ZN(n1232) );
XOR2_X1 U911 ( .A(n1255), .B(n1256), .Z(G36) );
NOR2_X1 U912 ( .A1(KEYINPUT47), .A2(n1257), .ZN(n1256) );
XOR2_X1 U913 ( .A(KEYINPUT2), .B(G134), .Z(n1257) );
NAND4_X1 U914 ( .A1(n1239), .A2(n1234), .A3(n1258), .A4(n1251), .ZN(n1255) );
XNOR2_X1 U915 ( .A(KEYINPUT1), .B(n1082), .ZN(n1258) );
XNOR2_X1 U916 ( .A(G131), .B(n1108), .ZN(G33) );
NAND3_X1 U917 ( .A1(n1170), .A2(n1240), .A3(n1223), .ZN(n1108) );
AND3_X1 U918 ( .A1(n1234), .A2(n1251), .A3(n1059), .ZN(n1240) );
INV_X1 U919 ( .A(n1082), .ZN(n1059) );
NAND2_X1 U920 ( .A1(n1073), .A2(n1259), .ZN(n1082) );
XOR2_X1 U921 ( .A(G128), .B(n1260), .Z(G30) );
NOR2_X1 U922 ( .A1(n1040), .A2(n1245), .ZN(n1260) );
NAND3_X1 U923 ( .A1(n1251), .A2(n1254), .A3(n1253), .ZN(n1245) );
NAND2_X1 U924 ( .A1(n1171), .A2(n1226), .ZN(n1040) );
INV_X1 U925 ( .A(n1061), .ZN(n1226) );
XNOR2_X1 U926 ( .A(n1261), .B(n1262), .ZN(G3) );
NOR2_X1 U927 ( .A1(n1068), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U928 ( .A(G125), .B(n1109), .ZN(G27) );
NAND4_X1 U929 ( .A1(n1264), .A2(n1227), .A3(n1212), .A4(n1251), .ZN(n1109) );
NAND2_X1 U930 ( .A1(n1265), .A2(n1266), .ZN(n1251) );
NAND4_X1 U931 ( .A1(n1267), .A2(G953), .A3(n1050), .A4(n1268), .ZN(n1266) );
INV_X1 U932 ( .A(G900), .ZN(n1268) );
XNOR2_X1 U933 ( .A(G902), .B(KEYINPUT5), .ZN(n1267) );
INV_X1 U934 ( .A(n1067), .ZN(n1227) );
XNOR2_X1 U935 ( .A(G122), .B(n1208), .ZN(G24) );
NAND4_X1 U936 ( .A1(n1269), .A2(n1037), .A3(n1252), .A4(n1250), .ZN(n1208) );
NOR2_X1 U937 ( .A1(n1254), .A2(n1253), .ZN(n1037) );
XNOR2_X1 U938 ( .A(G119), .B(n1209), .ZN(G21) );
NAND4_X1 U939 ( .A1(n1269), .A2(n1062), .A3(n1253), .A4(n1254), .ZN(n1209) );
INV_X1 U940 ( .A(n1270), .ZN(n1253) );
XNOR2_X1 U941 ( .A(G116), .B(n1210), .ZN(G18) );
NAND2_X1 U942 ( .A1(n1269), .A2(n1239), .ZN(n1210) );
NOR2_X1 U943 ( .A1(n1068), .A2(n1061), .ZN(n1239) );
NAND2_X1 U944 ( .A1(n1078), .A2(n1252), .ZN(n1061) );
INV_X1 U945 ( .A(n1223), .ZN(n1068) );
AND4_X1 U946 ( .A1(n1212), .A2(n1055), .A3(n1054), .A4(n1039), .ZN(n1269) );
XNOR2_X1 U947 ( .A(n1271), .B(n1272), .ZN(G15) );
NOR2_X1 U948 ( .A1(n1070), .A2(n1213), .ZN(n1272) );
NAND3_X1 U949 ( .A1(n1223), .A2(n1039), .A3(n1264), .ZN(n1213) );
AND3_X1 U950 ( .A1(n1055), .A2(n1054), .A3(n1170), .ZN(n1264) );
NOR2_X1 U951 ( .A1(n1252), .A2(n1078), .ZN(n1170) );
INV_X1 U952 ( .A(n1250), .ZN(n1078) );
NOR2_X1 U953 ( .A1(n1270), .A2(n1254), .ZN(n1223) );
XOR2_X1 U954 ( .A(G110), .B(n1273), .Z(G12) );
NOR2_X1 U955 ( .A1(n1067), .A2(n1263), .ZN(n1273) );
NAND3_X1 U956 ( .A1(n1171), .A2(n1039), .A3(n1062), .ZN(n1263) );
NOR2_X1 U957 ( .A1(n1250), .A2(n1252), .ZN(n1062) );
XOR2_X1 U958 ( .A(n1274), .B(n1275), .Z(n1252) );
XOR2_X1 U959 ( .A(KEYINPUT19), .B(n1087), .Z(n1275) );
NOR2_X1 U960 ( .A1(n1160), .A2(G902), .ZN(n1087) );
XNOR2_X1 U961 ( .A(n1276), .B(n1277), .ZN(n1160) );
XOR2_X1 U962 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U963 ( .A(G122), .B(G116), .Z(n1279) );
XOR2_X1 U964 ( .A(KEYINPUT62), .B(G134), .Z(n1278) );
XOR2_X1 U965 ( .A(n1280), .B(n1281), .Z(n1276) );
NOR2_X1 U966 ( .A1(KEYINPUT13), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U967 ( .A(G143), .B(n1283), .ZN(n1282) );
XOR2_X1 U968 ( .A(n1284), .B(G107), .Z(n1280) );
NAND3_X1 U969 ( .A1(G217), .A2(n1042), .A3(n1285), .ZN(n1284) );
NAND2_X1 U970 ( .A1(KEYINPUT44), .A2(n1086), .ZN(n1274) );
INV_X1 U971 ( .A(G478), .ZN(n1086) );
XNOR2_X1 U972 ( .A(n1286), .B(G475), .ZN(n1250) );
NAND2_X1 U973 ( .A1(n1165), .A2(n1287), .ZN(n1286) );
XNOR2_X1 U974 ( .A(n1288), .B(n1289), .ZN(n1165) );
XOR2_X1 U975 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U976 ( .A(n1292), .B(n1293), .Z(n1291) );
NAND2_X1 U977 ( .A1(G214), .A2(n1294), .ZN(n1293) );
NAND3_X1 U978 ( .A1(n1295), .A2(n1296), .A3(n1118), .ZN(n1292) );
NAND2_X1 U979 ( .A1(n1116), .A2(n1297), .ZN(n1296) );
INV_X1 U980 ( .A(KEYINPUT26), .ZN(n1297) );
NAND2_X1 U981 ( .A1(KEYINPUT26), .A2(G125), .ZN(n1295) );
XOR2_X1 U982 ( .A(n1298), .B(n1299), .Z(n1288) );
XOR2_X1 U983 ( .A(G131), .B(G122), .Z(n1299) );
XNOR2_X1 U984 ( .A(G113), .B(G104), .ZN(n1298) );
NAND2_X1 U985 ( .A1(n1265), .A2(n1300), .ZN(n1039) );
NAND3_X1 U986 ( .A1(n1132), .A2(n1050), .A3(G902), .ZN(n1300) );
NOR2_X1 U987 ( .A1(G898), .A2(n1042), .ZN(n1132) );
NAND3_X1 U988 ( .A1(G952), .A2(n1042), .A3(n1301), .ZN(n1265) );
XOR2_X1 U989 ( .A(n1050), .B(KEYINPUT8), .Z(n1301) );
NAND2_X1 U990 ( .A1(G237), .A2(G234), .ZN(n1050) );
NOR2_X1 U991 ( .A1(n1070), .A2(n1076), .ZN(n1171) );
INV_X1 U992 ( .A(n1234), .ZN(n1076) );
NOR2_X1 U993 ( .A1(n1055), .A2(n1077), .ZN(n1234) );
INV_X1 U994 ( .A(n1054), .ZN(n1077) );
NAND2_X1 U995 ( .A1(G221), .A2(n1302), .ZN(n1054) );
XOR2_X1 U996 ( .A(n1089), .B(n1303), .Z(n1055) );
NOR2_X1 U997 ( .A1(KEYINPUT37), .A2(n1304), .ZN(n1303) );
INV_X1 U998 ( .A(n1090), .ZN(n1304) );
XOR2_X1 U999 ( .A(G469), .B(KEYINPUT16), .Z(n1090) );
AND2_X1 U1000 ( .A1(n1305), .A2(n1287), .ZN(n1089) );
XNOR2_X1 U1001 ( .A(n1306), .B(n1190), .ZN(n1305) );
NAND2_X1 U1002 ( .A1(G227), .A2(n1042), .ZN(n1190) );
XOR2_X1 U1003 ( .A(n1307), .B(n1308), .Z(n1306) );
NOR2_X1 U1004 ( .A1(n1194), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1005 ( .A(n1310), .B(KEYINPUT33), .Z(n1309) );
NAND2_X1 U1006 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1007 ( .A(KEYINPUT46), .B(G110), .Z(n1312) );
XNOR2_X1 U1008 ( .A(KEYINPUT32), .B(n1195), .ZN(n1311) );
AND2_X1 U1009 ( .A1(G110), .A2(n1195), .ZN(n1194) );
INV_X1 U1010 ( .A(G140), .ZN(n1195) );
NAND3_X1 U1011 ( .A1(n1313), .A2(n1314), .A3(n1197), .ZN(n1307) );
NAND2_X1 U1012 ( .A1(n1315), .A2(n1316), .ZN(n1197) );
NAND2_X1 U1013 ( .A1(KEYINPUT17), .A2(n1317), .ZN(n1314) );
NAND3_X1 U1014 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n1317) );
INV_X1 U1015 ( .A(n1315), .ZN(n1320) );
NOR2_X1 U1016 ( .A1(n1127), .A2(n1126), .ZN(n1315) );
NAND2_X1 U1017 ( .A1(n1321), .A2(n1316), .ZN(n1319) );
NAND3_X1 U1018 ( .A1(n1126), .A2(n1127), .A3(n1322), .ZN(n1318) );
OR2_X1 U1019 ( .A1(n1196), .A2(KEYINPUT17), .ZN(n1313) );
AND2_X1 U1020 ( .A1(n1323), .A2(n1324), .ZN(n1196) );
NAND2_X1 U1021 ( .A1(n1325), .A2(n1127), .ZN(n1324) );
XNOR2_X1 U1022 ( .A(n1126), .B(n1316), .ZN(n1325) );
NAND3_X1 U1023 ( .A1(n1126), .A2(n1322), .A3(n1321), .ZN(n1323) );
INV_X1 U1024 ( .A(n1316), .ZN(n1322) );
XOR2_X1 U1025 ( .A(n1326), .B(n1327), .Z(n1316) );
NOR2_X1 U1026 ( .A1(G104), .A2(KEYINPUT63), .ZN(n1327) );
INV_X1 U1027 ( .A(n1122), .ZN(n1126) );
NAND2_X1 U1028 ( .A1(n1328), .A2(n1329), .ZN(n1122) );
NAND2_X1 U1029 ( .A1(n1283), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1030 ( .A(KEYINPUT60), .B(n1331), .Z(n1328) );
NOR2_X1 U1031 ( .A1(n1283), .A2(n1330), .ZN(n1331) );
XOR2_X1 U1032 ( .A(n1290), .B(KEYINPUT28), .Z(n1330) );
XNOR2_X1 U1033 ( .A(G143), .B(n1332), .ZN(n1290) );
INV_X1 U1034 ( .A(n1212), .ZN(n1070) );
NOR2_X1 U1035 ( .A1(n1073), .A2(n1072), .ZN(n1212) );
INV_X1 U1036 ( .A(n1259), .ZN(n1072) );
NAND2_X1 U1037 ( .A1(G214), .A2(n1333), .ZN(n1259) );
XOR2_X1 U1038 ( .A(n1334), .B(n1204), .Z(n1073) );
AND2_X1 U1039 ( .A1(G210), .A2(n1333), .ZN(n1204) );
NAND2_X1 U1040 ( .A1(n1335), .A2(n1287), .ZN(n1333) );
INV_X1 U1041 ( .A(G237), .ZN(n1335) );
NAND2_X1 U1042 ( .A1(n1336), .A2(n1287), .ZN(n1334) );
XNOR2_X1 U1043 ( .A(n1200), .B(n1337), .ZN(n1336) );
NOR2_X1 U1044 ( .A1(KEYINPUT52), .A2(n1338), .ZN(n1337) );
INV_X1 U1045 ( .A(n1203), .ZN(n1338) );
XOR2_X1 U1046 ( .A(n1144), .B(n1339), .Z(n1203) );
NOR2_X1 U1047 ( .A1(KEYINPUT22), .A2(n1141), .ZN(n1339) );
XNOR2_X1 U1048 ( .A(G122), .B(G110), .ZN(n1141) );
XOR2_X1 U1049 ( .A(n1146), .B(n1147), .Z(n1144) );
XOR2_X1 U1050 ( .A(G104), .B(n1326), .Z(n1146) );
XOR2_X1 U1051 ( .A(G101), .B(G107), .Z(n1326) );
XNOR2_X1 U1052 ( .A(n1340), .B(n1341), .ZN(n1200) );
XOR2_X1 U1053 ( .A(G125), .B(n1342), .Z(n1341) );
AND2_X1 U1054 ( .A1(n1042), .A2(G224), .ZN(n1342) );
NAND2_X1 U1055 ( .A1(n1270), .A2(n1254), .ZN(n1067) );
NAND2_X1 U1056 ( .A1(n1343), .A2(n1344), .ZN(n1254) );
NAND2_X1 U1057 ( .A1(n1098), .A2(n1345), .ZN(n1344) );
XNOR2_X1 U1058 ( .A(n1095), .B(KEYINPUT21), .ZN(n1343) );
NOR2_X1 U1059 ( .A1(n1345), .A2(n1098), .ZN(n1095) );
INV_X1 U1060 ( .A(n1154), .ZN(n1098) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1302), .ZN(n1154) );
NAND2_X1 U1062 ( .A1(G234), .A2(n1287), .ZN(n1302) );
INV_X1 U1063 ( .A(n1096), .ZN(n1345) );
NOR2_X1 U1064 ( .A1(n1346), .A2(G902), .ZN(n1096) );
INV_X1 U1065 ( .A(n1150), .ZN(n1346) );
XNOR2_X1 U1066 ( .A(n1347), .B(n1348), .ZN(n1150) );
XOR2_X1 U1067 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1068 ( .A(G137), .B(G119), .Z(n1350) );
XNOR2_X1 U1069 ( .A(KEYINPUT56), .B(n1332), .ZN(n1349) );
XOR2_X1 U1070 ( .A(n1351), .B(n1352), .Z(n1347) );
XOR2_X1 U1071 ( .A(n1353), .B(n1283), .Z(n1352) );
NAND3_X1 U1072 ( .A1(n1354), .A2(n1355), .A3(n1118), .ZN(n1353) );
NAND2_X1 U1073 ( .A1(G140), .A2(G125), .ZN(n1118) );
NAND2_X1 U1074 ( .A1(n1116), .A2(n1356), .ZN(n1355) );
INV_X1 U1075 ( .A(KEYINPUT42), .ZN(n1356) );
NOR2_X1 U1076 ( .A1(G140), .A2(G125), .ZN(n1116) );
NAND2_X1 U1077 ( .A1(KEYINPUT42), .A2(G125), .ZN(n1354) );
XOR2_X1 U1078 ( .A(n1357), .B(G110), .Z(n1351) );
NAND3_X1 U1079 ( .A1(n1285), .A2(n1042), .A3(G221), .ZN(n1357) );
INV_X1 U1080 ( .A(G953), .ZN(n1042) );
XNOR2_X1 U1081 ( .A(G234), .B(KEYINPUT11), .ZN(n1285) );
XNOR2_X1 U1082 ( .A(n1091), .B(n1358), .ZN(n1270) );
XNOR2_X1 U1083 ( .A(KEYINPUT39), .B(n1093), .ZN(n1358) );
INV_X1 U1084 ( .A(G472), .ZN(n1093) );
NAND2_X1 U1085 ( .A1(n1359), .A2(n1287), .ZN(n1091) );
INV_X1 U1086 ( .A(G902), .ZN(n1287) );
XNOR2_X1 U1087 ( .A(n1181), .B(n1360), .ZN(n1359) );
INV_X1 U1088 ( .A(n1174), .ZN(n1360) );
XOR2_X1 U1089 ( .A(n1361), .B(n1261), .Z(n1174) );
INV_X1 U1090 ( .A(G101), .ZN(n1261) );
NAND2_X1 U1091 ( .A1(G210), .A2(n1294), .ZN(n1361) );
NOR2_X1 U1092 ( .A1(G953), .A2(G237), .ZN(n1294) );
XOR2_X1 U1093 ( .A(n1362), .B(n1147), .Z(n1181) );
XNOR2_X1 U1094 ( .A(n1271), .B(n1363), .ZN(n1147) );
XOR2_X1 U1095 ( .A(G119), .B(G116), .Z(n1363) );
INV_X1 U1096 ( .A(G113), .ZN(n1271) );
XNOR2_X1 U1097 ( .A(n1340), .B(n1321), .ZN(n1362) );
INV_X1 U1098 ( .A(n1127), .ZN(n1321) );
XOR2_X1 U1099 ( .A(G131), .B(n1364), .Z(n1127) );
XOR2_X1 U1100 ( .A(G137), .B(G134), .Z(n1364) );
XNOR2_X1 U1101 ( .A(n1365), .B(n1283), .ZN(n1340) );
XNOR2_X1 U1102 ( .A(G128), .B(KEYINPUT20), .ZN(n1283) );
NAND4_X1 U1103 ( .A1(KEYINPUT48), .A2(n1366), .A3(n1367), .A4(n1368), .ZN(n1365) );
NAND3_X1 U1104 ( .A1(n1369), .A2(n1370), .A3(n1332), .ZN(n1368) );
INV_X1 U1105 ( .A(KEYINPUT35), .ZN(n1370) );
OR2_X1 U1106 ( .A1(n1332), .A2(n1369), .ZN(n1367) );
NOR2_X1 U1107 ( .A1(G143), .A2(KEYINPUT29), .ZN(n1369) );
INV_X1 U1108 ( .A(G146), .ZN(n1332) );
NAND2_X1 U1109 ( .A1(KEYINPUT35), .A2(G143), .ZN(n1366) );
endmodule


