//Key = 1100100010101110011111110101111011110101100111000101001111111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391;

XNOR2_X1 U760 ( .A(n1054), .B(n1055), .ZN(G9) );
NOR2_X1 U761 ( .A1(KEYINPUT53), .A2(n1056), .ZN(n1055) );
NOR2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(G75) );
NOR4_X1 U763 ( .A1(n1059), .A2(n1060), .A3(G953), .A4(n1061), .ZN(n1058) );
NOR4_X1 U764 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1060) );
NOR2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1062) );
NAND3_X1 U768 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1059) );
NAND2_X1 U769 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND2_X1 U770 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U771 ( .A1(n1070), .A2(n1079), .ZN(n1078) );
NAND2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND3_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
NAND2_X1 U774 ( .A1(n1071), .A2(n1085), .ZN(n1080) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U776 ( .A1(n1084), .A2(n1088), .ZN(n1087) );
OR2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U778 ( .A1(n1082), .A2(n1091), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U780 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
XOR2_X1 U781 ( .A(n1096), .B(KEYINPUT3), .Z(n1077) );
NAND4_X1 U782 ( .A1(n1097), .A2(n1070), .A3(n1098), .A4(n1099), .ZN(n1096) );
NOR2_X1 U783 ( .A1(n1065), .A2(n1063), .ZN(n1098) );
INV_X1 U784 ( .A(n1084), .ZN(n1063) );
INV_X1 U785 ( .A(n1100), .ZN(n1070) );
XOR2_X1 U786 ( .A(KEYINPUT52), .B(n1101), .Z(n1072) );
NOR3_X1 U787 ( .A1(n1061), .A2(G953), .A3(G952), .ZN(n1057) );
AND4_X1 U788 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1061) );
NOR3_X1 U789 ( .A1(n1106), .A2(n1107), .A3(n1097), .ZN(n1105) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(n1106) );
NOR2_X1 U791 ( .A1(G469), .A2(KEYINPUT36), .ZN(n1109) );
XOR2_X1 U792 ( .A(n1110), .B(KEYINPUT39), .Z(n1104) );
NAND4_X1 U793 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1110) );
NOR3_X1 U794 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
AND3_X1 U795 ( .A1(KEYINPUT51), .A2(n1118), .A3(n1119), .ZN(n1117) );
NOR2_X1 U796 ( .A1(KEYINPUT51), .A2(n1119), .ZN(n1116) );
XOR2_X1 U797 ( .A(n1120), .B(n1121), .Z(n1115) );
NAND2_X1 U798 ( .A1(KEYINPUT19), .A2(G472), .ZN(n1121) );
XOR2_X1 U799 ( .A(n1122), .B(n1123), .Z(n1111) );
NAND2_X1 U800 ( .A1(n1124), .A2(KEYINPUT34), .ZN(n1123) );
XNOR2_X1 U801 ( .A(G478), .B(KEYINPUT41), .ZN(n1124) );
NAND2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(n1103) );
XOR2_X1 U803 ( .A(n1127), .B(KEYINPUT16), .Z(n1125) );
NAND2_X1 U804 ( .A1(n1128), .A2(n1129), .ZN(n1102) );
XOR2_X1 U805 ( .A(n1127), .B(KEYINPUT4), .Z(n1128) );
XNOR2_X1 U806 ( .A(n1130), .B(KEYINPUT17), .ZN(n1127) );
XOR2_X1 U807 ( .A(n1131), .B(n1132), .Z(G72) );
NOR2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
AND2_X1 U809 ( .A1(G227), .A2(G900), .ZN(n1133) );
NAND2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1131) );
NAND3_X1 U811 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
INV_X1 U812 ( .A(n1140), .ZN(n1138) );
OR2_X1 U813 ( .A1(n1137), .A2(n1139), .ZN(n1135) );
NAND3_X1 U814 ( .A1(n1141), .A2(n1142), .A3(n1134), .ZN(n1139) );
NAND2_X1 U815 ( .A1(n1101), .A2(n1143), .ZN(n1142) );
INV_X1 U816 ( .A(KEYINPUT47), .ZN(n1143) );
NAND3_X1 U817 ( .A1(n1144), .A2(n1145), .A3(KEYINPUT47), .ZN(n1141) );
INV_X1 U818 ( .A(n1146), .ZN(n1145) );
XOR2_X1 U819 ( .A(n1147), .B(n1148), .Z(n1137) );
XOR2_X1 U820 ( .A(KEYINPUT9), .B(n1149), .Z(n1147) );
NAND2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(G69) );
NAND2_X1 U822 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
INV_X1 U823 ( .A(n1154), .ZN(n1153) );
NAND3_X1 U824 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1152) );
XOR2_X1 U825 ( .A(KEYINPUT24), .B(n1074), .Z(n1157) );
INV_X1 U826 ( .A(n1158), .ZN(n1156) );
NAND2_X1 U827 ( .A1(G953), .A2(n1159), .ZN(n1155) );
NAND2_X1 U828 ( .A1(n1154), .A2(n1160), .ZN(n1150) );
NAND2_X1 U829 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U830 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
INV_X1 U831 ( .A(KEYINPUT24), .ZN(n1164) );
NAND2_X1 U832 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
NAND2_X1 U833 ( .A1(n1074), .A2(n1134), .ZN(n1166) );
NAND2_X1 U834 ( .A1(G953), .A2(G224), .ZN(n1165) );
NAND2_X1 U835 ( .A1(KEYINPUT24), .A2(n1167), .ZN(n1161) );
NOR4_X1 U836 ( .A1(n1168), .A2(n1169), .A3(KEYINPUT11), .A4(n1158), .ZN(n1154) );
XOR2_X1 U837 ( .A(n1170), .B(KEYINPUT13), .Z(n1169) );
NAND2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U839 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
NOR2_X1 U840 ( .A1(n1173), .A2(n1174), .ZN(G66) );
XOR2_X1 U841 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U842 ( .A(KEYINPUT38), .B(n1177), .Z(n1176) );
NOR2_X1 U843 ( .A1(n1118), .A2(n1178), .ZN(n1177) );
NOR2_X1 U844 ( .A1(n1173), .A2(n1179), .ZN(G63) );
XOR2_X1 U845 ( .A(n1180), .B(n1181), .Z(n1179) );
XNOR2_X1 U846 ( .A(KEYINPUT40), .B(n1182), .ZN(n1181) );
NAND3_X1 U847 ( .A1(n1183), .A2(G478), .A3(KEYINPUT20), .ZN(n1180) );
NOR2_X1 U848 ( .A1(n1173), .A2(n1184), .ZN(G60) );
XNOR2_X1 U849 ( .A(n1185), .B(n1186), .ZN(n1184) );
AND2_X1 U850 ( .A1(G475), .A2(n1183), .ZN(n1186) );
XOR2_X1 U851 ( .A(n1187), .B(n1188), .Z(G6) );
NOR2_X1 U852 ( .A1(KEYINPUT15), .A2(n1189), .ZN(n1188) );
NOR2_X1 U853 ( .A1(n1173), .A2(n1190), .ZN(G57) );
XOR2_X1 U854 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U855 ( .A(n1193), .B(n1194), .Z(n1192) );
NAND2_X1 U856 ( .A1(KEYINPUT57), .A2(n1195), .ZN(n1194) );
NAND3_X1 U857 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1193) );
NAND2_X1 U858 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
OR3_X1 U859 ( .A1(n1200), .A2(n1199), .A3(n1201), .ZN(n1197) );
XOR2_X1 U860 ( .A(n1202), .B(KEYINPUT56), .Z(n1199) );
OR2_X1 U861 ( .A1(KEYINPUT26), .A2(n1148), .ZN(n1200) );
NAND2_X1 U862 ( .A1(n1148), .A2(n1201), .ZN(n1196) );
INV_X1 U863 ( .A(KEYINPUT18), .ZN(n1201) );
XNOR2_X1 U864 ( .A(n1203), .B(n1204), .ZN(n1191) );
AND2_X1 U865 ( .A1(G472), .A2(n1183), .ZN(n1204) );
NOR3_X1 U866 ( .A1(n1173), .A2(n1205), .A3(n1206), .ZN(G54) );
NOR2_X1 U867 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U868 ( .A(n1209), .B(n1210), .Z(n1207) );
NAND2_X1 U869 ( .A1(KEYINPUT21), .A2(n1211), .ZN(n1209) );
NOR2_X1 U870 ( .A1(n1212), .A2(n1213), .ZN(n1205) );
XOR2_X1 U871 ( .A(n1214), .B(n1210), .Z(n1213) );
XOR2_X1 U872 ( .A(n1215), .B(n1216), .Z(n1210) );
XOR2_X1 U873 ( .A(n1217), .B(n1218), .Z(n1215) );
AND2_X1 U874 ( .A1(G469), .A2(n1183), .ZN(n1218) );
INV_X1 U875 ( .A(n1178), .ZN(n1183) );
NAND2_X1 U876 ( .A1(G902), .A2(n1219), .ZN(n1178) );
NAND2_X1 U877 ( .A1(KEYINPUT49), .A2(n1220), .ZN(n1217) );
NAND2_X1 U878 ( .A1(KEYINPUT21), .A2(n1221), .ZN(n1214) );
INV_X1 U879 ( .A(n1211), .ZN(n1221) );
XOR2_X1 U880 ( .A(n1222), .B(G110), .Z(n1211) );
NAND2_X1 U881 ( .A1(KEYINPUT22), .A2(n1223), .ZN(n1222) );
INV_X1 U882 ( .A(G140), .ZN(n1223) );
NOR2_X1 U883 ( .A1(n1173), .A2(n1224), .ZN(G51) );
NOR3_X1 U884 ( .A1(n1130), .A2(n1225), .A3(n1226), .ZN(n1224) );
NOR3_X1 U885 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1226) );
AND2_X1 U886 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
NAND2_X1 U887 ( .A1(n1129), .A2(n1230), .ZN(n1227) );
XNOR2_X1 U888 ( .A(KEYINPUT12), .B(n1219), .ZN(n1230) );
NAND2_X1 U889 ( .A1(n1074), .A2(n1101), .ZN(n1219) );
NOR2_X1 U890 ( .A1(n1146), .A2(n1144), .ZN(n1101) );
NOR2_X1 U891 ( .A1(n1231), .A2(n1232), .ZN(n1144) );
XOR2_X1 U892 ( .A(KEYINPUT31), .B(n1233), .Z(n1232) );
NAND4_X1 U893 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1146) );
AND4_X1 U894 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1237) );
NAND2_X1 U895 ( .A1(n1242), .A2(n1067), .ZN(n1236) );
XOR2_X1 U896 ( .A(n1243), .B(KEYINPUT37), .Z(n1242) );
NAND3_X1 U897 ( .A1(n1083), .A2(n1089), .A3(n1244), .ZN(n1234) );
INV_X1 U898 ( .A(n1167), .ZN(n1074) );
NAND4_X1 U899 ( .A1(n1245), .A2(n1054), .A3(n1246), .A4(n1247), .ZN(n1167) );
NOR4_X1 U900 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1247) );
INV_X1 U901 ( .A(n1252), .ZN(n1250) );
NOR2_X1 U902 ( .A1(n1253), .A2(n1187), .ZN(n1246) );
AND3_X1 U903 ( .A1(n1084), .A2(n1254), .A3(n1090), .ZN(n1187) );
INV_X1 U904 ( .A(n1255), .ZN(n1253) );
NAND3_X1 U905 ( .A1(n1254), .A2(n1089), .A3(n1084), .ZN(n1054) );
INV_X1 U906 ( .A(n1126), .ZN(n1129) );
NOR2_X1 U907 ( .A1(n1134), .A2(G952), .ZN(n1173) );
XNOR2_X1 U908 ( .A(n1256), .B(n1235), .ZN(G48) );
NAND3_X1 U909 ( .A1(n1090), .A2(n1083), .A3(n1244), .ZN(n1235) );
NOR2_X1 U910 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U911 ( .A(KEYINPUT7), .B(KEYINPUT59), .ZN(n1257) );
XOR2_X1 U912 ( .A(G143), .B(n1259), .Z(G45) );
NOR2_X1 U913 ( .A1(n1260), .A2(n1243), .ZN(n1259) );
NAND3_X1 U914 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1243) );
NAND2_X1 U915 ( .A1(n1264), .A2(n1265), .ZN(G42) );
NAND2_X1 U916 ( .A1(G140), .A2(n1241), .ZN(n1265) );
XOR2_X1 U917 ( .A(KEYINPUT29), .B(n1266), .Z(n1264) );
NOR2_X1 U918 ( .A1(G140), .A2(n1241), .ZN(n1266) );
NAND3_X1 U919 ( .A1(n1075), .A2(n1083), .A3(n1267), .ZN(n1241) );
XOR2_X1 U920 ( .A(n1240), .B(n1268), .Z(G39) );
NAND2_X1 U921 ( .A1(KEYINPUT32), .A2(G137), .ZN(n1268) );
NAND4_X1 U922 ( .A1(n1269), .A2(n1270), .A3(n1083), .A4(n1271), .ZN(n1240) );
NOR2_X1 U923 ( .A1(n1065), .A2(n1233), .ZN(n1271) );
XNOR2_X1 U924 ( .A(G134), .B(n1239), .ZN(G36) );
NAND3_X1 U925 ( .A1(n1075), .A2(n1089), .A3(n1263), .ZN(n1239) );
XOR2_X1 U926 ( .A(G131), .B(n1272), .Z(G33) );
NOR2_X1 U927 ( .A1(n1233), .A2(n1231), .ZN(n1272) );
NAND2_X1 U928 ( .A1(n1263), .A2(n1090), .ZN(n1231) );
AND3_X1 U929 ( .A1(n1083), .A2(n1270), .A3(n1273), .ZN(n1263) );
INV_X1 U930 ( .A(n1075), .ZN(n1233) );
NOR2_X1 U931 ( .A1(n1068), .A2(n1107), .ZN(n1075) );
INV_X1 U932 ( .A(n1069), .ZN(n1107) );
XNOR2_X1 U933 ( .A(G128), .B(n1274), .ZN(G30) );
NAND3_X1 U934 ( .A1(n1244), .A2(n1089), .A3(n1275), .ZN(n1274) );
XNOR2_X1 U935 ( .A(n1083), .B(KEYINPUT35), .ZN(n1275) );
AND3_X1 U936 ( .A1(n1269), .A2(n1270), .A3(n1067), .ZN(n1244) );
XOR2_X1 U937 ( .A(n1195), .B(n1255), .Z(G3) );
NAND3_X1 U938 ( .A1(n1254), .A2(n1082), .A3(n1273), .ZN(n1255) );
INV_X1 U939 ( .A(G101), .ZN(n1195) );
XNOR2_X1 U940 ( .A(n1238), .B(n1276), .ZN(G27) );
NOR2_X1 U941 ( .A1(KEYINPUT50), .A2(n1277), .ZN(n1276) );
NAND3_X1 U942 ( .A1(n1071), .A2(n1067), .A3(n1267), .ZN(n1238) );
AND4_X1 U943 ( .A1(n1090), .A2(n1094), .A3(n1270), .A4(n1095), .ZN(n1267) );
NAND2_X1 U944 ( .A1(n1100), .A2(n1278), .ZN(n1270) );
NAND3_X1 U945 ( .A1(G902), .A2(n1279), .A3(n1140), .ZN(n1278) );
NOR2_X1 U946 ( .A1(n1134), .A2(G900), .ZN(n1140) );
XNOR2_X1 U947 ( .A(n1251), .B(n1280), .ZN(G24) );
XNOR2_X1 U948 ( .A(G122), .B(KEYINPUT48), .ZN(n1280) );
AND4_X1 U949 ( .A1(n1281), .A2(n1084), .A3(n1261), .A4(n1262), .ZN(n1251) );
NOR2_X1 U950 ( .A1(n1282), .A2(n1095), .ZN(n1084) );
XOR2_X1 U951 ( .A(G119), .B(n1283), .Z(G21) );
NOR2_X1 U952 ( .A1(KEYINPUT2), .A2(n1252), .ZN(n1283) );
NAND3_X1 U953 ( .A1(n1082), .A2(n1269), .A3(n1281), .ZN(n1252) );
NAND2_X1 U954 ( .A1(n1284), .A2(n1285), .ZN(n1269) );
OR2_X1 U955 ( .A1(n1092), .A2(KEYINPUT10), .ZN(n1285) );
INV_X1 U956 ( .A(n1273), .ZN(n1092) );
NAND3_X1 U957 ( .A1(n1095), .A2(n1282), .A3(KEYINPUT10), .ZN(n1284) );
XOR2_X1 U958 ( .A(G116), .B(n1249), .Z(G18) );
AND3_X1 U959 ( .A1(n1273), .A2(n1089), .A3(n1281), .ZN(n1249) );
NAND2_X1 U960 ( .A1(n1286), .A2(n1287), .ZN(n1089) );
OR2_X1 U961 ( .A1(n1065), .A2(KEYINPUT54), .ZN(n1287) );
INV_X1 U962 ( .A(n1082), .ZN(n1065) );
NAND3_X1 U963 ( .A1(n1262), .A2(n1113), .A3(KEYINPUT54), .ZN(n1286) );
XOR2_X1 U964 ( .A(G113), .B(n1248), .Z(G15) );
AND3_X1 U965 ( .A1(n1090), .A2(n1273), .A3(n1281), .ZN(n1248) );
AND2_X1 U966 ( .A1(n1071), .A2(n1288), .ZN(n1281) );
NOR2_X1 U967 ( .A1(n1289), .A2(n1097), .ZN(n1071) );
NOR2_X1 U968 ( .A1(n1095), .A2(n1094), .ZN(n1273) );
NOR2_X1 U969 ( .A1(n1262), .A2(n1113), .ZN(n1090) );
XOR2_X1 U970 ( .A(n1290), .B(n1245), .Z(G12) );
NAND4_X1 U971 ( .A1(n1254), .A2(n1082), .A3(n1094), .A4(n1095), .ZN(n1245) );
NAND3_X1 U972 ( .A1(n1291), .A2(n1292), .A3(n1112), .ZN(n1095) );
NAND2_X1 U973 ( .A1(n1293), .A2(n1294), .ZN(n1112) );
OR3_X1 U974 ( .A1(n1294), .A2(n1293), .A3(KEYINPUT62), .ZN(n1292) );
INV_X1 U975 ( .A(n1118), .ZN(n1293) );
NAND2_X1 U976 ( .A1(G217), .A2(n1295), .ZN(n1118) );
NAND2_X1 U977 ( .A1(KEYINPUT62), .A2(n1294), .ZN(n1291) );
INV_X1 U978 ( .A(n1119), .ZN(n1294) );
NOR2_X1 U979 ( .A1(n1175), .A2(G902), .ZN(n1119) );
XNOR2_X1 U980 ( .A(n1296), .B(n1297), .ZN(n1175) );
XOR2_X1 U981 ( .A(G137), .B(n1298), .Z(n1297) );
XOR2_X1 U982 ( .A(G146), .B(G140), .Z(n1298) );
XOR2_X1 U983 ( .A(n1299), .B(n1300), .Z(n1296) );
XOR2_X1 U984 ( .A(n1301), .B(n1302), .Z(n1300) );
NAND2_X1 U985 ( .A1(KEYINPUT44), .A2(n1277), .ZN(n1302) );
NAND2_X1 U986 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
NAND2_X1 U987 ( .A1(G110), .A2(n1305), .ZN(n1304) );
XOR2_X1 U988 ( .A(KEYINPUT1), .B(n1306), .Z(n1303) );
NOR2_X1 U989 ( .A1(G110), .A2(n1305), .ZN(n1306) );
XOR2_X1 U990 ( .A(G128), .B(G119), .Z(n1305) );
NAND3_X1 U991 ( .A1(G221), .A2(n1134), .A3(G234), .ZN(n1299) );
INV_X1 U992 ( .A(n1282), .ZN(n1094) );
NAND3_X1 U993 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1282) );
NAND2_X1 U994 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND2_X1 U995 ( .A1(KEYINPUT33), .A2(n1312), .ZN(n1311) );
XOR2_X1 U996 ( .A(KEYINPUT6), .B(n1313), .Z(n1312) );
NAND3_X1 U997 ( .A1(KEYINPUT33), .A2(n1314), .A3(n1313), .ZN(n1308) );
INV_X1 U998 ( .A(n1310), .ZN(n1314) );
XNOR2_X1 U999 ( .A(G472), .B(KEYINPUT45), .ZN(n1310) );
OR2_X1 U1000 ( .A1(n1313), .A2(KEYINPUT33), .ZN(n1307) );
INV_X1 U1001 ( .A(n1120), .ZN(n1313) );
NAND2_X1 U1002 ( .A1(n1315), .A2(n1229), .ZN(n1120) );
XOR2_X1 U1003 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1004 ( .A(n1148), .B(n1202), .ZN(n1317) );
XOR2_X1 U1005 ( .A(n1318), .B(n1319), .Z(n1202) );
XNOR2_X1 U1006 ( .A(G113), .B(G119), .ZN(n1318) );
XOR2_X1 U1007 ( .A(n1216), .B(n1320), .Z(n1148) );
XOR2_X1 U1008 ( .A(n1321), .B(G101), .Z(n1316) );
NAND2_X1 U1009 ( .A1(KEYINPUT60), .A2(n1203), .ZN(n1321) );
AND3_X1 U1010 ( .A1(n1322), .A2(n1134), .A3(G210), .ZN(n1203) );
NOR2_X1 U1011 ( .A1(n1262), .A2(n1261), .ZN(n1082) );
INV_X1 U1012 ( .A(n1113), .ZN(n1261) );
XOR2_X1 U1013 ( .A(n1323), .B(G475), .Z(n1113) );
NAND2_X1 U1014 ( .A1(n1185), .A2(n1229), .ZN(n1323) );
XNOR2_X1 U1015 ( .A(n1324), .B(n1325), .ZN(n1185) );
XOR2_X1 U1016 ( .A(n1326), .B(G122), .Z(n1324) );
NAND2_X1 U1017 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1018 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1019 ( .A(KEYINPUT14), .B(n1331), .Z(n1327) );
NOR2_X1 U1020 ( .A1(n1329), .A2(n1330), .ZN(n1331) );
NAND3_X1 U1021 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1330) );
NAND2_X1 U1022 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND2_X1 U1023 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
INV_X1 U1024 ( .A(KEYINPUT58), .ZN(n1338) );
NAND2_X1 U1025 ( .A1(n1339), .A2(n1340), .ZN(n1337) );
XOR2_X1 U1026 ( .A(KEYINPUT25), .B(n1336), .Z(n1340) );
INV_X1 U1027 ( .A(n1341), .ZN(n1336) );
NAND2_X1 U1028 ( .A1(KEYINPUT58), .A2(n1342), .ZN(n1332) );
NAND2_X1 U1029 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NAND3_X1 U1030 ( .A1(KEYINPUT25), .A2(n1339), .A3(n1341), .ZN(n1344) );
INV_X1 U1031 ( .A(n1335), .ZN(n1339) );
NAND2_X1 U1032 ( .A1(n1345), .A2(n1346), .ZN(n1335) );
NAND2_X1 U1033 ( .A1(KEYINPUT55), .A2(n1149), .ZN(n1346) );
XNOR2_X1 U1034 ( .A(G125), .B(G140), .ZN(n1149) );
OR3_X1 U1035 ( .A1(n1277), .A2(G140), .A3(KEYINPUT55), .ZN(n1345) );
OR2_X1 U1036 ( .A1(n1341), .A2(KEYINPUT25), .ZN(n1343) );
XOR2_X1 U1037 ( .A(n1258), .B(KEYINPUT23), .Z(n1341) );
XOR2_X1 U1038 ( .A(n1347), .B(n1348), .Z(n1329) );
XOR2_X1 U1039 ( .A(G143), .B(G131), .Z(n1348) );
NAND3_X1 U1040 ( .A1(n1322), .A2(n1134), .A3(G214), .ZN(n1347) );
XNOR2_X1 U1041 ( .A(G478), .B(n1122), .ZN(n1262) );
NAND2_X1 U1042 ( .A1(n1229), .A2(n1182), .ZN(n1122) );
NAND2_X1 U1043 ( .A1(n1349), .A2(n1350), .ZN(n1182) );
NAND2_X1 U1044 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XOR2_X1 U1045 ( .A(KEYINPUT30), .B(n1353), .Z(n1349) );
NOR2_X1 U1046 ( .A1(n1351), .A2(n1352), .ZN(n1353) );
XOR2_X1 U1047 ( .A(n1354), .B(n1355), .Z(n1352) );
XNOR2_X1 U1048 ( .A(n1356), .B(n1357), .ZN(n1355) );
NAND2_X1 U1049 ( .A1(n1358), .A2(KEYINPUT8), .ZN(n1356) );
XOR2_X1 U1050 ( .A(n1359), .B(G122), .Z(n1358) );
NAND2_X1 U1051 ( .A1(KEYINPUT0), .A2(n1360), .ZN(n1359) );
INV_X1 U1052 ( .A(G116), .ZN(n1360) );
XOR2_X1 U1053 ( .A(n1056), .B(G134), .Z(n1354) );
INV_X1 U1054 ( .A(G107), .ZN(n1056) );
AND3_X1 U1055 ( .A1(G234), .A2(n1361), .A3(G217), .ZN(n1351) );
XOR2_X1 U1056 ( .A(KEYINPUT27), .B(G953), .Z(n1361) );
AND2_X1 U1057 ( .A1(n1288), .A2(n1083), .ZN(n1254) );
NOR2_X1 U1058 ( .A1(n1099), .A2(n1097), .ZN(n1083) );
AND2_X1 U1059 ( .A1(G221), .A2(n1295), .ZN(n1097) );
NAND2_X1 U1060 ( .A1(n1362), .A2(n1229), .ZN(n1295) );
INV_X1 U1061 ( .A(n1289), .ZN(n1099) );
NAND2_X1 U1062 ( .A1(n1363), .A2(n1364), .ZN(n1289) );
OR2_X1 U1063 ( .A1(n1108), .A2(G469), .ZN(n1364) );
XOR2_X1 U1064 ( .A(n1365), .B(KEYINPUT46), .Z(n1363) );
NAND2_X1 U1065 ( .A1(G469), .A2(n1108), .ZN(n1365) );
NAND2_X1 U1066 ( .A1(n1366), .A2(n1229), .ZN(n1108) );
XOR2_X1 U1067 ( .A(n1367), .B(n1368), .Z(n1366) );
XOR2_X1 U1068 ( .A(n1369), .B(n1212), .Z(n1368) );
INV_X1 U1069 ( .A(n1208), .ZN(n1212) );
NAND2_X1 U1070 ( .A1(G227), .A2(n1134), .ZN(n1208) );
NAND2_X1 U1071 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1072 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
INV_X1 U1073 ( .A(KEYINPUT28), .ZN(n1373) );
XOR2_X1 U1074 ( .A(n1374), .B(n1216), .Z(n1372) );
NAND2_X1 U1075 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
NAND2_X1 U1076 ( .A1(KEYINPUT28), .A2(n1377), .ZN(n1370) );
XOR2_X1 U1077 ( .A(n1220), .B(n1216), .Z(n1377) );
XOR2_X1 U1078 ( .A(G131), .B(n1378), .Z(n1216) );
XOR2_X1 U1079 ( .A(G137), .B(G134), .Z(n1378) );
XNOR2_X1 U1080 ( .A(n1375), .B(n1376), .ZN(n1220) );
XNOR2_X1 U1081 ( .A(n1320), .B(n1379), .ZN(n1376) );
XOR2_X1 U1082 ( .A(KEYINPUT9), .B(KEYINPUT63), .Z(n1379) );
XOR2_X1 U1083 ( .A(n1189), .B(n1380), .Z(n1375) );
INV_X1 U1084 ( .A(G104), .ZN(n1189) );
XOR2_X1 U1085 ( .A(n1290), .B(G140), .Z(n1367) );
AND2_X1 U1086 ( .A1(n1067), .A2(n1381), .ZN(n1288) );
NAND2_X1 U1087 ( .A1(n1100), .A2(n1382), .ZN(n1381) );
NAND3_X1 U1088 ( .A1(n1158), .A2(n1279), .A3(G902), .ZN(n1382) );
NOR2_X1 U1089 ( .A1(G898), .A2(n1134), .ZN(n1158) );
NAND3_X1 U1090 ( .A1(n1279), .A2(n1134), .A3(G952), .ZN(n1100) );
INV_X1 U1091 ( .A(G953), .ZN(n1134) );
NAND2_X1 U1092 ( .A1(G237), .A2(n1362), .ZN(n1279) );
XOR2_X1 U1093 ( .A(G234), .B(KEYINPUT61), .Z(n1362) );
INV_X1 U1094 ( .A(n1260), .ZN(n1067) );
NAND2_X1 U1095 ( .A1(n1068), .A2(n1069), .ZN(n1260) );
NAND2_X1 U1096 ( .A1(G214), .A2(n1383), .ZN(n1069) );
XNOR2_X1 U1097 ( .A(n1126), .B(n1130), .ZN(n1068) );
AND2_X1 U1098 ( .A1(n1228), .A2(n1229), .ZN(n1130) );
XOR2_X1 U1099 ( .A(n1384), .B(n1385), .Z(n1228) );
XNOR2_X1 U1100 ( .A(n1320), .B(n1172), .ZN(n1385) );
XOR2_X1 U1101 ( .A(G122), .B(n1290), .Z(n1172) );
XNOR2_X1 U1102 ( .A(n1258), .B(n1357), .ZN(n1320) );
XOR2_X1 U1103 ( .A(G143), .B(G128), .Z(n1357) );
INV_X1 U1104 ( .A(G146), .ZN(n1258) );
XOR2_X1 U1105 ( .A(n1386), .B(n1387), .Z(n1384) );
NOR2_X1 U1106 ( .A1(KEYINPUT42), .A2(n1171), .ZN(n1387) );
XOR2_X1 U1107 ( .A(n1388), .B(n1389), .Z(n1171) );
XOR2_X1 U1108 ( .A(n1325), .B(n1380), .Z(n1389) );
XOR2_X1 U1109 ( .A(G107), .B(G101), .Z(n1380) );
XOR2_X1 U1110 ( .A(G104), .B(G113), .Z(n1325) );
XOR2_X1 U1111 ( .A(n1390), .B(G119), .Z(n1388) );
NAND2_X1 U1112 ( .A1(KEYINPUT43), .A2(n1319), .ZN(n1390) );
XNOR2_X1 U1113 ( .A(G116), .B(KEYINPUT5), .ZN(n1319) );
XOR2_X1 U1114 ( .A(n1277), .B(n1391), .Z(n1386) );
NOR2_X1 U1115 ( .A1(G953), .A2(n1159), .ZN(n1391) );
INV_X1 U1116 ( .A(G224), .ZN(n1159) );
INV_X1 U1117 ( .A(G125), .ZN(n1277) );
NAND2_X1 U1118 ( .A1(G210), .A2(n1383), .ZN(n1126) );
NAND2_X1 U1119 ( .A1(n1229), .A2(n1322), .ZN(n1383) );
INV_X1 U1120 ( .A(G237), .ZN(n1322) );
INV_X1 U1121 ( .A(G902), .ZN(n1229) );
INV_X1 U1122 ( .A(G110), .ZN(n1290) );
endmodule


