//Key = 1001000010110100100101010001011001011000101101011100010011000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378;

XOR2_X1 U768 ( .A(G107), .B(n1052), .Z(G9) );
NOR2_X1 U769 ( .A1(KEYINPUT41), .A2(n1053), .ZN(n1052) );
NOR2_X1 U770 ( .A1(n1054), .A2(n1055), .ZN(G75) );
NOR3_X1 U771 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND3_X1 U772 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1056) );
NAND2_X1 U773 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U774 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND3_X1 U775 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NAND2_X1 U776 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND2_X1 U777 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
OR2_X1 U778 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U779 ( .A1(n1075), .A2(n1076), .ZN(n1069) );
XOR2_X1 U780 ( .A(n1077), .B(n1078), .Z(n1076) );
NAND3_X1 U781 ( .A1(n1071), .A2(n1079), .A3(n1075), .ZN(n1064) );
NAND2_X1 U782 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U783 ( .A1(n1068), .A2(n1082), .ZN(n1081) );
NAND2_X1 U784 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U785 ( .A1(n1066), .A2(n1085), .ZN(n1080) );
NAND2_X1 U786 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U787 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR3_X1 U788 ( .A1(n1090), .A2(G953), .A3(n1091), .ZN(n1054) );
INV_X1 U789 ( .A(n1059), .ZN(n1091) );
NAND4_X1 U790 ( .A1(n1092), .A2(n1071), .A3(n1093), .A4(n1094), .ZN(n1059) );
NOR4_X1 U791 ( .A1(n1095), .A2(n1088), .A3(n1096), .A4(n1097), .ZN(n1094) );
XOR2_X1 U792 ( .A(n1098), .B(KEYINPUT30), .Z(n1096) );
NOR3_X1 U793 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1093) );
NOR3_X1 U794 ( .A1(n1102), .A2(KEYINPUT31), .A3(n1103), .ZN(n1101) );
AND2_X1 U795 ( .A1(n1102), .A2(KEYINPUT31), .ZN(n1100) );
XOR2_X1 U796 ( .A(G475), .B(n1104), .Z(n1099) );
XOR2_X1 U797 ( .A(n1105), .B(n1106), .Z(n1092) );
XOR2_X1 U798 ( .A(n1057), .B(KEYINPUT13), .Z(n1090) );
INV_X1 U799 ( .A(G952), .ZN(n1057) );
XOR2_X1 U800 ( .A(n1107), .B(n1108), .Z(G72) );
XOR2_X1 U801 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR3_X1 U802 ( .A1(n1111), .A2(KEYINPUT12), .A3(G953), .ZN(n1110) );
NOR2_X1 U803 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
XOR2_X1 U804 ( .A(KEYINPUT43), .B(G953), .Z(n1113) );
AND2_X1 U805 ( .A1(G227), .A2(G900), .ZN(n1112) );
NOR2_X1 U806 ( .A1(n1114), .A2(n1115), .ZN(n1107) );
XOR2_X1 U807 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U808 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U809 ( .A(n1120), .B(KEYINPUT35), .Z(n1119) );
NAND2_X1 U810 ( .A1(KEYINPUT8), .A2(n1121), .ZN(n1118) );
XOR2_X1 U811 ( .A(G137), .B(G134), .Z(n1121) );
XNOR2_X1 U812 ( .A(n1122), .B(n1123), .ZN(n1116) );
XOR2_X1 U813 ( .A(n1124), .B(n1125), .Z(G69) );
NOR2_X1 U814 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NOR2_X1 U815 ( .A1(n1060), .A2(n1128), .ZN(n1127) );
XOR2_X1 U816 ( .A(KEYINPUT20), .B(n1129), .Z(n1128) );
NOR2_X1 U817 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U818 ( .A1(G953), .A2(n1132), .ZN(n1126) );
NAND2_X1 U819 ( .A1(n1133), .A2(n1134), .ZN(n1124) );
NAND2_X1 U820 ( .A1(G953), .A2(n1131), .ZN(n1134) );
XOR2_X1 U821 ( .A(n1135), .B(n1136), .Z(n1133) );
XOR2_X1 U822 ( .A(n1137), .B(KEYINPUT56), .Z(n1135) );
NAND2_X1 U823 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U824 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U825 ( .A(KEYINPUT6), .B(n1142), .Z(n1141) );
XOR2_X1 U826 ( .A(KEYINPUT14), .B(n1143), .Z(n1140) );
NAND2_X1 U827 ( .A1(n1144), .A2(n1145), .ZN(n1138) );
XOR2_X1 U828 ( .A(n1146), .B(KEYINPUT14), .Z(n1145) );
XOR2_X1 U829 ( .A(n1147), .B(KEYINPUT34), .Z(n1144) );
NOR2_X1 U830 ( .A1(n1148), .A2(n1149), .ZN(G66) );
XOR2_X1 U831 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U832 ( .A1(KEYINPUT58), .A2(n1152), .ZN(n1151) );
XOR2_X1 U833 ( .A(n1153), .B(KEYINPUT19), .Z(n1152) );
NAND2_X1 U834 ( .A1(n1154), .A2(n1155), .ZN(n1150) );
NOR2_X1 U835 ( .A1(n1148), .A2(n1156), .ZN(G63) );
XNOR2_X1 U836 ( .A(n1157), .B(n1158), .ZN(n1156) );
AND2_X1 U837 ( .A1(G478), .A2(n1154), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1159), .A2(n1160), .ZN(G60) );
XOR2_X1 U839 ( .A(KEYINPUT15), .B(n1148), .Z(n1160) );
XOR2_X1 U840 ( .A(n1161), .B(n1162), .Z(n1159) );
AND2_X1 U841 ( .A1(G475), .A2(n1154), .ZN(n1162) );
XOR2_X1 U842 ( .A(n1163), .B(n1164), .Z(G6) );
NOR2_X1 U843 ( .A1(n1148), .A2(n1165), .ZN(G57) );
XOR2_X1 U844 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U845 ( .A(KEYINPUT2), .B(n1168), .Z(n1167) );
NOR3_X1 U846 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1168) );
NOR3_X1 U847 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
INV_X1 U848 ( .A(n1175), .ZN(n1174) );
NOR2_X1 U849 ( .A1(n1176), .A2(n1175), .ZN(n1170) );
NAND2_X1 U850 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
XOR2_X1 U851 ( .A(n1179), .B(KEYINPUT61), .Z(n1177) );
INV_X1 U852 ( .A(n1180), .ZN(n1169) );
XOR2_X1 U853 ( .A(n1181), .B(n1182), .Z(n1166) );
AND2_X1 U854 ( .A1(G472), .A2(n1154), .ZN(n1182) );
NOR2_X1 U855 ( .A1(n1148), .A2(n1183), .ZN(G54) );
XOR2_X1 U856 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U857 ( .A1(KEYINPUT4), .A2(n1186), .ZN(n1185) );
XOR2_X1 U858 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U859 ( .A(G110), .B(n1189), .ZN(n1188) );
XOR2_X1 U860 ( .A(n1190), .B(n1191), .Z(n1187) );
NOR2_X1 U861 ( .A1(G140), .A2(KEYINPUT60), .ZN(n1191) );
NAND2_X1 U862 ( .A1(n1154), .A2(G469), .ZN(n1184) );
INV_X1 U863 ( .A(n1192), .ZN(n1154) );
NOR2_X1 U864 ( .A1(n1148), .A2(n1193), .ZN(G51) );
XOR2_X1 U865 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U866 ( .A1(n1106), .A2(n1192), .ZN(n1194) );
NAND2_X1 U867 ( .A1(G902), .A2(n1058), .ZN(n1192) );
NAND2_X1 U868 ( .A1(n1111), .A2(n1132), .ZN(n1058) );
AND4_X1 U869 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1132) );
AND4_X1 U870 ( .A1(n1200), .A2(n1201), .A3(n1164), .A4(n1053), .ZN(n1199) );
NAND3_X1 U871 ( .A1(n1074), .A2(n1066), .A3(n1202), .ZN(n1053) );
NAND3_X1 U872 ( .A1(n1202), .A2(n1066), .A3(n1073), .ZN(n1164) );
NAND2_X1 U873 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
XOR2_X1 U874 ( .A(KEYINPUT24), .B(n1075), .Z(n1204) );
NAND2_X1 U875 ( .A1(n1205), .A2(n1206), .ZN(n1196) );
NAND2_X1 U876 ( .A1(n1207), .A2(n1083), .ZN(n1206) );
XOR2_X1 U877 ( .A(n1084), .B(KEYINPUT18), .Z(n1207) );
AND4_X1 U878 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1111) );
NOR3_X1 U879 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
NOR2_X1 U880 ( .A1(n1215), .A2(n1216), .ZN(n1212) );
NOR2_X1 U881 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
XNOR2_X1 U882 ( .A(KEYINPUT37), .B(n1219), .ZN(n1218) );
NOR2_X1 U883 ( .A1(n1220), .A2(n1221), .ZN(n1217) );
NOR2_X1 U884 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
XOR2_X1 U885 ( .A(n1084), .B(KEYINPUT29), .Z(n1223) );
NOR2_X1 U886 ( .A1(n1060), .A2(G952), .ZN(n1148) );
XOR2_X1 U887 ( .A(G146), .B(n1214), .Z(G48) );
AND3_X1 U888 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1214) );
NAND3_X1 U889 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(G45) );
OR2_X1 U890 ( .A1(n1213), .A2(KEYINPUT53), .ZN(n1229) );
NAND3_X1 U891 ( .A1(KEYINPUT53), .A2(n1213), .A3(n1230), .ZN(n1228) );
NAND2_X1 U892 ( .A1(G143), .A2(n1231), .ZN(n1227) );
NAND2_X1 U893 ( .A1(n1232), .A2(KEYINPUT53), .ZN(n1231) );
XNOR2_X1 U894 ( .A(n1213), .B(KEYINPUT49), .ZN(n1232) );
AND3_X1 U895 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1213) );
NOR3_X1 U896 ( .A1(n1086), .A2(n1236), .A3(n1098), .ZN(n1235) );
INV_X1 U897 ( .A(n1225), .ZN(n1086) );
XOR2_X1 U898 ( .A(G140), .B(n1237), .Z(G42) );
NOR3_X1 U899 ( .A1(n1221), .A2(n1238), .A3(n1216), .ZN(n1237) );
XOR2_X1 U900 ( .A(n1083), .B(KEYINPUT25), .Z(n1238) );
INV_X1 U901 ( .A(n1222), .ZN(n1083) );
NAND2_X1 U902 ( .A1(n1239), .A2(n1240), .ZN(G39) );
NAND2_X1 U903 ( .A1(KEYINPUT22), .A2(G137), .ZN(n1240) );
XOR2_X1 U904 ( .A(n1241), .B(n1242), .Z(n1239) );
NOR2_X1 U905 ( .A1(n1216), .A2(n1219), .ZN(n1242) );
NAND3_X1 U906 ( .A1(n1233), .A2(n1224), .A3(n1075), .ZN(n1219) );
NOR2_X1 U907 ( .A1(G137), .A2(KEYINPUT22), .ZN(n1241) );
XOR2_X1 U908 ( .A(n1243), .B(n1210), .Z(G36) );
NAND4_X1 U909 ( .A1(n1068), .A2(n1233), .A3(n1074), .A4(n1234), .ZN(n1210) );
NAND2_X1 U910 ( .A1(n1244), .A2(n1245), .ZN(G33) );
NAND2_X1 U911 ( .A1(G131), .A2(n1246), .ZN(n1245) );
XOR2_X1 U912 ( .A(KEYINPUT16), .B(n1247), .Z(n1244) );
NOR2_X1 U913 ( .A1(G131), .A2(n1246), .ZN(n1247) );
NAND3_X1 U914 ( .A1(n1068), .A2(n1234), .A3(n1226), .ZN(n1246) );
INV_X1 U915 ( .A(n1221), .ZN(n1226) );
NAND2_X1 U916 ( .A1(n1233), .A2(n1073), .ZN(n1221) );
INV_X1 U917 ( .A(n1216), .ZN(n1068) );
NAND2_X1 U918 ( .A1(n1089), .A2(n1248), .ZN(n1216) );
XNOR2_X1 U919 ( .A(G128), .B(n1208), .ZN(G30) );
NAND4_X1 U920 ( .A1(n1233), .A2(n1224), .A3(n1074), .A4(n1225), .ZN(n1208) );
AND3_X1 U921 ( .A1(n1249), .A2(n1077), .A3(n1250), .ZN(n1233) );
XNOR2_X1 U922 ( .A(G101), .B(n1251), .ZN(G3) );
NAND2_X1 U923 ( .A1(n1205), .A2(n1234), .ZN(n1251) );
XOR2_X1 U924 ( .A(n1252), .B(n1209), .Z(G27) );
NAND4_X1 U925 ( .A1(n1222), .A2(n1073), .A3(n1253), .A4(n1071), .ZN(n1209) );
AND2_X1 U926 ( .A1(n1249), .A2(n1225), .ZN(n1253) );
NAND2_X1 U927 ( .A1(n1254), .A2(n1255), .ZN(n1249) );
NAND3_X1 U928 ( .A1(G902), .A2(n1063), .A3(n1114), .ZN(n1255) );
NOR2_X1 U929 ( .A1(n1060), .A2(G900), .ZN(n1114) );
XOR2_X1 U930 ( .A(n1256), .B(n1201), .Z(G24) );
NAND4_X1 U931 ( .A1(n1257), .A2(n1066), .A3(n1258), .A4(n1259), .ZN(n1201) );
NAND2_X1 U932 ( .A1(n1260), .A2(n1261), .ZN(n1066) );
OR2_X1 U933 ( .A1(n1084), .A2(KEYINPUT23), .ZN(n1261) );
NAND3_X1 U934 ( .A1(n1262), .A2(n1263), .A3(KEYINPUT23), .ZN(n1260) );
XOR2_X1 U935 ( .A(n1264), .B(n1265), .Z(G21) );
NAND2_X1 U936 ( .A1(n1203), .A2(n1075), .ZN(n1265) );
AND2_X1 U937 ( .A1(n1257), .A2(n1224), .ZN(n1203) );
NOR2_X1 U938 ( .A1(n1263), .A2(n1262), .ZN(n1224) );
XNOR2_X1 U939 ( .A(G116), .B(n1200), .ZN(G18) );
NAND3_X1 U940 ( .A1(n1074), .A2(n1234), .A3(n1257), .ZN(n1200) );
NOR2_X1 U941 ( .A1(n1259), .A2(n1098), .ZN(n1074) );
XOR2_X1 U942 ( .A(n1266), .B(n1198), .Z(G15) );
NAND3_X1 U943 ( .A1(n1073), .A2(n1234), .A3(n1257), .ZN(n1198) );
AND3_X1 U944 ( .A1(n1225), .A2(n1267), .A3(n1071), .ZN(n1257) );
AND2_X1 U945 ( .A1(n1078), .A2(n1077), .ZN(n1071) );
INV_X1 U946 ( .A(n1084), .ZN(n1234) );
NAND2_X1 U947 ( .A1(n1262), .A2(n1097), .ZN(n1084) );
NOR2_X1 U948 ( .A1(n1258), .A2(n1236), .ZN(n1073) );
XNOR2_X1 U949 ( .A(G110), .B(n1268), .ZN(G12) );
NAND2_X1 U950 ( .A1(n1205), .A2(n1222), .ZN(n1268) );
NOR2_X1 U951 ( .A1(n1097), .A2(n1262), .ZN(n1222) );
NOR2_X1 U952 ( .A1(n1269), .A2(n1095), .ZN(n1262) );
NOR2_X1 U953 ( .A1(n1270), .A2(n1155), .ZN(n1095) );
INV_X1 U954 ( .A(n1102), .ZN(n1155) );
NOR2_X1 U955 ( .A1(n1102), .A2(n1103), .ZN(n1269) );
INV_X1 U956 ( .A(n1270), .ZN(n1103) );
NAND2_X1 U957 ( .A1(n1153), .A2(n1271), .ZN(n1270) );
XOR2_X1 U958 ( .A(n1272), .B(n1273), .Z(n1153) );
XOR2_X1 U959 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U960 ( .A(G110), .B(n1276), .Z(n1275) );
NOR2_X1 U961 ( .A1(KEYINPUT50), .A2(n1277), .ZN(n1276) );
XOR2_X1 U962 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U963 ( .A(G146), .B(G125), .Z(n1279) );
NOR2_X1 U964 ( .A1(KEYINPUT7), .A2(n1280), .ZN(n1278) );
NOR2_X1 U965 ( .A1(n1281), .A2(n1282), .ZN(n1274) );
INV_X1 U966 ( .A(G221), .ZN(n1281) );
XOR2_X1 U967 ( .A(n1264), .B(n1283), .Z(n1272) );
XOR2_X1 U968 ( .A(G137), .B(G128), .Z(n1283) );
NAND2_X1 U969 ( .A1(G217), .A2(n1284), .ZN(n1102) );
INV_X1 U970 ( .A(n1263), .ZN(n1097) );
XOR2_X1 U971 ( .A(n1285), .B(G472), .Z(n1263) );
NAND2_X1 U972 ( .A1(n1286), .A2(n1271), .ZN(n1285) );
XOR2_X1 U973 ( .A(n1287), .B(n1288), .Z(n1286) );
INV_X1 U974 ( .A(n1181), .ZN(n1288) );
XOR2_X1 U975 ( .A(n1289), .B(G101), .Z(n1181) );
NAND2_X1 U976 ( .A1(n1290), .A2(G210), .ZN(n1289) );
XOR2_X1 U977 ( .A(n1291), .B(KEYINPUT21), .Z(n1287) );
NAND3_X1 U978 ( .A1(n1292), .A2(n1293), .A3(n1180), .ZN(n1291) );
NAND2_X1 U979 ( .A1(n1173), .A2(n1172), .ZN(n1180) );
NOR2_X1 U980 ( .A1(n1178), .A2(n1179), .ZN(n1173) );
NAND2_X1 U981 ( .A1(n1294), .A2(n1179), .ZN(n1293) );
XOR2_X1 U982 ( .A(n1176), .B(n1178), .Z(n1294) );
NAND3_X1 U983 ( .A1(n1176), .A2(n1178), .A3(n1295), .ZN(n1292) );
INV_X1 U984 ( .A(n1172), .ZN(n1176) );
XOR2_X1 U985 ( .A(n1296), .B(n1297), .Z(n1172) );
XOR2_X1 U986 ( .A(n1264), .B(n1298), .Z(n1297) );
NAND2_X1 U987 ( .A1(KEYINPUT40), .A2(n1299), .ZN(n1298) );
XOR2_X1 U988 ( .A(KEYINPUT3), .B(G116), .Z(n1299) );
INV_X1 U989 ( .A(G119), .ZN(n1264) );
NAND2_X1 U990 ( .A1(KEYINPUT48), .A2(n1266), .ZN(n1296) );
AND2_X1 U991 ( .A1(n1075), .A2(n1202), .ZN(n1205) );
AND4_X1 U992 ( .A1(n1225), .A2(n1250), .A3(n1077), .A4(n1267), .ZN(n1202) );
NAND2_X1 U993 ( .A1(n1300), .A2(n1254), .ZN(n1267) );
NAND3_X1 U994 ( .A1(n1063), .A2(n1060), .A3(n1301), .ZN(n1254) );
XOR2_X1 U995 ( .A(KEYINPUT17), .B(G952), .Z(n1301) );
XOR2_X1 U996 ( .A(n1302), .B(KEYINPUT55), .Z(n1300) );
NAND4_X1 U997 ( .A1(G953), .A2(G902), .A3(n1063), .A4(n1131), .ZN(n1302) );
INV_X1 U998 ( .A(G898), .ZN(n1131) );
NAND2_X1 U999 ( .A1(G237), .A2(G234), .ZN(n1063) );
NAND2_X1 U1000 ( .A1(G221), .A2(n1284), .ZN(n1077) );
NAND2_X1 U1001 ( .A1(G234), .A2(n1271), .ZN(n1284) );
INV_X1 U1002 ( .A(n1078), .ZN(n1250) );
XOR2_X1 U1003 ( .A(n1303), .B(G469), .Z(n1078) );
NAND2_X1 U1004 ( .A1(n1304), .A2(n1271), .ZN(n1303) );
XOR2_X1 U1005 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1006 ( .A(n1307), .B(KEYINPUT33), .ZN(n1306) );
NAND2_X1 U1007 ( .A1(n1308), .A2(KEYINPUT36), .ZN(n1307) );
XOR2_X1 U1008 ( .A(n1309), .B(n1310), .Z(n1308) );
NOR2_X1 U1009 ( .A1(KEYINPUT9), .A2(n1189), .ZN(n1310) );
NAND2_X1 U1010 ( .A1(G227), .A2(n1060), .ZN(n1189) );
XNOR2_X1 U1011 ( .A(G110), .B(n1311), .ZN(n1309) );
NOR2_X1 U1012 ( .A1(G140), .A2(KEYINPUT28), .ZN(n1311) );
INV_X1 U1013 ( .A(n1190), .ZN(n1305) );
XOR2_X1 U1014 ( .A(n1312), .B(n1313), .Z(n1190) );
XNOR2_X1 U1015 ( .A(n1123), .B(n1314), .ZN(n1313) );
XNOR2_X1 U1016 ( .A(n1315), .B(n1178), .ZN(n1314) );
XOR2_X1 U1017 ( .A(n1316), .B(n1317), .Z(n1178) );
NOR2_X1 U1018 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NOR2_X1 U1019 ( .A1(n1320), .A2(n1243), .ZN(n1319) );
NOR2_X1 U1020 ( .A1(KEYINPUT52), .A2(n1321), .ZN(n1320) );
NOR2_X1 U1021 ( .A1(KEYINPUT32), .A2(n1322), .ZN(n1321) );
INV_X1 U1022 ( .A(G137), .ZN(n1322) );
NOR2_X1 U1023 ( .A1(G137), .A2(n1323), .ZN(n1318) );
NOR2_X1 U1024 ( .A1(n1324), .A2(KEYINPUT32), .ZN(n1323) );
NOR2_X1 U1025 ( .A1(KEYINPUT52), .A2(G134), .ZN(n1324) );
NAND2_X1 U1026 ( .A1(KEYINPUT10), .A2(n1120), .ZN(n1316) );
XNOR2_X1 U1027 ( .A(n1325), .B(n1326), .ZN(n1123) );
XNOR2_X1 U1028 ( .A(G128), .B(KEYINPUT44), .ZN(n1325) );
XOR2_X1 U1029 ( .A(n1163), .B(n1327), .Z(n1312) );
XOR2_X1 U1030 ( .A(KEYINPUT38), .B(G107), .Z(n1327) );
NOR2_X1 U1031 ( .A1(n1089), .A2(n1088), .ZN(n1225) );
INV_X1 U1032 ( .A(n1248), .ZN(n1088) );
NAND2_X1 U1033 ( .A1(G214), .A2(n1328), .ZN(n1248) );
XNOR2_X1 U1034 ( .A(n1106), .B(n1329), .ZN(n1089) );
NOR2_X1 U1035 ( .A1(n1105), .A2(KEYINPUT39), .ZN(n1329) );
AND2_X1 U1036 ( .A1(n1330), .A2(n1271), .ZN(n1105) );
XOR2_X1 U1037 ( .A(KEYINPUT57), .B(n1195), .Z(n1330) );
XNOR2_X1 U1038 ( .A(n1331), .B(n1332), .ZN(n1195) );
XOR2_X1 U1039 ( .A(n1295), .B(n1136), .Z(n1332) );
XOR2_X1 U1040 ( .A(G110), .B(G122), .Z(n1136) );
INV_X1 U1041 ( .A(n1179), .ZN(n1295) );
XOR2_X1 U1042 ( .A(n1333), .B(n1326), .Z(n1179) );
XOR2_X1 U1043 ( .A(G146), .B(G143), .Z(n1326) );
XNOR2_X1 U1044 ( .A(KEYINPUT54), .B(n1334), .ZN(n1333) );
NOR2_X1 U1045 ( .A1(G128), .A2(KEYINPUT5), .ZN(n1334) );
XOR2_X1 U1046 ( .A(n1335), .B(n1336), .Z(n1331) );
NOR2_X1 U1047 ( .A1(G953), .A2(n1130), .ZN(n1336) );
INV_X1 U1048 ( .A(G224), .ZN(n1130) );
XOR2_X1 U1049 ( .A(n1337), .B(G125), .Z(n1335) );
NAND2_X1 U1050 ( .A1(KEYINPUT0), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1051 ( .A(n1339), .B(n1142), .Z(n1338) );
INV_X1 U1052 ( .A(n1147), .ZN(n1142) );
XOR2_X1 U1053 ( .A(n1340), .B(n1341), .Z(n1147) );
XOR2_X1 U1054 ( .A(KEYINPUT51), .B(G119), .Z(n1341) );
XOR2_X1 U1055 ( .A(n1266), .B(G116), .Z(n1340) );
NOR2_X1 U1056 ( .A1(KEYINPUT1), .A2(n1143), .ZN(n1339) );
INV_X1 U1057 ( .A(n1146), .ZN(n1143) );
NAND2_X1 U1058 ( .A1(n1342), .A2(n1343), .ZN(n1146) );
NAND2_X1 U1059 ( .A1(G107), .A2(n1344), .ZN(n1343) );
NAND2_X1 U1060 ( .A1(n1345), .A2(n1346), .ZN(n1342) );
XNOR2_X1 U1061 ( .A(KEYINPUT26), .B(n1344), .ZN(n1345) );
XOR2_X1 U1062 ( .A(G104), .B(n1315), .Z(n1344) );
XNOR2_X1 U1063 ( .A(G101), .B(KEYINPUT46), .ZN(n1315) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1328), .ZN(n1106) );
NAND2_X1 U1065 ( .A1(n1347), .A2(n1271), .ZN(n1328) );
INV_X1 U1066 ( .A(G902), .ZN(n1271) );
INV_X1 U1067 ( .A(G237), .ZN(n1347) );
NOR2_X1 U1068 ( .A1(n1258), .A2(n1259), .ZN(n1075) );
INV_X1 U1069 ( .A(n1236), .ZN(n1259) );
XOR2_X1 U1070 ( .A(n1348), .B(n1104), .Z(n1236) );
NOR2_X1 U1071 ( .A1(n1161), .A2(G902), .ZN(n1104) );
XOR2_X1 U1072 ( .A(n1349), .B(n1350), .Z(n1161) );
NOR2_X1 U1073 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XOR2_X1 U1074 ( .A(n1353), .B(KEYINPUT11), .Z(n1352) );
NAND2_X1 U1075 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NOR2_X1 U1076 ( .A1(n1355), .A2(n1354), .ZN(n1351) );
XNOR2_X1 U1077 ( .A(G146), .B(n1122), .ZN(n1354) );
XOR2_X1 U1078 ( .A(n1252), .B(n1280), .Z(n1122) );
INV_X1 U1079 ( .A(G140), .ZN(n1280) );
INV_X1 U1080 ( .A(G125), .ZN(n1252) );
AND2_X1 U1081 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1082 ( .A1(n1358), .A2(n1120), .ZN(n1357) );
XOR2_X1 U1083 ( .A(KEYINPUT42), .B(n1359), .Z(n1356) );
NOR2_X1 U1084 ( .A1(n1358), .A2(n1120), .ZN(n1359) );
INV_X1 U1085 ( .A(G131), .ZN(n1120) );
AND2_X1 U1086 ( .A1(n1360), .A2(n1361), .ZN(n1358) );
NAND2_X1 U1087 ( .A1(n1362), .A2(n1230), .ZN(n1361) );
INV_X1 U1088 ( .A(G143), .ZN(n1230) );
NAND2_X1 U1089 ( .A1(n1290), .A2(G214), .ZN(n1362) );
NAND3_X1 U1090 ( .A1(n1290), .A2(G214), .A3(G143), .ZN(n1360) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1290) );
NAND2_X1 U1092 ( .A1(n1363), .A2(n1364), .ZN(n1349) );
NAND2_X1 U1093 ( .A1(n1365), .A2(n1163), .ZN(n1364) );
XOR2_X1 U1094 ( .A(KEYINPUT27), .B(n1366), .Z(n1363) );
NOR2_X1 U1095 ( .A1(n1163), .A2(n1365), .ZN(n1366) );
XOR2_X1 U1096 ( .A(n1266), .B(n1367), .Z(n1365) );
NAND2_X1 U1097 ( .A1(KEYINPUT45), .A2(n1256), .ZN(n1367) );
INV_X1 U1098 ( .A(G122), .ZN(n1256) );
INV_X1 U1099 ( .A(G113), .ZN(n1266) );
INV_X1 U1100 ( .A(G104), .ZN(n1163) );
NAND2_X1 U1101 ( .A1(KEYINPUT47), .A2(G475), .ZN(n1348) );
INV_X1 U1102 ( .A(n1098), .ZN(n1258) );
XOR2_X1 U1103 ( .A(n1368), .B(G478), .Z(n1098) );
NAND2_X1 U1104 ( .A1(n1158), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1105 ( .A(KEYINPUT62), .B(G902), .Z(n1369) );
XOR2_X1 U1106 ( .A(n1370), .B(n1371), .Z(n1158) );
XOR2_X1 U1107 ( .A(n1372), .B(n1373), .Z(n1371) );
NOR2_X1 U1108 ( .A1(n1282), .A2(n1374), .ZN(n1373) );
INV_X1 U1109 ( .A(G217), .ZN(n1374) );
NAND2_X1 U1110 ( .A1(G234), .A2(n1060), .ZN(n1282) );
INV_X1 U1111 ( .A(G953), .ZN(n1060) );
NOR2_X1 U1112 ( .A1(KEYINPUT59), .A2(n1375), .ZN(n1372) );
XOR2_X1 U1113 ( .A(n1243), .B(n1376), .Z(n1375) );
NOR2_X1 U1114 ( .A1(KEYINPUT63), .A2(n1377), .ZN(n1376) );
XOR2_X1 U1115 ( .A(G143), .B(G128), .Z(n1377) );
INV_X1 U1116 ( .A(G134), .ZN(n1243) );
XOR2_X1 U1117 ( .A(n1346), .B(n1378), .Z(n1370) );
XOR2_X1 U1118 ( .A(G122), .B(G116), .Z(n1378) );
INV_X1 U1119 ( .A(G107), .ZN(n1346) );
endmodule


