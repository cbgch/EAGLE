//Key = 0110011011011000010100000110101101101110001101000010000100110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324;

XNOR2_X1 U733 ( .A(G107), .B(n1018), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR2_X1 U735 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND4_X1 U736 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
NAND2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XOR2_X1 U738 ( .A(KEYINPUT13), .B(n1029), .Z(n1028) );
NAND2_X1 U739 ( .A1(n1030), .A2(n1031), .ZN(n1025) );
NAND2_X1 U740 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U741 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
XNOR2_X1 U742 ( .A(n1036), .B(KEYINPUT26), .ZN(n1034) );
NAND2_X1 U743 ( .A1(n1037), .A2(n1036), .ZN(n1032) );
NAND4_X1 U744 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1021) );
NAND4_X1 U745 ( .A1(n1042), .A2(n1043), .A3(n1036), .A4(n1044), .ZN(n1039) );
NAND3_X1 U746 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NAND2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XNOR2_X1 U748 ( .A(n1050), .B(n1051), .ZN(n1048) );
NOR2_X1 U749 ( .A1(KEYINPUT60), .A2(n1052), .ZN(n1051) );
NAND3_X1 U750 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1045) );
NAND3_X1 U751 ( .A1(n1056), .A2(n1057), .A3(n1029), .ZN(n1038) );
AND2_X1 U752 ( .A1(n1030), .A2(n1043), .ZN(n1029) );
AND3_X1 U753 ( .A1(n1049), .A2(n1053), .A3(n1042), .ZN(n1030) );
INV_X1 U754 ( .A(n1058), .ZN(n1042) );
NOR3_X1 U755 ( .A1(n1059), .A2(G953), .A3(G952), .ZN(n1019) );
INV_X1 U756 ( .A(n1040), .ZN(n1059) );
NAND4_X1 U757 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1040) );
NOR4_X1 U758 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
XOR2_X1 U759 ( .A(G469), .B(n1068), .Z(n1067) );
XOR2_X1 U760 ( .A(KEYINPUT32), .B(n1069), .Z(n1066) );
NOR2_X1 U761 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR3_X1 U762 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1062) );
NAND2_X1 U763 ( .A1(n1070), .A2(n1071), .ZN(n1061) );
XOR2_X1 U764 ( .A(G472), .B(n1075), .Z(n1060) );
NOR2_X1 U765 ( .A1(n1076), .A2(KEYINPUT24), .ZN(n1075) );
XOR2_X1 U766 ( .A(n1077), .B(n1078), .Z(G72) );
XOR2_X1 U767 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U768 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U769 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U770 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U771 ( .A1(KEYINPUT44), .A2(n1087), .ZN(n1085) );
XOR2_X1 U772 ( .A(n1088), .B(n1089), .Z(n1083) );
XNOR2_X1 U773 ( .A(n1090), .B(G125), .ZN(n1089) );
NAND2_X1 U774 ( .A1(KEYINPUT19), .A2(n1091), .ZN(n1088) );
NOR2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1081) );
NAND2_X1 U776 ( .A1(n1041), .A2(n1094), .ZN(n1079) );
NAND2_X1 U777 ( .A1(G953), .A2(n1095), .ZN(n1077) );
NAND2_X1 U778 ( .A1(G900), .A2(G227), .ZN(n1095) );
XOR2_X1 U779 ( .A(n1096), .B(n1097), .Z(G69) );
XOR2_X1 U780 ( .A(n1098), .B(n1099), .Z(n1097) );
OR2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U782 ( .A1(G953), .A2(n1102), .ZN(n1098) );
NAND2_X1 U783 ( .A1(G898), .A2(G224), .ZN(n1102) );
NOR2_X1 U784 ( .A1(n1023), .A2(G953), .ZN(n1096) );
NOR2_X1 U785 ( .A1(n1103), .A2(n1104), .ZN(G66) );
XOR2_X1 U786 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U787 ( .A1(KEYINPUT3), .A2(n1107), .ZN(n1106) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1070), .ZN(n1105) );
NOR2_X1 U789 ( .A1(n1103), .A2(n1109), .ZN(G63) );
XNOR2_X1 U790 ( .A(n1110), .B(n1111), .ZN(n1109) );
AND2_X1 U791 ( .A1(G478), .A2(n1108), .ZN(n1111) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1112), .ZN(G60) );
XNOR2_X1 U793 ( .A(n1113), .B(n1114), .ZN(n1112) );
NAND3_X1 U794 ( .A1(n1115), .A2(n1116), .A3(G475), .ZN(n1113) );
XNOR2_X1 U795 ( .A(KEYINPUT7), .B(n1117), .ZN(n1115) );
XOR2_X1 U796 ( .A(G104), .B(n1118), .Z(G6) );
NOR2_X1 U797 ( .A1(n1103), .A2(n1119), .ZN(G57) );
XOR2_X1 U798 ( .A(n1120), .B(n1121), .Z(n1119) );
XOR2_X1 U799 ( .A(n1122), .B(n1123), .Z(n1121) );
AND2_X1 U800 ( .A1(G472), .A2(n1108), .ZN(n1123) );
NOR2_X1 U801 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
XOR2_X1 U802 ( .A(KEYINPUT10), .B(n1126), .Z(n1125) );
NOR2_X1 U803 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
AND2_X1 U804 ( .A1(n1128), .A2(n1127), .ZN(n1124) );
XOR2_X1 U805 ( .A(n1129), .B(G116), .Z(n1127) );
XOR2_X1 U806 ( .A(n1130), .B(n1131), .Z(n1128) );
NAND2_X1 U807 ( .A1(KEYINPUT11), .A2(n1132), .ZN(n1120) );
XNOR2_X1 U808 ( .A(G101), .B(n1133), .ZN(n1132) );
NOR2_X1 U809 ( .A1(n1103), .A2(n1134), .ZN(G54) );
XOR2_X1 U810 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U811 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U812 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U813 ( .A1(KEYINPUT14), .A2(n1141), .ZN(n1140) );
AND2_X1 U814 ( .A1(G469), .A2(n1108), .ZN(n1139) );
XNOR2_X1 U815 ( .A(G110), .B(n1142), .ZN(n1135) );
XNOR2_X1 U816 ( .A(KEYINPUT45), .B(KEYINPUT31), .ZN(n1142) );
NOR2_X1 U817 ( .A1(n1103), .A2(n1143), .ZN(G51) );
XNOR2_X1 U818 ( .A(n1144), .B(n1145), .ZN(n1143) );
XNOR2_X1 U819 ( .A(n1146), .B(n1147), .ZN(n1145) );
NOR2_X1 U820 ( .A1(KEYINPUT35), .A2(n1148), .ZN(n1147) );
NOR3_X1 U821 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
AND3_X1 U823 ( .A1(n1153), .A2(n1154), .A3(n1152), .ZN(n1150) );
INV_X1 U824 ( .A(KEYINPUT23), .ZN(n1153) );
NAND2_X1 U825 ( .A1(KEYINPUT50), .A2(n1155), .ZN(n1146) );
NAND2_X1 U826 ( .A1(n1108), .A2(n1156), .ZN(n1155) );
AND2_X1 U827 ( .A1(G902), .A2(n1116), .ZN(n1108) );
NAND2_X1 U828 ( .A1(n1023), .A2(n1024), .ZN(n1116) );
INV_X1 U829 ( .A(n1094), .ZN(n1024) );
NAND4_X1 U830 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1094) );
AND4_X1 U831 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
NAND2_X1 U832 ( .A1(n1027), .A2(n1165), .ZN(n1164) );
NOR2_X1 U833 ( .A1(n1166), .A2(n1167), .ZN(n1159) );
AND4_X1 U834 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1023) );
NOR4_X1 U835 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
INV_X1 U836 ( .A(n1176), .ZN(n1175) );
INV_X1 U837 ( .A(n1018), .ZN(n1172) );
NAND3_X1 U838 ( .A1(n1035), .A2(n1049), .A3(n1177), .ZN(n1018) );
NOR2_X1 U839 ( .A1(n1178), .A2(n1118), .ZN(n1170) );
AND3_X1 U840 ( .A1(n1177), .A2(n1049), .A3(n1037), .ZN(n1118) );
AND3_X1 U841 ( .A1(n1037), .A2(n1179), .A3(n1180), .ZN(n1178) );
NOR2_X1 U842 ( .A1(n1041), .A2(G952), .ZN(n1103) );
XOR2_X1 U843 ( .A(n1157), .B(n1181), .Z(G48) );
NAND2_X1 U844 ( .A1(KEYINPUT25), .A2(G146), .ZN(n1181) );
NAND4_X1 U845 ( .A1(n1182), .A2(n1037), .A3(n1055), .A4(n1027), .ZN(n1157) );
XNOR2_X1 U846 ( .A(G143), .B(n1158), .ZN(G45) );
NAND3_X1 U847 ( .A1(n1182), .A2(n1027), .A3(n1183), .ZN(n1158) );
AND3_X1 U848 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1183) );
XOR2_X1 U849 ( .A(G140), .B(n1167), .Z(G42) );
AND3_X1 U850 ( .A1(n1036), .A2(n1187), .A3(n1188), .ZN(n1167) );
XOR2_X1 U851 ( .A(G137), .B(n1189), .Z(G39) );
NOR2_X1 U852 ( .A1(KEYINPUT56), .A2(n1163), .ZN(n1189) );
NAND3_X1 U853 ( .A1(n1190), .A2(n1036), .A3(n1182), .ZN(n1163) );
XNOR2_X1 U854 ( .A(G134), .B(n1162), .ZN(G36) );
NAND2_X1 U855 ( .A1(n1191), .A2(n1035), .ZN(n1162) );
NAND2_X1 U856 ( .A1(n1192), .A2(n1193), .ZN(G33) );
NAND2_X1 U857 ( .A1(n1194), .A2(n1161), .ZN(n1193) );
XOR2_X1 U858 ( .A(KEYINPUT53), .B(n1195), .Z(n1194) );
XOR2_X1 U859 ( .A(KEYINPUT33), .B(n1196), .Z(n1192) );
NOR2_X1 U860 ( .A1(n1161), .A2(n1197), .ZN(n1196) );
XOR2_X1 U861 ( .A(KEYINPUT61), .B(n1195), .Z(n1197) );
XOR2_X1 U862 ( .A(G131), .B(KEYINPUT63), .Z(n1195) );
NAND2_X1 U863 ( .A1(n1191), .A2(n1037), .ZN(n1161) );
AND3_X1 U864 ( .A1(n1036), .A2(n1186), .A3(n1182), .ZN(n1191) );
INV_X1 U865 ( .A(n1064), .ZN(n1036) );
NAND2_X1 U866 ( .A1(n1056), .A2(n1198), .ZN(n1064) );
XNOR2_X1 U867 ( .A(G128), .B(n1199), .ZN(G30) );
NAND2_X1 U868 ( .A1(n1200), .A2(n1027), .ZN(n1199) );
XNOR2_X1 U869 ( .A(n1165), .B(KEYINPUT62), .ZN(n1200) );
AND3_X1 U870 ( .A1(n1055), .A2(n1035), .A3(n1182), .ZN(n1165) );
AND3_X1 U871 ( .A1(n1187), .A2(n1201), .A3(n1202), .ZN(n1182) );
XNOR2_X1 U872 ( .A(G101), .B(n1168), .ZN(G3) );
NAND4_X1 U873 ( .A1(n1202), .A2(n1043), .A3(n1177), .A4(n1186), .ZN(n1168) );
XOR2_X1 U874 ( .A(G125), .B(n1166), .Z(G27) );
AND3_X1 U875 ( .A1(n1027), .A2(n1053), .A3(n1188), .ZN(n1166) );
AND4_X1 U876 ( .A1(n1055), .A2(n1037), .A3(n1054), .A4(n1201), .ZN(n1188) );
NAND2_X1 U877 ( .A1(n1058), .A2(n1203), .ZN(n1201) );
NAND4_X1 U878 ( .A1(n1204), .A2(G902), .A3(n1205), .A4(n1206), .ZN(n1203) );
INV_X1 U879 ( .A(n1093), .ZN(n1205) );
XOR2_X1 U880 ( .A(n1092), .B(KEYINPUT12), .Z(n1204) );
XNOR2_X1 U881 ( .A(G900), .B(KEYINPUT9), .ZN(n1092) );
XNOR2_X1 U882 ( .A(G122), .B(n1169), .ZN(G24) );
NAND4_X1 U883 ( .A1(n1053), .A2(n1185), .A3(n1184), .A4(n1207), .ZN(n1169) );
AND2_X1 U884 ( .A1(n1179), .A2(n1049), .ZN(n1207) );
NOR2_X1 U885 ( .A1(n1202), .A2(n1055), .ZN(n1049) );
XOR2_X1 U886 ( .A(n1065), .B(KEYINPUT46), .Z(n1184) );
NAND2_X1 U887 ( .A1(n1208), .A2(n1209), .ZN(G21) );
NAND2_X1 U888 ( .A1(G119), .A2(n1176), .ZN(n1209) );
XOR2_X1 U889 ( .A(KEYINPUT58), .B(n1210), .Z(n1208) );
NOR2_X1 U890 ( .A1(G119), .A2(n1176), .ZN(n1210) );
NAND4_X1 U891 ( .A1(n1202), .A2(n1190), .A3(n1179), .A4(n1053), .ZN(n1176) );
XOR2_X1 U892 ( .A(G116), .B(n1174), .Z(G18) );
AND3_X1 U893 ( .A1(n1035), .A2(n1179), .A3(n1180), .ZN(n1174) );
NOR2_X1 U894 ( .A1(n1185), .A2(n1211), .ZN(n1035) );
INV_X1 U895 ( .A(n1065), .ZN(n1211) );
XNOR2_X1 U896 ( .A(G113), .B(n1212), .ZN(G15) );
NAND4_X1 U897 ( .A1(n1213), .A2(n1037), .A3(n1180), .A4(n1027), .ZN(n1212) );
INV_X1 U898 ( .A(n1046), .ZN(n1180) );
NAND3_X1 U899 ( .A1(n1053), .A2(n1186), .A3(n1202), .ZN(n1046) );
INV_X1 U900 ( .A(n1054), .ZN(n1202) );
NAND2_X1 U901 ( .A1(n1214), .A2(n1215), .ZN(n1053) );
OR3_X1 U902 ( .A1(n1216), .A2(n1074), .A3(KEYINPUT60), .ZN(n1215) );
INV_X1 U903 ( .A(n1050), .ZN(n1216) );
NAND2_X1 U904 ( .A1(KEYINPUT60), .A2(n1187), .ZN(n1214) );
NOR2_X1 U905 ( .A1(n1065), .A2(n1217), .ZN(n1037) );
XOR2_X1 U906 ( .A(n1218), .B(KEYINPUT16), .Z(n1213) );
XNOR2_X1 U907 ( .A(n1219), .B(n1173), .ZN(G12) );
AND3_X1 U908 ( .A1(n1177), .A2(n1054), .A3(n1190), .ZN(n1173) );
AND2_X1 U909 ( .A1(n1043), .A2(n1055), .ZN(n1190) );
INV_X1 U910 ( .A(n1186), .ZN(n1055) );
XNOR2_X1 U911 ( .A(n1071), .B(n1220), .ZN(n1186) );
NOR2_X1 U912 ( .A1(n1070), .A2(KEYINPUT54), .ZN(n1220) );
AND2_X1 U913 ( .A1(G217), .A2(n1221), .ZN(n1070) );
OR2_X1 U914 ( .A1(n1107), .A2(G902), .ZN(n1071) );
XNOR2_X1 U915 ( .A(n1222), .B(n1223), .ZN(n1107) );
XOR2_X1 U916 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U917 ( .A(n1226), .B(n1227), .ZN(n1225) );
NOR2_X1 U918 ( .A1(KEYINPUT47), .A2(n1228), .ZN(n1227) );
XOR2_X1 U919 ( .A(n1229), .B(KEYINPUT2), .Z(n1228) );
NOR2_X1 U920 ( .A1(KEYINPUT15), .A2(n1230), .ZN(n1226) );
NOR2_X1 U921 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NOR2_X1 U922 ( .A1(n1233), .A2(n1219), .ZN(n1232) );
NOR2_X1 U923 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NOR2_X1 U924 ( .A1(n1236), .A2(n1237), .ZN(n1234) );
NOR2_X1 U925 ( .A1(n1238), .A2(n1239), .ZN(n1231) );
INV_X1 U926 ( .A(n1237), .ZN(n1239) );
XNOR2_X1 U927 ( .A(G119), .B(n1240), .ZN(n1237) );
NOR2_X1 U928 ( .A1(n1241), .A2(n1236), .ZN(n1238) );
INV_X1 U929 ( .A(KEYINPUT5), .ZN(n1236) );
NOR2_X1 U930 ( .A1(G110), .A2(n1235), .ZN(n1241) );
INV_X1 U931 ( .A(KEYINPUT59), .ZN(n1235) );
NAND2_X1 U932 ( .A1(n1242), .A2(G221), .ZN(n1224) );
XNOR2_X1 U933 ( .A(G137), .B(n1243), .ZN(n1222) );
XNOR2_X1 U934 ( .A(KEYINPUT36), .B(n1244), .ZN(n1243) );
NOR2_X1 U935 ( .A1(n1065), .A2(n1185), .ZN(n1043) );
INV_X1 U936 ( .A(n1217), .ZN(n1185) );
NOR2_X1 U937 ( .A1(n1245), .A2(n1073), .ZN(n1217) );
NOR3_X1 U938 ( .A1(G475), .A2(G902), .A3(n1114), .ZN(n1073) );
XOR2_X1 U939 ( .A(n1072), .B(KEYINPUT20), .Z(n1245) );
AND2_X1 U940 ( .A1(G475), .A2(n1246), .ZN(n1072) );
OR2_X1 U941 ( .A1(n1114), .A2(G902), .ZN(n1246) );
XNOR2_X1 U942 ( .A(n1247), .B(n1248), .ZN(n1114) );
XNOR2_X1 U943 ( .A(n1249), .B(n1250), .ZN(n1248) );
INV_X1 U944 ( .A(n1251), .ZN(n1250) );
NOR2_X1 U945 ( .A1(KEYINPUT57), .A2(n1229), .ZN(n1249) );
XOR2_X1 U946 ( .A(G125), .B(n1087), .Z(n1229) );
XNOR2_X1 U947 ( .A(n1252), .B(n1244), .ZN(n1247) );
NAND3_X1 U948 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1252) );
NAND2_X1 U949 ( .A1(KEYINPUT27), .A2(n1256), .ZN(n1255) );
NAND3_X1 U950 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1254) );
INV_X1 U951 ( .A(KEYINPUT27), .ZN(n1258) );
OR2_X1 U952 ( .A1(n1259), .A2(n1257), .ZN(n1253) );
NOR2_X1 U953 ( .A1(KEYINPUT22), .A2(n1256), .ZN(n1257) );
XNOR2_X1 U954 ( .A(n1260), .B(G143), .ZN(n1256) );
NAND2_X1 U955 ( .A1(n1261), .A2(G214), .ZN(n1260) );
XNOR2_X1 U956 ( .A(n1262), .B(G478), .ZN(n1065) );
NAND2_X1 U957 ( .A1(n1110), .A2(n1117), .ZN(n1262) );
XNOR2_X1 U958 ( .A(n1263), .B(n1264), .ZN(n1110) );
NOR2_X1 U959 ( .A1(KEYINPUT41), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U960 ( .A(n1266), .B(n1267), .ZN(n1265) );
XOR2_X1 U961 ( .A(G122), .B(G116), .Z(n1267) );
XOR2_X1 U962 ( .A(n1268), .B(n1269), .Z(n1263) );
AND2_X1 U963 ( .A1(n1242), .A2(G217), .ZN(n1269) );
AND2_X1 U964 ( .A1(G234), .A2(n1041), .ZN(n1242) );
NAND3_X1 U965 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1268) );
NAND2_X1 U966 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U967 ( .A1(KEYINPUT55), .A2(n1275), .ZN(n1274) );
XNOR2_X1 U968 ( .A(KEYINPUT1), .B(n1090), .ZN(n1273) );
NAND4_X1 U969 ( .A1(n1276), .A2(KEYINPUT55), .A3(KEYINPUT37), .A4(n1275), .ZN(n1271) );
XNOR2_X1 U970 ( .A(KEYINPUT1), .B(G134), .ZN(n1276) );
OR2_X1 U971 ( .A1(n1275), .A2(KEYINPUT37), .ZN(n1270) );
XNOR2_X1 U972 ( .A(n1240), .B(n1277), .ZN(n1275) );
INV_X1 U973 ( .A(G128), .ZN(n1240) );
XOR2_X1 U974 ( .A(n1076), .B(n1278), .Z(n1054) );
XOR2_X1 U975 ( .A(KEYINPUT42), .B(G472), .Z(n1278) );
AND2_X1 U976 ( .A1(n1279), .A2(n1117), .ZN(n1076) );
XOR2_X1 U977 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U978 ( .A(n1129), .B(n1282), .Z(n1281) );
XNOR2_X1 U979 ( .A(G113), .B(n1283), .ZN(n1129) );
XNOR2_X1 U980 ( .A(KEYINPUT28), .B(n1284), .ZN(n1283) );
XOR2_X1 U981 ( .A(n1130), .B(n1285), .Z(n1280) );
XNOR2_X1 U982 ( .A(n1286), .B(n1287), .ZN(n1285) );
NOR2_X1 U983 ( .A1(KEYINPUT49), .A2(n1133), .ZN(n1287) );
NAND2_X1 U984 ( .A1(n1261), .A2(G210), .ZN(n1133) );
AND2_X1 U985 ( .A1(n1288), .A2(n1041), .ZN(n1261) );
XNOR2_X1 U986 ( .A(G237), .B(KEYINPUT0), .ZN(n1288) );
NAND2_X1 U987 ( .A1(KEYINPUT38), .A2(n1131), .ZN(n1286) );
INV_X1 U988 ( .A(n1141), .ZN(n1131) );
AND2_X1 U989 ( .A1(n1179), .A2(n1187), .ZN(n1177) );
NOR2_X1 U990 ( .A1(n1050), .A2(n1074), .ZN(n1187) );
INV_X1 U991 ( .A(n1052), .ZN(n1074) );
NAND2_X1 U992 ( .A1(G221), .A2(n1221), .ZN(n1052) );
NAND2_X1 U993 ( .A1(G234), .A2(n1117), .ZN(n1221) );
XOR2_X1 U994 ( .A(G469), .B(n1289), .Z(n1050) );
NOR2_X1 U995 ( .A1(n1068), .A2(KEYINPUT4), .ZN(n1289) );
AND2_X1 U996 ( .A1(n1290), .A2(n1117), .ZN(n1068) );
XOR2_X1 U997 ( .A(n1291), .B(n1137), .Z(n1290) );
XNOR2_X1 U998 ( .A(n1292), .B(n1293), .ZN(n1137) );
XOR2_X1 U999 ( .A(n1087), .B(n1091), .Z(n1293) );
XOR2_X1 U1000 ( .A(n1294), .B(n1295), .Z(n1091) );
XNOR2_X1 U1001 ( .A(n1277), .B(n1296), .ZN(n1295) );
NOR2_X1 U1002 ( .A1(KEYINPUT39), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U1003 ( .A(KEYINPUT51), .B(n1244), .ZN(n1297) );
INV_X1 U1004 ( .A(G146), .ZN(n1244) );
INV_X1 U1005 ( .A(G143), .ZN(n1277) );
XNOR2_X1 U1006 ( .A(G140), .B(KEYINPUT34), .ZN(n1087) );
XOR2_X1 U1007 ( .A(n1298), .B(n1299), .Z(n1292) );
AND2_X1 U1008 ( .A1(n1041), .A2(G227), .ZN(n1299) );
NAND3_X1 U1009 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1298) );
NAND2_X1 U1010 ( .A1(KEYINPUT52), .A2(n1303), .ZN(n1302) );
OR3_X1 U1011 ( .A1(n1304), .A2(KEYINPUT52), .A3(G101), .ZN(n1301) );
NAND2_X1 U1012 ( .A1(G101), .A2(n1304), .ZN(n1300) );
NAND2_X1 U1013 ( .A1(KEYINPUT8), .A2(n1305), .ZN(n1304) );
INV_X1 U1014 ( .A(n1303), .ZN(n1305) );
XOR2_X1 U1015 ( .A(G104), .B(n1266), .Z(n1303) );
INV_X1 U1016 ( .A(G107), .ZN(n1266) );
XNOR2_X1 U1017 ( .A(n1141), .B(n1306), .ZN(n1291) );
NOR2_X1 U1018 ( .A1(G110), .A2(KEYINPUT29), .ZN(n1306) );
XNOR2_X1 U1019 ( .A(n1307), .B(n1086), .ZN(n1141) );
XNOR2_X1 U1020 ( .A(G137), .B(n1259), .ZN(n1086) );
XNOR2_X1 U1021 ( .A(G131), .B(KEYINPUT21), .ZN(n1259) );
NAND2_X1 U1022 ( .A1(KEYINPUT43), .A2(n1090), .ZN(n1307) );
INV_X1 U1023 ( .A(G134), .ZN(n1090) );
AND2_X1 U1024 ( .A1(n1027), .A2(n1218), .ZN(n1179) );
NAND2_X1 U1025 ( .A1(n1058), .A2(n1308), .ZN(n1218) );
NAND3_X1 U1026 ( .A1(n1101), .A2(n1206), .A3(G902), .ZN(n1308) );
NOR2_X1 U1027 ( .A1(n1093), .A2(G898), .ZN(n1101) );
XOR2_X1 U1028 ( .A(G953), .B(KEYINPUT17), .Z(n1093) );
NAND3_X1 U1029 ( .A1(n1206), .A2(n1041), .A3(G952), .ZN(n1058) );
NAND2_X1 U1030 ( .A1(G237), .A2(G234), .ZN(n1206) );
NOR2_X1 U1031 ( .A1(n1056), .A2(n1057), .ZN(n1027) );
INV_X1 U1032 ( .A(n1198), .ZN(n1057) );
NAND2_X1 U1033 ( .A1(G214), .A2(n1309), .ZN(n1198) );
XNOR2_X1 U1034 ( .A(n1156), .B(n1310), .ZN(n1056) );
NOR2_X1 U1035 ( .A1(G902), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U1036 ( .A(n1312), .B(n1100), .ZN(n1311) );
INV_X1 U1037 ( .A(n1144), .ZN(n1100) );
XNOR2_X1 U1038 ( .A(n1313), .B(n1314), .ZN(n1144) );
XOR2_X1 U1039 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1040 ( .A(G107), .B(G110), .ZN(n1316) );
NAND2_X1 U1041 ( .A1(KEYINPUT30), .A2(n1284), .ZN(n1315) );
INV_X1 U1042 ( .A(G119), .ZN(n1284) );
XNOR2_X1 U1043 ( .A(n1251), .B(n1282), .ZN(n1313) );
XOR2_X1 U1044 ( .A(G101), .B(G116), .Z(n1282) );
XOR2_X1 U1045 ( .A(G104), .B(n1317), .Z(n1251) );
XOR2_X1 U1046 ( .A(G122), .B(G113), .Z(n1317) );
NAND2_X1 U1047 ( .A1(n1318), .A2(n1319), .ZN(n1312) );
NAND2_X1 U1048 ( .A1(n1152), .A2(n1154), .ZN(n1319) );
INV_X1 U1049 ( .A(n1149), .ZN(n1318) );
NOR2_X1 U1050 ( .A1(n1154), .A2(n1152), .ZN(n1149) );
XOR2_X1 U1051 ( .A(n1130), .B(G125), .Z(n1152) );
XOR2_X1 U1052 ( .A(n1294), .B(n1320), .Z(n1130) );
NOR2_X1 U1053 ( .A1(KEYINPUT40), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1054 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1055 ( .A(G146), .B(KEYINPUT48), .ZN(n1323) );
NAND2_X1 U1056 ( .A1(KEYINPUT6), .A2(G143), .ZN(n1322) );
XNOR2_X1 U1057 ( .A(G128), .B(KEYINPUT18), .ZN(n1294) );
NAND2_X1 U1058 ( .A1(G224), .A2(n1041), .ZN(n1154) );
INV_X1 U1059 ( .A(G953), .ZN(n1041) );
AND2_X1 U1060 ( .A1(G210), .A2(n1309), .ZN(n1156) );
NAND2_X1 U1061 ( .A1(n1324), .A2(n1117), .ZN(n1309) );
INV_X1 U1062 ( .A(G902), .ZN(n1117) );
INV_X1 U1063 ( .A(G237), .ZN(n1324) );
INV_X1 U1064 ( .A(G110), .ZN(n1219) );
endmodule


