//Key = 1010001100000111010111000000011011011111010011010000011101010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U739 ( .A(G107), .B(n1017), .ZN(G9) );
NOR2_X1 U740 ( .A1(n1018), .A2(n1019), .ZN(G75) );
XOR2_X1 U741 ( .A(KEYINPUT4), .B(n1020), .Z(n1019) );
NOR3_X1 U742 ( .A1(n1021), .A2(G953), .A3(G952), .ZN(n1020) );
INV_X1 U743 ( .A(n1022), .ZN(n1021) );
NOR2_X1 U744 ( .A1(n1023), .A2(n1024), .ZN(n1018) );
NAND4_X1 U745 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
XOR2_X1 U746 ( .A(n1029), .B(KEYINPUT27), .Z(n1025) );
NAND2_X1 U747 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U748 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U749 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1032) );
NAND2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND4_X1 U752 ( .A1(n1041), .A2(n1034), .A3(n1042), .A4(n1043), .ZN(n1040) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1048), .A2(n1049), .ZN(n1042) );
NAND3_X1 U756 ( .A1(n1050), .A2(n1036), .A3(n1051), .ZN(n1039) );
NAND4_X1 U757 ( .A1(G952), .A2(n1052), .A3(n1053), .A4(n1022), .ZN(n1023) );
NAND4_X1 U758 ( .A1(n1041), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1022) );
NOR4_X1 U759 ( .A1(n1057), .A2(n1058), .A3(n1051), .A4(n1059), .ZN(n1056) );
NOR3_X1 U760 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1058) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
AND3_X1 U762 ( .A1(n1064), .A2(n1065), .A3(n1063), .ZN(n1061) );
NOR2_X1 U763 ( .A1(n1066), .A2(KEYINPUT23), .ZN(n1063) );
INV_X1 U764 ( .A(n1067), .ZN(n1066) );
NOR2_X1 U765 ( .A1(n1067), .A2(n1065), .ZN(n1060) );
INV_X1 U766 ( .A(KEYINPUT42), .ZN(n1065) );
NAND3_X1 U767 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1057) );
NOR3_X1 U768 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1055) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1072) );
NOR2_X1 U771 ( .A1(G902), .A2(n1078), .ZN(n1076) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(n1071) );
NOR2_X1 U773 ( .A1(n1081), .A2(KEYINPUT5), .ZN(n1080) );
INV_X1 U774 ( .A(n1082), .ZN(n1081) );
XOR2_X1 U775 ( .A(KEYINPUT54), .B(n1083), .Z(n1054) );
AND2_X1 U776 ( .A1(n1075), .A2(n1074), .ZN(n1083) );
NAND2_X1 U777 ( .A1(n1030), .A2(n1084), .ZN(n1053) );
NAND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND4_X1 U779 ( .A1(n1037), .A2(n1034), .A3(n1044), .A4(n1087), .ZN(n1086) );
NAND2_X1 U780 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U781 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U782 ( .A1(n1036), .A2(n1092), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U784 ( .A1(n1034), .A2(n1095), .ZN(n1094) );
NAND2_X1 U785 ( .A1(n1037), .A2(n1096), .ZN(n1093) );
INV_X1 U786 ( .A(n1097), .ZN(n1030) );
XNOR2_X1 U787 ( .A(KEYINPUT29), .B(n1098), .ZN(n1052) );
XOR2_X1 U788 ( .A(n1099), .B(n1100), .Z(G72) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND4_X1 U790 ( .A1(n1103), .A2(n1026), .A3(n1104), .A4(n1105), .ZN(n1102) );
XOR2_X1 U791 ( .A(n1106), .B(n1107), .Z(n1103) );
NAND3_X1 U792 ( .A1(n1108), .A2(n1098), .A3(n1109), .ZN(n1101) );
XNOR2_X1 U793 ( .A(n1107), .B(n1106), .ZN(n1109) );
NAND2_X1 U794 ( .A1(n1026), .A2(n1104), .ZN(n1108) );
NAND2_X1 U795 ( .A1(n1105), .A2(n1110), .ZN(n1099) );
NAND2_X1 U796 ( .A1(G953), .A2(n1111), .ZN(n1110) );
INV_X1 U797 ( .A(n1112), .ZN(n1105) );
NAND2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(G69) );
NAND3_X1 U799 ( .A1(n1115), .A2(n1116), .A3(G953), .ZN(n1114) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1115) );
NAND2_X1 U801 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
OR2_X1 U802 ( .A1(n1098), .A2(G224), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1116), .B(n1119), .Z(n1117) );
NAND2_X1 U804 ( .A1(KEYINPUT44), .A2(n1120), .ZN(n1119) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1116) );
NAND2_X1 U806 ( .A1(G953), .A2(n1123), .ZN(n1122) );
XOR2_X1 U807 ( .A(n1124), .B(n1125), .Z(n1121) );
NAND2_X1 U808 ( .A1(KEYINPUT41), .A2(n1126), .ZN(n1124) );
NOR2_X1 U809 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U811 ( .A1(n1082), .A2(n1131), .ZN(n1130) );
NOR2_X1 U812 ( .A1(n1127), .A2(n1132), .ZN(G63) );
XOR2_X1 U813 ( .A(KEYINPUT28), .B(n1133), .Z(n1132) );
NOR3_X1 U814 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
INV_X1 U816 ( .A(n1139), .ZN(n1138) );
NOR2_X1 U817 ( .A1(KEYINPUT49), .A2(n1140), .ZN(n1137) );
XNOR2_X1 U818 ( .A(n1141), .B(KEYINPUT24), .ZN(n1140) );
NOR3_X1 U819 ( .A1(n1139), .A2(KEYINPUT49), .A3(n1078), .ZN(n1135) );
NOR2_X1 U820 ( .A1(n1131), .A2(n1077), .ZN(n1139) );
AND2_X1 U821 ( .A1(n1078), .A2(KEYINPUT49), .ZN(n1134) );
INV_X1 U822 ( .A(n1141), .ZN(n1078) );
NOR2_X1 U823 ( .A1(n1127), .A2(n1142), .ZN(G60) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR3_X1 U825 ( .A1(n1131), .A2(KEYINPUT58), .A3(n1075), .ZN(n1143) );
XNOR2_X1 U826 ( .A(G104), .B(n1145), .ZN(G6) );
NAND2_X1 U827 ( .A1(n1146), .A2(n1096), .ZN(n1145) );
XOR2_X1 U828 ( .A(n1147), .B(KEYINPUT57), .Z(n1146) );
NOR2_X1 U829 ( .A1(n1127), .A2(n1148), .ZN(G57) );
XOR2_X1 U830 ( .A(n1149), .B(n1150), .Z(n1148) );
XNOR2_X1 U831 ( .A(n1151), .B(n1152), .ZN(n1150) );
NOR2_X1 U832 ( .A1(n1153), .A2(n1131), .ZN(n1151) );
NOR2_X1 U833 ( .A1(n1154), .A2(n1155), .ZN(n1149) );
AND2_X1 U834 ( .A1(KEYINPUT31), .A2(n1156), .ZN(n1155) );
NOR2_X1 U835 ( .A1(KEYINPUT10), .A2(n1156), .ZN(n1154) );
NAND3_X1 U836 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
OR2_X1 U837 ( .A1(G101), .A2(KEYINPUT30), .ZN(n1158) );
NAND2_X1 U838 ( .A1(n1160), .A2(KEYINPUT30), .ZN(n1157) );
NOR2_X1 U839 ( .A1(n1127), .A2(n1161), .ZN(G54) );
XOR2_X1 U840 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U841 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U842 ( .A1(n1166), .A2(n1131), .ZN(n1165) );
NOR2_X1 U843 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
XOR2_X1 U844 ( .A(KEYINPUT25), .B(n1169), .Z(n1168) );
NOR2_X1 U845 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
AND2_X1 U846 ( .A1(n1170), .A2(n1171), .ZN(n1167) );
XOR2_X1 U847 ( .A(n1172), .B(G110), .Z(n1171) );
NAND2_X1 U848 ( .A1(n1173), .A2(KEYINPUT33), .ZN(n1172) );
XNOR2_X1 U849 ( .A(G140), .B(KEYINPUT32), .ZN(n1173) );
NOR2_X1 U850 ( .A1(n1127), .A2(n1174), .ZN(G51) );
XOR2_X1 U851 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR3_X1 U852 ( .A1(n1177), .A2(KEYINPUT22), .A3(n1178), .ZN(n1176) );
NOR2_X1 U853 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U854 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
INV_X1 U855 ( .A(KEYINPUT47), .ZN(n1182) );
AND2_X1 U856 ( .A1(n1183), .A2(KEYINPUT20), .ZN(n1181) );
NOR2_X1 U857 ( .A1(n1184), .A2(n1183), .ZN(n1177) );
XOR2_X1 U858 ( .A(n1125), .B(n1185), .Z(n1183) );
XNOR2_X1 U859 ( .A(G110), .B(G122), .ZN(n1125) );
NOR2_X1 U860 ( .A1(n1186), .A2(n1187), .ZN(n1184) );
INV_X1 U861 ( .A(KEYINPUT20), .ZN(n1187) );
AND2_X1 U862 ( .A1(KEYINPUT47), .A2(n1180), .ZN(n1186) );
XOR2_X1 U863 ( .A(n1188), .B(n1189), .Z(n1180) );
XOR2_X1 U864 ( .A(KEYINPUT61), .B(G146), .Z(n1189) );
OR2_X1 U865 ( .A1(n1131), .A2(n1067), .ZN(n1175) );
NAND2_X1 U866 ( .A1(n1190), .A2(n1191), .ZN(n1131) );
NAND3_X1 U867 ( .A1(n1027), .A2(n1028), .A3(n1026), .ZN(n1191) );
AND4_X1 U868 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1026) );
INV_X1 U869 ( .A(n1120), .ZN(n1028) );
NAND4_X1 U870 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1120) );
NOR4_X1 U871 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NOR2_X1 U872 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NOR2_X1 U873 ( .A1(n1017), .A2(n1206), .ZN(n1205) );
NAND3_X1 U874 ( .A1(n1035), .A2(n1207), .A3(n1096), .ZN(n1017) );
NAND4_X1 U875 ( .A1(n1207), .A2(n1206), .A3(n1035), .A4(n1208), .ZN(n1197) );
INV_X1 U876 ( .A(KEYINPUT35), .ZN(n1206) );
NAND2_X1 U877 ( .A1(n1096), .A2(n1209), .ZN(n1196) );
NAND2_X1 U878 ( .A1(n1210), .A2(n1147), .ZN(n1209) );
NAND2_X1 U879 ( .A1(n1095), .A2(n1207), .ZN(n1147) );
NOR3_X1 U880 ( .A1(n1048), .A2(n1211), .A3(n1088), .ZN(n1207) );
XNOR2_X1 U881 ( .A(n1104), .B(KEYINPUT53), .ZN(n1027) );
AND4_X1 U882 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1104) );
XNOR2_X1 U883 ( .A(KEYINPUT16), .B(n1216), .ZN(n1190) );
NOR2_X1 U884 ( .A1(n1098), .A2(G952), .ZN(n1127) );
XNOR2_X1 U885 ( .A(G146), .B(n1212), .ZN(G48) );
NAND3_X1 U886 ( .A1(n1095), .A2(n1096), .A3(n1217), .ZN(n1212) );
NAND3_X1 U887 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(G45) );
NAND2_X1 U888 ( .A1(KEYINPUT48), .A2(n1213), .ZN(n1220) );
OR3_X1 U889 ( .A1(n1213), .A2(KEYINPUT48), .A3(G143), .ZN(n1219) );
NAND2_X1 U890 ( .A1(G143), .A2(n1221), .ZN(n1218) );
NAND2_X1 U891 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
INV_X1 U892 ( .A(KEYINPUT48), .ZN(n1223) );
XOR2_X1 U893 ( .A(n1213), .B(KEYINPUT45), .Z(n1222) );
NAND4_X1 U894 ( .A1(n1224), .A2(n1096), .A3(n1225), .A4(n1226), .ZN(n1213) );
XNOR2_X1 U895 ( .A(G140), .B(n1214), .ZN(G42) );
NAND3_X1 U896 ( .A1(n1227), .A2(n1228), .A3(n1034), .ZN(n1214) );
XOR2_X1 U897 ( .A(G137), .B(n1229), .Z(G39) );
NOR2_X1 U898 ( .A1(KEYINPUT63), .A2(n1215), .ZN(n1229) );
NAND3_X1 U899 ( .A1(n1034), .A2(n1217), .A3(n1037), .ZN(n1215) );
XNOR2_X1 U900 ( .A(G134), .B(n1192), .ZN(G36) );
NAND3_X1 U901 ( .A1(n1224), .A2(n1035), .A3(n1034), .ZN(n1192) );
XNOR2_X1 U902 ( .A(n1230), .B(n1193), .ZN(G33) );
NAND3_X1 U903 ( .A1(n1224), .A2(n1095), .A3(n1034), .ZN(n1193) );
NOR2_X1 U904 ( .A1(n1231), .A2(n1051), .ZN(n1034) );
AND4_X1 U905 ( .A1(n1228), .A2(n1044), .A3(n1091), .A4(n1232), .ZN(n1224) );
XNOR2_X1 U906 ( .A(G131), .B(KEYINPUT7), .ZN(n1230) );
XNOR2_X1 U907 ( .A(G128), .B(n1233), .ZN(G30) );
NAND2_X1 U908 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
INV_X1 U909 ( .A(n1194), .ZN(n1235) );
NAND3_X1 U910 ( .A1(n1096), .A2(n1035), .A3(n1217), .ZN(n1194) );
AND4_X1 U911 ( .A1(n1048), .A2(n1228), .A3(n1091), .A4(n1232), .ZN(n1217) );
XNOR2_X1 U912 ( .A(KEYINPUT8), .B(KEYINPUT52), .ZN(n1234) );
XNOR2_X1 U913 ( .A(n1204), .B(n1236), .ZN(G3) );
NAND2_X1 U914 ( .A1(KEYINPUT38), .A2(G101), .ZN(n1236) );
AND3_X1 U915 ( .A1(n1037), .A2(n1228), .A3(n1237), .ZN(n1204) );
XNOR2_X1 U916 ( .A(G125), .B(n1195), .ZN(G27) );
NAND3_X1 U917 ( .A1(n1227), .A2(n1096), .A3(n1090), .ZN(n1195) );
AND4_X1 U918 ( .A1(n1048), .A2(n1095), .A3(n1041), .A4(n1232), .ZN(n1227) );
NAND2_X1 U919 ( .A1(n1097), .A2(n1238), .ZN(n1232) );
NAND3_X1 U920 ( .A1(G902), .A2(n1239), .A3(n1112), .ZN(n1238) );
NOR2_X1 U921 ( .A1(G900), .A2(n1098), .ZN(n1112) );
XOR2_X1 U922 ( .A(G122), .B(n1203), .Z(G24) );
AND3_X1 U923 ( .A1(n1036), .A2(n1096), .A3(n1240), .ZN(n1203) );
NOR3_X1 U924 ( .A1(n1241), .A2(n1242), .A3(n1211), .ZN(n1240) );
NOR3_X1 U925 ( .A1(n1091), .A2(n1048), .A3(n1049), .ZN(n1036) );
XNOR2_X1 U926 ( .A(n1243), .B(n1244), .ZN(G21) );
NOR2_X1 U927 ( .A1(n1245), .A2(n1208), .ZN(n1244) );
XOR2_X1 U928 ( .A(n1210), .B(KEYINPUT12), .Z(n1245) );
OR3_X1 U929 ( .A1(n1049), .A2(n1041), .A3(n1246), .ZN(n1210) );
XNOR2_X1 U930 ( .A(G116), .B(n1247), .ZN(G18) );
NAND2_X1 U931 ( .A1(KEYINPUT13), .A2(n1202), .ZN(n1247) );
AND3_X1 U932 ( .A1(n1090), .A2(n1035), .A3(n1237), .ZN(n1202) );
NOR2_X1 U933 ( .A1(n1225), .A2(n1242), .ZN(n1035) );
INV_X1 U934 ( .A(n1226), .ZN(n1242) );
XOR2_X1 U935 ( .A(G113), .B(n1201), .Z(G15) );
AND3_X1 U936 ( .A1(n1090), .A2(n1095), .A3(n1237), .ZN(n1201) );
NOR4_X1 U937 ( .A1(n1208), .A2(n1048), .A3(n1041), .A4(n1211), .ZN(n1237) );
INV_X1 U938 ( .A(n1248), .ZN(n1211) );
NOR2_X1 U939 ( .A1(n1226), .A2(n1241), .ZN(n1095) );
INV_X1 U940 ( .A(n1049), .ZN(n1090) );
NAND2_X1 U941 ( .A1(n1047), .A2(n1069), .ZN(n1049) );
XOR2_X1 U942 ( .A(n1200), .B(n1249), .Z(G12) );
NOR2_X1 U943 ( .A1(KEYINPUT46), .A2(n1250), .ZN(n1249) );
NOR3_X1 U944 ( .A1(n1208), .A2(n1088), .A3(n1246), .ZN(n1200) );
NAND3_X1 U945 ( .A1(n1048), .A2(n1248), .A3(n1037), .ZN(n1246) );
NOR2_X1 U946 ( .A1(n1226), .A2(n1225), .ZN(n1037) );
INV_X1 U947 ( .A(n1241), .ZN(n1225) );
XOR2_X1 U948 ( .A(n1074), .B(n1075), .Z(n1241) );
INV_X1 U949 ( .A(G475), .ZN(n1075) );
NOR2_X1 U950 ( .A1(n1144), .A2(n1251), .ZN(n1074) );
XNOR2_X1 U951 ( .A(KEYINPUT2), .B(G902), .ZN(n1251) );
XNOR2_X1 U952 ( .A(n1252), .B(n1253), .ZN(n1144) );
XOR2_X1 U953 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U954 ( .A(G104), .B(n1256), .Z(n1255) );
AND3_X1 U955 ( .A1(n1257), .A2(n1258), .A3(G214), .ZN(n1256) );
INV_X1 U956 ( .A(KEYINPUT3), .ZN(n1258) );
XOR2_X1 U957 ( .A(G143), .B(G122), .Z(n1254) );
XNOR2_X1 U958 ( .A(n1259), .B(n1260), .ZN(n1252) );
XNOR2_X1 U959 ( .A(n1261), .B(n1262), .ZN(n1260) );
NOR2_X1 U960 ( .A1(KEYINPUT51), .A2(n1263), .ZN(n1262) );
NAND2_X1 U961 ( .A1(KEYINPUT59), .A2(n1107), .ZN(n1261) );
NAND2_X1 U962 ( .A1(n1264), .A2(n1068), .ZN(n1226) );
NAND3_X1 U963 ( .A1(n1077), .A2(n1216), .A3(n1141), .ZN(n1068) );
INV_X1 U964 ( .A(G478), .ZN(n1077) );
NAND2_X1 U965 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U966 ( .A1(n1141), .A2(n1216), .ZN(n1266) );
XNOR2_X1 U967 ( .A(n1267), .B(n1268), .ZN(n1141) );
XOR2_X1 U968 ( .A(n1269), .B(n1270), .Z(n1268) );
NAND2_X1 U969 ( .A1(G217), .A2(n1271), .ZN(n1270) );
NAND2_X1 U970 ( .A1(n1272), .A2(n1273), .ZN(n1269) );
NAND2_X1 U971 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U972 ( .A(KEYINPUT36), .B(n1276), .Z(n1272) );
NOR2_X1 U973 ( .A1(n1274), .A2(n1275), .ZN(n1276) );
INV_X1 U974 ( .A(G134), .ZN(n1275) );
XOR2_X1 U975 ( .A(G143), .B(n1277), .Z(n1274) );
NOR2_X1 U976 ( .A1(G128), .A2(KEYINPUT26), .ZN(n1277) );
XOR2_X1 U977 ( .A(n1278), .B(n1279), .Z(n1267) );
XOR2_X1 U978 ( .A(G122), .B(G116), .Z(n1279) );
NAND2_X1 U979 ( .A1(KEYINPUT17), .A2(G107), .ZN(n1278) );
XNOR2_X1 U980 ( .A(G478), .B(KEYINPUT0), .ZN(n1265) );
NAND2_X1 U981 ( .A1(n1097), .A2(n1280), .ZN(n1248) );
NAND4_X1 U982 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1123), .ZN(n1280) );
INV_X1 U983 ( .A(G898), .ZN(n1123) );
NAND3_X1 U984 ( .A1(n1239), .A2(n1098), .A3(G952), .ZN(n1097) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1239) );
INV_X1 U986 ( .A(n1044), .ZN(n1048) );
XOR2_X1 U987 ( .A(n1281), .B(n1082), .Z(n1044) );
NAND2_X1 U988 ( .A1(G217), .A2(n1282), .ZN(n1082) );
NAND2_X1 U989 ( .A1(KEYINPUT21), .A2(n1079), .ZN(n1281) );
NAND2_X1 U990 ( .A1(n1129), .A2(n1216), .ZN(n1079) );
XNOR2_X1 U991 ( .A(n1283), .B(n1284), .ZN(n1129) );
XNOR2_X1 U992 ( .A(n1107), .B(n1285), .ZN(n1284) );
XOR2_X1 U993 ( .A(n1286), .B(n1287), .Z(n1285) );
NAND2_X1 U994 ( .A1(G221), .A2(n1271), .ZN(n1286) );
AND2_X1 U995 ( .A1(G234), .A2(n1098), .ZN(n1271) );
XOR2_X1 U996 ( .A(G140), .B(n1288), .Z(n1107) );
XOR2_X1 U997 ( .A(n1289), .B(n1290), .Z(n1283) );
NOR2_X1 U998 ( .A1(KEYINPUT9), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U999 ( .A(G128), .B(n1292), .ZN(n1291) );
NOR2_X1 U1000 ( .A1(KEYINPUT1), .A2(n1243), .ZN(n1292) );
XNOR2_X1 U1001 ( .A(G137), .B(KEYINPUT56), .ZN(n1289) );
NAND2_X1 U1002 ( .A1(n1228), .A2(n1041), .ZN(n1088) );
INV_X1 U1003 ( .A(n1091), .ZN(n1041) );
XOR2_X1 U1004 ( .A(n1293), .B(n1153), .Z(n1091) );
INV_X1 U1005 ( .A(G472), .ZN(n1153) );
NAND3_X1 U1006 ( .A1(n1294), .A2(n1295), .A3(n1216), .ZN(n1293) );
NAND2_X1 U1007 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
INV_X1 U1008 ( .A(KEYINPUT11), .ZN(n1297) );
XNOR2_X1 U1009 ( .A(n1298), .B(n1299), .ZN(n1296) );
NOR2_X1 U1010 ( .A1(KEYINPUT34), .A2(n1152), .ZN(n1299) );
NAND3_X1 U1011 ( .A1(n1298), .A2(n1152), .A3(KEYINPUT11), .ZN(n1294) );
XOR2_X1 U1012 ( .A(n1300), .B(n1301), .Z(n1152) );
XNOR2_X1 U1013 ( .A(n1243), .B(G116), .ZN(n1301) );
XNOR2_X1 U1014 ( .A(n1302), .B(n1263), .ZN(n1300) );
INV_X1 U1015 ( .A(n1303), .ZN(n1263) );
AND2_X1 U1016 ( .A1(n1304), .A2(n1159), .ZN(n1298) );
NAND2_X1 U1017 ( .A1(n1305), .A2(n1306), .ZN(n1159) );
NAND2_X1 U1018 ( .A1(n1257), .A2(G210), .ZN(n1306) );
INV_X1 U1019 ( .A(G101), .ZN(n1305) );
XOR2_X1 U1020 ( .A(KEYINPUT55), .B(n1160), .Z(n1304) );
AND3_X1 U1021 ( .A1(G210), .A2(G101), .A3(n1257), .ZN(n1160) );
NOR2_X1 U1022 ( .A1(G237), .A2(G953), .ZN(n1257) );
NOR2_X1 U1023 ( .A1(n1047), .A2(n1046), .ZN(n1228) );
INV_X1 U1024 ( .A(n1069), .ZN(n1046) );
NAND2_X1 U1025 ( .A1(G221), .A2(n1282), .ZN(n1069) );
NAND2_X1 U1026 ( .A1(n1307), .A2(G234), .ZN(n1282) );
XNOR2_X1 U1027 ( .A(G902), .B(KEYINPUT60), .ZN(n1307) );
AND2_X1 U1028 ( .A1(n1308), .A2(n1070), .ZN(n1047) );
NAND3_X1 U1029 ( .A1(n1166), .A2(n1216), .A3(n1309), .ZN(n1070) );
INV_X1 U1030 ( .A(G469), .ZN(n1166) );
XOR2_X1 U1031 ( .A(KEYINPUT37), .B(n1059), .Z(n1308) );
AND2_X1 U1032 ( .A1(G469), .A2(n1310), .ZN(n1059) );
NAND2_X1 U1033 ( .A1(n1309), .A2(n1216), .ZN(n1310) );
XNOR2_X1 U1034 ( .A(n1311), .B(n1312), .ZN(n1309) );
XNOR2_X1 U1035 ( .A(n1313), .B(G110), .ZN(n1312) );
INV_X1 U1036 ( .A(G140), .ZN(n1313) );
XNOR2_X1 U1037 ( .A(n1162), .B(n1170), .ZN(n1311) );
NOR2_X1 U1038 ( .A1(n1111), .A2(G953), .ZN(n1170) );
INV_X1 U1039 ( .A(G227), .ZN(n1111) );
XNOR2_X1 U1040 ( .A(n1314), .B(n1315), .ZN(n1162) );
XOR2_X1 U1041 ( .A(n1302), .B(n1316), .Z(n1314) );
NOR2_X1 U1042 ( .A1(G101), .A2(KEYINPUT18), .ZN(n1316) );
XOR2_X1 U1043 ( .A(n1106), .B(n1317), .Z(n1302) );
XOR2_X1 U1044 ( .A(KEYINPUT50), .B(KEYINPUT15), .Z(n1317) );
XOR2_X1 U1045 ( .A(n1318), .B(n1319), .Z(n1106) );
XOR2_X1 U1046 ( .A(n1320), .B(n1259), .Z(n1319) );
XOR2_X1 U1047 ( .A(G131), .B(G146), .Z(n1259) );
XNOR2_X1 U1048 ( .A(G137), .B(G134), .ZN(n1318) );
INV_X1 U1049 ( .A(n1096), .ZN(n1208) );
NOR2_X1 U1050 ( .A1(n1050), .A2(n1051), .ZN(n1096) );
AND2_X1 U1051 ( .A1(G214), .A2(n1321), .ZN(n1051) );
INV_X1 U1052 ( .A(n1231), .ZN(n1050) );
XOR2_X1 U1053 ( .A(n1064), .B(n1067), .Z(n1231) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1321), .ZN(n1067) );
NAND2_X1 U1055 ( .A1(n1322), .A2(n1216), .ZN(n1321) );
INV_X1 U1056 ( .A(G237), .ZN(n1322) );
NAND2_X1 U1057 ( .A1(n1323), .A2(n1216), .ZN(n1064) );
INV_X1 U1058 ( .A(G902), .ZN(n1216) );
XOR2_X1 U1059 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U1060 ( .A(G122), .B(n1287), .Z(n1325) );
XNOR2_X1 U1061 ( .A(n1250), .B(G146), .ZN(n1287) );
INV_X1 U1062 ( .A(G110), .ZN(n1250) );
XOR2_X1 U1063 ( .A(n1188), .B(n1185), .Z(n1324) );
XOR2_X1 U1064 ( .A(n1126), .B(KEYINPUT43), .Z(n1185) );
XOR2_X1 U1065 ( .A(n1315), .B(n1326), .Z(n1126) );
XNOR2_X1 U1066 ( .A(G101), .B(n1327), .ZN(n1326) );
NAND3_X1 U1067 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1327) );
NAND2_X1 U1068 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
INV_X1 U1069 ( .A(KEYINPUT6), .ZN(n1332) );
NAND3_X1 U1070 ( .A1(KEYINPUT6), .A2(n1333), .A3(n1334), .ZN(n1329) );
OR2_X1 U1071 ( .A1(n1334), .A2(n1333), .ZN(n1328) );
NOR2_X1 U1072 ( .A1(n1335), .A2(n1331), .ZN(n1333) );
XOR2_X1 U1073 ( .A(n1303), .B(KEYINPUT39), .Z(n1331) );
XOR2_X1 U1074 ( .A(G113), .B(KEYINPUT62), .Z(n1303) );
INV_X1 U1075 ( .A(KEYINPUT19), .ZN(n1335) );
NAND2_X1 U1076 ( .A1(n1336), .A2(n1337), .ZN(n1334) );
NAND2_X1 U1077 ( .A1(G116), .A2(n1243), .ZN(n1337) );
XOR2_X1 U1078 ( .A(KEYINPUT14), .B(n1338), .Z(n1336) );
NOR2_X1 U1079 ( .A1(G116), .A2(n1243), .ZN(n1338) );
INV_X1 U1080 ( .A(G119), .ZN(n1243) );
XOR2_X1 U1081 ( .A(G104), .B(G107), .Z(n1315) );
XOR2_X1 U1082 ( .A(n1339), .B(n1320), .Z(n1188) );
XNOR2_X1 U1083 ( .A(n1340), .B(G143), .ZN(n1320) );
INV_X1 U1084 ( .A(G128), .ZN(n1340) );
XOR2_X1 U1085 ( .A(n1341), .B(n1288), .Z(n1339) );
XOR2_X1 U1086 ( .A(G125), .B(KEYINPUT40), .Z(n1288) );
NAND2_X1 U1087 ( .A1(G224), .A2(n1098), .ZN(n1341) );
INV_X1 U1088 ( .A(G953), .ZN(n1098) );
endmodule


