//Key = 0111011011011000011101000011001001111111010010100100010000110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343;

XNOR2_X1 U734 ( .A(G107), .B(n1014), .ZN(G9) );
NAND3_X1 U735 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(G75) );
NAND2_X1 U736 ( .A1(G952), .A2(n1018), .ZN(n1017) );
NAND4_X1 U737 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NOR4_X1 U738 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n1022) );
NOR4_X1 U739 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1024) );
NAND3_X1 U740 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1028) );
NOR2_X1 U741 ( .A1(n1034), .A2(n1035), .ZN(n1023) );
NOR3_X1 U742 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1034) );
NOR2_X1 U743 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
INV_X1 U744 ( .A(n1041), .ZN(n1039) );
NOR3_X1 U745 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1037) );
NOR2_X1 U746 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U747 ( .A1(n1047), .A2(n1029), .ZN(n1046) );
NOR2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U749 ( .A(KEYINPUT32), .B(n1050), .Z(n1049) );
NOR2_X1 U750 ( .A1(n1030), .A2(n1032), .ZN(n1048) );
INV_X1 U751 ( .A(KEYINPUT39), .ZN(n1032) );
NOR2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1045) );
NOR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
XOR2_X1 U755 ( .A(KEYINPUT43), .B(n1057), .Z(n1036) );
NOR2_X1 U756 ( .A1(n1058), .A2(n1040), .ZN(n1057) );
NAND2_X1 U757 ( .A1(n1059), .A2(n1060), .ZN(n1021) );
XOR2_X1 U758 ( .A(KEYINPUT57), .B(n1061), .Z(n1060) );
NAND3_X1 U759 ( .A1(n1062), .A2(n1061), .A3(n1063), .ZN(n1019) );
NOR2_X1 U760 ( .A1(n1040), .A2(n1042), .ZN(n1061) );
NAND3_X1 U761 ( .A1(n1064), .A2(n1031), .A3(n1065), .ZN(n1040) );
NAND4_X1 U762 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1015) );
NOR4_X1 U763 ( .A1(n1070), .A2(n1071), .A3(n1035), .A4(n1072), .ZN(n1069) );
NOR2_X1 U764 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
INV_X1 U765 ( .A(n1056), .ZN(n1070) );
NOR2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1068) );
XOR2_X1 U767 ( .A(KEYINPUT14), .B(n1055), .Z(n1076) );
XOR2_X1 U768 ( .A(KEYINPUT56), .B(n1077), .Z(n1075) );
NOR2_X1 U769 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U770 ( .A(n1080), .B(n1081), .Z(n1067) );
XOR2_X1 U771 ( .A(n1082), .B(KEYINPUT48), .Z(n1066) );
XOR2_X1 U772 ( .A(n1083), .B(n1084), .Z(G72) );
NOR2_X1 U773 ( .A1(n1085), .A2(n1016), .ZN(n1084) );
AND2_X1 U774 ( .A1(G227), .A2(G900), .ZN(n1085) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1083) );
NAND2_X1 U776 ( .A1(n1088), .A2(n1016), .ZN(n1087) );
XNOR2_X1 U777 ( .A(n1025), .B(n1089), .ZN(n1088) );
OR3_X1 U778 ( .A1(n1090), .A2(n1089), .A3(n1016), .ZN(n1086) );
XNOR2_X1 U779 ( .A(n1091), .B(n1092), .ZN(n1089) );
XOR2_X1 U780 ( .A(G131), .B(n1093), .Z(n1092) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1091) );
XOR2_X1 U782 ( .A(n1096), .B(n1097), .Z(G69) );
XOR2_X1 U783 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U785 ( .A1(G953), .A2(n1102), .ZN(n1101) );
XOR2_X1 U786 ( .A(n1103), .B(KEYINPUT7), .Z(n1100) );
NAND2_X1 U787 ( .A1(n1016), .A2(n1104), .ZN(n1098) );
NAND2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U789 ( .A(KEYINPUT38), .B(n1020), .ZN(n1106) );
NOR2_X1 U790 ( .A1(n1107), .A2(n1016), .ZN(n1096) );
NOR2_X1 U791 ( .A1(n1108), .A2(n1102), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1109), .A2(n1110), .ZN(G66) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U794 ( .A1(KEYINPUT50), .A2(n1113), .ZN(n1112) );
NAND2_X1 U795 ( .A1(n1114), .A2(n1078), .ZN(n1111) );
INV_X1 U796 ( .A(n1074), .ZN(n1078) );
NOR2_X1 U797 ( .A1(n1109), .A2(n1115), .ZN(G63) );
XNOR2_X1 U798 ( .A(n1116), .B(n1117), .ZN(n1115) );
AND2_X1 U799 ( .A1(G478), .A2(n1114), .ZN(n1117) );
NOR2_X1 U800 ( .A1(n1109), .A2(n1118), .ZN(G60) );
NOR3_X1 U801 ( .A1(n1080), .A2(n1119), .A3(n1120), .ZN(n1118) );
AND3_X1 U802 ( .A1(n1121), .A2(G475), .A3(n1114), .ZN(n1120) );
NOR2_X1 U803 ( .A1(n1122), .A2(n1121), .ZN(n1119) );
NOR2_X1 U804 ( .A1(n1123), .A2(n1081), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(G6) );
NAND2_X1 U806 ( .A1(G104), .A2(n1126), .ZN(n1125) );
XOR2_X1 U807 ( .A(KEYINPUT27), .B(n1127), .Z(n1124) );
NOR2_X1 U808 ( .A1(G104), .A2(n1126), .ZN(n1127) );
NAND3_X1 U809 ( .A1(n1128), .A2(n1033), .A3(n1129), .ZN(n1126) );
NOR2_X1 U810 ( .A1(n1109), .A2(n1130), .ZN(G57) );
XOR2_X1 U811 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U812 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U813 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U814 ( .A1(KEYINPUT23), .A2(n1137), .ZN(n1136) );
AND2_X1 U815 ( .A1(G472), .A2(n1114), .ZN(n1135) );
XOR2_X1 U816 ( .A(n1138), .B(n1139), .Z(n1131) );
NOR2_X1 U817 ( .A1(n1109), .A2(n1140), .ZN(G54) );
XOR2_X1 U818 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U819 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U820 ( .A(n1145), .B(n1146), .ZN(n1143) );
AND2_X1 U821 ( .A1(G469), .A2(n1114), .ZN(n1146) );
XOR2_X1 U822 ( .A(n1147), .B(n1148), .Z(n1141) );
XNOR2_X1 U823 ( .A(KEYINPUT53), .B(n1149), .ZN(n1148) );
NAND2_X1 U824 ( .A1(KEYINPUT37), .A2(n1150), .ZN(n1147) );
NOR2_X1 U825 ( .A1(n1109), .A2(n1151), .ZN(G51) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U827 ( .A(n1154), .B(n1103), .Z(n1153) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1152) );
XNOR2_X1 U829 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR3_X1 U830 ( .A1(n1159), .A2(KEYINPUT15), .A3(n1160), .ZN(n1158) );
INV_X1 U831 ( .A(n1114), .ZN(n1159) );
NOR2_X1 U832 ( .A1(n1161), .A2(n1123), .ZN(n1114) );
AND3_X1 U833 ( .A1(n1105), .A2(n1020), .A3(n1162), .ZN(n1123) );
XOR2_X1 U834 ( .A(n1025), .B(KEYINPUT30), .Z(n1162) );
NAND4_X1 U835 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1025) );
AND4_X1 U836 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
NOR2_X1 U837 ( .A1(n1171), .A2(n1172), .ZN(n1165) );
NOR2_X1 U838 ( .A1(n1035), .A2(n1173), .ZN(n1172) );
NOR3_X1 U839 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1171) );
NOR2_X1 U840 ( .A1(n1050), .A2(n1129), .ZN(n1176) );
NAND2_X1 U841 ( .A1(n1177), .A2(n1178), .ZN(n1164) );
OR3_X1 U842 ( .A1(n1179), .A2(n1180), .A3(n1178), .ZN(n1163) );
INV_X1 U843 ( .A(KEYINPUT60), .ZN(n1178) );
INV_X1 U844 ( .A(n1026), .ZN(n1105) );
NAND4_X1 U845 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1026) );
AND4_X1 U846 ( .A1(n1014), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1184) );
NAND3_X1 U847 ( .A1(n1033), .A2(n1050), .A3(n1128), .ZN(n1014) );
NAND2_X1 U848 ( .A1(n1188), .A2(n1189), .ZN(n1183) );
NAND4_X1 U849 ( .A1(n1190), .A2(n1129), .A3(n1191), .A4(n1033), .ZN(n1181) );
NOR2_X1 U850 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U851 ( .A(n1179), .B(KEYINPUT8), .Z(n1190) );
NAND2_X1 U852 ( .A1(KEYINPUT17), .A2(n1194), .ZN(n1155) );
NOR2_X1 U853 ( .A1(n1016), .A2(G952), .ZN(n1109) );
XOR2_X1 U854 ( .A(n1195), .B(n1196), .Z(G48) );
NAND3_X1 U855 ( .A1(n1129), .A2(n1197), .A3(n1198), .ZN(n1196) );
XOR2_X1 U856 ( .A(KEYINPUT49), .B(n1175), .Z(n1197) );
XNOR2_X1 U857 ( .A(G143), .B(n1170), .ZN(G45) );
NAND4_X1 U858 ( .A1(n1199), .A2(n1200), .A3(n1041), .A4(n1201), .ZN(n1170) );
NOR3_X1 U859 ( .A1(n1202), .A2(n1179), .A3(n1193), .ZN(n1201) );
XOR2_X1 U860 ( .A(n1203), .B(n1169), .Z(G42) );
NAND3_X1 U861 ( .A1(n1129), .A2(n1204), .A3(n1205), .ZN(n1169) );
XOR2_X1 U862 ( .A(G137), .B(n1206), .Z(G39) );
NOR2_X1 U863 ( .A1(KEYINPUT20), .A2(n1168), .ZN(n1206) );
NAND3_X1 U864 ( .A1(n1207), .A2(n1064), .A3(n1205), .ZN(n1168) );
XOR2_X1 U865 ( .A(n1208), .B(n1167), .Z(G36) );
NAND2_X1 U866 ( .A1(n1205), .A2(n1188), .ZN(n1167) );
NOR3_X1 U867 ( .A1(n1193), .A2(n1175), .A3(n1035), .ZN(n1205) );
XOR2_X1 U868 ( .A(n1209), .B(n1210), .Z(G33) );
NAND2_X1 U869 ( .A1(n1211), .A2(n1027), .ZN(n1210) );
INV_X1 U870 ( .A(n1035), .ZN(n1027) );
NAND2_X1 U871 ( .A1(n1062), .A2(n1212), .ZN(n1035) );
XOR2_X1 U872 ( .A(n1173), .B(KEYINPUT18), .Z(n1211) );
NAND4_X1 U873 ( .A1(n1129), .A2(n1054), .A3(n1041), .A4(n1200), .ZN(n1173) );
XOR2_X1 U874 ( .A(n1213), .B(n1214), .Z(G30) );
NAND3_X1 U875 ( .A1(n1198), .A2(n1050), .A3(n1215), .ZN(n1214) );
XOR2_X1 U876 ( .A(n1200), .B(KEYINPUT51), .Z(n1215) );
INV_X1 U877 ( .A(n1174), .ZN(n1198) );
NAND3_X1 U878 ( .A1(n1054), .A2(n1059), .A3(n1207), .ZN(n1174) );
INV_X1 U879 ( .A(n1193), .ZN(n1054) );
XNOR2_X1 U880 ( .A(G101), .B(n1020), .ZN(G3) );
NAND3_X1 U881 ( .A1(n1128), .A2(n1041), .A3(n1064), .ZN(n1020) );
XOR2_X1 U882 ( .A(n1177), .B(n1216), .Z(G27) );
NOR2_X1 U883 ( .A1(KEYINPUT54), .A2(n1194), .ZN(n1216) );
AND2_X1 U884 ( .A1(n1180), .A2(n1059), .ZN(n1177) );
NOR4_X1 U885 ( .A1(n1030), .A2(n1029), .A3(n1058), .A4(n1175), .ZN(n1180) );
INV_X1 U886 ( .A(n1200), .ZN(n1175) );
NAND2_X1 U887 ( .A1(n1217), .A2(n1218), .ZN(n1200) );
NAND2_X1 U888 ( .A1(n1219), .A2(n1090), .ZN(n1218) );
INV_X1 U889 ( .A(G900), .ZN(n1090) );
XNOR2_X1 U890 ( .A(G122), .B(n1182), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1220), .A2(n1189), .A3(n1033), .A4(n1199), .ZN(n1182) );
INV_X1 U892 ( .A(n1082), .ZN(n1199) );
NAND2_X1 U893 ( .A1(n1221), .A2(n1222), .ZN(G21) );
OR2_X1 U894 ( .A1(n1187), .A2(G119), .ZN(n1222) );
XOR2_X1 U895 ( .A(n1223), .B(KEYINPUT16), .Z(n1221) );
NAND2_X1 U896 ( .A1(G119), .A2(n1187), .ZN(n1223) );
NAND3_X1 U897 ( .A1(n1189), .A2(n1064), .A3(n1207), .ZN(n1187) );
AND2_X1 U898 ( .A1(n1224), .A2(n1225), .ZN(n1207) );
XNOR2_X1 U899 ( .A(KEYINPUT33), .B(n1072), .ZN(n1225) );
XOR2_X1 U900 ( .A(n1226), .B(KEYINPUT1), .Z(n1224) );
XNOR2_X1 U901 ( .A(G116), .B(n1227), .ZN(G18) );
NAND4_X1 U902 ( .A1(n1188), .A2(n1065), .A3(n1228), .A4(n1229), .ZN(n1227) );
XOR2_X1 U903 ( .A(KEYINPUT55), .B(n1059), .Z(n1228) );
INV_X1 U904 ( .A(n1029), .ZN(n1065) );
AND2_X1 U905 ( .A1(n1050), .A2(n1041), .ZN(n1188) );
NOR2_X1 U906 ( .A1(n1220), .A2(n1082), .ZN(n1050) );
XNOR2_X1 U907 ( .A(G113), .B(n1186), .ZN(G15) );
NAND3_X1 U908 ( .A1(n1129), .A2(n1041), .A3(n1189), .ZN(n1186) );
NOR3_X1 U909 ( .A1(n1179), .A2(n1192), .A3(n1029), .ZN(n1189) );
NAND2_X1 U910 ( .A1(n1230), .A2(n1056), .ZN(n1029) );
NAND2_X1 U911 ( .A1(n1231), .A2(n1232), .ZN(n1041) );
OR2_X1 U912 ( .A1(n1042), .A2(KEYINPUT33), .ZN(n1232) );
INV_X1 U913 ( .A(n1033), .ZN(n1042) );
NOR2_X1 U914 ( .A1(n1072), .A2(n1233), .ZN(n1033) );
NAND3_X1 U915 ( .A1(n1072), .A2(n1226), .A3(KEYINPUT33), .ZN(n1231) );
INV_X1 U916 ( .A(n1030), .ZN(n1129) );
NAND2_X1 U917 ( .A1(n1220), .A2(n1082), .ZN(n1030) );
XNOR2_X1 U918 ( .A(G110), .B(n1185), .ZN(G12) );
NAND3_X1 U919 ( .A1(n1204), .A2(n1128), .A3(n1064), .ZN(n1185) );
INV_X1 U920 ( .A(n1052), .ZN(n1064) );
NAND2_X1 U921 ( .A1(n1082), .A2(n1202), .ZN(n1052) );
INV_X1 U922 ( .A(n1220), .ZN(n1202) );
XOR2_X1 U923 ( .A(n1234), .B(n1235), .Z(n1220) );
NOR2_X1 U924 ( .A1(KEYINPUT31), .A2(n1080), .ZN(n1235) );
NOR2_X1 U925 ( .A1(n1121), .A2(G902), .ZN(n1080) );
XNOR2_X1 U926 ( .A(n1236), .B(n1237), .ZN(n1121) );
XOR2_X1 U927 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U928 ( .A(n1209), .B(n1240), .Z(n1239) );
NAND2_X1 U929 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
NAND2_X1 U930 ( .A1(G104), .A2(n1243), .ZN(n1242) );
NAND2_X1 U931 ( .A1(KEYINPUT46), .A2(n1244), .ZN(n1243) );
NAND2_X1 U932 ( .A1(KEYINPUT26), .A2(n1245), .ZN(n1244) );
INV_X1 U933 ( .A(n1246), .ZN(n1245) );
NAND2_X1 U934 ( .A1(n1246), .A2(n1247), .ZN(n1241) );
NAND2_X1 U935 ( .A1(KEYINPUT26), .A2(n1248), .ZN(n1247) );
NAND2_X1 U936 ( .A1(KEYINPUT46), .A2(n1249), .ZN(n1248) );
NOR2_X1 U937 ( .A1(KEYINPUT45), .A2(n1250), .ZN(n1238) );
XOR2_X1 U938 ( .A(n1203), .B(n1251), .Z(n1250) );
NAND2_X1 U939 ( .A1(KEYINPUT62), .A2(n1194), .ZN(n1251) );
XNOR2_X1 U940 ( .A(n1252), .B(n1253), .ZN(n1236) );
AND2_X1 U941 ( .A1(G214), .A2(n1254), .ZN(n1253) );
XOR2_X1 U942 ( .A(n1081), .B(KEYINPUT40), .Z(n1234) );
INV_X1 U943 ( .A(G475), .ZN(n1081) );
XOR2_X1 U944 ( .A(n1255), .B(G478), .Z(n1082) );
NAND2_X1 U945 ( .A1(n1116), .A2(n1161), .ZN(n1255) );
XNOR2_X1 U946 ( .A(n1256), .B(n1257), .ZN(n1116) );
XOR2_X1 U947 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U948 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U949 ( .A1(KEYINPUT52), .A2(n1262), .ZN(n1261) );
XOR2_X1 U950 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U951 ( .A(G122), .B(KEYINPUT2), .ZN(n1263) );
NAND2_X1 U952 ( .A1(n1265), .A2(G217), .ZN(n1260) );
XOR2_X1 U953 ( .A(n1213), .B(n1266), .Z(n1256) );
XOR2_X1 U954 ( .A(KEYINPUT41), .B(G134), .Z(n1266) );
INV_X1 U955 ( .A(G128), .ZN(n1213) );
NOR3_X1 U956 ( .A1(n1179), .A2(n1192), .A3(n1193), .ZN(n1128) );
NAND2_X1 U957 ( .A1(n1055), .A2(n1056), .ZN(n1193) );
NAND2_X1 U958 ( .A1(G221), .A2(n1267), .ZN(n1056) );
INV_X1 U959 ( .A(n1230), .ZN(n1055) );
XOR2_X1 U960 ( .A(n1268), .B(G469), .Z(n1230) );
NAND2_X1 U961 ( .A1(n1269), .A2(n1161), .ZN(n1268) );
XNOR2_X1 U962 ( .A(n1150), .B(n1270), .ZN(n1269) );
XOR2_X1 U963 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U964 ( .A1(KEYINPUT4), .A2(n1145), .ZN(n1272) );
XNOR2_X1 U965 ( .A(n1273), .B(n1094), .ZN(n1145) );
XOR2_X1 U966 ( .A(n1252), .B(n1274), .Z(n1094) );
XOR2_X1 U967 ( .A(KEYINPUT13), .B(G128), .Z(n1274) );
NAND2_X1 U968 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
XOR2_X1 U970 ( .A(n1279), .B(KEYINPUT0), .Z(n1275) );
OR2_X1 U971 ( .A1(n1278), .A2(n1277), .ZN(n1279) );
XOR2_X1 U972 ( .A(G107), .B(G104), .Z(n1277) );
NAND3_X1 U973 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1271) );
OR2_X1 U974 ( .A1(n1149), .A2(n1144), .ZN(n1282) );
NAND2_X1 U975 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
INV_X1 U976 ( .A(KEYINPUT35), .ZN(n1284) );
NAND2_X1 U977 ( .A1(n1285), .A2(n1149), .ZN(n1283) );
XOR2_X1 U978 ( .A(KEYINPUT61), .B(n1286), .Z(n1285) );
INV_X1 U979 ( .A(n1144), .ZN(n1286) );
NAND2_X1 U980 ( .A1(KEYINPUT35), .A2(n1287), .ZN(n1280) );
NAND2_X1 U981 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
OR2_X1 U982 ( .A1(n1144), .A2(KEYINPUT61), .ZN(n1289) );
NAND3_X1 U983 ( .A1(n1144), .A2(n1149), .A3(KEYINPUT61), .ZN(n1288) );
NAND2_X1 U984 ( .A1(G227), .A2(n1016), .ZN(n1149) );
XOR2_X1 U985 ( .A(G110), .B(G140), .Z(n1144) );
INV_X1 U986 ( .A(n1229), .ZN(n1192) );
NAND2_X1 U987 ( .A1(n1217), .A2(n1290), .ZN(n1229) );
NAND2_X1 U988 ( .A1(n1219), .A2(n1102), .ZN(n1290) );
INV_X1 U989 ( .A(G898), .ZN(n1102) );
NOR3_X1 U990 ( .A1(n1161), .A2(n1043), .A3(n1016), .ZN(n1219) );
NAND3_X1 U991 ( .A1(n1291), .A2(n1016), .A3(G952), .ZN(n1217) );
XOR2_X1 U992 ( .A(KEYINPUT58), .B(n1043), .Z(n1291) );
INV_X1 U993 ( .A(n1031), .ZN(n1043) );
NAND2_X1 U994 ( .A1(G237), .A2(G234), .ZN(n1031) );
INV_X1 U995 ( .A(n1059), .ZN(n1179) );
NOR2_X1 U996 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
INV_X1 U997 ( .A(n1212), .ZN(n1063) );
NAND2_X1 U998 ( .A1(G214), .A2(n1292), .ZN(n1212) );
XNOR2_X1 U999 ( .A(n1293), .B(n1160), .ZN(n1062) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1292), .ZN(n1160) );
NAND2_X1 U1001 ( .A1(n1294), .A2(n1161), .ZN(n1292) );
INV_X1 U1002 ( .A(G237), .ZN(n1294) );
NAND4_X1 U1003 ( .A1(n1295), .A2(n1161), .A3(n1296), .A4(n1297), .ZN(n1293) );
NAND2_X1 U1004 ( .A1(KEYINPUT42), .A2(n1298), .ZN(n1297) );
NAND2_X1 U1005 ( .A1(n1103), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U1006 ( .A(KEYINPUT9), .B(n1300), .ZN(n1299) );
NAND2_X1 U1007 ( .A1(n1301), .A2(n1302), .ZN(n1296) );
INV_X1 U1008 ( .A(KEYINPUT42), .ZN(n1302) );
NAND2_X1 U1009 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
NAND3_X1 U1010 ( .A1(KEYINPUT9), .A2(n1103), .A3(n1300), .ZN(n1304) );
OR2_X1 U1011 ( .A1(n1300), .A2(KEYINPUT9), .ZN(n1303) );
OR2_X1 U1012 ( .A1(n1300), .A2(n1103), .ZN(n1295) );
XOR2_X1 U1013 ( .A(n1305), .B(n1306), .Z(n1103) );
XOR2_X1 U1014 ( .A(n1278), .B(n1307), .Z(n1306) );
XOR2_X1 U1015 ( .A(n1246), .B(n1308), .Z(n1307) );
XOR2_X1 U1016 ( .A(G113), .B(G122), .Z(n1246) );
XOR2_X1 U1017 ( .A(n1139), .B(KEYINPUT63), .Z(n1278) );
XOR2_X1 U1018 ( .A(n1309), .B(n1310), .Z(n1305) );
XOR2_X1 U1019 ( .A(KEYINPUT47), .B(KEYINPUT22), .Z(n1310) );
XOR2_X1 U1020 ( .A(n1249), .B(n1264), .Z(n1309) );
XOR2_X1 U1021 ( .A(G107), .B(G116), .Z(n1264) );
INV_X1 U1022 ( .A(G104), .ZN(n1249) );
XOR2_X1 U1023 ( .A(n1311), .B(n1312), .Z(n1300) );
INV_X1 U1024 ( .A(n1154), .ZN(n1312) );
XOR2_X1 U1025 ( .A(n1313), .B(n1314), .Z(n1311) );
NOR2_X1 U1026 ( .A1(KEYINPUT10), .A2(n1194), .ZN(n1314) );
NAND2_X1 U1027 ( .A1(KEYINPUT19), .A2(n1157), .ZN(n1313) );
NOR2_X1 U1028 ( .A1(n1108), .A2(G953), .ZN(n1157) );
INV_X1 U1029 ( .A(G224), .ZN(n1108) );
INV_X1 U1030 ( .A(n1058), .ZN(n1204) );
NAND2_X1 U1031 ( .A1(n1315), .A2(n1233), .ZN(n1058) );
INV_X1 U1032 ( .A(n1226), .ZN(n1233) );
NAND3_X1 U1033 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1226) );
NAND2_X1 U1034 ( .A1(n1073), .A2(n1319), .ZN(n1318) );
NAND3_X1 U1035 ( .A1(n1320), .A2(n1079), .A3(KEYINPUT59), .ZN(n1317) );
INV_X1 U1036 ( .A(n1073), .ZN(n1079) );
NOR2_X1 U1037 ( .A1(n1113), .A2(G902), .ZN(n1073) );
XNOR2_X1 U1038 ( .A(n1321), .B(n1322), .ZN(n1113) );
XNOR2_X1 U1039 ( .A(n1323), .B(n1093), .ZN(n1322) );
XOR2_X1 U1040 ( .A(n1194), .B(n1203), .Z(n1093) );
INV_X1 U1041 ( .A(G140), .ZN(n1203) );
INV_X1 U1042 ( .A(G125), .ZN(n1194) );
NAND2_X1 U1043 ( .A1(KEYINPUT3), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1044 ( .A(G128), .B(n1308), .Z(n1324) );
XOR2_X1 U1045 ( .A(G110), .B(G119), .Z(n1308) );
XOR2_X1 U1046 ( .A(n1325), .B(G146), .Z(n1321) );
NAND2_X1 U1047 ( .A1(n1326), .A2(KEYINPUT21), .ZN(n1325) );
XOR2_X1 U1048 ( .A(n1327), .B(G137), .Z(n1326) );
NAND2_X1 U1049 ( .A1(n1265), .A2(G221), .ZN(n1327) );
AND2_X1 U1050 ( .A1(G234), .A2(n1016), .ZN(n1265) );
INV_X1 U1051 ( .A(G953), .ZN(n1016) );
INV_X1 U1052 ( .A(n1319), .ZN(n1320) );
NAND2_X1 U1053 ( .A1(KEYINPUT36), .A2(n1074), .ZN(n1319) );
OR2_X1 U1054 ( .A1(n1074), .A2(KEYINPUT59), .ZN(n1316) );
NAND2_X1 U1055 ( .A1(G217), .A2(n1267), .ZN(n1074) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1161), .ZN(n1267) );
XNOR2_X1 U1057 ( .A(n1072), .B(KEYINPUT25), .ZN(n1315) );
XNOR2_X1 U1058 ( .A(n1328), .B(G472), .ZN(n1072) );
NAND2_X1 U1059 ( .A1(n1329), .A2(n1161), .ZN(n1328) );
INV_X1 U1060 ( .A(G902), .ZN(n1161) );
XOR2_X1 U1061 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1062 ( .A(n1137), .B(n1139), .ZN(n1331) );
XOR2_X1 U1063 ( .A(G101), .B(KEYINPUT5), .Z(n1139) );
NAND2_X1 U1064 ( .A1(n1254), .A2(G210), .ZN(n1137) );
NOR2_X1 U1065 ( .A1(G953), .A2(G237), .ZN(n1254) );
XOR2_X1 U1066 ( .A(n1332), .B(KEYINPUT34), .Z(n1330) );
NAND3_X1 U1067 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1332) );
OR2_X1 U1068 ( .A1(n1138), .A2(n1336), .ZN(n1335) );
NAND3_X1 U1069 ( .A1(n1336), .A2(n1138), .A3(KEYINPUT6), .ZN(n1334) );
XOR2_X1 U1070 ( .A(n1150), .B(n1154), .Z(n1138) );
XOR2_X1 U1071 ( .A(n1337), .B(G128), .Z(n1154) );
NAND2_X1 U1072 ( .A1(KEYINPUT11), .A2(n1252), .ZN(n1337) );
XOR2_X1 U1073 ( .A(n1195), .B(n1258), .Z(n1252) );
XNOR2_X1 U1074 ( .A(G143), .B(KEYINPUT29), .ZN(n1258) );
INV_X1 U1075 ( .A(G146), .ZN(n1195) );
XNOR2_X1 U1076 ( .A(n1209), .B(n1338), .ZN(n1150) );
NOR2_X1 U1077 ( .A1(KEYINPUT24), .A2(n1095), .ZN(n1338) );
XOR2_X1 U1078 ( .A(n1208), .B(G137), .Z(n1095) );
INV_X1 U1079 ( .A(G134), .ZN(n1208) );
INV_X1 U1080 ( .A(G131), .ZN(n1209) );
NOR2_X1 U1081 ( .A1(KEYINPUT28), .A2(n1133), .ZN(n1336) );
NAND2_X1 U1082 ( .A1(n1133), .A2(n1339), .ZN(n1333) );
INV_X1 U1083 ( .A(KEYINPUT6), .ZN(n1339) );
XNOR2_X1 U1084 ( .A(n1340), .B(n1341), .ZN(n1133) );
XNOR2_X1 U1085 ( .A(G116), .B(n1342), .ZN(n1341) );
NAND2_X1 U1086 ( .A1(n1343), .A2(KEYINPUT12), .ZN(n1342) );
XNOR2_X1 U1087 ( .A(G113), .B(KEYINPUT22), .ZN(n1343) );
NAND2_X1 U1088 ( .A1(KEYINPUT44), .A2(G119), .ZN(n1340) );
endmodule


