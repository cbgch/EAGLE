//Key = 0100010110011100110101010011111100101010001011110100011000001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
n1401, n1402, n1403;

XNOR2_X1 U763 ( .A(G107), .B(n1061), .ZN(G9) );
NOR2_X1 U764 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR3_X1 U765 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NOR3_X1 U766 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1065) );
NOR2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR3_X1 U768 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NOR2_X1 U769 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U770 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR3_X1 U771 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NOR2_X1 U772 ( .A1(KEYINPUT61), .A2(n1082), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1077) );
NOR2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U775 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U776 ( .A1(n1089), .A2(n1090), .ZN(n1073) );
AND3_X1 U777 ( .A1(KEYINPUT61), .A2(n1083), .A3(n1091), .ZN(n1090) );
INV_X1 U778 ( .A(n1075), .ZN(n1089) );
NOR2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1070) );
INV_X1 U780 ( .A(n1094), .ZN(n1093) );
NOR2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NOR2_X1 U782 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NAND3_X1 U783 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1064) );
NAND3_X1 U784 ( .A1(n1102), .A2(n1103), .A3(n1094), .ZN(n1101) );
NOR3_X1 U785 ( .A1(n1079), .A2(n1086), .A3(n1075), .ZN(n1094) );
NAND2_X1 U786 ( .A1(KEYINPUT54), .A2(n1104), .ZN(n1075) );
INV_X1 U787 ( .A(n1105), .ZN(n1086) );
NOR3_X1 U788 ( .A1(n1106), .A2(G953), .A3(G952), .ZN(n1062) );
INV_X1 U789 ( .A(n1099), .ZN(n1106) );
NAND4_X1 U790 ( .A1(n1088), .A2(n1098), .A3(n1107), .A4(n1108), .ZN(n1099) );
NOR2_X1 U791 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U792 ( .A(G469), .B(n1111), .ZN(n1110) );
XOR2_X1 U793 ( .A(n1112), .B(KEYINPUT35), .Z(n1109) );
NAND4_X1 U794 ( .A1(n1113), .A2(n1105), .A3(n1114), .A4(n1115), .ZN(n1112) );
NAND2_X1 U795 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U796 ( .A(KEYINPUT58), .B(n1118), .ZN(n1116) );
XOR2_X1 U797 ( .A(KEYINPUT45), .B(n1119), .Z(n1114) );
NOR2_X1 U798 ( .A1(n1120), .A2(n1117), .ZN(n1119) );
XNOR2_X1 U799 ( .A(G472), .B(KEYINPUT11), .ZN(n1120) );
XNOR2_X1 U800 ( .A(n1121), .B(n1122), .ZN(n1107) );
NAND2_X1 U801 ( .A1(KEYINPUT30), .A2(n1123), .ZN(n1122) );
XOR2_X1 U802 ( .A(n1124), .B(n1125), .Z(G72) );
XOR2_X1 U803 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U804 ( .A1(n1128), .A2(n1100), .ZN(n1127) );
AND2_X1 U805 ( .A1(G227), .A2(G900), .ZN(n1128) );
NOR2_X1 U806 ( .A1(KEYINPUT50), .A2(n1129), .ZN(n1126) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U808 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND2_X1 U809 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NAND3_X1 U810 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
XOR2_X1 U811 ( .A(KEYINPUT49), .B(n1139), .Z(n1134) );
NOR2_X1 U812 ( .A1(n1140), .A2(n1138), .ZN(n1139) );
AND2_X1 U813 ( .A1(n1137), .A2(n1136), .ZN(n1140) );
XNOR2_X1 U814 ( .A(n1141), .B(KEYINPUT34), .ZN(n1136) );
NAND2_X1 U815 ( .A1(G131), .A2(n1142), .ZN(n1141) );
OR2_X1 U816 ( .A1(n1142), .A2(G131), .ZN(n1137) );
NAND3_X1 U817 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
NAND2_X1 U818 ( .A1(G134), .A2(n1146), .ZN(n1145) );
NAND2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
INV_X1 U820 ( .A(KEYINPUT53), .ZN(n1148) );
NAND2_X1 U821 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
XNOR2_X1 U822 ( .A(KEYINPUT8), .B(G137), .ZN(n1149) );
NAND2_X1 U823 ( .A1(KEYINPUT53), .A2(n1151), .ZN(n1143) );
NAND2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
OR2_X1 U825 ( .A1(G137), .A2(KEYINPUT8), .ZN(n1153) );
NAND3_X1 U826 ( .A1(G137), .A2(n1150), .A3(KEYINPUT8), .ZN(n1152) );
NOR2_X1 U827 ( .A1(n1154), .A2(n1155), .ZN(n1130) );
XOR2_X1 U828 ( .A(KEYINPUT2), .B(G900), .Z(n1155) );
NAND2_X1 U829 ( .A1(n1100), .A2(n1156), .ZN(n1124) );
XOR2_X1 U830 ( .A(n1157), .B(n1158), .Z(G69) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U832 ( .A1(n1161), .A2(n1100), .ZN(n1160) );
NOR2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1159) );
XOR2_X1 U834 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U835 ( .A(n1166), .B(n1167), .ZN(n1165) );
NOR2_X1 U836 ( .A1(G898), .A2(n1154), .ZN(n1162) );
INV_X1 U837 ( .A(n1168), .ZN(n1154) );
NOR2_X1 U838 ( .A1(n1169), .A2(n1100), .ZN(n1157) );
NOR2_X1 U839 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(G66) );
XNOR2_X1 U841 ( .A(n1174), .B(n1175), .ZN(n1173) );
NOR2_X1 U842 ( .A1(n1176), .A2(n1177), .ZN(n1174) );
NOR2_X1 U843 ( .A1(n1172), .A2(n1178), .ZN(G63) );
XOR2_X1 U844 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U845 ( .A1(n1181), .A2(n1177), .ZN(n1179) );
NOR2_X1 U846 ( .A1(n1172), .A2(n1182), .ZN(G60) );
XOR2_X1 U847 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1177), .ZN(n1183) );
XOR2_X1 U849 ( .A(n1186), .B(n1187), .Z(G6) );
XNOR2_X1 U850 ( .A(G104), .B(KEYINPUT41), .ZN(n1187) );
NOR2_X1 U851 ( .A1(n1172), .A2(n1188), .ZN(G57) );
XNOR2_X1 U852 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND2_X1 U853 ( .A1(KEYINPUT16), .A2(n1191), .ZN(n1189) );
XOR2_X1 U854 ( .A(n1192), .B(n1193), .Z(n1191) );
NOR2_X1 U855 ( .A1(KEYINPUT51), .A2(n1194), .ZN(n1193) );
NOR2_X1 U856 ( .A1(n1118), .A2(n1177), .ZN(n1192) );
NOR2_X1 U857 ( .A1(n1172), .A2(n1195), .ZN(G54) );
XOR2_X1 U858 ( .A(n1196), .B(n1197), .Z(n1195) );
NOR2_X1 U859 ( .A1(n1198), .A2(n1177), .ZN(n1197) );
NAND3_X1 U860 ( .A1(n1199), .A2(n1200), .A3(KEYINPUT28), .ZN(n1196) );
NAND2_X1 U861 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND2_X1 U862 ( .A1(KEYINPUT29), .A2(n1203), .ZN(n1202) );
OR2_X1 U863 ( .A1(n1204), .A2(KEYINPUT56), .ZN(n1203) );
NAND2_X1 U864 ( .A1(n1205), .A2(n1204), .ZN(n1199) );
NAND3_X1 U865 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1204) );
NAND2_X1 U866 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
OR3_X1 U867 ( .A1(n1210), .A2(n1209), .A3(n1211), .ZN(n1207) );
NOR2_X1 U868 ( .A1(KEYINPUT24), .A2(n1212), .ZN(n1209) );
NAND2_X1 U869 ( .A1(n1213), .A2(n1211), .ZN(n1206) );
INV_X1 U870 ( .A(KEYINPUT26), .ZN(n1211) );
NAND2_X1 U871 ( .A1(n1214), .A2(n1212), .ZN(n1213) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1216), .ZN(n1205) );
NAND2_X1 U873 ( .A1(n1217), .A2(KEYINPUT29), .ZN(n1216) );
INV_X1 U874 ( .A(n1201), .ZN(n1217) );
XNOR2_X1 U875 ( .A(n1218), .B(n1219), .ZN(n1201) );
NAND2_X1 U876 ( .A1(n1220), .A2(KEYINPUT17), .ZN(n1218) );
XNOR2_X1 U877 ( .A(n1221), .B(n1222), .ZN(n1220) );
INV_X1 U878 ( .A(KEYINPUT56), .ZN(n1215) );
NOR2_X1 U879 ( .A1(n1172), .A2(n1223), .ZN(G51) );
NOR3_X1 U880 ( .A1(n1121), .A2(n1224), .A3(n1225), .ZN(n1223) );
NOR3_X1 U881 ( .A1(n1226), .A2(n1123), .A3(n1177), .ZN(n1225) );
NAND2_X1 U882 ( .A1(G902), .A2(n1066), .ZN(n1177) );
INV_X1 U883 ( .A(n1227), .ZN(n1066) );
NOR2_X1 U884 ( .A1(n1228), .A2(n1229), .ZN(n1224) );
NOR2_X1 U885 ( .A1(n1227), .A2(n1123), .ZN(n1228) );
NOR2_X1 U886 ( .A1(n1161), .A2(n1156), .ZN(n1227) );
NAND4_X1 U887 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1156) );
NOR3_X1 U888 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
INV_X1 U889 ( .A(n1237), .ZN(n1235) );
NAND2_X1 U890 ( .A1(n1091), .A2(n1238), .ZN(n1232) );
NAND2_X1 U891 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NAND2_X1 U892 ( .A1(n1241), .A2(n1103), .ZN(n1240) );
OR2_X1 U893 ( .A1(n1242), .A2(n1243), .ZN(n1103) );
NAND2_X1 U894 ( .A1(n1244), .A2(n1245), .ZN(n1239) );
NAND3_X1 U895 ( .A1(n1244), .A2(n1246), .A3(n1247), .ZN(n1230) );
XNOR2_X1 U896 ( .A(n1243), .B(KEYINPUT47), .ZN(n1247) );
NAND4_X1 U897 ( .A1(n1248), .A2(n1186), .A3(n1249), .A4(n1250), .ZN(n1161) );
AND4_X1 U898 ( .A1(n1061), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1250) );
NAND3_X1 U899 ( .A1(n1113), .A2(n1080), .A3(n1254), .ZN(n1061) );
NAND2_X1 U900 ( .A1(n1255), .A2(n1256), .ZN(n1249) );
NAND2_X1 U901 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U902 ( .A(n1091), .B(KEYINPUT40), .ZN(n1257) );
INV_X1 U903 ( .A(n1259), .ZN(n1255) );
NAND3_X1 U904 ( .A1(n1113), .A2(n1254), .A3(n1091), .ZN(n1186) );
NOR2_X1 U905 ( .A1(n1100), .A2(G952), .ZN(n1172) );
XNOR2_X1 U906 ( .A(G146), .B(n1260), .ZN(G48) );
NAND3_X1 U907 ( .A1(n1091), .A2(n1261), .A3(n1244), .ZN(n1260) );
XOR2_X1 U908 ( .A(KEYINPUT4), .B(n1245), .Z(n1261) );
XNOR2_X1 U909 ( .A(G143), .B(n1262), .ZN(G45) );
NAND3_X1 U910 ( .A1(n1243), .A2(n1246), .A3(n1244), .ZN(n1262) );
XOR2_X1 U911 ( .A(n1263), .B(G140), .Z(G42) );
NAND2_X1 U912 ( .A1(KEYINPUT7), .A2(n1264), .ZN(n1263) );
NAND3_X1 U913 ( .A1(n1241), .A2(n1091), .A3(n1242), .ZN(n1264) );
XNOR2_X1 U914 ( .A(n1146), .B(n1234), .ZN(G39) );
AND3_X1 U915 ( .A1(n1245), .A2(n1105), .A3(n1241), .ZN(n1234) );
XNOR2_X1 U916 ( .A(n1150), .B(n1236), .ZN(G36) );
AND3_X1 U917 ( .A1(n1243), .A2(n1080), .A3(n1241), .ZN(n1236) );
AND2_X1 U918 ( .A1(n1102), .A2(n1265), .ZN(n1241) );
NAND2_X1 U919 ( .A1(n1266), .A2(n1267), .ZN(G33) );
NAND2_X1 U920 ( .A1(G131), .A2(n1268), .ZN(n1267) );
XOR2_X1 U921 ( .A(n1269), .B(KEYINPUT20), .Z(n1266) );
OR2_X1 U922 ( .A1(n1268), .A2(G131), .ZN(n1269) );
NAND4_X1 U923 ( .A1(n1265), .A2(n1091), .A3(n1243), .A4(n1270), .ZN(n1268) );
XNOR2_X1 U924 ( .A(KEYINPUT15), .B(n1072), .ZN(n1270) );
INV_X1 U925 ( .A(n1102), .ZN(n1072) );
NOR2_X1 U926 ( .A1(n1097), .A2(n1271), .ZN(n1102) );
INV_X1 U927 ( .A(n1098), .ZN(n1271) );
XNOR2_X1 U928 ( .A(G128), .B(n1237), .ZN(G30) );
NAND3_X1 U929 ( .A1(n1245), .A2(n1080), .A3(n1244), .ZN(n1237) );
AND2_X1 U930 ( .A1(n1265), .A2(n1096), .ZN(n1244) );
AND3_X1 U931 ( .A1(n1272), .A2(n1088), .A3(n1273), .ZN(n1265) );
NAND2_X1 U932 ( .A1(n1274), .A2(n1275), .ZN(n1272) );
INV_X1 U933 ( .A(n1258), .ZN(n1080) );
XOR2_X1 U934 ( .A(n1253), .B(n1276), .Z(G3) );
XNOR2_X1 U935 ( .A(G101), .B(KEYINPUT22), .ZN(n1276) );
NAND4_X1 U936 ( .A1(n1277), .A2(n1105), .A3(n1273), .A4(n1088), .ZN(n1253) );
INV_X1 U937 ( .A(n1087), .ZN(n1273) );
XNOR2_X1 U938 ( .A(G125), .B(n1231), .ZN(G27) );
NAND4_X1 U939 ( .A1(n1242), .A2(n1091), .A3(n1278), .A4(n1083), .ZN(n1231) );
NOR2_X1 U940 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
AND2_X1 U941 ( .A1(n1275), .A2(n1274), .ZN(n1279) );
NAND4_X1 U942 ( .A1(n1281), .A2(G902), .A3(n1168), .A4(n1104), .ZN(n1274) );
XNOR2_X1 U943 ( .A(G900), .B(KEYINPUT2), .ZN(n1281) );
NOR2_X1 U944 ( .A1(n1069), .A2(n1113), .ZN(n1242) );
XOR2_X1 U945 ( .A(n1282), .B(G122), .Z(G24) );
NAND2_X1 U946 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
OR2_X1 U947 ( .A1(n1248), .A2(KEYINPUT59), .ZN(n1284) );
OR2_X1 U948 ( .A1(n1285), .A2(n1280), .ZN(n1248) );
NAND3_X1 U949 ( .A1(n1096), .A2(n1285), .A3(KEYINPUT59), .ZN(n1283) );
NAND3_X1 U950 ( .A1(n1113), .A2(n1083), .A3(n1286), .ZN(n1285) );
AND3_X1 U951 ( .A1(n1287), .A2(n1288), .A3(n1246), .ZN(n1286) );
NAND2_X1 U952 ( .A1(n1289), .A2(n1290), .ZN(n1246) );
OR2_X1 U953 ( .A1(n1082), .A2(KEYINPUT46), .ZN(n1290) );
NAND3_X1 U954 ( .A1(n1291), .A2(n1292), .A3(KEYINPUT46), .ZN(n1289) );
INV_X1 U955 ( .A(n1280), .ZN(n1096) );
XNOR2_X1 U956 ( .A(G119), .B(n1252), .ZN(G21) );
NAND4_X1 U957 ( .A1(n1083), .A2(n1245), .A3(n1293), .A4(n1105), .ZN(n1252) );
NOR2_X1 U958 ( .A1(n1294), .A2(n1280), .ZN(n1293) );
NOR2_X1 U959 ( .A1(n1113), .A2(n1287), .ZN(n1245) );
INV_X1 U960 ( .A(n1067), .ZN(n1113) );
XOR2_X1 U961 ( .A(n1295), .B(n1296), .Z(G18) );
XNOR2_X1 U962 ( .A(KEYINPUT33), .B(n1297), .ZN(n1296) );
NOR2_X1 U963 ( .A1(n1258), .A2(n1259), .ZN(n1295) );
NAND2_X1 U964 ( .A1(n1298), .A2(n1299), .ZN(n1258) );
XNOR2_X1 U965 ( .A(n1292), .B(KEYINPUT9), .ZN(n1299) );
XNOR2_X1 U966 ( .A(KEYINPUT46), .B(n1291), .ZN(n1298) );
XNOR2_X1 U967 ( .A(n1300), .B(n1301), .ZN(G15) );
NOR2_X1 U968 ( .A1(n1082), .A2(n1259), .ZN(n1301) );
NAND2_X1 U969 ( .A1(n1277), .A2(n1083), .ZN(n1259) );
INV_X1 U970 ( .A(n1079), .ZN(n1083) );
NAND2_X1 U971 ( .A1(n1087), .A2(n1088), .ZN(n1079) );
NOR3_X1 U972 ( .A1(n1280), .A2(n1294), .A3(n1302), .ZN(n1277) );
INV_X1 U973 ( .A(n1243), .ZN(n1302) );
NOR2_X1 U974 ( .A1(n1067), .A2(n1287), .ZN(n1243) );
INV_X1 U975 ( .A(n1288), .ZN(n1294) );
INV_X1 U976 ( .A(n1091), .ZN(n1082) );
NOR2_X1 U977 ( .A1(n1291), .A2(n1303), .ZN(n1091) );
INV_X1 U978 ( .A(n1292), .ZN(n1303) );
NAND2_X1 U979 ( .A1(n1304), .A2(n1305), .ZN(G12) );
NAND2_X1 U980 ( .A1(G110), .A2(n1251), .ZN(n1305) );
XOR2_X1 U981 ( .A(KEYINPUT60), .B(n1306), .Z(n1304) );
NOR2_X1 U982 ( .A1(G110), .A2(n1251), .ZN(n1306) );
NAND3_X1 U983 ( .A1(n1254), .A2(n1067), .A3(n1105), .ZN(n1251) );
NOR2_X1 U984 ( .A1(n1291), .A2(n1292), .ZN(n1105) );
XOR2_X1 U985 ( .A(n1307), .B(n1185), .Z(n1292) );
INV_X1 U986 ( .A(G475), .ZN(n1185) );
OR2_X1 U987 ( .A1(n1184), .A2(G902), .ZN(n1307) );
XNOR2_X1 U988 ( .A(n1308), .B(n1309), .ZN(n1184) );
XOR2_X1 U989 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U990 ( .A(n1300), .B(G104), .ZN(n1311) );
XNOR2_X1 U991 ( .A(n1312), .B(G122), .ZN(n1310) );
XNOR2_X1 U992 ( .A(n1313), .B(n1314), .ZN(n1308) );
XOR2_X1 U993 ( .A(n1315), .B(n1316), .Z(n1313) );
NOR2_X1 U994 ( .A1(G131), .A2(KEYINPUT43), .ZN(n1316) );
NAND2_X1 U995 ( .A1(n1317), .A2(G214), .ZN(n1315) );
XOR2_X1 U996 ( .A(n1318), .B(n1181), .Z(n1291) );
INV_X1 U997 ( .A(G478), .ZN(n1181) );
OR2_X1 U998 ( .A1(n1180), .A2(G902), .ZN(n1318) );
XNOR2_X1 U999 ( .A(n1319), .B(KEYINPUT25), .ZN(n1180) );
XOR2_X1 U1000 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1001 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1002 ( .A(n1324), .B(G122), .ZN(n1323) );
XNOR2_X1 U1003 ( .A(KEYINPUT1), .B(n1150), .ZN(n1322) );
INV_X1 U1004 ( .A(G134), .ZN(n1150) );
XOR2_X1 U1005 ( .A(n1325), .B(n1326), .Z(n1320) );
XOR2_X1 U1006 ( .A(n1327), .B(n1328), .Z(n1326) );
NAND2_X1 U1007 ( .A1(KEYINPUT42), .A2(n1312), .ZN(n1328) );
NAND2_X1 U1008 ( .A1(KEYINPUT38), .A2(n1329), .ZN(n1327) );
XNOR2_X1 U1009 ( .A(n1330), .B(n1297), .ZN(n1325) );
NAND2_X1 U1010 ( .A1(G217), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1011 ( .A(n1332), .B(n1176), .Z(n1067) );
NAND2_X1 U1012 ( .A1(G217), .A2(n1333), .ZN(n1176) );
NAND2_X1 U1013 ( .A1(n1334), .A2(n1175), .ZN(n1332) );
XOR2_X1 U1014 ( .A(n1335), .B(n1336), .Z(n1175) );
XNOR2_X1 U1015 ( .A(G137), .B(n1337), .ZN(n1336) );
NAND2_X1 U1016 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NAND2_X1 U1017 ( .A1(n1340), .A2(n1314), .ZN(n1339) );
XOR2_X1 U1018 ( .A(KEYINPUT44), .B(n1341), .Z(n1338) );
NOR2_X1 U1019 ( .A1(n1340), .A2(n1314), .ZN(n1341) );
XNOR2_X1 U1020 ( .A(G146), .B(n1133), .ZN(n1314) );
XOR2_X1 U1021 ( .A(G125), .B(G140), .Z(n1133) );
AND2_X1 U1022 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1023 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XNOR2_X1 U1024 ( .A(G119), .B(n1346), .ZN(n1344) );
NAND2_X1 U1025 ( .A1(n1347), .A2(n1348), .ZN(n1342) );
XNOR2_X1 U1026 ( .A(n1349), .B(n1346), .ZN(n1348) );
NOR2_X1 U1027 ( .A1(KEYINPUT14), .A2(n1324), .ZN(n1346) );
INV_X1 U1028 ( .A(G128), .ZN(n1324) );
XNOR2_X1 U1029 ( .A(G110), .B(KEYINPUT12), .ZN(n1347) );
NAND2_X1 U1030 ( .A1(n1331), .A2(G221), .ZN(n1335) );
AND2_X1 U1031 ( .A1(G234), .A2(n1100), .ZN(n1331) );
XNOR2_X1 U1032 ( .A(G902), .B(KEYINPUT62), .ZN(n1334) );
AND4_X1 U1033 ( .A1(n1288), .A2(n1088), .A3(n1287), .A4(n1350), .ZN(n1254) );
NOR2_X1 U1034 ( .A1(n1280), .A2(n1087), .ZN(n1350) );
XOR2_X1 U1035 ( .A(n1351), .B(n1198), .Z(n1087) );
INV_X1 U1036 ( .A(G469), .ZN(n1198) );
NAND2_X1 U1037 ( .A1(n1352), .A2(KEYINPUT23), .ZN(n1351) );
XOR2_X1 U1038 ( .A(n1111), .B(KEYINPUT37), .Z(n1352) );
NAND2_X1 U1039 ( .A1(n1353), .A2(n1354), .ZN(n1111) );
XNOR2_X1 U1040 ( .A(n1355), .B(n1356), .ZN(n1353) );
INV_X1 U1041 ( .A(n1221), .ZN(n1356) );
XNOR2_X1 U1042 ( .A(n1357), .B(n1358), .ZN(n1221) );
NAND2_X1 U1043 ( .A1(KEYINPUT36), .A2(n1329), .ZN(n1357) );
INV_X1 U1044 ( .A(G107), .ZN(n1329) );
XNOR2_X1 U1045 ( .A(n1359), .B(n1360), .ZN(n1355) );
NOR2_X1 U1046 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
XOR2_X1 U1047 ( .A(n1363), .B(KEYINPUT63), .Z(n1362) );
NAND2_X1 U1048 ( .A1(n1364), .A2(n1212), .ZN(n1363) );
NOR2_X1 U1049 ( .A1(n1364), .A2(n1212), .ZN(n1361) );
NAND2_X1 U1050 ( .A1(n1365), .A2(n1100), .ZN(n1212) );
XOR2_X1 U1051 ( .A(KEYINPUT39), .B(G227), .Z(n1365) );
XNOR2_X1 U1052 ( .A(KEYINPUT13), .B(n1214), .ZN(n1364) );
INV_X1 U1053 ( .A(n1210), .ZN(n1214) );
XOR2_X1 U1054 ( .A(G140), .B(n1345), .Z(n1210) );
INV_X1 U1055 ( .A(G110), .ZN(n1345) );
NAND2_X1 U1056 ( .A1(n1097), .A2(n1098), .ZN(n1280) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1366), .ZN(n1098) );
NAND2_X1 U1058 ( .A1(n1367), .A2(n1368), .ZN(n1097) );
NAND2_X1 U1059 ( .A1(n1121), .A2(n1123), .ZN(n1368) );
XOR2_X1 U1060 ( .A(n1369), .B(KEYINPUT32), .Z(n1367) );
OR2_X1 U1061 ( .A1(n1123), .A2(n1121), .ZN(n1369) );
NOR2_X1 U1062 ( .A1(n1229), .A2(G902), .ZN(n1121) );
INV_X1 U1063 ( .A(n1226), .ZN(n1229) );
XNOR2_X1 U1064 ( .A(n1370), .B(n1371), .ZN(n1226) );
XOR2_X1 U1065 ( .A(n1167), .B(n1372), .Z(n1371) );
XNOR2_X1 U1066 ( .A(n1373), .B(n1374), .ZN(n1372) );
NOR2_X1 U1067 ( .A1(KEYINPUT57), .A2(n1375), .ZN(n1374) );
XNOR2_X1 U1068 ( .A(KEYINPUT19), .B(n1376), .ZN(n1375) );
INV_X1 U1069 ( .A(n1166), .ZN(n1376) );
XNOR2_X1 U1070 ( .A(n1377), .B(n1358), .ZN(n1166) );
XOR2_X1 U1071 ( .A(G101), .B(G104), .Z(n1358) );
XNOR2_X1 U1072 ( .A(G107), .B(KEYINPUT3), .ZN(n1377) );
INV_X1 U1073 ( .A(G125), .ZN(n1373) );
AND2_X1 U1074 ( .A1(n1378), .A2(n1379), .ZN(n1167) );
NAND2_X1 U1075 ( .A1(n1380), .A2(n1300), .ZN(n1379) );
XOR2_X1 U1076 ( .A(KEYINPUT21), .B(n1381), .Z(n1378) );
NOR2_X1 U1077 ( .A1(n1380), .A2(n1300), .ZN(n1381) );
XNOR2_X1 U1078 ( .A(G116), .B(G119), .ZN(n1380) );
XNOR2_X1 U1079 ( .A(n1382), .B(n1138), .ZN(n1370) );
XOR2_X1 U1080 ( .A(n1383), .B(n1384), .Z(n1382) );
NOR2_X1 U1081 ( .A1(G953), .A2(n1170), .ZN(n1384) );
INV_X1 U1082 ( .A(G224), .ZN(n1170) );
NAND2_X1 U1083 ( .A1(KEYINPUT5), .A2(n1164), .ZN(n1383) );
XNOR2_X1 U1084 ( .A(G122), .B(G110), .ZN(n1164) );
NAND2_X1 U1085 ( .A1(G210), .A2(n1366), .ZN(n1123) );
NAND2_X1 U1086 ( .A1(n1385), .A2(n1354), .ZN(n1366) );
XNOR2_X1 U1087 ( .A(G237), .B(KEYINPUT0), .ZN(n1385) );
INV_X1 U1088 ( .A(n1069), .ZN(n1287) );
XOR2_X1 U1089 ( .A(n1117), .B(n1118), .Z(n1069) );
INV_X1 U1090 ( .A(G472), .ZN(n1118) );
NAND2_X1 U1091 ( .A1(n1386), .A2(n1354), .ZN(n1117) );
XOR2_X1 U1092 ( .A(n1387), .B(n1388), .Z(n1386) );
XNOR2_X1 U1093 ( .A(n1194), .B(n1389), .ZN(n1388) );
INV_X1 U1094 ( .A(n1190), .ZN(n1389) );
XNOR2_X1 U1095 ( .A(n1390), .B(G101), .ZN(n1190) );
NAND2_X1 U1096 ( .A1(n1317), .A2(G210), .ZN(n1390) );
NOR2_X1 U1097 ( .A1(G953), .A2(G237), .ZN(n1317) );
XOR2_X1 U1098 ( .A(n1391), .B(n1359), .Z(n1194) );
XNOR2_X1 U1099 ( .A(n1219), .B(n1138), .ZN(n1359) );
INV_X1 U1100 ( .A(n1222), .ZN(n1138) );
XNOR2_X1 U1101 ( .A(n1392), .B(n1393), .ZN(n1222) );
XNOR2_X1 U1102 ( .A(n1312), .B(G128), .ZN(n1393) );
INV_X1 U1103 ( .A(G143), .ZN(n1312) );
XNOR2_X1 U1104 ( .A(G146), .B(KEYINPUT27), .ZN(n1392) );
XNOR2_X1 U1105 ( .A(n1394), .B(n1395), .ZN(n1219) );
XNOR2_X1 U1106 ( .A(KEYINPUT55), .B(n1146), .ZN(n1395) );
INV_X1 U1107 ( .A(G137), .ZN(n1146) );
XNOR2_X1 U1108 ( .A(G131), .B(G134), .ZN(n1394) );
XNOR2_X1 U1109 ( .A(n1396), .B(n1300), .ZN(n1391) );
INV_X1 U1110 ( .A(G113), .ZN(n1300) );
NAND3_X1 U1111 ( .A1(n1397), .A2(n1398), .A3(n1399), .ZN(n1396) );
NAND2_X1 U1112 ( .A1(KEYINPUT6), .A2(n1400), .ZN(n1399) );
NAND3_X1 U1113 ( .A1(n1401), .A2(n1402), .A3(n1297), .ZN(n1398) );
INV_X1 U1114 ( .A(KEYINPUT6), .ZN(n1402) );
OR2_X1 U1115 ( .A1(n1297), .A2(n1401), .ZN(n1397) );
NOR2_X1 U1116 ( .A1(KEYINPUT48), .A2(n1400), .ZN(n1401) );
XNOR2_X1 U1117 ( .A(n1349), .B(KEYINPUT10), .ZN(n1400) );
INV_X1 U1118 ( .A(G119), .ZN(n1349) );
INV_X1 U1119 ( .A(G116), .ZN(n1297) );
XNOR2_X1 U1120 ( .A(KEYINPUT52), .B(KEYINPUT31), .ZN(n1387) );
NAND2_X1 U1121 ( .A1(G221), .A2(n1333), .ZN(n1088) );
NAND2_X1 U1122 ( .A1(G234), .A2(n1354), .ZN(n1333) );
INV_X1 U1123 ( .A(G902), .ZN(n1354) );
NAND2_X1 U1124 ( .A1(n1275), .A2(n1403), .ZN(n1288) );
NAND4_X1 U1125 ( .A1(G902), .A2(n1168), .A3(n1104), .A4(n1171), .ZN(n1403) );
INV_X1 U1126 ( .A(G898), .ZN(n1171) );
XOR2_X1 U1127 ( .A(G953), .B(KEYINPUT18), .Z(n1168) );
NAND3_X1 U1128 ( .A1(n1104), .A2(n1100), .A3(G952), .ZN(n1275) );
INV_X1 U1129 ( .A(G953), .ZN(n1100) );
NAND2_X1 U1130 ( .A1(G237), .A2(G234), .ZN(n1104) );
endmodule


