//Key = 0011001110100101001001011011011101011011010000011001100110011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389;

XNOR2_X1 U767 ( .A(G107), .B(n1073), .ZN(G9) );
NOR2_X1 U768 ( .A1(n1074), .A2(n1075), .ZN(G75) );
NOR3_X1 U769 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1075) );
NAND3_X1 U770 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1076) );
NAND2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND4_X1 U773 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1085) );
NAND2_X1 U774 ( .A1(n1090), .A2(n1091), .ZN(n1084) );
NAND2_X1 U775 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND3_X1 U776 ( .A1(n1088), .A2(n1094), .A3(n1086), .ZN(n1093) );
NAND2_X1 U777 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U778 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
INV_X1 U779 ( .A(n1099), .ZN(n1095) );
NAND2_X1 U780 ( .A1(n1087), .A2(n1100), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NAND2_X1 U782 ( .A1(n1086), .A2(n1103), .ZN(n1102) );
NAND2_X1 U783 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U784 ( .A1(n1088), .A2(n1106), .ZN(n1101) );
NAND2_X1 U785 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U786 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U787 ( .A(n1111), .ZN(n1082) );
NOR3_X1 U788 ( .A1(n1112), .A2(G953), .A3(G952), .ZN(n1074) );
INV_X1 U789 ( .A(n1079), .ZN(n1112) );
NAND4_X1 U790 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1079) );
NOR4_X1 U791 ( .A1(n1109), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1116) );
XOR2_X1 U792 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U793 ( .A(KEYINPUT23), .B(n1122), .ZN(n1121) );
NOR2_X1 U794 ( .A1(n1123), .A2(KEYINPUT12), .ZN(n1120) );
XNOR2_X1 U795 ( .A(n1124), .B(KEYINPUT38), .ZN(n1117) );
INV_X1 U796 ( .A(n1125), .ZN(n1109) );
XOR2_X1 U797 ( .A(n1126), .B(n1127), .Z(n1115) );
XOR2_X1 U798 ( .A(KEYINPUT18), .B(G475), .Z(n1127) );
NAND2_X1 U799 ( .A1(KEYINPUT8), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U800 ( .A(n1129), .B(KEYINPUT1), .ZN(n1114) );
XOR2_X1 U801 ( .A(n1130), .B(n1131), .Z(n1113) );
XOR2_X1 U802 ( .A(KEYINPUT17), .B(G472), .Z(n1131) );
XOR2_X1 U803 ( .A(n1132), .B(n1133), .Z(G72) );
XOR2_X1 U804 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U805 ( .A1(n1136), .A2(n1080), .ZN(n1135) );
AND2_X1 U806 ( .A1(G227), .A2(G900), .ZN(n1136) );
NAND2_X1 U807 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
XOR2_X1 U808 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U809 ( .A(n1141), .B(n1142), .ZN(n1140) );
NAND2_X1 U810 ( .A1(KEYINPUT26), .A2(n1143), .ZN(n1141) );
XOR2_X1 U811 ( .A(KEYINPUT32), .B(n1144), .Z(n1139) );
NOR2_X1 U812 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U813 ( .A(n1147), .B(KEYINPUT29), .Z(n1146) );
NAND2_X1 U814 ( .A1(n1148), .A2(G131), .ZN(n1147) );
XOR2_X1 U815 ( .A(n1149), .B(KEYINPUT22), .Z(n1148) );
NOR2_X1 U816 ( .A1(G131), .A2(n1149), .ZN(n1145) );
XOR2_X1 U817 ( .A(n1150), .B(G134), .Z(n1149) );
NAND2_X1 U818 ( .A1(KEYINPUT47), .A2(n1151), .ZN(n1150) );
XOR2_X1 U819 ( .A(KEYINPUT52), .B(n1152), .Z(n1137) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1080), .ZN(n1152) );
XNOR2_X1 U821 ( .A(G900), .B(KEYINPUT15), .ZN(n1153) );
NAND2_X1 U822 ( .A1(n1080), .A2(n1077), .ZN(n1132) );
NAND3_X1 U823 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(G69) );
XOR2_X1 U824 ( .A(n1157), .B(KEYINPUT14), .Z(n1156) );
NAND2_X1 U825 ( .A1(G953), .A2(n1158), .ZN(n1157) );
NAND2_X1 U826 ( .A1(G898), .A2(n1159), .ZN(n1158) );
OR2_X1 U827 ( .A1(n1160), .A2(G224), .ZN(n1159) );
NAND2_X1 U828 ( .A1(n1161), .A2(n1080), .ZN(n1155) );
XNOR2_X1 U829 ( .A(n1078), .B(n1162), .ZN(n1161) );
NAND4_X1 U830 ( .A1(n1160), .A2(G224), .A3(G898), .A4(G953), .ZN(n1154) );
NOR2_X1 U831 ( .A1(n1163), .A2(n1164), .ZN(G66) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1165) );
NOR2_X1 U834 ( .A1(n1163), .A2(n1169), .ZN(G63) );
NOR2_X1 U835 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U836 ( .A(n1172), .B(n1173), .Z(n1171) );
NAND2_X1 U837 ( .A1(n1167), .A2(G478), .ZN(n1173) );
NAND2_X1 U838 ( .A1(KEYINPUT63), .A2(n1174), .ZN(n1172) );
NOR2_X1 U839 ( .A1(KEYINPUT63), .A2(n1174), .ZN(n1170) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1175), .ZN(G60) );
XOR2_X1 U841 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U842 ( .A1(KEYINPUT50), .A2(n1178), .ZN(n1177) );
XOR2_X1 U843 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U844 ( .A1(n1167), .A2(G475), .ZN(n1176) );
XNOR2_X1 U845 ( .A(G104), .B(n1181), .ZN(G6) );
NOR2_X1 U846 ( .A1(n1163), .A2(n1182), .ZN(G57) );
XOR2_X1 U847 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U848 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U849 ( .A(n1187), .B(KEYINPUT53), .Z(n1186) );
NAND3_X1 U850 ( .A1(G472), .A2(n1188), .A3(n1189), .ZN(n1187) );
XNOR2_X1 U851 ( .A(G902), .B(KEYINPUT2), .ZN(n1189) );
NAND2_X1 U852 ( .A1(KEYINPUT13), .A2(n1190), .ZN(n1185) );
XOR2_X1 U853 ( .A(n1191), .B(n1192), .Z(n1183) );
NOR2_X1 U854 ( .A1(n1163), .A2(n1193), .ZN(G54) );
NOR2_X1 U855 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U856 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U857 ( .A(KEYINPUT43), .B(n1198), .Z(n1197) );
XOR2_X1 U858 ( .A(KEYINPUT40), .B(n1199), .Z(n1196) );
AND2_X1 U859 ( .A1(G469), .A2(n1167), .ZN(n1199) );
AND3_X1 U860 ( .A1(n1167), .A2(n1198), .A3(G469), .ZN(n1194) );
XNOR2_X1 U861 ( .A(n1200), .B(n1201), .ZN(n1198) );
XOR2_X1 U862 ( .A(n1202), .B(n1203), .Z(n1200) );
NOR2_X1 U863 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
XOR2_X1 U864 ( .A(KEYINPUT28), .B(n1206), .Z(n1205) );
NOR3_X1 U865 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1206) );
NOR2_X1 U866 ( .A1(n1210), .A2(n1211), .ZN(n1204) );
INV_X1 U867 ( .A(n1209), .ZN(n1211) );
NOR2_X1 U868 ( .A1(n1208), .A2(n1207), .ZN(n1210) );
NAND2_X1 U869 ( .A1(n1212), .A2(n1213), .ZN(n1207) );
NAND2_X1 U870 ( .A1(KEYINPUT45), .A2(n1143), .ZN(n1213) );
NAND2_X1 U871 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
INV_X1 U872 ( .A(KEYINPUT45), .ZN(n1215) );
NAND2_X1 U873 ( .A1(n1216), .A2(n1217), .ZN(n1202) );
NAND2_X1 U874 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U875 ( .A(n1220), .B(KEYINPUT0), .Z(n1216) );
OR2_X1 U876 ( .A1(n1219), .A2(n1218), .ZN(n1220) );
XNOR2_X1 U877 ( .A(n1221), .B(KEYINPUT30), .ZN(n1219) );
INV_X1 U878 ( .A(n1222), .ZN(n1167) );
NOR3_X1 U879 ( .A1(n1163), .A2(n1223), .A3(n1224), .ZN(G51) );
NOR2_X1 U880 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U881 ( .A(n1227), .B(n1228), .Z(n1226) );
NOR2_X1 U882 ( .A1(KEYINPUT19), .A2(n1229), .ZN(n1228) );
INV_X1 U883 ( .A(n1230), .ZN(n1229) );
NOR2_X1 U884 ( .A1(n1231), .A2(n1232), .ZN(n1223) );
XOR2_X1 U885 ( .A(n1227), .B(n1233), .Z(n1232) );
NOR2_X1 U886 ( .A1(KEYINPUT19), .A2(n1230), .ZN(n1233) );
XNOR2_X1 U887 ( .A(n1234), .B(n1235), .ZN(n1230) );
XNOR2_X1 U888 ( .A(KEYINPUT27), .B(n1236), .ZN(n1235) );
NAND2_X1 U889 ( .A1(KEYINPUT51), .A2(n1221), .ZN(n1234) );
XNOR2_X1 U890 ( .A(n1237), .B(n1160), .ZN(n1227) );
OR2_X1 U891 ( .A1(n1222), .A2(n1122), .ZN(n1237) );
NAND2_X1 U892 ( .A1(G902), .A2(n1188), .ZN(n1222) );
NAND2_X1 U893 ( .A1(n1238), .A2(n1239), .ZN(n1188) );
INV_X1 U894 ( .A(n1077), .ZN(n1239) );
NAND4_X1 U895 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1077) );
NOR3_X1 U896 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
INV_X1 U897 ( .A(n1247), .ZN(n1244) );
NAND2_X1 U898 ( .A1(n1248), .A2(n1249), .ZN(n1242) );
INV_X1 U899 ( .A(KEYINPUT11), .ZN(n1249) );
NAND3_X1 U900 ( .A1(n1086), .A2(n1089), .A3(n1250), .ZN(n1241) );
OR2_X1 U901 ( .A1(n1251), .A2(n1252), .ZN(n1089) );
NAND2_X1 U902 ( .A1(n1253), .A2(n1254), .ZN(n1240) );
NAND2_X1 U903 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
NAND3_X1 U904 ( .A1(n1129), .A2(n1257), .A3(n1250), .ZN(n1256) );
NAND2_X1 U905 ( .A1(n1251), .A2(n1258), .ZN(n1255) );
NAND2_X1 U906 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NAND4_X1 U907 ( .A1(KEYINPUT11), .A2(n1087), .A3(n1261), .A4(n1104), .ZN(n1260) );
INV_X1 U908 ( .A(n1262), .ZN(n1104) );
INV_X1 U909 ( .A(n1078), .ZN(n1238) );
NAND4_X1 U910 ( .A1(n1263), .A2(n1181), .A3(n1264), .A4(n1265), .ZN(n1078) );
AND4_X1 U911 ( .A1(n1073), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1265) );
NAND3_X1 U912 ( .A1(n1252), .A2(n1088), .A3(n1269), .ZN(n1073) );
NOR2_X1 U913 ( .A1(n1270), .A2(n1271), .ZN(n1264) );
NOR2_X1 U914 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XNOR2_X1 U915 ( .A(KEYINPUT7), .B(n1274), .ZN(n1273) );
NAND3_X1 U916 ( .A1(n1269), .A2(n1088), .A3(n1251), .ZN(n1181) );
NAND2_X1 U917 ( .A1(n1253), .A2(n1275), .ZN(n1263) );
XNOR2_X1 U918 ( .A(KEYINPUT4), .B(n1276), .ZN(n1275) );
INV_X1 U919 ( .A(n1225), .ZN(n1231) );
NOR2_X1 U920 ( .A1(n1080), .A2(G952), .ZN(n1163) );
NAND2_X1 U921 ( .A1(n1277), .A2(n1278), .ZN(G48) );
NAND2_X1 U922 ( .A1(G146), .A2(n1279), .ZN(n1278) );
XOR2_X1 U923 ( .A(KEYINPUT59), .B(n1280), .Z(n1277) );
NOR2_X1 U924 ( .A1(G146), .A2(n1279), .ZN(n1280) );
NAND3_X1 U925 ( .A1(n1251), .A2(n1253), .A3(n1281), .ZN(n1279) );
XNOR2_X1 U926 ( .A(G143), .B(n1282), .ZN(G45) );
NAND3_X1 U927 ( .A1(KEYINPUT3), .A2(n1250), .A3(n1283), .ZN(n1282) );
NOR3_X1 U928 ( .A1(n1107), .A2(n1284), .A3(n1285), .ZN(n1283) );
XNOR2_X1 U929 ( .A(n1143), .B(n1286), .ZN(G42) );
NOR2_X1 U930 ( .A1(KEYINPUT9), .A2(n1247), .ZN(n1286) );
NAND3_X1 U931 ( .A1(n1086), .A2(n1099), .A3(n1287), .ZN(n1247) );
XNOR2_X1 U932 ( .A(n1151), .B(n1246), .ZN(G39) );
AND3_X1 U933 ( .A1(n1281), .A2(n1090), .A3(n1086), .ZN(n1246) );
XNOR2_X1 U934 ( .A(G134), .B(n1288), .ZN(G36) );
NAND3_X1 U935 ( .A1(n1250), .A2(n1252), .A3(n1289), .ZN(n1288) );
XNOR2_X1 U936 ( .A(n1086), .B(KEYINPUT21), .ZN(n1289) );
XNOR2_X1 U937 ( .A(G131), .B(n1290), .ZN(G33) );
NAND3_X1 U938 ( .A1(n1250), .A2(n1086), .A3(n1291), .ZN(n1290) );
XNOR2_X1 U939 ( .A(n1251), .B(KEYINPUT41), .ZN(n1291) );
AND2_X1 U940 ( .A1(n1110), .A2(n1125), .ZN(n1086) );
AND3_X1 U941 ( .A1(n1099), .A2(n1261), .A3(n1292), .ZN(n1250) );
XOR2_X1 U942 ( .A(n1293), .B(n1245), .Z(G30) );
AND3_X1 U943 ( .A1(n1252), .A2(n1253), .A3(n1281), .ZN(n1245) );
INV_X1 U944 ( .A(n1259), .ZN(n1281) );
NAND4_X1 U945 ( .A1(n1099), .A2(n1124), .A3(n1261), .A4(n1294), .ZN(n1259) );
NAND2_X1 U946 ( .A1(KEYINPUT55), .A2(n1295), .ZN(n1293) );
XOR2_X1 U947 ( .A(G101), .B(n1270), .Z(G3) );
AND3_X1 U948 ( .A1(n1090), .A2(n1269), .A3(n1292), .ZN(n1270) );
XNOR2_X1 U949 ( .A(n1236), .B(n1248), .ZN(G27) );
AND3_X1 U950 ( .A1(n1087), .A2(n1253), .A3(n1287), .ZN(n1248) );
AND3_X1 U951 ( .A1(n1262), .A2(n1261), .A3(n1251), .ZN(n1287) );
NAND2_X1 U952 ( .A1(n1111), .A2(n1296), .ZN(n1261) );
NAND4_X1 U953 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1298), .ZN(n1296) );
INV_X1 U954 ( .A(G900), .ZN(n1298) );
XNOR2_X1 U955 ( .A(G122), .B(n1299), .ZN(G24) );
NAND2_X1 U956 ( .A1(KEYINPUT39), .A2(n1300), .ZN(n1299) );
INV_X1 U957 ( .A(n1268), .ZN(n1300) );
NAND4_X1 U958 ( .A1(n1301), .A2(n1088), .A3(n1129), .A4(n1257), .ZN(n1268) );
NOR2_X1 U959 ( .A1(n1294), .A2(n1124), .ZN(n1088) );
XNOR2_X1 U960 ( .A(G119), .B(n1267), .ZN(G21) );
NAND4_X1 U961 ( .A1(n1301), .A2(n1090), .A3(n1124), .A4(n1294), .ZN(n1267) );
XOR2_X1 U962 ( .A(G116), .B(n1302), .Z(G18) );
NOR2_X1 U963 ( .A1(n1107), .A2(n1276), .ZN(n1302) );
NAND4_X1 U964 ( .A1(n1292), .A2(n1087), .A3(n1252), .A4(n1303), .ZN(n1276) );
NOR2_X1 U965 ( .A1(n1257), .A2(n1285), .ZN(n1252) );
INV_X1 U966 ( .A(n1129), .ZN(n1285) );
INV_X1 U967 ( .A(n1253), .ZN(n1107) );
XNOR2_X1 U968 ( .A(n1304), .B(n1305), .ZN(G15) );
NOR2_X1 U969 ( .A1(n1274), .A2(n1272), .ZN(n1305) );
NAND2_X1 U970 ( .A1(n1292), .A2(n1301), .ZN(n1272) );
AND3_X1 U971 ( .A1(n1253), .A2(n1303), .A3(n1087), .ZN(n1301) );
INV_X1 U972 ( .A(n1118), .ZN(n1087) );
NAND2_X1 U973 ( .A1(n1098), .A2(n1306), .ZN(n1118) );
INV_X1 U974 ( .A(n1105), .ZN(n1292) );
NAND2_X1 U975 ( .A1(n1307), .A2(n1294), .ZN(n1105) );
INV_X1 U976 ( .A(n1251), .ZN(n1274) );
NOR2_X1 U977 ( .A1(n1129), .A2(n1284), .ZN(n1251) );
INV_X1 U978 ( .A(n1257), .ZN(n1284) );
XNOR2_X1 U979 ( .A(G110), .B(n1266), .ZN(G12) );
NAND3_X1 U980 ( .A1(n1262), .A2(n1269), .A3(n1090), .ZN(n1266) );
NOR2_X1 U981 ( .A1(n1129), .A2(n1257), .ZN(n1090) );
XNOR2_X1 U982 ( .A(n1128), .B(G475), .ZN(n1257) );
NAND2_X1 U983 ( .A1(n1308), .A2(n1309), .ZN(n1128) );
XNOR2_X1 U984 ( .A(n1180), .B(n1179), .ZN(n1308) );
NOR2_X1 U985 ( .A1(KEYINPUT61), .A2(n1310), .ZN(n1179) );
XOR2_X1 U986 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U987 ( .A(G143), .B(G131), .Z(n1312) );
XOR2_X1 U988 ( .A(n1313), .B(n1314), .Z(n1311) );
NOR2_X1 U989 ( .A1(KEYINPUT34), .A2(n1315), .ZN(n1314) );
XOR2_X1 U990 ( .A(n1316), .B(n1317), .Z(n1315) );
NOR2_X1 U991 ( .A1(G140), .A2(KEYINPUT5), .ZN(n1317) );
XNOR2_X1 U992 ( .A(G125), .B(G146), .ZN(n1316) );
NAND2_X1 U993 ( .A1(n1318), .A2(G214), .ZN(n1313) );
XOR2_X1 U994 ( .A(G104), .B(n1319), .Z(n1180) );
XNOR2_X1 U995 ( .A(G122), .B(n1304), .ZN(n1319) );
XNOR2_X1 U996 ( .A(n1320), .B(G478), .ZN(n1129) );
NAND2_X1 U997 ( .A1(n1174), .A2(n1309), .ZN(n1320) );
XNOR2_X1 U998 ( .A(n1321), .B(n1322), .ZN(n1174) );
XOR2_X1 U999 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1000 ( .A(G122), .B(G116), .Z(n1324) );
XOR2_X1 U1001 ( .A(KEYINPUT42), .B(G134), .Z(n1323) );
XOR2_X1 U1002 ( .A(n1325), .B(n1326), .Z(n1321) );
XOR2_X1 U1003 ( .A(n1327), .B(n1328), .Z(n1325) );
AND2_X1 U1004 ( .A1(n1329), .A2(G217), .ZN(n1328) );
NAND2_X1 U1005 ( .A1(n1330), .A2(KEYINPUT24), .ZN(n1327) );
XNOR2_X1 U1006 ( .A(G107), .B(KEYINPUT48), .ZN(n1330) );
AND3_X1 U1007 ( .A1(n1253), .A2(n1303), .A3(n1099), .ZN(n1269) );
NOR2_X1 U1008 ( .A1(n1098), .A2(n1097), .ZN(n1099) );
INV_X1 U1009 ( .A(n1306), .ZN(n1097) );
NAND2_X1 U1010 ( .A1(G221), .A2(n1331), .ZN(n1306) );
XOR2_X1 U1011 ( .A(n1332), .B(G469), .Z(n1098) );
NAND2_X1 U1012 ( .A1(n1333), .A2(n1309), .ZN(n1332) );
XOR2_X1 U1013 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1014 ( .A(n1336), .B(n1201), .Z(n1335) );
NOR2_X1 U1015 ( .A1(n1214), .A2(n1208), .ZN(n1336) );
AND2_X1 U1016 ( .A1(G110), .A2(n1143), .ZN(n1208) );
NOR2_X1 U1017 ( .A1(n1143), .A2(G110), .ZN(n1214) );
INV_X1 U1018 ( .A(G140), .ZN(n1143) );
XNOR2_X1 U1019 ( .A(n1337), .B(n1209), .ZN(n1334) );
NAND2_X1 U1020 ( .A1(G227), .A2(n1080), .ZN(n1209) );
NAND2_X1 U1021 ( .A1(KEYINPUT33), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1022 ( .A(n1221), .B(n1218), .Z(n1338) );
XOR2_X1 U1023 ( .A(n1339), .B(n1340), .Z(n1218) );
XNOR2_X1 U1024 ( .A(KEYINPUT54), .B(n1341), .ZN(n1340) );
INV_X1 U1025 ( .A(G107), .ZN(n1341) );
XNOR2_X1 U1026 ( .A(G104), .B(n1342), .ZN(n1339) );
NOR2_X1 U1027 ( .A1(KEYINPUT37), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1028 ( .A1(n1111), .A2(n1344), .ZN(n1303) );
NAND4_X1 U1029 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1345), .ZN(n1344) );
INV_X1 U1030 ( .A(G898), .ZN(n1345) );
NAND3_X1 U1031 ( .A1(n1297), .A2(n1080), .A3(G952), .ZN(n1111) );
NAND2_X1 U1032 ( .A1(G237), .A2(G234), .ZN(n1297) );
NOR2_X1 U1033 ( .A1(n1346), .A2(n1110), .ZN(n1253) );
XNOR2_X1 U1034 ( .A(n1347), .B(n1123), .ZN(n1110) );
AND2_X1 U1035 ( .A1(n1348), .A2(n1309), .ZN(n1123) );
XNOR2_X1 U1036 ( .A(n1160), .B(n1349), .ZN(n1348) );
XNOR2_X1 U1037 ( .A(n1225), .B(n1142), .ZN(n1349) );
XNOR2_X1 U1038 ( .A(G125), .B(n1221), .ZN(n1142) );
NAND2_X1 U1039 ( .A1(G224), .A2(n1080), .ZN(n1225) );
INV_X1 U1040 ( .A(n1162), .ZN(n1160) );
XNOR2_X1 U1041 ( .A(n1350), .B(n1351), .ZN(n1162) );
XOR2_X1 U1042 ( .A(n1343), .B(n1352), .Z(n1351) );
XOR2_X1 U1043 ( .A(n1353), .B(n1354), .Z(n1352) );
NAND3_X1 U1044 ( .A1(n1355), .A2(n1356), .A3(n1357), .ZN(n1353) );
NAND2_X1 U1045 ( .A1(G104), .A2(n1358), .ZN(n1357) );
OR3_X1 U1046 ( .A1(n1358), .A2(n1359), .A3(G107), .ZN(n1356) );
INV_X1 U1047 ( .A(KEYINPUT36), .ZN(n1358) );
NAND2_X1 U1048 ( .A1(G107), .A2(n1359), .ZN(n1355) );
NAND2_X1 U1049 ( .A1(KEYINPUT35), .A2(n1360), .ZN(n1359) );
INV_X1 U1050 ( .A(G104), .ZN(n1360) );
XNOR2_X1 U1051 ( .A(G101), .B(KEYINPUT58), .ZN(n1343) );
XOR2_X1 U1052 ( .A(n1361), .B(n1362), .Z(n1350) );
XNOR2_X1 U1053 ( .A(KEYINPUT44), .B(n1304), .ZN(n1362) );
XOR2_X1 U1054 ( .A(n1363), .B(G110), .Z(n1361) );
NAND2_X1 U1055 ( .A1(KEYINPUT60), .A2(G122), .ZN(n1363) );
NAND2_X1 U1056 ( .A1(KEYINPUT6), .A2(n1122), .ZN(n1347) );
NAND2_X1 U1057 ( .A1(G210), .A2(n1364), .ZN(n1122) );
XNOR2_X1 U1058 ( .A(n1125), .B(KEYINPUT25), .ZN(n1346) );
NAND2_X1 U1059 ( .A1(G214), .A2(n1364), .ZN(n1125) );
NAND2_X1 U1060 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
INV_X1 U1061 ( .A(G237), .ZN(n1366) );
NOR2_X1 U1062 ( .A1(n1294), .A2(n1307), .ZN(n1262) );
INV_X1 U1063 ( .A(n1124), .ZN(n1307) );
XNOR2_X1 U1064 ( .A(n1367), .B(n1168), .ZN(n1124) );
AND2_X1 U1065 ( .A1(G217), .A2(n1331), .ZN(n1168) );
NAND2_X1 U1066 ( .A1(G234), .A2(n1365), .ZN(n1331) );
XNOR2_X1 U1067 ( .A(G902), .B(KEYINPUT49), .ZN(n1365) );
NAND2_X1 U1068 ( .A1(n1166), .A2(n1309), .ZN(n1367) );
XOR2_X1 U1069 ( .A(n1368), .B(n1369), .Z(n1166) );
XOR2_X1 U1070 ( .A(n1370), .B(n1371), .Z(n1369) );
XNOR2_X1 U1071 ( .A(n1236), .B(G119), .ZN(n1371) );
INV_X1 U1072 ( .A(G125), .ZN(n1236) );
XNOR2_X1 U1073 ( .A(G146), .B(n1295), .ZN(n1370) );
XOR2_X1 U1074 ( .A(n1372), .B(n1373), .Z(n1368) );
XNOR2_X1 U1075 ( .A(n1374), .B(n1375), .ZN(n1373) );
NOR2_X1 U1076 ( .A1(G140), .A2(KEYINPUT57), .ZN(n1375) );
NAND2_X1 U1077 ( .A1(KEYINPUT31), .A2(G137), .ZN(n1374) );
XOR2_X1 U1078 ( .A(n1376), .B(G110), .Z(n1372) );
NAND2_X1 U1079 ( .A1(n1329), .A2(G221), .ZN(n1376) );
AND2_X1 U1080 ( .A1(G234), .A2(n1080), .ZN(n1329) );
INV_X1 U1081 ( .A(G953), .ZN(n1080) );
NAND2_X1 U1082 ( .A1(n1377), .A2(n1378), .ZN(n1294) );
OR2_X1 U1083 ( .A1(n1130), .A2(G472), .ZN(n1378) );
XOR2_X1 U1084 ( .A(n1379), .B(KEYINPUT62), .Z(n1377) );
NAND2_X1 U1085 ( .A1(G472), .A2(n1130), .ZN(n1379) );
NAND2_X1 U1086 ( .A1(n1380), .A2(n1309), .ZN(n1130) );
INV_X1 U1087 ( .A(G902), .ZN(n1309) );
XOR2_X1 U1088 ( .A(n1381), .B(n1192), .Z(n1380) );
XNOR2_X1 U1089 ( .A(n1382), .B(G101), .ZN(n1192) );
NAND2_X1 U1090 ( .A1(n1318), .A2(G210), .ZN(n1382) );
NOR2_X1 U1091 ( .A1(G953), .A2(G237), .ZN(n1318) );
XNOR2_X1 U1092 ( .A(KEYINPUT56), .B(n1383), .ZN(n1381) );
NOR2_X1 U1093 ( .A1(KEYINPUT20), .A2(n1384), .ZN(n1383) );
XOR2_X1 U1094 ( .A(n1190), .B(n1385), .Z(n1384) );
NOR2_X1 U1095 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
AND2_X1 U1096 ( .A1(KEYINPUT16), .A2(n1191), .ZN(n1387) );
NOR2_X1 U1097 ( .A1(KEYINPUT46), .A2(n1191), .ZN(n1386) );
XOR2_X1 U1098 ( .A(n1388), .B(n1354), .Z(n1191) );
XOR2_X1 U1099 ( .A(G116), .B(G119), .Z(n1354) );
NAND2_X1 U1100 ( .A1(KEYINPUT10), .A2(n1304), .ZN(n1388) );
INV_X1 U1101 ( .A(G113), .ZN(n1304) );
XOR2_X1 U1102 ( .A(n1201), .B(n1221), .Z(n1190) );
XNOR2_X1 U1103 ( .A(G146), .B(n1326), .ZN(n1221) );
XNOR2_X1 U1104 ( .A(n1295), .B(G143), .ZN(n1326) );
INV_X1 U1105 ( .A(G128), .ZN(n1295) );
XOR2_X1 U1106 ( .A(G131), .B(n1389), .Z(n1201) );
XNOR2_X1 U1107 ( .A(n1151), .B(G134), .ZN(n1389) );
INV_X1 U1108 ( .A(G137), .ZN(n1151) );
endmodule


