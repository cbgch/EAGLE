//Key = 1110000011000101100001111110110101010110000111001101110110000101


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267;

INV_X2 U1279 ( .A(n1862), .ZN(n1848) );
INV_X2 U1280 ( .A(U280), .ZN(n1849) );
INV_X1 U1281 ( .A(n1708), .ZN(U375) );
NAND2_X1 U1282 ( .A1(n1709), .A2(n1710), .ZN(U344) );
NAND2_X1 U1283 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1711), .ZN(n1710) );
NAND2_X1 U1284 ( .A1(n1712), .A2(DATA_IN_7_), .ZN(n1709) );
NAND2_X1 U1285 ( .A1(n1713), .A2(n1714), .ZN(U343) );
NAND2_X1 U1286 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1711), .ZN(n1714) );
XOR2_X1 U1287 ( .A(n1715), .B(KEYINPUT30), .Z(n1713) );
NAND2_X1 U1288 ( .A1(n1712), .A2(DATA_IN_6_), .ZN(n1715) );
NAND2_X1 U1289 ( .A1(n1716), .A2(n1717), .ZN(U342) );
NAND2_X1 U1290 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1711), .ZN(n1717) );
NAND2_X1 U1291 ( .A1(n1712), .A2(DATA_IN_5_), .ZN(n1716) );
NAND2_X1 U1292 ( .A1(n1718), .A2(n1719), .ZN(U341) );
NAND2_X1 U1293 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1711), .ZN(n1719) );
XOR2_X1 U1294 ( .A(KEYINPUT55), .B(n1720), .Z(n1718) );
NOR2_X1 U1295 ( .A1(n1721), .A2(n1711), .ZN(n1720) );
NAND2_X1 U1296 ( .A1(n1722), .A2(n1723), .ZN(U340) );
NAND2_X1 U1297 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1711), .ZN(n1723) );
NAND2_X1 U1298 ( .A1(n1712), .A2(DATA_IN_3_), .ZN(n1722) );
NAND2_X1 U1299 ( .A1(n1724), .A2(n1725), .ZN(U339) );
NAND2_X1 U1300 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1711), .ZN(n1725) );
NAND2_X1 U1301 ( .A1(n1712), .A2(DATA_IN_2_), .ZN(n1724) );
NAND2_X1 U1302 ( .A1(n1726), .A2(n1727), .ZN(U338) );
NAND2_X1 U1303 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1711), .ZN(n1727) );
NAND2_X1 U1304 ( .A1(n1712), .A2(DATA_IN_1_), .ZN(n1726) );
NAND2_X1 U1305 ( .A1(n1728), .A2(n1729), .ZN(U337) );
NAND2_X1 U1306 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1711), .ZN(n1729) );
NAND2_X1 U1307 ( .A1(n1712), .A2(DATA_IN_0_), .ZN(n1728) );
INV_X1 U1308 ( .A(n1711), .ZN(n1712) );
NAND2_X1 U1309 ( .A1(n1708), .A2(n1730), .ZN(n1711) );
NAND3_X1 U1310 ( .A1(n1731), .A2(n1732), .A3(n1733), .ZN(n1730) );
NAND2_X1 U1311 ( .A1(n1734), .A2(n1735), .ZN(U336) );
NAND2_X1 U1312 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1736), .ZN(n1735) );
NAND2_X1 U1313 ( .A1(n1737), .A2(DATA_IN_7_), .ZN(n1734) );
NAND2_X1 U1314 ( .A1(n1738), .A2(n1739), .ZN(U335) );
NAND2_X1 U1315 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1736), .ZN(n1739) );
NAND2_X1 U1316 ( .A1(n1737), .A2(DATA_IN_6_), .ZN(n1738) );
NAND2_X1 U1317 ( .A1(n1740), .A2(n1741), .ZN(U334) );
NAND2_X1 U1318 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1736), .ZN(n1741) );
NAND2_X1 U1319 ( .A1(n1737), .A2(DATA_IN_5_), .ZN(n1740) );
NAND2_X1 U1320 ( .A1(n1742), .A2(n1743), .ZN(U333) );
NAND2_X1 U1321 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1736), .ZN(n1743) );
NAND2_X1 U1322 ( .A1(n1737), .A2(DATA_IN_4_), .ZN(n1742) );
NAND2_X1 U1323 ( .A1(n1744), .A2(n1745), .ZN(U332) );
NAND2_X1 U1324 ( .A1(n1737), .A2(DATA_IN_3_), .ZN(n1745) );
NAND2_X1 U1325 ( .A1(n1746), .A2(n1736), .ZN(n1744) );
XOR2_X1 U1326 ( .A(n1747), .B(KEYINPUT48), .Z(n1746) );
NAND2_X1 U1327 ( .A1(n1748), .A2(n1749), .ZN(U331) );
NAND2_X1 U1328 ( .A1(n1737), .A2(DATA_IN_2_), .ZN(n1749) );
NAND2_X1 U1329 ( .A1(n1750), .A2(n1736), .ZN(n1748) );
XOR2_X1 U1330 ( .A(n1751), .B(KEYINPUT61), .Z(n1750) );
NAND2_X1 U1331 ( .A1(n1752), .A2(n1753), .ZN(U330) );
NAND2_X1 U1332 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1736), .ZN(n1753) );
NAND2_X1 U1333 ( .A1(n1737), .A2(DATA_IN_1_), .ZN(n1752) );
NAND2_X1 U1334 ( .A1(n1754), .A2(n1755), .ZN(U329) );
NAND2_X1 U1335 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1736), .ZN(n1755) );
NAND2_X1 U1336 ( .A1(n1737), .A2(DATA_IN_0_), .ZN(n1754) );
INV_X1 U1337 ( .A(n1736), .ZN(n1737) );
NAND2_X1 U1338 ( .A1(n1708), .A2(n1756), .ZN(n1736) );
NAND2_X1 U1339 ( .A1(n1757), .A2(n1732), .ZN(n1756) );
NAND3_X1 U1340 ( .A1(n1733), .A2(n1731), .A3(n1758), .ZN(n1757) );
NAND2_X1 U1341 ( .A1(n1759), .A2(n1760), .ZN(n1758) );
NAND3_X1 U1342 ( .A1(n1761), .A2(n1762), .A3(n1763), .ZN(n1760) );
OR2_X1 U1343 ( .A1(n1764), .A2(DATA_IN_7_), .ZN(n1763) );
NAND3_X1 U1344 ( .A1(n1765), .A2(n1766), .A3(n1767), .ZN(n1762) );
NAND2_X1 U1345 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1768), .ZN(n1767) );
NAND3_X1 U1346 ( .A1(n1769), .A2(n1770), .A3(n1771), .ZN(n1766) );
NAND2_X1 U1347 ( .A1(DATA_IN_5_), .A2(n1772), .ZN(n1771) );
NAND3_X1 U1348 ( .A1(n1773), .A2(n1774), .A3(n1775), .ZN(n1770) );
NAND2_X1 U1349 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1721), .ZN(n1775) );
NAND3_X1 U1350 ( .A1(n1776), .A2(n1777), .A3(n1778), .ZN(n1774) );
NAND2_X1 U1351 ( .A1(DATA_IN_3_), .A2(n1747), .ZN(n1778) );
NAND3_X1 U1352 ( .A1(n1779), .A2(n1780), .A3(n1781), .ZN(n1777) );
NAND2_X1 U1353 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1782), .ZN(n1781) );
NAND3_X1 U1354 ( .A1(n1783), .A2(n1784), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1780) );
INV_X1 U1355 ( .A(DATA_IN_0_), .ZN(n1784) );
NAND2_X1 U1356 ( .A1(DATA_IN_1_), .A2(n1785), .ZN(n1783) );
NAND2_X1 U1357 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1786), .ZN(n1779) );
NAND2_X1 U1358 ( .A1(DATA_IN_2_), .A2(n1751), .ZN(n1776) );
NAND2_X1 U1359 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1787), .ZN(n1773) );
NAND2_X1 U1360 ( .A1(DATA_IN_4_), .A2(n1788), .ZN(n1769) );
NAND2_X1 U1361 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1789), .ZN(n1765) );
XOR2_X1 U1362 ( .A(KEYINPUT51), .B(DATA_IN_5_), .Z(n1789) );
NAND2_X1 U1363 ( .A1(n1790), .A2(DATA_IN_6_), .ZN(n1761) );
XOR2_X1 U1364 ( .A(n1791), .B(KEYINPUT40), .Z(n1790) );
NAND2_X1 U1365 ( .A1(DATA_IN_7_), .A2(n1764), .ZN(n1759) );
NAND2_X1 U1366 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1792), .ZN(n1731) );
XOR2_X1 U1367 ( .A(KEYINPUT26), .B(DATA_IN_7_), .Z(n1792) );
NAND3_X1 U1368 ( .A1(n1793), .A2(n1794), .A3(n1795), .ZN(n1733) );
NAND2_X1 U1369 ( .A1(DATA_IN_7_), .A2(n1796), .ZN(n1795) );
NAND3_X1 U1370 ( .A1(n1797), .A2(n1798), .A3(n1799), .ZN(n1794) );
NAND2_X1 U1371 ( .A1(DATA_IN_6_), .A2(n1800), .ZN(n1799) );
NAND3_X1 U1372 ( .A1(n1801), .A2(n1802), .A3(n1803), .ZN(n1798) );
NAND2_X1 U1373 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1804), .ZN(n1803) );
NAND3_X1 U1374 ( .A1(n1805), .A2(n1806), .A3(n1807), .ZN(n1802) );
NAND2_X1 U1375 ( .A1(DATA_IN_4_), .A2(n1808), .ZN(n1807) );
NAND3_X1 U1376 ( .A1(n1809), .A2(n1810), .A3(n1811), .ZN(n1806) );
NAND2_X1 U1377 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1812), .ZN(n1811) );
XOR2_X1 U1378 ( .A(KEYINPUT43), .B(DATA_IN_3_), .Z(n1812) );
NAND3_X1 U1379 ( .A1(n1813), .A2(n1814), .A3(n1815), .ZN(n1810) );
NAND2_X1 U1380 ( .A1(DATA_IN_2_), .A2(n1816), .ZN(n1815) );
NAND3_X1 U1381 ( .A1(n1817), .A2(n1818), .A3(DATA_IN_0_), .ZN(n1814) );
INV_X1 U1382 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1818) );
NAND2_X1 U1383 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1786), .ZN(n1817) );
NAND2_X1 U1384 ( .A1(DATA_IN_1_), .A2(n1819), .ZN(n1813) );
NAND2_X1 U1385 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1820), .ZN(n1809) );
XOR2_X1 U1386 ( .A(KEYINPUT0), .B(DATA_IN_2_), .Z(n1820) );
NAND2_X1 U1387 ( .A1(DATA_IN_3_), .A2(n1821), .ZN(n1805) );
NAND2_X1 U1388 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1721), .ZN(n1801) );
NAND2_X1 U1389 ( .A1(DATA_IN_5_), .A2(n1822), .ZN(n1797) );
NAND2_X1 U1390 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1768), .ZN(n1793) );
NAND2_X1 U1391 ( .A1(n1823), .A2(n1824), .ZN(U328) );
NAND2_X1 U1392 ( .A1(n1825), .A2(DATA_IN_7_), .ZN(n1824) );
NAND2_X1 U1393 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1826), .ZN(n1823) );
NAND2_X1 U1394 ( .A1(n1827), .A2(n1828), .ZN(U327) );
NAND2_X1 U1395 ( .A1(n1825), .A2(DATA_IN_6_), .ZN(n1828) );
NAND2_X1 U1396 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1826), .ZN(n1827) );
NAND2_X1 U1397 ( .A1(n1829), .A2(n1830), .ZN(U326) );
NAND2_X1 U1398 ( .A1(n1825), .A2(DATA_IN_5_), .ZN(n1830) );
NAND2_X1 U1399 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1826), .ZN(n1829) );
NAND2_X1 U1400 ( .A1(n1831), .A2(n1832), .ZN(U325) );
NAND2_X1 U1401 ( .A1(n1825), .A2(DATA_IN_4_), .ZN(n1832) );
NAND2_X1 U1402 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1826), .ZN(n1831) );
NAND2_X1 U1403 ( .A1(n1833), .A2(n1834), .ZN(U324) );
NAND2_X1 U1404 ( .A1(n1825), .A2(DATA_IN_3_), .ZN(n1834) );
NAND2_X1 U1405 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1826), .ZN(n1833) );
NAND2_X1 U1406 ( .A1(n1835), .A2(n1836), .ZN(U323) );
NAND2_X1 U1407 ( .A1(n1825), .A2(DATA_IN_2_), .ZN(n1836) );
XOR2_X1 U1408 ( .A(n1837), .B(KEYINPUT10), .Z(n1835) );
NAND2_X1 U1409 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1826), .ZN(n1837) );
NAND2_X1 U1410 ( .A1(n1838), .A2(n1839), .ZN(U322) );
NAND2_X1 U1411 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1826), .ZN(n1839) );
XOR2_X1 U1412 ( .A(n1840), .B(KEYINPUT11), .Z(n1838) );
NAND2_X1 U1413 ( .A1(n1825), .A2(DATA_IN_1_), .ZN(n1840) );
NAND2_X1 U1414 ( .A1(n1841), .A2(n1842), .ZN(U321) );
NAND2_X1 U1415 ( .A1(n1825), .A2(DATA_IN_0_), .ZN(n1842) );
AND2_X1 U1416 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1843), .ZN(n1825) );
NAND2_X1 U1417 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1826), .ZN(n1841) );
NAND2_X1 U1418 ( .A1(n1708), .A2(n1843), .ZN(n1826) );
NAND2_X1 U1419 ( .A1(n1732), .A2(n1844), .ZN(n1843) );
NAND2_X1 U1420 ( .A1(n1732), .A2(n1845), .ZN(n1708) );
NAND2_X1 U1421 ( .A1(n1846), .A2(n1847), .ZN(U320) );
NAND2_X1 U1422 ( .A1(n1848), .A2(DATA_IN_7_), .ZN(n1847) );
NAND2_X1 U1423 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1849), .ZN(n1846) );
NAND2_X1 U1424 ( .A1(n1850), .A2(n1851), .ZN(U319) );
NAND2_X1 U1425 ( .A1(n1848), .A2(DATA_IN_6_), .ZN(n1851) );
NAND2_X1 U1426 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1849), .ZN(n1850) );
NAND2_X1 U1427 ( .A1(n1852), .A2(n1853), .ZN(U318) );
NAND2_X1 U1428 ( .A1(DATA_IN_5_), .A2(n1854), .ZN(n1853) );
XOR2_X1 U1429 ( .A(KEYINPUT62), .B(n1848), .Z(n1854) );
NAND2_X1 U1430 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1849), .ZN(n1852) );
NAND2_X1 U1431 ( .A1(n1855), .A2(n1856), .ZN(U317) );
NAND2_X1 U1432 ( .A1(n1848), .A2(DATA_IN_4_), .ZN(n1856) );
NAND2_X1 U1433 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1849), .ZN(n1855) );
NAND2_X1 U1434 ( .A1(n1857), .A2(n1858), .ZN(U316) );
NAND2_X1 U1435 ( .A1(n1848), .A2(DATA_IN_3_), .ZN(n1858) );
NAND2_X1 U1436 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1849), .ZN(n1857) );
NAND2_X1 U1437 ( .A1(n1859), .A2(n1860), .ZN(U315) );
NAND2_X1 U1438 ( .A1(n1861), .A2(DATA_IN_2_), .ZN(n1860) );
XOR2_X1 U1439 ( .A(n1862), .B(KEYINPUT8), .Z(n1861) );
NAND2_X1 U1440 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1863), .ZN(n1859) );
XOR2_X1 U1441 ( .A(KEYINPUT46), .B(n1849), .Z(n1863) );
NAND2_X1 U1442 ( .A1(n1864), .A2(n1865), .ZN(U314) );
NAND2_X1 U1443 ( .A1(n1848), .A2(DATA_IN_1_), .ZN(n1865) );
NAND2_X1 U1444 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1849), .ZN(n1864) );
NAND2_X1 U1445 ( .A1(n1866), .A2(n1867), .ZN(U313) );
NAND2_X1 U1446 ( .A1(n1848), .A2(DATA_IN_0_), .ZN(n1867) );
NAND2_X1 U1447 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1849), .ZN(n1866) );
NAND2_X1 U1448 ( .A1(n1868), .A2(n1869), .ZN(U312) );
NAND2_X1 U1449 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1848), .ZN(n1869) );
NAND2_X1 U1450 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1849), .ZN(n1868) );
NAND2_X1 U1451 ( .A1(n1870), .A2(n1871), .ZN(U311) );
NAND2_X1 U1452 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1848), .ZN(n1871) );
NAND2_X1 U1453 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1849), .ZN(n1870) );
NAND2_X1 U1454 ( .A1(n1872), .A2(n1873), .ZN(U310) );
NAND2_X1 U1455 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1848), .ZN(n1873) );
NAND2_X1 U1456 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1849), .ZN(n1872) );
NAND2_X1 U1457 ( .A1(n1874), .A2(n1875), .ZN(U309) );
NAND2_X1 U1458 ( .A1(n1876), .A2(n1849), .ZN(n1875) );
XOR2_X1 U1459 ( .A(REG2_REG_4__SCAN_IN), .B(KEYINPUT39), .Z(n1876) );
NAND2_X1 U1460 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1848), .ZN(n1874) );
NAND2_X1 U1461 ( .A1(n1877), .A2(n1878), .ZN(U308) );
NAND2_X1 U1462 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1848), .ZN(n1878) );
XOR2_X1 U1463 ( .A(KEYINPUT29), .B(n1879), .Z(n1877) );
AND2_X1 U1464 ( .A1(n1849), .A2(REG2_REG_3__SCAN_IN), .ZN(n1879) );
NAND2_X1 U1465 ( .A1(n1880), .A2(n1881), .ZN(U307) );
NAND2_X1 U1466 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1848), .ZN(n1881) );
NAND2_X1 U1467 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1849), .ZN(n1880) );
NAND2_X1 U1468 ( .A1(n1882), .A2(n1883), .ZN(U306) );
NAND2_X1 U1469 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1848), .ZN(n1883) );
NAND2_X1 U1470 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1849), .ZN(n1882) );
NAND2_X1 U1471 ( .A1(n1884), .A2(n1885), .ZN(U305) );
NAND2_X1 U1472 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1848), .ZN(n1885) );
NAND2_X1 U1473 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1849), .ZN(n1884) );
NAND2_X1 U1474 ( .A1(n1886), .A2(n1887), .ZN(U304) );
NAND2_X1 U1475 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1888), .ZN(n1887) );
XOR2_X1 U1476 ( .A(KEYINPUT60), .B(n1849), .Z(n1888) );
NAND2_X1 U1477 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1848), .ZN(n1886) );
NAND2_X1 U1478 ( .A1(n1889), .A2(n1890), .ZN(U303) );
NAND2_X1 U1479 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1848), .ZN(n1890) );
NAND2_X1 U1480 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1849), .ZN(n1889) );
NAND2_X1 U1481 ( .A1(n1891), .A2(n1892), .ZN(U302) );
NAND2_X1 U1482 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1848), .ZN(n1892) );
NAND2_X1 U1483 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1849), .ZN(n1891) );
NAND2_X1 U1484 ( .A1(n1893), .A2(n1894), .ZN(U301) );
NAND2_X1 U1485 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1848), .ZN(n1894) );
NAND2_X1 U1486 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1849), .ZN(n1893) );
NAND2_X1 U1487 ( .A1(n1895), .A2(n1896), .ZN(U300) );
NAND2_X1 U1488 ( .A1(n1848), .A2(n1897), .ZN(n1896) );
XOR2_X1 U1489 ( .A(REG2_REG_3__SCAN_IN), .B(KEYINPUT27), .Z(n1897) );
NAND2_X1 U1490 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1849), .ZN(n1895) );
NAND2_X1 U1491 ( .A1(n1898), .A2(n1899), .ZN(U299) );
NAND2_X1 U1492 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1848), .ZN(n1899) );
NAND2_X1 U1493 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1849), .ZN(n1898) );
NAND2_X1 U1494 ( .A1(n1900), .A2(n1901), .ZN(U298) );
NAND2_X1 U1495 ( .A1(n1902), .A2(n1849), .ZN(n1901) );
XOR2_X1 U1496 ( .A(REG3_REG_1__SCAN_IN), .B(KEYINPUT20), .Z(n1902) );
NAND2_X1 U1497 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1848), .ZN(n1900) );
NAND2_X1 U1498 ( .A1(n1903), .A2(n1904), .ZN(U297) );
NAND2_X1 U1499 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1848), .ZN(n1904) );
NAND2_X1 U1500 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1849), .ZN(n1903) );
NAND2_X1 U1501 ( .A1(n1905), .A2(n1906), .ZN(U296) );
NAND2_X1 U1502 ( .A1(n1907), .A2(REG3_REG_7__SCAN_IN), .ZN(n1906) );
XOR2_X1 U1503 ( .A(n1862), .B(KEYINPUT56), .Z(n1907) );
NAND2_X1 U1504 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1849), .ZN(n1905) );
NAND2_X1 U1505 ( .A1(n1908), .A2(n1909), .ZN(U295) );
NAND2_X1 U1506 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1910), .ZN(n1909) );
XOR2_X1 U1507 ( .A(KEYINPUT4), .B(n1848), .Z(n1910) );
NAND2_X1 U1508 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1849), .ZN(n1908) );
NAND2_X1 U1509 ( .A1(n1911), .A2(n1912), .ZN(U294) );
NAND2_X1 U1510 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1848), .ZN(n1912) );
NAND2_X1 U1511 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1849), .ZN(n1911) );
NAND2_X1 U1512 ( .A1(n1913), .A2(n1914), .ZN(U293) );
NAND2_X1 U1513 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1849), .ZN(n1914) );
XOR2_X1 U1514 ( .A(KEYINPUT35), .B(n1915), .Z(n1913) );
AND2_X1 U1515 ( .A1(n1848), .A2(REG3_REG_4__SCAN_IN), .ZN(n1915) );
NAND2_X1 U1516 ( .A1(n1916), .A2(n1917), .ZN(U292) );
NAND2_X1 U1517 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1918), .ZN(n1917) );
XOR2_X1 U1518 ( .A(KEYINPUT32), .B(n1849), .Z(n1918) );
NAND2_X1 U1519 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1848), .ZN(n1916) );
NAND2_X1 U1520 ( .A1(n1919), .A2(n1920), .ZN(U291) );
NAND2_X1 U1521 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1849), .ZN(n1920) );
XOR2_X1 U1522 ( .A(KEYINPUT44), .B(n1921), .Z(n1919) );
AND2_X1 U1523 ( .A1(n1848), .A2(REG3_REG_2__SCAN_IN), .ZN(n1921) );
NAND2_X1 U1524 ( .A1(n1922), .A2(n1923), .ZN(U290) );
NAND2_X1 U1525 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1848), .ZN(n1923) );
NAND2_X1 U1526 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1849), .ZN(n1922) );
NAND2_X1 U1527 ( .A1(n1924), .A2(n1925), .ZN(U289) );
NAND2_X1 U1528 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1848), .ZN(n1925) );
XOR2_X1 U1529 ( .A(n1926), .B(KEYINPUT5), .Z(n1924) );
NAND2_X1 U1530 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1849), .ZN(n1926) );
NAND4_X1 U1531 ( .A1(n1927), .A2(n1928), .A3(n1929), .A4(n1930), .ZN(U288));
NAND2_X1 U1532 ( .A1(n1931), .A2(n1932), .ZN(n1930) );
XNOR2_X1 U1533 ( .A(n1933), .B(KEYINPUT63), .ZN(n1931) );
NAND2_X1 U1534 ( .A1(n1934), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1929) );
NAND2_X1 U1535 ( .A1(n1935), .A2(REG4_REG_7__SCAN_IN), .ZN(n1928) );
NAND2_X1 U1536 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1849), .ZN(n1927) );
NAND4_X1 U1537 ( .A1(n1936), .A2(n1937), .A3(n1938), .A4(n1939), .ZN(U287));
NAND2_X1 U1538 ( .A1(n1934), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1939) );
NOR2_X1 U1539 ( .A1(n1940), .A2(n1941), .ZN(n1938) );
NOR2_X1 U1540 ( .A1(n1942), .A2(n1943), .ZN(n1941) );
NOR2_X1 U1541 ( .A1(n1933), .A2(n1944), .ZN(n1942) );
XOR2_X1 U1542 ( .A(KEYINPUT18), .B(n1945), .Z(n1944) );
NOR2_X1 U1543 ( .A1(n1946), .A2(n1947), .ZN(n1945) );
AND2_X1 U1544 ( .A1(n1948), .A2(n1947), .ZN(n1933) );
XOR2_X1 U1545 ( .A(n1949), .B(KEYINPUT13), .Z(n1948) );
AND4_X1 U1546 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(n1940));
NAND2_X1 U1547 ( .A1(n1935), .A2(REG4_REG_6__SCAN_IN), .ZN(n1937) );
NAND2_X1 U1548 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1849), .ZN(n1936) );
NAND4_X1 U1549 ( .A1(n1954), .A2(n1955), .A3(n1956), .A4(n1957), .ZN(U286));
NOR3_X1 U1550 ( .A1(n1958), .A2(n1959), .A3(n1960), .ZN(n1957) );
NOR2_X1 U1551 ( .A1(n1961), .A2(n1962), .ZN(n1960) );
XOR2_X1 U1552 ( .A(n1963), .B(n1950), .Z(n1962) );
XOR2_X1 U1553 ( .A(n1964), .B(n1965), .Z(n1950) );
NAND2_X1 U1554 ( .A1(KEYINPUT2), .A2(n1951), .ZN(n1964) );
NOR2_X1 U1555 ( .A1(n1952), .A2(KEYINPUT57), .ZN(n1963) );
NOR3_X1 U1556 ( .A1(n1943), .A2(n1966), .A3(n1967), .ZN(n1959) );
NOR3_X1 U1557 ( .A1(n1968), .A2(n1969), .A3(n1946), .ZN(n1967) );
AND2_X1 U1558 ( .A1(n1970), .A2(n1951), .ZN(n1968) );
INV_X1 U1559 ( .A(n1947), .ZN(n1966) );
NAND2_X1 U1560 ( .A1(n1969), .A2(n1971), .ZN(n1947) );
NAND2_X1 U1561 ( .A1(n1972), .A2(n1949), .ZN(n1971) );
INV_X1 U1562 ( .A(n1946), .ZN(n1949) );
NOR2_X1 U1563 ( .A1(n1970), .A2(n1951), .ZN(n1946) );
NAND2_X1 U1564 ( .A1(n1951), .A2(n1970), .ZN(n1972) );
INV_X1 U1565 ( .A(n1973), .ZN(n1951) );
NOR2_X1 U1566 ( .A1(n1973), .A2(n1974), .ZN(n1958) );
NAND2_X1 U1567 ( .A1(n1975), .A2(n1976), .ZN(n1973) );
NAND2_X1 U1568 ( .A1(n1977), .A2(n1978), .ZN(n1976) );
NAND2_X1 U1569 ( .A1(n1979), .A2(n1980), .ZN(n1978) );
XNOR2_X1 U1570 ( .A(n1981), .B(KEYINPUT38), .ZN(n1980) );
NAND2_X1 U1571 ( .A1(n1982), .A2(n1983), .ZN(n1977) );
NAND2_X1 U1572 ( .A1(n1984), .A2(n1985), .ZN(n1983) );
XNOR2_X1 U1573 ( .A(KEYINPUT42), .B(n1986), .ZN(n1984) );
NAND4_X1 U1574 ( .A1(n1979), .A2(n1981), .A3(n1987), .A4(n1982), .ZN(n1975));
NAND2_X1 U1575 ( .A1(n1988), .A2(n1989), .ZN(n1982) );
NAND2_X1 U1576 ( .A1(n1986), .A2(n1990), .ZN(n1988) );
OR2_X1 U1577 ( .A1(n1990), .A2(n1986), .ZN(n1987) );
AND2_X1 U1578 ( .A1(n1991), .A2(n1992), .ZN(n1981) );
NAND3_X1 U1579 ( .A1(DATA_IN_6_), .A2(n1993), .A3(n1994), .ZN(n1992) );
NAND3_X1 U1580 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1791), .A3(RESTART), .ZN(n1991) );
AND2_X1 U1581 ( .A1(n1995), .A2(n1996), .ZN(n1979) );
NAND3_X1 U1582 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1768), .A3(n1994), .ZN(n1996) );
NAND3_X1 U1583 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1800), .A3(RESTART), .ZN(n1995) );
NAND2_X1 U1584 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1849), .ZN(n1956) );
NAND2_X1 U1585 ( .A1(n1934), .A2(RLAST_REG_5__SCAN_IN), .ZN(n1955) );
NAND2_X1 U1586 ( .A1(n1935), .A2(REG4_REG_5__SCAN_IN), .ZN(n1954) );
NAND4_X1 U1587 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(U285));
NOR3_X1 U1588 ( .A1(n2001), .A2(n2002), .A3(n2003), .ZN(n2000) );
NOR3_X1 U1589 ( .A1(n1961), .A2(n2004), .A3(n1952), .ZN(n2003) );
AND3_X1 U1590 ( .A1(n2005), .A2(n2006), .A3(n2007), .ZN(n1952) );
NAND2_X1 U1591 ( .A1(n2008), .A2(n1965), .ZN(n2005) );
NAND2_X1 U1592 ( .A1(n2009), .A2(n2010), .ZN(n1965) );
XOR2_X1 U1593 ( .A(KEYINPUT54), .B(n2011), .Z(n2010) );
NOR2_X1 U1594 ( .A1(n2012), .A2(n2013), .ZN(n2004) );
INV_X1 U1595 ( .A(n2008), .ZN(n2013) );
NAND2_X1 U1596 ( .A1(n2014), .A2(n2015), .ZN(n2008) );
NOR2_X1 U1597 ( .A1(n2016), .A2(n2017), .ZN(n2012) );
XOR2_X1 U1598 ( .A(n2006), .B(KEYINPUT28), .Z(n2016) );
NOR3_X1 U1599 ( .A1(n1943), .A2(n1969), .A3(n2018), .ZN(n2002) );
NOR2_X1 U1600 ( .A1(n2019), .A2(n2020), .ZN(n2018) );
AND2_X1 U1601 ( .A1(n2021), .A2(n2022), .ZN(n2019) );
AND3_X1 U1602 ( .A1(n2020), .A2(n2021), .A3(n2022), .ZN(n1969) );
NAND2_X1 U1603 ( .A1(n1970), .A2(n2023), .ZN(n2020) );
NAND2_X1 U1604 ( .A1(n2014), .A2(n2024), .ZN(n2023) );
NAND3_X1 U1605 ( .A1(n2025), .A2(n2011), .A3(n2026), .ZN(n1970) );
NOR2_X1 U1606 ( .A1(n2011), .A2(n1974), .ZN(n2001) );
INV_X1 U1607 ( .A(n2014), .ZN(n2011) );
XOR2_X1 U1608 ( .A(n2027), .B(n2028), .Z(n2014) );
NOR2_X1 U1609 ( .A1(KEYINPUT47), .A2(n1986), .ZN(n2028) );
NAND2_X1 U1610 ( .A1(n2029), .A2(n2030), .ZN(n1986) );
NAND2_X1 U1611 ( .A1(RESTART), .A2(n1772), .ZN(n2030) );
NAND2_X1 U1612 ( .A1(n2031), .A2(n1994), .ZN(n2029) );
XOR2_X1 U1613 ( .A(n1989), .B(n1985), .Z(n2027) );
INV_X1 U1614 ( .A(n1990), .ZN(n1985) );
NAND2_X1 U1615 ( .A1(n2032), .A2(n2033), .ZN(n1990) );
NAND2_X1 U1616 ( .A1(n2034), .A2(n1994), .ZN(n2033) );
NAND2_X1 U1617 ( .A1(KEYINPUT45), .A2(DATA_IN_5_), .ZN(n2034) );
NAND2_X1 U1618 ( .A1(n2035), .A2(n1822), .ZN(n2032) );
NAND2_X1 U1619 ( .A1(DATA_IN_5_), .A2(n2036), .ZN(n2035) );
NAND2_X1 U1620 ( .A1(KEYINPUT45), .A2(RESTART), .ZN(n2036) );
NAND2_X1 U1621 ( .A1(n2037), .A2(n2038), .ZN(n1989) );
NAND2_X1 U1622 ( .A1(n2039), .A2(n2040), .ZN(n2038) );
NAND2_X1 U1623 ( .A1(n2041), .A2(n2042), .ZN(n2040) );
NAND2_X1 U1624 ( .A1(n2043), .A2(n2044), .ZN(n2037) );
NAND2_X1 U1625 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1849), .ZN(n1999) );
NAND2_X1 U1626 ( .A1(n1934), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1998) );
NAND2_X1 U1627 ( .A1(n1935), .A2(REG4_REG_4__SCAN_IN), .ZN(n1997) );
NAND4_X1 U1628 ( .A1(n2045), .A2(n2046), .A3(n2047), .A4(n2048), .ZN(U284));
NOR3_X1 U1629 ( .A1(n2049), .A2(n2050), .A3(n2051), .ZN(n2048) );
NOR2_X1 U1630 ( .A1(n1961), .A2(n2052), .ZN(n2051) );
XOR2_X1 U1631 ( .A(n2017), .B(n2006), .Z(n2052) );
NAND2_X1 U1632 ( .A1(n2015), .A2(n2053), .ZN(n2006) );
NAND2_X1 U1633 ( .A1(n2054), .A2(n2055), .ZN(n2053) );
INV_X1 U1634 ( .A(n2009), .ZN(n2015) );
NOR2_X1 U1635 ( .A1(n2054), .A2(n2055), .ZN(n2009) );
NOR2_X1 U1636 ( .A1(n1943), .A2(n2056), .ZN(n2050) );
XNOR2_X1 U1637 ( .A(n2022), .B(n2021), .ZN(n2056) );
NAND2_X1 U1638 ( .A1(n2057), .A2(n2024), .ZN(n2021) );
NAND2_X1 U1639 ( .A1(n2026), .A2(n2025), .ZN(n2024) );
XOR2_X1 U1640 ( .A(n2058), .B(KEYINPUT17), .Z(n2057) );
OR2_X1 U1641 ( .A1(n2026), .A2(n2025), .ZN(n2058) );
NOR2_X1 U1642 ( .A1(n2025), .A2(n1974), .ZN(n2049) );
INV_X1 U1643 ( .A(n2055), .ZN(n2025) );
NAND2_X1 U1644 ( .A1(n2059), .A2(n2060), .ZN(n2055) );
NAND4_X1 U1645 ( .A1(n2043), .A2(n2061), .A3(n2062), .A4(n2063), .ZN(n2060));
OR2_X1 U1646 ( .A1(n2064), .A2(KEYINPUT23), .ZN(n2063) );
NAND3_X1 U1647 ( .A1(n2064), .A2(n2044), .A3(KEYINPUT23), .ZN(n2062) );
INV_X1 U1648 ( .A(n2041), .ZN(n2044) );
XOR2_X1 U1649 ( .A(KEYINPUT15), .B(n2065), .Z(n2059) );
NOR2_X1 U1650 ( .A1(n2043), .A2(n2066), .ZN(n2065) );
NOR2_X1 U1651 ( .A1(n2067), .A2(n2068), .ZN(n2066) );
INV_X1 U1652 ( .A(n2061), .ZN(n2068) );
NAND2_X1 U1653 ( .A1(n2039), .A2(n2041), .ZN(n2061) );
INV_X1 U1654 ( .A(n2064), .ZN(n2039) );
NOR2_X1 U1655 ( .A1(n2041), .A2(n2069), .ZN(n2067) );
XOR2_X1 U1656 ( .A(n2064), .B(KEYINPUT23), .Z(n2069) );
NAND2_X1 U1657 ( .A1(n2070), .A2(n2071), .ZN(n2064) );
NAND2_X1 U1658 ( .A1(RESTART), .A2(n1788), .ZN(n2071) );
OR2_X1 U1659 ( .A1(REG4_REG_4__SCAN_IN), .A2(RESTART), .ZN(n2070) );
NAND2_X1 U1660 ( .A1(n2072), .A2(n2073), .ZN(n2041) );
NAND2_X1 U1661 ( .A1(RESTART), .A2(n1808), .ZN(n2073) );
NAND2_X1 U1662 ( .A1(n1721), .A2(n1994), .ZN(n2072) );
INV_X1 U1663 ( .A(n2042), .ZN(n2043) );
NAND2_X1 U1664 ( .A1(n2074), .A2(n2075), .ZN(n2042) );
NAND2_X1 U1665 ( .A1(n2076), .A2(n2077), .ZN(n2075) );
NAND2_X1 U1666 ( .A1(n2078), .A2(n2079), .ZN(n2076) );
INV_X1 U1667 ( .A(n2080), .ZN(n2079) );
XNOR2_X1 U1668 ( .A(KEYINPUT36), .B(n2081), .ZN(n2078) );
NAND2_X1 U1669 ( .A1(n2081), .A2(n2080), .ZN(n2074) );
NAND2_X1 U1670 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1849), .ZN(n2047) );
NAND2_X1 U1671 ( .A1(n1934), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2046) );
NAND2_X1 U1672 ( .A1(n1935), .A2(REG4_REG_3__SCAN_IN), .ZN(n2045) );
NAND4_X1 U1673 ( .A1(n2082), .A2(n2083), .A3(n2084), .A4(n2085), .ZN(U283));
NOR3_X1 U1674 ( .A1(n2086), .A2(n2087), .A3(n2088), .ZN(n2085) );
NOR3_X1 U1675 ( .A1(n1961), .A2(n2007), .A3(n2089), .ZN(n2088) );
NOR2_X1 U1676 ( .A1(n2090), .A2(n2091), .ZN(n2089) );
NOR2_X1 U1677 ( .A1(n2092), .A2(n2093), .ZN(n2090) );
XOR2_X1 U1678 ( .A(n2094), .B(KEYINPUT49), .Z(n2093) );
INV_X1 U1679 ( .A(n2017), .ZN(n2007) );
NAND3_X1 U1680 ( .A1(n2095), .A2(n2094), .A3(n2091), .ZN(n2017) );
NAND3_X1 U1681 ( .A1(n2096), .A2(n2097), .A3(n2054), .ZN(n2091) );
NAND2_X1 U1682 ( .A1(n2098), .A2(n2099), .ZN(n2054) );
OR2_X1 U1683 ( .A1(n2100), .A2(KEYINPUT53), .ZN(n2097) );
NAND3_X1 U1684 ( .A1(n2100), .A2(n2101), .A3(KEYINPUT53), .ZN(n2096) );
NOR3_X1 U1685 ( .A1(n1943), .A2(n2022), .A3(n2102), .ZN(n2087) );
NOR3_X1 U1686 ( .A1(n2100), .A2(n2026), .A3(n2103), .ZN(n2102) );
AND2_X1 U1687 ( .A1(n2094), .A2(n2104), .ZN(n2103) );
NOR2_X1 U1688 ( .A1(n2100), .A2(n2105), .ZN(n2026) );
AND4_X1 U1689 ( .A1(n2104), .A2(n2094), .A3(n2106), .A4(n2107), .ZN(n2022));
NAND2_X1 U1690 ( .A1(n2099), .A2(n2100), .ZN(n2107) );
INV_X1 U1691 ( .A(n2098), .ZN(n2100) );
NAND2_X1 U1692 ( .A1(n2098), .A2(n2105), .ZN(n2106) );
XNOR2_X1 U1693 ( .A(n2099), .B(KEYINPUT34), .ZN(n2105) );
NOR2_X1 U1694 ( .A1(n2108), .A2(n2109), .ZN(n2086) );
XOR2_X1 U1695 ( .A(REG4_REG_2__SCAN_IN), .B(KEYINPUT37), .Z(n2109) );
NAND2_X1 U1696 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1849), .ZN(n2084) );
NAND2_X1 U1697 ( .A1(n2110), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2083) );
XNOR2_X1 U1698 ( .A(n1934), .B(KEYINPUT52), .ZN(n2110) );
OR2_X1 U1699 ( .A1(n1974), .A2(n2098), .ZN(n2082) );
XOR2_X1 U1700 ( .A(n2080), .B(n2111), .Z(n2098) );
NOR2_X1 U1701 ( .A1(n2112), .A2(n2113), .ZN(n2111) );
NOR3_X1 U1702 ( .A1(n2077), .A2(KEYINPUT19), .A3(n2081), .ZN(n2113) );
AND2_X1 U1703 ( .A1(n2077), .A2(n2081), .ZN(n2112) );
NAND2_X1 U1704 ( .A1(n2114), .A2(n2115), .ZN(n2081) );
NAND2_X1 U1705 ( .A1(RESTART), .A2(n1821), .ZN(n2115) );
NAND2_X1 U1706 ( .A1(n1787), .A2(n1994), .ZN(n2114) );
NAND2_X1 U1707 ( .A1(n2116), .A2(n2117), .ZN(n2077) );
NAND2_X1 U1708 ( .A1(n2118), .A2(n2119), .ZN(n2117) );
NAND2_X1 U1709 ( .A1(n2120), .A2(n2121), .ZN(n2116) );
NAND2_X1 U1710 ( .A1(n2122), .A2(n2123), .ZN(n2080) );
NAND2_X1 U1711 ( .A1(RESTART), .A2(n1747), .ZN(n2123) );
NAND2_X1 U1712 ( .A1(n2124), .A2(n1994), .ZN(n2122) );
NAND4_X1 U1713 ( .A1(n2125), .A2(n2126), .A3(n2127), .A4(n2128), .ZN(U282));
NOR3_X1 U1714 ( .A1(n2129), .A2(n2130), .A3(n2131), .ZN(n2128) );
NOR2_X1 U1715 ( .A1(n1961), .A2(n2132), .ZN(n2131) );
XNOR2_X1 U1716 ( .A(n2094), .B(n2133), .ZN(n2132) );
NOR2_X1 U1717 ( .A1(n2092), .A2(KEYINPUT50), .ZN(n2133) );
INV_X1 U1718 ( .A(n2095), .ZN(n2092) );
NAND2_X1 U1719 ( .A1(n2101), .A2(n2134), .ZN(n2095) );
NAND2_X1 U1720 ( .A1(n2135), .A2(n2136), .ZN(n2134) );
XOR2_X1 U1721 ( .A(n2137), .B(KEYINPUT31), .Z(n2135) );
NOR2_X1 U1722 ( .A1(n2138), .A2(n1943), .ZN(n2130) );
XNOR2_X1 U1723 ( .A(n2104), .B(n2094), .ZN(n2138) );
NAND2_X1 U1724 ( .A1(n2101), .A2(n2139), .ZN(n2104) );
NAND2_X1 U1725 ( .A1(n2140), .A2(n2136), .ZN(n2139) );
INV_X1 U1726 ( .A(n2099), .ZN(n2101) );
NOR2_X1 U1727 ( .A1(n2136), .A2(n2140), .ZN(n2099) );
INV_X1 U1728 ( .A(n2137), .ZN(n2140) );
NOR2_X1 U1729 ( .A1(n2137), .A2(n1974), .ZN(n2129) );
XNOR2_X1 U1730 ( .A(n2141), .B(n2118), .ZN(n2137) );
NAND2_X1 U1731 ( .A1(n2142), .A2(n2143), .ZN(n2118) );
NAND2_X1 U1732 ( .A1(RESTART), .A2(n1751), .ZN(n2143) );
INV_X1 U1733 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1751) );
NAND2_X1 U1734 ( .A1(n2144), .A2(n1994), .ZN(n2142) );
NAND2_X1 U1735 ( .A1(n2119), .A2(n2145), .ZN(n2141) );
NAND2_X1 U1736 ( .A1(n2146), .A2(n2121), .ZN(n2145) );
NAND2_X1 U1737 ( .A1(KEYINPUT16), .A2(n2147), .ZN(n2146) );
NAND2_X1 U1738 ( .A1(n2147), .A2(n2148), .ZN(n2119) );
INV_X1 U1739 ( .A(n2121), .ZN(n2148) );
NAND2_X1 U1740 ( .A1(n2149), .A2(n2150), .ZN(n2121) );
OR2_X1 U1741 ( .A1(n2151), .A2(n2152), .ZN(n2150) );
NAND2_X1 U1742 ( .A1(n2153), .A2(n2154), .ZN(n2149) );
INV_X1 U1743 ( .A(n2120), .ZN(n2147) );
NAND2_X1 U1744 ( .A1(n2155), .A2(n2156), .ZN(n2120) );
NAND2_X1 U1745 ( .A1(RESTART), .A2(n1816), .ZN(n2156) );
NAND2_X1 U1746 ( .A1(n1782), .A2(n1994), .ZN(n2155) );
NAND2_X1 U1747 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1849), .ZN(n2127) );
NAND2_X1 U1748 ( .A1(n1934), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2126) );
NAND2_X1 U1749 ( .A1(n1935), .A2(REG4_REG_1__SCAN_IN), .ZN(n2125) );
NAND3_X1 U1750 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(U281) );
NOR3_X1 U1751 ( .A1(n2160), .A2(n2161), .A3(n2162), .ZN(n2159) );
AND2_X1 U1752 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1934), .ZN(n2162) );
AND3_X1 U1753 ( .A1(n1844), .A2(n1994), .A3(n2163), .ZN(n1934) );
INV_X1 U1754 ( .A(ENABLE), .ZN(n1844) );
NOR2_X1 U1755 ( .A1(n2164), .A2(n2094), .ZN(n2161) );
NAND2_X1 U1756 ( .A1(n2136), .A2(n2165), .ZN(n2094) );
NAND3_X1 U1757 ( .A1(n2166), .A2(n2167), .A3(n2168), .ZN(n2165) );
NAND2_X1 U1758 ( .A1(n2169), .A2(n2170), .ZN(n2136) );
NAND2_X1 U1759 ( .A1(n2168), .A2(n2166), .ZN(n2170) );
NAND2_X1 U1760 ( .A1(KEYINPUT9), .A2(n2171), .ZN(n2166) );
NAND2_X1 U1761 ( .A1(n2172), .A2(n2173), .ZN(n2168) );
NAND2_X1 U1762 ( .A1(RESTART), .A2(n2174), .ZN(n2173) );
NAND2_X1 U1763 ( .A1(n2175), .A2(n2176), .ZN(n2174) );
NAND2_X1 U1764 ( .A1(KEYINPUT9), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2176) );
INV_X1 U1765 ( .A(RMIN_REG_0__SCAN_IN), .ZN(n2175) );
NAND2_X1 U1766 ( .A1(n2177), .A2(n1994), .ZN(n2172) );
NAND2_X1 U1767 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
NAND2_X1 U1768 ( .A1(KEYINPUT9), .A2(DATA_IN_0_), .ZN(n2179) );
INV_X1 U1769 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2178) );
NOR2_X1 U1770 ( .A1(n1932), .A2(n1953), .ZN(n2164) );
INV_X1 U1771 ( .A(n1961), .ZN(n1953) );
NAND3_X1 U1772 ( .A1(n2163), .A2(n2180), .A3(RESTART), .ZN(n1961) );
INV_X1 U1773 ( .A(n1943), .ZN(n1932) );
NAND3_X1 U1774 ( .A1(n2181), .A2(n2182), .A3(n2183), .ZN(n1943) );
XOR2_X1 U1775 ( .A(KEYINPUT33), .B(n2184), .Z(n2181) );
NOR2_X1 U1776 ( .A1(n2169), .A2(n1974), .ZN(n2160) );
NAND3_X1 U1777 ( .A1(n2185), .A2(n2186), .A3(n2163), .ZN(n1974) );
NAND2_X1 U1778 ( .A1(n2187), .A2(n1994), .ZN(n2186) );
NAND4_X1 U1779 ( .A1(n2184), .A2(ENABLE), .A3(n2188), .A4(n2182), .ZN(n2187));
INV_X1 U1780 ( .A(AVERAGE), .ZN(n2182) );
NAND2_X1 U1781 ( .A1(n2180), .A2(n2189), .ZN(n2188) );
INV_X1 U1782 ( .A(KEYINPUT25), .ZN(n2189) );
AND2_X1 U1783 ( .A1(n2190), .A2(n2191), .ZN(n2184) );
NAND2_X1 U1784 ( .A1(n2192), .A2(DATA_IN_7_), .ZN(n2191) );
XNOR2_X1 U1785 ( .A(REG4_REG_7__SCAN_IN), .B(KEYINPUT21), .ZN(n2192) );
XOR2_X1 U1786 ( .A(n2193), .B(KEYINPUT6), .Z(n2190) );
NAND3_X1 U1787 ( .A1(n2194), .A2(n2195), .A3(n2196), .ZN(n2193) );
OR2_X1 U1788 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2196) );
NAND3_X1 U1789 ( .A1(n2197), .A2(n2198), .A3(n2199), .ZN(n2195) );
NAND2_X1 U1790 ( .A1(n1768), .A2(n1993), .ZN(n2199) );
INV_X1 U1791 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1993) );
INV_X1 U1792 ( .A(DATA_IN_6_), .ZN(n1768) );
NAND3_X1 U1793 ( .A1(n2200), .A2(n2201), .A3(n2202), .ZN(n2198) );
NAND2_X1 U1794 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2202) );
NAND3_X1 U1795 ( .A1(n2203), .A2(n2204), .A3(n2205), .ZN(n2201) );
NAND2_X1 U1796 ( .A1(n1787), .A2(n2124), .ZN(n2205) );
INV_X1 U1797 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2124) );
INV_X1 U1798 ( .A(DATA_IN_3_), .ZN(n1787) );
NAND3_X1 U1799 ( .A1(n2206), .A2(n2207), .A3(n2208), .ZN(n2204) );
NAND2_X1 U1800 ( .A1(REG4_REG_3__SCAN_IN), .A2(DATA_IN_3_), .ZN(n2208) );
NAND3_X1 U1801 ( .A1(n2209), .A2(n2210), .A3(n2211), .ZN(n2207) );
NAND2_X1 U1802 ( .A1(n1782), .A2(n2144), .ZN(n2211) );
INV_X1 U1803 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2144) );
INV_X1 U1804 ( .A(DATA_IN_2_), .ZN(n1782) );
NAND2_X1 U1805 ( .A1(n2212), .A2(n2213), .ZN(n2210) );
OR2_X1 U1806 ( .A1(n2214), .A2(n1786), .ZN(n2212) );
NAND2_X1 U1807 ( .A1(n2214), .A2(n1786), .ZN(n2209) );
NAND2_X1 U1808 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2206) );
NAND2_X1 U1809 ( .A1(n2215), .A2(n1721), .ZN(n2203) );
INV_X1 U1810 ( .A(DATA_IN_4_), .ZN(n1721) );
XOR2_X1 U1811 ( .A(REG4_REG_4__SCAN_IN), .B(KEYINPUT1), .Z(n2215) );
NAND2_X1 U1812 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2200) );
NAND2_X1 U1813 ( .A1(n1804), .A2(n2031), .ZN(n2197) );
INV_X1 U1814 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2031) );
INV_X1 U1815 ( .A(DATA_IN_5_), .ZN(n1804) );
NAND2_X1 U1816 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2194) );
NAND3_X1 U1817 ( .A1(KEYINPUT25), .A2(n2180), .A3(RESTART), .ZN(n2185) );
XNOR2_X1 U1818 ( .A(n2216), .B(KEYINPUT14), .ZN(n2180) );
NAND2_X1 U1819 ( .A1(n2217), .A2(n2218), .ZN(n2216) );
NAND2_X1 U1820 ( .A1(n2219), .A2(n1764), .ZN(n2218) );
INV_X1 U1821 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1764) );
OR2_X1 U1822 ( .A1(n2220), .A2(n1796), .ZN(n2219) );
NAND2_X1 U1823 ( .A1(n2220), .A2(n1796), .ZN(n2217) );
INV_X1 U1824 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1796) );
NAND2_X1 U1825 ( .A1(n2221), .A2(n2222), .ZN(n2220) );
NAND2_X1 U1826 ( .A1(n2223), .A2(n2224), .ZN(n2222) );
NAND2_X1 U1827 ( .A1(n1791), .A2(n1800), .ZN(n2224) );
INV_X1 U1828 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1800) );
INV_X1 U1829 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1791) );
NAND2_X1 U1830 ( .A1(n2225), .A2(n2226), .ZN(n2223) );
NAND2_X1 U1831 ( .A1(RMIN_REG_5__SCAN_IN), .A2(RMAX_REG_5__SCAN_IN), .ZN(n2226) );
NAND2_X1 U1832 ( .A1(n2227), .A2(n2228), .ZN(n2225) );
NAND2_X1 U1833 ( .A1(n2229), .A2(n2230), .ZN(n2228) );
NAND3_X1 U1834 ( .A1(n2231), .A2(n2232), .A3(n2233), .ZN(n2230) );
NAND2_X1 U1835 ( .A1(n1808), .A2(n1788), .ZN(n2233) );
INV_X1 U1836 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1788) );
INV_X1 U1837 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1808) );
NAND3_X1 U1838 ( .A1(n2234), .A2(n2235), .A3(n2236), .ZN(n2232) );
NAND2_X1 U1839 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2236) );
NAND3_X1 U1840 ( .A1(n2237), .A2(n2238), .A3(n2239), .ZN(n2235) );
NAND2_X1 U1841 ( .A1(n1819), .A2(n1785), .ZN(n2239) );
NAND2_X1 U1842 ( .A1(n2240), .A2(n2241), .ZN(n2238) );
NAND2_X1 U1843 ( .A1(RMIN_REG_1__SCAN_IN), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2241) );
XOR2_X1 U1844 ( .A(n2242), .B(KEYINPUT58), .Z(n2240) );
NAND2_X1 U1845 ( .A1(n2243), .A2(n1816), .ZN(n2237) );
INV_X1 U1846 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1816) );
XOR2_X1 U1847 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT24), .Z(n2243) );
NAND2_X1 U1848 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2234) );
NAND2_X1 U1849 ( .A1(n1821), .A2(n1747), .ZN(n2231) );
INV_X1 U1850 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1747) );
INV_X1 U1851 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1821) );
XOR2_X1 U1852 ( .A(n2244), .B(KEYINPUT3), .Z(n2229) );
NAND2_X1 U1853 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2244) );
NAND2_X1 U1854 ( .A1(n2245), .A2(n1772), .ZN(n2227) );
INV_X1 U1855 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1772) );
XOR2_X1 U1856 ( .A(n1822), .B(KEYINPUT59), .Z(n2245) );
INV_X1 U1857 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1822) );
NAND2_X1 U1858 ( .A1(RMIN_REG_6__SCAN_IN), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2221) );
INV_X1 U1859 ( .A(n2167), .ZN(n2169) );
NAND3_X1 U1860 ( .A1(n2246), .A2(n2247), .A3(n2248), .ZN(n2167) );
NAND2_X1 U1861 ( .A1(n2153), .A2(n2249), .ZN(n2248) );
NAND2_X1 U1862 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
NAND2_X1 U1863 ( .A1(n2154), .A2(n2252), .ZN(n2251) );
INV_X1 U1864 ( .A(KEYINPUT22), .ZN(n2252) );
XOR2_X1 U1865 ( .A(n2253), .B(n2254), .Z(n2250) );
NOR2_X1 U1866 ( .A1(KEYINPUT41), .A2(n2154), .ZN(n2254) );
NAND2_X1 U1867 ( .A1(n2253), .A2(n2255), .ZN(n2247) );
NAND2_X1 U1868 ( .A1(n2256), .A2(n2257), .ZN(n2255) );
NAND3_X1 U1869 ( .A1(n2171), .A2(n2154), .A3(KEYINPUT22), .ZN(n2257) );
NAND2_X1 U1870 ( .A1(KEYINPUT12), .A2(n2152), .ZN(n2256) );
NAND3_X1 U1871 ( .A1(n2152), .A2(n2258), .A3(n2151), .ZN(n2246) );
INV_X1 U1872 ( .A(n2253), .ZN(n2151) );
NAND2_X1 U1873 ( .A1(n2259), .A2(n2260), .ZN(n2253) );
NAND2_X1 U1874 ( .A1(RESTART), .A2(n1785), .ZN(n2260) );
INV_X1 U1875 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1785) );
NAND2_X1 U1876 ( .A1(n2213), .A2(n1994), .ZN(n2259) );
INV_X1 U1877 ( .A(REG4_REG_1__SCAN_IN), .ZN(n2213) );
INV_X1 U1878 ( .A(KEYINPUT12), .ZN(n2258) );
NOR2_X1 U1879 ( .A1(n2154), .A2(n2261), .ZN(n2152) );
XOR2_X1 U1880 ( .A(n2171), .B(KEYINPUT22), .Z(n2261) );
INV_X1 U1881 ( .A(n2153), .ZN(n2171) );
NAND2_X1 U1882 ( .A1(n2262), .A2(n2263), .ZN(n2153) );
NAND2_X1 U1883 ( .A1(n2214), .A2(n1994), .ZN(n2263) );
NAND2_X1 U1884 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2214) );
NAND2_X1 U1885 ( .A1(RESTART), .A2(n2242), .ZN(n2262) );
NAND2_X1 U1886 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2242) );
NAND2_X1 U1887 ( .A1(n2264), .A2(n2265), .ZN(n2154) );
NAND2_X1 U1888 ( .A1(RESTART), .A2(n1819), .ZN(n2265) );
INV_X1 U1889 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1819) );
NAND2_X1 U1890 ( .A1(n2266), .A2(n1994), .ZN(n2264) );
XOR2_X1 U1891 ( .A(n1786), .B(KEYINPUT7), .Z(n2266) );
INV_X1 U1892 ( .A(DATA_IN_1_), .ZN(n1786) );
NAND2_X1 U1893 ( .A1(n1935), .A2(REG4_REG_0__SCAN_IN), .ZN(n2158) );
INV_X1 U1894 ( .A(n2108), .ZN(n1935) );
NAND2_X1 U1895 ( .A1(AVERAGE), .A2(n2183), .ZN(n2108) );
AND3_X1 U1896 ( .A1(n2163), .A2(n1994), .A3(ENABLE), .ZN(n2183) );
INV_X1 U1897 ( .A(RESTART), .ZN(n1994) );
NOR2_X1 U1898 ( .A1(n1845), .A2(n1849), .ZN(n2163) );
NAND2_X1 U1899 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1849), .ZN(n2157) );
NAND2_X1 U1900 ( .A1(n1862), .A2(n2267), .ZN(U280) );
NAND2_X1 U1901 ( .A1(STATO_REG_0__SCAN_IN), .A2(n1845), .ZN(n2267) );
INV_X1 U1902 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1845) );
NAND2_X1 U1903 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1732), .ZN(n1862) );
INV_X1 U1904 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1732) );
endmodule


