//Key = 1000100000100101100100000111011100111001010010101000001101000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;

XNOR2_X1 U743 ( .A(n1027), .B(n1028), .ZN(G9) );
XNOR2_X1 U744 ( .A(G107), .B(KEYINPUT18), .ZN(n1028) );
NOR2_X1 U745 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U746 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
XOR2_X1 U747 ( .A(n1035), .B(KEYINPUT12), .Z(n1034) );
NAND2_X1 U748 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U749 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND2_X1 U750 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND2_X1 U751 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1036) );
AND2_X1 U757 ( .A1(n1055), .A2(n1053), .ZN(n1033) );
AND3_X1 U758 ( .A1(n1051), .A2(n1043), .A3(n1040), .ZN(n1053) );
NAND3_X1 U759 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1031) );
NAND3_X1 U760 ( .A1(n1038), .A2(n1059), .A3(n1040), .ZN(n1058) );
INV_X1 U761 ( .A(n1060), .ZN(n1040) );
NAND2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND4_X1 U763 ( .A1(n1051), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1062) );
INV_X1 U764 ( .A(KEYINPUT47), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1043), .A2(n1066), .ZN(n1061) );
NAND3_X1 U766 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
NAND2_X1 U767 ( .A1(KEYINPUT47), .A2(n1051), .ZN(n1069) );
AND2_X1 U768 ( .A1(n1048), .A2(n1049), .ZN(n1051) );
NAND3_X1 U769 ( .A1(n1070), .A2(n1071), .A3(n1048), .ZN(n1068) );
NAND3_X1 U770 ( .A1(n1072), .A2(n1049), .A3(n1073), .ZN(n1067) );
AND3_X1 U771 ( .A1(n1056), .A2(n1057), .A3(n1074), .ZN(n1029) );
NAND4_X1 U772 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1056) );
NOR4_X1 U773 ( .A1(n1079), .A2(n1063), .A3(n1080), .A4(n1081), .ZN(n1078) );
XOR2_X1 U774 ( .A(n1082), .B(n1083), .Z(n1081) );
NAND2_X1 U775 ( .A1(KEYINPUT48), .A2(n1084), .ZN(n1082) );
NOR2_X1 U776 ( .A1(n1085), .A2(n1086), .ZN(n1080) );
INV_X1 U777 ( .A(n1087), .ZN(n1063) );
INV_X1 U778 ( .A(n1088), .ZN(n1079) );
NOR2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1077) );
XOR2_X1 U780 ( .A(n1091), .B(n1092), .Z(n1089) );
NAND2_X1 U781 ( .A1(KEYINPUT25), .A2(n1093), .ZN(n1091) );
XOR2_X1 U782 ( .A(n1094), .B(n1095), .Z(n1076) );
XNOR2_X1 U783 ( .A(n1096), .B(KEYINPUT41), .ZN(n1094) );
XOR2_X1 U784 ( .A(n1097), .B(KEYINPUT28), .Z(n1075) );
XOR2_X1 U785 ( .A(n1098), .B(n1099), .Z(G72) );
NOR2_X1 U786 ( .A1(n1057), .A2(n1100), .ZN(n1099) );
XOR2_X1 U787 ( .A(KEYINPUT23), .B(n1101), .Z(n1100) );
AND2_X1 U788 ( .A1(G227), .A2(G900), .ZN(n1101) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
NAND3_X1 U790 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1103) );
INV_X1 U791 ( .A(n1107), .ZN(n1105) );
OR2_X1 U792 ( .A1(n1106), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U793 ( .A(n1108), .B(n1109), .ZN(n1104) );
XNOR2_X1 U794 ( .A(n1110), .B(n1111), .ZN(n1108) );
NOR3_X1 U795 ( .A1(KEYINPUT20), .A2(n1112), .A3(n1113), .ZN(n1111) );
NOR3_X1 U796 ( .A1(G131), .A2(n1114), .A3(n1115), .ZN(n1113) );
NOR2_X1 U797 ( .A1(n1116), .A2(n1117), .ZN(n1112) );
NOR2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(n1116) );
NAND2_X1 U799 ( .A1(n1057), .A2(n1118), .ZN(n1106) );
NAND4_X1 U800 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U802 ( .A1(n1125), .A2(n1126), .ZN(G69) );
NAND2_X1 U803 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND3_X1 U804 ( .A1(n1129), .A2(n1130), .A3(G953), .ZN(n1128) );
NAND2_X1 U805 ( .A1(G898), .A2(G224), .ZN(n1129) );
NAND3_X1 U806 ( .A1(n1131), .A2(n1130), .A3(n1132), .ZN(n1125) );
INV_X1 U807 ( .A(n1127), .ZN(n1132) );
XNOR2_X1 U808 ( .A(n1133), .B(n1134), .ZN(n1127) );
NOR2_X1 U809 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XNOR2_X1 U810 ( .A(KEYINPUT58), .B(n1057), .ZN(n1136) );
NAND2_X1 U811 ( .A1(n1137), .A2(n1138), .ZN(n1133) );
XNOR2_X1 U812 ( .A(KEYINPUT60), .B(n1139), .ZN(n1137) );
INV_X1 U813 ( .A(n1140), .ZN(n1139) );
INV_X1 U814 ( .A(KEYINPUT9), .ZN(n1130) );
NAND2_X1 U815 ( .A1(n1138), .A2(n1141), .ZN(n1131) );
OR2_X1 U816 ( .A1(n1057), .A2(G224), .ZN(n1141) );
INV_X1 U817 ( .A(n1142), .ZN(n1138) );
NOR3_X1 U818 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(G66) );
NOR3_X1 U819 ( .A1(n1146), .A2(n1057), .A3(n1074), .ZN(n1145) );
INV_X1 U820 ( .A(G952), .ZN(n1074) );
AND2_X1 U821 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
INV_X1 U822 ( .A(KEYINPUT2), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1148), .B(n1149), .Z(n1143) );
NOR2_X1 U824 ( .A1(n1150), .A2(KEYINPUT24), .ZN(n1149) );
OR2_X1 U825 ( .A1(n1151), .A2(n1086), .ZN(n1148) );
NOR2_X1 U826 ( .A1(n1147), .A2(n1152), .ZN(G63) );
NOR3_X1 U827 ( .A1(n1092), .A2(n1153), .A3(n1154), .ZN(n1152) );
NOR3_X1 U828 ( .A1(n1155), .A2(n1093), .A3(n1151), .ZN(n1154) );
NOR2_X1 U829 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
NOR2_X1 U830 ( .A1(n1158), .A2(n1093), .ZN(n1156) );
NOR2_X1 U831 ( .A1(n1147), .A2(n1159), .ZN(G60) );
NOR3_X1 U832 ( .A1(n1096), .A2(n1160), .A3(n1161), .ZN(n1159) );
NOR3_X1 U833 ( .A1(n1162), .A2(n1163), .A3(n1151), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
NOR2_X1 U835 ( .A1(n1158), .A2(n1163), .ZN(n1164) );
INV_X1 U836 ( .A(n1032), .ZN(n1158) );
XNOR2_X1 U837 ( .A(G104), .B(n1166), .ZN(G6) );
NOR2_X1 U838 ( .A1(n1147), .A2(n1167), .ZN(G57) );
XOR2_X1 U839 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U840 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U841 ( .A(n1172), .B(n1173), .Z(n1168) );
XOR2_X1 U842 ( .A(KEYINPUT61), .B(n1174), .Z(n1173) );
NOR2_X1 U843 ( .A1(n1084), .A2(n1151), .ZN(n1174) );
INV_X1 U844 ( .A(G472), .ZN(n1084) );
NOR2_X1 U845 ( .A1(n1147), .A2(n1175), .ZN(G54) );
XOR2_X1 U846 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U847 ( .A(n1178), .B(n1179), .ZN(n1177) );
NAND3_X1 U848 ( .A1(n1180), .A2(n1181), .A3(KEYINPUT16), .ZN(n1178) );
NAND2_X1 U849 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XOR2_X1 U850 ( .A(KEYINPUT30), .B(n1184), .Z(n1180) );
NOR2_X1 U851 ( .A1(n1182), .A2(n1183), .ZN(n1184) );
XNOR2_X1 U852 ( .A(n1185), .B(n1186), .ZN(n1183) );
NOR2_X1 U853 ( .A1(KEYINPUT37), .A2(n1187), .ZN(n1186) );
XNOR2_X1 U854 ( .A(n1188), .B(KEYINPUT42), .ZN(n1182) );
XOR2_X1 U855 ( .A(n1189), .B(n1190), .Z(n1176) );
NOR2_X1 U856 ( .A1(KEYINPUT52), .A2(n1191), .ZN(n1190) );
NOR2_X1 U857 ( .A1(n1192), .A2(n1151), .ZN(n1189) );
NOR2_X1 U858 ( .A1(n1147), .A2(n1193), .ZN(G51) );
XNOR2_X1 U859 ( .A(n1140), .B(n1194), .ZN(n1193) );
XOR2_X1 U860 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U861 ( .A1(n1197), .A2(n1151), .ZN(n1196) );
NAND2_X1 U862 ( .A1(G902), .A2(n1032), .ZN(n1151) );
NAND4_X1 U863 ( .A1(n1198), .A2(n1199), .A3(n1135), .A4(n1200), .ZN(n1032) );
NOR3_X1 U864 ( .A1(n1123), .A2(n1201), .A3(n1202), .ZN(n1200) );
AND3_X1 U865 ( .A1(n1203), .A2(n1055), .A3(n1204), .ZN(n1123) );
XNOR2_X1 U866 ( .A(n1050), .B(KEYINPUT10), .ZN(n1204) );
AND4_X1 U867 ( .A1(n1166), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1135) );
NOR4_X1 U868 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1027), .ZN(n1207) );
AND4_X1 U869 ( .A1(n1052), .A2(n1211), .A3(n1049), .A4(n1055), .ZN(n1027) );
NAND3_X1 U870 ( .A1(n1211), .A2(n1212), .A3(n1043), .ZN(n1206) );
NAND2_X1 U871 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U872 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XNOR2_X1 U873 ( .A(n1049), .B(KEYINPUT57), .ZN(n1215) );
NAND2_X1 U874 ( .A1(n1047), .A2(n1054), .ZN(n1213) );
NAND4_X1 U875 ( .A1(n1052), .A2(n1211), .A3(n1049), .A4(n1054), .ZN(n1166) );
XNOR2_X1 U876 ( .A(KEYINPUT0), .B(n1119), .ZN(n1199) );
XNOR2_X1 U877 ( .A(KEYINPUT59), .B(n1124), .ZN(n1198) );
NAND4_X1 U878 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1124) );
NAND3_X1 U879 ( .A1(n1216), .A2(n1221), .A3(n1222), .ZN(n1217) );
XOR2_X1 U880 ( .A(KEYINPUT38), .B(n1050), .Z(n1221) );
NOR3_X1 U881 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1195) );
NOR2_X1 U882 ( .A1(KEYINPUT17), .A2(n1226), .ZN(n1225) );
NOR2_X1 U883 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
AND3_X1 U884 ( .A1(KEYINPUT27), .A2(n1229), .A3(n1230), .ZN(n1228) );
NOR2_X1 U885 ( .A1(KEYINPUT27), .A2(n1229), .ZN(n1227) );
NOR2_X1 U886 ( .A1(n1231), .A2(n1232), .ZN(n1224) );
INV_X1 U887 ( .A(KEYINPUT17), .ZN(n1232) );
NOR2_X1 U888 ( .A1(n1233), .A2(n1234), .ZN(n1231) );
XOR2_X1 U889 ( .A(KEYINPUT27), .B(n1229), .Z(n1234) );
NOR2_X1 U890 ( .A1(n1230), .A2(n1229), .ZN(n1223) );
XOR2_X1 U891 ( .A(G125), .B(n1171), .Z(n1229) );
NOR2_X1 U892 ( .A1(n1057), .A2(G952), .ZN(n1147) );
XNOR2_X1 U893 ( .A(G146), .B(n1218), .ZN(G48) );
NAND2_X1 U894 ( .A1(n1235), .A2(n1054), .ZN(n1218) );
XOR2_X1 U895 ( .A(n1236), .B(n1237), .Z(G45) );
XOR2_X1 U896 ( .A(KEYINPUT15), .B(G143), .Z(n1237) );
NAND3_X1 U897 ( .A1(n1216), .A2(n1050), .A3(n1222), .ZN(n1236) );
XNOR2_X1 U898 ( .A(G140), .B(n1219), .ZN(G42) );
NAND3_X1 U899 ( .A1(n1048), .A2(n1052), .A3(n1238), .ZN(n1219) );
XNOR2_X1 U900 ( .A(G137), .B(n1220), .ZN(G39) );
NAND3_X1 U901 ( .A1(n1203), .A2(n1048), .A3(n1038), .ZN(n1220) );
XNOR2_X1 U902 ( .A(G134), .B(n1239), .ZN(G36) );
NAND2_X1 U903 ( .A1(KEYINPUT62), .A2(n1202), .ZN(n1239) );
INV_X1 U904 ( .A(n1121), .ZN(n1202) );
NAND3_X1 U905 ( .A1(n1048), .A2(n1055), .A3(n1222), .ZN(n1121) );
XNOR2_X1 U906 ( .A(G131), .B(n1119), .ZN(G33) );
NAND3_X1 U907 ( .A1(n1048), .A2(n1054), .A3(n1222), .ZN(n1119) );
AND3_X1 U908 ( .A1(n1052), .A2(n1240), .A3(n1047), .ZN(n1222) );
INV_X1 U909 ( .A(n1090), .ZN(n1048) );
NAND2_X1 U910 ( .A1(n1072), .A2(n1241), .ZN(n1090) );
XNOR2_X1 U911 ( .A(G128), .B(n1242), .ZN(G30) );
NAND2_X1 U912 ( .A1(n1235), .A2(n1055), .ZN(n1242) );
AND2_X1 U913 ( .A1(n1203), .A2(n1050), .ZN(n1235) );
AND4_X1 U914 ( .A1(n1243), .A2(n1052), .A3(n1240), .A4(n1071), .ZN(n1203) );
XNOR2_X1 U915 ( .A(G101), .B(n1205), .ZN(G3) );
NAND3_X1 U916 ( .A1(n1038), .A2(n1052), .A3(n1244), .ZN(n1205) );
NAND2_X1 U917 ( .A1(n1245), .A2(n1246), .ZN(G27) );
NAND2_X1 U918 ( .A1(n1201), .A2(n1247), .ZN(n1246) );
XOR2_X1 U919 ( .A(KEYINPUT36), .B(n1248), .Z(n1245) );
NOR2_X1 U920 ( .A1(n1201), .A2(n1247), .ZN(n1248) );
INV_X1 U921 ( .A(G125), .ZN(n1247) );
INV_X1 U922 ( .A(n1120), .ZN(n1201) );
NAND3_X1 U923 ( .A1(n1238), .A2(n1050), .A3(n1043), .ZN(n1120) );
AND4_X1 U924 ( .A1(n1054), .A2(n1070), .A3(n1240), .A4(n1071), .ZN(n1238) );
NAND2_X1 U925 ( .A1(n1060), .A2(n1249), .ZN(n1240) );
NAND3_X1 U926 ( .A1(n1250), .A2(n1251), .A3(n1107), .ZN(n1249) );
NOR2_X1 U927 ( .A1(n1057), .A2(G900), .ZN(n1107) );
XNOR2_X1 U928 ( .A(KEYINPUT63), .B(n1252), .ZN(n1250) );
XOR2_X1 U929 ( .A(n1253), .B(G122), .Z(G24) );
NAND2_X1 U930 ( .A1(KEYINPUT54), .A2(n1254), .ZN(n1253) );
NAND4_X1 U931 ( .A1(n1043), .A2(n1211), .A3(n1049), .A4(n1216), .ZN(n1254) );
NOR2_X1 U932 ( .A1(n1071), .A2(n1243), .ZN(n1049) );
XOR2_X1 U933 ( .A(G119), .B(n1210), .Z(G21) );
AND3_X1 U934 ( .A1(n1243), .A2(n1043), .A3(n1255), .ZN(n1210) );
INV_X1 U935 ( .A(n1070), .ZN(n1243) );
XNOR2_X1 U936 ( .A(n1256), .B(n1209), .ZN(G18) );
AND3_X1 U937 ( .A1(n1043), .A2(n1055), .A3(n1244), .ZN(n1209) );
NAND2_X1 U938 ( .A1(n1257), .A2(n1258), .ZN(n1055) );
OR3_X1 U939 ( .A1(n1259), .A2(n1260), .A3(KEYINPUT49), .ZN(n1258) );
NAND2_X1 U940 ( .A1(KEYINPUT49), .A2(n1216), .ZN(n1257) );
XNOR2_X1 U941 ( .A(G113), .B(n1261), .ZN(G15) );
NAND3_X1 U942 ( .A1(n1244), .A2(n1054), .A3(n1262), .ZN(n1261) );
XNOR2_X1 U943 ( .A(n1043), .B(KEYINPUT35), .ZN(n1262) );
AND2_X1 U944 ( .A1(n1064), .A2(n1087), .ZN(n1043) );
XOR2_X1 U945 ( .A(n1263), .B(KEYINPUT6), .Z(n1064) );
NAND2_X1 U946 ( .A1(n1264), .A2(n1265), .ZN(n1054) );
NAND2_X1 U947 ( .A1(n1216), .A2(n1266), .ZN(n1265) );
INV_X1 U948 ( .A(KEYINPUT13), .ZN(n1266) );
AND2_X1 U949 ( .A1(n1267), .A2(n1260), .ZN(n1216) );
NAND3_X1 U950 ( .A1(n1260), .A2(n1259), .A3(KEYINPUT13), .ZN(n1264) );
AND2_X1 U951 ( .A1(n1047), .A2(n1211), .ZN(n1244) );
NOR2_X1 U952 ( .A1(n1070), .A2(n1071), .ZN(n1047) );
XNOR2_X1 U953 ( .A(n1185), .B(n1208), .ZN(G12) );
AND3_X1 U954 ( .A1(n1052), .A2(n1070), .A3(n1255), .ZN(n1208) );
AND3_X1 U955 ( .A1(n1211), .A2(n1071), .A3(n1038), .ZN(n1255) );
NOR2_X1 U956 ( .A1(n1267), .A2(n1260), .ZN(n1038) );
XOR2_X1 U957 ( .A(n1096), .B(n1268), .Z(n1260) );
NOR2_X1 U958 ( .A1(KEYINPUT43), .A2(n1095), .ZN(n1268) );
XNOR2_X1 U959 ( .A(n1163), .B(KEYINPUT4), .ZN(n1095) );
INV_X1 U960 ( .A(G475), .ZN(n1163) );
NOR2_X1 U961 ( .A1(n1165), .A2(G902), .ZN(n1096) );
INV_X1 U962 ( .A(n1162), .ZN(n1165) );
XNOR2_X1 U963 ( .A(n1269), .B(n1270), .ZN(n1162) );
XNOR2_X1 U964 ( .A(n1271), .B(n1272), .ZN(n1270) );
NOR2_X1 U965 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U966 ( .A(n1275), .B(KEYINPUT34), .Z(n1274) );
NAND2_X1 U967 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NOR2_X1 U968 ( .A1(n1277), .A2(n1276), .ZN(n1273) );
XNOR2_X1 U969 ( .A(n1278), .B(KEYINPUT32), .ZN(n1276) );
XOR2_X1 U970 ( .A(n1279), .B(n1280), .Z(n1277) );
XNOR2_X1 U971 ( .A(G143), .B(n1117), .ZN(n1280) );
NAND2_X1 U972 ( .A1(n1281), .A2(G214), .ZN(n1279) );
INV_X1 U973 ( .A(G104), .ZN(n1271) );
XNOR2_X1 U974 ( .A(G113), .B(G122), .ZN(n1269) );
INV_X1 U975 ( .A(n1259), .ZN(n1267) );
XOR2_X1 U976 ( .A(n1092), .B(n1093), .Z(n1259) );
INV_X1 U977 ( .A(G478), .ZN(n1093) );
NOR2_X1 U978 ( .A1(n1157), .A2(G902), .ZN(n1092) );
INV_X1 U979 ( .A(n1155), .ZN(n1157) );
XOR2_X1 U980 ( .A(n1282), .B(n1283), .Z(n1155) );
XNOR2_X1 U981 ( .A(n1284), .B(n1285), .ZN(n1283) );
NAND2_X1 U982 ( .A1(n1286), .A2(n1287), .ZN(n1284) );
NAND2_X1 U983 ( .A1(G107), .A2(n1288), .ZN(n1287) );
XOR2_X1 U984 ( .A(n1289), .B(KEYINPUT51), .Z(n1286) );
OR2_X1 U985 ( .A1(n1288), .A2(G107), .ZN(n1289) );
XOR2_X1 U986 ( .A(G116), .B(G122), .Z(n1288) );
XOR2_X1 U987 ( .A(n1290), .B(n1291), .Z(n1282) );
XNOR2_X1 U988 ( .A(G143), .B(n1292), .ZN(n1291) );
NAND3_X1 U989 ( .A1(G234), .A2(n1057), .A3(G217), .ZN(n1290) );
NAND3_X1 U990 ( .A1(n1293), .A2(n1294), .A3(n1088), .ZN(n1071) );
NAND2_X1 U991 ( .A1(n1085), .A2(n1086), .ZN(n1088) );
NAND2_X1 U992 ( .A1(KEYINPUT11), .A2(n1086), .ZN(n1294) );
OR3_X1 U993 ( .A1(n1085), .A2(KEYINPUT11), .A3(n1086), .ZN(n1293) );
NAND2_X1 U994 ( .A1(G217), .A2(n1295), .ZN(n1086) );
NOR2_X1 U995 ( .A1(G902), .A2(n1150), .ZN(n1085) );
AND3_X1 U996 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1150) );
NAND2_X1 U997 ( .A1(KEYINPUT53), .A2(n1299), .ZN(n1298) );
OR3_X1 U998 ( .A1(n1299), .A2(KEYINPUT53), .A3(n1300), .ZN(n1297) );
NAND2_X1 U999 ( .A1(n1300), .A2(n1301), .ZN(n1296) );
NAND2_X1 U1000 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
INV_X1 U1001 ( .A(KEYINPUT53), .ZN(n1303) );
XNOR2_X1 U1002 ( .A(n1299), .B(KEYINPUT40), .ZN(n1302) );
XNOR2_X1 U1003 ( .A(n1304), .B(n1305), .ZN(n1299) );
NOR2_X1 U1004 ( .A1(KEYINPUT7), .A2(n1306), .ZN(n1305) );
NAND3_X1 U1005 ( .A1(n1307), .A2(n1057), .A3(G221), .ZN(n1304) );
XOR2_X1 U1006 ( .A(KEYINPUT21), .B(G234), .Z(n1307) );
XOR2_X1 U1007 ( .A(n1308), .B(n1278), .Z(n1300) );
XOR2_X1 U1008 ( .A(G146), .B(n1110), .Z(n1278) );
XOR2_X1 U1009 ( .A(G125), .B(G140), .Z(n1110) );
XNOR2_X1 U1010 ( .A(G110), .B(n1309), .ZN(n1308) );
NOR2_X1 U1011 ( .A1(KEYINPUT22), .A2(n1310), .ZN(n1309) );
NOR2_X1 U1012 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1013 ( .A(n1313), .B(KEYINPUT19), .Z(n1312) );
NAND2_X1 U1014 ( .A1(G119), .A2(n1285), .ZN(n1313) );
NOR2_X1 U1015 ( .A1(G119), .A2(n1285), .ZN(n1311) );
AND2_X1 U1016 ( .A1(n1050), .A2(n1314), .ZN(n1211) );
NAND2_X1 U1017 ( .A1(n1060), .A2(n1315), .ZN(n1314) );
NAND3_X1 U1018 ( .A1(n1142), .A2(n1251), .A3(G902), .ZN(n1315) );
NOR2_X1 U1019 ( .A1(n1057), .A2(G898), .ZN(n1142) );
NAND3_X1 U1020 ( .A1(n1251), .A2(n1057), .A3(G952), .ZN(n1060) );
NAND2_X1 U1021 ( .A1(G237), .A2(G234), .ZN(n1251) );
NOR2_X1 U1022 ( .A1(n1072), .A2(n1073), .ZN(n1050) );
INV_X1 U1023 ( .A(n1241), .ZN(n1073) );
NAND2_X1 U1024 ( .A1(G214), .A2(n1316), .ZN(n1241) );
XNOR2_X1 U1025 ( .A(n1317), .B(n1197), .ZN(n1072) );
NAND2_X1 U1026 ( .A1(G210), .A2(n1316), .ZN(n1197) );
NAND2_X1 U1027 ( .A1(n1318), .A2(n1252), .ZN(n1316) );
INV_X1 U1028 ( .A(G237), .ZN(n1318) );
NAND2_X1 U1029 ( .A1(n1319), .A2(n1252), .ZN(n1317) );
XOR2_X1 U1030 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1031 ( .A(n1322), .B(n1171), .Z(n1321) );
NOR2_X1 U1032 ( .A1(G125), .A2(KEYINPUT56), .ZN(n1322) );
XOR2_X1 U1033 ( .A(n1323), .B(n1324), .Z(n1320) );
NOR2_X1 U1034 ( .A1(KEYINPUT45), .A2(n1140), .ZN(n1324) );
XNOR2_X1 U1035 ( .A(n1325), .B(n1326), .ZN(n1140) );
XOR2_X1 U1036 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1037 ( .A1(G104), .A2(KEYINPUT14), .ZN(n1327) );
XNOR2_X1 U1038 ( .A(G107), .B(n1329), .ZN(n1325) );
XNOR2_X1 U1039 ( .A(G122), .B(n1185), .ZN(n1329) );
XNOR2_X1 U1040 ( .A(n1230), .B(KEYINPUT26), .ZN(n1323) );
INV_X1 U1041 ( .A(n1233), .ZN(n1230) );
NAND2_X1 U1042 ( .A1(G224), .A2(n1057), .ZN(n1233) );
XOR2_X1 U1043 ( .A(G472), .B(n1330), .Z(n1070) );
NOR2_X1 U1044 ( .A1(n1083), .A2(KEYINPUT5), .ZN(n1330) );
AND2_X1 U1045 ( .A1(n1331), .A2(n1252), .ZN(n1083) );
XNOR2_X1 U1046 ( .A(n1332), .B(n1172), .ZN(n1331) );
XNOR2_X1 U1047 ( .A(n1333), .B(n1328), .ZN(n1172) );
XNOR2_X1 U1048 ( .A(n1334), .B(n1335), .ZN(n1328) );
XNOR2_X1 U1049 ( .A(G119), .B(n1256), .ZN(n1335) );
INV_X1 U1050 ( .A(G116), .ZN(n1256) );
XNOR2_X1 U1051 ( .A(G101), .B(G113), .ZN(n1334) );
NAND2_X1 U1052 ( .A1(n1281), .A2(G210), .ZN(n1333) );
NOR2_X1 U1053 ( .A1(G953), .A2(G237), .ZN(n1281) );
NAND2_X1 U1054 ( .A1(KEYINPUT31), .A2(n1336), .ZN(n1332) );
XNOR2_X1 U1055 ( .A(n1337), .B(n1170), .ZN(n1336) );
NAND2_X1 U1056 ( .A1(KEYINPUT39), .A2(n1171), .ZN(n1337) );
XOR2_X1 U1057 ( .A(n1338), .B(n1339), .Z(n1171) );
AND2_X1 U1058 ( .A1(n1340), .A2(n1087), .ZN(n1052) );
NAND2_X1 U1059 ( .A1(G221), .A2(n1295), .ZN(n1087) );
NAND2_X1 U1060 ( .A1(G234), .A2(n1252), .ZN(n1295) );
XOR2_X1 U1061 ( .A(n1263), .B(KEYINPUT46), .Z(n1340) );
XOR2_X1 U1062 ( .A(n1097), .B(KEYINPUT8), .Z(n1263) );
XNOR2_X1 U1063 ( .A(n1341), .B(n1192), .ZN(n1097) );
INV_X1 U1064 ( .A(G469), .ZN(n1192) );
NAND2_X1 U1065 ( .A1(n1342), .A2(n1252), .ZN(n1341) );
INV_X1 U1066 ( .A(G902), .ZN(n1252) );
XOR2_X1 U1067 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1068 ( .A(n1345), .B(n1191), .ZN(n1344) );
XNOR2_X1 U1069 ( .A(n1346), .B(n1347), .ZN(n1191) );
NOR2_X1 U1070 ( .A1(KEYINPUT33), .A2(G101), .ZN(n1347) );
XNOR2_X1 U1071 ( .A(G104), .B(G107), .ZN(n1346) );
INV_X1 U1072 ( .A(n1179), .ZN(n1345) );
XOR2_X1 U1073 ( .A(n1170), .B(n1109), .Z(n1179) );
XNOR2_X1 U1074 ( .A(n1348), .B(n1339), .ZN(n1109) );
XOR2_X1 U1075 ( .A(G146), .B(n1285), .Z(n1339) );
XOR2_X1 U1076 ( .A(G128), .B(KEYINPUT55), .Z(n1285) );
XNOR2_X1 U1077 ( .A(KEYINPUT29), .B(n1349), .ZN(n1348) );
NOR2_X1 U1078 ( .A1(KEYINPUT3), .A2(n1338), .ZN(n1349) );
XOR2_X1 U1079 ( .A(G143), .B(KEYINPUT50), .Z(n1338) );
XOR2_X1 U1080 ( .A(n1350), .B(n1117), .Z(n1170) );
INV_X1 U1081 ( .A(G131), .ZN(n1117) );
NAND3_X1 U1082 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1350) );
INV_X1 U1083 ( .A(n1115), .ZN(n1353) );
NOR2_X1 U1084 ( .A1(n1306), .A2(G134), .ZN(n1115) );
INV_X1 U1085 ( .A(G137), .ZN(n1306) );
OR2_X1 U1086 ( .A1(G134), .A2(KEYINPUT44), .ZN(n1352) );
NAND2_X1 U1087 ( .A1(n1114), .A2(KEYINPUT44), .ZN(n1351) );
NOR2_X1 U1088 ( .A1(n1292), .A2(G137), .ZN(n1114) );
INV_X1 U1089 ( .A(G134), .ZN(n1292) );
XOR2_X1 U1090 ( .A(n1354), .B(n1355), .Z(n1343) );
XNOR2_X1 U1091 ( .A(n1187), .B(n1188), .ZN(n1355) );
AND2_X1 U1092 ( .A1(G227), .A2(n1057), .ZN(n1188) );
INV_X1 U1093 ( .A(G953), .ZN(n1057) );
INV_X1 U1094 ( .A(G140), .ZN(n1187) );
NOR2_X1 U1095 ( .A1(KEYINPUT1), .A2(G110), .ZN(n1354) );
INV_X1 U1096 ( .A(G110), .ZN(n1185) );
endmodule


