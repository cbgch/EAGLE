//Key = 1000111111001110000100010111010011101001101010011100010101111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351;

XNOR2_X1 U747 ( .A(n1029), .B(n1030), .ZN(G9) );
NAND4_X1 U748 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(G75) );
NAND4_X1 U749 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1033) );
NOR4_X1 U750 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1038) );
XOR2_X1 U751 ( .A(n1043), .B(KEYINPUT63), .Z(n1042) );
NAND2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U753 ( .A1(G475), .A2(n1046), .ZN(n1045) );
XOR2_X1 U754 ( .A(n1047), .B(KEYINPUT19), .Z(n1041) );
XOR2_X1 U755 ( .A(n1048), .B(n1049), .Z(n1040) );
NOR2_X1 U756 ( .A1(n1050), .A2(KEYINPUT31), .ZN(n1049) );
XNOR2_X1 U757 ( .A(n1051), .B(n1052), .ZN(n1036) );
NOR2_X1 U758 ( .A1(KEYINPUT15), .A2(n1053), .ZN(n1051) );
XOR2_X1 U759 ( .A(KEYINPUT11), .B(G472), .Z(n1053) );
NAND2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1032) );
NAND2_X1 U761 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND3_X1 U762 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
NAND2_X1 U763 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND2_X1 U764 ( .A1(n1037), .A2(n1063), .ZN(n1062) );
OR2_X1 U765 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(n1061) );
NAND2_X1 U767 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND3_X1 U769 ( .A1(n1037), .A2(n1072), .A3(n1066), .ZN(n1056) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U771 ( .A1(n1060), .A2(n1075), .ZN(n1074) );
NAND2_X1 U772 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U773 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U774 ( .A1(n1058), .A2(n1080), .ZN(n1073) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U776 ( .A1(n1039), .A2(n1083), .ZN(n1082) );
INV_X1 U777 ( .A(n1084), .ZN(n1081) );
INV_X1 U778 ( .A(n1085), .ZN(n1054) );
XOR2_X1 U779 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U780 ( .A1(n1088), .A2(n1034), .ZN(n1087) );
AND2_X1 U781 ( .A1(G227), .A2(G900), .ZN(n1088) );
NAND2_X1 U782 ( .A1(n1089), .A2(n1090), .ZN(n1086) );
NAND2_X1 U783 ( .A1(n1091), .A2(n1034), .ZN(n1090) );
XOR2_X1 U784 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
XNOR2_X1 U786 ( .A(n1096), .B(KEYINPUT10), .ZN(n1094) );
NAND3_X1 U787 ( .A1(G900), .A2(n1093), .A3(G953), .ZN(n1089) );
XNOR2_X1 U788 ( .A(n1097), .B(n1098), .ZN(n1093) );
NOR2_X1 U789 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U790 ( .A(n1101), .B(KEYINPUT25), .Z(n1100) );
NAND2_X1 U791 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U792 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
AND2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U795 ( .A(n1108), .B(n1109), .ZN(n1106) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1104) );
XNOR2_X1 U797 ( .A(G134), .B(n1109), .ZN(n1111) );
NOR2_X1 U798 ( .A1(G137), .A2(KEYINPUT3), .ZN(n1109) );
XNOR2_X1 U799 ( .A(G131), .B(KEYINPUT29), .ZN(n1110) );
NAND2_X1 U800 ( .A1(KEYINPUT53), .A2(n1112), .ZN(n1097) );
XOR2_X1 U801 ( .A(KEYINPUT37), .B(n1113), .Z(n1112) );
NOR2_X1 U802 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U803 ( .A(n1116), .B(KEYINPUT5), .Z(n1115) );
NAND2_X1 U804 ( .A1(G140), .A2(n1117), .ZN(n1116) );
NOR2_X1 U805 ( .A1(G140), .A2(n1118), .ZN(n1114) );
XNOR2_X1 U806 ( .A(G125), .B(KEYINPUT20), .ZN(n1118) );
XOR2_X1 U807 ( .A(n1119), .B(n1120), .Z(G69) );
NOR2_X1 U808 ( .A1(n1121), .A2(n1034), .ZN(n1120) );
NOR2_X1 U809 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U810 ( .A1(n1124), .A2(n1125), .ZN(n1119) );
OR3_X1 U811 ( .A1(n1126), .A2(G953), .A3(n1127), .ZN(n1125) );
NAND3_X1 U812 ( .A1(n1128), .A2(n1129), .A3(n1127), .ZN(n1124) );
XNOR2_X1 U813 ( .A(n1130), .B(n1131), .ZN(n1127) );
XOR2_X1 U814 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U816 ( .A(n1136), .B(KEYINPUT27), .Z(n1135) );
NAND2_X1 U817 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NOR2_X1 U818 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
XNOR2_X1 U819 ( .A(n1139), .B(G116), .ZN(n1137) );
XNOR2_X1 U820 ( .A(G122), .B(KEYINPUT38), .ZN(n1130) );
NAND2_X1 U821 ( .A1(G953), .A2(n1123), .ZN(n1129) );
XOR2_X1 U822 ( .A(KEYINPUT1), .B(n1126), .Z(n1128) );
NOR2_X1 U823 ( .A1(n1140), .A2(n1141), .ZN(G66) );
XOR2_X1 U824 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U825 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
NOR2_X1 U826 ( .A1(n1140), .A2(n1146), .ZN(G63) );
XOR2_X1 U827 ( .A(n1147), .B(n1148), .Z(n1146) );
AND2_X1 U828 ( .A1(G478), .A2(n1149), .ZN(n1147) );
NOR2_X1 U829 ( .A1(n1140), .A2(n1150), .ZN(G60) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U831 ( .A(KEYINPUT4), .B(n1153), .ZN(n1151) );
NOR3_X1 U832 ( .A1(n1145), .A2(KEYINPUT46), .A3(n1154), .ZN(n1153) );
XNOR2_X1 U833 ( .A(G104), .B(n1155), .ZN(G6) );
NOR2_X1 U834 ( .A1(n1140), .A2(n1156), .ZN(G57) );
XOR2_X1 U835 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U836 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U837 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U838 ( .A1(n1163), .A2(n1164), .ZN(n1159) );
XOR2_X1 U839 ( .A(n1162), .B(KEYINPUT8), .Z(n1164) );
XOR2_X1 U840 ( .A(n1165), .B(n1166), .Z(n1162) );
XOR2_X1 U841 ( .A(n1167), .B(n1168), .Z(n1165) );
NAND2_X1 U842 ( .A1(KEYINPUT60), .A2(n1169), .ZN(n1167) );
INV_X1 U843 ( .A(n1161), .ZN(n1163) );
NAND2_X1 U844 ( .A1(n1170), .A2(n1149), .ZN(n1161) );
XNOR2_X1 U845 ( .A(G472), .B(KEYINPUT49), .ZN(n1170) );
NOR2_X1 U846 ( .A1(KEYINPUT50), .A2(n1171), .ZN(n1157) );
NOR2_X1 U847 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XNOR2_X1 U848 ( .A(n1174), .B(KEYINPUT13), .ZN(n1173) );
NOR3_X1 U849 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(G54) );
AND3_X1 U850 ( .A1(KEYINPUT18), .A2(G953), .A3(G952), .ZN(n1177) );
NOR2_X1 U851 ( .A1(KEYINPUT18), .A2(n1178), .ZN(n1176) );
INV_X1 U852 ( .A(n1140), .ZN(n1178) );
NOR3_X1 U853 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1175) );
NOR3_X1 U854 ( .A1(n1182), .A2(KEYINPUT28), .A3(n1183), .ZN(n1181) );
INV_X1 U855 ( .A(n1184), .ZN(n1182) );
NOR2_X1 U856 ( .A1(n1185), .A2(n1184), .ZN(n1180) );
XNOR2_X1 U857 ( .A(n1186), .B(n1187), .ZN(n1184) );
NAND2_X1 U858 ( .A1(KEYINPUT36), .A2(n1188), .ZN(n1186) );
NOR2_X1 U859 ( .A1(KEYINPUT28), .A2(n1189), .ZN(n1185) );
XOR2_X1 U860 ( .A(KEYINPUT62), .B(n1183), .Z(n1189) );
AND2_X1 U861 ( .A1(n1183), .A2(KEYINPUT28), .ZN(n1179) );
AND2_X1 U862 ( .A1(n1149), .A2(G469), .ZN(n1183) );
NOR2_X1 U863 ( .A1(n1140), .A2(n1190), .ZN(G51) );
XOR2_X1 U864 ( .A(n1191), .B(n1192), .Z(n1190) );
XNOR2_X1 U865 ( .A(n1117), .B(n1193), .ZN(n1192) );
NOR2_X1 U866 ( .A1(n1048), .A2(n1145), .ZN(n1193) );
INV_X1 U867 ( .A(n1149), .ZN(n1145) );
NOR2_X1 U868 ( .A1(n1194), .A2(n1031), .ZN(n1149) );
AND3_X1 U869 ( .A1(n1095), .A2(n1195), .A3(n1126), .ZN(n1031) );
AND2_X1 U870 ( .A1(n1196), .A2(n1197), .ZN(n1126) );
NOR4_X1 U871 ( .A1(n1198), .A2(n1030), .A3(n1199), .A4(n1200), .ZN(n1197) );
INV_X1 U872 ( .A(n1201), .ZN(n1200) );
AND3_X1 U873 ( .A1(n1065), .A2(n1058), .A3(n1202), .ZN(n1030) );
AND4_X1 U874 ( .A1(n1203), .A2(n1204), .A3(n1155), .A4(n1205), .ZN(n1196) );
NAND3_X1 U875 ( .A1(n1206), .A2(n1207), .A3(n1065), .ZN(n1205) );
NAND3_X1 U876 ( .A1(n1202), .A2(n1058), .A3(n1064), .ZN(n1155) );
AND4_X1 U877 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1095) );
AND3_X1 U878 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
OR2_X1 U879 ( .A1(n1215), .A2(n1216), .ZN(n1212) );
NOR2_X1 U880 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
NOR2_X1 U881 ( .A1(n1034), .A2(G952), .ZN(n1140) );
XNOR2_X1 U882 ( .A(n1219), .B(n1210), .ZN(G48) );
NAND4_X1 U883 ( .A1(n1220), .A2(n1064), .A3(n1084), .A4(n1221), .ZN(n1210) );
NAND2_X1 U884 ( .A1(KEYINPUT6), .A2(n1222), .ZN(n1219) );
XNOR2_X1 U885 ( .A(G143), .B(n1214), .ZN(G45) );
NAND4_X1 U886 ( .A1(n1223), .A2(n1084), .A3(n1224), .A4(n1225), .ZN(n1214) );
XNOR2_X1 U887 ( .A(G140), .B(n1226), .ZN(G42) );
NAND3_X1 U888 ( .A1(n1218), .A2(n1227), .A3(KEYINPUT44), .ZN(n1226) );
XNOR2_X1 U889 ( .A(KEYINPUT30), .B(n1216), .ZN(n1227) );
AND3_X1 U890 ( .A1(n1078), .A2(n1064), .A3(n1220), .ZN(n1218) );
NAND3_X1 U891 ( .A1(n1228), .A2(n1229), .A3(n1230), .ZN(G39) );
OR2_X1 U892 ( .A1(n1096), .A2(KEYINPUT32), .ZN(n1230) );
NAND3_X1 U893 ( .A1(KEYINPUT32), .A2(n1096), .A3(n1231), .ZN(n1229) );
NAND2_X1 U894 ( .A1(G137), .A2(n1232), .ZN(n1228) );
NAND2_X1 U895 ( .A1(n1233), .A2(KEYINPUT32), .ZN(n1232) );
XNOR2_X1 U896 ( .A(n1096), .B(KEYINPUT23), .ZN(n1233) );
INV_X1 U897 ( .A(n1195), .ZN(n1096) );
NAND4_X1 U898 ( .A1(n1060), .A2(n1220), .A3(n1066), .A4(n1221), .ZN(n1195) );
AND3_X1 U899 ( .A1(n1079), .A2(n1234), .A3(n1235), .ZN(n1220) );
XNOR2_X1 U900 ( .A(G134), .B(n1236), .ZN(G36) );
NAND2_X1 U901 ( .A1(n1060), .A2(n1237), .ZN(n1236) );
XOR2_X1 U902 ( .A(KEYINPUT54), .B(n1217), .Z(n1237) );
AND2_X1 U903 ( .A1(n1223), .A2(n1065), .ZN(n1217) );
XNOR2_X1 U904 ( .A(G131), .B(n1213), .ZN(G33) );
NAND3_X1 U905 ( .A1(n1060), .A2(n1064), .A3(n1223), .ZN(n1213) );
AND3_X1 U906 ( .A1(n1235), .A2(n1234), .A3(n1207), .ZN(n1223) );
INV_X1 U907 ( .A(n1216), .ZN(n1060) );
NAND2_X1 U908 ( .A1(n1083), .A2(n1238), .ZN(n1216) );
XNOR2_X1 U909 ( .A(G128), .B(n1208), .ZN(G30) );
NAND4_X1 U910 ( .A1(n1239), .A2(n1065), .A3(n1221), .A4(n1240), .ZN(n1208) );
XNOR2_X1 U911 ( .A(G101), .B(n1204), .ZN(G3) );
NAND3_X1 U912 ( .A1(n1202), .A2(n1207), .A3(n1066), .ZN(n1204) );
XNOR2_X1 U913 ( .A(G125), .B(n1209), .ZN(G27) );
NAND4_X1 U914 ( .A1(n1239), .A2(n1064), .A3(n1078), .A4(n1037), .ZN(n1209) );
INV_X1 U915 ( .A(n1241), .ZN(n1064) );
AND3_X1 U916 ( .A1(n1079), .A2(n1234), .A3(n1084), .ZN(n1239) );
NAND2_X1 U917 ( .A1(n1085), .A2(n1242), .ZN(n1234) );
NAND2_X1 U918 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
INV_X1 U919 ( .A(G900), .ZN(n1244) );
XNOR2_X1 U920 ( .A(G122), .B(n1203), .ZN(G24) );
NAND4_X1 U921 ( .A1(n1206), .A2(n1058), .A3(n1224), .A4(n1225), .ZN(n1203) );
NAND2_X1 U922 ( .A1(n1245), .A2(n1246), .ZN(n1058) );
NAND3_X1 U923 ( .A1(n1047), .A2(n1078), .A3(n1247), .ZN(n1246) );
INV_X1 U924 ( .A(KEYINPUT2), .ZN(n1247) );
NAND2_X1 U925 ( .A1(KEYINPUT2), .A2(n1207), .ZN(n1245) );
NAND2_X1 U926 ( .A1(n1248), .A2(n1249), .ZN(G21) );
OR2_X1 U927 ( .A1(n1201), .A2(G119), .ZN(n1249) );
XOR2_X1 U928 ( .A(n1250), .B(KEYINPUT43), .Z(n1248) );
NAND2_X1 U929 ( .A1(G119), .A2(n1201), .ZN(n1250) );
NAND4_X1 U930 ( .A1(n1066), .A2(n1206), .A3(n1079), .A4(n1221), .ZN(n1201) );
INV_X1 U931 ( .A(n1251), .ZN(n1206) );
XNOR2_X1 U932 ( .A(G116), .B(n1252), .ZN(G18) );
NAND3_X1 U933 ( .A1(n1253), .A2(n1037), .A3(n1254), .ZN(n1252) );
AND3_X1 U934 ( .A1(n1065), .A2(n1255), .A3(n1207), .ZN(n1254) );
INV_X1 U935 ( .A(n1076), .ZN(n1207) );
NOR2_X1 U936 ( .A1(n1225), .A2(n1035), .ZN(n1065) );
XNOR2_X1 U937 ( .A(n1084), .B(KEYINPUT26), .ZN(n1253) );
XOR2_X1 U938 ( .A(n1256), .B(n1198), .Z(G15) );
NOR3_X1 U939 ( .A1(n1251), .A2(n1076), .A3(n1241), .ZN(n1198) );
NAND2_X1 U940 ( .A1(n1035), .A2(n1225), .ZN(n1241) );
INV_X1 U941 ( .A(n1224), .ZN(n1035) );
NAND2_X1 U942 ( .A1(n1047), .A2(n1221), .ZN(n1076) );
INV_X1 U943 ( .A(n1078), .ZN(n1221) );
NAND3_X1 U944 ( .A1(n1084), .A2(n1255), .A3(n1037), .ZN(n1251) );
NOR2_X1 U945 ( .A1(n1257), .A2(n1070), .ZN(n1037) );
NAND2_X1 U946 ( .A1(KEYINPUT61), .A2(n1258), .ZN(n1256) );
XOR2_X1 U947 ( .A(G110), .B(n1199), .Z(G12) );
AND4_X1 U948 ( .A1(n1066), .A2(n1202), .A3(n1078), .A4(n1079), .ZN(n1199) );
XNOR2_X1 U949 ( .A(n1047), .B(KEYINPUT51), .ZN(n1079) );
XNOR2_X1 U950 ( .A(n1259), .B(n1144), .ZN(n1047) );
NAND2_X1 U951 ( .A1(G217), .A2(n1260), .ZN(n1144) );
OR2_X1 U952 ( .A1(n1143), .A2(G902), .ZN(n1259) );
XNOR2_X1 U953 ( .A(n1261), .B(n1262), .ZN(n1143) );
XOR2_X1 U954 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U955 ( .A(n1231), .B(G128), .ZN(n1264) );
INV_X1 U956 ( .A(G137), .ZN(n1231) );
XNOR2_X1 U957 ( .A(KEYINPUT58), .B(n1222), .ZN(n1263) );
XOR2_X1 U958 ( .A(n1265), .B(n1266), .Z(n1261) );
XNOR2_X1 U959 ( .A(n1117), .B(G119), .ZN(n1266) );
XNOR2_X1 U960 ( .A(n1267), .B(n1268), .ZN(n1265) );
NAND2_X1 U961 ( .A1(n1269), .A2(G221), .ZN(n1267) );
XOR2_X1 U962 ( .A(n1052), .B(G472), .Z(n1078) );
NAND2_X1 U963 ( .A1(n1270), .A2(n1194), .ZN(n1052) );
XOR2_X1 U964 ( .A(n1168), .B(n1271), .Z(n1270) );
XOR2_X1 U965 ( .A(n1272), .B(n1273), .Z(n1271) );
NOR2_X1 U966 ( .A1(KEYINPUT21), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U967 ( .A(n1169), .B(n1166), .ZN(n1274) );
XNOR2_X1 U968 ( .A(n1275), .B(KEYINPUT40), .ZN(n1166) );
NOR2_X1 U969 ( .A1(n1174), .A2(n1172), .ZN(n1272) );
NOR2_X1 U970 ( .A1(G101), .A2(n1276), .ZN(n1172) );
NOR2_X1 U971 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NOR3_X1 U972 ( .A1(n1277), .A2(n1279), .A3(n1278), .ZN(n1174) );
INV_X1 U973 ( .A(n1280), .ZN(n1278) );
INV_X1 U974 ( .A(G210), .ZN(n1277) );
XNOR2_X1 U975 ( .A(n1281), .B(n1282), .ZN(n1168) );
XNOR2_X1 U976 ( .A(G119), .B(n1258), .ZN(n1282) );
NAND2_X1 U977 ( .A1(KEYINPUT12), .A2(n1283), .ZN(n1281) );
INV_X1 U978 ( .A(G116), .ZN(n1283) );
AND3_X1 U979 ( .A1(n1240), .A2(n1255), .A3(n1084), .ZN(n1202) );
NOR2_X1 U980 ( .A1(n1083), .A2(n1039), .ZN(n1084) );
INV_X1 U981 ( .A(n1238), .ZN(n1039) );
NAND2_X1 U982 ( .A1(G214), .A2(n1284), .ZN(n1238) );
XOR2_X1 U983 ( .A(n1050), .B(n1048), .Z(n1083) );
NAND2_X1 U984 ( .A1(G210), .A2(n1284), .ZN(n1048) );
NAND2_X1 U985 ( .A1(n1285), .A2(n1194), .ZN(n1284) );
INV_X1 U986 ( .A(G237), .ZN(n1285) );
AND2_X1 U987 ( .A1(n1286), .A2(n1194), .ZN(n1050) );
XNOR2_X1 U988 ( .A(n1191), .B(n1287), .ZN(n1286) );
NOR2_X1 U989 ( .A1(KEYINPUT45), .A2(n1117), .ZN(n1287) );
INV_X1 U990 ( .A(G125), .ZN(n1117) );
XNOR2_X1 U991 ( .A(n1288), .B(n1289), .ZN(n1191) );
XOR2_X1 U992 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U993 ( .A(n1275), .B(n1292), .Z(n1291) );
NOR2_X1 U994 ( .A1(G953), .A2(n1122), .ZN(n1292) );
INV_X1 U995 ( .A(G224), .ZN(n1122) );
XNOR2_X1 U996 ( .A(G128), .B(n1293), .ZN(n1275) );
XNOR2_X1 U997 ( .A(n1132), .B(KEYINPUT48), .ZN(n1290) );
NOR2_X1 U998 ( .A1(KEYINPUT16), .A2(G110), .ZN(n1132) );
XNOR2_X1 U999 ( .A(n1294), .B(n1295), .ZN(n1288) );
INV_X1 U1000 ( .A(n1139), .ZN(n1295) );
XNOR2_X1 U1001 ( .A(n1296), .B(G119), .ZN(n1139) );
NAND2_X1 U1002 ( .A1(KEYINPUT47), .A2(G113), .ZN(n1296) );
XNOR2_X1 U1003 ( .A(n1138), .B(n1297), .ZN(n1294) );
XNOR2_X1 U1004 ( .A(n1298), .B(n1299), .ZN(n1138) );
NAND2_X1 U1005 ( .A1(n1300), .A2(KEYINPUT39), .ZN(n1298) );
XNOR2_X1 U1006 ( .A(n1301), .B(KEYINPUT55), .ZN(n1300) );
NAND2_X1 U1007 ( .A1(n1085), .A2(n1302), .ZN(n1255) );
NAND2_X1 U1008 ( .A1(n1243), .A2(n1123), .ZN(n1302) );
INV_X1 U1009 ( .A(G898), .ZN(n1123) );
AND3_X1 U1010 ( .A1(G953), .A2(n1303), .A3(n1304), .ZN(n1243) );
XNOR2_X1 U1011 ( .A(G902), .B(KEYINPUT9), .ZN(n1304) );
NAND3_X1 U1012 ( .A1(n1303), .A2(n1034), .A3(G952), .ZN(n1085) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1303) );
XNOR2_X1 U1014 ( .A(n1068), .B(KEYINPUT35), .ZN(n1240) );
INV_X1 U1015 ( .A(n1235), .ZN(n1068) );
NOR2_X1 U1016 ( .A1(n1071), .A2(n1070), .ZN(n1235) );
AND2_X1 U1017 ( .A1(G221), .A2(n1260), .ZN(n1070) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1194), .ZN(n1260) );
INV_X1 U1019 ( .A(n1257), .ZN(n1071) );
XNOR2_X1 U1020 ( .A(n1305), .B(n1306), .ZN(n1257) );
XOR2_X1 U1021 ( .A(KEYINPUT22), .B(G469), .Z(n1306) );
NAND2_X1 U1022 ( .A1(n1307), .A2(n1194), .ZN(n1305) );
INV_X1 U1023 ( .A(G902), .ZN(n1194) );
XNOR2_X1 U1024 ( .A(n1188), .B(n1308), .ZN(n1307) );
XOR2_X1 U1025 ( .A(KEYINPUT52), .B(n1309), .Z(n1308) );
NOR2_X1 U1026 ( .A1(KEYINPUT24), .A2(n1187), .ZN(n1309) );
AND2_X1 U1027 ( .A1(n1310), .A2(n1311), .ZN(n1187) );
NAND2_X1 U1028 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1029 ( .A1(G227), .A2(n1034), .ZN(n1313) );
INV_X1 U1030 ( .A(n1268), .ZN(n1312) );
NAND3_X1 U1031 ( .A1(G227), .A2(n1034), .A3(n1268), .ZN(n1310) );
XOR2_X1 U1032 ( .A(G110), .B(n1314), .Z(n1268) );
INV_X1 U1033 ( .A(G140), .ZN(n1314) );
XNOR2_X1 U1034 ( .A(n1315), .B(n1316), .ZN(n1188) );
XNOR2_X1 U1035 ( .A(n1317), .B(n1299), .ZN(n1316) );
XNOR2_X1 U1036 ( .A(n1279), .B(n1318), .ZN(n1299) );
XNOR2_X1 U1037 ( .A(KEYINPUT17), .B(n1029), .ZN(n1318) );
INV_X1 U1038 ( .A(G101), .ZN(n1279) );
INV_X1 U1039 ( .A(n1301), .ZN(n1317) );
XOR2_X1 U1040 ( .A(G104), .B(KEYINPUT42), .Z(n1301) );
XNOR2_X1 U1041 ( .A(n1319), .B(n1103), .ZN(n1315) );
XOR2_X1 U1042 ( .A(n1320), .B(n1293), .Z(n1103) );
XNOR2_X1 U1043 ( .A(n1321), .B(G146), .ZN(n1293) );
NAND2_X1 U1044 ( .A1(KEYINPUT7), .A2(n1322), .ZN(n1320) );
INV_X1 U1045 ( .A(G128), .ZN(n1322) );
XNOR2_X1 U1046 ( .A(n1169), .B(KEYINPUT57), .ZN(n1319) );
AND2_X1 U1047 ( .A1(n1323), .A2(n1324), .ZN(n1169) );
OR2_X1 U1048 ( .A1(n1325), .A2(G131), .ZN(n1324) );
XOR2_X1 U1049 ( .A(n1326), .B(KEYINPUT56), .Z(n1323) );
NAND2_X1 U1050 ( .A1(G131), .A2(n1325), .ZN(n1326) );
XNOR2_X1 U1051 ( .A(G137), .B(n1108), .ZN(n1325) );
INV_X1 U1052 ( .A(G134), .ZN(n1108) );
NOR2_X1 U1053 ( .A1(n1224), .A2(n1225), .ZN(n1066) );
NAND3_X1 U1054 ( .A1(n1327), .A2(n1328), .A3(n1044), .ZN(n1225) );
NAND2_X1 U1055 ( .A1(n1329), .A2(n1154), .ZN(n1044) );
INV_X1 U1056 ( .A(G475), .ZN(n1154) );
OR2_X1 U1057 ( .A1(G475), .A2(KEYINPUT14), .ZN(n1328) );
NAND3_X1 U1058 ( .A1(G475), .A2(n1046), .A3(KEYINPUT14), .ZN(n1327) );
INV_X1 U1059 ( .A(n1329), .ZN(n1046) );
NOR2_X1 U1060 ( .A1(n1152), .A2(G902), .ZN(n1329) );
XNOR2_X1 U1061 ( .A(n1330), .B(n1331), .ZN(n1152) );
XOR2_X1 U1062 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1063 ( .A(n1334), .B(n1335), .ZN(n1333) );
NAND2_X1 U1064 ( .A1(KEYINPUT59), .A2(n1222), .ZN(n1335) );
INV_X1 U1065 ( .A(G146), .ZN(n1222) );
NAND2_X1 U1066 ( .A1(n1336), .A2(KEYINPUT33), .ZN(n1334) );
XNOR2_X1 U1067 ( .A(n1337), .B(n1258), .ZN(n1336) );
INV_X1 U1068 ( .A(G113), .ZN(n1258) );
NAND2_X1 U1069 ( .A1(KEYINPUT34), .A2(n1338), .ZN(n1337) );
XOR2_X1 U1070 ( .A(n1339), .B(G104), .Z(n1332) );
NAND2_X1 U1071 ( .A1(n1280), .A2(G214), .ZN(n1339) );
NOR2_X1 U1072 ( .A1(G953), .A2(G237), .ZN(n1280) );
XOR2_X1 U1073 ( .A(n1340), .B(n1341), .Z(n1330) );
XNOR2_X1 U1074 ( .A(n1107), .B(G125), .ZN(n1341) );
INV_X1 U1075 ( .A(G131), .ZN(n1107) );
XNOR2_X1 U1076 ( .A(G140), .B(G143), .ZN(n1340) );
XNOR2_X1 U1077 ( .A(n1342), .B(G478), .ZN(n1224) );
OR2_X1 U1078 ( .A1(n1148), .A2(G902), .ZN(n1342) );
XNOR2_X1 U1079 ( .A(n1343), .B(n1344), .ZN(n1148) );
XNOR2_X1 U1080 ( .A(n1345), .B(n1297), .ZN(n1344) );
XNOR2_X1 U1081 ( .A(G116), .B(n1338), .ZN(n1297) );
INV_X1 U1082 ( .A(G122), .ZN(n1338) );
NAND2_X1 U1083 ( .A1(G217), .A2(n1269), .ZN(n1345) );
AND2_X1 U1084 ( .A1(G234), .A2(n1034), .ZN(n1269) );
INV_X1 U1085 ( .A(G953), .ZN(n1034) );
XOR2_X1 U1086 ( .A(n1346), .B(n1347), .Z(n1343) );
NOR2_X1 U1087 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1088 ( .A(KEYINPUT41), .B(n1350), .Z(n1349) );
NOR2_X1 U1089 ( .A1(G134), .A2(n1351), .ZN(n1350) );
AND2_X1 U1090 ( .A1(n1351), .A2(G134), .ZN(n1348) );
XNOR2_X1 U1091 ( .A(G128), .B(n1321), .ZN(n1351) );
INV_X1 U1092 ( .A(G143), .ZN(n1321) );
NAND2_X1 U1093 ( .A1(KEYINPUT0), .A2(n1029), .ZN(n1346) );
INV_X1 U1094 ( .A(G107), .ZN(n1029) );
endmodule


