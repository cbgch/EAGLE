//Key = 0000111011000111111011101000001001110100000100011001010101010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
n1436, n1437, n1438, n1439, n1440;

XNOR2_X1 U796 ( .A(G107), .B(n1096), .ZN(G9) );
NAND4_X1 U797 ( .A1(KEYINPUT57), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1096) );
NOR2_X1 U798 ( .A1(n1100), .A2(n1101), .ZN(G75) );
NOR3_X1 U799 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NOR2_X1 U800 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
INV_X1 U801 ( .A(n1107), .ZN(n1106) );
NOR2_X1 U802 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NOR2_X1 U803 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
AND4_X1 U804 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1110) );
NOR4_X1 U805 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1108) );
INV_X1 U806 ( .A(n1098), .ZN(n1117) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1121), .ZN(n1116) );
NOR2_X1 U808 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NAND3_X1 U809 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1102) );
NAND3_X1 U810 ( .A1(n1114), .A2(n1127), .A3(n1115), .ZN(n1126) );
INV_X1 U811 ( .A(n1119), .ZN(n1115) );
NAND2_X1 U812 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U813 ( .A1(n1107), .A2(n1130), .ZN(n1129) );
NAND2_X1 U814 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U815 ( .A1(n1133), .A2(n1098), .ZN(n1132) );
NAND2_X1 U816 ( .A1(n1113), .A2(n1134), .ZN(n1128) );
NAND2_X1 U817 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND3_X1 U818 ( .A1(n1107), .A2(n1111), .A3(n1112), .ZN(n1136) );
INV_X1 U819 ( .A(KEYINPUT1), .ZN(n1111) );
NAND2_X1 U820 ( .A1(n1098), .A2(n1137), .ZN(n1135) );
NAND2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U822 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR3_X1 U823 ( .A1(n1142), .A2(G953), .A3(G952), .ZN(n1100) );
INV_X1 U824 ( .A(n1124), .ZN(n1142) );
NAND4_X1 U825 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1124) );
NOR3_X1 U826 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
XNOR2_X1 U827 ( .A(n1150), .B(n1151), .ZN(n1149) );
NAND2_X1 U828 ( .A1(KEYINPUT37), .A2(n1152), .ZN(n1150) );
NOR2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1148) );
NAND3_X1 U830 ( .A1(n1123), .A2(n1155), .A3(n1156), .ZN(n1147) );
NOR3_X1 U831 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1145) );
XOR2_X1 U832 ( .A(n1160), .B(KEYINPUT24), .Z(n1158) );
NAND2_X1 U833 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XNOR2_X1 U834 ( .A(KEYINPUT49), .B(n1163), .ZN(n1161) );
XNOR2_X1 U835 ( .A(n1164), .B(n1165), .ZN(n1157) );
NAND2_X1 U836 ( .A1(KEYINPUT15), .A2(G475), .ZN(n1165) );
XOR2_X1 U837 ( .A(n1166), .B(KEYINPUT50), .Z(n1144) );
NAND2_X1 U838 ( .A1(n1153), .A2(n1154), .ZN(n1166) );
XNOR2_X1 U839 ( .A(n1167), .B(n1141), .ZN(n1143) );
XNOR2_X1 U840 ( .A(KEYINPUT7), .B(KEYINPUT44), .ZN(n1167) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(G72) );
NOR2_X1 U842 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XOR2_X1 U843 ( .A(n1172), .B(KEYINPUT9), .Z(n1171) );
NAND3_X1 U844 ( .A1(n1173), .A2(n1125), .A3(n1174), .ZN(n1172) );
NOR3_X1 U845 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1170) );
AND2_X1 U846 ( .A1(n1125), .A2(n1173), .ZN(n1176) );
NAND2_X1 U847 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
XNOR2_X1 U848 ( .A(KEYINPUT16), .B(n1179), .ZN(n1178) );
NOR2_X1 U849 ( .A1(G900), .A2(n1125), .ZN(n1175) );
XOR2_X1 U850 ( .A(n1180), .B(n1181), .Z(n1174) );
XNOR2_X1 U851 ( .A(n1182), .B(n1183), .ZN(n1181) );
NAND2_X1 U852 ( .A1(KEYINPUT43), .A2(G140), .ZN(n1182) );
XOR2_X1 U853 ( .A(n1184), .B(n1185), .Z(n1180) );
XNOR2_X1 U854 ( .A(G125), .B(n1186), .ZN(n1185) );
NAND2_X1 U855 ( .A1(KEYINPUT17), .A2(G131), .ZN(n1184) );
NAND2_X1 U856 ( .A1(G953), .A2(n1187), .ZN(n1168) );
NAND2_X1 U857 ( .A1(G900), .A2(G227), .ZN(n1187) );
XOR2_X1 U858 ( .A(n1188), .B(n1189), .Z(G69) );
NOR2_X1 U859 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XOR2_X1 U860 ( .A(n1192), .B(KEYINPUT28), .Z(n1191) );
NAND2_X1 U861 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NAND2_X1 U862 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U863 ( .A(n1197), .B(KEYINPUT11), .Z(n1193) );
OR2_X1 U864 ( .A1(n1196), .A2(n1195), .ZN(n1197) );
XNOR2_X1 U865 ( .A(n1198), .B(n1199), .ZN(n1196) );
NAND3_X1 U866 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1188) );
NAND2_X1 U867 ( .A1(KEYINPUT21), .A2(n1203), .ZN(n1202) );
NAND2_X1 U868 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
OR2_X1 U869 ( .A1(n1125), .A2(G224), .ZN(n1205) );
INV_X1 U870 ( .A(n1190), .ZN(n1204) );
NAND4_X1 U871 ( .A1(G224), .A2(n1206), .A3(G898), .A4(G953), .ZN(n1201) );
INV_X1 U872 ( .A(KEYINPUT21), .ZN(n1206) );
NAND2_X1 U873 ( .A1(n1207), .A2(n1125), .ZN(n1200) );
NAND2_X1 U874 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NOR2_X1 U875 ( .A1(n1210), .A2(n1211), .ZN(G66) );
XOR2_X1 U876 ( .A(n1212), .B(n1213), .Z(n1211) );
NOR2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
NOR2_X1 U878 ( .A1(n1210), .A2(n1216), .ZN(G63) );
XOR2_X1 U879 ( .A(n1217), .B(n1218), .Z(n1216) );
XOR2_X1 U880 ( .A(KEYINPUT19), .B(n1219), .Z(n1218) );
NOR2_X1 U881 ( .A1(n1163), .A2(n1215), .ZN(n1219) );
INV_X1 U882 ( .A(G478), .ZN(n1163) );
NOR2_X1 U883 ( .A1(KEYINPUT56), .A2(n1220), .ZN(n1217) );
NOR2_X1 U884 ( .A1(n1210), .A2(n1221), .ZN(G60) );
NOR3_X1 U885 ( .A1(n1164), .A2(n1222), .A3(n1223), .ZN(n1221) );
NOR3_X1 U886 ( .A1(n1224), .A2(n1225), .A3(n1215), .ZN(n1223) );
INV_X1 U887 ( .A(n1226), .ZN(n1224) );
NOR2_X1 U888 ( .A1(n1227), .A2(n1226), .ZN(n1222) );
AND2_X1 U889 ( .A1(n1104), .A2(G475), .ZN(n1227) );
XNOR2_X1 U890 ( .A(G104), .B(n1228), .ZN(G6) );
NOR2_X1 U891 ( .A1(n1229), .A2(n1230), .ZN(G57) );
XOR2_X1 U892 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U893 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U894 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U895 ( .A1(n1154), .A2(n1215), .ZN(n1236) );
INV_X1 U896 ( .A(G472), .ZN(n1154) );
NAND2_X1 U897 ( .A1(KEYINPUT8), .A2(n1237), .ZN(n1235) );
NAND2_X1 U898 ( .A1(KEYINPUT63), .A2(n1238), .ZN(n1233) );
XOR2_X1 U899 ( .A(n1239), .B(n1240), .Z(n1231) );
NOR2_X1 U900 ( .A1(n1125), .A2(n1241), .ZN(n1229) );
XOR2_X1 U901 ( .A(KEYINPUT31), .B(G952), .Z(n1241) );
NOR2_X1 U902 ( .A1(n1210), .A2(n1242), .ZN(G54) );
XOR2_X1 U903 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U904 ( .A(n1245), .B(n1237), .Z(n1244) );
NAND2_X1 U905 ( .A1(KEYINPUT20), .A2(n1246), .ZN(n1245) );
INV_X1 U906 ( .A(n1247), .ZN(n1246) );
XOR2_X1 U907 ( .A(n1248), .B(n1249), .Z(n1243) );
XNOR2_X1 U908 ( .A(n1186), .B(n1250), .ZN(n1249) );
NOR3_X1 U909 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1250) );
NOR2_X1 U910 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NOR2_X1 U911 ( .A1(G953), .A2(KEYINPUT40), .ZN(n1254) );
NOR2_X1 U912 ( .A1(KEYINPUT40), .A2(n1256), .ZN(n1251) );
NOR2_X1 U913 ( .A1(n1151), .A2(n1215), .ZN(n1248) );
NAND2_X1 U914 ( .A1(G902), .A2(n1104), .ZN(n1215) );
NOR2_X1 U915 ( .A1(n1210), .A2(n1257), .ZN(G51) );
XOR2_X1 U916 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U917 ( .A(n1260), .B(n1261), .Z(n1259) );
NAND3_X1 U918 ( .A1(n1262), .A2(n1104), .A3(n1263), .ZN(n1260) );
XNOR2_X1 U919 ( .A(G902), .B(KEYINPUT53), .ZN(n1263) );
NAND4_X1 U920 ( .A1(n1264), .A2(n1177), .A3(n1208), .A4(n1179), .ZN(n1104) );
AND4_X1 U921 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1208) );
NOR3_X1 U922 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1268) );
NOR2_X1 U923 ( .A1(n1131), .A2(n1272), .ZN(n1271) );
INV_X1 U924 ( .A(n1099), .ZN(n1272) );
AND2_X1 U925 ( .A1(n1273), .A2(n1274), .ZN(n1131) );
NAND2_X1 U926 ( .A1(n1097), .A2(n1098), .ZN(n1274) );
NAND2_X1 U927 ( .A1(n1275), .A2(n1113), .ZN(n1273) );
INV_X1 U928 ( .A(n1228), .ZN(n1270) );
NAND3_X1 U929 ( .A1(n1098), .A2(n1099), .A3(n1133), .ZN(n1228) );
NOR2_X1 U930 ( .A1(n1138), .A2(n1276), .ZN(n1269) );
AND4_X1 U931 ( .A1(n1277), .A2(n1278), .A3(n1279), .A4(n1280), .ZN(n1177) );
AND4_X1 U932 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1280) );
NAND2_X1 U933 ( .A1(n1285), .A2(n1286), .ZN(n1279) );
XNOR2_X1 U934 ( .A(n1275), .B(KEYINPUT30), .ZN(n1285) );
NAND3_X1 U935 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1277) );
XNOR2_X1 U936 ( .A(n1121), .B(KEYINPUT6), .ZN(n1289) );
INV_X1 U937 ( .A(n1290), .ZN(n1121) );
XOR2_X1 U938 ( .A(n1209), .B(KEYINPUT0), .Z(n1264) );
NAND2_X1 U939 ( .A1(KEYINPUT35), .A2(n1291), .ZN(n1258) );
NOR2_X1 U940 ( .A1(n1125), .A2(G952), .ZN(n1210) );
XNOR2_X1 U941 ( .A(G146), .B(n1292), .ZN(G48) );
NAND2_X1 U942 ( .A1(n1287), .A2(n1293), .ZN(n1292) );
AND2_X1 U943 ( .A1(n1133), .A2(n1294), .ZN(n1287) );
XNOR2_X1 U944 ( .A(G143), .B(n1278), .ZN(G45) );
NAND3_X1 U945 ( .A1(n1112), .A2(n1293), .A3(n1295), .ZN(n1278) );
XNOR2_X1 U946 ( .A(G140), .B(n1296), .ZN(G42) );
NAND2_X1 U947 ( .A1(n1275), .A2(n1286), .ZN(n1296) );
XNOR2_X1 U948 ( .A(G137), .B(n1284), .ZN(G39) );
NAND4_X1 U949 ( .A1(n1113), .A2(n1297), .A3(n1298), .A4(n1159), .ZN(n1284) );
XNOR2_X1 U950 ( .A(G134), .B(n1283), .ZN(G36) );
NAND3_X1 U951 ( .A1(n1297), .A2(n1097), .A3(n1112), .ZN(n1283) );
NAND2_X1 U952 ( .A1(n1299), .A2(n1300), .ZN(G33) );
NAND2_X1 U953 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U954 ( .A1(G131), .A2(n1303), .ZN(n1302) );
OR2_X1 U955 ( .A1(n1304), .A2(KEYINPUT5), .ZN(n1303) );
INV_X1 U956 ( .A(n1282), .ZN(n1301) );
NAND3_X1 U957 ( .A1(n1305), .A2(n1306), .A3(KEYINPUT5), .ZN(n1299) );
NAND2_X1 U958 ( .A1(G131), .A2(n1304), .ZN(n1306) );
INV_X1 U959 ( .A(KEYINPUT18), .ZN(n1304) );
NAND2_X1 U960 ( .A1(KEYINPUT18), .A2(n1307), .ZN(n1305) );
NAND2_X1 U961 ( .A1(G131), .A2(n1282), .ZN(n1307) );
NAND2_X1 U962 ( .A1(n1112), .A2(n1286), .ZN(n1282) );
AND2_X1 U963 ( .A1(n1133), .A2(n1297), .ZN(n1286) );
AND2_X1 U964 ( .A1(n1107), .A2(n1293), .ZN(n1297) );
NOR2_X1 U965 ( .A1(n1308), .A2(n1140), .ZN(n1107) );
XNOR2_X1 U966 ( .A(n1309), .B(n1310), .ZN(G30) );
NOR2_X1 U967 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NOR2_X1 U968 ( .A1(KEYINPUT39), .A2(n1313), .ZN(n1312) );
INV_X1 U969 ( .A(n1281), .ZN(n1313) );
NOR2_X1 U970 ( .A1(KEYINPUT59), .A2(n1281), .ZN(n1311) );
NAND3_X1 U971 ( .A1(n1294), .A2(n1097), .A3(n1293), .ZN(n1281) );
NOR2_X1 U972 ( .A1(n1290), .A2(n1314), .ZN(n1293) );
XNOR2_X1 U973 ( .A(n1238), .B(n1315), .ZN(G3) );
NOR2_X1 U974 ( .A1(KEYINPUT36), .A2(n1209), .ZN(n1315) );
NAND3_X1 U975 ( .A1(n1112), .A2(n1099), .A3(n1113), .ZN(n1209) );
NOR3_X1 U976 ( .A1(n1290), .A2(n1316), .A3(n1138), .ZN(n1099) );
XNOR2_X1 U977 ( .A(G125), .B(n1179), .ZN(G27) );
NAND4_X1 U978 ( .A1(n1114), .A2(n1275), .A3(n1317), .A4(n1133), .ZN(n1179) );
NOR2_X1 U979 ( .A1(n1314), .A2(n1138), .ZN(n1317) );
INV_X1 U980 ( .A(n1288), .ZN(n1314) );
NAND2_X1 U981 ( .A1(n1119), .A2(n1318), .ZN(n1288) );
NAND4_X1 U982 ( .A1(G902), .A2(G953), .A3(n1319), .A4(n1320), .ZN(n1318) );
INV_X1 U983 ( .A(G900), .ZN(n1320) );
XNOR2_X1 U984 ( .A(G122), .B(n1267), .ZN(G24) );
NAND3_X1 U985 ( .A1(n1295), .A2(n1098), .A3(n1321), .ZN(n1267) );
NOR2_X1 U986 ( .A1(n1159), .A2(n1298), .ZN(n1098) );
NOR3_X1 U987 ( .A1(n1138), .A2(n1322), .A3(n1323), .ZN(n1295) );
INV_X1 U988 ( .A(n1324), .ZN(n1138) );
XOR2_X1 U989 ( .A(n1265), .B(n1325), .Z(G21) );
XNOR2_X1 U990 ( .A(KEYINPUT4), .B(n1326), .ZN(n1325) );
NAND3_X1 U991 ( .A1(n1113), .A2(n1294), .A3(n1321), .ZN(n1265) );
AND3_X1 U992 ( .A1(n1324), .A2(n1159), .A3(n1298), .ZN(n1294) );
INV_X1 U993 ( .A(n1327), .ZN(n1298) );
XNOR2_X1 U994 ( .A(G116), .B(n1266), .ZN(G18) );
NAND4_X1 U995 ( .A1(n1321), .A2(n1112), .A3(n1097), .A4(n1324), .ZN(n1266) );
AND2_X1 U996 ( .A1(n1323), .A2(n1328), .ZN(n1097) );
NAND2_X1 U997 ( .A1(n1329), .A2(n1330), .ZN(G15) );
NAND2_X1 U998 ( .A1(G113), .A2(n1331), .ZN(n1330) );
XOR2_X1 U999 ( .A(n1332), .B(KEYINPUT54), .Z(n1329) );
OR2_X1 U1000 ( .A1(n1331), .A2(G113), .ZN(n1332) );
NAND2_X1 U1001 ( .A1(n1333), .A2(n1324), .ZN(n1331) );
XOR2_X1 U1002 ( .A(n1276), .B(KEYINPUT62), .Z(n1333) );
NAND3_X1 U1003 ( .A1(n1112), .A2(n1133), .A3(n1321), .ZN(n1276) );
AND2_X1 U1004 ( .A1(n1114), .A2(n1334), .ZN(n1321) );
NOR2_X1 U1005 ( .A1(n1122), .A2(n1335), .ZN(n1114) );
INV_X1 U1006 ( .A(n1123), .ZN(n1335) );
NOR2_X1 U1007 ( .A1(n1328), .A2(n1323), .ZN(n1133) );
NOR2_X1 U1008 ( .A1(n1327), .A2(n1159), .ZN(n1112) );
XNOR2_X1 U1009 ( .A(G110), .B(n1336), .ZN(G12) );
NAND4_X1 U1010 ( .A1(n1275), .A2(n1113), .A3(n1337), .A4(n1338), .ZN(n1336) );
NOR3_X1 U1011 ( .A1(n1290), .A2(KEYINPUT46), .A3(n1316), .ZN(n1338) );
INV_X1 U1012 ( .A(n1334), .ZN(n1316) );
NAND2_X1 U1013 ( .A1(n1339), .A2(n1119), .ZN(n1334) );
NAND3_X1 U1014 ( .A1(n1319), .A2(n1125), .A3(G952), .ZN(n1119) );
NAND3_X1 U1015 ( .A1(n1190), .A2(n1319), .A3(G902), .ZN(n1339) );
NAND2_X1 U1016 ( .A1(G237), .A2(n1340), .ZN(n1319) );
NOR2_X1 U1017 ( .A1(n1125), .A2(G898), .ZN(n1190) );
NAND2_X1 U1018 ( .A1(n1122), .A2(n1123), .ZN(n1290) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1341), .ZN(n1123) );
XOR2_X1 U1020 ( .A(n1152), .B(n1151), .Z(n1122) );
INV_X1 U1021 ( .A(G469), .ZN(n1151) );
NAND2_X1 U1022 ( .A1(n1342), .A2(n1343), .ZN(n1152) );
XOR2_X1 U1023 ( .A(n1237), .B(n1344), .Z(n1342) );
XOR2_X1 U1024 ( .A(n1345), .B(n1346), .Z(n1344) );
NAND2_X1 U1025 ( .A1(n1347), .A2(n1256), .ZN(n1346) );
NAND3_X1 U1026 ( .A1(n1255), .A2(n1125), .A3(G227), .ZN(n1256) );
INV_X1 U1027 ( .A(n1252), .ZN(n1347) );
NOR2_X1 U1028 ( .A1(n1255), .A2(G227), .ZN(n1252) );
XOR2_X1 U1029 ( .A(G140), .B(n1348), .Z(n1255) );
NAND3_X1 U1030 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1345) );
OR2_X1 U1031 ( .A1(n1186), .A2(n1247), .ZN(n1351) );
NAND2_X1 U1032 ( .A1(KEYINPUT38), .A2(n1352), .ZN(n1350) );
NAND2_X1 U1033 ( .A1(n1353), .A2(n1186), .ZN(n1352) );
XNOR2_X1 U1034 ( .A(KEYINPUT61), .B(n1247), .ZN(n1353) );
NAND2_X1 U1035 ( .A1(n1354), .A2(n1355), .ZN(n1349) );
INV_X1 U1036 ( .A(KEYINPUT38), .ZN(n1355) );
NAND2_X1 U1037 ( .A1(n1356), .A2(n1357), .ZN(n1354) );
OR2_X1 U1038 ( .A1(n1247), .A2(KEYINPUT61), .ZN(n1357) );
NAND3_X1 U1039 ( .A1(n1247), .A2(n1186), .A3(KEYINPUT61), .ZN(n1356) );
NAND3_X1 U1040 ( .A1(n1358), .A2(n1359), .A3(n1360), .ZN(n1186) );
NAND2_X1 U1041 ( .A1(KEYINPUT3), .A2(n1361), .ZN(n1360) );
NAND3_X1 U1042 ( .A1(n1362), .A2(n1363), .A3(n1309), .ZN(n1359) );
INV_X1 U1043 ( .A(KEYINPUT3), .ZN(n1363) );
OR2_X1 U1044 ( .A1(n1309), .A2(n1362), .ZN(n1358) );
NOR2_X1 U1045 ( .A1(KEYINPUT10), .A2(n1361), .ZN(n1362) );
XNOR2_X1 U1046 ( .A(n1364), .B(n1365), .ZN(n1247) );
NOR2_X1 U1047 ( .A1(KEYINPUT27), .A2(n1366), .ZN(n1365) );
XNOR2_X1 U1048 ( .A(G101), .B(G107), .ZN(n1364) );
XNOR2_X1 U1049 ( .A(n1324), .B(KEYINPUT47), .ZN(n1337) );
NOR2_X1 U1050 ( .A1(n1141), .A2(n1140), .ZN(n1324) );
INV_X1 U1051 ( .A(n1156), .ZN(n1140) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1367), .ZN(n1156) );
INV_X1 U1053 ( .A(n1308), .ZN(n1141) );
XNOR2_X1 U1054 ( .A(n1368), .B(n1262), .ZN(n1308) );
AND2_X1 U1055 ( .A1(G210), .A2(n1367), .ZN(n1262) );
NAND2_X1 U1056 ( .A1(n1369), .A2(n1343), .ZN(n1367) );
INV_X1 U1057 ( .A(G237), .ZN(n1369) );
NAND2_X1 U1058 ( .A1(n1370), .A2(n1343), .ZN(n1368) );
XOR2_X1 U1059 ( .A(n1371), .B(n1291), .Z(n1370) );
XOR2_X1 U1060 ( .A(n1372), .B(n1195), .Z(n1291) );
XNOR2_X1 U1061 ( .A(G122), .B(n1348), .ZN(n1195) );
NAND3_X1 U1062 ( .A1(n1373), .A2(n1374), .A3(n1375), .ZN(n1372) );
NAND2_X1 U1063 ( .A1(KEYINPUT45), .A2(n1198), .ZN(n1375) );
NAND3_X1 U1064 ( .A1(n1376), .A2(n1377), .A3(n1199), .ZN(n1374) );
INV_X1 U1065 ( .A(KEYINPUT45), .ZN(n1377) );
OR2_X1 U1066 ( .A1(n1199), .A2(n1376), .ZN(n1373) );
NOR2_X1 U1067 ( .A1(KEYINPUT23), .A2(n1198), .ZN(n1376) );
XNOR2_X1 U1068 ( .A(n1378), .B(n1379), .ZN(n1198) );
XNOR2_X1 U1069 ( .A(KEYINPUT41), .B(n1380), .ZN(n1379) );
INV_X1 U1070 ( .A(G107), .ZN(n1380) );
XNOR2_X1 U1071 ( .A(G101), .B(G104), .ZN(n1378) );
NAND2_X1 U1072 ( .A1(KEYINPUT14), .A2(n1261), .ZN(n1371) );
AND2_X1 U1073 ( .A1(n1381), .A2(n1382), .ZN(n1261) );
NAND3_X1 U1074 ( .A1(n1383), .A2(n1125), .A3(n1384), .ZN(n1382) );
XNOR2_X1 U1075 ( .A(n1385), .B(n1240), .ZN(n1383) );
NAND2_X1 U1076 ( .A1(n1386), .A2(n1387), .ZN(n1381) );
NAND2_X1 U1077 ( .A1(n1384), .A2(n1125), .ZN(n1387) );
XNOR2_X1 U1078 ( .A(KEYINPUT13), .B(G224), .ZN(n1384) );
XNOR2_X1 U1079 ( .A(G125), .B(n1240), .ZN(n1386) );
INV_X1 U1080 ( .A(n1118), .ZN(n1113) );
NAND2_X1 U1081 ( .A1(n1322), .A2(n1323), .ZN(n1118) );
NAND3_X1 U1082 ( .A1(n1388), .A2(n1389), .A3(n1390), .ZN(n1323) );
NAND2_X1 U1083 ( .A1(KEYINPUT32), .A2(n1164), .ZN(n1390) );
NAND3_X1 U1084 ( .A1(n1391), .A2(n1392), .A3(n1225), .ZN(n1389) );
INV_X1 U1085 ( .A(KEYINPUT32), .ZN(n1392) );
OR2_X1 U1086 ( .A1(n1225), .A2(n1391), .ZN(n1388) );
NOR2_X1 U1087 ( .A1(n1164), .A2(KEYINPUT12), .ZN(n1391) );
NOR2_X1 U1088 ( .A1(n1226), .A2(G902), .ZN(n1164) );
XNOR2_X1 U1089 ( .A(n1393), .B(n1394), .ZN(n1226) );
XNOR2_X1 U1090 ( .A(n1366), .B(n1395), .ZN(n1394) );
NOR2_X1 U1091 ( .A1(KEYINPUT58), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1092 ( .A(n1397), .B(n1398), .Z(n1396) );
XNOR2_X1 U1093 ( .A(n1361), .B(n1399), .ZN(n1398) );
INV_X1 U1094 ( .A(n1400), .ZN(n1361) );
XNOR2_X1 U1095 ( .A(G131), .B(n1401), .ZN(n1397) );
NAND2_X1 U1096 ( .A1(G214), .A2(n1402), .ZN(n1401) );
INV_X1 U1097 ( .A(G104), .ZN(n1366) );
XNOR2_X1 U1098 ( .A(G113), .B(G122), .ZN(n1393) );
INV_X1 U1099 ( .A(G475), .ZN(n1225) );
INV_X1 U1100 ( .A(n1328), .ZN(n1322) );
NAND2_X1 U1101 ( .A1(n1403), .A2(n1155), .ZN(n1328) );
OR2_X1 U1102 ( .A1(n1162), .A2(G478), .ZN(n1155) );
NAND2_X1 U1103 ( .A1(G478), .A2(n1162), .ZN(n1403) );
NAND2_X1 U1104 ( .A1(n1220), .A2(n1343), .ZN(n1162) );
XOR2_X1 U1105 ( .A(n1404), .B(n1405), .Z(n1220) );
XNOR2_X1 U1106 ( .A(n1406), .B(n1407), .ZN(n1405) );
XOR2_X1 U1107 ( .A(n1408), .B(n1409), .Z(n1407) );
NOR2_X1 U1108 ( .A1(n1410), .A2(n1411), .ZN(n1409) );
XOR2_X1 U1109 ( .A(n1412), .B(KEYINPUT55), .Z(n1411) );
NAND2_X1 U1110 ( .A1(n1413), .A2(n1414), .ZN(n1412) );
NOR2_X1 U1111 ( .A1(n1413), .A2(n1414), .ZN(n1410) );
XNOR2_X1 U1112 ( .A(G128), .B(n1415), .ZN(n1413) );
XNOR2_X1 U1113 ( .A(KEYINPUT29), .B(n1416), .ZN(n1415) );
INV_X1 U1114 ( .A(G143), .ZN(n1416) );
NAND2_X1 U1115 ( .A1(G217), .A2(n1417), .ZN(n1408) );
XNOR2_X1 U1116 ( .A(G107), .B(n1418), .ZN(n1404) );
XNOR2_X1 U1117 ( .A(KEYINPUT52), .B(n1419), .ZN(n1418) );
INV_X1 U1118 ( .A(G122), .ZN(n1419) );
AND2_X1 U1119 ( .A1(n1159), .A2(n1327), .ZN(n1275) );
XOR2_X1 U1120 ( .A(n1153), .B(n1420), .Z(n1327) );
NOR2_X1 U1121 ( .A1(G472), .A2(KEYINPUT26), .ZN(n1420) );
AND2_X1 U1122 ( .A1(n1421), .A2(n1343), .ZN(n1153) );
XOR2_X1 U1123 ( .A(n1422), .B(n1423), .Z(n1421) );
XOR2_X1 U1124 ( .A(n1424), .B(n1239), .Z(n1423) );
XNOR2_X1 U1125 ( .A(n1425), .B(n1199), .ZN(n1239) );
XOR2_X1 U1126 ( .A(n1426), .B(n1406), .Z(n1199) );
XOR2_X1 U1127 ( .A(G116), .B(KEYINPUT34), .Z(n1406) );
XNOR2_X1 U1128 ( .A(G119), .B(G113), .ZN(n1426) );
XOR2_X1 U1129 ( .A(n1427), .B(KEYINPUT25), .Z(n1425) );
NAND2_X1 U1130 ( .A1(G210), .A2(n1402), .ZN(n1427) );
NOR2_X1 U1131 ( .A1(G953), .A2(G237), .ZN(n1402) );
NAND2_X1 U1132 ( .A1(n1428), .A2(n1429), .ZN(n1424) );
NAND2_X1 U1133 ( .A1(n1237), .A2(n1240), .ZN(n1429) );
XOR2_X1 U1134 ( .A(n1430), .B(KEYINPUT2), .Z(n1428) );
OR2_X1 U1135 ( .A1(n1240), .A2(n1237), .ZN(n1430) );
XNOR2_X1 U1136 ( .A(G131), .B(n1183), .ZN(n1237) );
XNOR2_X1 U1137 ( .A(G137), .B(n1414), .ZN(n1183) );
INV_X1 U1138 ( .A(G134), .ZN(n1414) );
XOR2_X1 U1139 ( .A(n1400), .B(n1431), .Z(n1240) );
NOR2_X1 U1140 ( .A1(G128), .A2(KEYINPUT42), .ZN(n1431) );
XOR2_X1 U1141 ( .A(G143), .B(G146), .Z(n1400) );
XNOR2_X1 U1142 ( .A(KEYINPUT33), .B(n1238), .ZN(n1422) );
INV_X1 U1143 ( .A(G101), .ZN(n1238) );
XOR2_X1 U1144 ( .A(n1432), .B(n1214), .Z(n1159) );
NAND2_X1 U1145 ( .A1(G217), .A2(n1341), .ZN(n1214) );
NAND2_X1 U1146 ( .A1(n1340), .A2(n1343), .ZN(n1341) );
INV_X1 U1147 ( .A(G902), .ZN(n1343) );
XOR2_X1 U1148 ( .A(G234), .B(KEYINPUT60), .Z(n1340) );
OR2_X1 U1149 ( .A1(n1213), .A2(G902), .ZN(n1432) );
XNOR2_X1 U1150 ( .A(n1433), .B(G137), .ZN(n1213) );
XOR2_X1 U1151 ( .A(n1434), .B(n1435), .Z(n1433) );
XOR2_X1 U1152 ( .A(n1436), .B(n1437), .Z(n1435) );
XNOR2_X1 U1153 ( .A(G146), .B(n1309), .ZN(n1437) );
INV_X1 U1154 ( .A(G128), .ZN(n1309) );
XOR2_X1 U1155 ( .A(KEYINPUT51), .B(KEYINPUT48), .Z(n1436) );
XOR2_X1 U1156 ( .A(n1438), .B(n1439), .Z(n1434) );
XOR2_X1 U1157 ( .A(n1348), .B(n1399), .Z(n1439) );
XNOR2_X1 U1158 ( .A(n1385), .B(G140), .ZN(n1399) );
INV_X1 U1159 ( .A(G125), .ZN(n1385) );
XOR2_X1 U1160 ( .A(G110), .B(KEYINPUT22), .Z(n1348) );
XNOR2_X1 U1161 ( .A(n1440), .B(n1326), .ZN(n1438) );
INV_X1 U1162 ( .A(G119), .ZN(n1326) );
NAND2_X1 U1163 ( .A1(G221), .A2(n1417), .ZN(n1440) );
AND2_X1 U1164 ( .A1(G234), .A2(n1125), .ZN(n1417) );
INV_X1 U1165 ( .A(G953), .ZN(n1125) );
endmodule


