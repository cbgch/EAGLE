//Key = 0100000001001111100011111110000000010111011000001100110110001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347;

XNOR2_X1 U745 ( .A(G107), .B(n1025), .ZN(G9) );
NAND3_X1 U746 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(G75) );
NAND2_X1 U747 ( .A1(G952), .A2(n1029), .ZN(n1028) );
NAND3_X1 U748 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
XOR2_X1 U749 ( .A(n1033), .B(KEYINPUT45), .Z(n1032) );
NAND2_X1 U750 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U751 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U752 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U755 ( .A1(n1045), .A2(n1046), .ZN(n1041) );
NAND3_X1 U756 ( .A1(n1044), .A2(n1047), .A3(n1045), .ZN(n1036) );
NAND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1050), .A2(n1040), .ZN(n1049) );
NAND2_X1 U759 ( .A1(n1038), .A2(n1051), .ZN(n1048) );
NAND2_X1 U760 ( .A1(n1034), .A2(n1052), .ZN(n1031) );
NAND2_X1 U761 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U762 ( .A1(n1055), .A2(n1038), .A3(n1056), .ZN(n1054) );
NAND2_X1 U763 ( .A1(n1045), .A2(n1057), .ZN(n1053) );
NAND2_X1 U764 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U765 ( .A1(n1038), .A2(n1060), .ZN(n1059) );
NAND2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND3_X1 U767 ( .A1(n1063), .A2(n1040), .A3(n1064), .ZN(n1062) );
NAND3_X1 U768 ( .A1(n1065), .A2(n1044), .A3(n1066), .ZN(n1061) );
NAND2_X1 U769 ( .A1(n1067), .A2(n1056), .ZN(n1058) );
XOR2_X1 U770 ( .A(n1068), .B(KEYINPUT47), .Z(n1034) );
NAND4_X1 U771 ( .A1(n1069), .A2(n1070), .A3(n1056), .A4(n1071), .ZN(n1026) );
NOR3_X1 U772 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
AND2_X1 U773 ( .A1(n1075), .A2(G478), .ZN(n1074) );
XOR2_X1 U774 ( .A(n1076), .B(n1077), .Z(n1072) );
NOR2_X1 U775 ( .A1(G475), .A2(KEYINPUT46), .ZN(n1077) );
AND2_X1 U776 ( .A1(n1044), .A2(n1040), .ZN(n1056) );
XNOR2_X1 U777 ( .A(n1078), .B(n1079), .ZN(n1070) );
NOR2_X1 U778 ( .A1(G472), .A2(KEYINPUT27), .ZN(n1079) );
XOR2_X1 U779 ( .A(n1080), .B(n1081), .Z(G72) );
NOR2_X1 U780 ( .A1(n1082), .A2(n1027), .ZN(n1081) );
AND2_X1 U781 ( .A1(G227), .A2(G900), .ZN(n1082) );
NAND2_X1 U782 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
NAND2_X1 U783 ( .A1(n1085), .A2(n1027), .ZN(n1084) );
XOR2_X1 U784 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND2_X1 U785 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
XOR2_X1 U786 ( .A(n1090), .B(KEYINPUT21), .Z(n1088) );
NAND3_X1 U787 ( .A1(n1087), .A2(n1091), .A3(G953), .ZN(n1083) );
INV_X1 U788 ( .A(n1092), .ZN(n1091) );
XOR2_X1 U789 ( .A(n1093), .B(n1094), .Z(n1087) );
XOR2_X1 U790 ( .A(n1095), .B(n1096), .Z(G69) );
NOR2_X1 U791 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
AND3_X1 U792 ( .A1(KEYINPUT63), .A2(n1099), .A3(G953), .ZN(n1098) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1099) );
NOR3_X1 U794 ( .A1(G953), .A2(KEYINPUT62), .A3(n1100), .ZN(n1097) );
NAND2_X1 U795 ( .A1(n1101), .A2(n1102), .ZN(n1095) );
NAND2_X1 U796 ( .A1(G953), .A2(n1103), .ZN(n1102) );
XOR2_X1 U797 ( .A(n1104), .B(n1105), .Z(n1101) );
NOR2_X1 U798 ( .A1(n1106), .A2(n1107), .ZN(G66) );
XNOR2_X1 U799 ( .A(n1108), .B(n1109), .ZN(n1107) );
XOR2_X1 U800 ( .A(KEYINPUT17), .B(n1110), .Z(n1109) );
NOR2_X1 U801 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U802 ( .A1(n1106), .A2(n1113), .ZN(G63) );
XOR2_X1 U803 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U804 ( .A1(KEYINPUT1), .A2(n1116), .ZN(n1114) );
NAND2_X1 U805 ( .A1(n1117), .A2(G478), .ZN(n1116) );
NOR3_X1 U806 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(G60) );
AND4_X1 U807 ( .A1(n1121), .A2(KEYINPUT56), .A3(G475), .A4(n1117), .ZN(n1120) );
NOR2_X1 U808 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
NOR3_X1 U809 ( .A1(n1112), .A2(n1123), .A3(n1124), .ZN(n1122) );
NOR2_X1 U810 ( .A1(KEYINPUT56), .A2(n1125), .ZN(n1123) );
AND2_X1 U811 ( .A1(KEYINPUT35), .A2(n1125), .ZN(n1121) );
NOR2_X1 U812 ( .A1(n1126), .A2(n1127), .ZN(n1118) );
XNOR2_X1 U813 ( .A(G952), .B(KEYINPUT15), .ZN(n1126) );
XNOR2_X1 U814 ( .A(G104), .B(n1128), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1106), .A2(n1129), .ZN(G57) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U817 ( .A(n1132), .B(n1133), .Z(n1131) );
AND2_X1 U818 ( .A1(G472), .A2(n1117), .ZN(n1133) );
XNOR2_X1 U819 ( .A(G101), .B(n1134), .ZN(n1130) );
NOR2_X1 U820 ( .A1(KEYINPUT11), .A2(n1135), .ZN(n1134) );
NOR2_X1 U821 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
XOR2_X1 U822 ( .A(n1138), .B(KEYINPUT39), .Z(n1137) );
NAND2_X1 U823 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
XNOR2_X1 U825 ( .A(n1141), .B(KEYINPUT23), .ZN(n1140) );
NOR2_X1 U826 ( .A1(n1106), .A2(n1142), .ZN(G54) );
XOR2_X1 U827 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U828 ( .A(n1145), .B(n1146), .Z(n1144) );
AND2_X1 U829 ( .A1(G469), .A2(n1117), .ZN(n1145) );
XNOR2_X1 U830 ( .A(G101), .B(n1147), .ZN(n1143) );
NOR2_X1 U831 ( .A1(KEYINPUT40), .A2(n1148), .ZN(n1147) );
XNOR2_X1 U832 ( .A(G110), .B(G140), .ZN(n1148) );
NOR2_X1 U833 ( .A1(n1106), .A2(n1149), .ZN(G51) );
XOR2_X1 U834 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U835 ( .A(n1152), .B(n1153), .Z(n1151) );
NOR2_X1 U836 ( .A1(n1154), .A2(n1112), .ZN(n1153) );
INV_X1 U837 ( .A(n1117), .ZN(n1112) );
NOR2_X1 U838 ( .A1(n1155), .A2(n1030), .ZN(n1117) );
AND3_X1 U839 ( .A1(n1100), .A2(n1089), .A3(n1156), .ZN(n1030) );
XOR2_X1 U840 ( .A(n1090), .B(KEYINPUT13), .Z(n1156) );
NAND4_X1 U841 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1090) );
NAND3_X1 U842 ( .A1(n1055), .A2(n1161), .A3(n1162), .ZN(n1157) );
XOR2_X1 U843 ( .A(KEYINPUT10), .B(n1050), .Z(n1161) );
AND4_X1 U844 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1089) );
NOR2_X1 U845 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
OR2_X1 U846 ( .A1(n1169), .A2(KEYINPUT32), .ZN(n1164) );
NAND3_X1 U847 ( .A1(n1170), .A2(n1171), .A3(KEYINPUT32), .ZN(n1163) );
AND4_X1 U848 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1100) );
AND4_X1 U849 ( .A1(n1128), .A2(n1025), .A3(n1176), .A4(n1177), .ZN(n1175) );
NAND3_X1 U850 ( .A1(n1055), .A2(n1038), .A3(n1178), .ZN(n1025) );
NAND3_X1 U851 ( .A1(n1178), .A2(n1038), .A3(n1043), .ZN(n1128) );
AND2_X1 U852 ( .A1(n1179), .A2(n1180), .ZN(n1174) );
NAND3_X1 U853 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1173) );
NAND2_X1 U854 ( .A1(KEYINPUT53), .A2(n1184), .ZN(n1182) );
OR2_X1 U855 ( .A1(n1185), .A2(KEYINPUT53), .ZN(n1181) );
NAND2_X1 U856 ( .A1(n1186), .A2(KEYINPUT20), .ZN(n1152) );
XOR2_X1 U857 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U858 ( .A1(n1189), .A2(KEYINPUT9), .ZN(n1187) );
XOR2_X1 U859 ( .A(n1190), .B(KEYINPUT7), .Z(n1189) );
NOR2_X1 U860 ( .A1(n1127), .A2(G952), .ZN(n1106) );
XOR2_X1 U861 ( .A(G953), .B(KEYINPUT37), .Z(n1127) );
XNOR2_X1 U862 ( .A(G146), .B(n1165), .ZN(G48) );
NAND2_X1 U863 ( .A1(n1191), .A2(n1043), .ZN(n1165) );
NAND2_X1 U864 ( .A1(n1192), .A2(n1193), .ZN(G45) );
OR2_X1 U865 ( .A1(n1169), .A2(G143), .ZN(n1193) );
XOR2_X1 U866 ( .A(n1194), .B(KEYINPUT8), .Z(n1192) );
NAND2_X1 U867 ( .A1(G143), .A2(n1169), .ZN(n1194) );
NAND2_X1 U868 ( .A1(n1171), .A2(n1195), .ZN(n1169) );
AND3_X1 U869 ( .A1(n1050), .A2(n1046), .A3(n1196), .ZN(n1171) );
NOR3_X1 U870 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
XOR2_X1 U871 ( .A(n1168), .B(n1200), .Z(G42) );
XNOR2_X1 U872 ( .A(KEYINPUT61), .B(n1201), .ZN(n1200) );
AND3_X1 U873 ( .A1(n1067), .A2(n1043), .A3(n1162), .ZN(n1168) );
XNOR2_X1 U874 ( .A(n1202), .B(n1167), .ZN(G39) );
AND2_X1 U875 ( .A1(n1162), .A2(n1183), .ZN(n1167) );
XNOR2_X1 U876 ( .A(G134), .B(n1203), .ZN(G36) );
NAND2_X1 U877 ( .A1(n1204), .A2(n1055), .ZN(n1203) );
XNOR2_X1 U878 ( .A(G131), .B(n1158), .ZN(G33) );
NAND2_X1 U879 ( .A1(n1204), .A2(n1043), .ZN(n1158) );
AND2_X1 U880 ( .A1(n1162), .A2(n1050), .ZN(n1204) );
AND3_X1 U881 ( .A1(n1046), .A2(n1195), .A3(n1040), .ZN(n1162) );
NOR2_X1 U882 ( .A1(n1205), .A2(n1066), .ZN(n1040) );
XNOR2_X1 U883 ( .A(G128), .B(n1159), .ZN(G30) );
NAND2_X1 U884 ( .A1(n1191), .A2(n1055), .ZN(n1159) );
AND3_X1 U885 ( .A1(n1046), .A2(n1051), .A3(n1206), .ZN(n1191) );
NOR3_X1 U886 ( .A1(n1069), .A2(n1170), .A3(n1207), .ZN(n1206) );
XNOR2_X1 U887 ( .A(G101), .B(n1180), .ZN(G3) );
NAND3_X1 U888 ( .A1(n1050), .A2(n1178), .A3(n1045), .ZN(n1180) );
XOR2_X1 U889 ( .A(n1160), .B(n1208), .Z(G27) );
NAND2_X1 U890 ( .A1(KEYINPUT38), .A2(G125), .ZN(n1208) );
NAND4_X1 U891 ( .A1(n1067), .A2(n1043), .A3(n1209), .A4(n1044), .ZN(n1160) );
NOR2_X1 U892 ( .A1(n1170), .A2(n1197), .ZN(n1209) );
INV_X1 U893 ( .A(n1195), .ZN(n1170) );
NAND2_X1 U894 ( .A1(n1210), .A2(n1211), .ZN(n1195) );
NAND2_X1 U895 ( .A1(n1212), .A2(n1092), .ZN(n1210) );
XOR2_X1 U896 ( .A(G900), .B(KEYINPUT26), .Z(n1092) );
NAND2_X1 U897 ( .A1(n1213), .A2(n1214), .ZN(G24) );
NAND3_X1 U898 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
NAND2_X1 U899 ( .A1(n1218), .A2(n1219), .ZN(n1216) );
NAND2_X1 U900 ( .A1(G122), .A2(n1220), .ZN(n1215) );
NAND3_X1 U901 ( .A1(n1221), .A2(n1222), .A3(n1219), .ZN(n1220) );
INV_X1 U902 ( .A(KEYINPUT29), .ZN(n1219) );
OR2_X1 U903 ( .A1(n1172), .A2(KEYINPUT3), .ZN(n1222) );
NAND2_X1 U904 ( .A1(n1223), .A2(n1224), .ZN(n1172) );
NAND3_X1 U905 ( .A1(n1185), .A2(n1223), .A3(KEYINPUT3), .ZN(n1221) );
AND3_X1 U906 ( .A1(n1225), .A2(n1197), .A3(n1044), .ZN(n1185) );
INV_X1 U907 ( .A(n1051), .ZN(n1197) );
NAND3_X1 U908 ( .A1(n1223), .A2(n1044), .A3(n1226), .ZN(n1213) );
NOR3_X1 U909 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1226) );
NOR2_X1 U910 ( .A1(n1230), .A2(n1218), .ZN(n1229) );
NOR2_X1 U911 ( .A1(KEYINPUT29), .A2(n1217), .ZN(n1230) );
INV_X1 U912 ( .A(KEYINPUT44), .ZN(n1217) );
INV_X1 U913 ( .A(n1225), .ZN(n1228) );
XNOR2_X1 U914 ( .A(n1051), .B(KEYINPUT3), .ZN(n1227) );
AND3_X1 U915 ( .A1(n1231), .A2(n1232), .A3(n1038), .ZN(n1223) );
NOR2_X1 U916 ( .A1(n1233), .A2(n1234), .ZN(n1038) );
XNOR2_X1 U917 ( .A(G119), .B(n1235), .ZN(G21) );
NAND3_X1 U918 ( .A1(n1183), .A2(n1224), .A3(KEYINPUT22), .ZN(n1235) );
AND3_X1 U919 ( .A1(n1234), .A2(n1233), .A3(n1045), .ZN(n1183) );
XNOR2_X1 U920 ( .A(G116), .B(n1179), .ZN(G18) );
NAND3_X1 U921 ( .A1(n1224), .A2(n1055), .A3(n1050), .ZN(n1179) );
AND2_X1 U922 ( .A1(n1236), .A2(n1232), .ZN(n1055) );
NAND2_X1 U923 ( .A1(n1237), .A2(n1238), .ZN(G15) );
NAND2_X1 U924 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NAND2_X1 U925 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
NAND2_X1 U926 ( .A1(KEYINPUT50), .A2(n1177), .ZN(n1242) );
NAND2_X1 U927 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
INV_X1 U928 ( .A(KEYINPUT50), .ZN(n1244) );
OR2_X1 U929 ( .A1(n1243), .A2(n1240), .ZN(n1237) );
NAND2_X1 U930 ( .A1(KEYINPUT41), .A2(n1177), .ZN(n1243) );
NAND3_X1 U931 ( .A1(n1050), .A2(n1224), .A3(n1043), .ZN(n1177) );
NOR2_X1 U932 ( .A1(n1232), .A2(n1199), .ZN(n1043) );
INV_X1 U933 ( .A(n1198), .ZN(n1232) );
INV_X1 U934 ( .A(n1184), .ZN(n1224) );
NAND3_X1 U935 ( .A1(n1051), .A2(n1225), .A3(n1044), .ZN(n1184) );
NOR2_X1 U936 ( .A1(n1245), .A2(n1064), .ZN(n1044) );
NOR2_X1 U937 ( .A1(n1234), .A2(n1207), .ZN(n1050) );
INV_X1 U938 ( .A(n1233), .ZN(n1207) );
XNOR2_X1 U939 ( .A(G110), .B(n1176), .ZN(G12) );
NAND3_X1 U940 ( .A1(n1045), .A2(n1178), .A3(n1067), .ZN(n1176) );
NOR2_X1 U941 ( .A1(n1233), .A2(n1069), .ZN(n1067) );
INV_X1 U942 ( .A(n1234), .ZN(n1069) );
XOR2_X1 U943 ( .A(n1246), .B(n1111), .Z(n1234) );
NAND2_X1 U944 ( .A1(G217), .A2(n1247), .ZN(n1111) );
NAND2_X1 U945 ( .A1(n1108), .A2(n1155), .ZN(n1246) );
XNOR2_X1 U946 ( .A(n1248), .B(n1249), .ZN(n1108) );
XOR2_X1 U947 ( .A(n1250), .B(n1251), .Z(n1249) );
XOR2_X1 U948 ( .A(n1252), .B(n1253), .Z(n1251) );
NOR2_X1 U949 ( .A1(KEYINPUT28), .A2(n1202), .ZN(n1253) );
NAND2_X1 U950 ( .A1(n1254), .A2(G221), .ZN(n1252) );
XNOR2_X1 U951 ( .A(G119), .B(KEYINPUT34), .ZN(n1250) );
XNOR2_X1 U952 ( .A(n1255), .B(n1256), .ZN(n1248) );
XOR2_X1 U953 ( .A(n1257), .B(n1094), .Z(n1256) );
NOR2_X1 U954 ( .A1(KEYINPUT51), .A2(n1258), .ZN(n1257) );
NAND2_X1 U955 ( .A1(n1259), .A2(n1260), .ZN(n1233) );
NAND2_X1 U956 ( .A1(G472), .A2(n1078), .ZN(n1260) );
XOR2_X1 U957 ( .A(n1261), .B(KEYINPUT58), .Z(n1259) );
OR2_X1 U958 ( .A1(n1078), .A2(G472), .ZN(n1261) );
NAND2_X1 U959 ( .A1(n1262), .A2(n1155), .ZN(n1078) );
XOR2_X1 U960 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U961 ( .A(n1265), .B(n1132), .ZN(n1264) );
NAND2_X1 U962 ( .A1(n1266), .A2(G210), .ZN(n1132) );
NAND2_X1 U963 ( .A1(n1267), .A2(KEYINPUT48), .ZN(n1265) );
XOR2_X1 U964 ( .A(n1268), .B(KEYINPUT18), .Z(n1267) );
NAND3_X1 U965 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1268) );
NAND2_X1 U966 ( .A1(n1139), .A2(n1272), .ZN(n1271) );
INV_X1 U967 ( .A(KEYINPUT16), .ZN(n1272) );
NAND3_X1 U968 ( .A1(KEYINPUT16), .A2(n1273), .A3(n1141), .ZN(n1270) );
OR2_X1 U969 ( .A1(n1141), .A2(n1273), .ZN(n1269) );
NOR2_X1 U970 ( .A1(KEYINPUT59), .A2(n1139), .ZN(n1273) );
XOR2_X1 U971 ( .A(n1274), .B(n1275), .Z(n1139) );
XNOR2_X1 U972 ( .A(G119), .B(G113), .ZN(n1274) );
XNOR2_X1 U973 ( .A(n1190), .B(n1276), .ZN(n1141) );
NAND2_X1 U974 ( .A1(KEYINPUT25), .A2(G101), .ZN(n1263) );
AND3_X1 U975 ( .A1(n1051), .A2(n1225), .A3(n1046), .ZN(n1178) );
NOR2_X1 U976 ( .A1(n1063), .A2(n1064), .ZN(n1046) );
AND2_X1 U977 ( .A1(G221), .A2(n1247), .ZN(n1064) );
NAND2_X1 U978 ( .A1(G234), .A2(n1155), .ZN(n1247) );
INV_X1 U979 ( .A(n1245), .ZN(n1063) );
XNOR2_X1 U980 ( .A(n1277), .B(G469), .ZN(n1245) );
NAND2_X1 U981 ( .A1(n1278), .A2(n1155), .ZN(n1277) );
XNOR2_X1 U982 ( .A(n1146), .B(n1279), .ZN(n1278) );
XNOR2_X1 U983 ( .A(G140), .B(n1280), .ZN(n1279) );
XNOR2_X1 U984 ( .A(n1281), .B(n1282), .ZN(n1146) );
XNOR2_X1 U985 ( .A(n1283), .B(G104), .ZN(n1282) );
XOR2_X1 U986 ( .A(n1093), .B(n1284), .Z(n1281) );
NOR2_X1 U987 ( .A1(G953), .A2(n1285), .ZN(n1284) );
XOR2_X1 U988 ( .A(KEYINPUT52), .B(G227), .Z(n1285) );
NAND2_X1 U989 ( .A1(n1286), .A2(n1287), .ZN(n1093) );
NAND2_X1 U990 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
INV_X1 U991 ( .A(G128), .ZN(n1289) );
XNOR2_X1 U992 ( .A(n1290), .B(KEYINPUT0), .ZN(n1288) );
NAND2_X1 U993 ( .A1(n1291), .A2(G128), .ZN(n1286) );
XNOR2_X1 U994 ( .A(KEYINPUT36), .B(n1292), .ZN(n1291) );
INV_X1 U995 ( .A(n1290), .ZN(n1292) );
XNOR2_X1 U996 ( .A(n1293), .B(n1294), .ZN(n1290) );
XOR2_X1 U997 ( .A(KEYINPUT57), .B(G146), .Z(n1294) );
XOR2_X1 U998 ( .A(n1276), .B(G143), .Z(n1293) );
XNOR2_X1 U999 ( .A(G131), .B(n1295), .ZN(n1276) );
XNOR2_X1 U1000 ( .A(n1202), .B(G134), .ZN(n1295) );
INV_X1 U1001 ( .A(G137), .ZN(n1202) );
NAND2_X1 U1002 ( .A1(n1211), .A2(n1296), .ZN(n1225) );
NAND2_X1 U1003 ( .A1(n1212), .A2(n1103), .ZN(n1296) );
INV_X1 U1004 ( .A(G898), .ZN(n1103) );
AND3_X1 U1005 ( .A1(G902), .A2(n1068), .A3(G953), .ZN(n1212) );
NAND3_X1 U1006 ( .A1(n1297), .A2(n1027), .A3(G952), .ZN(n1211) );
XNOR2_X1 U1007 ( .A(KEYINPUT55), .B(n1068), .ZN(n1297) );
NAND2_X1 U1008 ( .A1(G237), .A2(G234), .ZN(n1068) );
NOR2_X1 U1009 ( .A1(n1065), .A2(n1066), .ZN(n1051) );
AND2_X1 U1010 ( .A1(G214), .A2(n1298), .ZN(n1066) );
INV_X1 U1011 ( .A(n1205), .ZN(n1065) );
XOR2_X1 U1012 ( .A(n1299), .B(n1154), .Z(n1205) );
NAND2_X1 U1013 ( .A1(G210), .A2(n1298), .ZN(n1154) );
NAND2_X1 U1014 ( .A1(n1300), .A2(n1155), .ZN(n1298) );
INV_X1 U1015 ( .A(G237), .ZN(n1300) );
NAND2_X1 U1016 ( .A1(n1301), .A2(n1155), .ZN(n1299) );
XOR2_X1 U1017 ( .A(n1150), .B(n1302), .Z(n1301) );
XNOR2_X1 U1018 ( .A(n1190), .B(n1188), .ZN(n1302) );
XOR2_X1 U1019 ( .A(G125), .B(n1303), .Z(n1188) );
AND2_X1 U1020 ( .A1(n1027), .A2(G224), .ZN(n1303) );
XNOR2_X1 U1021 ( .A(n1304), .B(n1305), .ZN(n1190) );
INV_X1 U1022 ( .A(n1255), .ZN(n1305) );
XOR2_X1 U1023 ( .A(G128), .B(G146), .Z(n1255) );
NAND2_X1 U1024 ( .A1(KEYINPUT42), .A2(G143), .ZN(n1304) );
XOR2_X1 U1025 ( .A(n1306), .B(n1105), .Z(n1150) );
XOR2_X1 U1026 ( .A(n1280), .B(n1307), .Z(n1105) );
XNOR2_X1 U1027 ( .A(n1218), .B(n1308), .ZN(n1307) );
NOR4_X1 U1028 ( .A1(n1309), .A2(n1310), .A3(KEYINPUT54), .A4(n1311), .ZN(n1308) );
NOR2_X1 U1029 ( .A1(KEYINPUT12), .A2(n1312), .ZN(n1311) );
NOR2_X1 U1030 ( .A1(n1313), .A2(n1283), .ZN(n1310) );
AND2_X1 U1031 ( .A1(n1312), .A2(KEYINPUT49), .ZN(n1313) );
AND4_X1 U1032 ( .A1(n1283), .A2(KEYINPUT12), .A3(n1312), .A4(KEYINPUT49), .ZN(n1309) );
INV_X1 U1033 ( .A(G104), .ZN(n1312) );
INV_X1 U1034 ( .A(G107), .ZN(n1283) );
XNOR2_X1 U1035 ( .A(G101), .B(n1258), .ZN(n1280) );
INV_X1 U1036 ( .A(G110), .ZN(n1258) );
NAND2_X1 U1037 ( .A1(KEYINPUT14), .A2(n1104), .ZN(n1306) );
NAND2_X1 U1038 ( .A1(n1314), .A2(n1315), .ZN(n1104) );
NAND2_X1 U1039 ( .A1(n1316), .A2(n1240), .ZN(n1315) );
XOR2_X1 U1040 ( .A(KEYINPUT24), .B(n1317), .Z(n1314) );
NOR2_X1 U1041 ( .A1(n1316), .A2(n1240), .ZN(n1317) );
INV_X1 U1042 ( .A(G113), .ZN(n1240) );
XNOR2_X1 U1043 ( .A(n1318), .B(n1319), .ZN(n1316) );
NOR2_X1 U1044 ( .A1(KEYINPUT30), .A2(n1275), .ZN(n1319) );
XNOR2_X1 U1045 ( .A(n1320), .B(KEYINPUT6), .ZN(n1275) );
INV_X1 U1046 ( .A(G119), .ZN(n1318) );
AND2_X1 U1047 ( .A1(n1198), .A2(n1321), .ZN(n1045) );
XOR2_X1 U1048 ( .A(KEYINPUT33), .B(n1236), .Z(n1321) );
XNOR2_X1 U1049 ( .A(n1199), .B(KEYINPUT60), .ZN(n1236) );
INV_X1 U1050 ( .A(n1231), .ZN(n1199) );
XOR2_X1 U1051 ( .A(n1076), .B(n1124), .Z(n1231) );
INV_X1 U1052 ( .A(G475), .ZN(n1124) );
NAND2_X1 U1053 ( .A1(n1125), .A2(n1155), .ZN(n1076) );
INV_X1 U1054 ( .A(G902), .ZN(n1155) );
XOR2_X1 U1055 ( .A(n1322), .B(n1323), .Z(n1125) );
XNOR2_X1 U1056 ( .A(n1094), .B(n1324), .ZN(n1323) );
XOR2_X1 U1057 ( .A(n1325), .B(n1326), .Z(n1324) );
NOR2_X1 U1058 ( .A1(G146), .A2(KEYINPUT4), .ZN(n1326) );
NAND2_X1 U1059 ( .A1(n1266), .A2(G214), .ZN(n1325) );
NOR2_X1 U1060 ( .A1(G953), .A2(G237), .ZN(n1266) );
XNOR2_X1 U1061 ( .A(G125), .B(n1201), .ZN(n1094) );
INV_X1 U1062 ( .A(G140), .ZN(n1201) );
XOR2_X1 U1063 ( .A(n1327), .B(n1328), .Z(n1322) );
XOR2_X1 U1064 ( .A(G143), .B(G131), .Z(n1328) );
NAND3_X1 U1065 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1327) );
NAND2_X1 U1066 ( .A1(KEYINPUT43), .A2(G104), .ZN(n1331) );
OR3_X1 U1067 ( .A1(G104), .A2(KEYINPUT43), .A3(n1332), .ZN(n1330) );
NAND2_X1 U1068 ( .A1(n1332), .A2(n1333), .ZN(n1329) );
NAND2_X1 U1069 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
INV_X1 U1070 ( .A(KEYINPUT43), .ZN(n1335) );
XNOR2_X1 U1071 ( .A(G104), .B(KEYINPUT31), .ZN(n1334) );
XNOR2_X1 U1072 ( .A(G113), .B(n1218), .ZN(n1332) );
NOR2_X1 U1073 ( .A1(n1336), .A2(n1073), .ZN(n1198) );
NOR2_X1 U1074 ( .A1(n1075), .A2(G478), .ZN(n1073) );
AND2_X1 U1075 ( .A1(n1337), .A2(n1075), .ZN(n1336) );
OR2_X1 U1076 ( .A1(n1115), .A2(G902), .ZN(n1075) );
XNOR2_X1 U1077 ( .A(n1338), .B(n1339), .ZN(n1115) );
XOR2_X1 U1078 ( .A(n1340), .B(n1341), .Z(n1339) );
NAND2_X1 U1079 ( .A1(G217), .A2(n1254), .ZN(n1341) );
AND2_X1 U1080 ( .A1(G234), .A2(n1027), .ZN(n1254) );
INV_X1 U1081 ( .A(G953), .ZN(n1027) );
NAND2_X1 U1082 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1083 ( .A1(G122), .A2(n1320), .ZN(n1343) );
INV_X1 U1084 ( .A(G116), .ZN(n1320) );
XOR2_X1 U1085 ( .A(n1344), .B(KEYINPUT19), .Z(n1342) );
NAND2_X1 U1086 ( .A1(G116), .A2(n1218), .ZN(n1344) );
INV_X1 U1087 ( .A(G122), .ZN(n1218) );
XOR2_X1 U1088 ( .A(n1345), .B(n1346), .Z(n1338) );
NOR2_X1 U1089 ( .A1(KEYINPUT5), .A2(n1347), .ZN(n1346) );
XNOR2_X1 U1090 ( .A(G128), .B(G143), .ZN(n1347) );
XNOR2_X1 U1091 ( .A(G134), .B(G107), .ZN(n1345) );
XOR2_X1 U1092 ( .A(KEYINPUT2), .B(G478), .Z(n1337) );
endmodule


