//Key = 0011001001011100011000010011111101101110000111011000000110000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339;

XNOR2_X1 U744 ( .A(G107), .B(n1014), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR4_X1 U746 ( .A1(G953), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1016) );
INV_X1 U747 ( .A(n1020), .ZN(n1019) );
NOR3_X1 U748 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1018) );
INV_X1 U749 ( .A(n1024), .ZN(n1023) );
NOR2_X1 U750 ( .A1(n1025), .A2(n1026), .ZN(n1022) );
NOR2_X1 U751 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U752 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U753 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U754 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U755 ( .A1(n1035), .A2(n1036), .ZN(n1029) );
NOR2_X1 U756 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U757 ( .A1(n1036), .A2(n1039), .A3(n1032), .ZN(n1025) );
NOR2_X1 U758 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
XOR2_X1 U759 ( .A(n1042), .B(KEYINPUT55), .Z(n1041) );
NAND2_X1 U760 ( .A1(KEYINPUT48), .A2(n1043), .ZN(n1042) );
NOR4_X1 U761 ( .A1(n1044), .A2(n1032), .A3(n1036), .A4(n1028), .ZN(n1017) );
NOR2_X1 U762 ( .A1(n1045), .A2(n1024), .ZN(n1044) );
NOR2_X1 U763 ( .A1(n1046), .A2(n1021), .ZN(n1045) );
NOR2_X1 U764 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR3_X1 U765 ( .A1(n1049), .A2(G953), .A3(G952), .ZN(n1015) );
XOR2_X1 U766 ( .A(n1050), .B(n1051), .Z(G72) );
NOR2_X1 U767 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XNOR2_X1 U768 ( .A(G953), .B(KEYINPUT20), .ZN(n1053) );
AND2_X1 U769 ( .A1(G227), .A2(G900), .ZN(n1052) );
NAND2_X1 U770 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
NAND2_X1 U771 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XOR2_X1 U772 ( .A(n1058), .B(n1059), .Z(n1056) );
NAND3_X1 U773 ( .A1(G900), .A2(n1059), .A3(G953), .ZN(n1054) );
XNOR2_X1 U774 ( .A(n1060), .B(n1061), .ZN(n1059) );
NAND2_X1 U775 ( .A1(n1062), .A2(KEYINPUT34), .ZN(n1060) );
XOR2_X1 U776 ( .A(n1063), .B(n1064), .Z(n1062) );
XNOR2_X1 U777 ( .A(n1065), .B(G134), .ZN(n1064) );
XOR2_X1 U778 ( .A(n1066), .B(G131), .Z(n1063) );
NAND2_X1 U779 ( .A1(n1067), .A2(n1068), .ZN(G69) );
NAND2_X1 U780 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U781 ( .A1(n1071), .A2(n1072), .ZN(n1067) );
NAND2_X1 U782 ( .A1(n1073), .A2(n1070), .ZN(n1072) );
NAND2_X1 U783 ( .A1(G953), .A2(n1074), .ZN(n1070) );
INV_X1 U784 ( .A(n1075), .ZN(n1073) );
INV_X1 U785 ( .A(n1069), .ZN(n1071) );
XNOR2_X1 U786 ( .A(n1076), .B(n1077), .ZN(n1069) );
NOR2_X1 U787 ( .A1(n1075), .A2(n1078), .ZN(n1077) );
XNOR2_X1 U788 ( .A(n1079), .B(n1080), .ZN(n1078) );
NAND3_X1 U789 ( .A1(n1081), .A2(n1057), .A3(KEYINPUT18), .ZN(n1076) );
NOR2_X1 U790 ( .A1(n1082), .A2(n1083), .ZN(G66) );
XOR2_X1 U791 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U792 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U793 ( .A1(n1088), .A2(n1089), .ZN(G63) );
XOR2_X1 U794 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U795 ( .A1(n1086), .A2(n1092), .ZN(n1090) );
XOR2_X1 U796 ( .A(KEYINPUT10), .B(G478), .Z(n1092) );
NOR2_X1 U797 ( .A1(G952), .A2(n1093), .ZN(n1088) );
XNOR2_X1 U798 ( .A(KEYINPUT3), .B(n1057), .ZN(n1093) );
NOR2_X1 U799 ( .A1(n1082), .A2(n1094), .ZN(G60) );
XOR2_X1 U800 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND3_X1 U801 ( .A1(n1097), .A2(n1098), .A3(G475), .ZN(n1095) );
OR2_X1 U802 ( .A1(n1099), .A2(n1086), .ZN(n1098) );
NAND2_X1 U803 ( .A1(n1100), .A2(n1099), .ZN(n1097) );
INV_X1 U804 ( .A(KEYINPUT13), .ZN(n1099) );
NAND2_X1 U805 ( .A1(n1020), .A2(G902), .ZN(n1100) );
XNOR2_X1 U806 ( .A(n1101), .B(n1102), .ZN(G6) );
NAND2_X1 U807 ( .A1(KEYINPUT31), .A2(G104), .ZN(n1102) );
NOR2_X1 U808 ( .A1(n1103), .A2(n1104), .ZN(G57) );
XOR2_X1 U809 ( .A(n1105), .B(n1106), .Z(n1104) );
XNOR2_X1 U810 ( .A(n1107), .B(n1108), .ZN(n1106) );
XNOR2_X1 U811 ( .A(n1109), .B(n1110), .ZN(n1105) );
NAND2_X1 U812 ( .A1(n1086), .A2(G472), .ZN(n1109) );
NOR2_X1 U813 ( .A1(G952), .A2(n1111), .ZN(n1103) );
XNOR2_X1 U814 ( .A(G953), .B(KEYINPUT21), .ZN(n1111) );
NOR2_X1 U815 ( .A1(n1082), .A2(n1112), .ZN(G54) );
XOR2_X1 U816 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U817 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U818 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND2_X1 U819 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NAND2_X1 U820 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XNOR2_X1 U821 ( .A(KEYINPUT0), .B(n1123), .ZN(n1122) );
INV_X1 U822 ( .A(n1124), .ZN(n1119) );
NAND2_X1 U823 ( .A1(n1125), .A2(n1126), .ZN(n1115) );
NAND3_X1 U824 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
NAND2_X1 U825 ( .A1(KEYINPUT0), .A2(n1124), .ZN(n1129) );
NOR2_X1 U826 ( .A1(n1130), .A2(n1121), .ZN(n1124) );
OR3_X1 U827 ( .A1(n1121), .A2(KEYINPUT0), .A3(n1123), .ZN(n1128) );
NAND2_X1 U828 ( .A1(n1121), .A2(n1123), .ZN(n1127) );
INV_X1 U829 ( .A(n1130), .ZN(n1123) );
XNOR2_X1 U830 ( .A(n1131), .B(KEYINPUT56), .ZN(n1121) );
INV_X1 U831 ( .A(n1118), .ZN(n1125) );
NAND2_X1 U832 ( .A1(KEYINPUT36), .A2(n1132), .ZN(n1118) );
NAND2_X1 U833 ( .A1(n1086), .A2(G469), .ZN(n1113) );
NOR2_X1 U834 ( .A1(n1082), .A2(n1133), .ZN(G51) );
XOR2_X1 U835 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U836 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U837 ( .A1(KEYINPUT44), .A2(n1138), .ZN(n1137) );
NAND3_X1 U838 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
NAND2_X1 U839 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U840 ( .A1(KEYINPUT9), .A2(n1144), .ZN(n1143) );
XNOR2_X1 U841 ( .A(KEYINPUT39), .B(n1145), .ZN(n1144) );
XNOR2_X1 U842 ( .A(n1108), .B(n1146), .ZN(n1142) );
OR2_X1 U843 ( .A1(n1147), .A2(KEYINPUT9), .ZN(n1140) );
NAND3_X1 U844 ( .A1(n1147), .A2(n1148), .A3(KEYINPUT9), .ZN(n1139) );
XNOR2_X1 U845 ( .A(n1146), .B(n1149), .ZN(n1148) );
AND2_X1 U846 ( .A1(KEYINPUT6), .A2(n1150), .ZN(n1146) );
NAND2_X1 U847 ( .A1(n1151), .A2(n1086), .ZN(n1136) );
NOR2_X1 U848 ( .A1(n1152), .A2(n1020), .ZN(n1086) );
NOR2_X1 U849 ( .A1(n1081), .A2(n1058), .ZN(n1020) );
NAND4_X1 U850 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1058) );
NOR4_X1 U851 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
NOR2_X1 U852 ( .A1(KEYINPUT58), .A2(n1161), .ZN(n1160) );
NOR2_X1 U853 ( .A1(n1162), .A2(n1163), .ZN(n1159) );
NOR2_X1 U854 ( .A1(n1164), .A2(n1165), .ZN(n1158) );
AND3_X1 U855 ( .A1(n1166), .A2(n1037), .A3(n1047), .ZN(n1157) );
AND3_X1 U856 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1155) );
NAND3_X1 U857 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(n1153) );
NAND2_X1 U858 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND3_X1 U859 ( .A1(n1049), .A2(n1163), .A3(n1175), .ZN(n1174) );
INV_X1 U860 ( .A(KEYINPUT62), .ZN(n1163) );
NAND4_X1 U861 ( .A1(KEYINPUT58), .A2(n1176), .A3(n1037), .A4(n1040), .ZN(n1173) );
NAND4_X1 U862 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1081) );
NOR4_X1 U863 ( .A1(n1181), .A2(n1101), .A3(n1182), .A4(n1183), .ZN(n1180) );
NOR2_X1 U864 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
INV_X1 U865 ( .A(KEYINPUT12), .ZN(n1185) );
NOR4_X1 U866 ( .A1(n1186), .A2(n1187), .A3(n1164), .A4(n1036), .ZN(n1182) );
AND2_X1 U867 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U868 ( .A1(n1190), .A2(n1188), .ZN(n1186) );
NOR3_X1 U869 ( .A1(n1191), .A2(KEYINPUT12), .A3(n1032), .ZN(n1190) );
AND3_X1 U870 ( .A1(n1192), .A2(n1024), .A3(n1038), .ZN(n1101) );
INV_X1 U871 ( .A(n1193), .ZN(n1181) );
AND2_X1 U872 ( .A1(n1014), .A2(n1194), .ZN(n1179) );
NAND3_X1 U873 ( .A1(n1024), .A2(n1037), .A3(n1192), .ZN(n1014) );
XOR2_X1 U874 ( .A(n1195), .B(KEYINPUT37), .Z(n1151) );
NOR2_X1 U875 ( .A1(n1057), .A2(G952), .ZN(n1082) );
XOR2_X1 U876 ( .A(G146), .B(n1196), .Z(G48) );
NOR2_X1 U877 ( .A1(n1197), .A2(n1164), .ZN(n1196) );
XOR2_X1 U878 ( .A(n1165), .B(KEYINPUT4), .Z(n1197) );
NAND3_X1 U879 ( .A1(n1176), .A2(n1038), .A3(n1198), .ZN(n1165) );
XOR2_X1 U880 ( .A(n1154), .B(n1199), .Z(G45) );
NAND2_X1 U881 ( .A1(KEYINPUT61), .A2(G143), .ZN(n1199) );
NAND3_X1 U882 ( .A1(n1198), .A2(n1047), .A3(n1200), .ZN(n1154) );
NOR3_X1 U883 ( .A1(n1164), .A2(n1201), .A3(n1202), .ZN(n1200) );
INV_X1 U884 ( .A(n1040), .ZN(n1164) );
XNOR2_X1 U885 ( .A(G140), .B(n1167), .ZN(G42) );
NAND2_X1 U886 ( .A1(n1166), .A2(n1203), .ZN(n1167) );
XNOR2_X1 U887 ( .A(G137), .B(n1169), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1176), .A2(n1204), .A3(n1166), .ZN(n1169) );
NAND2_X1 U889 ( .A1(n1205), .A2(n1206), .ZN(G36) );
NAND3_X1 U890 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1206) );
NAND2_X1 U891 ( .A1(n1210), .A2(G134), .ZN(n1205) );
NAND2_X1 U892 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND2_X1 U893 ( .A1(KEYINPUT50), .A2(n1207), .ZN(n1212) );
NAND2_X1 U894 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
INV_X1 U895 ( .A(KEYINPUT50), .ZN(n1214) );
NAND2_X1 U896 ( .A1(n1207), .A2(n1208), .ZN(n1213) );
INV_X1 U897 ( .A(KEYINPUT57), .ZN(n1208) );
AND3_X1 U898 ( .A1(n1047), .A2(n1215), .A3(n1166), .ZN(n1207) );
XOR2_X1 U899 ( .A(KEYINPUT53), .B(n1037), .Z(n1215) );
XOR2_X1 U900 ( .A(n1162), .B(n1216), .Z(G33) );
NAND2_X1 U901 ( .A1(KEYINPUT11), .A2(n1217), .ZN(n1216) );
XOR2_X1 U902 ( .A(KEYINPUT46), .B(G131), .Z(n1217) );
NAND2_X1 U903 ( .A1(n1175), .A2(n1166), .ZN(n1162) );
AND2_X1 U904 ( .A1(n1049), .A2(n1198), .ZN(n1166) );
INV_X1 U905 ( .A(n1028), .ZN(n1049) );
NAND2_X1 U906 ( .A1(n1043), .A2(n1218), .ZN(n1028) );
INV_X1 U907 ( .A(n1189), .ZN(n1175) );
XNOR2_X1 U908 ( .A(G128), .B(n1161), .ZN(G30) );
NAND4_X1 U909 ( .A1(n1198), .A2(n1176), .A3(n1037), .A4(n1040), .ZN(n1161) );
AND2_X1 U910 ( .A1(n1033), .A2(n1170), .ZN(n1198) );
XOR2_X1 U911 ( .A(n1219), .B(G101), .Z(G3) );
NAND2_X1 U912 ( .A1(KEYINPUT43), .A2(n1193), .ZN(n1219) );
NAND3_X1 U913 ( .A1(n1204), .A2(n1192), .A3(n1047), .ZN(n1193) );
XNOR2_X1 U914 ( .A(G125), .B(n1168), .ZN(G27) );
NAND4_X1 U915 ( .A1(n1203), .A2(n1220), .A3(n1040), .A4(n1170), .ZN(n1168) );
NAND2_X1 U916 ( .A1(n1021), .A2(n1221), .ZN(n1170) );
NAND4_X1 U917 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1223), .ZN(n1221) );
INV_X1 U918 ( .A(G900), .ZN(n1223) );
AND3_X1 U919 ( .A1(n1048), .A2(n1224), .A3(n1038), .ZN(n1203) );
XNOR2_X1 U920 ( .A(G122), .B(n1194), .ZN(G24) );
NAND3_X1 U921 ( .A1(n1220), .A2(n1024), .A3(n1225), .ZN(n1194) );
NOR3_X1 U922 ( .A1(n1226), .A2(n1201), .A3(n1202), .ZN(n1225) );
NOR2_X1 U923 ( .A1(n1227), .A2(n1224), .ZN(n1024) );
XNOR2_X1 U924 ( .A(G119), .B(n1184), .ZN(G21) );
NAND4_X1 U925 ( .A1(n1176), .A2(n1220), .A3(n1204), .A4(n1228), .ZN(n1184) );
INV_X1 U926 ( .A(n1191), .ZN(n1176) );
NAND2_X1 U927 ( .A1(n1224), .A2(n1227), .ZN(n1191) );
XNOR2_X1 U928 ( .A(G116), .B(n1177), .ZN(G18) );
NAND4_X1 U929 ( .A1(n1220), .A2(n1047), .A3(n1037), .A4(n1228), .ZN(n1177) );
INV_X1 U930 ( .A(n1226), .ZN(n1228) );
AND2_X1 U931 ( .A1(n1229), .A2(n1230), .ZN(n1037) );
XOR2_X1 U932 ( .A(n1202), .B(KEYINPUT59), .Z(n1229) );
XOR2_X1 U933 ( .A(G113), .B(n1231), .Z(G15) );
NOR3_X1 U934 ( .A1(n1189), .A2(n1232), .A3(n1226), .ZN(n1231) );
XNOR2_X1 U935 ( .A(n1220), .B(KEYINPUT52), .ZN(n1232) );
INV_X1 U936 ( .A(n1036), .ZN(n1220) );
NAND2_X1 U937 ( .A1(n1034), .A2(n1233), .ZN(n1036) );
NAND2_X1 U938 ( .A1(G221), .A2(n1234), .ZN(n1233) );
NAND2_X1 U939 ( .A1(n1038), .A2(n1047), .ZN(n1189) );
NOR2_X1 U940 ( .A1(n1224), .A2(n1048), .ZN(n1047) );
NOR2_X1 U941 ( .A1(n1230), .A2(n1202), .ZN(n1038) );
XNOR2_X1 U942 ( .A(n1178), .B(n1235), .ZN(G12) );
NOR2_X1 U943 ( .A1(KEYINPUT40), .A2(n1236), .ZN(n1235) );
INV_X1 U944 ( .A(G110), .ZN(n1236) );
NAND4_X1 U945 ( .A1(n1204), .A2(n1192), .A3(n1048), .A4(n1224), .ZN(n1178) );
XNOR2_X1 U946 ( .A(n1237), .B(n1087), .ZN(n1224) );
AND2_X1 U947 ( .A1(G217), .A2(n1234), .ZN(n1087) );
NAND2_X1 U948 ( .A1(n1085), .A2(n1238), .ZN(n1237) );
XNOR2_X1 U949 ( .A(n1239), .B(n1240), .ZN(n1085) );
XOR2_X1 U950 ( .A(n1241), .B(n1242), .Z(n1240) );
XNOR2_X1 U951 ( .A(G137), .B(n1243), .ZN(n1242) );
NOR2_X1 U952 ( .A1(KEYINPUT24), .A2(n1244), .ZN(n1243) );
XNOR2_X1 U953 ( .A(G110), .B(n1245), .ZN(n1244) );
XOR2_X1 U954 ( .A(G128), .B(G119), .Z(n1245) );
NAND2_X1 U955 ( .A1(KEYINPUT17), .A2(n1246), .ZN(n1241) );
XNOR2_X1 U956 ( .A(n1061), .B(n1247), .ZN(n1239) );
NOR2_X1 U957 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
INV_X1 U958 ( .A(G221), .ZN(n1248) );
INV_X1 U959 ( .A(n1227), .ZN(n1048) );
XNOR2_X1 U960 ( .A(n1250), .B(G472), .ZN(n1227) );
NAND2_X1 U961 ( .A1(n1251), .A2(n1238), .ZN(n1250) );
XOR2_X1 U962 ( .A(n1107), .B(n1252), .Z(n1251) );
XNOR2_X1 U963 ( .A(KEYINPUT2), .B(n1253), .ZN(n1252) );
NOR2_X1 U964 ( .A1(KEYINPUT1), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U965 ( .A(n1255), .B(n1149), .ZN(n1254) );
INV_X1 U966 ( .A(n1108), .ZN(n1149) );
NOR2_X1 U967 ( .A1(KEYINPUT51), .A2(n1110), .ZN(n1255) );
XNOR2_X1 U968 ( .A(n1256), .B(n1257), .ZN(n1107) );
XOR2_X1 U969 ( .A(n1258), .B(G101), .Z(n1256) );
NAND3_X1 U970 ( .A1(G210), .A2(n1057), .A3(n1259), .ZN(n1258) );
XNOR2_X1 U971 ( .A(G237), .B(KEYINPUT16), .ZN(n1259) );
NOR2_X1 U972 ( .A1(n1171), .A2(n1226), .ZN(n1192) );
NAND2_X1 U973 ( .A1(n1040), .A2(n1188), .ZN(n1226) );
NAND2_X1 U974 ( .A1(n1021), .A2(n1260), .ZN(n1188) );
NAND3_X1 U975 ( .A1(G902), .A2(n1222), .A3(n1075), .ZN(n1260) );
NOR2_X1 U976 ( .A1(G898), .A2(n1057), .ZN(n1075) );
NAND3_X1 U977 ( .A1(n1222), .A2(n1057), .A3(G952), .ZN(n1021) );
NAND2_X1 U978 ( .A1(G237), .A2(G234), .ZN(n1222) );
NOR2_X1 U979 ( .A1(n1043), .A2(n1261), .ZN(n1040) );
INV_X1 U980 ( .A(n1218), .ZN(n1261) );
NAND2_X1 U981 ( .A1(G214), .A2(n1262), .ZN(n1218) );
XNOR2_X1 U982 ( .A(n1263), .B(n1195), .ZN(n1043) );
NAND2_X1 U983 ( .A1(G210), .A2(n1262), .ZN(n1195) );
NAND2_X1 U984 ( .A1(n1264), .A2(n1152), .ZN(n1262) );
NAND2_X1 U985 ( .A1(n1265), .A2(n1238), .ZN(n1263) );
XOR2_X1 U986 ( .A(n1266), .B(n1134), .Z(n1265) );
XNOR2_X1 U987 ( .A(n1267), .B(n1079), .ZN(n1134) );
XNOR2_X1 U988 ( .A(n1268), .B(n1269), .ZN(n1079) );
XOR2_X1 U989 ( .A(n1270), .B(n1271), .Z(n1269) );
NOR2_X1 U990 ( .A1(KEYINPUT60), .A2(n1272), .ZN(n1270) );
XNOR2_X1 U991 ( .A(G110), .B(n1273), .ZN(n1268) );
XNOR2_X1 U992 ( .A(KEYINPUT5), .B(n1274), .ZN(n1273) );
NAND2_X1 U993 ( .A1(KEYINPUT26), .A2(n1080), .ZN(n1267) );
XNOR2_X1 U994 ( .A(n1257), .B(KEYINPUT29), .ZN(n1080) );
XNOR2_X1 U995 ( .A(G113), .B(n1275), .ZN(n1257) );
XOR2_X1 U996 ( .A(G119), .B(G116), .Z(n1275) );
NAND3_X1 U997 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1266) );
NAND2_X1 U998 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
OR3_X1 U999 ( .A1(n1280), .A2(n1279), .A3(KEYINPUT63), .ZN(n1277) );
XOR2_X1 U1000 ( .A(n1281), .B(n1108), .Z(n1279) );
XNOR2_X1 U1001 ( .A(n1282), .B(n1246), .ZN(n1108) );
XOR2_X1 U1002 ( .A(n1283), .B(G143), .Z(n1282) );
NAND2_X1 U1003 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1283) );
NAND2_X1 U1004 ( .A1(KEYINPUT27), .A2(n1284), .ZN(n1281) );
OR2_X1 U1005 ( .A1(KEYINPUT41), .A2(n1145), .ZN(n1280) );
NAND2_X1 U1006 ( .A1(KEYINPUT63), .A2(n1145), .ZN(n1276) );
INV_X1 U1007 ( .A(n1147), .ZN(n1145) );
NOR2_X1 U1008 ( .A1(n1074), .A2(G953), .ZN(n1147) );
INV_X1 U1009 ( .A(G224), .ZN(n1074) );
INV_X1 U1010 ( .A(n1033), .ZN(n1171) );
NOR2_X1 U1011 ( .A1(n1034), .A2(n1285), .ZN(n1033) );
AND2_X1 U1012 ( .A1(G221), .A2(n1234), .ZN(n1285) );
NAND2_X1 U1013 ( .A1(G234), .A2(n1152), .ZN(n1234) );
INV_X1 U1014 ( .A(G902), .ZN(n1152) );
XOR2_X1 U1015 ( .A(n1286), .B(G469), .Z(n1034) );
NAND2_X1 U1016 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
XNOR2_X1 U1017 ( .A(n1289), .B(n1130), .ZN(n1288) );
XNOR2_X1 U1018 ( .A(n1290), .B(n1291), .ZN(n1130) );
XNOR2_X1 U1019 ( .A(n1292), .B(G110), .ZN(n1291) );
INV_X1 U1020 ( .A(G140), .ZN(n1292) );
NAND2_X1 U1021 ( .A1(G227), .A2(n1057), .ZN(n1290) );
NAND3_X1 U1022 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1289) );
NAND2_X1 U1023 ( .A1(n1132), .A2(n1110), .ZN(n1295) );
INV_X1 U1024 ( .A(n1296), .ZN(n1132) );
NAND2_X1 U1025 ( .A1(KEYINPUT14), .A2(n1297), .ZN(n1294) );
NAND2_X1 U1026 ( .A1(n1298), .A2(n1131), .ZN(n1297) );
XNOR2_X1 U1027 ( .A(n1296), .B(KEYINPUT45), .ZN(n1298) );
NAND2_X1 U1028 ( .A1(n1299), .A2(n1300), .ZN(n1293) );
INV_X1 U1029 ( .A(KEYINPUT14), .ZN(n1300) );
NAND2_X1 U1030 ( .A1(n1301), .A2(n1302), .ZN(n1299) );
OR2_X1 U1031 ( .A1(n1296), .A2(KEYINPUT45), .ZN(n1302) );
NAND3_X1 U1032 ( .A1(n1131), .A2(n1296), .A3(KEYINPUT45), .ZN(n1301) );
XNOR2_X1 U1033 ( .A(n1303), .B(n1304), .ZN(n1296) );
XNOR2_X1 U1034 ( .A(KEYINPUT19), .B(n1272), .ZN(n1304) );
INV_X1 U1035 ( .A(G107), .ZN(n1272) );
XOR2_X1 U1036 ( .A(n1066), .B(n1271), .Z(n1303) );
XNOR2_X1 U1037 ( .A(G101), .B(n1305), .ZN(n1271) );
XOR2_X1 U1038 ( .A(n1306), .B(n1307), .Z(n1066) );
XOR2_X1 U1039 ( .A(n1308), .B(n1246), .Z(n1307) );
NOR2_X1 U1040 ( .A1(G128), .A2(KEYINPUT49), .ZN(n1308) );
XNOR2_X1 U1041 ( .A(G143), .B(KEYINPUT38), .ZN(n1306) );
INV_X1 U1042 ( .A(n1110), .ZN(n1131) );
NAND2_X1 U1043 ( .A1(n1309), .A2(n1310), .ZN(n1110) );
NAND2_X1 U1044 ( .A1(G131), .A2(n1311), .ZN(n1310) );
XOR2_X1 U1045 ( .A(n1312), .B(KEYINPUT35), .Z(n1309) );
OR2_X1 U1046 ( .A1(n1311), .A2(G131), .ZN(n1312) );
NAND2_X1 U1047 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NAND2_X1 U1048 ( .A1(G134), .A2(n1065), .ZN(n1314) );
XOR2_X1 U1049 ( .A(KEYINPUT33), .B(n1315), .Z(n1313) );
NOR2_X1 U1050 ( .A1(G134), .A2(n1065), .ZN(n1315) );
INV_X1 U1051 ( .A(G137), .ZN(n1065) );
XNOR2_X1 U1052 ( .A(n1238), .B(KEYINPUT47), .ZN(n1287) );
INV_X1 U1053 ( .A(n1032), .ZN(n1204) );
NAND2_X1 U1054 ( .A1(n1201), .A2(n1202), .ZN(n1032) );
XOR2_X1 U1055 ( .A(n1316), .B(G475), .Z(n1202) );
NAND2_X1 U1056 ( .A1(n1096), .A2(n1238), .ZN(n1316) );
XOR2_X1 U1057 ( .A(n1317), .B(n1318), .Z(n1096) );
XOR2_X1 U1058 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1059 ( .A(n1274), .B(G113), .ZN(n1320) );
INV_X1 U1060 ( .A(G122), .ZN(n1274) );
NOR2_X1 U1061 ( .A1(KEYINPUT54), .A2(n1321), .ZN(n1319) );
NOR2_X1 U1062 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1063 ( .A(KEYINPUT8), .B(n1324), .Z(n1323) );
NOR2_X1 U1064 ( .A1(G131), .A2(n1325), .ZN(n1324) );
AND2_X1 U1065 ( .A1(G131), .A2(n1325), .ZN(n1322) );
XNOR2_X1 U1066 ( .A(G143), .B(n1326), .ZN(n1325) );
AND3_X1 U1067 ( .A1(G214), .A2(n1057), .A3(n1264), .ZN(n1326) );
INV_X1 U1068 ( .A(G237), .ZN(n1264) );
XOR2_X1 U1069 ( .A(n1327), .B(n1061), .Z(n1317) );
XNOR2_X1 U1070 ( .A(G140), .B(n1150), .ZN(n1061) );
INV_X1 U1071 ( .A(n1284), .ZN(n1150) );
XOR2_X1 U1072 ( .A(G125), .B(KEYINPUT42), .Z(n1284) );
XOR2_X1 U1073 ( .A(n1328), .B(n1246), .Z(n1327) );
XOR2_X1 U1074 ( .A(G146), .B(KEYINPUT15), .Z(n1246) );
NAND2_X1 U1075 ( .A1(KEYINPUT30), .A2(n1305), .ZN(n1328) );
INV_X1 U1076 ( .A(G104), .ZN(n1305) );
INV_X1 U1077 ( .A(n1230), .ZN(n1201) );
XNOR2_X1 U1078 ( .A(n1329), .B(G478), .ZN(n1230) );
NAND2_X1 U1079 ( .A1(n1091), .A2(n1238), .ZN(n1329) );
XOR2_X1 U1080 ( .A(G902), .B(KEYINPUT28), .Z(n1238) );
XOR2_X1 U1081 ( .A(n1330), .B(n1331), .Z(n1091) );
XOR2_X1 U1082 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1083 ( .A(n1334), .B(n1335), .ZN(n1333) );
NOR3_X1 U1084 ( .A1(n1249), .A2(KEYINPUT32), .A3(n1336), .ZN(n1335) );
INV_X1 U1085 ( .A(G217), .ZN(n1336) );
NAND2_X1 U1086 ( .A1(n1337), .A2(n1057), .ZN(n1249) );
INV_X1 U1087 ( .A(G953), .ZN(n1057) );
XOR2_X1 U1088 ( .A(KEYINPUT25), .B(G234), .Z(n1337) );
NOR2_X1 U1089 ( .A1(KEYINPUT22), .A2(G143), .ZN(n1334) );
XNOR2_X1 U1090 ( .A(G116), .B(G107), .ZN(n1332) );
XOR2_X1 U1091 ( .A(n1338), .B(n1339), .Z(n1330) );
XNOR2_X1 U1092 ( .A(KEYINPUT7), .B(n1209), .ZN(n1339) );
INV_X1 U1093 ( .A(G134), .ZN(n1209) );
XNOR2_X1 U1094 ( .A(G122), .B(G128), .ZN(n1338) );
endmodule


