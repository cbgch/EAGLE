//Key = 0111100110000011000111010100010110110011101001100000101100101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310;

XOR2_X1 U711 ( .A(n1007), .B(n1008), .Z(G9) );
NOR2_X1 U712 ( .A1(n1009), .A2(n1010), .ZN(G75) );
XOR2_X1 U713 ( .A(n1011), .B(KEYINPUT38), .Z(n1010) );
NAND4_X1 U714 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
NAND3_X1 U715 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
INV_X1 U716 ( .A(n1019), .ZN(n1018) );
NAND2_X1 U717 ( .A1(n1020), .A2(n1021), .ZN(n1017) );
NAND4_X1 U718 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
OR2_X1 U719 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U720 ( .A1(n1028), .A2(n1029), .ZN(n1020) );
NAND2_X1 U721 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND3_X1 U722 ( .A1(n1032), .A2(n1033), .A3(n1022), .ZN(n1031) );
NAND2_X1 U723 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND3_X1 U724 ( .A1(n1036), .A2(n1037), .A3(n1024), .ZN(n1032) );
NAND2_X1 U725 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NAND2_X1 U726 ( .A1(n1040), .A2(n1023), .ZN(n1030) );
NAND4_X1 U727 ( .A1(n1024), .A2(n1041), .A3(n1022), .A4(n1042), .ZN(n1014) );
NOR3_X1 U728 ( .A1(n1019), .A2(n1035), .A3(n1043), .ZN(n1042) );
NAND2_X1 U729 ( .A1(n1044), .A2(n1045), .ZN(n1041) );
NAND2_X1 U730 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
XOR2_X1 U731 ( .A(n1048), .B(KEYINPUT37), .Z(n1046) );
INV_X1 U732 ( .A(n1049), .ZN(n1013) );
NOR2_X1 U733 ( .A1(G952), .A2(n1049), .ZN(n1009) );
NAND2_X1 U734 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND4_X1 U735 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
NOR3_X1 U736 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
AND2_X1 U737 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U738 ( .A(n1061), .B(KEYINPUT31), .Z(n1054) );
NAND3_X1 U739 ( .A1(n1023), .A2(n1062), .A3(n1063), .ZN(n1061) );
XOR2_X1 U740 ( .A(n1064), .B(n1065), .Z(n1063) );
XOR2_X1 U741 ( .A(G472), .B(n1066), .Z(n1053) );
NOR2_X1 U742 ( .A1(n1067), .A2(KEYINPUT9), .ZN(n1066) );
XOR2_X1 U743 ( .A(n1068), .B(n1069), .Z(G72) );
XOR2_X1 U744 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND2_X1 U745 ( .A1(G953), .A2(n1072), .ZN(n1071) );
NAND2_X1 U746 ( .A1(G900), .A2(G227), .ZN(n1072) );
NAND2_X1 U747 ( .A1(n1073), .A2(n1074), .ZN(n1070) );
NAND2_X1 U748 ( .A1(G953), .A2(n1075), .ZN(n1074) );
XOR2_X1 U749 ( .A(n1076), .B(n1077), .Z(n1073) );
XOR2_X1 U750 ( .A(n1078), .B(n1079), .Z(n1077) );
XNOR2_X1 U751 ( .A(n1080), .B(n1081), .ZN(n1078) );
XOR2_X1 U752 ( .A(n1082), .B(n1083), .Z(n1076) );
NOR2_X1 U753 ( .A1(G131), .A2(KEYINPUT6), .ZN(n1083) );
XOR2_X1 U754 ( .A(n1084), .B(KEYINPUT62), .Z(n1082) );
NAND2_X1 U755 ( .A1(KEYINPUT21), .A2(n1085), .ZN(n1084) );
NOR2_X1 U756 ( .A1(n1086), .A2(G953), .ZN(n1068) );
NAND2_X1 U757 ( .A1(n1087), .A2(n1088), .ZN(G69) );
NAND2_X1 U758 ( .A1(G953), .A2(n1089), .ZN(n1088) );
XOR2_X1 U759 ( .A(n1090), .B(n1091), .Z(n1087) );
NOR2_X1 U760 ( .A1(KEYINPUT33), .A2(n1092), .ZN(n1091) );
XOR2_X1 U761 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U762 ( .A(n1095), .B(n1096), .Z(n1093) );
NAND2_X1 U763 ( .A1(KEYINPUT29), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U764 ( .A(G101), .B(n1098), .ZN(n1097) );
NAND2_X1 U765 ( .A1(n1099), .A2(n1100), .ZN(n1090) );
NAND3_X1 U766 ( .A1(n1101), .A2(n1102), .A3(n1050), .ZN(n1100) );
XOR2_X1 U767 ( .A(n1103), .B(KEYINPUT44), .Z(n1102) );
NAND2_X1 U768 ( .A1(G953), .A2(G224), .ZN(n1099) );
NOR2_X1 U769 ( .A1(n1104), .A2(n1105), .ZN(G66) );
XOR2_X1 U770 ( .A(n1106), .B(n1107), .Z(n1105) );
NAND2_X1 U771 ( .A1(n1108), .A2(n1060), .ZN(n1106) );
NOR2_X1 U772 ( .A1(n1104), .A2(n1109), .ZN(G63) );
XOR2_X1 U773 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U774 ( .A1(n1108), .A2(G478), .ZN(n1110) );
NOR2_X1 U775 ( .A1(n1104), .A2(n1112), .ZN(G60) );
XNOR2_X1 U776 ( .A(n1113), .B(n1114), .ZN(n1112) );
NAND2_X1 U777 ( .A1(n1108), .A2(G475), .ZN(n1113) );
XOR2_X1 U778 ( .A(n1115), .B(n1116), .Z(G6) );
NAND2_X1 U779 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U780 ( .A(n1119), .B(KEYINPUT46), .Z(n1117) );
NOR2_X1 U781 ( .A1(n1104), .A2(n1120), .ZN(G57) );
XOR2_X1 U782 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U783 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U784 ( .A(n1125), .B(n1080), .Z(n1123) );
NAND3_X1 U785 ( .A1(n1108), .A2(G472), .A3(KEYINPUT23), .ZN(n1125) );
XNOR2_X1 U786 ( .A(n1126), .B(n1127), .ZN(n1121) );
XNOR2_X1 U787 ( .A(G101), .B(KEYINPUT7), .ZN(n1126) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1128), .ZN(G54) );
XOR2_X1 U789 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U790 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U791 ( .A(G110), .B(n1133), .Z(n1132) );
NOR2_X1 U792 ( .A1(KEYINPUT0), .A2(n1134), .ZN(n1133) );
XNOR2_X1 U793 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U794 ( .A(KEYINPUT57), .B(G140), .Z(n1131) );
XOR2_X1 U795 ( .A(n1137), .B(n1138), .Z(n1129) );
XOR2_X1 U796 ( .A(n1139), .B(n1140), .Z(n1137) );
NAND2_X1 U797 ( .A1(n1108), .A2(G469), .ZN(n1139) );
NOR2_X1 U798 ( .A1(n1104), .A2(n1141), .ZN(G51) );
XOR2_X1 U799 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U800 ( .A1(n1108), .A2(G210), .ZN(n1142) );
NOR2_X1 U801 ( .A1(n1144), .A2(n1012), .ZN(n1108) );
AND3_X1 U802 ( .A1(n1101), .A2(n1103), .A3(n1086), .ZN(n1012) );
AND4_X1 U803 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1086) );
AND4_X1 U804 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
NAND2_X1 U805 ( .A1(n1026), .A2(n1153), .ZN(n1147) );
NAND2_X1 U806 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND3_X1 U807 ( .A1(n1156), .A2(n1023), .A3(n1157), .ZN(n1154) );
XOR2_X1 U808 ( .A(n1158), .B(KEYINPUT22), .Z(n1157) );
AND4_X1 U809 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1101) );
AND3_X1 U810 ( .A1(n1008), .A2(n1163), .A3(n1164), .ZN(n1162) );
NAND4_X1 U811 ( .A1(n1165), .A2(n1118), .A3(n1027), .A4(n1166), .ZN(n1008) );
NAND2_X1 U812 ( .A1(n1118), .A2(n1167), .ZN(n1161) );
NAND2_X1 U813 ( .A1(n1168), .A2(n1119), .ZN(n1167) );
NAND3_X1 U814 ( .A1(n1165), .A2(n1166), .A3(n1026), .ZN(n1119) );
XOR2_X1 U815 ( .A(KEYINPUT35), .B(n1169), .Z(n1168) );
NOR2_X1 U816 ( .A1(n1050), .A2(G952), .ZN(n1104) );
NAND2_X1 U817 ( .A1(n1170), .A2(n1171), .ZN(G48) );
NAND2_X1 U818 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U819 ( .A(KEYINPUT1), .B(n1174), .Z(n1170) );
NOR2_X1 U820 ( .A1(n1172), .A2(n1173), .ZN(n1174) );
INV_X1 U821 ( .A(n1146), .ZN(n1172) );
NAND3_X1 U822 ( .A1(n1175), .A2(n1118), .A3(n1026), .ZN(n1146) );
XOR2_X1 U823 ( .A(n1176), .B(n1145), .Z(G45) );
NAND3_X1 U824 ( .A1(n1156), .A2(n1158), .A3(n1177), .ZN(n1145) );
XOR2_X1 U825 ( .A(n1178), .B(n1152), .Z(G42) );
NAND4_X1 U826 ( .A1(n1165), .A2(n1158), .A3(n1023), .A4(n1179), .ZN(n1152) );
NOR2_X1 U827 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U828 ( .A(n1151), .B(n1182), .Z(G39) );
NAND2_X1 U829 ( .A1(KEYINPUT61), .A2(G137), .ZN(n1182) );
NAND3_X1 U830 ( .A1(n1175), .A2(n1023), .A3(n1028), .ZN(n1151) );
XOR2_X1 U831 ( .A(n1150), .B(n1183), .Z(G36) );
XOR2_X1 U832 ( .A(KEYINPUT2), .B(G134), .Z(n1183) );
NAND4_X1 U833 ( .A1(n1156), .A2(n1023), .A3(n1027), .A4(n1158), .ZN(n1150) );
XOR2_X1 U834 ( .A(n1184), .B(n1185), .Z(G33) );
NAND4_X1 U835 ( .A1(n1026), .A2(n1156), .A3(n1023), .A4(n1158), .ZN(n1185) );
INV_X1 U836 ( .A(n1035), .ZN(n1023) );
NAND2_X1 U837 ( .A1(n1039), .A2(n1186), .ZN(n1035) );
XNOR2_X1 U838 ( .A(G128), .B(n1149), .ZN(G30) );
NAND3_X1 U839 ( .A1(n1118), .A2(n1027), .A3(n1175), .ZN(n1149) );
AND4_X1 U840 ( .A1(n1034), .A2(n1165), .A3(n1158), .A4(n1187), .ZN(n1175) );
XOR2_X1 U841 ( .A(n1159), .B(n1188), .Z(G3) );
NAND2_X1 U842 ( .A1(KEYINPUT19), .A2(G101), .ZN(n1188) );
NAND2_X1 U843 ( .A1(n1189), .A2(n1156), .ZN(n1159) );
AND3_X1 U844 ( .A1(n1022), .A2(n1165), .A3(n1034), .ZN(n1156) );
XOR2_X1 U845 ( .A(n1190), .B(n1191), .Z(G27) );
NAND2_X1 U846 ( .A1(KEYINPUT54), .A2(G125), .ZN(n1191) );
NAND2_X1 U847 ( .A1(n1192), .A2(n1193), .ZN(n1190) );
INV_X1 U848 ( .A(n1155), .ZN(n1193) );
NAND4_X1 U849 ( .A1(n1016), .A2(n1040), .A3(n1118), .A4(n1158), .ZN(n1155) );
NAND2_X1 U850 ( .A1(n1019), .A2(n1194), .ZN(n1158) );
NAND4_X1 U851 ( .A1(G953), .A2(G902), .A3(n1195), .A4(n1075), .ZN(n1194) );
INV_X1 U852 ( .A(G900), .ZN(n1075) );
XOR2_X1 U853 ( .A(n1181), .B(KEYINPUT20), .Z(n1192) );
XNOR2_X1 U854 ( .A(G122), .B(n1103), .ZN(G24) );
NAND3_X1 U855 ( .A1(n1177), .A2(n1166), .A3(n1016), .ZN(n1103) );
AND3_X1 U856 ( .A1(n1024), .A2(n1196), .A3(n1022), .ZN(n1166) );
NOR3_X1 U857 ( .A1(n1037), .A2(n1052), .A3(n1197), .ZN(n1177) );
INV_X1 U858 ( .A(n1118), .ZN(n1037) );
XNOR2_X1 U859 ( .A(G119), .B(n1160), .ZN(G21) );
NAND4_X1 U860 ( .A1(n1189), .A2(n1016), .A3(n1034), .A4(n1187), .ZN(n1160) );
XOR2_X1 U861 ( .A(n1198), .B(n1199), .Z(G18) );
XOR2_X1 U862 ( .A(KEYINPUT55), .B(G116), .Z(n1199) );
NAND2_X1 U863 ( .A1(n1169), .A2(n1118), .ZN(n1198) );
AND2_X1 U864 ( .A1(n1200), .A2(n1027), .ZN(n1169) );
NOR2_X1 U865 ( .A1(n1056), .A2(n1052), .ZN(n1027) );
XNOR2_X1 U866 ( .A(G113), .B(n1164), .ZN(G15) );
NAND3_X1 U867 ( .A1(n1026), .A2(n1118), .A3(n1200), .ZN(n1164) );
AND4_X1 U868 ( .A1(n1034), .A2(n1016), .A3(n1022), .A4(n1196), .ZN(n1200) );
XOR2_X1 U869 ( .A(n1187), .B(KEYINPUT8), .Z(n1022) );
NOR2_X1 U870 ( .A1(n1201), .A2(n1047), .ZN(n1016) );
INV_X1 U871 ( .A(n1062), .ZN(n1047) );
INV_X1 U872 ( .A(n1181), .ZN(n1026) );
NAND2_X1 U873 ( .A1(n1056), .A2(n1202), .ZN(n1181) );
XOR2_X1 U874 ( .A(n1203), .B(n1163), .Z(G12) );
NAND3_X1 U875 ( .A1(n1040), .A2(n1165), .A3(n1189), .ZN(n1163) );
AND3_X1 U876 ( .A1(n1118), .A2(n1196), .A3(n1028), .ZN(n1189) );
INV_X1 U877 ( .A(n1043), .ZN(n1028) );
NAND2_X1 U878 ( .A1(n1202), .A2(n1197), .ZN(n1043) );
INV_X1 U879 ( .A(n1056), .ZN(n1197) );
XOR2_X1 U880 ( .A(n1204), .B(n1205), .Z(n1056) );
NOR2_X1 U881 ( .A1(n1206), .A2(n1114), .ZN(n1205) );
XNOR2_X1 U882 ( .A(n1207), .B(n1208), .ZN(n1114) );
XOR2_X1 U883 ( .A(n1209), .B(n1210), .Z(n1208) );
NAND2_X1 U884 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND2_X1 U885 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NAND2_X1 U886 ( .A1(KEYINPUT14), .A2(n1215), .ZN(n1213) );
NAND2_X1 U887 ( .A1(KEYINPUT4), .A2(n1184), .ZN(n1215) );
NAND2_X1 U888 ( .A1(G131), .A2(n1216), .ZN(n1211) );
NAND2_X1 U889 ( .A1(KEYINPUT4), .A2(n1217), .ZN(n1216) );
NAND2_X1 U890 ( .A1(n1218), .A2(KEYINPUT14), .ZN(n1217) );
INV_X1 U891 ( .A(n1214), .ZN(n1218) );
NAND2_X1 U892 ( .A1(n1219), .A2(n1220), .ZN(n1214) );
NAND2_X1 U893 ( .A1(n1221), .A2(n1176), .ZN(n1220) );
XOR2_X1 U894 ( .A(KEYINPUT60), .B(n1222), .Z(n1219) );
NOR2_X1 U895 ( .A1(n1176), .A2(n1221), .ZN(n1222) );
NAND3_X1 U896 ( .A1(n1223), .A2(n1050), .A3(G214), .ZN(n1221) );
INV_X1 U897 ( .A(G143), .ZN(n1176) );
NAND2_X1 U898 ( .A1(n1224), .A2(n1225), .ZN(n1209) );
NAND2_X1 U899 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U900 ( .A(KEYINPUT45), .B(n1228), .Z(n1224) );
NOR2_X1 U901 ( .A1(n1227), .A2(n1226), .ZN(n1228) );
XOR2_X1 U902 ( .A(KEYINPUT26), .B(G104), .Z(n1226) );
XOR2_X1 U903 ( .A(G113), .B(G122), .Z(n1227) );
XOR2_X1 U904 ( .A(n1229), .B(G146), .Z(n1207) );
NAND3_X1 U905 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1229) );
OR2_X1 U906 ( .A1(n1178), .A2(KEYINPUT34), .ZN(n1232) );
NAND3_X1 U907 ( .A1(KEYINPUT34), .A2(n1178), .A3(G125), .ZN(n1231) );
NAND2_X1 U908 ( .A1(n1233), .A2(n1234), .ZN(n1230) );
INV_X1 U909 ( .A(G125), .ZN(n1234) );
NAND2_X1 U910 ( .A1(n1235), .A2(KEYINPUT34), .ZN(n1233) );
XOR2_X1 U911 ( .A(n1178), .B(KEYINPUT18), .Z(n1235) );
XOR2_X1 U912 ( .A(n1144), .B(KEYINPUT42), .Z(n1206) );
XNOR2_X1 U913 ( .A(G475), .B(KEYINPUT15), .ZN(n1204) );
XNOR2_X1 U914 ( .A(n1052), .B(KEYINPUT40), .ZN(n1202) );
XNOR2_X1 U915 ( .A(G478), .B(n1236), .ZN(n1052) );
AND2_X1 U916 ( .A1(n1144), .A2(n1111), .ZN(n1236) );
XNOR2_X1 U917 ( .A(n1237), .B(n1238), .ZN(n1111) );
NOR2_X1 U918 ( .A1(n1239), .A2(KEYINPUT47), .ZN(n1238) );
NOR2_X1 U919 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
INV_X1 U920 ( .A(G217), .ZN(n1241) );
NAND2_X1 U921 ( .A1(n1242), .A2(n1243), .ZN(n1237) );
NAND2_X1 U922 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U923 ( .A(n1246), .B(KEYINPUT5), .Z(n1242) );
NAND2_X1 U924 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
INV_X1 U925 ( .A(n1244), .ZN(n1248) );
XOR2_X1 U926 ( .A(n1249), .B(n1250), .Z(n1244) );
XOR2_X1 U927 ( .A(G107), .B(n1251), .Z(n1250) );
NOR2_X1 U928 ( .A1(G116), .A2(KEYINPUT63), .ZN(n1251) );
XNOR2_X1 U929 ( .A(G122), .B(KEYINPUT59), .ZN(n1249) );
XNOR2_X1 U930 ( .A(n1245), .B(KEYINPUT53), .ZN(n1247) );
XNOR2_X1 U931 ( .A(n1252), .B(n1253), .ZN(n1245) );
NOR2_X1 U932 ( .A1(G143), .A2(KEYINPUT30), .ZN(n1253) );
XOR2_X1 U933 ( .A(n1254), .B(G128), .Z(n1252) );
INV_X1 U934 ( .A(G134), .ZN(n1254) );
NAND2_X1 U935 ( .A1(n1019), .A2(n1255), .ZN(n1196) );
NAND4_X1 U936 ( .A1(G953), .A2(G902), .A3(n1195), .A4(n1089), .ZN(n1255) );
INV_X1 U937 ( .A(G898), .ZN(n1089) );
NAND3_X1 U938 ( .A1(n1195), .A2(n1050), .A3(G952), .ZN(n1019) );
NAND2_X1 U939 ( .A1(G237), .A2(G234), .ZN(n1195) );
NOR2_X1 U940 ( .A1(n1039), .A2(n1038), .ZN(n1118) );
INV_X1 U941 ( .A(n1186), .ZN(n1038) );
NAND2_X1 U942 ( .A1(G214), .A2(n1256), .ZN(n1186) );
XOR2_X1 U943 ( .A(n1257), .B(n1258), .Z(n1039) );
NOR2_X1 U944 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U945 ( .A(KEYINPUT52), .B(G210), .Z(n1260) );
INV_X1 U946 ( .A(n1256), .ZN(n1259) );
NAND2_X1 U947 ( .A1(n1144), .A2(n1223), .ZN(n1256) );
NAND2_X1 U948 ( .A1(n1261), .A2(n1144), .ZN(n1257) );
XOR2_X1 U949 ( .A(KEYINPUT3), .B(n1262), .Z(n1261) );
INV_X1 U950 ( .A(n1143), .ZN(n1262) );
XOR2_X1 U951 ( .A(n1263), .B(n1264), .Z(n1143) );
XOR2_X1 U952 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U953 ( .A(G125), .B(n1267), .Z(n1266) );
NOR2_X1 U954 ( .A1(KEYINPUT56), .A2(n1096), .ZN(n1267) );
AND2_X1 U955 ( .A1(n1050), .A2(G224), .ZN(n1265) );
XOR2_X1 U956 ( .A(n1268), .B(n1098), .Z(n1263) );
AND2_X1 U957 ( .A1(n1269), .A2(n1270), .ZN(n1098) );
NAND2_X1 U958 ( .A1(KEYINPUT32), .A2(n1136), .ZN(n1270) );
OR3_X1 U959 ( .A1(n1115), .A2(G107), .A3(KEYINPUT32), .ZN(n1269) );
INV_X1 U960 ( .A(G104), .ZN(n1115) );
XOR2_X1 U961 ( .A(n1135), .B(n1094), .Z(n1268) );
XOR2_X1 U962 ( .A(G110), .B(G122), .Z(n1094) );
INV_X1 U963 ( .A(n1045), .ZN(n1165) );
NAND2_X1 U964 ( .A1(n1201), .A2(n1062), .ZN(n1045) );
NAND2_X1 U965 ( .A1(G221), .A2(n1271), .ZN(n1062) );
INV_X1 U966 ( .A(n1048), .ZN(n1201) );
XNOR2_X1 U967 ( .A(n1065), .B(n1272), .ZN(n1048) );
NOR2_X1 U968 ( .A1(KEYINPUT10), .A2(n1273), .ZN(n1272) );
XOR2_X1 U969 ( .A(n1064), .B(KEYINPUT36), .Z(n1273) );
NAND2_X1 U970 ( .A1(n1274), .A2(n1144), .ZN(n1064) );
XOR2_X1 U971 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U972 ( .A(n1136), .B(n1138), .ZN(n1276) );
XOR2_X1 U973 ( .A(n1277), .B(KEYINPUT43), .Z(n1138) );
XOR2_X1 U974 ( .A(G104), .B(n1007), .Z(n1136) );
INV_X1 U975 ( .A(G107), .ZN(n1007) );
XOR2_X1 U976 ( .A(n1278), .B(n1279), .Z(n1275) );
XNOR2_X1 U977 ( .A(G101), .B(n1280), .ZN(n1279) );
NAND2_X1 U978 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U979 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U980 ( .A(G140), .B(n1285), .Z(n1283) );
XOR2_X1 U981 ( .A(n1286), .B(KEYINPUT11), .Z(n1281) );
NAND2_X1 U982 ( .A1(n1287), .A2(n1140), .ZN(n1286) );
INV_X1 U983 ( .A(n1284), .ZN(n1140) );
NAND2_X1 U984 ( .A1(G227), .A2(n1050), .ZN(n1284) );
XOR2_X1 U985 ( .A(n1178), .B(n1285), .Z(n1287) );
NOR2_X1 U986 ( .A1(KEYINPUT50), .A2(n1203), .ZN(n1285) );
INV_X1 U987 ( .A(G140), .ZN(n1178) );
NAND2_X1 U988 ( .A1(KEYINPUT39), .A2(n1080), .ZN(n1278) );
XOR2_X1 U989 ( .A(G469), .B(KEYINPUT41), .Z(n1065) );
INV_X1 U990 ( .A(n1180), .ZN(n1040) );
NAND2_X1 U991 ( .A1(n1288), .A2(n1024), .ZN(n1180) );
INV_X1 U992 ( .A(n1034), .ZN(n1024) );
XNOR2_X1 U993 ( .A(G472), .B(n1289), .ZN(n1034) );
NOR2_X1 U994 ( .A1(KEYINPUT12), .A2(n1290), .ZN(n1289) );
XOR2_X1 U995 ( .A(KEYINPUT27), .B(n1067), .Z(n1290) );
AND2_X1 U996 ( .A1(n1291), .A2(n1144), .ZN(n1067) );
XOR2_X1 U997 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U998 ( .A(n1135), .B(n1124), .Z(n1293) );
XOR2_X1 U999 ( .A(n1096), .B(n1277), .Z(n1124) );
XNOR2_X1 U1000 ( .A(n1294), .B(n1081), .ZN(n1277) );
XOR2_X1 U1001 ( .A(G134), .B(KEYINPUT13), .Z(n1081) );
XOR2_X1 U1002 ( .A(n1184), .B(G137), .Z(n1294) );
INV_X1 U1003 ( .A(G131), .ZN(n1184) );
XOR2_X1 U1004 ( .A(G113), .B(n1295), .Z(n1096) );
XOR2_X1 U1005 ( .A(G119), .B(G116), .Z(n1295) );
XNOR2_X1 U1006 ( .A(n1080), .B(G101), .ZN(n1135) );
XOR2_X1 U1007 ( .A(G128), .B(n1296), .Z(n1080) );
XOR2_X1 U1008 ( .A(G146), .B(G143), .Z(n1296) );
XOR2_X1 U1009 ( .A(n1127), .B(KEYINPUT17), .Z(n1292) );
NAND3_X1 U1010 ( .A1(G210), .A2(n1223), .A3(n1297), .ZN(n1127) );
XOR2_X1 U1011 ( .A(n1050), .B(KEYINPUT28), .Z(n1297) );
INV_X1 U1012 ( .A(G237), .ZN(n1223) );
XOR2_X1 U1013 ( .A(n1187), .B(KEYINPUT51), .Z(n1288) );
NAND2_X1 U1014 ( .A1(n1298), .A2(n1299), .ZN(n1187) );
NAND2_X1 U1015 ( .A1(n1060), .A2(n1059), .ZN(n1299) );
XOR2_X1 U1016 ( .A(KEYINPUT58), .B(n1057), .Z(n1298) );
NOR2_X1 U1017 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
AND2_X1 U1018 ( .A1(G217), .A2(n1271), .ZN(n1060) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1144), .ZN(n1271) );
NAND2_X1 U1020 ( .A1(n1107), .A2(n1144), .ZN(n1059) );
INV_X1 U1021 ( .A(G902), .ZN(n1144) );
XNOR2_X1 U1022 ( .A(n1300), .B(n1301), .ZN(n1107) );
XOR2_X1 U1023 ( .A(n1302), .B(n1079), .Z(n1301) );
XOR2_X1 U1024 ( .A(G125), .B(G140), .Z(n1079) );
NOR2_X1 U1025 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
XNOR2_X1 U1026 ( .A(KEYINPUT25), .B(KEYINPUT24), .ZN(n1304) );
XOR2_X1 U1027 ( .A(n1085), .B(n1305), .Z(n1303) );
NOR3_X1 U1028 ( .A1(n1240), .A2(KEYINPUT48), .A3(n1306), .ZN(n1305) );
INV_X1 U1029 ( .A(G221), .ZN(n1306) );
NAND2_X1 U1030 ( .A1(G234), .A2(n1050), .ZN(n1240) );
INV_X1 U1031 ( .A(G953), .ZN(n1050) );
INV_X1 U1032 ( .A(G137), .ZN(n1085) );
XOR2_X1 U1033 ( .A(n1307), .B(n1308), .Z(n1300) );
NOR2_X1 U1034 ( .A1(KEYINPUT16), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1035 ( .A(n1203), .B(n1310), .Z(n1309) );
XOR2_X1 U1036 ( .A(G128), .B(G119), .Z(n1310) );
XOR2_X1 U1037 ( .A(n1173), .B(KEYINPUT49), .Z(n1307) );
INV_X1 U1038 ( .A(G146), .ZN(n1173) );
INV_X1 U1039 ( .A(G110), .ZN(n1203) );
endmodule


