//Key = 0100001010010100011010010000000100110100100100001101001101011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300;

XOR2_X1 U709 ( .A(n984), .B(n985), .Z(G9) );
NAND2_X1 U710 ( .A1(KEYINPUT63), .A2(n986), .ZN(n984) );
NOR2_X1 U711 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR4_X1 U712 ( .A1(n989), .A2(n990), .A3(n991), .A4(n992), .ZN(n988) );
INV_X1 U713 ( .A(G952), .ZN(n991) );
NAND4_X1 U714 ( .A1(n993), .A2(n994), .A3(n995), .A4(n996), .ZN(n989) );
NAND2_X1 U715 ( .A1(n997), .A2(n998), .ZN(n994) );
NAND2_X1 U716 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND4_X1 U717 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
NAND2_X1 U718 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U719 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND3_X1 U720 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1003) );
NAND2_X1 U721 ( .A1(n1007), .A2(n1012), .ZN(n1010) );
NAND2_X1 U722 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U723 ( .A1(n1008), .A2(n1015), .ZN(n1009) );
NAND2_X1 U724 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U725 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND4_X1 U726 ( .A1(n1020), .A2(n1021), .A3(n1007), .A4(n1022), .ZN(n999) );
NOR2_X1 U727 ( .A1(n1005), .A2(n1023), .ZN(n1022) );
NAND2_X1 U728 ( .A1(n1024), .A2(n1025), .ZN(n1021) );
NAND3_X1 U729 ( .A1(n1026), .A2(n1027), .A3(n1002), .ZN(n1020) );
INV_X1 U730 ( .A(n1028), .ZN(n997) );
XNOR2_X1 U731 ( .A(KEYINPUT39), .B(n1029), .ZN(n993) );
NOR3_X1 U732 ( .A1(n1030), .A2(G953), .A3(n1031), .ZN(n987) );
INV_X1 U733 ( .A(n995), .ZN(n1031) );
NAND4_X1 U734 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n995) );
NOR4_X1 U735 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
XOR2_X1 U736 ( .A(n1040), .B(n1041), .Z(n1036) );
NOR2_X1 U737 ( .A1(G472), .A2(KEYINPUT7), .ZN(n1041) );
NOR3_X1 U738 ( .A1(n1005), .A2(n1042), .A3(n1018), .ZN(n1034) );
INV_X1 U739 ( .A(n1011), .ZN(n1005) );
NAND2_X1 U740 ( .A1(n1043), .A2(n1044), .ZN(n1033) );
XOR2_X1 U741 ( .A(n1045), .B(n1046), .Z(n1032) );
NOR2_X1 U742 ( .A1(n1047), .A2(KEYINPUT26), .ZN(n1046) );
XOR2_X1 U743 ( .A(KEYINPUT46), .B(G952), .Z(n1030) );
XOR2_X1 U744 ( .A(n1048), .B(n1049), .Z(G72) );
XOR2_X1 U745 ( .A(n1050), .B(n1051), .Z(n1049) );
NOR2_X1 U746 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U747 ( .A(n996), .B(KEYINPUT30), .Z(n1053) );
AND2_X1 U748 ( .A1(G227), .A2(G900), .ZN(n1052) );
NAND2_X1 U749 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
INV_X1 U750 ( .A(n1056), .ZN(n1055) );
XNOR2_X1 U751 ( .A(n1057), .B(n1058), .ZN(n1054) );
NAND2_X1 U752 ( .A1(n1059), .A2(KEYINPUT8), .ZN(n1057) );
XOR2_X1 U753 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR2_X1 U754 ( .A1(KEYINPUT25), .A2(n1062), .ZN(n1061) );
NAND2_X1 U755 ( .A1(n1063), .A2(n1064), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
INV_X1 U757 ( .A(n990), .ZN(n1065) );
XOR2_X1 U758 ( .A(n996), .B(KEYINPUT28), .Z(n1063) );
NAND2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(G69) );
NAND2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U761 ( .A1(G953), .A2(n1071), .ZN(n1070) );
NAND3_X1 U762 ( .A1(n1072), .A2(n1073), .A3(G953), .ZN(n1067) );
NAND2_X1 U763 ( .A1(G898), .A2(G224), .ZN(n1073) );
XOR2_X1 U764 ( .A(KEYINPUT57), .B(n1069), .Z(n1072) );
XNOR2_X1 U765 ( .A(n1074), .B(n1075), .ZN(n1069) );
NOR2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U767 ( .A(n1078), .B(n1079), .Z(n1077) );
XNOR2_X1 U768 ( .A(KEYINPUT13), .B(n1080), .ZN(n1078) );
NOR3_X1 U769 ( .A1(n1081), .A2(KEYINPUT16), .A3(n1082), .ZN(n1080) );
AND2_X1 U770 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U771 ( .A(KEYINPUT32), .B(n1085), .Z(n1081) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1083), .ZN(n1085) );
NOR2_X1 U773 ( .A1(G898), .A2(n996), .ZN(n1076) );
NAND2_X1 U774 ( .A1(n996), .A2(n1029), .ZN(n1074) );
NOR2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(G66) );
XOR2_X1 U776 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1092), .ZN(G63) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR3_X1 U780 ( .A1(n1095), .A2(KEYINPUT22), .A3(n1096), .ZN(n1093) );
INV_X1 U781 ( .A(G478), .ZN(n1096) );
NOR2_X1 U782 ( .A1(n1086), .A2(n1097), .ZN(G60) );
XOR2_X1 U783 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U784 ( .A1(n1090), .A2(G475), .ZN(n1098) );
XOR2_X1 U785 ( .A(G104), .B(n1100), .Z(G6) );
NOR2_X1 U786 ( .A1(n1086), .A2(n1101), .ZN(G57) );
XOR2_X1 U787 ( .A(n1102), .B(n1103), .Z(n1101) );
XNOR2_X1 U788 ( .A(n1104), .B(n1105), .ZN(n1103) );
NAND2_X1 U789 ( .A1(KEYINPUT35), .A2(n1106), .ZN(n1105) );
NAND2_X1 U790 ( .A1(n1107), .A2(KEYINPUT34), .ZN(n1104) );
XOR2_X1 U791 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U792 ( .A(n1110), .B(n1111), .Z(n1102) );
NAND2_X1 U793 ( .A1(n1090), .A2(G472), .ZN(n1110) );
NOR2_X1 U794 ( .A1(n1086), .A2(n1112), .ZN(G54) );
XOR2_X1 U795 ( .A(n1113), .B(n1114), .Z(n1112) );
XOR2_X1 U796 ( .A(n1115), .B(n1062), .Z(n1114) );
XOR2_X1 U797 ( .A(n1116), .B(n1117), .Z(n1113) );
NOR2_X1 U798 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
XOR2_X1 U799 ( .A(n1120), .B(KEYINPUT18), .Z(n1119) );
NAND2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
NAND2_X1 U802 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NAND2_X1 U803 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U804 ( .A(KEYINPUT31), .B(n1127), .Z(n1123) );
NOR2_X1 U805 ( .A1(n1125), .A2(n1126), .ZN(n1127) );
XNOR2_X1 U806 ( .A(KEYINPUT48), .B(G110), .ZN(n1125) );
XNOR2_X1 U807 ( .A(KEYINPUT21), .B(n1128), .ZN(n1121) );
NAND2_X1 U808 ( .A1(n1090), .A2(G469), .ZN(n1116) );
NOR2_X1 U809 ( .A1(n1086), .A2(n1129), .ZN(G51) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR3_X1 U811 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NOR3_X1 U813 ( .A1(n1137), .A2(KEYINPUT45), .A3(n1138), .ZN(n1133) );
INV_X1 U814 ( .A(n1135), .ZN(n1138) );
NOR2_X1 U815 ( .A1(KEYINPUT5), .A2(n1139), .ZN(n1135) );
AND2_X1 U816 ( .A1(n1139), .A2(KEYINPUT45), .ZN(n1132) );
XOR2_X1 U817 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U818 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
OR2_X1 U819 ( .A1(n1144), .A2(KEYINPUT29), .ZN(n1143) );
NAND3_X1 U820 ( .A1(n1109), .A2(n1145), .A3(KEYINPUT29), .ZN(n1142) );
NAND2_X1 U821 ( .A1(n1090), .A2(n1045), .ZN(n1130) );
INV_X1 U822 ( .A(n1095), .ZN(n1090) );
NAND2_X1 U823 ( .A1(G902), .A2(n1146), .ZN(n1095) );
OR3_X1 U824 ( .A1(n992), .A2(n1029), .A3(n990), .ZN(n1146) );
NAND4_X1 U825 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n990) );
AND4_X1 U826 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
NAND4_X1 U827 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1029) );
NOR4_X1 U828 ( .A1(n1159), .A2(n1160), .A3(n985), .A4(n1100), .ZN(n1158) );
NOR3_X1 U829 ( .A1(n1023), .A2(n1161), .A3(n1026), .ZN(n1100) );
NOR3_X1 U830 ( .A1(n1023), .A2(n1161), .A3(n1027), .ZN(n985) );
INV_X1 U831 ( .A(n1008), .ZN(n1023) );
NOR2_X1 U832 ( .A1(n1162), .A2(n1163), .ZN(n1157) );
NOR2_X1 U833 ( .A1(n1164), .A2(n1016), .ZN(n1163) );
XOR2_X1 U834 ( .A(n1165), .B(KEYINPUT50), .Z(n1164) );
NOR3_X1 U835 ( .A1(n1013), .A2(n1166), .A3(n1161), .ZN(n1162) );
XOR2_X1 U836 ( .A(n1024), .B(KEYINPUT2), .Z(n1166) );
XNOR2_X1 U837 ( .A(n1066), .B(KEYINPUT27), .ZN(n992) );
NOR2_X1 U838 ( .A1(n996), .A2(G952), .ZN(n1086) );
XNOR2_X1 U839 ( .A(G146), .B(n1147), .ZN(G48) );
NAND3_X1 U840 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1147) );
XOR2_X1 U841 ( .A(n1170), .B(n1148), .Z(G45) );
NAND4_X1 U842 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1148) );
XOR2_X1 U843 ( .A(n1175), .B(n1039), .Z(n1171) );
XOR2_X1 U844 ( .A(n1126), .B(n1176), .Z(G42) );
NAND2_X1 U845 ( .A1(KEYINPUT37), .A2(n1177), .ZN(n1176) );
INV_X1 U846 ( .A(n1149), .ZN(n1177) );
NAND4_X1 U847 ( .A1(n1167), .A2(n1007), .A3(n1168), .A4(n1178), .ZN(n1149) );
XNOR2_X1 U848 ( .A(G137), .B(n1153), .ZN(G39) );
NAND4_X1 U849 ( .A1(n1167), .A2(n1001), .A3(n1179), .A4(n1007), .ZN(n1153) );
XNOR2_X1 U850 ( .A(G134), .B(n1152), .ZN(G36) );
NAND3_X1 U851 ( .A1(n1007), .A2(n1180), .A3(n1172), .ZN(n1152) );
XNOR2_X1 U852 ( .A(G131), .B(n1066), .ZN(G33) );
NAND3_X1 U853 ( .A1(n1007), .A2(n1168), .A3(n1172), .ZN(n1066) );
AND2_X1 U854 ( .A1(n1181), .A2(n1182), .ZN(n1172) );
NOR2_X1 U855 ( .A1(n1183), .A2(n1018), .ZN(n1007) );
INV_X1 U856 ( .A(n1184), .ZN(n1018) );
NAND2_X1 U857 ( .A1(n1185), .A2(n1186), .ZN(G30) );
NAND2_X1 U858 ( .A1(G128), .A2(n1154), .ZN(n1186) );
XOR2_X1 U859 ( .A(KEYINPUT20), .B(n1187), .Z(n1185) );
NOR2_X1 U860 ( .A1(G128), .A2(n1154), .ZN(n1187) );
NAND3_X1 U861 ( .A1(n1167), .A2(n1180), .A3(n1169), .ZN(n1154) );
AND2_X1 U862 ( .A1(n1181), .A2(n1038), .ZN(n1167) );
AND3_X1 U863 ( .A1(n1011), .A2(n1188), .A3(n1025), .ZN(n1181) );
XOR2_X1 U864 ( .A(G101), .B(n1189), .Z(G3) );
NOR3_X1 U865 ( .A1(n1024), .A2(n1161), .A3(n1013), .ZN(n1189) );
XNOR2_X1 U866 ( .A(n1151), .B(n1190), .ZN(G27) );
NOR2_X1 U867 ( .A1(KEYINPUT10), .A2(n1145), .ZN(n1190) );
NAND4_X1 U868 ( .A1(n1011), .A2(n1188), .A3(n1173), .A4(n1191), .ZN(n1151) );
NOR3_X1 U869 ( .A1(n1014), .A2(n1026), .A3(n1025), .ZN(n1191) );
NAND2_X1 U870 ( .A1(n1192), .A2(n1028), .ZN(n1188) );
NAND3_X1 U871 ( .A1(G902), .A2(n1193), .A3(n1056), .ZN(n1192) );
NOR2_X1 U872 ( .A1(n996), .A2(G900), .ZN(n1056) );
XOR2_X1 U873 ( .A(G122), .B(n1160), .Z(G24) );
AND3_X1 U874 ( .A1(n1008), .A2(n1173), .A3(n1194), .ZN(n1160) );
NOR3_X1 U875 ( .A1(n1195), .A2(n1196), .A3(n1197), .ZN(n1194) );
NOR2_X1 U876 ( .A1(n1198), .A2(n1175), .ZN(n1197) );
INV_X1 U877 ( .A(KEYINPUT11), .ZN(n1175) );
NOR2_X1 U878 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
NOR2_X1 U879 ( .A1(KEYINPUT11), .A2(n1168), .ZN(n1196) );
NOR2_X1 U880 ( .A1(n1038), .A2(n1179), .ZN(n1008) );
XNOR2_X1 U881 ( .A(G119), .B(n1155), .ZN(G21) );
NAND4_X1 U882 ( .A1(n1201), .A2(n1169), .A3(n1001), .A4(n1038), .ZN(n1155) );
INV_X1 U883 ( .A(n1024), .ZN(n1001) );
NOR2_X1 U884 ( .A1(n1178), .A2(n1016), .ZN(n1169) );
XOR2_X1 U885 ( .A(n1202), .B(n1203), .Z(G18) );
NOR2_X1 U886 ( .A1(KEYINPUT19), .A2(n1204), .ZN(n1203) );
INV_X1 U887 ( .A(G116), .ZN(n1204) );
NOR2_X1 U888 ( .A1(n1205), .A2(n1165), .ZN(n1202) );
NAND3_X1 U889 ( .A1(n1182), .A2(n1180), .A3(n1201), .ZN(n1165) );
INV_X1 U890 ( .A(n1027), .ZN(n1180) );
NAND2_X1 U891 ( .A1(n1200), .A2(n1039), .ZN(n1027) );
INV_X1 U892 ( .A(n1199), .ZN(n1039) );
XOR2_X1 U893 ( .A(n1016), .B(KEYINPUT33), .Z(n1205) );
XOR2_X1 U894 ( .A(n1206), .B(n1156), .Z(G15) );
NAND4_X1 U895 ( .A1(n1201), .A2(n1182), .A3(n1168), .A4(n1173), .ZN(n1156) );
INV_X1 U896 ( .A(n1026), .ZN(n1168) );
NAND2_X1 U897 ( .A1(n1199), .A2(n1174), .ZN(n1026) );
INV_X1 U898 ( .A(n1200), .ZN(n1174) );
INV_X1 U899 ( .A(n1013), .ZN(n1182) );
NAND2_X1 U900 ( .A1(n1179), .A2(n1207), .ZN(n1013) );
XOR2_X1 U901 ( .A(KEYINPUT49), .B(n1038), .Z(n1207) );
INV_X1 U902 ( .A(n1195), .ZN(n1201) );
NAND3_X1 U903 ( .A1(n1208), .A2(n1011), .A3(n1002), .ZN(n1195) );
INV_X1 U904 ( .A(n1025), .ZN(n1002) );
XOR2_X1 U905 ( .A(G110), .B(n1159), .Z(G12) );
NOR3_X1 U906 ( .A1(n1014), .A2(n1161), .A3(n1024), .ZN(n1159) );
NAND2_X1 U907 ( .A1(n1199), .A2(n1200), .ZN(n1024) );
XNOR2_X1 U908 ( .A(n1037), .B(KEYINPUT61), .ZN(n1200) );
XNOR2_X1 U909 ( .A(n1209), .B(G475), .ZN(n1037) );
NAND2_X1 U910 ( .A1(n1099), .A2(n1210), .ZN(n1209) );
XNOR2_X1 U911 ( .A(n1211), .B(n1212), .ZN(n1099) );
XOR2_X1 U912 ( .A(n1213), .B(n1214), .Z(n1212) );
XOR2_X1 U913 ( .A(G122), .B(G113), .Z(n1214) );
XOR2_X1 U914 ( .A(G146), .B(G131), .Z(n1213) );
XOR2_X1 U915 ( .A(n1215), .B(n1058), .Z(n1211) );
XNOR2_X1 U916 ( .A(G104), .B(n1216), .ZN(n1215) );
NOR2_X1 U917 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U918 ( .A(n1219), .B(KEYINPUT6), .Z(n1218) );
NAND2_X1 U919 ( .A1(n1170), .A2(n1220), .ZN(n1219) );
NOR2_X1 U920 ( .A1(n1170), .A2(n1220), .ZN(n1217) );
NAND3_X1 U921 ( .A1(n1221), .A2(n996), .A3(G214), .ZN(n1220) );
XOR2_X1 U922 ( .A(n1222), .B(G478), .Z(n1199) );
OR2_X1 U923 ( .A1(n1094), .A2(G902), .ZN(n1222) );
XNOR2_X1 U924 ( .A(n1223), .B(n1224), .ZN(n1094) );
XOR2_X1 U925 ( .A(n1225), .B(n1226), .Z(n1224) );
AND2_X1 U926 ( .A1(n1227), .A2(G217), .ZN(n1226) );
NOR2_X1 U927 ( .A1(KEYINPUT24), .A2(n1228), .ZN(n1225) );
XOR2_X1 U928 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U929 ( .A(G116), .B(G107), .Z(n1230) );
NOR2_X1 U930 ( .A1(KEYINPUT4), .A2(n1231), .ZN(n1229) );
XOR2_X1 U931 ( .A(KEYINPUT9), .B(G122), .Z(n1231) );
XOR2_X1 U932 ( .A(n1232), .B(n1233), .Z(n1223) );
NOR2_X1 U933 ( .A1(KEYINPUT47), .A2(G128), .ZN(n1233) );
XOR2_X1 U934 ( .A(G134), .B(n1170), .Z(n1232) );
NAND4_X1 U935 ( .A1(n1173), .A2(n1025), .A3(n1208), .A4(n1011), .ZN(n1161) );
NAND2_X1 U936 ( .A1(G221), .A2(n1234), .ZN(n1011) );
NAND2_X1 U937 ( .A1(n1028), .A2(n1235), .ZN(n1208) );
NAND4_X1 U938 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1237), .ZN(n1235) );
INV_X1 U939 ( .A(G898), .ZN(n1237) );
XNOR2_X1 U940 ( .A(KEYINPUT55), .B(n1193), .ZN(n1236) );
NAND3_X1 U941 ( .A1(n1193), .A2(n996), .A3(G952), .ZN(n1028) );
NAND2_X1 U942 ( .A1(G237), .A2(G234), .ZN(n1193) );
NAND3_X1 U943 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1025) );
INV_X1 U944 ( .A(n1042), .ZN(n1240) );
NOR2_X1 U945 ( .A1(n1044), .A2(n1043), .ZN(n1042) );
NAND3_X1 U946 ( .A1(n1043), .A2(n1044), .A3(n1241), .ZN(n1239) );
NAND2_X1 U947 ( .A1(n1242), .A2(n1210), .ZN(n1044) );
XOR2_X1 U948 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U949 ( .A(n1128), .B(n1245), .Z(n1244) );
AND2_X1 U950 ( .A1(G227), .A2(n996), .ZN(n1128) );
XOR2_X1 U951 ( .A(n1246), .B(n1247), .Z(n1243) );
NOR2_X1 U952 ( .A1(KEYINPUT58), .A2(n1115), .ZN(n1247) );
XNOR2_X1 U953 ( .A(n1248), .B(n1249), .ZN(n1115) );
XOR2_X1 U954 ( .A(G101), .B(n1109), .Z(n1249) );
XOR2_X1 U955 ( .A(G104), .B(n986), .Z(n1248) );
INV_X1 U956 ( .A(G107), .ZN(n986) );
XOR2_X1 U957 ( .A(n1126), .B(G110), .Z(n1246) );
INV_X1 U958 ( .A(G140), .ZN(n1126) );
OR2_X1 U959 ( .A1(n1241), .A2(n1043), .ZN(n1238) );
XNOR2_X1 U960 ( .A(G469), .B(KEYINPUT43), .ZN(n1043) );
INV_X1 U961 ( .A(KEYINPUT38), .ZN(n1241) );
INV_X1 U962 ( .A(n1016), .ZN(n1173) );
NAND2_X1 U963 ( .A1(n1250), .A2(n1184), .ZN(n1016) );
NAND2_X1 U964 ( .A1(G214), .A2(n1251), .ZN(n1184) );
XOR2_X1 U965 ( .A(KEYINPUT14), .B(n1183), .Z(n1250) );
INV_X1 U966 ( .A(n1019), .ZN(n1183) );
XOR2_X1 U967 ( .A(n1252), .B(n1045), .Z(n1019) );
AND2_X1 U968 ( .A1(G210), .A2(n1251), .ZN(n1045) );
NAND2_X1 U969 ( .A1(n1221), .A2(n1210), .ZN(n1251) );
XNOR2_X1 U970 ( .A(n1047), .B(KEYINPUT12), .ZN(n1252) );
AND2_X1 U971 ( .A1(n1253), .A2(n1210), .ZN(n1047) );
XOR2_X1 U972 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U973 ( .A(n1137), .B(n1144), .Z(n1255) );
XOR2_X1 U974 ( .A(n1145), .B(n1060), .Z(n1144) );
INV_X1 U975 ( .A(n1136), .ZN(n1137) );
XOR2_X1 U976 ( .A(n1256), .B(n1257), .Z(n1136) );
XNOR2_X1 U977 ( .A(n1084), .B(n1079), .ZN(n1257) );
XOR2_X1 U978 ( .A(G110), .B(n1258), .Z(n1079) );
XOR2_X1 U979 ( .A(KEYINPUT0), .B(G122), .Z(n1258) );
XOR2_X1 U980 ( .A(n1259), .B(n1260), .Z(n1084) );
XOR2_X1 U981 ( .A(G107), .B(n1261), .Z(n1260) );
NOR2_X1 U982 ( .A1(G104), .A2(KEYINPUT15), .ZN(n1261) );
NAND2_X1 U983 ( .A1(KEYINPUT60), .A2(n1106), .ZN(n1259) );
XOR2_X1 U984 ( .A(n1083), .B(KEYINPUT17), .Z(n1256) );
NAND2_X1 U985 ( .A1(n1262), .A2(n1263), .ZN(n1083) );
NAND2_X1 U986 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U987 ( .A(KEYINPUT3), .B(n1266), .Z(n1265) );
XOR2_X1 U988 ( .A(KEYINPUT56), .B(G113), .Z(n1264) );
XOR2_X1 U989 ( .A(n1267), .B(KEYINPUT53), .Z(n1262) );
NAND2_X1 U990 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U991 ( .A(KEYINPUT3), .B(n1266), .ZN(n1269) );
XOR2_X1 U992 ( .A(KEYINPUT56), .B(n1206), .Z(n1268) );
XOR2_X1 U993 ( .A(KEYINPUT1), .B(n1141), .Z(n1254) );
NOR2_X1 U994 ( .A1(n1071), .A2(G953), .ZN(n1141) );
INV_X1 U995 ( .A(G224), .ZN(n1071) );
NAND2_X1 U996 ( .A1(n1038), .A2(n1178), .ZN(n1014) );
INV_X1 U997 ( .A(n1179), .ZN(n1178) );
XOR2_X1 U998 ( .A(n1270), .B(G472), .Z(n1179) );
NAND2_X1 U999 ( .A1(KEYINPUT40), .A2(n1040), .ZN(n1270) );
NAND2_X1 U1000 ( .A1(n1271), .A2(n1210), .ZN(n1040) );
XOR2_X1 U1001 ( .A(n1272), .B(KEYINPUT44), .Z(n1271) );
NAND2_X1 U1002 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
OR2_X1 U1003 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
XOR2_X1 U1004 ( .A(n1277), .B(KEYINPUT52), .Z(n1273) );
NAND2_X1 U1005 ( .A1(n1276), .A2(n1275), .ZN(n1277) );
XNOR2_X1 U1006 ( .A(n1278), .B(n1279), .ZN(n1275) );
INV_X1 U1007 ( .A(n1108), .ZN(n1279) );
XOR2_X1 U1008 ( .A(n1280), .B(n1245), .Z(n1108) );
INV_X1 U1009 ( .A(n1062), .ZN(n1245) );
XNOR2_X1 U1010 ( .A(G131), .B(n1281), .ZN(n1062) );
XOR2_X1 U1011 ( .A(G137), .B(G134), .Z(n1281) );
NAND2_X1 U1012 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
NAND2_X1 U1013 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U1014 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U1015 ( .A1(KEYINPUT59), .A2(n1206), .ZN(n1287) );
INV_X1 U1016 ( .A(G113), .ZN(n1206) );
INV_X1 U1017 ( .A(KEYINPUT41), .ZN(n1286) );
NAND2_X1 U1018 ( .A1(G113), .A2(n1288), .ZN(n1282) );
NAND2_X1 U1019 ( .A1(KEYINPUT59), .A2(n1289), .ZN(n1288) );
OR2_X1 U1020 ( .A1(n1284), .A2(KEYINPUT41), .ZN(n1289) );
XNOR2_X1 U1021 ( .A(n1266), .B(KEYINPUT23), .ZN(n1284) );
XOR2_X1 U1022 ( .A(G116), .B(G119), .Z(n1266) );
NAND2_X1 U1023 ( .A1(n1290), .A2(n1291), .ZN(n1278) );
XOR2_X1 U1024 ( .A(KEYINPUT54), .B(n1109), .Z(n1291) );
INV_X1 U1025 ( .A(n1060), .ZN(n1109) );
XOR2_X1 U1026 ( .A(n1170), .B(n1292), .Z(n1060) );
INV_X1 U1027 ( .A(G143), .ZN(n1170) );
XNOR2_X1 U1028 ( .A(KEYINPUT62), .B(KEYINPUT42), .ZN(n1290) );
XNOR2_X1 U1029 ( .A(n1293), .B(n1111), .ZN(n1276) );
AND3_X1 U1030 ( .A1(n1221), .A2(n996), .A3(G210), .ZN(n1111) );
INV_X1 U1031 ( .A(G237), .ZN(n1221) );
NAND2_X1 U1032 ( .A1(KEYINPUT51), .A2(n1106), .ZN(n1293) );
INV_X1 U1033 ( .A(G101), .ZN(n1106) );
XNOR2_X1 U1034 ( .A(n1294), .B(n1091), .ZN(n1038) );
AND2_X1 U1035 ( .A1(G217), .A2(n1234), .ZN(n1091) );
NAND2_X1 U1036 ( .A1(G234), .A2(n1210), .ZN(n1234) );
NAND2_X1 U1037 ( .A1(n1089), .A2(n1210), .ZN(n1294) );
INV_X1 U1038 ( .A(G902), .ZN(n1210) );
XNOR2_X1 U1039 ( .A(n1295), .B(n1296), .ZN(n1089) );
XOR2_X1 U1040 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1041 ( .A(G119), .B(G110), .Z(n1298) );
XOR2_X1 U1042 ( .A(KEYINPUT36), .B(G137), .Z(n1297) );
XOR2_X1 U1043 ( .A(n1299), .B(n1058), .Z(n1295) );
XNOR2_X1 U1044 ( .A(n1145), .B(G140), .ZN(n1058) );
INV_X1 U1045 ( .A(G125), .ZN(n1145) );
XOR2_X1 U1046 ( .A(n1300), .B(n1292), .Z(n1299) );
XOR2_X1 U1047 ( .A(G146), .B(G128), .Z(n1292) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1227), .ZN(n1300) );
AND2_X1 U1049 ( .A1(G234), .A2(n996), .ZN(n1227) );
INV_X1 U1050 ( .A(G953), .ZN(n996) );
endmodule


