//Key = 0111001010110011101111100010100010010001011101000101110011101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370;

XNOR2_X1 U757 ( .A(G107), .B(n1040), .ZN(G9) );
NOR2_X1 U758 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U759 ( .A1(n1043), .A2(n1044), .A3(G953), .A4(n1045), .ZN(n1042) );
NOR3_X1 U760 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1044) );
NAND2_X1 U761 ( .A1(n1049), .A2(n1050), .ZN(n1043) );
NAND3_X1 U762 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NAND2_X1 U763 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NAND2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XNOR2_X1 U765 ( .A(n1058), .B(KEYINPUT28), .ZN(n1056) );
NAND4_X1 U766 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1051) );
NAND2_X1 U767 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NAND3_X1 U768 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND2_X1 U769 ( .A1(KEYINPUT1), .A2(n1068), .ZN(n1067) );
NAND2_X1 U770 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
NAND2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U772 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1065) );
XNOR2_X1 U774 ( .A(KEYINPUT29), .B(n1077), .ZN(n1076) );
NAND2_X1 U775 ( .A1(n1057), .A2(n1078), .ZN(n1060) );
NAND2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U777 ( .A(n1046), .ZN(n1057) );
NAND3_X1 U778 ( .A1(n1069), .A2(n1081), .A3(n1082), .ZN(n1046) );
NAND2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1059) );
INV_X1 U780 ( .A(KEYINPUT1), .ZN(n1084) );
NAND2_X1 U781 ( .A1(n1063), .A2(n1068), .ZN(n1083) );
AND2_X1 U782 ( .A1(n1058), .A2(n1081), .ZN(n1063) );
NOR3_X1 U783 ( .A1(n1045), .A2(G953), .A3(G952), .ZN(n1041) );
AND4_X1 U784 ( .A1(n1085), .A2(n1082), .A3(n1086), .A4(n1087), .ZN(n1045) );
NOR4_X1 U785 ( .A1(n1088), .A2(n1054), .A3(n1089), .A4(n1090), .ZN(n1087) );
XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U787 ( .A1(KEYINPUT60), .A2(n1093), .ZN(n1091) );
NOR2_X1 U788 ( .A1(n1094), .A2(n1095), .ZN(n1089) );
XNOR2_X1 U789 ( .A(n1096), .B(KEYINPUT4), .ZN(n1095) );
INV_X1 U790 ( .A(n1097), .ZN(n1088) );
NOR2_X1 U791 ( .A1(n1098), .A2(n1099), .ZN(n1086) );
XOR2_X1 U792 ( .A(n1100), .B(n1101), .Z(G72) );
XOR2_X1 U793 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U794 ( .A1(n1104), .A2(KEYINPUT17), .ZN(n1103) );
AND2_X1 U795 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NOR2_X1 U796 ( .A1(n1107), .A2(n1108), .ZN(n1102) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1108) );
XNOR2_X1 U798 ( .A(G131), .B(n1111), .ZN(n1110) );
NAND3_X1 U799 ( .A1(n1112), .A2(n1113), .A3(KEYINPUT8), .ZN(n1111) );
OR2_X1 U800 ( .A1(n1114), .A2(KEYINPUT23), .ZN(n1113) );
NAND3_X1 U801 ( .A1(G134), .A2(n1115), .A3(KEYINPUT23), .ZN(n1112) );
XOR2_X1 U802 ( .A(n1116), .B(n1117), .Z(n1109) );
NAND2_X1 U803 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NAND2_X1 U804 ( .A1(G125), .A2(n1120), .ZN(n1119) );
XOR2_X1 U805 ( .A(KEYINPUT3), .B(n1121), .Z(n1118) );
NOR2_X1 U806 ( .A1(G125), .A2(n1120), .ZN(n1121) );
NOR2_X1 U807 ( .A1(G900), .A2(n1105), .ZN(n1107) );
NAND2_X1 U808 ( .A1(G953), .A2(n1122), .ZN(n1100) );
NAND2_X1 U809 ( .A1(G900), .A2(G227), .ZN(n1122) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(G69) );
XOR2_X1 U811 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U813 ( .A1(G898), .A2(n1129), .ZN(n1127) );
XNOR2_X1 U814 ( .A(G953), .B(KEYINPUT37), .ZN(n1129) );
NAND2_X1 U815 ( .A1(n1105), .A2(n1130), .ZN(n1125) );
NAND2_X1 U816 ( .A1(G953), .A2(n1131), .ZN(n1123) );
NAND2_X1 U817 ( .A1(G224), .A2(G898), .ZN(n1131) );
NOR2_X1 U818 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XOR2_X1 U819 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U820 ( .A(n1136), .B(KEYINPUT10), .Z(n1135) );
NAND2_X1 U821 ( .A1(n1137), .A2(n1096), .ZN(n1136) );
INV_X1 U822 ( .A(n1138), .ZN(n1096) );
XNOR2_X1 U823 ( .A(n1139), .B(KEYINPUT6), .ZN(n1132) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1140), .ZN(G63) );
NOR3_X1 U825 ( .A1(n1092), .A2(n1141), .A3(n1142), .ZN(n1140) );
AND4_X1 U826 ( .A1(n1143), .A2(n1137), .A3(n1144), .A4(G478), .ZN(n1142) );
INV_X1 U827 ( .A(KEYINPUT61), .ZN(n1144) );
NOR2_X1 U828 ( .A1(n1145), .A2(n1143), .ZN(n1141) );
NOR3_X1 U829 ( .A1(n1093), .A2(KEYINPUT61), .A3(n1049), .ZN(n1145) );
INV_X1 U830 ( .A(G478), .ZN(n1093) );
NOR2_X1 U831 ( .A1(n1139), .A2(n1146), .ZN(G60) );
XOR2_X1 U832 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND2_X1 U833 ( .A1(n1137), .A2(G475), .ZN(n1148) );
XOR2_X1 U834 ( .A(n1149), .B(n1150), .Z(G6) );
NAND2_X1 U835 ( .A1(KEYINPUT32), .A2(n1151), .ZN(n1149) );
NOR2_X1 U836 ( .A1(n1139), .A2(n1152), .ZN(G57) );
XNOR2_X1 U837 ( .A(n1153), .B(n1154), .ZN(n1152) );
XOR2_X1 U838 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U839 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U840 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U841 ( .A1(KEYINPUT30), .A2(n1161), .ZN(n1159) );
NOR2_X1 U842 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NOR2_X1 U843 ( .A1(n1164), .A2(n1165), .ZN(n1157) );
NOR2_X1 U844 ( .A1(n1166), .A2(n1163), .ZN(n1164) );
INV_X1 U845 ( .A(KEYINPUT22), .ZN(n1163) );
NOR2_X1 U846 ( .A1(KEYINPUT30), .A2(n1167), .ZN(n1166) );
NAND2_X1 U847 ( .A1(n1137), .A2(G472), .ZN(n1155) );
NOR2_X1 U848 ( .A1(n1139), .A2(n1168), .ZN(G54) );
XOR2_X1 U849 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U850 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U851 ( .A(n1173), .B(n1174), .ZN(n1169) );
NAND2_X1 U852 ( .A1(n1137), .A2(G469), .ZN(n1173) );
NOR2_X1 U853 ( .A1(n1139), .A2(n1175), .ZN(G51) );
XOR2_X1 U854 ( .A(n1128), .B(n1176), .Z(n1175) );
XOR2_X1 U855 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U856 ( .A1(n1137), .A2(G210), .ZN(n1178) );
NOR2_X1 U857 ( .A1(n1179), .A2(n1049), .ZN(n1137) );
NOR2_X1 U858 ( .A1(n1106), .A2(n1130), .ZN(n1049) );
NAND4_X1 U859 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1130) );
NOR4_X1 U860 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
INV_X1 U861 ( .A(n1040), .ZN(n1187) );
NAND3_X1 U862 ( .A1(n1188), .A2(n1069), .A3(n1189), .ZN(n1040) );
NOR2_X1 U863 ( .A1(n1150), .A2(n1190), .ZN(n1182) );
NOR4_X1 U864 ( .A1(n1191), .A2(n1192), .A3(n1077), .A4(n1079), .ZN(n1190) );
XNOR2_X1 U865 ( .A(n1193), .B(KEYINPUT12), .ZN(n1191) );
AND3_X1 U866 ( .A1(n1189), .A2(n1069), .A3(n1194), .ZN(n1150) );
NAND3_X1 U867 ( .A1(n1189), .A2(n1195), .A3(n1075), .ZN(n1181) );
XNOR2_X1 U868 ( .A(KEYINPUT36), .B(n1048), .ZN(n1195) );
NAND2_X1 U869 ( .A1(n1196), .A2(n1197), .ZN(n1180) );
XOR2_X1 U870 ( .A(n1198), .B(KEYINPUT42), .Z(n1196) );
NAND4_X1 U871 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1106) );
NOR4_X1 U872 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
NAND2_X1 U873 ( .A1(n1207), .A2(n1208), .ZN(n1201) );
NAND2_X1 U874 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U875 ( .A1(n1211), .A2(n1058), .ZN(n1210) );
XNOR2_X1 U876 ( .A(n1212), .B(KEYINPUT16), .ZN(n1211) );
NAND2_X1 U877 ( .A1(n1075), .A2(n1194), .ZN(n1209) );
INV_X1 U878 ( .A(n1213), .ZN(n1207) );
NAND2_X1 U879 ( .A1(n1214), .A2(KEYINPUT11), .ZN(n1177) );
XOR2_X1 U880 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U881 ( .A(n1217), .B(n1218), .ZN(n1216) );
NOR2_X1 U882 ( .A1(n1105), .A2(G952), .ZN(n1139) );
XNOR2_X1 U883 ( .A(G146), .B(n1199), .ZN(G48) );
NAND3_X1 U884 ( .A1(n1219), .A2(n1194), .A3(n1212), .ZN(n1199) );
NAND2_X1 U885 ( .A1(n1220), .A2(n1221), .ZN(G45) );
NAND2_X1 U886 ( .A1(n1222), .A2(n1200), .ZN(n1221) );
NAND2_X1 U887 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NAND2_X1 U888 ( .A1(KEYINPUT48), .A2(n1225), .ZN(n1224) );
NAND3_X1 U889 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1220) );
INV_X1 U890 ( .A(KEYINPUT48), .ZN(n1228) );
NAND2_X1 U891 ( .A1(G143), .A2(n1225), .ZN(n1227) );
INV_X1 U892 ( .A(KEYINPUT38), .ZN(n1225) );
NAND2_X1 U893 ( .A1(n1229), .A2(n1223), .ZN(n1226) );
OR2_X1 U894 ( .A1(n1200), .A2(KEYINPUT38), .ZN(n1229) );
NAND4_X1 U895 ( .A1(n1193), .A2(n1219), .A3(n1230), .A4(n1231), .ZN(n1200) );
XNOR2_X1 U896 ( .A(n1120), .B(n1232), .ZN(G42) );
NOR4_X1 U897 ( .A1(KEYINPUT25), .A2(n1079), .A3(n1233), .A4(n1213), .ZN(n1232) );
XNOR2_X1 U898 ( .A(n1115), .B(n1234), .ZN(G39) );
NOR2_X1 U899 ( .A1(n1213), .A2(n1235), .ZN(n1234) );
XNOR2_X1 U900 ( .A(n1236), .B(n1206), .ZN(G36) );
NOR3_X1 U901 ( .A1(n1237), .A2(n1080), .A3(n1213), .ZN(n1206) );
XNOR2_X1 U902 ( .A(n1238), .B(n1205), .ZN(G33) );
NOR3_X1 U903 ( .A1(n1237), .A2(n1079), .A3(n1213), .ZN(n1205) );
NAND4_X1 U904 ( .A1(n1053), .A2(n1239), .A3(n1062), .A4(n1240), .ZN(n1213) );
XNOR2_X1 U905 ( .A(n1085), .B(KEYINPUT14), .ZN(n1053) );
XNOR2_X1 U906 ( .A(n1204), .B(n1241), .ZN(G30) );
NOR2_X1 U907 ( .A1(G128), .A2(KEYINPUT59), .ZN(n1241) );
AND3_X1 U908 ( .A1(n1219), .A2(n1188), .A3(n1212), .ZN(n1204) );
INV_X1 U909 ( .A(n1080), .ZN(n1188) );
NOR3_X1 U910 ( .A1(n1047), .A2(n1242), .A3(n1071), .ZN(n1219) );
XNOR2_X1 U911 ( .A(n1243), .B(n1186), .ZN(G3) );
NOR3_X1 U912 ( .A1(n1237), .A2(n1244), .A3(n1048), .ZN(n1186) );
XNOR2_X1 U913 ( .A(n1203), .B(n1245), .ZN(G27) );
XNOR2_X1 U914 ( .A(G125), .B(KEYINPUT40), .ZN(n1245) );
AND3_X1 U915 ( .A1(n1075), .A2(n1194), .A3(n1246), .ZN(n1203) );
NOR3_X1 U916 ( .A1(n1077), .A2(n1242), .A3(n1047), .ZN(n1246) );
INV_X1 U917 ( .A(n1240), .ZN(n1242) );
NAND2_X1 U918 ( .A1(n1247), .A2(n1248), .ZN(n1240) );
NAND3_X1 U919 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1247) );
INV_X1 U920 ( .A(G900), .ZN(n1250) );
XNOR2_X1 U921 ( .A(KEYINPUT47), .B(n1179), .ZN(n1249) );
NAND2_X1 U922 ( .A1(n1252), .A2(n1253), .ZN(G24) );
NAND2_X1 U923 ( .A1(n1185), .A2(n1254), .ZN(n1253) );
XOR2_X1 U924 ( .A(KEYINPUT49), .B(n1255), .Z(n1252) );
NOR2_X1 U925 ( .A1(n1185), .A2(n1254), .ZN(n1255) );
INV_X1 U926 ( .A(G122), .ZN(n1254) );
AND4_X1 U927 ( .A1(n1082), .A2(n1069), .A3(n1256), .A4(n1230), .ZN(n1185) );
NOR2_X1 U928 ( .A1(n1257), .A2(n1192), .ZN(n1256) );
INV_X1 U929 ( .A(n1231), .ZN(n1257) );
NOR2_X1 U930 ( .A1(n1258), .A2(n1098), .ZN(n1069) );
XNOR2_X1 U931 ( .A(n1259), .B(n1260), .ZN(G21) );
NOR2_X1 U932 ( .A1(n1047), .A2(n1198), .ZN(n1260) );
NAND3_X1 U933 ( .A1(n1082), .A2(n1261), .A3(n1262), .ZN(n1198) );
INV_X1 U934 ( .A(n1235), .ZN(n1262) );
NAND2_X1 U935 ( .A1(n1058), .A2(n1212), .ZN(n1235) );
NOR2_X1 U936 ( .A1(n1263), .A2(n1264), .ZN(n1212) );
INV_X1 U937 ( .A(n1048), .ZN(n1058) );
INV_X1 U938 ( .A(n1077), .ZN(n1082) );
XOR2_X1 U939 ( .A(G116), .B(n1184), .Z(G18) );
NOR3_X1 U940 ( .A1(n1080), .A2(n1192), .A3(n1265), .ZN(n1184) );
INV_X1 U941 ( .A(n1068), .ZN(n1265) );
NAND2_X1 U942 ( .A1(n1266), .A2(n1230), .ZN(n1080) );
XOR2_X1 U943 ( .A(n1267), .B(KEYINPUT2), .Z(n1230) );
XOR2_X1 U944 ( .A(G113), .B(n1268), .Z(G15) );
NOR2_X1 U945 ( .A1(n1269), .A2(n1047), .ZN(n1268) );
INV_X1 U946 ( .A(n1197), .ZN(n1047) );
XOR2_X1 U947 ( .A(n1270), .B(KEYINPUT54), .Z(n1269) );
NAND3_X1 U948 ( .A1(n1194), .A2(n1261), .A3(n1068), .ZN(n1270) );
NOR2_X1 U949 ( .A1(n1237), .A2(n1077), .ZN(n1068) );
NAND2_X1 U950 ( .A1(n1074), .A2(n1271), .ZN(n1077) );
INV_X1 U951 ( .A(n1193), .ZN(n1237) );
NOR2_X1 U952 ( .A1(n1258), .A2(n1263), .ZN(n1193) );
INV_X1 U953 ( .A(n1098), .ZN(n1263) );
INV_X1 U954 ( .A(n1079), .ZN(n1194) );
NAND2_X1 U955 ( .A1(n1267), .A2(n1231), .ZN(n1079) );
XOR2_X1 U956 ( .A(n1099), .B(KEYINPUT63), .Z(n1231) );
XNOR2_X1 U957 ( .A(n1272), .B(n1273), .ZN(G12) );
NOR3_X1 U958 ( .A1(n1048), .A2(n1244), .A3(n1233), .ZN(n1273) );
INV_X1 U959 ( .A(n1075), .ZN(n1233) );
NOR2_X1 U960 ( .A1(n1098), .A2(n1264), .ZN(n1075) );
INV_X1 U961 ( .A(n1258), .ZN(n1264) );
NAND2_X1 U962 ( .A1(n1274), .A2(n1097), .ZN(n1258) );
NAND2_X1 U963 ( .A1(n1094), .A2(n1138), .ZN(n1097) );
OR2_X1 U964 ( .A1(n1138), .A2(n1094), .ZN(n1274) );
NOR2_X1 U965 ( .A1(n1134), .A2(G902), .ZN(n1094) );
XOR2_X1 U966 ( .A(n1275), .B(n1276), .Z(n1134) );
XNOR2_X1 U967 ( .A(n1115), .B(n1277), .ZN(n1276) );
NOR2_X1 U968 ( .A1(KEYINPUT50), .A2(n1278), .ZN(n1277) );
XOR2_X1 U969 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U970 ( .A(n1281), .B(n1282), .Z(n1280) );
NAND2_X1 U971 ( .A1(KEYINPUT62), .A2(n1272), .ZN(n1282) );
NAND2_X1 U972 ( .A1(KEYINPUT39), .A2(n1259), .ZN(n1281) );
XOR2_X1 U973 ( .A(G128), .B(n1283), .Z(n1279) );
NOR2_X1 U974 ( .A1(KEYINPUT7), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U975 ( .A(n1285), .B(n1286), .ZN(n1284) );
NOR2_X1 U976 ( .A1(G146), .A2(KEYINPUT34), .ZN(n1286) );
NAND2_X1 U977 ( .A1(n1287), .A2(G221), .ZN(n1275) );
NAND2_X1 U978 ( .A1(G217), .A2(n1288), .ZN(n1138) );
XNOR2_X1 U979 ( .A(n1289), .B(G472), .ZN(n1098) );
NAND2_X1 U980 ( .A1(n1290), .A2(n1179), .ZN(n1289) );
XNOR2_X1 U981 ( .A(n1291), .B(n1292), .ZN(n1290) );
INV_X1 U982 ( .A(n1153), .ZN(n1292) );
XOR2_X1 U983 ( .A(n1293), .B(n1243), .Z(n1153) );
INV_X1 U984 ( .A(G101), .ZN(n1243) );
NAND2_X1 U985 ( .A1(n1294), .A2(G210), .ZN(n1293) );
XOR2_X1 U986 ( .A(n1295), .B(KEYINPUT41), .Z(n1291) );
NAND2_X1 U987 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U988 ( .A1(n1165), .A2(n1160), .ZN(n1297) );
INV_X1 U989 ( .A(n1167), .ZN(n1160) );
INV_X1 U990 ( .A(n1162), .ZN(n1165) );
XOR2_X1 U991 ( .A(n1298), .B(KEYINPUT46), .Z(n1296) );
NAND2_X1 U992 ( .A1(n1167), .A2(n1162), .ZN(n1298) );
XOR2_X1 U993 ( .A(n1215), .B(n1299), .Z(n1162) );
INV_X1 U994 ( .A(n1300), .ZN(n1299) );
XNOR2_X1 U995 ( .A(n1301), .B(KEYINPUT20), .ZN(n1167) );
NAND2_X1 U996 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
NAND2_X1 U997 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
INV_X1 U998 ( .A(KEYINPUT0), .ZN(n1305) );
XOR2_X1 U999 ( .A(G113), .B(n1306), .Z(n1304) );
NAND3_X1 U1000 ( .A1(G113), .A2(n1306), .A3(KEYINPUT0), .ZN(n1302) );
INV_X1 U1001 ( .A(n1189), .ZN(n1244) );
NOR2_X1 U1002 ( .A1(n1071), .A2(n1192), .ZN(n1189) );
NAND2_X1 U1003 ( .A1(n1197), .A2(n1261), .ZN(n1192) );
NAND2_X1 U1004 ( .A1(n1248), .A2(n1307), .ZN(n1261) );
NAND3_X1 U1005 ( .A1(n1251), .A2(n1308), .A3(G902), .ZN(n1307) );
XOR2_X1 U1006 ( .A(KEYINPUT53), .B(G898), .Z(n1308) );
AND2_X1 U1007 ( .A1(G953), .A2(n1309), .ZN(n1251) );
NAND2_X1 U1008 ( .A1(n1310), .A2(n1081), .ZN(n1248) );
AND2_X1 U1009 ( .A1(n1311), .A2(n1309), .ZN(n1081) );
NAND2_X1 U1010 ( .A1(G237), .A2(G234), .ZN(n1309) );
XOR2_X1 U1011 ( .A(KEYINPUT24), .B(G952), .Z(n1311) );
XNOR2_X1 U1012 ( .A(G953), .B(KEYINPUT13), .ZN(n1310) );
NOR2_X1 U1013 ( .A1(n1054), .A2(n1085), .ZN(n1197) );
AND3_X1 U1014 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1085) );
OR2_X1 U1015 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND3_X1 U1016 ( .A1(n1316), .A2(n1315), .A3(n1179), .ZN(n1313) );
NAND2_X1 U1017 ( .A1(G210), .A2(G237), .ZN(n1315) );
XNOR2_X1 U1018 ( .A(n1317), .B(n1318), .ZN(n1316) );
XOR2_X1 U1019 ( .A(n1218), .B(n1319), .Z(n1318) );
XNOR2_X1 U1020 ( .A(KEYINPUT15), .B(n1217), .ZN(n1319) );
AND2_X1 U1021 ( .A1(G224), .A2(n1105), .ZN(n1218) );
XOR2_X1 U1022 ( .A(n1320), .B(n1128), .Z(n1317) );
XNOR2_X1 U1023 ( .A(n1321), .B(n1322), .ZN(n1128) );
XOR2_X1 U1024 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1025 ( .A(n1306), .B(n1325), .Z(n1324) );
XNOR2_X1 U1026 ( .A(G116), .B(n1259), .ZN(n1306) );
INV_X1 U1027 ( .A(G119), .ZN(n1259) );
XOR2_X1 U1028 ( .A(n1326), .B(n1327), .Z(n1321) );
XNOR2_X1 U1029 ( .A(KEYINPUT44), .B(n1272), .ZN(n1327) );
XNOR2_X1 U1030 ( .A(KEYINPUT9), .B(KEYINPUT57), .ZN(n1326) );
NAND2_X1 U1031 ( .A1(KEYINPUT52), .A2(n1215), .ZN(n1320) );
XNOR2_X1 U1032 ( .A(G146), .B(n1328), .ZN(n1215) );
INV_X1 U1033 ( .A(n1329), .ZN(n1328) );
NAND2_X1 U1034 ( .A1(G210), .A2(G902), .ZN(n1312) );
INV_X1 U1035 ( .A(n1062), .ZN(n1054) );
NAND2_X1 U1036 ( .A1(G214), .A2(n1330), .ZN(n1062) );
OR2_X1 U1037 ( .A1(G237), .A2(G902), .ZN(n1330) );
INV_X1 U1038 ( .A(n1239), .ZN(n1071) );
NOR2_X1 U1039 ( .A1(n1074), .A2(n1073), .ZN(n1239) );
INV_X1 U1040 ( .A(n1271), .ZN(n1073) );
NAND2_X1 U1041 ( .A1(G221), .A2(n1288), .ZN(n1271) );
NAND2_X1 U1042 ( .A1(G234), .A2(n1179), .ZN(n1288) );
XOR2_X1 U1043 ( .A(n1331), .B(G469), .Z(n1074) );
NAND2_X1 U1044 ( .A1(n1332), .A2(n1179), .ZN(n1331) );
XOR2_X1 U1045 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1046 ( .A(n1172), .B(KEYINPUT27), .ZN(n1334) );
XNOR2_X1 U1047 ( .A(n1335), .B(n1336), .ZN(n1172) );
XNOR2_X1 U1048 ( .A(n1120), .B(G110), .ZN(n1336) );
INV_X1 U1049 ( .A(G140), .ZN(n1120) );
NAND2_X1 U1050 ( .A1(G227), .A2(n1105), .ZN(n1335) );
NAND2_X1 U1051 ( .A1(n1337), .A2(n1338), .ZN(n1333) );
OR2_X1 U1052 ( .A1(n1339), .A2(n1171), .ZN(n1338) );
NAND2_X1 U1053 ( .A1(n1340), .A2(n1171), .ZN(n1337) );
XOR2_X1 U1054 ( .A(n1323), .B(KEYINPUT33), .Z(n1171) );
XNOR2_X1 U1055 ( .A(n1341), .B(n1342), .ZN(n1323) );
XNOR2_X1 U1056 ( .A(KEYINPUT58), .B(n1343), .ZN(n1342) );
INV_X1 U1057 ( .A(G107), .ZN(n1343) );
XNOR2_X1 U1058 ( .A(G101), .B(G104), .ZN(n1341) );
XNOR2_X1 U1059 ( .A(KEYINPUT35), .B(n1339), .ZN(n1340) );
INV_X1 U1060 ( .A(n1174), .ZN(n1339) );
XOR2_X1 U1061 ( .A(n1300), .B(n1117), .Z(n1174) );
XNOR2_X1 U1062 ( .A(n1329), .B(n1344), .ZN(n1117) );
NOR2_X1 U1063 ( .A1(KEYINPUT5), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1064 ( .A(n1346), .B(n1238), .Z(n1300) );
INV_X1 U1065 ( .A(G131), .ZN(n1238) );
NAND2_X1 U1066 ( .A1(KEYINPUT19), .A2(n1114), .ZN(n1346) );
XNOR2_X1 U1067 ( .A(G134), .B(n1115), .ZN(n1114) );
INV_X1 U1068 ( .A(G137), .ZN(n1115) );
NAND2_X1 U1069 ( .A1(n1267), .A2(n1347), .ZN(n1048) );
XNOR2_X1 U1070 ( .A(KEYINPUT21), .B(n1266), .ZN(n1347) );
INV_X1 U1071 ( .A(n1099), .ZN(n1266) );
XNOR2_X1 U1072 ( .A(n1348), .B(G475), .ZN(n1099) );
NAND2_X1 U1073 ( .A1(n1179), .A2(n1147), .ZN(n1348) );
NAND2_X1 U1074 ( .A1(n1349), .A2(n1350), .ZN(n1147) );
NAND2_X1 U1075 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
XOR2_X1 U1076 ( .A(KEYINPUT18), .B(n1353), .Z(n1349) );
NOR2_X1 U1077 ( .A1(n1351), .A2(n1352), .ZN(n1353) );
XNOR2_X1 U1078 ( .A(n1151), .B(n1325), .ZN(n1352) );
XOR2_X1 U1079 ( .A(G113), .B(G122), .Z(n1325) );
INV_X1 U1080 ( .A(G104), .ZN(n1151) );
XOR2_X1 U1081 ( .A(n1354), .B(n1355), .Z(n1351) );
XNOR2_X1 U1082 ( .A(n1356), .B(n1357), .ZN(n1355) );
AND2_X1 U1083 ( .A1(G214), .A2(n1294), .ZN(n1357) );
NOR2_X1 U1084 ( .A1(G953), .A2(G237), .ZN(n1294) );
NAND2_X1 U1085 ( .A1(KEYINPUT26), .A2(G131), .ZN(n1356) );
XOR2_X1 U1086 ( .A(n1358), .B(n1359), .Z(n1354) );
XNOR2_X1 U1087 ( .A(n1345), .B(G143), .ZN(n1359) );
INV_X1 U1088 ( .A(G146), .ZN(n1345) );
NAND2_X1 U1089 ( .A1(n1360), .A2(n1285), .ZN(n1358) );
XNOR2_X1 U1090 ( .A(G140), .B(n1217), .ZN(n1285) );
INV_X1 U1091 ( .A(G125), .ZN(n1217) );
XOR2_X1 U1092 ( .A(KEYINPUT55), .B(KEYINPUT45), .Z(n1360) );
INV_X1 U1093 ( .A(G902), .ZN(n1179) );
XNOR2_X1 U1094 ( .A(n1092), .B(G478), .ZN(n1267) );
NOR2_X1 U1095 ( .A1(n1143), .A2(G902), .ZN(n1092) );
XNOR2_X1 U1096 ( .A(n1361), .B(n1362), .ZN(n1143) );
XOR2_X1 U1097 ( .A(n1363), .B(n1364), .Z(n1362) );
NAND3_X1 U1098 ( .A1(G217), .A2(n1287), .A3(KEYINPUT51), .ZN(n1364) );
AND2_X1 U1099 ( .A1(G234), .A2(n1105), .ZN(n1287) );
INV_X1 U1100 ( .A(G953), .ZN(n1105) );
NAND2_X1 U1101 ( .A1(n1365), .A2(n1366), .ZN(n1363) );
NAND2_X1 U1102 ( .A1(n1329), .A2(n1236), .ZN(n1366) );
XOR2_X1 U1103 ( .A(KEYINPUT43), .B(n1367), .Z(n1365) );
NOR2_X1 U1104 ( .A1(n1329), .A2(n1236), .ZN(n1367) );
INV_X1 U1105 ( .A(G134), .ZN(n1236) );
XOR2_X1 U1106 ( .A(G128), .B(n1223), .Z(n1329) );
INV_X1 U1107 ( .A(G143), .ZN(n1223) );
XOR2_X1 U1108 ( .A(n1368), .B(n1369), .Z(n1361) );
NOR2_X1 U1109 ( .A1(KEYINPUT31), .A2(n1370), .ZN(n1369) );
XNOR2_X1 U1110 ( .A(G122), .B(KEYINPUT56), .ZN(n1370) );
XNOR2_X1 U1111 ( .A(G107), .B(G116), .ZN(n1368) );
INV_X1 U1112 ( .A(G110), .ZN(n1272) );
endmodule


