//Key = 0001111000111100011110001100111000101011111111110110100100100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399;

XOR2_X1 U768 ( .A(G107), .B(n1068), .Z(G9) );
NOR2_X1 U769 ( .A1(n1069), .A2(n1070), .ZN(G75) );
XOR2_X1 U770 ( .A(n1071), .B(KEYINPUT3), .Z(n1070) );
NAND3_X1 U771 ( .A1(n1072), .A2(G952), .A3(n1073), .ZN(n1071) );
NOR3_X1 U772 ( .A1(n1074), .A2(G953), .A3(n1075), .ZN(n1073) );
NOR2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR3_X1 U775 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NAND3_X1 U776 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1080) );
OR2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND3_X1 U778 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1084) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND3_X1 U780 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1096), .A2(n1097), .ZN(n1083) );
NAND2_X1 U782 ( .A1(n1091), .A2(n1094), .ZN(n1097) );
INV_X1 U783 ( .A(KEYINPUT48), .ZN(n1094) );
NOR4_X1 U784 ( .A1(n1096), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1078) );
NOR2_X1 U785 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NOR2_X1 U786 ( .A1(n1082), .A2(n1103), .ZN(n1102) );
NOR3_X1 U787 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1101) );
NOR3_X1 U788 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
NOR2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U790 ( .A1(n1112), .A2(n1113), .ZN(n1105) );
NOR3_X1 U791 ( .A1(n1114), .A2(G952), .A3(n1075), .ZN(n1069) );
AND4_X1 U792 ( .A1(n1115), .A2(n1093), .A3(n1116), .A4(n1117), .ZN(n1075) );
NOR4_X1 U793 ( .A1(n1118), .A2(n1082), .A3(n1119), .A4(n1120), .ZN(n1117) );
NOR3_X1 U794 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
INV_X1 U795 ( .A(KEYINPUT49), .ZN(n1121) );
NOR2_X1 U796 ( .A1(KEYINPUT49), .A2(G478), .ZN(n1119) );
NAND3_X1 U797 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1118) );
XNOR2_X1 U798 ( .A(G475), .B(n1127), .ZN(n1126) );
NAND2_X1 U799 ( .A1(KEYINPUT38), .A2(n1128), .ZN(n1127) );
NAND2_X1 U800 ( .A1(n1129), .A2(n1130), .ZN(n1125) );
XOR2_X1 U801 ( .A(KEYINPUT33), .B(G472), .Z(n1129) );
XOR2_X1 U802 ( .A(n1131), .B(n1132), .Z(n1124) );
NAND2_X1 U803 ( .A1(KEYINPUT39), .A2(n1133), .ZN(n1132) );
INV_X1 U804 ( .A(G469), .ZN(n1133) );
NOR3_X1 U805 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1116) );
INV_X1 U806 ( .A(n1137), .ZN(n1134) );
NAND2_X1 U807 ( .A1(n1138), .A2(n1139), .ZN(n1115) );
XOR2_X1 U808 ( .A(n1140), .B(KEYINPUT44), .Z(n1114) );
XOR2_X1 U809 ( .A(n1141), .B(n1142), .Z(G72) );
NOR2_X1 U810 ( .A1(n1143), .A2(n1140), .ZN(n1142) );
NOR2_X1 U811 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NAND2_X1 U812 ( .A1(n1146), .A2(n1147), .ZN(n1141) );
NAND2_X1 U813 ( .A1(n1148), .A2(n1140), .ZN(n1147) );
XOR2_X1 U814 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND3_X1 U815 ( .A1(G900), .A2(n1150), .A3(G953), .ZN(n1146) );
XNOR2_X1 U816 ( .A(n1151), .B(n1152), .ZN(n1150) );
XOR2_X1 U817 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U818 ( .A(n1155), .B(n1156), .Z(n1151) );
NAND2_X1 U819 ( .A1(KEYINPUT6), .A2(n1157), .ZN(n1155) );
NAND2_X1 U820 ( .A1(n1158), .A2(n1159), .ZN(G69) );
NAND2_X1 U821 ( .A1(n1160), .A2(n1140), .ZN(n1159) );
XNOR2_X1 U822 ( .A(n1161), .B(n1162), .ZN(n1160) );
NAND2_X1 U823 ( .A1(n1163), .A2(G953), .ZN(n1158) );
NAND2_X1 U824 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U825 ( .A1(n1162), .A2(n1166), .ZN(n1165) );
INV_X1 U826 ( .A(G224), .ZN(n1166) );
NAND2_X1 U827 ( .A1(G224), .A2(n1167), .ZN(n1164) );
NAND2_X1 U828 ( .A1(G898), .A2(n1162), .ZN(n1167) );
NAND2_X1 U829 ( .A1(n1168), .A2(n1169), .ZN(n1162) );
NAND2_X1 U830 ( .A1(G953), .A2(n1170), .ZN(n1169) );
XNOR2_X1 U831 ( .A(n1171), .B(n1172), .ZN(n1168) );
NOR2_X1 U832 ( .A1(KEYINPUT59), .A2(n1173), .ZN(n1172) );
XOR2_X1 U833 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U834 ( .A1(KEYINPUT0), .A2(n1176), .ZN(n1174) );
NOR2_X1 U835 ( .A1(n1177), .A2(n1178), .ZN(G66) );
NOR2_X1 U836 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U837 ( .A(n1181), .B(KEYINPUT58), .Z(n1180) );
NAND2_X1 U838 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U839 ( .A1(n1136), .A2(n1184), .ZN(n1183) );
NOR3_X1 U840 ( .A1(n1185), .A2(n1182), .A3(n1139), .ZN(n1179) );
NOR2_X1 U841 ( .A1(n1177), .A2(n1186), .ZN(G63) );
XOR2_X1 U842 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U843 ( .A(n1189), .B(KEYINPUT46), .Z(n1188) );
NAND2_X1 U844 ( .A1(n1190), .A2(G478), .ZN(n1189) );
NOR2_X1 U845 ( .A1(n1177), .A2(n1191), .ZN(G60) );
XOR2_X1 U846 ( .A(n1192), .B(n1193), .Z(n1191) );
NAND2_X1 U847 ( .A1(n1190), .A2(G475), .ZN(n1192) );
XNOR2_X1 U848 ( .A(G104), .B(n1194), .ZN(G6) );
NOR2_X1 U849 ( .A1(n1177), .A2(n1195), .ZN(G57) );
XOR2_X1 U850 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U851 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
NAND2_X1 U852 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U853 ( .A1(n1190), .A2(G472), .ZN(n1201) );
XOR2_X1 U854 ( .A(n1202), .B(KEYINPUT63), .Z(n1198) );
NAND3_X1 U855 ( .A1(n1190), .A2(G472), .A3(n1203), .ZN(n1202) );
INV_X1 U856 ( .A(n1200), .ZN(n1203) );
XOR2_X1 U857 ( .A(n1204), .B(n1205), .Z(n1200) );
NOR2_X1 U858 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U859 ( .A1(KEYINPUT55), .A2(n1208), .ZN(n1207) );
AND2_X1 U860 ( .A1(KEYINPUT43), .A2(n1208), .ZN(n1206) );
NAND2_X1 U861 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U862 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U863 ( .A(n1213), .B(KEYINPUT28), .Z(n1211) );
NAND2_X1 U864 ( .A1(n1214), .A2(n1215), .ZN(n1209) );
XOR2_X1 U865 ( .A(KEYINPUT10), .B(n1216), .Z(n1214) );
NOR2_X1 U866 ( .A1(n1177), .A2(n1217), .ZN(G54) );
XOR2_X1 U867 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U868 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U869 ( .A(n1222), .B(n1213), .Z(n1221) );
NAND2_X1 U870 ( .A1(KEYINPUT12), .A2(n1223), .ZN(n1222) );
XOR2_X1 U871 ( .A(n1224), .B(n1225), .Z(n1218) );
XOR2_X1 U872 ( .A(n1226), .B(n1227), .Z(n1225) );
NAND2_X1 U873 ( .A1(n1228), .A2(n1229), .ZN(n1226) );
NAND2_X1 U874 ( .A1(G110), .A2(n1157), .ZN(n1229) );
XOR2_X1 U875 ( .A(KEYINPUT62), .B(n1230), .Z(n1228) );
NOR2_X1 U876 ( .A1(G110), .A2(n1157), .ZN(n1230) );
NAND2_X1 U877 ( .A1(n1190), .A2(G469), .ZN(n1224) );
INV_X1 U878 ( .A(n1185), .ZN(n1190) );
NOR2_X1 U879 ( .A1(n1177), .A2(n1231), .ZN(G51) );
XOR2_X1 U880 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U881 ( .A(n1234), .B(n1235), .Z(n1233) );
NOR3_X1 U882 ( .A1(n1185), .A2(KEYINPUT27), .A3(n1236), .ZN(n1235) );
NAND2_X1 U883 ( .A1(G902), .A2(n1184), .ZN(n1185) );
INV_X1 U884 ( .A(n1072), .ZN(n1184) );
NOR2_X1 U885 ( .A1(n1149), .A2(n1161), .ZN(n1072) );
NAND4_X1 U886 ( .A1(n1194), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1161) );
NOR4_X1 U887 ( .A1(n1068), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1239) );
NOR3_X1 U888 ( .A1(n1243), .A2(n1081), .A3(n1088), .ZN(n1068) );
NOR2_X1 U889 ( .A1(n1244), .A2(n1245), .ZN(n1238) );
NOR2_X1 U890 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U891 ( .A(n1248), .B(KEYINPUT7), .Z(n1246) );
NOR3_X1 U892 ( .A1(n1099), .A2(n1249), .A3(n1243), .ZN(n1244) );
XOR2_X1 U893 ( .A(n1103), .B(KEYINPUT31), .Z(n1249) );
OR3_X1 U894 ( .A1(n1243), .A2(n1081), .A3(n1089), .ZN(n1194) );
NAND4_X1 U895 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1149) );
AND4_X1 U896 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1253) );
NOR3_X1 U897 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1252) );
NOR3_X1 U898 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1260) );
AND2_X1 U899 ( .A1(n1261), .A2(n1264), .ZN(n1259) );
INV_X1 U900 ( .A(KEYINPUT26), .ZN(n1261) );
NOR3_X1 U901 ( .A1(n1265), .A2(n1247), .A3(n1088), .ZN(n1258) );
NOR2_X1 U902 ( .A1(n1266), .A2(n1267), .ZN(n1234) );
XNOR2_X1 U903 ( .A(KEYINPUT53), .B(KEYINPUT30), .ZN(n1267) );
NOR2_X1 U904 ( .A1(n1140), .A2(G952), .ZN(n1177) );
XOR2_X1 U905 ( .A(n1268), .B(n1251), .Z(G48) );
OR3_X1 U906 ( .A1(n1265), .A2(n1247), .A3(n1089), .ZN(n1251) );
XOR2_X1 U907 ( .A(n1257), .B(n1269), .Z(G45) );
NAND2_X1 U908 ( .A1(KEYINPUT20), .A2(G143), .ZN(n1269) );
NAND4_X1 U909 ( .A1(n1270), .A2(n1271), .A3(n1108), .A4(n1272), .ZN(n1257) );
NOR2_X1 U910 ( .A1(n1103), .A2(n1273), .ZN(n1272) );
XOR2_X1 U911 ( .A(n1256), .B(n1274), .Z(G42) );
XOR2_X1 U912 ( .A(KEYINPUT45), .B(G140), .Z(n1274) );
NAND3_X1 U913 ( .A1(n1262), .A2(n1275), .A3(n1276), .ZN(n1256) );
NOR3_X1 U914 ( .A1(n1082), .A2(n1112), .A3(n1104), .ZN(n1276) );
XNOR2_X1 U915 ( .A(G137), .B(n1255), .ZN(G39) );
OR3_X1 U916 ( .A1(n1265), .A2(n1082), .A3(n1099), .ZN(n1255) );
XNOR2_X1 U917 ( .A(n1254), .B(n1277), .ZN(G36) );
NOR2_X1 U918 ( .A1(KEYINPUT21), .A2(n1278), .ZN(n1277) );
INV_X1 U919 ( .A(G134), .ZN(n1278) );
OR4_X1 U920 ( .A1(n1273), .A2(n1103), .A3(n1082), .A4(n1088), .ZN(n1254) );
NAND2_X1 U921 ( .A1(n1279), .A2(n1280), .ZN(G33) );
NAND2_X1 U922 ( .A1(G131), .A2(n1250), .ZN(n1280) );
XOR2_X1 U923 ( .A(KEYINPUT42), .B(n1281), .Z(n1279) );
NOR2_X1 U924 ( .A1(G131), .A2(n1250), .ZN(n1281) );
NAND4_X1 U925 ( .A1(n1262), .A2(n1275), .A3(n1282), .A4(n1113), .ZN(n1250) );
INV_X1 U926 ( .A(n1082), .ZN(n1113) );
NAND2_X1 U927 ( .A1(n1283), .A2(n1111), .ZN(n1082) );
INV_X1 U928 ( .A(n1103), .ZN(n1282) );
XNOR2_X1 U929 ( .A(G128), .B(n1284), .ZN(G30) );
NAND2_X1 U930 ( .A1(n1108), .A2(n1285), .ZN(n1284) );
XOR2_X1 U931 ( .A(KEYINPUT22), .B(n1286), .Z(n1285) );
NOR2_X1 U932 ( .A1(n1088), .A2(n1265), .ZN(n1286) );
NAND3_X1 U933 ( .A1(n1107), .A2(n1104), .A3(n1275), .ZN(n1265) );
INV_X1 U934 ( .A(n1273), .ZN(n1275) );
NAND2_X1 U935 ( .A1(n1287), .A2(n1288), .ZN(n1273) );
XOR2_X1 U936 ( .A(G101), .B(n1289), .Z(G3) );
NOR3_X1 U937 ( .A1(n1099), .A2(n1243), .A3(n1103), .ZN(n1289) );
NAND3_X1 U938 ( .A1(n1287), .A2(n1290), .A3(n1108), .ZN(n1243) );
INV_X1 U939 ( .A(n1247), .ZN(n1108) );
INV_X1 U940 ( .A(n1095), .ZN(n1287) );
XOR2_X1 U941 ( .A(G125), .B(n1264), .Z(G27) );
NOR2_X1 U942 ( .A1(n1263), .A2(n1089), .ZN(n1264) );
NAND4_X1 U943 ( .A1(n1291), .A2(n1292), .A3(n1288), .A4(n1107), .ZN(n1263) );
NAND2_X1 U944 ( .A1(n1077), .A2(n1293), .ZN(n1288) );
NAND2_X1 U945 ( .A1(n1294), .A2(n1145), .ZN(n1293) );
INV_X1 U946 ( .A(G900), .ZN(n1145) );
NAND2_X1 U947 ( .A1(n1295), .A2(n1296), .ZN(G24) );
NAND2_X1 U948 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U949 ( .A(n1237), .B(KEYINPUT25), .Z(n1297) );
NAND2_X1 U950 ( .A1(G122), .A2(n1299), .ZN(n1295) );
XOR2_X1 U951 ( .A(n1237), .B(KEYINPUT1), .Z(n1299) );
OR4_X1 U952 ( .A1(n1300), .A2(n1081), .A3(n1301), .A4(n1302), .ZN(n1237) );
INV_X1 U953 ( .A(n1271), .ZN(n1302) );
NAND2_X1 U954 ( .A1(n1292), .A2(n1112), .ZN(n1081) );
XOR2_X1 U955 ( .A(G119), .B(n1242), .Z(G21) );
NOR4_X1 U956 ( .A1(n1300), .A2(n1099), .A3(n1112), .A4(n1292), .ZN(n1242) );
XOR2_X1 U957 ( .A(G116), .B(n1241), .Z(G18) );
NOR3_X1 U958 ( .A1(n1103), .A2(n1088), .A3(n1300), .ZN(n1241) );
NAND2_X1 U959 ( .A1(n1301), .A2(n1303), .ZN(n1088) );
XNOR2_X1 U960 ( .A(KEYINPUT36), .B(n1271), .ZN(n1303) );
XOR2_X1 U961 ( .A(G113), .B(n1240), .Z(G15) );
NOR3_X1 U962 ( .A1(n1089), .A2(n1103), .A3(n1300), .ZN(n1240) );
NAND2_X1 U963 ( .A1(n1291), .A2(n1290), .ZN(n1300) );
NOR3_X1 U964 ( .A1(n1247), .A2(n1096), .A3(n1100), .ZN(n1291) );
INV_X1 U965 ( .A(n1093), .ZN(n1096) );
NAND2_X1 U966 ( .A1(n1112), .A2(n1104), .ZN(n1103) );
INV_X1 U967 ( .A(n1292), .ZN(n1104) );
INV_X1 U968 ( .A(n1262), .ZN(n1089) );
NOR2_X1 U969 ( .A1(n1271), .A2(n1301), .ZN(n1262) );
XOR2_X1 U970 ( .A(G110), .B(n1304), .Z(G12) );
NOR2_X1 U971 ( .A1(n1247), .A2(n1248), .ZN(n1304) );
NAND4_X1 U972 ( .A1(n1087), .A2(n1292), .A3(n1290), .A4(n1107), .ZN(n1248) );
INV_X1 U973 ( .A(n1112), .ZN(n1107) );
NOR2_X1 U974 ( .A1(n1305), .A2(n1136), .ZN(n1112) );
NOR2_X1 U975 ( .A1(n1139), .A2(n1138), .ZN(n1136) );
AND2_X1 U976 ( .A1(n1306), .A2(n1139), .ZN(n1305) );
NAND2_X1 U977 ( .A1(G217), .A2(n1307), .ZN(n1139) );
XNOR2_X1 U978 ( .A(n1138), .B(KEYINPUT50), .ZN(n1306) );
AND2_X1 U979 ( .A1(n1182), .A2(n1308), .ZN(n1138) );
XOR2_X1 U980 ( .A(n1309), .B(n1310), .Z(n1182) );
XOR2_X1 U981 ( .A(n1311), .B(n1312), .Z(n1310) );
XOR2_X1 U982 ( .A(G128), .B(n1313), .Z(n1312) );
NOR2_X1 U983 ( .A1(KEYINPUT15), .A2(n1314), .ZN(n1313) );
XOR2_X1 U984 ( .A(G140), .B(G137), .Z(n1311) );
XOR2_X1 U985 ( .A(n1315), .B(n1316), .Z(n1309) );
XNOR2_X1 U986 ( .A(n1317), .B(n1318), .ZN(n1316) );
NOR2_X1 U987 ( .A1(G146), .A2(KEYINPUT51), .ZN(n1318) );
NAND2_X1 U988 ( .A1(KEYINPUT19), .A2(n1319), .ZN(n1317) );
INV_X1 U989 ( .A(G119), .ZN(n1319) );
XOR2_X1 U990 ( .A(n1320), .B(n1156), .Z(n1315) );
NAND2_X1 U991 ( .A1(G221), .A2(n1321), .ZN(n1320) );
NAND2_X1 U992 ( .A1(n1077), .A2(n1322), .ZN(n1290) );
NAND2_X1 U993 ( .A1(n1294), .A2(n1170), .ZN(n1322) );
INV_X1 U994 ( .A(G898), .ZN(n1170) );
AND3_X1 U995 ( .A1(n1323), .A2(n1324), .A3(G953), .ZN(n1294) );
XOR2_X1 U996 ( .A(KEYINPUT60), .B(G902), .Z(n1323) );
NAND3_X1 U997 ( .A1(n1324), .A2(n1140), .A3(G952), .ZN(n1077) );
NAND2_X1 U998 ( .A1(G234), .A2(G237), .ZN(n1324) );
NOR2_X1 U999 ( .A1(n1325), .A2(n1135), .ZN(n1292) );
NOR2_X1 U1000 ( .A1(n1130), .A2(G472), .ZN(n1135) );
AND2_X1 U1001 ( .A1(G472), .A2(n1130), .ZN(n1325) );
NAND2_X1 U1002 ( .A1(n1326), .A2(n1308), .ZN(n1130) );
XNOR2_X1 U1003 ( .A(n1327), .B(n1197), .ZN(n1326) );
XNOR2_X1 U1004 ( .A(n1328), .B(n1329), .ZN(n1197) );
AND2_X1 U1005 ( .A1(n1330), .A2(G210), .ZN(n1329) );
NAND2_X1 U1006 ( .A1(n1331), .A2(n1332), .ZN(n1327) );
OR2_X1 U1007 ( .A1(n1153), .A2(n1204), .ZN(n1332) );
XOR2_X1 U1008 ( .A(n1333), .B(KEYINPUT2), .Z(n1331) );
NAND2_X1 U1009 ( .A1(n1204), .A2(n1153), .ZN(n1333) );
XOR2_X1 U1010 ( .A(n1213), .B(n1212), .Z(n1153) );
XOR2_X1 U1011 ( .A(n1334), .B(n1335), .Z(n1204) );
XOR2_X1 U1012 ( .A(KEYINPUT14), .B(G113), .Z(n1335) );
NAND2_X1 U1013 ( .A1(n1336), .A2(n1337), .ZN(n1334) );
NAND2_X1 U1014 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
XOR2_X1 U1015 ( .A(KEYINPUT40), .B(n1340), .Z(n1336) );
NOR2_X1 U1016 ( .A1(n1338), .A2(n1339), .ZN(n1340) );
XOR2_X1 U1017 ( .A(G119), .B(KEYINPUT9), .Z(n1339) );
XNOR2_X1 U1018 ( .A(KEYINPUT54), .B(G116), .ZN(n1338) );
NOR2_X1 U1019 ( .A1(n1099), .A2(n1095), .ZN(n1087) );
NAND2_X1 U1020 ( .A1(n1100), .A2(n1093), .ZN(n1095) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1307), .ZN(n1093) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1308), .ZN(n1307) );
INV_X1 U1023 ( .A(n1086), .ZN(n1100) );
XOR2_X1 U1024 ( .A(n1131), .B(G469), .Z(n1086) );
NAND2_X1 U1025 ( .A1(n1341), .A2(n1308), .ZN(n1131) );
XOR2_X1 U1026 ( .A(n1342), .B(n1343), .Z(n1341) );
XOR2_X1 U1027 ( .A(n1344), .B(n1345), .Z(n1343) );
NAND2_X1 U1028 ( .A1(KEYINPUT17), .A2(n1216), .ZN(n1345) );
INV_X1 U1029 ( .A(n1213), .ZN(n1216) );
XNOR2_X1 U1030 ( .A(G131), .B(n1346), .ZN(n1213) );
XOR2_X1 U1031 ( .A(G137), .B(G134), .Z(n1346) );
NAND2_X1 U1032 ( .A1(n1347), .A2(n1348), .ZN(n1344) );
NAND2_X1 U1033 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
XOR2_X1 U1034 ( .A(KEYINPUT41), .B(n1351), .Z(n1347) );
NOR2_X1 U1035 ( .A1(n1350), .A2(n1349), .ZN(n1351) );
XOR2_X1 U1036 ( .A(KEYINPUT37), .B(n1227), .Z(n1349) );
NOR2_X1 U1037 ( .A1(n1144), .A2(G953), .ZN(n1227) );
INV_X1 U1038 ( .A(G227), .ZN(n1144) );
XOR2_X1 U1039 ( .A(G110), .B(n1352), .Z(n1350) );
NOR2_X1 U1040 ( .A1(G140), .A2(KEYINPUT23), .ZN(n1352) );
XNOR2_X1 U1041 ( .A(n1223), .B(n1220), .ZN(n1342) );
XNOR2_X1 U1042 ( .A(n1353), .B(n1354), .ZN(n1220) );
XOR2_X1 U1043 ( .A(KEYINPUT18), .B(G107), .Z(n1354) );
XOR2_X1 U1044 ( .A(n1328), .B(G104), .Z(n1353) );
INV_X1 U1045 ( .A(G101), .ZN(n1328) );
XOR2_X1 U1046 ( .A(n1154), .B(n1215), .Z(n1223) );
INV_X1 U1047 ( .A(n1212), .ZN(n1215) );
XOR2_X1 U1048 ( .A(KEYINPUT57), .B(KEYINPUT47), .Z(n1154) );
INV_X1 U1049 ( .A(n1091), .ZN(n1099) );
NOR2_X1 U1050 ( .A1(n1270), .A2(n1271), .ZN(n1091) );
NAND3_X1 U1051 ( .A1(n1355), .A2(n1356), .A3(n1137), .ZN(n1271) );
NAND2_X1 U1052 ( .A1(n1122), .A2(n1123), .ZN(n1137) );
NAND2_X1 U1053 ( .A1(n1123), .A2(n1357), .ZN(n1356) );
OR3_X1 U1054 ( .A1(n1123), .A2(n1122), .A3(n1357), .ZN(n1355) );
INV_X1 U1055 ( .A(KEYINPUT11), .ZN(n1357) );
NOR2_X1 U1056 ( .A1(n1187), .A2(G902), .ZN(n1122) );
XOR2_X1 U1057 ( .A(n1358), .B(n1359), .Z(n1187) );
XOR2_X1 U1058 ( .A(G116), .B(n1360), .Z(n1359) );
XOR2_X1 U1059 ( .A(G134), .B(G122), .Z(n1360) );
XOR2_X1 U1060 ( .A(n1361), .B(n1362), .Z(n1358) );
XOR2_X1 U1061 ( .A(n1363), .B(G107), .Z(n1361) );
NAND3_X1 U1062 ( .A1(G217), .A2(n1321), .A3(KEYINPUT4), .ZN(n1363) );
AND2_X1 U1063 ( .A1(G234), .A2(n1140), .ZN(n1321) );
INV_X1 U1064 ( .A(G478), .ZN(n1123) );
INV_X1 U1065 ( .A(n1301), .ZN(n1270) );
XOR2_X1 U1066 ( .A(n1128), .B(G475), .Z(n1301) );
NAND2_X1 U1067 ( .A1(n1364), .A2(n1308), .ZN(n1128) );
XOR2_X1 U1068 ( .A(n1193), .B(KEYINPUT16), .Z(n1364) );
XOR2_X1 U1069 ( .A(n1365), .B(n1366), .Z(n1193) );
XOR2_X1 U1070 ( .A(n1367), .B(n1368), .Z(n1366) );
XOR2_X1 U1071 ( .A(n1369), .B(n1370), .Z(n1368) );
NOR3_X1 U1072 ( .A1(KEYINPUT35), .A2(n1371), .A3(n1372), .ZN(n1370) );
NOR2_X1 U1073 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XOR2_X1 U1074 ( .A(n1375), .B(KEYINPUT13), .Z(n1374) );
NOR2_X1 U1075 ( .A1(n1376), .A2(n1375), .ZN(n1371) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1330), .ZN(n1375) );
AND2_X1 U1077 ( .A1(n1377), .A2(n1140), .ZN(n1330) );
XOR2_X1 U1078 ( .A(KEYINPUT61), .B(G237), .Z(n1377) );
NAND2_X1 U1079 ( .A1(n1378), .A2(n1379), .ZN(n1369) );
NAND2_X1 U1080 ( .A1(n1380), .A2(n1157), .ZN(n1379) );
INV_X1 U1081 ( .A(G140), .ZN(n1157) );
XOR2_X1 U1082 ( .A(KEYINPUT5), .B(n1156), .Z(n1380) );
XOR2_X1 U1083 ( .A(n1381), .B(KEYINPUT8), .Z(n1378) );
NAND2_X1 U1084 ( .A1(G140), .A2(n1382), .ZN(n1381) );
XOR2_X1 U1085 ( .A(KEYINPUT56), .B(n1156), .Z(n1382) );
NAND2_X1 U1086 ( .A1(KEYINPUT24), .A2(n1383), .ZN(n1367) );
XOR2_X1 U1087 ( .A(n1384), .B(n1385), .Z(n1365) );
XOR2_X1 U1088 ( .A(G146), .B(G131), .Z(n1385) );
XOR2_X1 U1089 ( .A(G104), .B(n1298), .Z(n1384) );
NAND2_X1 U1090 ( .A1(n1110), .A2(n1111), .ZN(n1247) );
NAND2_X1 U1091 ( .A1(G214), .A2(n1386), .ZN(n1111) );
INV_X1 U1092 ( .A(n1283), .ZN(n1110) );
XNOR2_X1 U1093 ( .A(n1387), .B(n1236), .ZN(n1283) );
NAND2_X1 U1094 ( .A1(G210), .A2(n1386), .ZN(n1236) );
NAND2_X1 U1095 ( .A1(n1388), .A2(n1308), .ZN(n1386) );
INV_X1 U1096 ( .A(G237), .ZN(n1388) );
NAND2_X1 U1097 ( .A1(n1389), .A2(n1308), .ZN(n1387) );
INV_X1 U1098 ( .A(G902), .ZN(n1308) );
XOR2_X1 U1099 ( .A(n1266), .B(n1232), .Z(n1389) );
XOR2_X1 U1100 ( .A(n1390), .B(n1212), .Z(n1232) );
XOR2_X1 U1101 ( .A(n1268), .B(n1362), .Z(n1212) );
XOR2_X1 U1102 ( .A(G128), .B(n1376), .Z(n1362) );
INV_X1 U1103 ( .A(n1373), .ZN(n1376) );
XNOR2_X1 U1104 ( .A(G143), .B(KEYINPUT32), .ZN(n1373) );
INV_X1 U1105 ( .A(G146), .ZN(n1268) );
XOR2_X1 U1106 ( .A(n1391), .B(n1156), .Z(n1390) );
XOR2_X1 U1107 ( .A(G125), .B(KEYINPUT34), .Z(n1156) );
NAND2_X1 U1108 ( .A1(G224), .A2(n1140), .ZN(n1391) );
INV_X1 U1109 ( .A(G953), .ZN(n1140) );
XOR2_X1 U1110 ( .A(n1392), .B(n1175), .Z(n1266) );
XNOR2_X1 U1111 ( .A(n1393), .B(n1394), .ZN(n1175) );
XOR2_X1 U1112 ( .A(G119), .B(G116), .Z(n1394) );
NAND2_X1 U1113 ( .A1(KEYINPUT52), .A2(n1383), .ZN(n1393) );
INV_X1 U1114 ( .A(G113), .ZN(n1383) );
XNOR2_X1 U1115 ( .A(n1176), .B(n1171), .ZN(n1392) );
XOR2_X1 U1116 ( .A(n1298), .B(n1314), .Z(n1171) );
INV_X1 U1117 ( .A(G110), .ZN(n1314) );
INV_X1 U1118 ( .A(G122), .ZN(n1298) );
XNOR2_X1 U1119 ( .A(n1395), .B(G101), .ZN(n1176) );
NAND2_X1 U1120 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
NAND2_X1 U1121 ( .A1(G104), .A2(n1398), .ZN(n1397) );
XOR2_X1 U1122 ( .A(KEYINPUT29), .B(n1399), .Z(n1396) );
NOR2_X1 U1123 ( .A1(G104), .A2(n1398), .ZN(n1399) );
INV_X1 U1124 ( .A(G107), .ZN(n1398) );
endmodule


