//Key = 0110011011011100001001111101000100111111001110010111010010111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
n1478, n1479, n1480, n1481, n1482, n1483, n1484;

XOR2_X1 U804 ( .A(G107), .B(n1118), .Z(G9) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(G75) );
NOR4_X1 U806 ( .A1(G953), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1120) );
XOR2_X1 U807 ( .A(n1124), .B(KEYINPUT62), .Z(n1122) );
NAND2_X1 U808 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND4_X1 U809 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
NAND2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NAND2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
INV_X1 U812 ( .A(KEYINPUT61), .ZN(n1134) );
NAND4_X1 U813 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1129) );
NAND2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NAND2_X1 U815 ( .A1(n1141), .A2(n1142), .ZN(n1136) );
NAND2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U817 ( .A1(KEYINPUT61), .A2(n1133), .ZN(n1135) );
AND3_X1 U818 ( .A1(n1145), .A2(n1146), .A3(n1139), .ZN(n1133) );
NAND4_X1 U819 ( .A1(n1138), .A2(n1141), .A3(n1139), .A4(n1147), .ZN(n1125) );
NAND2_X1 U820 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U821 ( .A1(n1128), .A2(n1150), .ZN(n1149) );
NAND2_X1 U822 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND2_X1 U823 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U824 ( .A1(n1127), .A2(n1155), .ZN(n1148) );
NAND2_X1 U825 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
INV_X1 U826 ( .A(n1132), .ZN(n1138) );
NOR3_X1 U827 ( .A1(n1121), .A2(G953), .A3(G952), .ZN(n1119) );
AND4_X1 U828 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1121) );
NOR4_X1 U829 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1161) );
XOR2_X1 U830 ( .A(KEYINPUT28), .B(n1166), .Z(n1165) );
NOR2_X1 U831 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U832 ( .A(KEYINPUT56), .B(n1169), .Z(n1168) );
XNOR2_X1 U833 ( .A(n1170), .B(n1171), .ZN(n1163) );
XOR2_X1 U834 ( .A(KEYINPUT33), .B(n1172), .Z(n1171) );
NAND3_X1 U835 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1162) );
XNOR2_X1 U836 ( .A(n1176), .B(KEYINPUT3), .ZN(n1175) );
NAND2_X1 U837 ( .A1(KEYINPUT14), .A2(n1177), .ZN(n1174) );
OR2_X1 U838 ( .A1(n1127), .A2(KEYINPUT14), .ZN(n1173) );
NOR3_X1 U839 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1160) );
NOR2_X1 U840 ( .A1(G478), .A2(n1169), .ZN(n1178) );
XNOR2_X1 U841 ( .A(n1181), .B(KEYINPUT21), .ZN(n1169) );
NAND2_X1 U842 ( .A1(n1182), .A2(n1183), .ZN(n1159) );
XNOR2_X1 U843 ( .A(KEYINPUT9), .B(n1184), .ZN(n1158) );
XOR2_X1 U844 ( .A(n1185), .B(n1186), .Z(G72) );
NOR2_X1 U845 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U846 ( .A(n1189), .B(n1190), .Z(n1188) );
XNOR2_X1 U847 ( .A(n1191), .B(n1192), .ZN(n1190) );
XNOR2_X1 U848 ( .A(n1193), .B(n1194), .ZN(n1189) );
NAND3_X1 U849 ( .A1(n1195), .A2(n1196), .A3(KEYINPUT2), .ZN(n1193) );
NAND2_X1 U850 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
INV_X1 U851 ( .A(KEYINPUT51), .ZN(n1198) );
NAND2_X1 U852 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
OR3_X1 U853 ( .A1(G137), .A2(KEYINPUT63), .A3(G134), .ZN(n1200) );
NAND2_X1 U854 ( .A1(n1201), .A2(G134), .ZN(n1199) );
NAND2_X1 U855 ( .A1(n1202), .A2(KEYINPUT51), .ZN(n1195) );
XOR2_X1 U856 ( .A(G134), .B(n1201), .Z(n1202) );
NOR2_X1 U857 ( .A1(n1203), .A2(G137), .ZN(n1201) );
INV_X1 U858 ( .A(KEYINPUT63), .ZN(n1203) );
NOR2_X1 U859 ( .A1(G900), .A2(n1204), .ZN(n1187) );
NAND2_X1 U860 ( .A1(n1205), .A2(n1206), .ZN(n1185) );
NAND2_X1 U861 ( .A1(G953), .A2(n1207), .ZN(n1206) );
NAND2_X1 U862 ( .A1(G900), .A2(G227), .ZN(n1207) );
XOR2_X1 U863 ( .A(n1208), .B(n1209), .Z(G69) );
NOR2_X1 U864 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U865 ( .A(n1212), .B(KEYINPUT25), .Z(n1211) );
NAND3_X1 U866 ( .A1(n1213), .A2(n1204), .A3(n1214), .ZN(n1212) );
NOR3_X1 U867 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1210) );
AND2_X1 U868 ( .A1(n1204), .A2(n1213), .ZN(n1216) );
NAND2_X1 U869 ( .A1(n1217), .A2(n1218), .ZN(n1213) );
XOR2_X1 U870 ( .A(n1219), .B(KEYINPUT41), .Z(n1217) );
NOR2_X1 U871 ( .A1(G898), .A2(n1204), .ZN(n1215) );
NAND3_X1 U872 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1214) );
NAND2_X1 U873 ( .A1(KEYINPUT17), .A2(n1223), .ZN(n1222) );
OR3_X1 U874 ( .A1(n1223), .A2(KEYINPUT17), .A3(n1224), .ZN(n1221) );
NAND2_X1 U875 ( .A1(n1224), .A2(n1225), .ZN(n1220) );
NAND2_X1 U876 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
INV_X1 U877 ( .A(KEYINPUT17), .ZN(n1227) );
XOR2_X1 U878 ( .A(KEYINPUT39), .B(n1223), .Z(n1226) );
NAND2_X1 U879 ( .A1(G953), .A2(n1228), .ZN(n1208) );
NAND2_X1 U880 ( .A1(G898), .A2(G224), .ZN(n1228) );
NOR2_X1 U881 ( .A1(n1229), .A2(n1230), .ZN(G66) );
NOR3_X1 U882 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1230) );
AND3_X1 U883 ( .A1(n1234), .A2(n1182), .A3(n1235), .ZN(n1233) );
NOR2_X1 U884 ( .A1(n1236), .A2(n1234), .ZN(n1232) );
NOR2_X1 U885 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NOR2_X1 U886 ( .A1(n1229), .A2(n1239), .ZN(G63) );
XOR2_X1 U887 ( .A(n1240), .B(n1241), .Z(n1239) );
NOR2_X1 U888 ( .A1(n1242), .A2(KEYINPUT57), .ZN(n1241) );
INV_X1 U889 ( .A(n1243), .ZN(n1242) );
NAND3_X1 U890 ( .A1(G478), .A2(n1244), .A3(G902), .ZN(n1240) );
XNOR2_X1 U891 ( .A(KEYINPUT44), .B(n1123), .ZN(n1244) );
NOR2_X1 U892 ( .A1(n1229), .A2(n1245), .ZN(G60) );
XOR2_X1 U893 ( .A(n1246), .B(n1247), .Z(n1245) );
NAND2_X1 U894 ( .A1(KEYINPUT38), .A2(n1248), .ZN(n1247) );
NAND2_X1 U895 ( .A1(n1235), .A2(G475), .ZN(n1246) );
XNOR2_X1 U896 ( .A(n1249), .B(n1250), .ZN(G6) );
NOR3_X1 U897 ( .A1(n1251), .A2(n1229), .A3(n1252), .ZN(G57) );
NOR4_X1 U898 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1252) );
NOR2_X1 U899 ( .A1(n1257), .A2(n1258), .ZN(n1254) );
NOR2_X1 U900 ( .A1(n1259), .A2(n1260), .ZN(n1253) );
NOR3_X1 U901 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1251) );
NOR2_X1 U902 ( .A1(n1258), .A2(n1260), .ZN(n1263) );
XNOR2_X1 U903 ( .A(n1259), .B(n1264), .ZN(n1258) );
XOR2_X1 U904 ( .A(KEYINPUT40), .B(KEYINPUT29), .Z(n1264) );
NOR2_X1 U905 ( .A1(n1257), .A2(n1259), .ZN(n1262) );
XNOR2_X1 U906 ( .A(n1265), .B(KEYINPUT27), .ZN(n1259) );
INV_X1 U907 ( .A(n1260), .ZN(n1257) );
NAND2_X1 U908 ( .A1(n1235), .A2(G472), .ZN(n1260) );
NOR2_X1 U909 ( .A1(n1255), .A2(n1256), .ZN(n1261) );
INV_X1 U910 ( .A(KEYINPUT53), .ZN(n1256) );
NOR2_X1 U911 ( .A1(n1266), .A2(n1267), .ZN(G54) );
XOR2_X1 U912 ( .A(KEYINPUT46), .B(n1229), .Z(n1267) );
XOR2_X1 U913 ( .A(n1268), .B(n1269), .Z(n1266) );
XOR2_X1 U914 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U915 ( .A(n1272), .B(n1273), .Z(n1271) );
NAND3_X1 U916 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
INV_X1 U917 ( .A(n1277), .ZN(n1276) );
NAND2_X1 U918 ( .A1(n1278), .A2(n1279), .ZN(n1275) );
INV_X1 U919 ( .A(KEYINPUT59), .ZN(n1279) );
XNOR2_X1 U920 ( .A(n1280), .B(n1281), .ZN(n1278) );
NOR2_X1 U921 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U922 ( .A1(KEYINPUT59), .A2(n1284), .ZN(n1274) );
AND2_X1 U923 ( .A1(G469), .A2(n1235), .ZN(n1270) );
XNOR2_X1 U924 ( .A(G110), .B(n1285), .ZN(n1268) );
XNOR2_X1 U925 ( .A(KEYINPUT20), .B(n1286), .ZN(n1285) );
NOR2_X1 U926 ( .A1(n1229), .A2(n1287), .ZN(G51) );
XOR2_X1 U927 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U928 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U929 ( .A(G125), .B(n1292), .ZN(n1291) );
NOR2_X1 U930 ( .A1(n1170), .A2(n1293), .ZN(n1290) );
INV_X1 U931 ( .A(n1235), .ZN(n1293) );
NOR2_X1 U932 ( .A1(n1294), .A2(n1237), .ZN(n1235) );
INV_X1 U933 ( .A(n1123), .ZN(n1237) );
NAND3_X1 U934 ( .A1(n1205), .A2(n1219), .A3(n1218), .ZN(n1123) );
AND4_X1 U935 ( .A1(n1295), .A2(n1296), .A3(n1297), .A4(n1298), .ZN(n1218) );
NOR4_X1 U936 ( .A1(n1299), .A2(n1300), .A3(n1301), .A4(n1302), .ZN(n1298) );
NOR3_X1 U937 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1302) );
INV_X1 U938 ( .A(n1306), .ZN(n1301) );
AND2_X1 U939 ( .A1(KEYINPUT60), .A2(n1250), .ZN(n1300) );
AND2_X1 U940 ( .A1(n1307), .A2(n1308), .ZN(n1250) );
NOR4_X1 U941 ( .A1(KEYINPUT60), .A2(n1309), .A3(n1177), .A4(n1143), .ZN(n1299) );
INV_X1 U942 ( .A(n1310), .ZN(n1177) );
NAND3_X1 U943 ( .A1(n1311), .A2(n1312), .A3(n1128), .ZN(n1309) );
NOR2_X1 U944 ( .A1(n1118), .A2(n1313), .ZN(n1297) );
AND2_X1 U945 ( .A1(n1314), .A2(n1308), .ZN(n1118) );
AND4_X1 U946 ( .A1(n1310), .A2(n1140), .A3(n1128), .A4(n1311), .ZN(n1308) );
AND4_X1 U947 ( .A1(n1315), .A2(n1316), .A3(n1317), .A4(n1318), .ZN(n1205) );
AND4_X1 U948 ( .A1(n1319), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1318) );
NAND3_X1 U949 ( .A1(n1323), .A2(n1324), .A3(n1140), .ZN(n1317) );
NAND2_X1 U950 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
NAND4_X1 U951 ( .A1(n1327), .A2(n1328), .A3(n1329), .A4(n1164), .ZN(n1326) );
NAND3_X1 U952 ( .A1(n1127), .A2(n1330), .A3(n1307), .ZN(n1325) );
NAND3_X1 U953 ( .A1(n1331), .A2(n1332), .A3(n1333), .ZN(n1315) );
XNOR2_X1 U954 ( .A(n1140), .B(KEYINPUT12), .ZN(n1333) );
XOR2_X1 U955 ( .A(n1334), .B(n1335), .Z(n1288) );
NAND2_X1 U956 ( .A1(KEYINPUT8), .A2(n1336), .ZN(n1334) );
NOR2_X1 U957 ( .A1(n1204), .A2(G952), .ZN(n1229) );
XNOR2_X1 U958 ( .A(n1337), .B(n1338), .ZN(G48) );
AND2_X1 U959 ( .A1(n1331), .A2(n1339), .ZN(n1338) );
XNOR2_X1 U960 ( .A(G143), .B(n1340), .ZN(G45) );
NAND4_X1 U961 ( .A1(n1328), .A2(n1140), .A3(n1341), .A4(n1342), .ZN(n1340) );
AND3_X1 U962 ( .A1(n1329), .A2(n1324), .A3(n1164), .ZN(n1342) );
XNOR2_X1 U963 ( .A(n1151), .B(KEYINPUT52), .ZN(n1341) );
XOR2_X1 U964 ( .A(n1321), .B(n1343), .Z(G42) );
XNOR2_X1 U965 ( .A(G140), .B(KEYINPUT7), .ZN(n1343) );
NAND3_X1 U966 ( .A1(n1331), .A2(n1330), .A3(n1141), .ZN(n1321) );
XNOR2_X1 U967 ( .A(G137), .B(n1316), .ZN(G39) );
NAND3_X1 U968 ( .A1(n1327), .A2(n1141), .A3(n1344), .ZN(n1316) );
NOR3_X1 U969 ( .A1(n1303), .A2(n1345), .A3(n1304), .ZN(n1344) );
XNOR2_X1 U970 ( .A(G134), .B(n1320), .ZN(G36) );
NAND3_X1 U971 ( .A1(n1327), .A2(n1141), .A3(n1346), .ZN(n1320) );
NOR3_X1 U972 ( .A1(n1157), .A2(n1345), .A3(n1144), .ZN(n1346) );
INV_X1 U973 ( .A(n1151), .ZN(n1327) );
XNOR2_X1 U974 ( .A(G131), .B(n1319), .ZN(G33) );
NAND3_X1 U975 ( .A1(n1331), .A2(n1328), .A3(n1141), .ZN(n1319) );
AND2_X1 U976 ( .A1(n1146), .A2(n1184), .ZN(n1141) );
NOR3_X1 U977 ( .A1(n1143), .A2(n1345), .A3(n1151), .ZN(n1331) );
XOR2_X1 U978 ( .A(n1310), .B(KEYINPUT24), .Z(n1151) );
XNOR2_X1 U979 ( .A(G128), .B(n1322), .ZN(G30) );
NAND4_X1 U980 ( .A1(n1339), .A2(n1314), .A3(n1310), .A4(n1324), .ZN(n1322) );
XNOR2_X1 U981 ( .A(G101), .B(n1306), .ZN(G3) );
NAND3_X1 U982 ( .A1(n1347), .A2(n1140), .A3(n1328), .ZN(n1306) );
XOR2_X1 U983 ( .A(n1348), .B(n1349), .Z(G27) );
XNOR2_X1 U984 ( .A(KEYINPUT5), .B(n1350), .ZN(n1349) );
NOR2_X1 U985 ( .A1(KEYINPUT48), .A2(n1351), .ZN(n1348) );
NOR4_X1 U986 ( .A1(n1352), .A2(n1156), .A3(n1353), .A4(n1312), .ZN(n1351) );
XNOR2_X1 U987 ( .A(n1345), .B(KEYINPUT36), .ZN(n1353) );
INV_X1 U988 ( .A(n1324), .ZN(n1345) );
NAND2_X1 U989 ( .A1(n1132), .A2(n1354), .ZN(n1324) );
NAND4_X1 U990 ( .A1(G902), .A2(G953), .A3(n1355), .A4(n1356), .ZN(n1354) );
INV_X1 U991 ( .A(G900), .ZN(n1356) );
INV_X1 U992 ( .A(n1330), .ZN(n1156) );
NAND2_X1 U993 ( .A1(n1307), .A2(n1127), .ZN(n1352) );
INV_X1 U994 ( .A(n1143), .ZN(n1307) );
XNOR2_X1 U995 ( .A(G122), .B(n1295), .ZN(G24) );
NAND4_X1 U996 ( .A1(n1357), .A2(n1128), .A3(n1329), .A4(n1164), .ZN(n1295) );
NOR2_X1 U997 ( .A1(n1358), .A2(n1359), .ZN(n1128) );
XNOR2_X1 U998 ( .A(G119), .B(n1360), .ZN(G21) );
NAND4_X1 U999 ( .A1(n1339), .A2(n1139), .A3(n1361), .A4(n1311), .ZN(n1360) );
XOR2_X1 U1000 ( .A(KEYINPUT55), .B(n1127), .Z(n1361) );
NOR2_X1 U1001 ( .A1(n1303), .A2(n1312), .ZN(n1339) );
INV_X1 U1002 ( .A(n1332), .ZN(n1303) );
NOR2_X1 U1003 ( .A1(n1362), .A2(n1363), .ZN(n1332) );
XNOR2_X1 U1004 ( .A(G116), .B(n1296), .ZN(G18) );
NAND3_X1 U1005 ( .A1(n1357), .A2(n1314), .A3(n1328), .ZN(n1296) );
INV_X1 U1006 ( .A(n1144), .ZN(n1314) );
NAND2_X1 U1007 ( .A1(n1364), .A2(n1329), .ZN(n1144) );
XOR2_X1 U1008 ( .A(n1365), .B(KEYINPUT13), .Z(n1329) );
INV_X1 U1009 ( .A(n1305), .ZN(n1357) );
XNOR2_X1 U1010 ( .A(n1366), .B(n1313), .ZN(G15) );
NOR3_X1 U1011 ( .A1(n1305), .A2(n1143), .A3(n1157), .ZN(n1313) );
INV_X1 U1012 ( .A(n1328), .ZN(n1157) );
NOR2_X1 U1013 ( .A1(n1359), .A2(n1363), .ZN(n1328) );
INV_X1 U1014 ( .A(n1362), .ZN(n1359) );
NAND2_X1 U1015 ( .A1(n1367), .A2(n1164), .ZN(n1143) );
XOR2_X1 U1016 ( .A(n1365), .B(KEYINPUT0), .Z(n1367) );
NAND3_X1 U1017 ( .A1(n1140), .A2(n1311), .A3(n1127), .ZN(n1305) );
NOR2_X1 U1018 ( .A1(n1368), .A2(n1153), .ZN(n1127) );
XNOR2_X1 U1019 ( .A(G110), .B(n1369), .ZN(G12) );
NOR2_X1 U1020 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NOR3_X1 U1021 ( .A1(n1372), .A2(n1373), .A3(n1312), .ZN(n1371) );
INV_X1 U1022 ( .A(n1140), .ZN(n1312) );
INV_X1 U1023 ( .A(KEYINPUT30), .ZN(n1372) );
NOR2_X1 U1024 ( .A1(KEYINPUT30), .A2(n1219), .ZN(n1370) );
NAND2_X1 U1025 ( .A1(n1373), .A2(n1140), .ZN(n1219) );
NOR2_X1 U1026 ( .A1(n1146), .A2(n1145), .ZN(n1140) );
INV_X1 U1027 ( .A(n1184), .ZN(n1145) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1374), .ZN(n1184) );
XNOR2_X1 U1029 ( .A(n1375), .B(n1172), .ZN(n1146) );
AND3_X1 U1030 ( .A1(n1376), .A2(n1294), .A3(n1377), .ZN(n1172) );
XOR2_X1 U1031 ( .A(KEYINPUT49), .B(n1378), .Z(n1377) );
NOR2_X1 U1032 ( .A1(n1379), .A2(n1335), .ZN(n1378) );
NAND2_X1 U1033 ( .A1(n1379), .A2(n1335), .ZN(n1376) );
XOR2_X1 U1034 ( .A(n1223), .B(n1224), .Z(n1335) );
XNOR2_X1 U1035 ( .A(n1380), .B(n1381), .ZN(n1224) );
XNOR2_X1 U1036 ( .A(n1382), .B(n1383), .ZN(n1381) );
NAND2_X1 U1037 ( .A1(KEYINPUT22), .A2(n1249), .ZN(n1382) );
XNOR2_X1 U1038 ( .A(n1384), .B(n1366), .ZN(n1380) );
NAND3_X1 U1039 ( .A1(n1385), .A2(n1386), .A3(n1387), .ZN(n1384) );
OR2_X1 U1040 ( .A1(n1388), .A2(KEYINPUT1), .ZN(n1387) );
NAND3_X1 U1041 ( .A1(KEYINPUT1), .A2(n1388), .A3(G116), .ZN(n1386) );
NAND2_X1 U1042 ( .A1(n1389), .A2(n1390), .ZN(n1385) );
INV_X1 U1043 ( .A(G116), .ZN(n1390) );
NAND2_X1 U1044 ( .A1(KEYINPUT1), .A2(n1391), .ZN(n1389) );
XNOR2_X1 U1045 ( .A(KEYINPUT50), .B(n1388), .ZN(n1391) );
AND2_X1 U1046 ( .A1(n1392), .A2(n1393), .ZN(n1223) );
NAND2_X1 U1047 ( .A1(G122), .A2(n1394), .ZN(n1393) );
XOR2_X1 U1048 ( .A(n1395), .B(KEYINPUT10), .Z(n1392) );
OR2_X1 U1049 ( .A1(n1394), .A2(G122), .ZN(n1395) );
AND2_X1 U1050 ( .A1(n1396), .A2(n1397), .ZN(n1379) );
NAND2_X1 U1051 ( .A1(n1398), .A2(n1292), .ZN(n1397) );
XNOR2_X1 U1052 ( .A(n1399), .B(n1336), .ZN(n1398) );
INV_X1 U1053 ( .A(n1400), .ZN(n1336) );
NAND2_X1 U1054 ( .A1(n1401), .A2(n1402), .ZN(n1396) );
XNOR2_X1 U1055 ( .A(n1400), .B(n1399), .ZN(n1402) );
AND2_X1 U1056 ( .A1(KEYINPUT35), .A2(G125), .ZN(n1399) );
INV_X1 U1057 ( .A(n1292), .ZN(n1401) );
NAND2_X1 U1058 ( .A1(G224), .A2(n1403), .ZN(n1292) );
XNOR2_X1 U1059 ( .A(KEYINPUT11), .B(n1204), .ZN(n1403) );
NAND2_X1 U1060 ( .A1(KEYINPUT37), .A2(n1170), .ZN(n1375) );
NAND2_X1 U1061 ( .A1(G210), .A2(n1374), .ZN(n1170) );
NAND2_X1 U1062 ( .A1(n1404), .A2(n1294), .ZN(n1374) );
INV_X1 U1063 ( .A(G237), .ZN(n1404) );
AND2_X1 U1064 ( .A1(n1330), .A2(n1347), .ZN(n1373) );
AND3_X1 U1065 ( .A1(n1310), .A2(n1311), .A3(n1139), .ZN(n1347) );
INV_X1 U1066 ( .A(n1304), .ZN(n1139) );
NAND2_X1 U1067 ( .A1(n1364), .A2(n1365), .ZN(n1304) );
XNOR2_X1 U1068 ( .A(n1181), .B(n1167), .ZN(n1365) );
INV_X1 U1069 ( .A(G478), .ZN(n1167) );
NAND2_X1 U1070 ( .A1(n1294), .A2(n1243), .ZN(n1181) );
NAND2_X1 U1071 ( .A1(n1405), .A2(n1406), .ZN(n1243) );
NAND4_X1 U1072 ( .A1(G234), .A2(G217), .A3(n1407), .A4(n1204), .ZN(n1406) );
NAND2_X1 U1073 ( .A1(n1408), .A2(n1409), .ZN(n1405) );
NAND3_X1 U1074 ( .A1(G217), .A2(n1204), .A3(G234), .ZN(n1409) );
XOR2_X1 U1075 ( .A(KEYINPUT6), .B(n1407), .Z(n1408) );
XNOR2_X1 U1076 ( .A(n1410), .B(n1411), .ZN(n1407) );
XOR2_X1 U1077 ( .A(n1412), .B(n1413), .Z(n1411) );
XOR2_X1 U1078 ( .A(G107), .B(n1414), .Z(n1413) );
NOR2_X1 U1079 ( .A1(G128), .A2(KEYINPUT32), .ZN(n1414) );
XNOR2_X1 U1080 ( .A(G116), .B(n1415), .ZN(n1410) );
XOR2_X1 U1081 ( .A(G134), .B(G122), .Z(n1415) );
INV_X1 U1082 ( .A(n1164), .ZN(n1364) );
XNOR2_X1 U1083 ( .A(n1416), .B(G475), .ZN(n1164) );
OR2_X1 U1084 ( .A1(n1248), .A2(G902), .ZN(n1416) );
XNOR2_X1 U1085 ( .A(n1417), .B(n1418), .ZN(n1248) );
XOR2_X1 U1086 ( .A(n1419), .B(n1420), .Z(n1418) );
XNOR2_X1 U1087 ( .A(G122), .B(n1366), .ZN(n1420) );
XNOR2_X1 U1088 ( .A(KEYINPUT26), .B(n1194), .ZN(n1419) );
INV_X1 U1089 ( .A(G131), .ZN(n1194) );
XOR2_X1 U1090 ( .A(n1421), .B(n1422), .Z(n1417) );
XNOR2_X1 U1091 ( .A(n1249), .B(n1423), .ZN(n1422) );
XOR2_X1 U1092 ( .A(n1424), .B(n1425), .Z(n1421) );
AND2_X1 U1093 ( .A1(n1426), .A2(G214), .ZN(n1425) );
NAND2_X1 U1094 ( .A1(KEYINPUT34), .A2(n1192), .ZN(n1424) );
XNOR2_X1 U1095 ( .A(n1350), .B(G140), .ZN(n1192) );
NAND2_X1 U1096 ( .A1(n1132), .A2(n1427), .ZN(n1311) );
NAND4_X1 U1097 ( .A1(G902), .A2(G953), .A3(n1355), .A4(n1428), .ZN(n1427) );
INV_X1 U1098 ( .A(G898), .ZN(n1428) );
NAND3_X1 U1099 ( .A1(n1355), .A2(n1204), .A3(G952), .ZN(n1132) );
NAND2_X1 U1100 ( .A1(G237), .A2(n1429), .ZN(n1355) );
NOR2_X1 U1101 ( .A1(n1154), .A2(n1153), .ZN(n1310) );
AND2_X1 U1102 ( .A1(G221), .A2(n1430), .ZN(n1153) );
INV_X1 U1103 ( .A(n1368), .ZN(n1154) );
XNOR2_X1 U1104 ( .A(n1431), .B(G469), .ZN(n1368) );
NAND2_X1 U1105 ( .A1(n1432), .A2(n1294), .ZN(n1431) );
XOR2_X1 U1106 ( .A(n1433), .B(n1434), .Z(n1432) );
NOR2_X1 U1107 ( .A1(n1277), .A2(n1284), .ZN(n1434) );
NAND2_X1 U1108 ( .A1(n1435), .A2(n1436), .ZN(n1284) );
NAND3_X1 U1109 ( .A1(n1191), .A2(n1437), .A3(n1438), .ZN(n1436) );
INV_X1 U1110 ( .A(n1280), .ZN(n1438) );
NAND2_X1 U1111 ( .A1(n1439), .A2(n1280), .ZN(n1435) );
XNOR2_X1 U1112 ( .A(n1191), .B(n1282), .ZN(n1439) );
NOR3_X1 U1113 ( .A1(n1191), .A2(n1437), .A3(n1280), .ZN(n1277) );
INV_X1 U1114 ( .A(n1282), .ZN(n1437) );
XOR2_X1 U1115 ( .A(n1440), .B(n1441), .Z(n1282) );
INV_X1 U1116 ( .A(n1383), .ZN(n1441) );
XOR2_X1 U1117 ( .A(G101), .B(G107), .Z(n1383) );
NAND2_X1 U1118 ( .A1(KEYINPUT58), .A2(n1249), .ZN(n1440) );
INV_X1 U1119 ( .A(G104), .ZN(n1249) );
INV_X1 U1120 ( .A(n1283), .ZN(n1191) );
NAND2_X1 U1121 ( .A1(n1442), .A2(n1443), .ZN(n1283) );
NAND2_X1 U1122 ( .A1(G128), .A2(n1444), .ZN(n1443) );
NAND2_X1 U1123 ( .A1(n1445), .A2(n1446), .ZN(n1444) );
NAND2_X1 U1124 ( .A1(n1412), .A2(n1337), .ZN(n1446) );
XNOR2_X1 U1125 ( .A(n1447), .B(n1448), .ZN(n1445) );
NAND2_X1 U1126 ( .A1(n1449), .A2(n1450), .ZN(n1442) );
NAND2_X1 U1127 ( .A1(n1451), .A2(n1452), .ZN(n1449) );
NAND2_X1 U1128 ( .A1(n1448), .A2(n1447), .ZN(n1452) );
INV_X1 U1129 ( .A(KEYINPUT31), .ZN(n1447) );
NAND2_X1 U1130 ( .A1(n1423), .A2(KEYINPUT31), .ZN(n1451) );
XNOR2_X1 U1131 ( .A(n1453), .B(n1272), .ZN(n1433) );
NAND2_X1 U1132 ( .A1(G227), .A2(n1204), .ZN(n1272) );
NAND2_X1 U1133 ( .A1(n1454), .A2(n1455), .ZN(n1453) );
NAND2_X1 U1134 ( .A1(G140), .A2(n1394), .ZN(n1455) );
XOR2_X1 U1135 ( .A(KEYINPUT42), .B(n1456), .Z(n1454) );
NOR2_X1 U1136 ( .A1(G140), .A2(n1394), .ZN(n1456) );
NOR2_X1 U1137 ( .A1(n1358), .A2(n1362), .ZN(n1330) );
NOR2_X1 U1138 ( .A1(n1457), .A2(n1180), .ZN(n1362) );
NOR2_X1 U1139 ( .A1(n1183), .A2(n1182), .ZN(n1180) );
AND2_X1 U1140 ( .A1(n1182), .A2(n1458), .ZN(n1457) );
XNOR2_X1 U1141 ( .A(KEYINPUT47), .B(n1183), .ZN(n1458) );
INV_X1 U1142 ( .A(n1231), .ZN(n1183) );
NOR2_X1 U1143 ( .A1(n1234), .A2(G902), .ZN(n1231) );
XNOR2_X1 U1144 ( .A(n1459), .B(n1460), .ZN(n1234) );
XOR2_X1 U1145 ( .A(n1461), .B(n1462), .Z(n1460) );
NAND3_X1 U1146 ( .A1(G234), .A2(n1204), .A3(G221), .ZN(n1462) );
INV_X1 U1147 ( .A(G953), .ZN(n1204) );
NAND2_X1 U1148 ( .A1(n1463), .A2(n1464), .ZN(n1461) );
XNOR2_X1 U1149 ( .A(n1394), .B(n1465), .ZN(n1464) );
XNOR2_X1 U1150 ( .A(n1450), .B(G119), .ZN(n1465) );
INV_X1 U1151 ( .A(G128), .ZN(n1450) );
INV_X1 U1152 ( .A(G110), .ZN(n1394) );
XNOR2_X1 U1153 ( .A(KEYINPUT4), .B(KEYINPUT15), .ZN(n1463) );
XOR2_X1 U1154 ( .A(n1466), .B(n1467), .Z(n1459) );
XNOR2_X1 U1155 ( .A(n1337), .B(G137), .ZN(n1467) );
NAND2_X1 U1156 ( .A1(n1468), .A2(n1469), .ZN(n1466) );
NAND2_X1 U1157 ( .A1(G140), .A2(n1350), .ZN(n1469) );
INV_X1 U1158 ( .A(G125), .ZN(n1350) );
XOR2_X1 U1159 ( .A(n1470), .B(KEYINPUT16), .Z(n1468) );
NAND2_X1 U1160 ( .A1(G125), .A2(n1286), .ZN(n1470) );
INV_X1 U1161 ( .A(G140), .ZN(n1286) );
INV_X1 U1162 ( .A(n1238), .ZN(n1182) );
NAND2_X1 U1163 ( .A1(G217), .A2(n1430), .ZN(n1238) );
NAND2_X1 U1164 ( .A1(n1429), .A2(n1294), .ZN(n1430) );
INV_X1 U1165 ( .A(G902), .ZN(n1294) );
XNOR2_X1 U1166 ( .A(G234), .B(KEYINPUT43), .ZN(n1429) );
INV_X1 U1167 ( .A(n1363), .ZN(n1358) );
NOR2_X1 U1168 ( .A1(n1176), .A2(n1179), .ZN(n1363) );
NOR3_X1 U1169 ( .A1(G472), .A2(G902), .A3(n1471), .ZN(n1179) );
AND2_X1 U1170 ( .A1(G472), .A2(n1472), .ZN(n1176) );
OR2_X1 U1171 ( .A1(n1471), .A2(G902), .ZN(n1472) );
XOR2_X1 U1172 ( .A(n1255), .B(n1473), .Z(n1471) );
XNOR2_X1 U1173 ( .A(KEYINPUT23), .B(n1474), .ZN(n1473) );
INV_X1 U1174 ( .A(n1265), .ZN(n1474) );
XOR2_X1 U1175 ( .A(n1475), .B(n1476), .Z(n1265) );
INV_X1 U1176 ( .A(G101), .ZN(n1476) );
NAND2_X1 U1177 ( .A1(G210), .A2(n1426), .ZN(n1475) );
NOR2_X1 U1178 ( .A1(G953), .A2(G237), .ZN(n1426) );
XOR2_X1 U1179 ( .A(n1477), .B(n1478), .Z(n1255) );
XOR2_X1 U1180 ( .A(n1479), .B(n1480), .Z(n1478) );
XNOR2_X1 U1181 ( .A(G116), .B(n1481), .ZN(n1480) );
NOR2_X1 U1182 ( .A1(KEYINPUT19), .A2(n1366), .ZN(n1481) );
INV_X1 U1183 ( .A(G113), .ZN(n1366) );
NAND2_X1 U1184 ( .A1(KEYINPUT18), .A2(n1388), .ZN(n1479) );
INV_X1 U1185 ( .A(G119), .ZN(n1388) );
XNOR2_X1 U1186 ( .A(n1400), .B(n1280), .ZN(n1477) );
XOR2_X1 U1187 ( .A(G131), .B(n1482), .Z(n1280) );
XOR2_X1 U1188 ( .A(G137), .B(G134), .Z(n1482) );
XOR2_X1 U1189 ( .A(G128), .B(n1483), .Z(n1400) );
NOR2_X1 U1190 ( .A1(n1423), .A2(KEYINPUT54), .ZN(n1483) );
NOR2_X1 U1191 ( .A1(n1484), .A2(n1448), .ZN(n1423) );
NOR2_X1 U1192 ( .A1(n1337), .A2(n1412), .ZN(n1448) );
AND2_X1 U1193 ( .A1(n1412), .A2(n1337), .ZN(n1484) );
INV_X1 U1194 ( .A(G146), .ZN(n1337) );
XOR2_X1 U1195 ( .A(G143), .B(KEYINPUT45), .Z(n1412) );
endmodule


