//Key = 0110110110010011000010010011000110010100101110001110100010001010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383;

XOR2_X1 U763 ( .A(G107), .B(n1052), .Z(G9) );
NOR2_X1 U764 ( .A1(n1053), .A2(n1054), .ZN(G75) );
NOR3_X1 U765 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
INV_X1 U766 ( .A(n1058), .ZN(n1057) );
NOR2_X1 U767 ( .A1(n1059), .A2(n1060), .ZN(n1056) );
NOR2_X1 U768 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
XOR2_X1 U769 ( .A(KEYINPUT0), .B(n1063), .Z(n1062) );
AND3_X1 U770 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NOR3_X1 U771 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1061) );
INV_X1 U772 ( .A(n1065), .ZN(n1069) );
NOR2_X1 U773 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
AND2_X1 U774 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR3_X1 U775 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1070) );
INV_X1 U776 ( .A(n1077), .ZN(n1076) );
NOR2_X1 U777 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
NOR2_X1 U778 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NAND3_X1 U779 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1055) );
NAND3_X1 U780 ( .A1(n1077), .A2(n1085), .A3(n1064), .ZN(n1084) );
NOR3_X1 U781 ( .A1(n1074), .A2(n1086), .A3(n1067), .ZN(n1064) );
NAND3_X1 U782 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U784 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
XNOR2_X1 U785 ( .A(KEYINPUT41), .B(n1060), .ZN(n1093) );
NAND2_X1 U786 ( .A1(n1065), .A2(n1094), .ZN(n1087) );
NAND2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1099), .B(KEYINPUT51), .Z(n1097) );
AND3_X1 U790 ( .A1(n1082), .A2(n1083), .A3(n1100), .ZN(n1053) );
NAND4_X1 U791 ( .A1(n1101), .A2(n1080), .A3(n1102), .A4(n1103), .ZN(n1082) );
NOR4_X1 U792 ( .A1(n1098), .A2(n1066), .A3(n1104), .A4(n1105), .ZN(n1103) );
XNOR2_X1 U793 ( .A(n1106), .B(n1107), .ZN(n1105) );
NAND2_X1 U794 ( .A1(KEYINPUT37), .A2(n1108), .ZN(n1106) );
XNOR2_X1 U795 ( .A(n1109), .B(n1110), .ZN(n1104) );
XNOR2_X1 U796 ( .A(KEYINPUT50), .B(n1111), .ZN(n1110) );
INV_X1 U797 ( .A(n1112), .ZN(n1098) );
NOR2_X1 U798 ( .A1(n1113), .A2(n1114), .ZN(n1102) );
XNOR2_X1 U799 ( .A(n1115), .B(n1116), .ZN(n1114) );
NAND2_X1 U800 ( .A1(KEYINPUT56), .A2(n1117), .ZN(n1115) );
XNOR2_X1 U801 ( .A(n1118), .B(n1119), .ZN(n1113) );
NOR2_X1 U802 ( .A1(n1120), .A2(KEYINPUT39), .ZN(n1119) );
INV_X1 U803 ( .A(n1121), .ZN(n1080) );
XOR2_X1 U804 ( .A(n1122), .B(n1123), .Z(G72) );
NOR2_X1 U805 ( .A1(n1124), .A2(n1083), .ZN(n1123) );
AND2_X1 U806 ( .A1(G227), .A2(G900), .ZN(n1124) );
NAND2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
NAND3_X1 U808 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
NAND2_X1 U809 ( .A1(KEYINPUT33), .A2(n1130), .ZN(n1128) );
NAND2_X1 U810 ( .A1(G953), .A2(n1131), .ZN(n1130) );
NAND2_X1 U811 ( .A1(G900), .A2(n1132), .ZN(n1131) );
NAND2_X1 U812 ( .A1(n1133), .A2(n1134), .ZN(n1127) );
OR2_X1 U813 ( .A1(n1132), .A2(G953), .ZN(n1133) );
NAND2_X1 U814 ( .A1(n1132), .A2(n1135), .ZN(n1125) );
NAND3_X1 U815 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
OR2_X1 U816 ( .A1(n1129), .A2(n1139), .ZN(n1138) );
NAND2_X1 U817 ( .A1(KEYINPUT33), .A2(n1083), .ZN(n1137) );
NAND3_X1 U818 ( .A1(G900), .A2(n1134), .A3(G953), .ZN(n1136) );
INV_X1 U819 ( .A(KEYINPUT33), .ZN(n1134) );
XNOR2_X1 U820 ( .A(n1140), .B(n1141), .ZN(n1132) );
XNOR2_X1 U821 ( .A(G131), .B(n1142), .ZN(n1141) );
NAND2_X1 U822 ( .A1(KEYINPUT20), .A2(n1143), .ZN(n1142) );
XNOR2_X1 U823 ( .A(n1144), .B(n1145), .ZN(n1140) );
XOR2_X1 U824 ( .A(n1146), .B(n1147), .Z(G69) );
XOR2_X1 U825 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U826 ( .A1(n1150), .A2(n1083), .ZN(n1149) );
AND2_X1 U827 ( .A1(G224), .A2(G898), .ZN(n1150) );
NAND2_X1 U828 ( .A1(n1151), .A2(n1152), .ZN(n1148) );
NAND2_X1 U829 ( .A1(G953), .A2(n1153), .ZN(n1152) );
XOR2_X1 U830 ( .A(n1154), .B(n1155), .Z(n1151) );
NOR2_X1 U831 ( .A1(KEYINPUT55), .A2(n1156), .ZN(n1155) );
XOR2_X1 U832 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U833 ( .A(G101), .B(n1159), .ZN(n1157) );
NOR2_X1 U834 ( .A1(KEYINPUT19), .A2(n1160), .ZN(n1159) );
XNOR2_X1 U835 ( .A(G113), .B(n1161), .ZN(n1160) );
NAND2_X1 U836 ( .A1(n1083), .A2(n1162), .ZN(n1146) );
NOR2_X1 U837 ( .A1(n1163), .A2(n1164), .ZN(G66) );
XNOR2_X1 U838 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U839 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1169), .ZN(G63) );
XOR2_X1 U841 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U842 ( .A1(KEYINPUT23), .A2(n1172), .ZN(n1170) );
NAND2_X1 U843 ( .A1(n1173), .A2(G478), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1163), .A2(n1174), .ZN(G60) );
NOR3_X1 U845 ( .A1(n1109), .A2(n1175), .A3(n1176), .ZN(n1174) );
NOR3_X1 U846 ( .A1(n1177), .A2(n1111), .A3(n1168), .ZN(n1176) );
NOR2_X1 U847 ( .A1(n1178), .A2(n1179), .ZN(n1175) );
NOR2_X1 U848 ( .A1(n1058), .A2(n1111), .ZN(n1178) );
NAND2_X1 U849 ( .A1(n1180), .A2(n1181), .ZN(G6) );
OR2_X1 U850 ( .A1(n1182), .A2(G104), .ZN(n1181) );
XOR2_X1 U851 ( .A(n1183), .B(KEYINPUT13), .Z(n1180) );
NAND2_X1 U852 ( .A1(G104), .A2(n1182), .ZN(n1183) );
NOR2_X1 U853 ( .A1(n1163), .A2(n1184), .ZN(G57) );
XOR2_X1 U854 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U855 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U856 ( .A(n1189), .B(n1190), .Z(n1185) );
NOR2_X1 U857 ( .A1(n1117), .A2(n1168), .ZN(n1189) );
NOR3_X1 U858 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(G54) );
NOR3_X1 U859 ( .A1(n1194), .A2(n1083), .A3(n1100), .ZN(n1193) );
INV_X1 U860 ( .A(G952), .ZN(n1100) );
AND2_X1 U861 ( .A1(n1194), .A2(n1163), .ZN(n1192) );
NOR2_X1 U862 ( .A1(n1083), .A2(G952), .ZN(n1163) );
INV_X1 U863 ( .A(KEYINPUT57), .ZN(n1194) );
XOR2_X1 U864 ( .A(n1195), .B(n1196), .Z(n1191) );
NOR2_X1 U865 ( .A1(n1108), .A2(n1168), .ZN(n1195) );
NOR2_X1 U866 ( .A1(n1197), .A2(n1198), .ZN(G51) );
XOR2_X1 U867 ( .A(n1199), .B(n1200), .Z(n1198) );
XNOR2_X1 U868 ( .A(n1201), .B(n1202), .ZN(n1200) );
NAND3_X1 U869 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1201) );
NAND2_X1 U870 ( .A1(KEYINPUT10), .A2(n1206), .ZN(n1205) );
NAND3_X1 U871 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1204) );
INV_X1 U872 ( .A(KEYINPUT10), .ZN(n1208) );
OR2_X1 U873 ( .A1(n1209), .A2(n1207), .ZN(n1203) );
NOR2_X1 U874 ( .A1(KEYINPUT21), .A2(n1206), .ZN(n1207) );
XOR2_X1 U875 ( .A(n1210), .B(n1211), .Z(n1199) );
NOR2_X1 U876 ( .A1(n1212), .A2(n1168), .ZN(n1211) );
INV_X1 U877 ( .A(n1173), .ZN(n1168) );
NOR2_X1 U878 ( .A1(n1213), .A2(n1058), .ZN(n1173) );
NOR2_X1 U879 ( .A1(n1162), .A2(n1129), .ZN(n1058) );
NAND4_X1 U880 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1129) );
NOR4_X1 U881 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217) );
NOR2_X1 U882 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
INV_X1 U883 ( .A(KEYINPUT26), .ZN(n1223) );
NOR2_X1 U884 ( .A1(n1224), .A2(n1060), .ZN(n1220) );
NOR2_X1 U885 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XNOR2_X1 U886 ( .A(KEYINPUT53), .B(n1227), .ZN(n1226) );
NOR2_X1 U887 ( .A1(n1228), .A2(n1229), .ZN(n1225) );
XNOR2_X1 U888 ( .A(n1092), .B(KEYINPUT12), .ZN(n1228) );
NOR4_X1 U889 ( .A1(n1230), .A2(n1231), .A3(KEYINPUT42), .A4(n1232), .ZN(n1219) );
NOR2_X1 U890 ( .A1(n1233), .A2(n1095), .ZN(n1218) );
NOR3_X1 U891 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
AND3_X1 U892 ( .A1(KEYINPUT42), .A2(n1092), .A3(n1237), .ZN(n1236) );
NOR3_X1 U893 ( .A1(n1229), .A2(KEYINPUT26), .A3(n1238), .ZN(n1235) );
XNOR2_X1 U894 ( .A(n1239), .B(KEYINPUT7), .ZN(n1234) );
NAND4_X1 U895 ( .A1(n1240), .A2(n1182), .A3(n1241), .A4(n1242), .ZN(n1162) );
NOR4_X1 U896 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242) );
NOR2_X1 U897 ( .A1(n1247), .A2(n1052), .ZN(n1241) );
AND3_X1 U898 ( .A1(n1092), .A2(n1073), .A3(n1248), .ZN(n1052) );
NAND3_X1 U899 ( .A1(n1248), .A2(n1073), .A3(n1091), .ZN(n1182) );
NOR2_X1 U900 ( .A1(G952), .A2(n1249), .ZN(n1197) );
XNOR2_X1 U901 ( .A(KEYINPUT31), .B(n1083), .ZN(n1249) );
XNOR2_X1 U902 ( .A(G146), .B(n1250), .ZN(G48) );
NAND2_X1 U903 ( .A1(n1239), .A2(n1230), .ZN(n1250) );
AND2_X1 U904 ( .A1(n1237), .A2(n1091), .ZN(n1239) );
XNOR2_X1 U905 ( .A(G143), .B(n1222), .ZN(G45) );
NAND3_X1 U906 ( .A1(n1238), .A2(n1230), .A3(n1251), .ZN(n1222) );
XNOR2_X1 U907 ( .A(G140), .B(n1252), .ZN(G42) );
NOR2_X1 U908 ( .A1(n1253), .A2(KEYINPUT30), .ZN(n1252) );
NOR2_X1 U909 ( .A1(n1060), .A2(n1227), .ZN(n1253) );
NAND2_X1 U910 ( .A1(n1254), .A2(n1072), .ZN(n1227) );
XNOR2_X1 U911 ( .A(G137), .B(n1216), .ZN(G39) );
NAND3_X1 U912 ( .A1(n1090), .A2(n1065), .A3(n1237), .ZN(n1216) );
NAND2_X1 U913 ( .A1(n1255), .A2(n1256), .ZN(G36) );
OR2_X1 U914 ( .A1(n1143), .A2(n1257), .ZN(n1256) );
XOR2_X1 U915 ( .A(n1258), .B(KEYINPUT24), .Z(n1255) );
NAND2_X1 U916 ( .A1(n1257), .A2(n1143), .ZN(n1258) );
NOR3_X1 U917 ( .A1(n1060), .A2(n1232), .A3(n1229), .ZN(n1257) );
INV_X1 U918 ( .A(n1092), .ZN(n1232) );
XOR2_X1 U919 ( .A(n1214), .B(n1259), .Z(G33) );
XNOR2_X1 U920 ( .A(G131), .B(KEYINPUT36), .ZN(n1259) );
NAND3_X1 U921 ( .A1(n1090), .A2(n1091), .A3(n1251), .ZN(n1214) );
INV_X1 U922 ( .A(n1229), .ZN(n1251) );
NAND3_X1 U923 ( .A1(n1072), .A2(n1260), .A3(n1079), .ZN(n1229) );
INV_X1 U924 ( .A(n1060), .ZN(n1090) );
NAND2_X1 U925 ( .A1(n1099), .A2(n1112), .ZN(n1060) );
XOR2_X1 U926 ( .A(n1261), .B(KEYINPUT62), .Z(n1099) );
NAND4_X1 U927 ( .A1(n1262), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(G30) );
OR3_X1 U928 ( .A1(G128), .A2(KEYINPUT43), .A3(KEYINPUT58), .ZN(n1265) );
NAND2_X1 U929 ( .A1(n1266), .A2(KEYINPUT58), .ZN(n1264) );
XNOR2_X1 U930 ( .A(KEYINPUT43), .B(n1267), .ZN(n1266) );
NAND3_X1 U931 ( .A1(n1268), .A2(KEYINPUT43), .A3(n1269), .ZN(n1263) );
OR2_X1 U932 ( .A1(n1269), .A2(n1268), .ZN(n1262) );
NOR2_X1 U933 ( .A1(n1267), .A2(KEYINPUT58), .ZN(n1268) );
NAND3_X1 U934 ( .A1(n1092), .A2(n1230), .A3(n1237), .ZN(n1269) );
INV_X1 U935 ( .A(n1231), .ZN(n1237) );
NAND4_X1 U936 ( .A1(n1270), .A2(n1072), .A3(n1121), .A4(n1260), .ZN(n1231) );
XOR2_X1 U937 ( .A(G101), .B(n1247), .Z(G3) );
AND3_X1 U938 ( .A1(n1065), .A2(n1248), .A3(n1079), .ZN(n1247) );
XNOR2_X1 U939 ( .A(G125), .B(n1215), .ZN(G27) );
NAND4_X1 U940 ( .A1(n1271), .A2(n1254), .A3(n1230), .A4(n1077), .ZN(n1215) );
AND4_X1 U941 ( .A1(n1272), .A2(n1091), .A3(n1121), .A4(n1260), .ZN(n1254) );
NAND2_X1 U942 ( .A1(n1273), .A2(n1067), .ZN(n1260) );
NAND3_X1 U943 ( .A1(G902), .A2(n1274), .A3(n1139), .ZN(n1273) );
NOR2_X1 U944 ( .A1(n1083), .A2(G900), .ZN(n1139) );
XNOR2_X1 U945 ( .A(n1275), .B(n1246), .ZN(G24) );
AND3_X1 U946 ( .A1(n1276), .A2(n1073), .A3(n1238), .ZN(n1246) );
AND2_X1 U947 ( .A1(n1277), .A2(n1278), .ZN(n1238) );
INV_X1 U948 ( .A(n1086), .ZN(n1073) );
NAND2_X1 U949 ( .A1(n1279), .A2(n1272), .ZN(n1086) );
NAND3_X1 U950 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(G21) );
NAND2_X1 U951 ( .A1(G119), .A2(n1240), .ZN(n1282) );
NAND2_X1 U952 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
INV_X1 U953 ( .A(KEYINPUT15), .ZN(n1284) );
NAND2_X1 U954 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
XNOR2_X1 U955 ( .A(KEYINPUT11), .B(n1287), .ZN(n1286) );
NAND2_X1 U956 ( .A1(KEYINPUT15), .A2(n1288), .ZN(n1280) );
NAND2_X1 U957 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
OR2_X1 U958 ( .A1(n1287), .A2(KEYINPUT11), .ZN(n1290) );
NAND3_X1 U959 ( .A1(n1285), .A2(n1287), .A3(KEYINPUT11), .ZN(n1289) );
INV_X1 U960 ( .A(n1240), .ZN(n1285) );
NAND4_X1 U961 ( .A1(n1270), .A2(n1276), .A3(n1065), .A4(n1121), .ZN(n1240) );
XNOR2_X1 U962 ( .A(n1245), .B(n1291), .ZN(G18) );
NAND2_X1 U963 ( .A1(KEYINPUT4), .A2(G116), .ZN(n1291) );
AND3_X1 U964 ( .A1(n1079), .A2(n1092), .A3(n1276), .ZN(n1245) );
NOR2_X1 U965 ( .A1(n1278), .A2(n1101), .ZN(n1092) );
XOR2_X1 U966 ( .A(G113), .B(n1244), .Z(G15) );
AND3_X1 U967 ( .A1(n1079), .A2(n1091), .A3(n1276), .ZN(n1244) );
AND3_X1 U968 ( .A1(n1292), .A2(n1077), .A3(n1271), .ZN(n1276) );
XOR2_X1 U969 ( .A(n1066), .B(KEYINPUT49), .Z(n1077) );
AND2_X1 U970 ( .A1(n1101), .A2(n1278), .ZN(n1091) );
INV_X1 U971 ( .A(n1277), .ZN(n1101) );
AND2_X1 U972 ( .A1(n1279), .A2(n1270), .ZN(n1079) );
XNOR2_X1 U973 ( .A(n1081), .B(KEYINPUT1), .ZN(n1270) );
XNOR2_X1 U974 ( .A(KEYINPUT17), .B(n1121), .ZN(n1279) );
XNOR2_X1 U975 ( .A(n1243), .B(n1293), .ZN(G12) );
XNOR2_X1 U976 ( .A(G110), .B(KEYINPUT29), .ZN(n1293) );
AND4_X1 U977 ( .A1(n1065), .A2(n1248), .A3(n1272), .A4(n1121), .ZN(n1243) );
XOR2_X1 U978 ( .A(n1294), .B(n1167), .Z(n1121) );
NAND2_X1 U979 ( .A1(G217), .A2(n1295), .ZN(n1167) );
NAND2_X1 U980 ( .A1(n1165), .A2(n1213), .ZN(n1294) );
XNOR2_X1 U981 ( .A(n1296), .B(n1297), .ZN(n1165) );
XOR2_X1 U982 ( .A(G137), .B(n1298), .Z(n1297) );
NOR2_X1 U983 ( .A1(KEYINPUT25), .A2(n1299), .ZN(n1298) );
XOR2_X1 U984 ( .A(n1300), .B(n1145), .Z(n1299) );
NAND2_X1 U985 ( .A1(n1301), .A2(KEYINPUT60), .ZN(n1300) );
XNOR2_X1 U986 ( .A(G110), .B(n1302), .ZN(n1301) );
XNOR2_X1 U987 ( .A(n1267), .B(G119), .ZN(n1302) );
NAND2_X1 U988 ( .A1(n1303), .A2(G221), .ZN(n1296) );
INV_X1 U989 ( .A(n1081), .ZN(n1272) );
XOR2_X1 U990 ( .A(n1116), .B(n1117), .Z(n1081) );
INV_X1 U991 ( .A(G472), .ZN(n1117) );
NAND2_X1 U992 ( .A1(n1304), .A2(n1213), .ZN(n1116) );
XOR2_X1 U993 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U994 ( .A(G137), .B(n1307), .Z(n1306) );
NOR2_X1 U995 ( .A1(KEYINPUT54), .A2(n1206), .ZN(n1307) );
INV_X1 U996 ( .A(n1308), .ZN(n1206) );
XOR2_X1 U997 ( .A(n1187), .B(n1309), .Z(n1305) );
XOR2_X1 U998 ( .A(n1310), .B(n1311), .Z(n1187) );
XOR2_X1 U999 ( .A(n1312), .B(n1313), .Z(n1311) );
NOR3_X1 U1000 ( .A1(n1212), .A2(G953), .A3(G237), .ZN(n1312) );
INV_X1 U1001 ( .A(G210), .ZN(n1212) );
XNOR2_X1 U1002 ( .A(G116), .B(n1314), .ZN(n1310) );
XNOR2_X1 U1003 ( .A(KEYINPUT38), .B(n1287), .ZN(n1314) );
AND2_X1 U1004 ( .A1(n1292), .A2(n1072), .ZN(n1248) );
NOR2_X1 U1005 ( .A1(n1271), .A2(n1066), .ZN(n1072) );
AND2_X1 U1006 ( .A1(G221), .A2(n1295), .ZN(n1066) );
NAND2_X1 U1007 ( .A1(G234), .A2(n1213), .ZN(n1295) );
INV_X1 U1008 ( .A(n1074), .ZN(n1271) );
XNOR2_X1 U1009 ( .A(n1107), .B(n1315), .ZN(n1074) );
XNOR2_X1 U1010 ( .A(KEYINPUT22), .B(n1108), .ZN(n1315) );
INV_X1 U1011 ( .A(G469), .ZN(n1108) );
NAND2_X1 U1012 ( .A1(n1316), .A2(n1213), .ZN(n1107) );
XOR2_X1 U1013 ( .A(KEYINPUT40), .B(n1196), .Z(n1316) );
XNOR2_X1 U1014 ( .A(n1317), .B(n1318), .ZN(n1196) );
XOR2_X1 U1015 ( .A(n1319), .B(n1320), .Z(n1318) );
XNOR2_X1 U1016 ( .A(G101), .B(n1321), .ZN(n1320) );
NOR2_X1 U1017 ( .A1(G107), .A2(KEYINPUT45), .ZN(n1321) );
XNOR2_X1 U1018 ( .A(G110), .B(G104), .ZN(n1319) );
XOR2_X1 U1019 ( .A(n1188), .B(n1322), .Z(n1317) );
XOR2_X1 U1020 ( .A(n1323), .B(n1324), .Z(n1322) );
AND2_X1 U1021 ( .A1(n1083), .A2(G227), .ZN(n1323) );
XOR2_X1 U1022 ( .A(n1144), .B(n1309), .Z(n1188) );
XOR2_X1 U1023 ( .A(n1325), .B(n1326), .Z(n1309) );
NOR2_X1 U1024 ( .A1(G131), .A2(KEYINPUT47), .ZN(n1326) );
NOR2_X1 U1025 ( .A1(G134), .A2(KEYINPUT63), .ZN(n1325) );
XNOR2_X1 U1026 ( .A(G137), .B(n1327), .ZN(n1144) );
AND2_X1 U1027 ( .A1(n1230), .A2(n1328), .ZN(n1292) );
NAND2_X1 U1028 ( .A1(n1067), .A2(n1329), .ZN(n1328) );
NAND4_X1 U1029 ( .A1(G902), .A2(G953), .A3(n1274), .A4(n1153), .ZN(n1329) );
INV_X1 U1030 ( .A(G898), .ZN(n1153) );
NAND3_X1 U1031 ( .A1(n1274), .A2(n1083), .A3(G952), .ZN(n1067) );
NAND2_X1 U1032 ( .A1(G237), .A2(G234), .ZN(n1274) );
INV_X1 U1033 ( .A(n1095), .ZN(n1230) );
NAND2_X1 U1034 ( .A1(n1261), .A2(n1112), .ZN(n1095) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1330), .ZN(n1112) );
XNOR2_X1 U1036 ( .A(n1120), .B(n1331), .ZN(n1261) );
NOR2_X1 U1037 ( .A1(n1118), .A2(KEYINPUT3), .ZN(n1331) );
AND2_X1 U1038 ( .A1(n1332), .A2(n1213), .ZN(n1118) );
XOR2_X1 U1039 ( .A(KEYINPUT27), .B(n1333), .Z(n1332) );
NOR2_X1 U1040 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NOR2_X1 U1041 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XNOR2_X1 U1042 ( .A(KEYINPUT8), .B(n1338), .ZN(n1337) );
AND2_X1 U1043 ( .A1(n1338), .A2(n1336), .ZN(n1334) );
XNOR2_X1 U1044 ( .A(n1339), .B(n1340), .ZN(n1336) );
XNOR2_X1 U1045 ( .A(KEYINPUT44), .B(n1209), .ZN(n1340) );
INV_X1 U1046 ( .A(G125), .ZN(n1209) );
XNOR2_X1 U1047 ( .A(n1341), .B(n1210), .ZN(n1339) );
NAND2_X1 U1048 ( .A1(G224), .A2(n1342), .ZN(n1210) );
XNOR2_X1 U1049 ( .A(KEYINPUT2), .B(n1083), .ZN(n1342) );
NAND2_X1 U1050 ( .A1(KEYINPUT48), .A2(n1308), .ZN(n1341) );
XOR2_X1 U1051 ( .A(n1327), .B(n1190), .Z(n1308) );
XOR2_X1 U1052 ( .A(G146), .B(KEYINPUT35), .Z(n1190) );
INV_X1 U1053 ( .A(n1202), .ZN(n1338) );
XNOR2_X1 U1054 ( .A(n1343), .B(n1344), .ZN(n1202) );
XOR2_X1 U1055 ( .A(n1161), .B(n1345), .Z(n1344) );
NOR2_X1 U1056 ( .A1(KEYINPUT46), .A2(n1154), .ZN(n1345) );
XNOR2_X1 U1057 ( .A(n1346), .B(n1347), .ZN(n1154) );
INV_X1 U1058 ( .A(G110), .ZN(n1347) );
NAND2_X1 U1059 ( .A1(KEYINPUT5), .A2(n1275), .ZN(n1346) );
NOR3_X1 U1060 ( .A1(KEYINPUT59), .A2(n1348), .A3(n1349), .ZN(n1161) );
XOR2_X1 U1061 ( .A(n1350), .B(KEYINPUT32), .Z(n1349) );
NAND2_X1 U1062 ( .A1(G116), .A2(n1287), .ZN(n1350) );
NOR2_X1 U1063 ( .A1(G116), .A2(n1287), .ZN(n1348) );
INV_X1 U1064 ( .A(G119), .ZN(n1287) );
XNOR2_X1 U1065 ( .A(n1158), .B(n1313), .ZN(n1343) );
XOR2_X1 U1066 ( .A(G101), .B(G113), .Z(n1313) );
XNOR2_X1 U1067 ( .A(n1351), .B(G104), .ZN(n1158) );
NAND2_X1 U1068 ( .A1(KEYINPUT52), .A2(G107), .ZN(n1351) );
AND2_X1 U1069 ( .A1(n1352), .A2(G210), .ZN(n1120) );
XOR2_X1 U1070 ( .A(n1330), .B(KEYINPUT28), .Z(n1352) );
NAND2_X1 U1071 ( .A1(n1213), .A2(n1353), .ZN(n1330) );
INV_X1 U1072 ( .A(G902), .ZN(n1213) );
NOR2_X1 U1073 ( .A1(n1277), .A2(n1278), .ZN(n1065) );
NAND3_X1 U1074 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1278) );
NAND2_X1 U1075 ( .A1(G475), .A2(n1357), .ZN(n1356) );
INV_X1 U1076 ( .A(n1109), .ZN(n1357) );
NAND2_X1 U1077 ( .A1(KEYINPUT16), .A2(n1358), .ZN(n1355) );
NAND2_X1 U1078 ( .A1(n1359), .A2(n1111), .ZN(n1358) );
XNOR2_X1 U1079 ( .A(n1109), .B(KEYINPUT14), .ZN(n1359) );
NAND2_X1 U1080 ( .A1(n1360), .A2(n1361), .ZN(n1354) );
INV_X1 U1081 ( .A(KEYINPUT16), .ZN(n1361) );
NAND2_X1 U1082 ( .A1(n1362), .A2(n1363), .ZN(n1360) );
OR2_X1 U1083 ( .A1(n1109), .A2(KEYINPUT14), .ZN(n1363) );
NAND3_X1 U1084 ( .A1(n1109), .A2(n1111), .A3(KEYINPUT14), .ZN(n1362) );
INV_X1 U1085 ( .A(G475), .ZN(n1111) );
NOR2_X1 U1086 ( .A1(n1179), .A2(G902), .ZN(n1109) );
INV_X1 U1087 ( .A(n1177), .ZN(n1179) );
XNOR2_X1 U1088 ( .A(n1364), .B(n1365), .ZN(n1177) );
XOR2_X1 U1089 ( .A(n1366), .B(n1367), .Z(n1365) );
NOR2_X1 U1090 ( .A1(KEYINPUT61), .A2(n1145), .ZN(n1367) );
XNOR2_X1 U1091 ( .A(G125), .B(n1324), .ZN(n1145) );
XOR2_X1 U1092 ( .A(G140), .B(G146), .Z(n1324) );
NOR2_X1 U1093 ( .A1(n1368), .A2(n1369), .ZN(n1366) );
XOR2_X1 U1094 ( .A(KEYINPUT6), .B(n1370), .Z(n1369) );
NOR2_X1 U1095 ( .A1(G104), .A2(n1371), .ZN(n1370) );
INV_X1 U1096 ( .A(n1372), .ZN(n1371) );
NOR2_X1 U1097 ( .A1(n1372), .A2(n1373), .ZN(n1368) );
XNOR2_X1 U1098 ( .A(G104), .B(KEYINPUT34), .ZN(n1373) );
XOR2_X1 U1099 ( .A(G113), .B(n1275), .Z(n1372) );
XNOR2_X1 U1100 ( .A(G131), .B(n1374), .ZN(n1364) );
NOR2_X1 U1101 ( .A1(KEYINPUT18), .A2(n1375), .ZN(n1374) );
XNOR2_X1 U1102 ( .A(G143), .B(n1376), .ZN(n1375) );
AND3_X1 U1103 ( .A1(G214), .A2(n1083), .A3(n1353), .ZN(n1376) );
INV_X1 U1104 ( .A(G237), .ZN(n1353) );
XNOR2_X1 U1105 ( .A(n1377), .B(G478), .ZN(n1277) );
OR2_X1 U1106 ( .A1(n1171), .A2(G902), .ZN(n1377) );
XNOR2_X1 U1107 ( .A(n1378), .B(n1379), .ZN(n1171) );
XOR2_X1 U1108 ( .A(G107), .B(n1380), .Z(n1379) );
XNOR2_X1 U1109 ( .A(n1275), .B(G116), .ZN(n1380) );
INV_X1 U1110 ( .A(G122), .ZN(n1275) );
XOR2_X1 U1111 ( .A(n1381), .B(n1382), .Z(n1378) );
NOR2_X1 U1112 ( .A1(KEYINPUT9), .A2(n1383), .ZN(n1382) );
XNOR2_X1 U1113 ( .A(n1143), .B(n1327), .ZN(n1383) );
XNOR2_X1 U1114 ( .A(G143), .B(n1267), .ZN(n1327) );
INV_X1 U1115 ( .A(G128), .ZN(n1267) );
INV_X1 U1116 ( .A(G134), .ZN(n1143) );
NAND2_X1 U1117 ( .A1(G217), .A2(n1303), .ZN(n1381) );
AND2_X1 U1118 ( .A1(G234), .A2(n1083), .ZN(n1303) );
INV_X1 U1119 ( .A(G953), .ZN(n1083) );
endmodule


