//Key = 0100001000011011011111111111001011101111011000010000010000000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;

XNOR2_X1 U738 ( .A(n1010), .B(n1011), .ZN(G9) );
XOR2_X1 U739 ( .A(n1012), .B(KEYINPUT6), .Z(n1010) );
NAND3_X1 U740 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(G75) );
NOR3_X1 U741 ( .A1(n1016), .A2(G953), .A3(n1017), .ZN(n1015) );
NOR3_X1 U742 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NAND3_X1 U743 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1018) );
NAND2_X1 U744 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NAND2_X1 U745 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U746 ( .A1(n1028), .A2(n1029), .ZN(n1016) );
NOR2_X1 U747 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NOR4_X1 U748 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
XOR2_X1 U749 ( .A(n1036), .B(n1037), .Z(n1035) );
XNOR2_X1 U750 ( .A(KEYINPUT62), .B(n1038), .ZN(n1036) );
NOR2_X1 U751 ( .A1(KEYINPUT4), .A2(n1039), .ZN(n1038) );
XOR2_X1 U752 ( .A(n1040), .B(n1041), .Z(n1034) );
NOR2_X1 U753 ( .A1(G478), .A2(KEYINPUT52), .ZN(n1041) );
NAND3_X1 U754 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1032) );
XOR2_X1 U755 ( .A(KEYINPUT41), .B(n1045), .Z(n1044) );
NAND2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1042) );
NOR3_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1020), .ZN(n1030) );
NOR2_X1 U758 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND3_X1 U759 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1048) );
NAND2_X1 U760 ( .A1(n1055), .A2(n1033), .ZN(n1054) );
NAND4_X1 U761 ( .A1(n1043), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1053) );
NOR3_X1 U762 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NAND2_X1 U763 ( .A1(n1062), .A2(n1019), .ZN(n1052) );
NAND2_X1 U764 ( .A1(n1023), .A2(n1021), .ZN(n1062) );
INV_X1 U765 ( .A(n1063), .ZN(n1013) );
XOR2_X1 U766 ( .A(n1064), .B(n1065), .Z(G72) );
NAND2_X1 U767 ( .A1(G953), .A2(n1066), .ZN(n1065) );
NAND2_X1 U768 ( .A1(G900), .A2(G227), .ZN(n1066) );
NAND2_X1 U769 ( .A1(KEYINPUT33), .A2(n1067), .ZN(n1064) );
XOR2_X1 U770 ( .A(n1068), .B(n1069), .Z(n1067) );
NAND2_X1 U771 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U772 ( .A1(G953), .A2(n1072), .ZN(n1071) );
XOR2_X1 U773 ( .A(n1073), .B(n1074), .Z(n1070) );
XOR2_X1 U774 ( .A(KEYINPUT47), .B(n1075), .Z(n1074) );
NOR2_X1 U775 ( .A1(KEYINPUT63), .A2(n1076), .ZN(n1075) );
XOR2_X1 U776 ( .A(n1077), .B(n1078), .Z(n1073) );
NAND2_X1 U777 ( .A1(n1079), .A2(n1063), .ZN(n1068) );
XOR2_X1 U778 ( .A(n1080), .B(KEYINPUT5), .Z(n1079) );
XOR2_X1 U779 ( .A(n1081), .B(n1082), .Z(G69) );
XOR2_X1 U780 ( .A(n1083), .B(n1084), .Z(n1082) );
NAND2_X1 U781 ( .A1(G953), .A2(n1085), .ZN(n1084) );
NAND2_X1 U782 ( .A1(G898), .A2(G224), .ZN(n1085) );
NAND2_X1 U783 ( .A1(n1086), .A2(n1087), .ZN(n1083) );
NAND2_X1 U784 ( .A1(G953), .A2(n1088), .ZN(n1087) );
XOR2_X1 U785 ( .A(n1089), .B(n1090), .Z(n1086) );
XOR2_X1 U786 ( .A(n1091), .B(n1092), .Z(n1090) );
XOR2_X1 U787 ( .A(n1093), .B(n1094), .Z(n1089) );
NOR2_X1 U788 ( .A1(n1014), .A2(G953), .ZN(n1081) );
INV_X1 U789 ( .A(n1095), .ZN(n1014) );
NOR2_X1 U790 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XNOR2_X1 U791 ( .A(n1098), .B(n1099), .ZN(n1097) );
NOR4_X1 U792 ( .A1(n1100), .A2(n1101), .A3(KEYINPUT8), .A4(n1102), .ZN(n1099) );
NOR2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR3_X1 U794 ( .A1(n1105), .A2(n1106), .A3(n1095), .ZN(n1103) );
AND2_X1 U795 ( .A1(n1104), .A2(n1107), .ZN(n1100) );
INV_X1 U796 ( .A(KEYINPUT61), .ZN(n1104) );
NOR3_X1 U797 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(G63) );
AND3_X1 U798 ( .A1(KEYINPUT59), .A2(G953), .A3(G952), .ZN(n1110) );
NOR2_X1 U799 ( .A1(KEYINPUT59), .A2(n1111), .ZN(n1109) );
INV_X1 U800 ( .A(n1096), .ZN(n1111) );
XOR2_X1 U801 ( .A(n1112), .B(n1113), .Z(n1108) );
NOR2_X1 U802 ( .A1(n1114), .A2(n1107), .ZN(n1113) );
NAND2_X1 U803 ( .A1(KEYINPUT15), .A2(n1115), .ZN(n1112) );
NOR2_X1 U804 ( .A1(n1096), .A2(n1116), .ZN(G60) );
XOR2_X1 U805 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U806 ( .A1(n1047), .A2(n1107), .ZN(n1118) );
XNOR2_X1 U807 ( .A(G104), .B(n1119), .ZN(G6) );
NOR2_X1 U808 ( .A1(n1096), .A2(n1120), .ZN(G57) );
XOR2_X1 U809 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U811 ( .A1(KEYINPUT16), .A2(n1125), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1126), .A2(n1107), .ZN(n1123) );
INV_X1 U813 ( .A(G472), .ZN(n1126) );
XOR2_X1 U814 ( .A(n1127), .B(n1128), .Z(n1121) );
NOR2_X1 U815 ( .A1(n1096), .A2(n1129), .ZN(G54) );
XOR2_X1 U816 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U817 ( .A(n1132), .B(n1133), .Z(n1131) );
XNOR2_X1 U818 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR2_X1 U819 ( .A1(G110), .A2(n1136), .ZN(n1135) );
XOR2_X1 U820 ( .A(KEYINPUT29), .B(KEYINPUT13), .Z(n1136) );
XOR2_X1 U821 ( .A(n1137), .B(KEYINPUT28), .Z(n1132) );
XOR2_X1 U822 ( .A(n1138), .B(n1139), .Z(n1130) );
XOR2_X1 U823 ( .A(n1140), .B(n1078), .Z(n1139) );
NOR2_X1 U824 ( .A1(n1141), .A2(n1107), .ZN(n1140) );
INV_X1 U825 ( .A(G469), .ZN(n1141) );
NOR2_X1 U826 ( .A1(n1096), .A2(n1142), .ZN(G51) );
XOR2_X1 U827 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U828 ( .A1(n1145), .A2(n1107), .ZN(n1144) );
NAND2_X1 U829 ( .A1(G902), .A2(n1146), .ZN(n1107) );
OR2_X1 U830 ( .A1(n1105), .A2(n1095), .ZN(n1146) );
NAND4_X1 U831 ( .A1(n1147), .A2(n1011), .A3(n1148), .A4(n1149), .ZN(n1095) );
AND4_X1 U832 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1119), .ZN(n1149) );
NAND3_X1 U833 ( .A1(n1153), .A2(n1021), .A3(n1061), .ZN(n1119) );
INV_X1 U834 ( .A(n1154), .ZN(n1151) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1156), .ZN(n1148) );
NOR2_X1 U836 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U837 ( .A(n1159), .B(KEYINPUT60), .Z(n1157) );
NAND3_X1 U838 ( .A1(n1021), .A2(n1160), .A3(n1153), .ZN(n1011) );
XNOR2_X1 U839 ( .A(n1063), .B(KEYINPUT30), .ZN(n1105) );
NAND4_X1 U840 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1063) );
NOR4_X1 U841 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
INV_X1 U842 ( .A(n1169), .ZN(n1168) );
INV_X1 U843 ( .A(n1170), .ZN(n1165) );
NAND3_X1 U844 ( .A1(n1171), .A2(n1172), .A3(n1061), .ZN(n1163) );
NAND2_X1 U845 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
OR2_X1 U846 ( .A1(n1175), .A2(KEYINPUT18), .ZN(n1173) );
NAND3_X1 U847 ( .A1(n1176), .A2(n1177), .A3(n1059), .ZN(n1171) );
NAND3_X1 U848 ( .A1(n1050), .A2(n1178), .A3(n1179), .ZN(n1177) );
NAND2_X1 U849 ( .A1(KEYINPUT18), .A2(n1180), .ZN(n1176) );
NAND3_X1 U850 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(n1143) );
NAND2_X1 U851 ( .A1(KEYINPUT57), .A2(n1184), .ZN(n1183) );
INV_X1 U852 ( .A(n1185), .ZN(n1184) );
OR3_X1 U853 ( .A1(n1186), .A2(KEYINPUT57), .A3(n1187), .ZN(n1182) );
NAND2_X1 U854 ( .A1(n1187), .A2(n1186), .ZN(n1181) );
NAND2_X1 U855 ( .A1(KEYINPUT38), .A2(n1185), .ZN(n1186) );
NAND2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
NOR2_X1 U857 ( .A1(n1080), .A2(G952), .ZN(n1096) );
XOR2_X1 U858 ( .A(n1190), .B(n1161), .Z(G48) );
NAND3_X1 U859 ( .A1(n1191), .A2(n1192), .A3(n1061), .ZN(n1161) );
XNOR2_X1 U860 ( .A(G143), .B(n1162), .ZN(G45) );
NAND3_X1 U861 ( .A1(n1060), .A2(n1191), .A3(n1193), .ZN(n1162) );
XOR2_X1 U862 ( .A(G140), .B(n1194), .Z(G42) );
NOR3_X1 U863 ( .A1(n1174), .A2(n1175), .A3(n1159), .ZN(n1194) );
INV_X1 U864 ( .A(n1059), .ZN(n1174) );
XOR2_X1 U865 ( .A(n1195), .B(G137), .Z(G39) );
NAND2_X1 U866 ( .A1(KEYINPUT19), .A2(n1169), .ZN(n1195) );
NAND3_X1 U867 ( .A1(n1180), .A2(n1192), .A3(n1196), .ZN(n1169) );
XOR2_X1 U868 ( .A(n1167), .B(n1197), .Z(G36) );
NOR2_X1 U869 ( .A1(KEYINPUT56), .A2(n1198), .ZN(n1197) );
AND3_X1 U870 ( .A1(n1180), .A2(n1160), .A3(n1060), .ZN(n1167) );
XOR2_X1 U871 ( .A(n1199), .B(n1166), .Z(G33) );
AND3_X1 U872 ( .A1(n1061), .A2(n1180), .A3(n1060), .ZN(n1166) );
INV_X1 U873 ( .A(n1175), .ZN(n1180) );
NAND3_X1 U874 ( .A1(n1200), .A2(n1178), .A3(n1023), .ZN(n1175) );
INV_X1 U875 ( .A(n1055), .ZN(n1023) );
NAND2_X1 U876 ( .A1(n1051), .A2(n1043), .ZN(n1055) );
INV_X1 U877 ( .A(n1201), .ZN(n1051) );
XNOR2_X1 U878 ( .A(G131), .B(KEYINPUT24), .ZN(n1199) );
XOR2_X1 U879 ( .A(n1202), .B(n1170), .Z(G30) );
NAND3_X1 U880 ( .A1(n1192), .A2(n1160), .A3(n1191), .ZN(n1170) );
NOR3_X1 U881 ( .A1(n1056), .A2(n1203), .A3(n1024), .ZN(n1191) );
INV_X1 U882 ( .A(n1200), .ZN(n1024) );
INV_X1 U883 ( .A(n1057), .ZN(n1160) );
XNOR2_X1 U884 ( .A(n1155), .B(n1204), .ZN(G3) );
NAND2_X1 U885 ( .A1(G101), .A2(n1205), .ZN(n1204) );
XOR2_X1 U886 ( .A(KEYINPUT9), .B(KEYINPUT32), .Z(n1205) );
AND3_X1 U887 ( .A1(n1060), .A2(n1153), .A3(n1196), .ZN(n1155) );
XNOR2_X1 U888 ( .A(G125), .B(n1206), .ZN(G27) );
NAND3_X1 U889 ( .A1(n1207), .A2(n1059), .A3(n1208), .ZN(n1206) );
NOR3_X1 U890 ( .A1(n1029), .A2(n1203), .A3(n1056), .ZN(n1208) );
INV_X1 U891 ( .A(n1178), .ZN(n1203) );
NAND2_X1 U892 ( .A1(n1020), .A2(n1209), .ZN(n1178) );
NAND2_X1 U893 ( .A1(n1210), .A2(n1072), .ZN(n1209) );
INV_X1 U894 ( .A(G900), .ZN(n1072) );
XOR2_X1 U895 ( .A(n1159), .B(KEYINPUT1), .Z(n1207) );
XNOR2_X1 U896 ( .A(G122), .B(n1147), .ZN(G24) );
NAND4_X1 U897 ( .A1(n1179), .A2(n1193), .A3(n1021), .A4(n1211), .ZN(n1147) );
INV_X1 U898 ( .A(n1033), .ZN(n1021) );
NAND2_X1 U899 ( .A1(n1212), .A2(n1213), .ZN(n1033) );
AND2_X1 U900 ( .A1(n1214), .A2(n1215), .ZN(n1193) );
XOR2_X1 U901 ( .A(KEYINPUT21), .B(n1216), .Z(n1214) );
XOR2_X1 U902 ( .A(n1217), .B(n1152), .Z(G21) );
NAND4_X1 U903 ( .A1(n1179), .A2(n1196), .A3(n1192), .A4(n1211), .ZN(n1152) );
NOR2_X1 U904 ( .A1(n1213), .A2(n1212), .ZN(n1192) );
NAND2_X1 U905 ( .A1(n1218), .A2(n1219), .ZN(G18) );
NAND2_X1 U906 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NAND2_X1 U907 ( .A1(n1154), .A2(n1222), .ZN(n1221) );
NAND2_X1 U908 ( .A1(KEYINPUT51), .A2(KEYINPUT20), .ZN(n1222) );
OR3_X1 U909 ( .A1(n1223), .A2(KEYINPUT51), .A3(n1220), .ZN(n1218) );
XOR2_X1 U910 ( .A(G116), .B(KEYINPUT0), .Z(n1220) );
XOR2_X1 U911 ( .A(KEYINPUT20), .B(n1154), .Z(n1223) );
NOR2_X1 U912 ( .A1(n1158), .A2(n1057), .ZN(n1154) );
NAND2_X1 U913 ( .A1(n1216), .A2(n1215), .ZN(n1057) );
XOR2_X1 U914 ( .A(G113), .B(n1224), .Z(G15) );
NOR2_X1 U915 ( .A1(n1159), .A2(n1158), .ZN(n1224) );
NAND3_X1 U916 ( .A1(n1060), .A2(n1211), .A3(n1179), .ZN(n1158) );
INV_X1 U917 ( .A(n1029), .ZN(n1179) );
NAND2_X1 U918 ( .A1(n1027), .A2(n1225), .ZN(n1029) );
AND2_X1 U919 ( .A1(n1213), .A2(n1226), .ZN(n1060) );
INV_X1 U920 ( .A(n1061), .ZN(n1159) );
NOR2_X1 U921 ( .A1(n1215), .A2(n1216), .ZN(n1061) );
XOR2_X1 U922 ( .A(n1150), .B(n1227), .Z(G12) );
XOR2_X1 U923 ( .A(KEYINPUT25), .B(G110), .Z(n1227) );
NAND3_X1 U924 ( .A1(n1196), .A2(n1153), .A3(n1059), .ZN(n1150) );
NOR2_X1 U925 ( .A1(n1226), .A2(n1213), .ZN(n1059) );
XNOR2_X1 U926 ( .A(n1228), .B(n1102), .ZN(n1213) );
NAND2_X1 U927 ( .A1(G217), .A2(n1229), .ZN(n1102) );
NAND2_X1 U928 ( .A1(n1098), .A2(n1106), .ZN(n1228) );
XNOR2_X1 U929 ( .A(n1230), .B(n1231), .ZN(n1098) );
XOR2_X1 U930 ( .A(n1232), .B(n1076), .Z(n1231) );
NOR2_X1 U931 ( .A1(KEYINPUT7), .A2(n1233), .ZN(n1232) );
XOR2_X1 U932 ( .A(n1234), .B(n1235), .Z(n1233) );
XOR2_X1 U933 ( .A(KEYINPUT49), .B(G128), .Z(n1235) );
XOR2_X1 U934 ( .A(n1217), .B(G110), .Z(n1234) );
XOR2_X1 U935 ( .A(n1190), .B(n1236), .Z(n1230) );
NOR2_X1 U936 ( .A1(KEYINPUT2), .A2(n1237), .ZN(n1236) );
XOR2_X1 U937 ( .A(n1238), .B(n1239), .Z(n1237) );
AND2_X1 U938 ( .A1(G221), .A2(n1240), .ZN(n1239) );
INV_X1 U939 ( .A(G137), .ZN(n1238) );
INV_X1 U940 ( .A(n1212), .ZN(n1226) );
XOR2_X1 U941 ( .A(n1241), .B(G472), .Z(n1212) );
NAND2_X1 U942 ( .A1(n1242), .A2(n1106), .ZN(n1241) );
XOR2_X1 U943 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U944 ( .A(KEYINPUT31), .B(n1245), .Z(n1244) );
NOR2_X1 U945 ( .A1(KEYINPUT54), .A2(n1128), .ZN(n1245) );
XNOR2_X1 U946 ( .A(n1246), .B(n1247), .ZN(n1128) );
XOR2_X1 U947 ( .A(G119), .B(G116), .Z(n1247) );
NAND2_X1 U948 ( .A1(KEYINPUT53), .A2(n1248), .ZN(n1246) );
XNOR2_X1 U949 ( .A(n1127), .B(n1125), .ZN(n1243) );
XNOR2_X1 U950 ( .A(n1249), .B(n1250), .ZN(n1125) );
NAND3_X1 U951 ( .A1(n1251), .A2(n1252), .A3(G210), .ZN(n1249) );
XOR2_X1 U952 ( .A(n1253), .B(n1254), .Z(n1127) );
AND2_X1 U953 ( .A1(n1211), .A2(n1200), .ZN(n1153) );
NOR2_X1 U954 ( .A1(n1027), .A2(n1026), .ZN(n1200) );
INV_X1 U955 ( .A(n1225), .ZN(n1026) );
NAND2_X1 U956 ( .A1(G221), .A2(n1229), .ZN(n1225) );
NAND2_X1 U957 ( .A1(G234), .A2(n1106), .ZN(n1229) );
XOR2_X1 U958 ( .A(n1255), .B(G469), .Z(n1027) );
NAND2_X1 U959 ( .A1(n1256), .A2(n1106), .ZN(n1255) );
XOR2_X1 U960 ( .A(n1257), .B(n1258), .Z(n1256) );
XOR2_X1 U961 ( .A(n1259), .B(n1260), .Z(n1258) );
NAND3_X1 U962 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1260) );
NAND2_X1 U963 ( .A1(KEYINPUT46), .A2(n1134), .ZN(n1263) );
NAND3_X1 U964 ( .A1(n1264), .A2(n1265), .A3(n1078), .ZN(n1262) );
INV_X1 U965 ( .A(KEYINPUT46), .ZN(n1265) );
OR2_X1 U966 ( .A1(n1078), .A2(n1264), .ZN(n1261) );
NOR2_X1 U967 ( .A1(n1134), .A2(KEYINPUT58), .ZN(n1264) );
AND2_X1 U968 ( .A1(n1266), .A2(n1267), .ZN(n1134) );
NAND2_X1 U969 ( .A1(n1268), .A2(n1250), .ZN(n1267) );
XOR2_X1 U970 ( .A(G107), .B(n1269), .Z(n1268) );
NAND2_X1 U971 ( .A1(n1270), .A2(n1271), .ZN(n1266) );
XOR2_X1 U972 ( .A(n1012), .B(n1269), .Z(n1271) );
NOR2_X1 U973 ( .A1(KEYINPUT44), .A2(G104), .ZN(n1269) );
XOR2_X1 U974 ( .A(n1250), .B(KEYINPUT36), .Z(n1270) );
INV_X1 U975 ( .A(G101), .ZN(n1250) );
XNOR2_X1 U976 ( .A(n1272), .B(G128), .ZN(n1078) );
NAND2_X1 U977 ( .A1(KEYINPUT22), .A2(n1273), .ZN(n1272) );
XOR2_X1 U978 ( .A(G146), .B(G143), .Z(n1273) );
XOR2_X1 U979 ( .A(n1274), .B(n1275), .Z(n1257) );
INV_X1 U980 ( .A(n1138), .ZN(n1275) );
XOR2_X1 U981 ( .A(n1253), .B(n1276), .Z(n1138) );
AND2_X1 U982 ( .A1(n1251), .A2(G227), .ZN(n1276) );
XOR2_X1 U983 ( .A(n1077), .B(KEYINPUT26), .Z(n1253) );
XNOR2_X1 U984 ( .A(G131), .B(n1277), .ZN(n1077) );
XOR2_X1 U985 ( .A(G137), .B(G134), .Z(n1277) );
NAND2_X1 U986 ( .A1(KEYINPUT27), .A2(n1137), .ZN(n1274) );
INV_X1 U987 ( .A(G140), .ZN(n1137) );
AND2_X1 U988 ( .A1(n1050), .A2(n1278), .ZN(n1211) );
NAND2_X1 U989 ( .A1(n1020), .A2(n1279), .ZN(n1278) );
NAND2_X1 U990 ( .A1(n1210), .A2(n1088), .ZN(n1279) );
INV_X1 U991 ( .A(G898), .ZN(n1088) );
AND3_X1 U992 ( .A1(n1280), .A2(n1281), .A3(G953), .ZN(n1210) );
XOR2_X1 U993 ( .A(KEYINPUT10), .B(G902), .Z(n1280) );
NAND3_X1 U994 ( .A1(n1281), .A2(n1080), .A3(G952), .ZN(n1020) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1281) );
INV_X1 U996 ( .A(n1056), .ZN(n1050) );
NAND2_X1 U997 ( .A1(n1201), .A2(n1043), .ZN(n1056) );
NAND2_X1 U998 ( .A1(G214), .A2(n1282), .ZN(n1043) );
XOR2_X1 U999 ( .A(n1039), .B(n1283), .Z(n1201) );
NOR2_X1 U1000 ( .A1(n1037), .A2(KEYINPUT45), .ZN(n1283) );
INV_X1 U1001 ( .A(n1145), .ZN(n1037) );
NAND2_X1 U1002 ( .A1(G210), .A2(n1282), .ZN(n1145) );
NAND2_X1 U1003 ( .A1(n1252), .A2(n1106), .ZN(n1282) );
NAND2_X1 U1004 ( .A1(n1284), .A2(n1106), .ZN(n1039) );
XNOR2_X1 U1005 ( .A(n1285), .B(n1187), .ZN(n1284) );
XNOR2_X1 U1006 ( .A(n1286), .B(n1094), .ZN(n1187) );
NAND2_X1 U1007 ( .A1(n1287), .A2(n1288), .ZN(n1094) );
OR2_X1 U1008 ( .A1(n1259), .A2(G122), .ZN(n1288) );
XOR2_X1 U1009 ( .A(n1289), .B(KEYINPUT55), .Z(n1287) );
NAND2_X1 U1010 ( .A1(G122), .A2(n1259), .ZN(n1289) );
INV_X1 U1011 ( .A(G110), .ZN(n1259) );
NAND3_X1 U1012 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1286) );
NAND2_X1 U1013 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
NAND2_X1 U1014 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XOR2_X1 U1015 ( .A(n1093), .B(G113), .Z(n1293) );
NAND4_X1 U1016 ( .A1(n1297), .A2(n1296), .A3(KEYINPUT11), .A4(n1295), .ZN(n1291) );
INV_X1 U1017 ( .A(KEYINPUT48), .ZN(n1296) );
XOR2_X1 U1018 ( .A(n1248), .B(n1093), .Z(n1297) );
NAND2_X1 U1019 ( .A1(n1298), .A2(n1299), .ZN(n1093) );
NAND2_X1 U1020 ( .A1(n1300), .A2(n1217), .ZN(n1299) );
XNOR2_X1 U1021 ( .A(G116), .B(KEYINPUT42), .ZN(n1300) );
XOR2_X1 U1022 ( .A(KEYINPUT17), .B(n1301), .Z(n1298) );
NOR2_X1 U1023 ( .A1(n1302), .A2(n1217), .ZN(n1301) );
INV_X1 U1024 ( .A(G119), .ZN(n1217) );
XNOR2_X1 U1025 ( .A(G116), .B(KEYINPUT23), .ZN(n1302) );
OR2_X1 U1026 ( .A1(n1295), .A2(KEYINPUT11), .ZN(n1290) );
XOR2_X1 U1027 ( .A(n1092), .B(G104), .Z(n1295) );
XNOR2_X1 U1028 ( .A(n1303), .B(n1304), .ZN(n1092) );
NOR2_X1 U1029 ( .A1(KEYINPUT43), .A2(n1012), .ZN(n1304) );
NOR2_X1 U1030 ( .A1(G101), .A2(KEYINPUT35), .ZN(n1303) );
NAND2_X1 U1031 ( .A1(n1305), .A2(n1189), .ZN(n1285) );
NAND2_X1 U1032 ( .A1(n1306), .A2(n1307), .ZN(n1189) );
XNOR2_X1 U1033 ( .A(KEYINPUT34), .B(n1188), .ZN(n1305) );
OR2_X1 U1034 ( .A1(n1307), .A2(n1306), .ZN(n1188) );
XOR2_X1 U1035 ( .A(G125), .B(n1254), .Z(n1306) );
XOR2_X1 U1036 ( .A(n1190), .B(n1308), .Z(n1254) );
NAND2_X1 U1037 ( .A1(G224), .A2(n1251), .ZN(n1307) );
INV_X1 U1038 ( .A(n1019), .ZN(n1196) );
NAND2_X1 U1039 ( .A1(n1309), .A2(n1216), .ZN(n1019) );
NOR2_X1 U1040 ( .A1(n1310), .A2(n1045), .ZN(n1216) );
NOR2_X1 U1041 ( .A1(n1047), .A2(n1046), .ZN(n1045) );
AND2_X1 U1042 ( .A1(n1046), .A2(n1047), .ZN(n1310) );
INV_X1 U1043 ( .A(G475), .ZN(n1047) );
NOR2_X1 U1044 ( .A1(n1117), .A2(G902), .ZN(n1046) );
XOR2_X1 U1045 ( .A(n1091), .B(n1311), .Z(n1117) );
XOR2_X1 U1046 ( .A(G122), .B(n1312), .Z(n1311) );
NOR2_X1 U1047 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1048 ( .A(n1315), .B(KEYINPUT39), .Z(n1314) );
NAND3_X1 U1049 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1315) );
NAND2_X1 U1050 ( .A1(n1319), .A2(n1190), .ZN(n1316) );
INV_X1 U1051 ( .A(G146), .ZN(n1190) );
XNOR2_X1 U1052 ( .A(KEYINPUT40), .B(n1076), .ZN(n1319) );
NOR2_X1 U1053 ( .A1(n1320), .A2(n1318), .ZN(n1313) );
XNOR2_X1 U1054 ( .A(n1321), .B(n1322), .ZN(n1318) );
XOR2_X1 U1055 ( .A(G143), .B(G131), .Z(n1322) );
NAND3_X1 U1056 ( .A1(n1251), .A2(n1252), .A3(G214), .ZN(n1321) );
INV_X1 U1057 ( .A(G237), .ZN(n1252) );
NOR3_X1 U1058 ( .A1(n1323), .A2(n1324), .A3(n1325), .ZN(n1320) );
AND2_X1 U1059 ( .A1(n1076), .A2(KEYINPUT40), .ZN(n1325) );
NOR3_X1 U1060 ( .A1(KEYINPUT40), .A2(G146), .A3(n1076), .ZN(n1324) );
INV_X1 U1061 ( .A(n1317), .ZN(n1323) );
NAND2_X1 U1062 ( .A1(G146), .A2(n1076), .ZN(n1317) );
XOR2_X1 U1063 ( .A(G125), .B(G140), .Z(n1076) );
XOR2_X1 U1064 ( .A(G104), .B(n1248), .Z(n1091) );
INV_X1 U1065 ( .A(G113), .ZN(n1248) );
INV_X1 U1066 ( .A(n1215), .ZN(n1309) );
XOR2_X1 U1067 ( .A(n1114), .B(n1040), .Z(n1215) );
NAND2_X1 U1068 ( .A1(n1115), .A2(n1106), .ZN(n1040) );
INV_X1 U1069 ( .A(G902), .ZN(n1106) );
XNOR2_X1 U1070 ( .A(n1326), .B(n1327), .ZN(n1115) );
NOR2_X1 U1071 ( .A1(KEYINPUT3), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1072 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1073 ( .A(n1331), .B(n1332), .Z(n1330) );
NOR2_X1 U1074 ( .A1(G122), .A2(KEYINPUT50), .ZN(n1332) );
NAND3_X1 U1075 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1331) );
OR2_X1 U1076 ( .A1(n1308), .A2(KEYINPUT37), .ZN(n1335) );
NAND3_X1 U1077 ( .A1(KEYINPUT37), .A2(n1308), .A3(n1198), .ZN(n1334) );
INV_X1 U1078 ( .A(G134), .ZN(n1198) );
NAND2_X1 U1079 ( .A1(G134), .A2(n1336), .ZN(n1333) );
NAND2_X1 U1080 ( .A1(KEYINPUT37), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1081 ( .A(KEYINPUT14), .B(n1308), .ZN(n1337) );
XOR2_X1 U1082 ( .A(n1202), .B(G143), .Z(n1308) );
INV_X1 U1083 ( .A(G128), .ZN(n1202) );
XOR2_X1 U1084 ( .A(n1012), .B(G116), .Z(n1329) );
INV_X1 U1085 ( .A(G107), .ZN(n1012) );
NAND2_X1 U1086 ( .A1(n1240), .A2(G217), .ZN(n1326) );
AND2_X1 U1087 ( .A1(G234), .A2(n1251), .ZN(n1240) );
XNOR2_X1 U1088 ( .A(n1080), .B(KEYINPUT12), .ZN(n1251) );
INV_X1 U1089 ( .A(G953), .ZN(n1080) );
INV_X1 U1090 ( .A(G478), .ZN(n1114) );
endmodule


