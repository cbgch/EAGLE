//Key = 1100011001001110100111111010111101100100110110010001100001001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334;

XOR2_X1 U742 ( .A(G107), .B(n1020), .Z(G9) );
NOR2_X1 U743 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR4_X1 U744 ( .A1(G953), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1022) );
NOR2_X1 U745 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U746 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR3_X1 U747 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NOR2_X1 U748 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U749 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1033) );
NOR2_X1 U752 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR3_X1 U754 ( .A1(n1036), .A2(n1045), .A3(n1040), .ZN(n1028) );
INV_X1 U755 ( .A(n1046), .ZN(n1040) );
NOR3_X1 U756 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1045) );
NOR3_X1 U757 ( .A1(n1050), .A2(n1032), .A3(n1051), .ZN(n1049) );
INV_X1 U758 ( .A(n1052), .ZN(n1032) );
NOR2_X1 U759 ( .A1(n1053), .A2(n1030), .ZN(n1047) );
NOR2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR3_X1 U761 ( .A1(n1023), .A2(G953), .A3(G952), .ZN(n1021) );
AND4_X1 U762 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1023) );
NOR4_X1 U763 ( .A1(n1060), .A2(n1061), .A3(n1062), .A4(n1063), .ZN(n1059) );
NOR3_X1 U764 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
AND2_X1 U765 ( .A1(n1064), .A2(n1066), .ZN(n1062) );
INV_X1 U766 ( .A(KEYINPUT52), .ZN(n1064) );
XNOR2_X1 U767 ( .A(G478), .B(n1067), .ZN(n1061) );
NAND3_X1 U768 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1060) );
XOR2_X1 U769 ( .A(KEYINPUT22), .B(n1071), .Z(n1069) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
XOR2_X1 U771 ( .A(n1074), .B(n1075), .Z(n1068) );
XNOR2_X1 U772 ( .A(G472), .B(KEYINPUT36), .ZN(n1075) );
NAND2_X1 U773 ( .A1(n1076), .A2(KEYINPUT5), .ZN(n1074) );
XOR2_X1 U774 ( .A(n1077), .B(KEYINPUT58), .Z(n1076) );
AND3_X1 U775 ( .A1(n1050), .A2(n1078), .A3(n1043), .ZN(n1058) );
NAND2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(n1057) );
XNOR2_X1 U777 ( .A(KEYINPUT12), .B(n1073), .ZN(n1080) );
XNOR2_X1 U778 ( .A(n1072), .B(KEYINPUT43), .ZN(n1079) );
XNOR2_X1 U779 ( .A(KEYINPUT37), .B(n1081), .ZN(n1056) );
NAND2_X1 U780 ( .A1(n1082), .A2(n1083), .ZN(G72) );
NAND2_X1 U781 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U782 ( .A1(G953), .A2(n1086), .ZN(n1085) );
NAND2_X1 U783 ( .A1(G900), .A2(G227), .ZN(n1086) );
NAND2_X1 U784 ( .A1(n1087), .A2(n1088), .ZN(n1082) );
NAND2_X1 U785 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U786 ( .A1(G953), .A2(n1091), .ZN(n1090) );
INV_X1 U787 ( .A(n1092), .ZN(n1089) );
INV_X1 U788 ( .A(n1084), .ZN(n1087) );
XNOR2_X1 U789 ( .A(n1093), .B(n1094), .ZN(n1084) );
NOR4_X1 U790 ( .A1(n1095), .A2(n1096), .A3(KEYINPUT56), .A4(n1092), .ZN(n1094) );
NOR2_X1 U791 ( .A1(n1097), .A2(G900), .ZN(n1092) );
NOR2_X1 U792 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
XNOR2_X1 U793 ( .A(n1100), .B(KEYINPUT38), .ZN(n1099) );
INV_X1 U794 ( .A(n1101), .ZN(n1098) );
NOR2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(n1095) );
NAND2_X1 U796 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U797 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U798 ( .A(KEYINPUT34), .B(n1106), .Z(n1102) );
NOR2_X1 U799 ( .A1(n1105), .A2(n1104), .ZN(n1106) );
XOR2_X1 U800 ( .A(n1107), .B(KEYINPUT51), .Z(n1104) );
XNOR2_X1 U801 ( .A(n1108), .B(n1109), .ZN(n1100) );
XOR2_X1 U802 ( .A(KEYINPUT9), .B(KEYINPUT40), .Z(n1109) );
NAND2_X1 U803 ( .A1(n1110), .A2(n1111), .ZN(n1093) );
NAND3_X1 U804 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
XOR2_X1 U805 ( .A(KEYINPUT55), .B(n1115), .Z(n1112) );
XNOR2_X1 U806 ( .A(G953), .B(KEYINPUT2), .ZN(n1110) );
XOR2_X1 U807 ( .A(n1116), .B(n1117), .Z(G69) );
NOR2_X1 U808 ( .A1(n1118), .A2(n1097), .ZN(n1117) );
NOR2_X1 U809 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U810 ( .A1(n1121), .A2(n1122), .ZN(n1116) );
OR3_X1 U811 ( .A1(n1123), .A2(G953), .A3(n1124), .ZN(n1122) );
XOR2_X1 U812 ( .A(n1125), .B(KEYINPUT50), .Z(n1121) );
NAND3_X1 U813 ( .A1(n1124), .A2(n1126), .A3(n1127), .ZN(n1125) );
XOR2_X1 U814 ( .A(KEYINPUT10), .B(n1123), .Z(n1127) );
NAND2_X1 U815 ( .A1(G953), .A2(n1120), .ZN(n1126) );
XNOR2_X1 U816 ( .A(n1128), .B(n1129), .ZN(n1124) );
XOR2_X1 U817 ( .A(KEYINPUT32), .B(KEYINPUT13), .Z(n1129) );
NOR2_X1 U818 ( .A1(n1130), .A2(n1131), .ZN(G66) );
XOR2_X1 U819 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR3_X1 U820 ( .A1(n1134), .A2(KEYINPUT45), .A3(n1066), .ZN(n1133) );
NOR2_X1 U821 ( .A1(n1135), .A2(n1136), .ZN(G63) );
XNOR2_X1 U822 ( .A(n1130), .B(KEYINPUT61), .ZN(n1136) );
XNOR2_X1 U823 ( .A(n1137), .B(n1138), .ZN(n1135) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1134), .ZN(n1138) );
INV_X1 U825 ( .A(G478), .ZN(n1139) );
NOR3_X1 U826 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(G60) );
NOR3_X1 U827 ( .A1(n1143), .A2(G953), .A3(G952), .ZN(n1142) );
INV_X1 U828 ( .A(KEYINPUT15), .ZN(n1143) );
NOR2_X1 U829 ( .A1(KEYINPUT15), .A2(n1144), .ZN(n1141) );
INV_X1 U830 ( .A(n1130), .ZN(n1144) );
XNOR2_X1 U831 ( .A(n1145), .B(n1146), .ZN(n1140) );
NOR3_X1 U832 ( .A1(n1134), .A2(KEYINPUT53), .A3(n1147), .ZN(n1146) );
XOR2_X1 U833 ( .A(G104), .B(n1148), .Z(G6) );
NOR2_X1 U834 ( .A1(n1130), .A2(n1149), .ZN(G57) );
XOR2_X1 U835 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U836 ( .A1(n1152), .A2(n1134), .ZN(n1151) );
NOR2_X1 U837 ( .A1(n1153), .A2(n1154), .ZN(G54) );
XNOR2_X1 U838 ( .A(n1130), .B(KEYINPUT16), .ZN(n1154) );
XOR2_X1 U839 ( .A(n1155), .B(n1156), .Z(n1153) );
NOR2_X1 U840 ( .A1(n1073), .A2(n1134), .ZN(n1156) );
NAND2_X1 U841 ( .A1(n1157), .A2(KEYINPUT23), .ZN(n1155) );
XOR2_X1 U842 ( .A(n1158), .B(n1159), .Z(n1157) );
NAND2_X1 U843 ( .A1(KEYINPUT26), .A2(n1160), .ZN(n1158) );
NOR2_X1 U844 ( .A1(n1130), .A2(n1161), .ZN(G51) );
XNOR2_X1 U845 ( .A(n1162), .B(n1163), .ZN(n1161) );
XOR2_X1 U846 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U847 ( .A1(n1166), .A2(n1134), .ZN(n1165) );
NAND2_X1 U848 ( .A1(G902), .A2(n1025), .ZN(n1134) );
NAND4_X1 U849 ( .A1(n1123), .A2(n1115), .A3(n1114), .A4(n1113), .ZN(n1025) );
NAND4_X1 U850 ( .A1(n1054), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1113) );
NOR2_X1 U851 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XNOR2_X1 U852 ( .A(KEYINPUT25), .B(n1172), .ZN(n1171) );
AND3_X1 U853 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1114) );
NAND4_X1 U854 ( .A1(n1176), .A2(n1037), .A3(n1055), .A4(n1168), .ZN(n1175) );
NOR2_X1 U855 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NOR2_X1 U856 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
INV_X1 U857 ( .A(KEYINPUT46), .ZN(n1180) );
NOR2_X1 U858 ( .A1(n1167), .A2(n1181), .ZN(n1179) );
NOR2_X1 U859 ( .A1(KEYINPUT46), .A2(n1182), .ZN(n1177) );
AND3_X1 U860 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1115) );
NAND2_X1 U861 ( .A1(n1168), .A2(n1186), .ZN(n1185) );
NAND2_X1 U862 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND3_X1 U863 ( .A1(n1189), .A2(n1052), .A3(n1182), .ZN(n1188) );
AND4_X1 U864 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1123) );
NOR4_X1 U865 ( .A1(n1148), .A2(n1020), .A3(n1194), .A4(n1195), .ZN(n1193) );
INV_X1 U866 ( .A(n1196), .ZN(n1195) );
AND2_X1 U867 ( .A1(n1054), .A2(n1197), .ZN(n1020) );
AND2_X1 U868 ( .A1(n1055), .A2(n1197), .ZN(n1148) );
AND4_X1 U869 ( .A1(n1167), .A2(n1042), .A3(n1046), .A4(n1198), .ZN(n1197) );
NOR2_X1 U870 ( .A1(n1199), .A2(n1200), .ZN(n1192) );
NOR2_X1 U871 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NOR3_X1 U872 ( .A1(n1170), .A2(n1203), .A3(n1204), .ZN(n1199) );
NAND4_X1 U873 ( .A1(n1038), .A2(n1048), .A3(n1205), .A4(n1198), .ZN(n1190) );
XNOR2_X1 U874 ( .A(KEYINPUT27), .B(n1201), .ZN(n1205) );
NAND2_X1 U875 ( .A1(KEYINPUT14), .A2(n1128), .ZN(n1164) );
NOR2_X1 U876 ( .A1(n1097), .A2(G952), .ZN(n1130) );
NAND3_X1 U877 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(G48) );
NAND2_X1 U878 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND3_X1 U879 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
NAND2_X1 U880 ( .A1(KEYINPUT6), .A2(KEYINPUT39), .ZN(n1213) );
NAND2_X1 U881 ( .A1(n1214), .A2(n1215), .ZN(n1212) );
INV_X1 U882 ( .A(KEYINPUT8), .ZN(n1215) );
NAND2_X1 U883 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NAND2_X1 U884 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
NAND2_X1 U885 ( .A1(KEYINPUT8), .A2(n1216), .ZN(n1211) );
INV_X1 U886 ( .A(n1183), .ZN(n1209) );
NAND4_X1 U887 ( .A1(n1216), .A2(n1183), .A3(KEYINPUT6), .A4(n1218), .ZN(n1207) );
INV_X1 U888 ( .A(KEYINPUT39), .ZN(n1218) );
NAND2_X1 U889 ( .A1(KEYINPUT39), .A2(n1220), .ZN(n1206) );
NAND2_X1 U890 ( .A1(n1216), .A2(n1221), .ZN(n1220) );
NAND2_X1 U891 ( .A1(n1183), .A2(n1219), .ZN(n1221) );
INV_X1 U892 ( .A(KEYINPUT6), .ZN(n1219) );
NAND2_X1 U893 ( .A1(n1222), .A2(n1055), .ZN(n1183) );
XNOR2_X1 U894 ( .A(G146), .B(KEYINPUT28), .ZN(n1216) );
XNOR2_X1 U895 ( .A(G143), .B(n1184), .ZN(G45) );
NAND4_X1 U896 ( .A1(n1182), .A2(n1037), .A3(n1223), .A4(n1042), .ZN(n1184) );
NOR2_X1 U897 ( .A1(n1081), .A2(n1224), .ZN(n1223) );
XNOR2_X1 U898 ( .A(G140), .B(n1225), .ZN(G42) );
NAND2_X1 U899 ( .A1(n1226), .A2(n1168), .ZN(n1225) );
XOR2_X1 U900 ( .A(n1187), .B(KEYINPUT63), .Z(n1226) );
NAND3_X1 U901 ( .A1(n1038), .A2(n1055), .A3(n1182), .ZN(n1187) );
XNOR2_X1 U902 ( .A(G137), .B(n1227), .ZN(G39) );
NAND4_X1 U903 ( .A1(n1048), .A2(n1189), .A3(n1168), .A4(n1228), .ZN(n1227) );
XNOR2_X1 U904 ( .A(KEYINPUT44), .B(n1172), .ZN(n1228) );
XOR2_X1 U905 ( .A(G134), .B(n1229), .Z(G36) );
NOR2_X1 U906 ( .A1(n1203), .A2(n1230), .ZN(n1229) );
INV_X1 U907 ( .A(n1054), .ZN(n1203) );
XNOR2_X1 U908 ( .A(n1231), .B(n1232), .ZN(G33) );
NOR2_X1 U909 ( .A1(n1233), .A2(n1230), .ZN(n1232) );
NAND3_X1 U910 ( .A1(n1037), .A2(n1168), .A3(n1182), .ZN(n1230) );
INV_X1 U911 ( .A(n1036), .ZN(n1168) );
NAND2_X1 U912 ( .A1(n1070), .A2(n1234), .ZN(n1036) );
INV_X1 U913 ( .A(n1044), .ZN(n1070) );
XNOR2_X1 U914 ( .A(G128), .B(n1173), .ZN(G30) );
NAND2_X1 U915 ( .A1(n1222), .A2(n1054), .ZN(n1173) );
AND3_X1 U916 ( .A1(n1189), .A2(n1042), .A3(n1182), .ZN(n1222) );
AND2_X1 U917 ( .A1(n1167), .A2(n1172), .ZN(n1182) );
XNOR2_X1 U918 ( .A(G101), .B(n1235), .ZN(G3) );
NAND2_X1 U919 ( .A1(n1042), .A2(n1236), .ZN(n1235) );
XNOR2_X1 U920 ( .A(KEYINPUT59), .B(n1202), .ZN(n1236) );
NAND3_X1 U921 ( .A1(n1037), .A2(n1198), .A3(n1048), .ZN(n1202) );
XNOR2_X1 U922 ( .A(G125), .B(n1174), .ZN(G27) );
NAND3_X1 U923 ( .A1(n1038), .A2(n1055), .A3(n1237), .ZN(n1174) );
NOR3_X1 U924 ( .A1(n1030), .A2(n1181), .A3(n1201), .ZN(n1237) );
INV_X1 U925 ( .A(n1172), .ZN(n1181) );
NAND2_X1 U926 ( .A1(n1027), .A2(n1238), .ZN(n1172) );
NAND4_X1 U927 ( .A1(G902), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1238) );
INV_X1 U928 ( .A(G900), .ZN(n1241) );
XNOR2_X1 U929 ( .A(KEYINPUT49), .B(n1097), .ZN(n1239) );
XNOR2_X1 U930 ( .A(G122), .B(n1191), .ZN(G24) );
NAND4_X1 U931 ( .A1(n1242), .A2(n1046), .A3(n1243), .A4(n1244), .ZN(n1191) );
NOR2_X1 U932 ( .A1(n1245), .A2(n1246), .ZN(n1046) );
XOR2_X1 U933 ( .A(n1247), .B(G119), .Z(G21) );
NAND2_X1 U934 ( .A1(KEYINPUT1), .A2(n1196), .ZN(n1247) );
NAND3_X1 U935 ( .A1(n1242), .A2(n1052), .A3(n1189), .ZN(n1196) );
AND2_X1 U936 ( .A1(n1246), .A2(n1245), .ZN(n1189) );
INV_X1 U937 ( .A(n1248), .ZN(n1246) );
INV_X1 U938 ( .A(n1204), .ZN(n1242) );
XNOR2_X1 U939 ( .A(G116), .B(n1249), .ZN(G18) );
NAND4_X1 U940 ( .A1(n1054), .A2(n1198), .A3(n1250), .A4(n1251), .ZN(n1249) );
NOR2_X1 U941 ( .A1(n1170), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U942 ( .A(KEYINPUT21), .B(n1201), .ZN(n1252) );
NOR2_X1 U943 ( .A1(n1244), .A2(n1224), .ZN(n1054) );
INV_X1 U944 ( .A(n1243), .ZN(n1224) );
XOR2_X1 U945 ( .A(G113), .B(n1194), .Z(G15) );
NOR3_X1 U946 ( .A1(n1204), .A2(n1233), .A3(n1170), .ZN(n1194) );
INV_X1 U947 ( .A(n1037), .ZN(n1170) );
NOR2_X1 U948 ( .A1(n1248), .A2(n1245), .ZN(n1037) );
INV_X1 U949 ( .A(n1055), .ZN(n1233) );
NOR2_X1 U950 ( .A1(n1243), .A2(n1081), .ZN(n1055) );
INV_X1 U951 ( .A(n1244), .ZN(n1081) );
NAND3_X1 U952 ( .A1(n1042), .A2(n1198), .A3(n1250), .ZN(n1204) );
INV_X1 U953 ( .A(n1030), .ZN(n1250) );
NAND2_X1 U954 ( .A1(n1253), .A2(n1050), .ZN(n1030) );
INV_X1 U955 ( .A(n1051), .ZN(n1253) );
NAND2_X1 U956 ( .A1(n1254), .A2(n1255), .ZN(G12) );
NAND2_X1 U957 ( .A1(G110), .A2(n1256), .ZN(n1255) );
XOR2_X1 U958 ( .A(n1257), .B(KEYINPUT11), .Z(n1254) );
OR2_X1 U959 ( .A1(n1256), .A2(G110), .ZN(n1257) );
NAND4_X1 U960 ( .A1(n1038), .A2(n1048), .A3(n1042), .A4(n1198), .ZN(n1256) );
NAND2_X1 U961 ( .A1(n1027), .A2(n1258), .ZN(n1198) );
NAND4_X1 U962 ( .A1(G953), .A2(G902), .A3(n1240), .A4(n1120), .ZN(n1258) );
INV_X1 U963 ( .A(G898), .ZN(n1120) );
NAND3_X1 U964 ( .A1(n1240), .A2(n1097), .A3(G952), .ZN(n1027) );
NAND2_X1 U965 ( .A1(G237), .A2(G234), .ZN(n1240) );
INV_X1 U966 ( .A(n1201), .ZN(n1042) );
NAND2_X1 U967 ( .A1(n1234), .A2(n1044), .ZN(n1201) );
XOR2_X1 U968 ( .A(n1259), .B(n1166), .Z(n1044) );
NAND2_X1 U969 ( .A1(G210), .A2(n1260), .ZN(n1166) );
NAND2_X1 U970 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
XOR2_X1 U971 ( .A(n1128), .B(n1263), .Z(n1261) );
XNOR2_X1 U972 ( .A(KEYINPUT19), .B(n1264), .ZN(n1263) );
INV_X1 U973 ( .A(n1162), .ZN(n1264) );
XOR2_X1 U974 ( .A(n1265), .B(n1266), .Z(n1162) );
XNOR2_X1 U975 ( .A(n1267), .B(n1268), .ZN(n1266) );
NOR2_X1 U976 ( .A1(G953), .A2(n1119), .ZN(n1268) );
INV_X1 U977 ( .A(G224), .ZN(n1119) );
INV_X1 U978 ( .A(G125), .ZN(n1267) );
XOR2_X1 U979 ( .A(n1269), .B(n1270), .Z(n1128) );
XOR2_X1 U980 ( .A(n1271), .B(n1272), .Z(n1270) );
XOR2_X1 U981 ( .A(G110), .B(G101), .Z(n1272) );
NOR2_X1 U982 ( .A1(KEYINPUT4), .A2(n1273), .ZN(n1271) );
XNOR2_X1 U983 ( .A(G122), .B(KEYINPUT24), .ZN(n1273) );
XOR2_X1 U984 ( .A(n1274), .B(n1275), .Z(n1269) );
XOR2_X1 U985 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR2_X1 U986 ( .A1(G119), .A2(KEYINPUT35), .ZN(n1276) );
XNOR2_X1 U987 ( .A(n1043), .B(KEYINPUT62), .ZN(n1234) );
NAND2_X1 U988 ( .A1(n1278), .A2(n1260), .ZN(n1043) );
OR2_X1 U989 ( .A1(G902), .A2(G237), .ZN(n1260) );
XOR2_X1 U990 ( .A(KEYINPUT3), .B(G214), .Z(n1278) );
AND2_X1 U991 ( .A1(n1052), .A2(n1167), .ZN(n1048) );
AND2_X1 U992 ( .A1(n1051), .A2(n1050), .ZN(n1167) );
NAND2_X1 U993 ( .A1(G221), .A2(n1279), .ZN(n1050) );
XNOR2_X1 U994 ( .A(n1072), .B(n1073), .ZN(n1051) );
INV_X1 U995 ( .A(G469), .ZN(n1073) );
AND2_X1 U996 ( .A1(n1280), .A2(n1262), .ZN(n1072) );
XNOR2_X1 U997 ( .A(n1160), .B(n1159), .ZN(n1280) );
XNOR2_X1 U998 ( .A(n1281), .B(n1282), .ZN(n1159) );
XOR2_X1 U999 ( .A(G110), .B(n1283), .Z(n1282) );
NOR2_X1 U1000 ( .A1(G953), .A2(n1091), .ZN(n1283) );
INV_X1 U1001 ( .A(G227), .ZN(n1091) );
XOR2_X1 U1002 ( .A(n1107), .B(n1284), .Z(n1281) );
XOR2_X1 U1003 ( .A(n1285), .B(n1286), .Z(n1160) );
XNOR2_X1 U1004 ( .A(n1274), .B(n1105), .ZN(n1286) );
AND2_X1 U1005 ( .A1(n1287), .A2(n1288), .ZN(n1105) );
NAND2_X1 U1006 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
NAND2_X1 U1007 ( .A1(G143), .A2(n1291), .ZN(n1287) );
XOR2_X1 U1008 ( .A(n1289), .B(KEYINPUT20), .Z(n1291) );
XNOR2_X1 U1009 ( .A(G128), .B(G146), .ZN(n1289) );
XNOR2_X1 U1010 ( .A(G104), .B(G107), .ZN(n1274) );
XNOR2_X1 U1011 ( .A(KEYINPUT47), .B(n1292), .ZN(n1285) );
NOR2_X1 U1012 ( .A1(G101), .A2(KEYINPUT17), .ZN(n1292) );
NOR2_X1 U1013 ( .A1(n1243), .A2(n1244), .ZN(n1052) );
XOR2_X1 U1014 ( .A(n1293), .B(n1147), .Z(n1244) );
INV_X1 U1015 ( .A(G475), .ZN(n1147) );
NAND2_X1 U1016 ( .A1(n1145), .A2(n1262), .ZN(n1293) );
XNOR2_X1 U1017 ( .A(n1294), .B(n1295), .ZN(n1145) );
XOR2_X1 U1018 ( .A(n1296), .B(n1297), .Z(n1295) );
XNOR2_X1 U1019 ( .A(n1231), .B(G122), .ZN(n1297) );
INV_X1 U1020 ( .A(G131), .ZN(n1231) );
XNOR2_X1 U1021 ( .A(KEYINPUT31), .B(n1290), .ZN(n1296) );
INV_X1 U1022 ( .A(G143), .ZN(n1290) );
XOR2_X1 U1023 ( .A(n1298), .B(n1299), .Z(n1294) );
XOR2_X1 U1024 ( .A(G113), .B(G104), .Z(n1299) );
XOR2_X1 U1025 ( .A(n1300), .B(n1301), .Z(n1298) );
AND2_X1 U1026 ( .A1(n1302), .A2(G214), .ZN(n1301) );
NAND3_X1 U1027 ( .A1(n1303), .A2(n1304), .A3(KEYINPUT41), .ZN(n1300) );
OR2_X1 U1028 ( .A1(n1305), .A2(KEYINPUT18), .ZN(n1304) );
NAND3_X1 U1029 ( .A1(n1108), .A2(n1306), .A3(KEYINPUT18), .ZN(n1303) );
XOR2_X1 U1030 ( .A(G478), .B(n1307), .Z(n1243) );
NOR2_X1 U1031 ( .A1(KEYINPUT48), .A2(n1067), .ZN(n1307) );
NAND2_X1 U1032 ( .A1(n1137), .A2(n1262), .ZN(n1067) );
XNOR2_X1 U1033 ( .A(n1308), .B(n1309), .ZN(n1137) );
XOR2_X1 U1034 ( .A(n1310), .B(n1311), .Z(n1309) );
NOR2_X1 U1035 ( .A1(G116), .A2(KEYINPUT42), .ZN(n1311) );
AND3_X1 U1036 ( .A1(G234), .A2(n1097), .A3(G217), .ZN(n1310) );
XOR2_X1 U1037 ( .A(n1312), .B(n1313), .Z(n1308) );
NOR2_X1 U1038 ( .A1(KEYINPUT54), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1039 ( .A(G134), .B(n1315), .Z(n1314) );
XNOR2_X1 U1040 ( .A(G107), .B(G122), .ZN(n1312) );
AND2_X1 U1041 ( .A1(n1248), .A2(n1245), .ZN(n1038) );
NAND2_X1 U1042 ( .A1(n1316), .A2(n1078), .ZN(n1245) );
NAND2_X1 U1043 ( .A1(n1065), .A2(n1066), .ZN(n1078) );
OR2_X1 U1044 ( .A1(n1066), .A2(n1065), .ZN(n1316) );
NOR2_X1 U1045 ( .A1(n1132), .A2(G902), .ZN(n1065) );
XOR2_X1 U1046 ( .A(n1317), .B(n1318), .Z(n1132) );
XOR2_X1 U1047 ( .A(n1305), .B(n1319), .Z(n1318) );
XNOR2_X1 U1048 ( .A(n1320), .B(n1321), .ZN(n1319) );
NAND2_X1 U1049 ( .A1(KEYINPUT29), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U1050 ( .A(n1323), .B(G119), .ZN(n1322) );
NAND2_X1 U1051 ( .A1(KEYINPUT0), .A2(n1324), .ZN(n1320) );
XOR2_X1 U1052 ( .A(G137), .B(n1325), .Z(n1324) );
AND3_X1 U1053 ( .A1(G221), .A2(n1097), .A3(G234), .ZN(n1325) );
INV_X1 U1054 ( .A(G953), .ZN(n1097) );
XNOR2_X1 U1055 ( .A(n1108), .B(n1306), .ZN(n1305) );
INV_X1 U1056 ( .A(G146), .ZN(n1306) );
XNOR2_X1 U1057 ( .A(G125), .B(n1284), .ZN(n1108) );
XOR2_X1 U1058 ( .A(G140), .B(KEYINPUT7), .Z(n1284) );
XOR2_X1 U1059 ( .A(n1326), .B(G110), .Z(n1317) );
XNOR2_X1 U1060 ( .A(KEYINPUT60), .B(KEYINPUT30), .ZN(n1326) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1279), .ZN(n1066) );
NAND2_X1 U1062 ( .A1(G234), .A2(n1262), .ZN(n1279) );
XOR2_X1 U1063 ( .A(n1327), .B(n1077), .Z(n1248) );
NAND2_X1 U1064 ( .A1(n1328), .A2(n1262), .ZN(n1077) );
INV_X1 U1065 ( .A(G902), .ZN(n1262) );
XOR2_X1 U1066 ( .A(n1150), .B(KEYINPUT33), .Z(n1328) );
XOR2_X1 U1067 ( .A(n1329), .B(n1330), .Z(n1150) );
XOR2_X1 U1068 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1069 ( .A(G101), .B(G119), .ZN(n1332) );
NAND2_X1 U1070 ( .A1(G210), .A2(n1302), .ZN(n1331) );
NOR2_X1 U1071 ( .A1(G953), .A2(G237), .ZN(n1302) );
XOR2_X1 U1072 ( .A(n1333), .B(n1265), .Z(n1329) );
XOR2_X1 U1073 ( .A(G146), .B(n1315), .Z(n1265) );
XNOR2_X1 U1074 ( .A(n1323), .B(G143), .ZN(n1315) );
INV_X1 U1075 ( .A(G128), .ZN(n1323) );
XOR2_X1 U1076 ( .A(n1107), .B(n1277), .Z(n1333) );
XOR2_X1 U1077 ( .A(G113), .B(G116), .Z(n1277) );
XNOR2_X1 U1078 ( .A(G131), .B(n1334), .ZN(n1107) );
XOR2_X1 U1079 ( .A(G137), .B(G134), .Z(n1334) );
NAND2_X1 U1080 ( .A1(KEYINPUT57), .A2(n1152), .ZN(n1327) );
INV_X1 U1081 ( .A(G472), .ZN(n1152) );
endmodule


