//Key = 1100111010100111010111000110101101001010101010000100101101111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348;

XNOR2_X1 U747 ( .A(G107), .B(n1033), .ZN(G9) );
NAND3_X1 U748 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(G75) );
NAND2_X1 U749 ( .A1(G952), .A2(n1037), .ZN(n1035) );
NAND4_X1 U750 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1037) );
NAND2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(n1039) );
NAND2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NAND2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1049) );
OR2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND3_X1 U759 ( .A1(n1051), .A2(n1059), .A3(n1055), .ZN(n1044) );
NAND3_X1 U760 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NAND2_X1 U761 ( .A1(n1048), .A2(n1063), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U763 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U764 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1060) );
XOR2_X1 U765 ( .A(KEYINPUT50), .B(n1046), .Z(n1069) );
INV_X1 U766 ( .A(n1071), .ZN(n1042) );
NAND2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1034) );
XOR2_X1 U768 ( .A(n1040), .B(KEYINPUT6), .Z(n1072) );
NAND4_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1040) );
NOR4_X1 U770 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
NOR2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
INV_X1 U772 ( .A(KEYINPUT54), .ZN(n1083) );
NOR2_X1 U773 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
AND2_X1 U774 ( .A1(n1086), .A2(KEYINPUT41), .ZN(n1085) );
NOR3_X1 U775 ( .A1(KEYINPUT41), .A2(G472), .A3(n1086), .ZN(n1084) );
NOR2_X1 U776 ( .A1(KEYINPUT54), .A2(n1087), .ZN(n1080) );
NOR2_X1 U777 ( .A1(G472), .A2(n1088), .ZN(n1087) );
XOR2_X1 U778 ( .A(n1086), .B(KEYINPUT41), .Z(n1088) );
XOR2_X1 U779 ( .A(KEYINPUT3), .B(n1089), .Z(n1079) );
NAND3_X1 U780 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1078) );
XOR2_X1 U781 ( .A(n1093), .B(n1094), .Z(n1092) );
XOR2_X1 U782 ( .A(KEYINPUT53), .B(n1095), .Z(n1094) );
NAND2_X1 U783 ( .A1(KEYINPUT28), .A2(G475), .ZN(n1093) );
XNOR2_X1 U784 ( .A(n1096), .B(n1097), .ZN(n1091) );
NOR2_X1 U785 ( .A1(G469), .A2(KEYINPUT16), .ZN(n1097) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(n1090) );
XOR2_X1 U787 ( .A(KEYINPUT43), .B(G478), .Z(n1099) );
NOR3_X1 U788 ( .A1(n1100), .A2(n1070), .A3(n1066), .ZN(n1076) );
NAND2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1075) );
XOR2_X1 U790 ( .A(KEYINPUT35), .B(n1103), .Z(n1101) );
NAND2_X1 U791 ( .A1(G472), .A2(n1086), .ZN(n1074) );
XOR2_X1 U792 ( .A(n1104), .B(n1105), .Z(G72) );
NOR2_X1 U793 ( .A1(n1106), .A2(n1041), .ZN(n1105) );
AND2_X1 U794 ( .A1(G227), .A2(G900), .ZN(n1106) );
NAND2_X1 U795 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
NAND2_X1 U796 ( .A1(n1109), .A2(n1041), .ZN(n1108) );
XNOR2_X1 U797 ( .A(n1110), .B(n1111), .ZN(n1109) );
NAND3_X1 U798 ( .A1(G900), .A2(n1110), .A3(G953), .ZN(n1107) );
XNOR2_X1 U799 ( .A(n1112), .B(n1113), .ZN(n1110) );
NAND2_X1 U800 ( .A1(KEYINPUT20), .A2(n1114), .ZN(n1112) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U802 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U803 ( .A1(KEYINPUT52), .A2(n1119), .ZN(n1117) );
XOR2_X1 U804 ( .A(n1120), .B(n1121), .Z(G69) );
XOR2_X1 U805 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U806 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U808 ( .A1(KEYINPUT33), .A2(n1128), .ZN(n1127) );
XOR2_X1 U809 ( .A(n1129), .B(KEYINPUT42), .Z(n1124) );
NAND2_X1 U810 ( .A1(G953), .A2(n1130), .ZN(n1129) );
NOR2_X1 U811 ( .A1(n1131), .A2(G953), .ZN(n1122) );
NOR3_X1 U812 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
INV_X1 U813 ( .A(n1135), .ZN(n1133) );
XOR2_X1 U814 ( .A(KEYINPUT25), .B(n1136), .Z(n1132) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1041), .ZN(n1120) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1130), .ZN(n1137) );
NOR2_X1 U817 ( .A1(n1139), .A2(n1140), .ZN(G66) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U819 ( .A(n1143), .B(KEYINPUT1), .Z(n1142) );
NAND2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
AND4_X1 U822 ( .A1(n1146), .A2(G217), .A3(n1147), .A4(n1148), .ZN(n1144) );
XOR2_X1 U823 ( .A(n1149), .B(KEYINPUT55), .Z(n1146) );
NOR2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(G63) );
XOR2_X1 U825 ( .A(n1036), .B(KEYINPUT49), .Z(n1151) );
NOR3_X1 U826 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1150) );
NOR3_X1 U827 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1154) );
NOR2_X1 U828 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
NOR2_X1 U829 ( .A1(n1038), .A2(n1156), .ZN(n1158) );
INV_X1 U830 ( .A(n1148), .ZN(n1038) );
NOR2_X1 U831 ( .A1(n1139), .A2(n1160), .ZN(G60) );
XOR2_X1 U832 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND3_X1 U833 ( .A1(G475), .A2(n1148), .A3(n1163), .ZN(n1161) );
XOR2_X1 U834 ( .A(n1149), .B(KEYINPUT8), .Z(n1163) );
XNOR2_X1 U835 ( .A(G104), .B(n1164), .ZN(G6) );
NOR2_X1 U836 ( .A1(n1139), .A2(n1165), .ZN(G57) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U838 ( .A(n1168), .B(KEYINPUT60), .Z(n1167) );
NAND2_X1 U839 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
XNOR2_X1 U841 ( .A(n1171), .B(n1172), .ZN(n1170) );
NAND2_X1 U842 ( .A1(KEYINPUT5), .A2(G101), .ZN(n1171) );
XOR2_X1 U843 ( .A(n1173), .B(n1174), .Z(n1169) );
XNOR2_X1 U844 ( .A(n1175), .B(n1176), .ZN(n1174) );
NOR2_X1 U845 ( .A1(KEYINPUT23), .A2(n1177), .ZN(n1176) );
NAND2_X1 U846 ( .A1(KEYINPUT63), .A2(n1178), .ZN(n1175) );
NAND3_X1 U847 ( .A1(n1179), .A2(n1148), .A3(G472), .ZN(n1178) );
XOR2_X1 U848 ( .A(KEYINPUT11), .B(G902), .Z(n1179) );
NOR2_X1 U849 ( .A1(n1139), .A2(n1180), .ZN(G54) );
XOR2_X1 U850 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U851 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U852 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U853 ( .A(KEYINPUT47), .B(G140), .Z(n1183) );
XOR2_X1 U854 ( .A(n1187), .B(n1188), .Z(n1181) );
XOR2_X1 U855 ( .A(n1189), .B(n1190), .Z(n1187) );
NOR2_X1 U856 ( .A1(n1191), .A2(n1157), .ZN(n1190) );
INV_X1 U857 ( .A(G469), .ZN(n1191) );
NAND2_X1 U858 ( .A1(KEYINPUT31), .A2(n1192), .ZN(n1189) );
NOR3_X1 U859 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(G51) );
AND2_X1 U860 ( .A1(KEYINPUT21), .A2(n1139), .ZN(n1195) );
INV_X1 U861 ( .A(n1036), .ZN(n1139) );
NAND2_X1 U862 ( .A1(G953), .A2(n1073), .ZN(n1036) );
INV_X1 U863 ( .A(G952), .ZN(n1073) );
NOR3_X1 U864 ( .A1(KEYINPUT21), .A2(G953), .A3(G952), .ZN(n1194) );
NOR2_X1 U865 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
XOR2_X1 U866 ( .A(n1198), .B(KEYINPUT40), .Z(n1197) );
NAND2_X1 U867 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
OR2_X1 U868 ( .A1(n1157), .A2(n1201), .ZN(n1200) );
NOR3_X1 U869 ( .A1(n1199), .A2(n1201), .A3(n1157), .ZN(n1196) );
NAND2_X1 U870 ( .A1(G902), .A2(n1148), .ZN(n1157) );
NAND4_X1 U871 ( .A1(n1202), .A2(n1111), .A3(n1136), .A4(n1135), .ZN(n1148) );
AND4_X1 U872 ( .A1(n1164), .A2(n1203), .A3(n1204), .A4(n1033), .ZN(n1136) );
NAND3_X1 U873 ( .A1(n1051), .A2(n1205), .A3(n1206), .ZN(n1033) );
NAND3_X1 U874 ( .A1(n1206), .A2(n1051), .A3(n1207), .ZN(n1164) );
AND4_X1 U875 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1111) );
NOR4_X1 U876 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
INV_X1 U877 ( .A(n1216), .ZN(n1215) );
NAND2_X1 U878 ( .A1(n1217), .A2(n1218), .ZN(n1210) );
NAND2_X1 U879 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND4_X1 U880 ( .A1(n1221), .A2(n1205), .A3(n1222), .A4(n1223), .ZN(n1220) );
OR2_X1 U881 ( .A1(n1224), .A2(KEYINPUT56), .ZN(n1223) );
NAND2_X1 U882 ( .A1(KEYINPUT56), .A2(n1225), .ZN(n1222) );
NAND2_X1 U883 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XNOR2_X1 U884 ( .A(KEYINPUT19), .B(n1228), .ZN(n1219) );
NAND2_X1 U885 ( .A1(n1229), .A2(n1058), .ZN(n1208) );
INV_X1 U886 ( .A(n1134), .ZN(n1202) );
NAND3_X1 U887 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1134) );
XOR2_X1 U888 ( .A(n1233), .B(n1234), .Z(n1199) );
XOR2_X1 U889 ( .A(n1235), .B(n1236), .Z(n1234) );
NAND2_X1 U890 ( .A1(KEYINPUT44), .A2(n1237), .ZN(n1235) );
XOR2_X1 U891 ( .A(G146), .B(n1238), .Z(G48) );
NOR3_X1 U892 ( .A1(n1228), .A2(KEYINPUT2), .A3(n1239), .ZN(n1238) );
NAND3_X1 U893 ( .A1(n1221), .A2(n1207), .A3(n1224), .ZN(n1228) );
XOR2_X1 U894 ( .A(n1240), .B(n1209), .Z(G45) );
NAND4_X1 U895 ( .A1(n1217), .A2(n1057), .A3(n1241), .A4(n1242), .ZN(n1209) );
AND2_X1 U896 ( .A1(n1224), .A2(n1243), .ZN(n1242) );
XOR2_X1 U897 ( .A(n1244), .B(n1245), .Z(G42) );
NAND4_X1 U898 ( .A1(n1246), .A2(n1224), .A3(n1058), .A4(n1207), .ZN(n1245) );
XNOR2_X1 U899 ( .A(n1048), .B(KEYINPUT0), .ZN(n1246) );
NAND2_X1 U900 ( .A1(n1247), .A2(n1248), .ZN(G39) );
NAND2_X1 U901 ( .A1(n1214), .A2(n1249), .ZN(n1248) );
XOR2_X1 U902 ( .A(KEYINPUT14), .B(n1250), .Z(n1247) );
NOR2_X1 U903 ( .A1(n1214), .A2(n1249), .ZN(n1250) );
INV_X1 U904 ( .A(G137), .ZN(n1249) );
AND4_X1 U905 ( .A1(n1224), .A2(n1048), .A3(n1055), .A4(n1221), .ZN(n1214) );
XOR2_X1 U906 ( .A(G134), .B(n1251), .Z(G36) );
NOR2_X1 U907 ( .A1(KEYINPUT37), .A2(n1216), .ZN(n1251) );
NAND4_X1 U908 ( .A1(n1224), .A2(n1048), .A3(n1205), .A4(n1057), .ZN(n1216) );
XOR2_X1 U909 ( .A(n1252), .B(n1253), .Z(G33) );
NAND2_X1 U910 ( .A1(KEYINPUT17), .A2(n1213), .ZN(n1253) );
AND2_X1 U911 ( .A1(n1229), .A2(n1057), .ZN(n1213) );
AND3_X1 U912 ( .A1(n1048), .A2(n1207), .A3(n1224), .ZN(n1229) );
NOR2_X1 U913 ( .A1(n1089), .A2(n1070), .ZN(n1048) );
INV_X1 U914 ( .A(n1068), .ZN(n1089) );
XNOR2_X1 U915 ( .A(G128), .B(n1254), .ZN(G30) );
NAND4_X1 U916 ( .A1(n1255), .A2(n1224), .A3(n1256), .A4(n1221), .ZN(n1254) );
NOR2_X1 U917 ( .A1(KEYINPUT48), .A2(n1239), .ZN(n1256) );
NOR2_X1 U918 ( .A1(n1064), .A2(n1226), .ZN(n1224) );
INV_X1 U919 ( .A(n1227), .ZN(n1064) );
XOR2_X1 U920 ( .A(n1054), .B(KEYINPUT61), .Z(n1255) );
XNOR2_X1 U921 ( .A(G101), .B(n1203), .ZN(G3) );
NAND3_X1 U922 ( .A1(n1206), .A2(n1057), .A3(n1055), .ZN(n1203) );
XOR2_X1 U923 ( .A(G125), .B(n1212), .Z(G27) );
NOR4_X1 U924 ( .A1(n1257), .A2(n1061), .A3(n1053), .A4(n1226), .ZN(n1212) );
AND2_X1 U925 ( .A1(n1071), .A2(n1258), .ZN(n1226) );
NAND4_X1 U926 ( .A1(G953), .A2(G902), .A3(n1259), .A4(n1260), .ZN(n1258) );
INV_X1 U927 ( .A(G900), .ZN(n1260) );
INV_X1 U928 ( .A(n1207), .ZN(n1053) );
INV_X1 U929 ( .A(n1058), .ZN(n1257) );
XNOR2_X1 U930 ( .A(G122), .B(n1232), .ZN(G24) );
NAND4_X1 U931 ( .A1(n1243), .A2(n1261), .A3(n1241), .A4(n1051), .ZN(n1232) );
XNOR2_X1 U932 ( .A(G119), .B(n1230), .ZN(G21) );
NAND3_X1 U933 ( .A1(n1261), .A2(n1221), .A3(n1055), .ZN(n1230) );
NOR2_X1 U934 ( .A1(n1262), .A2(n1263), .ZN(n1221) );
XOR2_X1 U935 ( .A(n1264), .B(G116), .Z(G18) );
NAND2_X1 U936 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
OR2_X1 U937 ( .A1(n1135), .A2(KEYINPUT18), .ZN(n1266) );
NAND3_X1 U938 ( .A1(n1205), .A2(n1057), .A3(n1261), .ZN(n1135) );
INV_X1 U939 ( .A(n1054), .ZN(n1205) );
NAND4_X1 U940 ( .A1(n1057), .A2(n1054), .A3(n1261), .A4(KEYINPUT18), .ZN(n1265) );
NOR2_X1 U941 ( .A1(n1061), .A2(n1267), .ZN(n1261) );
INV_X1 U942 ( .A(n1268), .ZN(n1267) );
NAND2_X1 U943 ( .A1(n1046), .A2(n1217), .ZN(n1061) );
INV_X1 U944 ( .A(n1239), .ZN(n1217) );
XNOR2_X1 U945 ( .A(n1269), .B(KEYINPUT62), .ZN(n1239) );
NAND2_X1 U946 ( .A1(n1241), .A2(n1270), .ZN(n1054) );
XNOR2_X1 U947 ( .A(G113), .B(n1231), .ZN(G15) );
NAND4_X1 U948 ( .A1(n1057), .A2(n1268), .A3(n1269), .A4(n1271), .ZN(n1231) );
AND2_X1 U949 ( .A1(n1207), .A2(n1046), .ZN(n1271) );
NOR2_X1 U950 ( .A1(n1272), .A2(n1066), .ZN(n1046) );
INV_X1 U951 ( .A(n1067), .ZN(n1272) );
NOR2_X1 U952 ( .A1(n1270), .A2(n1241), .ZN(n1207) );
INV_X1 U953 ( .A(n1243), .ZN(n1270) );
NAND2_X1 U954 ( .A1(n1273), .A2(n1274), .ZN(n1057) );
NAND2_X1 U955 ( .A1(n1051), .A2(n1275), .ZN(n1274) );
INV_X1 U956 ( .A(KEYINPUT38), .ZN(n1275) );
AND2_X1 U957 ( .A1(n1263), .A2(n1262), .ZN(n1051) );
NAND3_X1 U958 ( .A1(n1263), .A2(n1276), .A3(KEYINPUT38), .ZN(n1273) );
XOR2_X1 U959 ( .A(n1185), .B(n1204), .Z(G12) );
NAND3_X1 U960 ( .A1(n1055), .A2(n1206), .A3(n1058), .ZN(n1204) );
NOR2_X1 U961 ( .A1(n1276), .A2(n1263), .ZN(n1058) );
NOR2_X1 U962 ( .A1(n1277), .A2(n1100), .ZN(n1263) );
NOR2_X1 U963 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
AND2_X1 U964 ( .A1(n1103), .A2(n1102), .ZN(n1277) );
OR2_X1 U965 ( .A1(n1145), .A2(G902), .ZN(n1102) );
XNOR2_X1 U966 ( .A(n1278), .B(n1279), .ZN(n1145) );
XOR2_X1 U967 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U968 ( .A(n1282), .B(n1283), .ZN(n1281) );
NOR2_X1 U969 ( .A1(KEYINPUT45), .A2(n1284), .ZN(n1283) );
XOR2_X1 U970 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U971 ( .A(KEYINPUT10), .B(G137), .Z(n1286) );
AND3_X1 U972 ( .A1(G221), .A2(n1041), .A3(G234), .ZN(n1285) );
NAND2_X1 U973 ( .A1(KEYINPUT4), .A2(n1244), .ZN(n1282) );
INV_X1 U974 ( .A(G140), .ZN(n1244) );
XOR2_X1 U975 ( .A(n1185), .B(n1287), .Z(n1278) );
XOR2_X1 U976 ( .A(G125), .B(G119), .Z(n1287) );
AND2_X1 U977 ( .A1(n1288), .A2(n1147), .ZN(n1103) );
XOR2_X1 U978 ( .A(KEYINPUT27), .B(G217), .Z(n1288) );
INV_X1 U979 ( .A(n1262), .ZN(n1276) );
XOR2_X1 U980 ( .A(n1086), .B(G472), .Z(n1262) );
NAND2_X1 U981 ( .A1(n1289), .A2(n1149), .ZN(n1086) );
XOR2_X1 U982 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U983 ( .A(n1172), .B(n1292), .Z(n1291) );
NOR2_X1 U984 ( .A1(G101), .A2(KEYINPUT12), .ZN(n1292) );
AND3_X1 U985 ( .A1(n1293), .A2(n1041), .A3(G210), .ZN(n1172) );
XOR2_X1 U986 ( .A(n1173), .B(n1177), .Z(n1290) );
INV_X1 U987 ( .A(n1294), .ZN(n1177) );
XNOR2_X1 U988 ( .A(n1192), .B(n1295), .ZN(n1173) );
AND3_X1 U989 ( .A1(n1269), .A2(n1268), .A3(n1227), .ZN(n1206) );
NOR2_X1 U990 ( .A1(n1067), .A2(n1066), .ZN(n1227) );
AND2_X1 U991 ( .A1(G221), .A2(n1147), .ZN(n1066) );
NAND2_X1 U992 ( .A1(G234), .A2(n1149), .ZN(n1147) );
XOR2_X1 U993 ( .A(n1096), .B(G469), .Z(n1067) );
NAND2_X1 U994 ( .A1(n1296), .A2(n1149), .ZN(n1096) );
XNOR2_X1 U995 ( .A(n1188), .B(n1297), .ZN(n1296) );
XNOR2_X1 U996 ( .A(n1298), .B(n1192), .ZN(n1297) );
XNOR2_X1 U997 ( .A(n1118), .B(n1299), .ZN(n1192) );
XOR2_X1 U998 ( .A(KEYINPUT32), .B(n1119), .Z(n1299) );
XOR2_X1 U999 ( .A(n1252), .B(G137), .Z(n1118) );
INV_X1 U1000 ( .A(G131), .ZN(n1252) );
NAND2_X1 U1001 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
NAND2_X1 U1002 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
XNOR2_X1 U1003 ( .A(KEYINPUT36), .B(n1186), .ZN(n1302) );
XOR2_X1 U1004 ( .A(KEYINPUT26), .B(n1304), .Z(n1300) );
NOR2_X1 U1005 ( .A1(n1186), .A2(n1303), .ZN(n1304) );
XOR2_X1 U1006 ( .A(n1185), .B(n1305), .Z(n1303) );
NAND2_X1 U1007 ( .A1(KEYINPUT58), .A2(G140), .ZN(n1305) );
NAND2_X1 U1008 ( .A1(G227), .A2(n1041), .ZN(n1186) );
XNOR2_X1 U1009 ( .A(n1306), .B(n1307), .ZN(n1188) );
XOR2_X1 U1010 ( .A(n1308), .B(n1115), .Z(n1307) );
XNOR2_X1 U1011 ( .A(n1309), .B(n1310), .ZN(n1115) );
NOR2_X1 U1012 ( .A1(G146), .A2(KEYINPUT9), .ZN(n1310) );
NOR2_X1 U1013 ( .A1(G107), .A2(KEYINPUT22), .ZN(n1308) );
XNOR2_X1 U1014 ( .A(G101), .B(G104), .ZN(n1306) );
NAND2_X1 U1015 ( .A1(n1071), .A2(n1311), .ZN(n1268) );
NAND4_X1 U1016 ( .A1(G953), .A2(G902), .A3(n1259), .A4(n1130), .ZN(n1311) );
INV_X1 U1017 ( .A(G898), .ZN(n1130) );
NAND3_X1 U1018 ( .A1(n1259), .A2(n1041), .A3(G952), .ZN(n1071) );
NAND2_X1 U1019 ( .A1(G237), .A2(G234), .ZN(n1259) );
NOR2_X1 U1020 ( .A1(n1068), .A2(n1070), .ZN(n1269) );
AND2_X1 U1021 ( .A1(G214), .A2(n1312), .ZN(n1070) );
XNOR2_X1 U1022 ( .A(n1313), .B(n1201), .ZN(n1068) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1312), .ZN(n1201) );
NAND2_X1 U1024 ( .A1(n1149), .A2(n1293), .ZN(n1312) );
NAND2_X1 U1025 ( .A1(n1314), .A2(n1149), .ZN(n1313) );
XOR2_X1 U1026 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1027 ( .A(n1317), .B(n1236), .Z(n1316) );
XOR2_X1 U1028 ( .A(n1295), .B(n1318), .Z(n1236) );
INV_X1 U1029 ( .A(G125), .ZN(n1318) );
XNOR2_X1 U1030 ( .A(n1240), .B(n1280), .ZN(n1295) );
XOR2_X1 U1031 ( .A(G128), .B(G146), .Z(n1280) );
NAND2_X1 U1032 ( .A1(KEYINPUT57), .A2(n1233), .ZN(n1317) );
XNOR2_X1 U1033 ( .A(n1128), .B(n1126), .ZN(n1233) );
NAND3_X1 U1034 ( .A1(n1319), .A2(n1320), .A3(n1321), .ZN(n1126) );
NAND2_X1 U1035 ( .A1(KEYINPUT7), .A2(G122), .ZN(n1321) );
OR3_X1 U1036 ( .A1(G122), .A2(KEYINPUT7), .A3(n1185), .ZN(n1320) );
NAND2_X1 U1037 ( .A1(n1322), .A2(n1185), .ZN(n1319) );
NAND2_X1 U1038 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
INV_X1 U1039 ( .A(KEYINPUT7), .ZN(n1324) );
XOR2_X1 U1040 ( .A(KEYINPUT30), .B(G122), .Z(n1323) );
XNOR2_X1 U1041 ( .A(n1325), .B(n1326), .ZN(n1128) );
XOR2_X1 U1042 ( .A(G107), .B(G101), .Z(n1326) );
XOR2_X1 U1043 ( .A(n1294), .B(n1327), .Z(n1325) );
NOR2_X1 U1044 ( .A1(G104), .A2(KEYINPUT51), .ZN(n1327) );
XNOR2_X1 U1045 ( .A(G113), .B(n1328), .ZN(n1294) );
XOR2_X1 U1046 ( .A(G119), .B(G116), .Z(n1328) );
XOR2_X1 U1047 ( .A(KEYINPUT39), .B(n1237), .Z(n1315) );
NOR2_X1 U1048 ( .A1(n1138), .A2(G953), .ZN(n1237) );
INV_X1 U1049 ( .A(G224), .ZN(n1138) );
NOR2_X1 U1050 ( .A1(n1243), .A2(n1241), .ZN(n1055) );
XOR2_X1 U1051 ( .A(n1329), .B(n1152), .Z(n1241) );
INV_X1 U1052 ( .A(n1098), .ZN(n1152) );
NAND2_X1 U1053 ( .A1(n1155), .A2(n1149), .ZN(n1098) );
INV_X1 U1054 ( .A(n1159), .ZN(n1155) );
XOR2_X1 U1055 ( .A(n1330), .B(n1331), .Z(n1159) );
XOR2_X1 U1056 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U1057 ( .A(G122), .B(n1334), .Z(n1333) );
AND3_X1 U1058 ( .A1(G217), .A2(n1041), .A3(G234), .ZN(n1334) );
NOR2_X1 U1059 ( .A1(KEYINPUT46), .A2(n1335), .ZN(n1332) );
INV_X1 U1060 ( .A(G116), .ZN(n1335) );
XOR2_X1 U1061 ( .A(n1336), .B(n1119), .Z(n1330) );
XOR2_X1 U1062 ( .A(G134), .B(KEYINPUT34), .Z(n1119) );
XNOR2_X1 U1063 ( .A(n1337), .B(n1309), .ZN(n1336) );
XOR2_X1 U1064 ( .A(G128), .B(n1240), .Z(n1309) );
INV_X1 U1065 ( .A(G143), .ZN(n1240) );
NAND2_X1 U1066 ( .A1(KEYINPUT59), .A2(G107), .ZN(n1337) );
NAND2_X1 U1067 ( .A1(KEYINPUT15), .A2(n1156), .ZN(n1329) );
INV_X1 U1068 ( .A(G478), .ZN(n1156) );
XOR2_X1 U1069 ( .A(n1338), .B(n1095), .Z(n1243) );
AND2_X1 U1070 ( .A1(n1162), .A2(n1149), .ZN(n1095) );
INV_X1 U1071 ( .A(G902), .ZN(n1149) );
XNOR2_X1 U1072 ( .A(n1339), .B(n1340), .ZN(n1162) );
XOR2_X1 U1073 ( .A(n1113), .B(n1341), .Z(n1340) );
XOR2_X1 U1074 ( .A(G104), .B(n1342), .Z(n1341) );
NOR2_X1 U1075 ( .A1(KEYINPUT29), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1076 ( .A(G131), .B(n1344), .Z(n1343) );
NOR2_X1 U1077 ( .A1(KEYINPUT24), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1078 ( .A(G143), .B(n1346), .Z(n1345) );
AND3_X1 U1079 ( .A1(G214), .A2(n1041), .A3(n1293), .ZN(n1346) );
INV_X1 U1080 ( .A(G237), .ZN(n1293) );
INV_X1 U1081 ( .A(G953), .ZN(n1041) );
XOR2_X1 U1082 ( .A(G125), .B(G140), .Z(n1113) );
XNOR2_X1 U1083 ( .A(G113), .B(n1347), .ZN(n1339) );
XOR2_X1 U1084 ( .A(G146), .B(G122), .Z(n1347) );
NAND2_X1 U1085 ( .A1(KEYINPUT13), .A2(n1348), .ZN(n1338) );
INV_X1 U1086 ( .A(G475), .ZN(n1348) );
INV_X1 U1087 ( .A(G110), .ZN(n1185) );
endmodule


