//Key = 0111110001100111100111001101010001001111111101011101100101010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412;

XNOR2_X1 U784 ( .A(n1077), .B(n1078), .ZN(G9) );
NOR2_X1 U785 ( .A1(n1079), .A2(n1080), .ZN(G75) );
NOR2_X1 U786 ( .A1(G952), .A2(n1081), .ZN(n1080) );
NOR3_X1 U787 ( .A1(n1082), .A2(n1083), .A3(n1081), .ZN(n1079) );
NAND2_X1 U788 ( .A1(n1084), .A2(n1085), .ZN(n1081) );
NAND4_X1 U789 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1085) );
NOR4_X1 U790 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
NOR3_X1 U791 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
NOR2_X1 U792 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
AND3_X1 U793 ( .A1(n1098), .A2(n1097), .A3(KEYINPUT39), .ZN(n1095) );
NOR2_X1 U794 ( .A1(n1099), .A2(KEYINPUT0), .ZN(n1097) );
NOR2_X1 U795 ( .A1(KEYINPUT39), .A2(n1100), .ZN(n1094) );
NOR2_X1 U796 ( .A1(n1101), .A2(n1102), .ZN(n1091) );
XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n1103), .ZN(n1102) );
INV_X1 U798 ( .A(n1104), .ZN(n1101) );
NOR2_X1 U799 ( .A1(n1105), .A2(n1106), .ZN(n1088) );
NOR2_X1 U800 ( .A1(n1107), .A2(n1108), .ZN(n1083) );
NOR2_X1 U801 ( .A1(n1109), .A2(n1110), .ZN(n1107) );
NOR3_X1 U802 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1110) );
NOR2_X1 U803 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR2_X1 U804 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U805 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NOR2_X1 U806 ( .A1(n1120), .A2(n1105), .ZN(n1118) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1114) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NOR3_X1 U809 ( .A1(n1117), .A2(n1125), .A3(n1122), .ZN(n1109) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1128), .A2(n1111), .ZN(n1127) );
NOR3_X1 U812 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
NOR2_X1 U813 ( .A1(KEYINPUT20), .A2(n1113), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1132), .A2(n1113), .ZN(n1126) );
NOR2_X1 U815 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR3_X1 U816 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1133) );
INV_X1 U817 ( .A(KEYINPUT20), .ZN(n1135) );
INV_X1 U818 ( .A(n1138), .ZN(n1117) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(G72) );
NOR2_X1 U820 ( .A1(n1141), .A2(n1084), .ZN(n1140) );
NOR2_X1 U821 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U822 ( .A1(n1144), .A2(n1145), .ZN(n1139) );
OR2_X1 U823 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U824 ( .A(n1148), .B(KEYINPUT32), .Z(n1144) );
NAND3_X1 U825 ( .A1(n1149), .A2(n1146), .A3(n1147), .ZN(n1148) );
XOR2_X1 U826 ( .A(n1150), .B(n1151), .Z(n1147) );
XOR2_X1 U827 ( .A(G131), .B(n1152), .Z(n1151) );
NOR2_X1 U828 ( .A1(KEYINPUT8), .A2(n1153), .ZN(n1152) );
XNOR2_X1 U829 ( .A(G137), .B(n1154), .ZN(n1153) );
NAND2_X1 U830 ( .A1(KEYINPUT29), .A2(n1155), .ZN(n1154) );
XNOR2_X1 U831 ( .A(n1156), .B(n1157), .ZN(n1150) );
NAND2_X1 U832 ( .A1(n1158), .A2(n1084), .ZN(n1146) );
NAND2_X1 U833 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XNOR2_X1 U834 ( .A(n1161), .B(KEYINPUT9), .ZN(n1159) );
NAND2_X1 U835 ( .A1(G953), .A2(n1143), .ZN(n1149) );
XOR2_X1 U836 ( .A(n1162), .B(n1163), .Z(G69) );
XOR2_X1 U837 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U838 ( .A1(G953), .A2(n1166), .ZN(n1165) );
NAND2_X1 U839 ( .A1(G898), .A2(G224), .ZN(n1166) );
NAND2_X1 U840 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
NAND2_X1 U841 ( .A1(G953), .A2(n1169), .ZN(n1168) );
XOR2_X1 U842 ( .A(n1170), .B(n1171), .Z(n1167) );
XNOR2_X1 U843 ( .A(n1172), .B(KEYINPUT50), .ZN(n1171) );
NAND2_X1 U844 ( .A1(KEYINPUT27), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U845 ( .A(n1174), .B(n1175), .ZN(n1170) );
NOR2_X1 U846 ( .A1(n1176), .A2(G953), .ZN(n1162) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1178), .ZN(G66) );
XNOR2_X1 U848 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U849 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U850 ( .A(n1103), .B(KEYINPUT23), .Z(n1181) );
NOR2_X1 U851 ( .A1(n1084), .A2(n1183), .ZN(n1177) );
XNOR2_X1 U852 ( .A(KEYINPUT43), .B(n1184), .ZN(n1183) );
NOR2_X1 U853 ( .A1(n1185), .A2(n1186), .ZN(G63) );
XOR2_X1 U854 ( .A(n1187), .B(n1188), .Z(n1186) );
AND2_X1 U855 ( .A1(G478), .A2(n1189), .ZN(n1187) );
NOR2_X1 U856 ( .A1(n1185), .A2(n1190), .ZN(G60) );
NOR3_X1 U857 ( .A1(n1099), .A2(n1191), .A3(n1192), .ZN(n1190) );
AND3_X1 U858 ( .A1(n1193), .A2(G475), .A3(n1189), .ZN(n1192) );
NOR2_X1 U859 ( .A1(n1194), .A2(n1193), .ZN(n1191) );
AND2_X1 U860 ( .A1(n1082), .A2(G475), .ZN(n1194) );
NAND2_X1 U861 ( .A1(n1195), .A2(n1196), .ZN(G6) );
NAND2_X1 U862 ( .A1(G104), .A2(n1197), .ZN(n1196) );
XOR2_X1 U863 ( .A(n1198), .B(KEYINPUT6), .Z(n1195) );
OR2_X1 U864 ( .A1(n1197), .A2(G104), .ZN(n1198) );
NAND4_X1 U865 ( .A1(n1199), .A2(n1119), .A3(n1200), .A4(n1201), .ZN(n1197) );
NOR2_X1 U866 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XNOR2_X1 U867 ( .A(KEYINPUT46), .B(n1204), .ZN(n1203) );
NOR2_X1 U868 ( .A1(n1185), .A2(n1205), .ZN(G57) );
NOR2_X1 U869 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XOR2_X1 U870 ( .A(n1208), .B(KEYINPUT48), .Z(n1207) );
NAND2_X1 U871 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NOR2_X1 U872 ( .A1(n1209), .A2(n1210), .ZN(n1206) );
XNOR2_X1 U873 ( .A(G101), .B(n1211), .ZN(n1210) );
NOR2_X1 U874 ( .A1(KEYINPUT18), .A2(n1212), .ZN(n1211) );
AND2_X1 U875 ( .A1(n1213), .A2(n1214), .ZN(n1209) );
NAND3_X1 U876 ( .A1(n1189), .A2(G472), .A3(n1215), .ZN(n1214) );
XOR2_X1 U877 ( .A(KEYINPUT25), .B(n1216), .Z(n1215) );
NAND2_X1 U878 ( .A1(n1217), .A2(n1218), .ZN(n1213) );
NAND2_X1 U879 ( .A1(n1189), .A2(G472), .ZN(n1218) );
XNOR2_X1 U880 ( .A(n1216), .B(KEYINPUT25), .ZN(n1217) );
NOR3_X1 U881 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(G54) );
NOR3_X1 U882 ( .A1(n1222), .A2(G953), .A3(n1184), .ZN(n1221) );
AND2_X1 U883 ( .A1(n1222), .A2(n1185), .ZN(n1220) );
INV_X1 U884 ( .A(KEYINPUT44), .ZN(n1222) );
XOR2_X1 U885 ( .A(n1223), .B(n1224), .Z(n1219) );
AND2_X1 U886 ( .A1(G469), .A2(n1189), .ZN(n1224) );
INV_X1 U887 ( .A(n1182), .ZN(n1189) );
NAND2_X1 U888 ( .A1(KEYINPUT21), .A2(n1225), .ZN(n1223) );
XOR2_X1 U889 ( .A(n1226), .B(n1227), .Z(n1225) );
XNOR2_X1 U890 ( .A(n1228), .B(n1229), .ZN(n1227) );
NOR2_X1 U891 ( .A1(KEYINPUT7), .A2(n1230), .ZN(n1229) );
XOR2_X1 U892 ( .A(n1231), .B(n1232), .Z(n1230) );
NOR2_X1 U893 ( .A1(KEYINPUT30), .A2(n1233), .ZN(n1232) );
XOR2_X1 U894 ( .A(n1234), .B(KEYINPUT53), .Z(n1226) );
NAND2_X1 U895 ( .A1(n1235), .A2(KEYINPUT49), .ZN(n1234) );
XOR2_X1 U896 ( .A(n1236), .B(n1237), .Z(n1235) );
XNOR2_X1 U897 ( .A(n1238), .B(n1239), .ZN(n1237) );
XNOR2_X1 U898 ( .A(G140), .B(KEYINPUT12), .ZN(n1236) );
NOR2_X1 U899 ( .A1(n1185), .A2(n1240), .ZN(G51) );
XOR2_X1 U900 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U901 ( .A1(n1243), .A2(n1182), .ZN(n1241) );
NAND2_X1 U902 ( .A1(G902), .A2(n1082), .ZN(n1182) );
NAND3_X1 U903 ( .A1(n1176), .A2(n1160), .A3(n1161), .ZN(n1082) );
AND4_X1 U904 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1161) );
AND4_X1 U905 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1160) );
NAND4_X1 U906 ( .A1(n1252), .A2(n1253), .A3(n1199), .A4(n1254), .ZN(n1248) );
INV_X1 U907 ( .A(n1255), .ZN(n1199) );
XNOR2_X1 U908 ( .A(n1123), .B(KEYINPUT37), .ZN(n1252) );
AND4_X1 U909 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1176) );
NOR4_X1 U910 ( .A1(n1078), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1259) );
NOR3_X1 U911 ( .A1(n1113), .A2(n1263), .A3(n1264), .ZN(n1078) );
INV_X1 U912 ( .A(n1123), .ZN(n1264) );
NOR3_X1 U913 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1258) );
NOR3_X1 U914 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1267) );
NOR4_X1 U915 ( .A1(n1271), .A2(n1255), .A3(n1113), .A4(n1202), .ZN(n1269) );
INV_X1 U916 ( .A(KEYINPUT62), .ZN(n1268) );
NOR4_X1 U917 ( .A1(KEYINPUT62), .A2(n1202), .A3(n1263), .A4(n1113), .ZN(n1266) );
INV_X1 U918 ( .A(n1272), .ZN(n1263) );
INV_X1 U919 ( .A(n1124), .ZN(n1202) );
NOR2_X1 U920 ( .A1(n1084), .A2(n1184), .ZN(n1185) );
XNOR2_X1 U921 ( .A(G952), .B(KEYINPUT63), .ZN(n1184) );
XNOR2_X1 U922 ( .A(G146), .B(n1244), .ZN(G48) );
NAND4_X1 U923 ( .A1(n1253), .A2(n1124), .A3(n1254), .A4(n1134), .ZN(n1244) );
XNOR2_X1 U924 ( .A(G143), .B(n1245), .ZN(G45) );
NAND3_X1 U925 ( .A1(n1130), .A2(n1253), .A3(n1273), .ZN(n1245) );
NOR3_X1 U926 ( .A1(n1274), .A2(n1275), .A3(n1086), .ZN(n1273) );
XNOR2_X1 U927 ( .A(G140), .B(n1246), .ZN(G42) );
NAND3_X1 U928 ( .A1(n1131), .A2(n1276), .A3(n1124), .ZN(n1246) );
XNOR2_X1 U929 ( .A(G137), .B(n1247), .ZN(G39) );
NAND3_X1 U930 ( .A1(n1276), .A2(n1138), .A3(n1254), .ZN(n1247) );
XNOR2_X1 U931 ( .A(G134), .B(n1249), .ZN(G36) );
NAND3_X1 U932 ( .A1(n1276), .A2(n1123), .A3(n1130), .ZN(n1249) );
XNOR2_X1 U933 ( .A(G131), .B(n1251), .ZN(G33) );
NAND3_X1 U934 ( .A1(n1124), .A2(n1276), .A3(n1130), .ZN(n1251) );
NOR3_X1 U935 ( .A1(n1274), .A2(n1277), .A3(n1122), .ZN(n1276) );
NAND2_X1 U936 ( .A1(n1278), .A2(n1279), .ZN(n1122) );
XNOR2_X1 U937 ( .A(n1092), .B(KEYINPUT22), .ZN(n1278) );
INV_X1 U938 ( .A(n1134), .ZN(n1274) );
XNOR2_X1 U939 ( .A(n1280), .B(KEYINPUT17), .ZN(n1134) );
XNOR2_X1 U940 ( .A(G128), .B(n1281), .ZN(G30) );
NAND4_X1 U941 ( .A1(n1253), .A2(n1254), .A3(n1282), .A4(n1123), .ZN(n1281) );
NOR2_X1 U942 ( .A1(KEYINPUT35), .A2(n1255), .ZN(n1282) );
XOR2_X1 U943 ( .A(G101), .B(n1265), .Z(G3) );
AND3_X1 U944 ( .A1(n1138), .A2(n1272), .A3(n1130), .ZN(n1265) );
XNOR2_X1 U945 ( .A(G125), .B(n1250), .ZN(G27) );
NAND4_X1 U946 ( .A1(n1087), .A2(n1253), .A3(n1124), .A4(n1131), .ZN(n1250) );
NOR2_X1 U947 ( .A1(n1270), .A2(n1277), .ZN(n1253) );
AND2_X1 U948 ( .A1(n1108), .A2(n1283), .ZN(n1277) );
NAND2_X1 U949 ( .A1(n1284), .A2(n1143), .ZN(n1283) );
INV_X1 U950 ( .A(G900), .ZN(n1143) );
XNOR2_X1 U951 ( .A(G122), .B(n1256), .ZN(G24) );
NAND4_X1 U952 ( .A1(n1285), .A2(n1200), .A3(n1286), .A4(n1287), .ZN(n1256) );
INV_X1 U953 ( .A(n1113), .ZN(n1200) );
NAND2_X1 U954 ( .A1(n1288), .A2(n1289), .ZN(n1113) );
INV_X1 U955 ( .A(n1106), .ZN(n1289) );
XNOR2_X1 U956 ( .A(G119), .B(n1257), .ZN(G21) );
NAND3_X1 U957 ( .A1(n1254), .A2(n1138), .A3(n1285), .ZN(n1257) );
AND2_X1 U958 ( .A1(n1290), .A2(n1106), .ZN(n1254) );
XOR2_X1 U959 ( .A(KEYINPUT15), .B(n1291), .Z(n1290) );
NAND3_X1 U960 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(G18) );
NAND2_X1 U961 ( .A1(G116), .A2(n1295), .ZN(n1294) );
NAND2_X1 U962 ( .A1(n1296), .A2(n1297), .ZN(n1293) );
INV_X1 U963 ( .A(KEYINPUT10), .ZN(n1297) );
NAND2_X1 U964 ( .A1(n1298), .A2(n1262), .ZN(n1296) );
INV_X1 U965 ( .A(n1295), .ZN(n1262) );
XNOR2_X1 U966 ( .A(KEYINPUT54), .B(G116), .ZN(n1298) );
NAND2_X1 U967 ( .A1(KEYINPUT10), .A2(n1299), .ZN(n1292) );
NAND2_X1 U968 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
OR3_X1 U969 ( .A1(n1295), .A2(G116), .A3(KEYINPUT54), .ZN(n1301) );
NAND3_X1 U970 ( .A1(n1130), .A2(n1123), .A3(n1285), .ZN(n1295) );
NOR2_X1 U971 ( .A1(n1287), .A2(n1086), .ZN(n1123) );
INV_X1 U972 ( .A(n1286), .ZN(n1086) );
NAND2_X1 U973 ( .A1(KEYINPUT54), .A2(G116), .ZN(n1300) );
XOR2_X1 U974 ( .A(G113), .B(n1261), .Z(G15) );
AND3_X1 U975 ( .A1(n1130), .A2(n1124), .A3(n1285), .ZN(n1261) );
NOR3_X1 U976 ( .A1(n1270), .A2(n1271), .A3(n1111), .ZN(n1285) );
INV_X1 U977 ( .A(n1087), .ZN(n1111) );
NOR2_X1 U978 ( .A1(n1137), .A2(n1302), .ZN(n1087) );
INV_X1 U979 ( .A(n1136), .ZN(n1302) );
NOR2_X1 U980 ( .A1(n1286), .A2(n1275), .ZN(n1124) );
AND2_X1 U981 ( .A1(n1288), .A2(n1106), .ZN(n1130) );
NAND3_X1 U982 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(G12) );
NAND2_X1 U983 ( .A1(G110), .A2(n1306), .ZN(n1305) );
NAND2_X1 U984 ( .A1(n1307), .A2(n1308), .ZN(n1304) );
INV_X1 U985 ( .A(KEYINPUT13), .ZN(n1308) );
NAND2_X1 U986 ( .A1(n1309), .A2(n1238), .ZN(n1307) );
XNOR2_X1 U987 ( .A(n1260), .B(KEYINPUT41), .ZN(n1309) );
NAND2_X1 U988 ( .A1(KEYINPUT13), .A2(n1310), .ZN(n1303) );
NAND2_X1 U989 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
OR2_X1 U990 ( .A1(n1260), .A2(KEYINPUT41), .ZN(n1312) );
NAND3_X1 U991 ( .A1(n1260), .A2(n1238), .A3(KEYINPUT41), .ZN(n1311) );
INV_X1 U992 ( .A(n1306), .ZN(n1260) );
NAND3_X1 U993 ( .A1(n1138), .A2(n1272), .A3(n1131), .ZN(n1306) );
NOR2_X1 U994 ( .A1(n1291), .A2(n1106), .ZN(n1131) );
XNOR2_X1 U995 ( .A(n1313), .B(G472), .ZN(n1106) );
NAND2_X1 U996 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XNOR2_X1 U997 ( .A(n1216), .B(n1316), .ZN(n1314) );
XOR2_X1 U998 ( .A(n1212), .B(n1317), .Z(n1316) );
NAND2_X1 U999 ( .A1(KEYINPUT14), .A2(G101), .ZN(n1317) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1318), .ZN(n1212) );
XNOR2_X1 U1001 ( .A(n1319), .B(n1320), .ZN(n1216) );
XNOR2_X1 U1002 ( .A(n1321), .B(n1174), .ZN(n1320) );
XOR2_X1 U1003 ( .A(n1288), .B(KEYINPUT26), .Z(n1291) );
NOR2_X1 U1004 ( .A1(n1322), .A2(n1090), .ZN(n1288) );
NOR2_X1 U1005 ( .A1(n1103), .A2(n1104), .ZN(n1090) );
AND2_X1 U1006 ( .A1(n1104), .A2(n1103), .ZN(n1322) );
NAND2_X1 U1007 ( .A1(G217), .A2(n1323), .ZN(n1103) );
NOR2_X1 U1008 ( .A1(n1324), .A2(G902), .ZN(n1104) );
INV_X1 U1009 ( .A(n1179), .ZN(n1324) );
XNOR2_X1 U1010 ( .A(n1325), .B(n1326), .ZN(n1179) );
XOR2_X1 U1011 ( .A(n1327), .B(n1156), .Z(n1326) );
XOR2_X1 U1012 ( .A(G125), .B(G140), .Z(n1156) );
NOR2_X1 U1013 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
INV_X1 U1014 ( .A(G221), .ZN(n1329) );
XOR2_X1 U1015 ( .A(n1330), .B(n1331), .Z(n1325) );
NOR2_X1 U1016 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XOR2_X1 U1017 ( .A(n1334), .B(KEYINPUT2), .Z(n1333) );
NAND2_X1 U1018 ( .A1(G110), .A2(n1335), .ZN(n1334) );
NOR2_X1 U1019 ( .A1(G110), .A2(n1335), .ZN(n1332) );
XOR2_X1 U1020 ( .A(n1336), .B(G128), .Z(n1335) );
NAND2_X1 U1021 ( .A1(KEYINPUT3), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1022 ( .A(G137), .B(G146), .ZN(n1330) );
NOR3_X1 U1023 ( .A1(n1255), .A2(n1271), .A3(n1270), .ZN(n1272) );
INV_X1 U1024 ( .A(n1119), .ZN(n1270) );
NOR2_X1 U1025 ( .A1(n1279), .A2(n1092), .ZN(n1119) );
INV_X1 U1026 ( .A(n1120), .ZN(n1092) );
NAND2_X1 U1027 ( .A1(G214), .A2(n1338), .ZN(n1120) );
INV_X1 U1028 ( .A(n1105), .ZN(n1279) );
XOR2_X1 U1029 ( .A(n1339), .B(n1243), .Z(n1105) );
NAND2_X1 U1030 ( .A1(G210), .A2(n1338), .ZN(n1243) );
NAND2_X1 U1031 ( .A1(n1340), .A2(n1315), .ZN(n1338) );
XNOR2_X1 U1032 ( .A(G237), .B(KEYINPUT60), .ZN(n1340) );
OR2_X1 U1033 ( .A1(n1242), .A2(G902), .ZN(n1339) );
XNOR2_X1 U1034 ( .A(n1341), .B(n1342), .ZN(n1242) );
XNOR2_X1 U1035 ( .A(n1175), .B(n1319), .ZN(n1342) );
NAND2_X1 U1036 ( .A1(n1343), .A2(n1344), .ZN(n1319) );
NAND2_X1 U1037 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
NAND2_X1 U1038 ( .A1(n1347), .A2(G146), .ZN(n1343) );
XOR2_X1 U1039 ( .A(KEYINPUT52), .B(n1345), .Z(n1347) );
XNOR2_X1 U1040 ( .A(G122), .B(n1238), .ZN(n1175) );
XOR2_X1 U1041 ( .A(n1348), .B(n1349), .Z(n1341) );
AND2_X1 U1042 ( .A1(n1084), .A2(G224), .ZN(n1349) );
XNOR2_X1 U1043 ( .A(n1350), .B(n1351), .ZN(n1348) );
NAND2_X1 U1044 ( .A1(n1352), .A2(n1353), .ZN(n1350) );
NAND2_X1 U1045 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XNOR2_X1 U1046 ( .A(KEYINPUT57), .B(n1356), .ZN(n1355) );
XOR2_X1 U1047 ( .A(KEYINPUT38), .B(n1357), .Z(n1352) );
NOR2_X1 U1048 ( .A1(n1356), .A2(n1354), .ZN(n1357) );
INV_X1 U1049 ( .A(n1173), .ZN(n1354) );
XNOR2_X1 U1050 ( .A(n1358), .B(n1359), .ZN(n1173) );
XNOR2_X1 U1051 ( .A(n1360), .B(G101), .ZN(n1359) );
NAND2_X1 U1052 ( .A1(KEYINPUT33), .A2(G107), .ZN(n1358) );
INV_X1 U1053 ( .A(n1174), .ZN(n1356) );
XOR2_X1 U1054 ( .A(G113), .B(n1361), .Z(n1174) );
XNOR2_X1 U1055 ( .A(n1337), .B(G116), .ZN(n1361) );
INV_X1 U1056 ( .A(G119), .ZN(n1337) );
INV_X1 U1057 ( .A(n1204), .ZN(n1271) );
NAND2_X1 U1058 ( .A1(n1108), .A2(n1362), .ZN(n1204) );
NAND2_X1 U1059 ( .A1(n1284), .A2(n1169), .ZN(n1362) );
INV_X1 U1060 ( .A(G898), .ZN(n1169) );
AND3_X1 U1061 ( .A1(n1363), .A2(n1364), .A3(G953), .ZN(n1284) );
XNOR2_X1 U1062 ( .A(KEYINPUT58), .B(n1315), .ZN(n1363) );
NAND3_X1 U1063 ( .A1(n1364), .A2(n1084), .A3(G952), .ZN(n1108) );
NAND2_X1 U1064 ( .A1(G237), .A2(G234), .ZN(n1364) );
XNOR2_X1 U1065 ( .A(n1280), .B(KEYINPUT4), .ZN(n1255) );
NAND2_X1 U1066 ( .A1(n1365), .A2(n1137), .ZN(n1280) );
XNOR2_X1 U1067 ( .A(n1366), .B(G469), .ZN(n1137) );
NAND2_X1 U1068 ( .A1(n1367), .A2(n1315), .ZN(n1366) );
XOR2_X1 U1069 ( .A(n1368), .B(n1369), .Z(n1367) );
XNOR2_X1 U1070 ( .A(n1370), .B(n1321), .ZN(n1369) );
INV_X1 U1071 ( .A(n1228), .ZN(n1321) );
XOR2_X1 U1072 ( .A(G131), .B(n1371), .Z(n1228) );
XNOR2_X1 U1073 ( .A(n1372), .B(G134), .ZN(n1371) );
INV_X1 U1074 ( .A(G137), .ZN(n1372) );
XNOR2_X1 U1075 ( .A(n1231), .B(n1233), .ZN(n1370) );
INV_X1 U1076 ( .A(n1157), .ZN(n1233) );
XNOR2_X1 U1077 ( .A(n1373), .B(n1374), .ZN(n1157) );
NOR2_X1 U1078 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
XOR2_X1 U1079 ( .A(n1377), .B(KEYINPUT16), .Z(n1376) );
NAND2_X1 U1080 ( .A1(G143), .A2(n1346), .ZN(n1377) );
NOR2_X1 U1081 ( .A1(G143), .A2(n1346), .ZN(n1375) );
NAND2_X1 U1082 ( .A1(n1378), .A2(KEYINPUT51), .ZN(n1373) );
XNOR2_X1 U1083 ( .A(G128), .B(KEYINPUT28), .ZN(n1378) );
XOR2_X1 U1084 ( .A(n1379), .B(n1380), .Z(n1231) );
XNOR2_X1 U1085 ( .A(n1077), .B(G101), .ZN(n1380) );
NAND2_X1 U1086 ( .A1(KEYINPUT40), .A2(n1360), .ZN(n1379) );
XOR2_X1 U1087 ( .A(n1381), .B(n1382), .Z(n1368) );
XOR2_X1 U1088 ( .A(KEYINPUT31), .B(G140), .Z(n1382) );
XOR2_X1 U1089 ( .A(n1383), .B(n1239), .Z(n1381) );
NOR2_X1 U1090 ( .A1(n1142), .A2(G953), .ZN(n1239) );
INV_X1 U1091 ( .A(G227), .ZN(n1142) );
NAND2_X1 U1092 ( .A1(KEYINPUT59), .A2(n1238), .ZN(n1383) );
INV_X1 U1093 ( .A(G110), .ZN(n1238) );
XNOR2_X1 U1094 ( .A(KEYINPUT19), .B(n1136), .ZN(n1365) );
NAND2_X1 U1095 ( .A1(G221), .A2(n1323), .ZN(n1136) );
NAND2_X1 U1096 ( .A1(G234), .A2(n1315), .ZN(n1323) );
INV_X1 U1097 ( .A(G902), .ZN(n1315) );
NOR2_X1 U1098 ( .A1(n1286), .A2(n1287), .ZN(n1138) );
INV_X1 U1099 ( .A(n1275), .ZN(n1287) );
XNOR2_X1 U1100 ( .A(n1100), .B(n1098), .ZN(n1275) );
INV_X1 U1101 ( .A(G475), .ZN(n1098) );
INV_X1 U1102 ( .A(n1099), .ZN(n1100) );
NOR2_X1 U1103 ( .A1(n1193), .A2(G902), .ZN(n1099) );
XOR2_X1 U1104 ( .A(n1384), .B(n1385), .Z(n1193) );
XNOR2_X1 U1105 ( .A(n1346), .B(n1386), .ZN(n1385) );
NOR2_X1 U1106 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
XOR2_X1 U1107 ( .A(n1389), .B(KEYINPUT47), .Z(n1388) );
NAND2_X1 U1108 ( .A1(G140), .A2(n1390), .ZN(n1389) );
NOR2_X1 U1109 ( .A1(G140), .A2(n1390), .ZN(n1387) );
XNOR2_X1 U1110 ( .A(KEYINPUT55), .B(n1351), .ZN(n1390) );
INV_X1 U1111 ( .A(G125), .ZN(n1351) );
INV_X1 U1112 ( .A(G146), .ZN(n1346) );
XNOR2_X1 U1113 ( .A(n1391), .B(n1392), .ZN(n1384) );
NAND2_X1 U1114 ( .A1(KEYINPUT24), .A2(n1393), .ZN(n1392) );
XOR2_X1 U1115 ( .A(n1394), .B(n1395), .Z(n1393) );
XNOR2_X1 U1116 ( .A(G131), .B(G143), .ZN(n1395) );
NAND2_X1 U1117 ( .A1(G214), .A2(n1318), .ZN(n1394) );
NOR2_X1 U1118 ( .A1(G953), .A2(G237), .ZN(n1318) );
NAND2_X1 U1119 ( .A1(n1396), .A2(KEYINPUT1), .ZN(n1391) );
XOR2_X1 U1120 ( .A(n1397), .B(n1398), .Z(n1396) );
XNOR2_X1 U1121 ( .A(n1360), .B(n1399), .ZN(n1398) );
NOR2_X1 U1122 ( .A1(G113), .A2(KEYINPUT56), .ZN(n1399) );
INV_X1 U1123 ( .A(G104), .ZN(n1360) );
XNOR2_X1 U1124 ( .A(G122), .B(KEYINPUT36), .ZN(n1397) );
XNOR2_X1 U1125 ( .A(n1400), .B(G478), .ZN(n1286) );
OR2_X1 U1126 ( .A1(n1188), .A2(G902), .ZN(n1400) );
XNOR2_X1 U1127 ( .A(n1401), .B(n1402), .ZN(n1188) );
XOR2_X1 U1128 ( .A(n1403), .B(n1404), .Z(n1402) );
NOR2_X1 U1129 ( .A1(n1328), .A2(n1405), .ZN(n1404) );
INV_X1 U1130 ( .A(G217), .ZN(n1405) );
NAND2_X1 U1131 ( .A1(n1406), .A2(n1084), .ZN(n1328) );
INV_X1 U1132 ( .A(G953), .ZN(n1084) );
XOR2_X1 U1133 ( .A(KEYINPUT34), .B(G234), .Z(n1406) );
NOR2_X1 U1134 ( .A1(KEYINPUT11), .A2(n1077), .ZN(n1403) );
INV_X1 U1135 ( .A(G107), .ZN(n1077) );
XOR2_X1 U1136 ( .A(n1407), .B(n1408), .Z(n1401) );
XNOR2_X1 U1137 ( .A(n1409), .B(G116), .ZN(n1408) );
INV_X1 U1138 ( .A(G122), .ZN(n1409) );
NAND2_X1 U1139 ( .A1(KEYINPUT45), .A2(n1410), .ZN(n1407) );
XNOR2_X1 U1140 ( .A(n1411), .B(n1345), .ZN(n1410) );
XOR2_X1 U1141 ( .A(G128), .B(G143), .Z(n1345) );
NAND2_X1 U1142 ( .A1(KEYINPUT5), .A2(n1412), .ZN(n1411) );
XNOR2_X1 U1143 ( .A(KEYINPUT42), .B(n1155), .ZN(n1412) );
INV_X1 U1144 ( .A(G134), .ZN(n1155) );
endmodule


