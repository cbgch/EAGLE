//Key = 1100011011010110000010000100100000110100010101110101011011110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380;

XNOR2_X1 U764 ( .A(n1049), .B(n1050), .ZN(G9) );
NOR2_X1 U765 ( .A1(n1051), .A2(n1052), .ZN(G75) );
NOR3_X1 U766 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NAND3_X1 U767 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1053) );
XOR2_X1 U768 ( .A(KEYINPUT54), .B(n1059), .Z(n1058) );
NAND2_X1 U769 ( .A1(n1060), .A2(n1061), .ZN(n1056) );
NAND2_X1 U770 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U771 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NAND2_X1 U772 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NAND2_X1 U773 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U774 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U775 ( .A1(n1073), .A2(n1074), .ZN(n1067) );
NAND2_X1 U776 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND3_X1 U778 ( .A1(n1073), .A2(n1079), .A3(n1069), .ZN(n1062) );
NAND3_X1 U779 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NAND2_X1 U780 ( .A1(n1064), .A2(n1083), .ZN(n1082) );
NAND2_X1 U781 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U782 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
INV_X1 U783 ( .A(n1088), .ZN(n1084) );
NAND2_X1 U784 ( .A1(n1066), .A2(n1089), .ZN(n1081) );
NAND2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U786 ( .A1(KEYINPUT43), .A2(n1092), .ZN(n1091) );
OR3_X1 U787 ( .A1(n1093), .A2(KEYINPUT43), .A3(n1066), .ZN(n1080) );
INV_X1 U788 ( .A(n1094), .ZN(n1060) );
NOR3_X1 U789 ( .A1(n1095), .A2(G953), .A3(n1059), .ZN(n1051) );
AND4_X1 U790 ( .A1(n1096), .A2(n1077), .A3(n1097), .A4(n1098), .ZN(n1059) );
NOR4_X1 U791 ( .A1(n1099), .A2(n1100), .A3(n1078), .A4(n1101), .ZN(n1098) );
INV_X1 U792 ( .A(n1102), .ZN(n1100) );
NAND2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1099) );
NOR3_X1 U794 ( .A1(n1105), .A2(n1087), .A3(n1106), .ZN(n1097) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(n1096) );
NOR2_X1 U796 ( .A1(KEYINPUT44), .A2(n1109), .ZN(n1108) );
XOR2_X1 U797 ( .A(KEYINPUT17), .B(n1110), .Z(n1109) );
XNOR2_X1 U798 ( .A(G478), .B(KEYINPUT9), .ZN(n1107) );
XNOR2_X1 U799 ( .A(KEYINPUT23), .B(n1054), .ZN(n1095) );
INV_X1 U800 ( .A(G952), .ZN(n1054) );
XOR2_X1 U801 ( .A(n1111), .B(n1112), .Z(G72) );
NOR2_X1 U802 ( .A1(n1113), .A2(n1057), .ZN(n1112) );
AND2_X1 U803 ( .A1(G227), .A2(G900), .ZN(n1113) );
NAND2_X1 U804 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U805 ( .A1(n1116), .A2(n1057), .ZN(n1115) );
XOR2_X1 U806 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U807 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
XNOR2_X1 U808 ( .A(n1121), .B(KEYINPUT51), .ZN(n1119) );
NAND3_X1 U809 ( .A1(n1118), .A2(G900), .A3(G953), .ZN(n1114) );
NOR2_X1 U810 ( .A1(KEYINPUT10), .A2(n1122), .ZN(n1118) );
XOR2_X1 U811 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U812 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U813 ( .A1(KEYINPUT20), .A2(n1127), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1128), .B(n1129), .Z(n1123) );
NOR2_X1 U815 ( .A1(KEYINPUT26), .A2(n1130), .ZN(n1129) );
NOR2_X1 U816 ( .A1(n1131), .A2(n1132), .ZN(n1128) );
XOR2_X1 U817 ( .A(KEYINPUT42), .B(n1133), .Z(n1132) );
NOR2_X1 U818 ( .A1(G140), .A2(n1134), .ZN(n1133) );
AND2_X1 U819 ( .A1(n1134), .A2(G140), .ZN(n1131) );
XOR2_X1 U820 ( .A(n1135), .B(n1136), .Z(G69) );
XOR2_X1 U821 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U822 ( .A1(G953), .A2(n1139), .ZN(n1138) );
OR2_X1 U823 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
NAND2_X1 U824 ( .A1(G953), .A2(n1142), .ZN(n1135) );
NAND2_X1 U825 ( .A1(G898), .A2(G224), .ZN(n1142) );
NOR2_X1 U826 ( .A1(n1143), .A2(n1144), .ZN(G66) );
XNOR2_X1 U827 ( .A(n1145), .B(n1146), .ZN(n1144) );
NOR2_X1 U828 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NOR2_X1 U829 ( .A1(n1143), .A2(n1149), .ZN(G63) );
NOR3_X1 U830 ( .A1(n1110), .A2(n1150), .A3(n1151), .ZN(n1149) );
NOR3_X1 U831 ( .A1(n1152), .A2(n1153), .A3(n1148), .ZN(n1151) );
NOR2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(n1150) );
AND2_X1 U833 ( .A1(n1055), .A2(G478), .ZN(n1154) );
NOR2_X1 U834 ( .A1(n1143), .A2(n1156), .ZN(G60) );
XNOR2_X1 U835 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR2_X1 U836 ( .A1(n1159), .A2(n1148), .ZN(n1158) );
XOR2_X1 U837 ( .A(n1160), .B(G104), .Z(G6) );
NAND2_X1 U838 ( .A1(KEYINPUT8), .A2(n1161), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1143), .A2(n1162), .ZN(G57) );
NOR2_X1 U840 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U841 ( .A(KEYINPUT2), .B(n1165), .Z(n1164) );
NOR2_X1 U842 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U843 ( .A(KEYINPUT22), .B(n1168), .Z(n1167) );
AND2_X1 U844 ( .A1(n1168), .A2(n1166), .ZN(n1163) );
XNOR2_X1 U845 ( .A(n1169), .B(n1170), .ZN(n1166) );
NOR2_X1 U846 ( .A1(n1171), .A2(n1148), .ZN(n1170) );
NOR2_X1 U847 ( .A1(n1143), .A2(n1172), .ZN(G54) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U849 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U850 ( .A1(KEYINPUT62), .A2(n1177), .ZN(n1175) );
XOR2_X1 U851 ( .A(KEYINPUT48), .B(n1178), .Z(n1173) );
NOR2_X1 U852 ( .A1(n1148), .A2(n1179), .ZN(n1178) );
XNOR2_X1 U853 ( .A(KEYINPUT53), .B(n1180), .ZN(n1179) );
NOR2_X1 U854 ( .A1(n1143), .A2(n1181), .ZN(G51) );
XOR2_X1 U855 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U856 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U857 ( .A1(n1186), .A2(n1148), .ZN(n1184) );
NAND2_X1 U858 ( .A1(G902), .A2(n1055), .ZN(n1148) );
NAND3_X1 U859 ( .A1(n1121), .A2(n1120), .A3(n1139), .ZN(n1055) );
AND2_X1 U860 ( .A1(n1187), .A2(n1188), .ZN(n1139) );
NOR4_X1 U861 ( .A1(n1189), .A2(n1050), .A3(n1190), .A4(n1191), .ZN(n1188) );
NOR4_X1 U862 ( .A1(n1192), .A2(n1193), .A3(n1072), .A4(n1093), .ZN(n1190) );
NOR2_X1 U863 ( .A1(KEYINPUT6), .A2(n1194), .ZN(n1193) );
NOR3_X1 U864 ( .A1(n1195), .A2(n1075), .A3(n1196), .ZN(n1194) );
NOR2_X1 U865 ( .A1(n1197), .A2(n1198), .ZN(n1192) );
INV_X1 U866 ( .A(KEYINPUT6), .ZN(n1198) );
AND3_X1 U867 ( .A1(n1073), .A2(n1199), .A3(n1200), .ZN(n1050) );
NOR4_X1 U868 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1187) );
NOR3_X1 U869 ( .A1(n1071), .A2(n1205), .A3(n1206), .ZN(n1204) );
INV_X1 U870 ( .A(n1207), .ZN(n1071) );
INV_X1 U871 ( .A(n1161), .ZN(n1203) );
NAND3_X1 U872 ( .A1(n1073), .A2(n1199), .A3(n1092), .ZN(n1161) );
INV_X1 U873 ( .A(n1205), .ZN(n1199) );
AND4_X1 U874 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1120) );
NAND2_X1 U875 ( .A1(n1212), .A2(n1069), .ZN(n1208) );
AND4_X1 U876 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1121) );
NAND3_X1 U877 ( .A1(n1069), .A2(n1088), .A3(n1217), .ZN(n1213) );
XOR2_X1 U878 ( .A(n1218), .B(n1219), .Z(n1182) );
XOR2_X1 U879 ( .A(n1220), .B(n1221), .Z(n1219) );
NOR2_X1 U880 ( .A1(KEYINPUT52), .A2(n1222), .ZN(n1221) );
NOR2_X1 U881 ( .A1(KEYINPUT30), .A2(n1140), .ZN(n1218) );
NOR2_X1 U882 ( .A1(n1057), .A2(G952), .ZN(n1143) );
NAND2_X1 U883 ( .A1(n1223), .A2(n1224), .ZN(G48) );
NAND2_X1 U884 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U885 ( .A(KEYINPUT59), .B(n1227), .Z(n1223) );
NOR2_X1 U886 ( .A1(n1225), .A2(n1226), .ZN(n1227) );
INV_X1 U887 ( .A(n1214), .ZN(n1225) );
NAND4_X1 U888 ( .A1(n1228), .A2(n1092), .A3(n1229), .A4(n1088), .ZN(n1214) );
XNOR2_X1 U889 ( .A(G143), .B(n1215), .ZN(G45) );
NAND4_X1 U890 ( .A1(n1230), .A2(n1229), .A3(n1231), .A4(n1106), .ZN(n1215) );
XNOR2_X1 U891 ( .A(G140), .B(n1232), .ZN(G42) );
NAND3_X1 U892 ( .A1(n1217), .A2(n1069), .A3(n1233), .ZN(n1232) );
XNOR2_X1 U893 ( .A(n1088), .B(KEYINPUT25), .ZN(n1233) );
XNOR2_X1 U894 ( .A(G137), .B(n1216), .ZN(G39) );
NAND4_X1 U895 ( .A1(n1069), .A2(n1228), .A3(n1064), .A4(n1088), .ZN(n1216) );
XNOR2_X1 U896 ( .A(G134), .B(n1209), .ZN(G36) );
NAND3_X1 U897 ( .A1(n1069), .A2(n1200), .A3(n1230), .ZN(n1209) );
NAND2_X1 U898 ( .A1(n1234), .A2(n1235), .ZN(G33) );
OR2_X1 U899 ( .A1(n1236), .A2(G131), .ZN(n1235) );
XOR2_X1 U900 ( .A(n1237), .B(KEYINPUT31), .Z(n1234) );
NAND2_X1 U901 ( .A1(G131), .A2(n1236), .ZN(n1237) );
NAND2_X1 U902 ( .A1(n1238), .A2(n1069), .ZN(n1236) );
AND2_X1 U903 ( .A1(n1077), .A2(n1239), .ZN(n1069) );
XOR2_X1 U904 ( .A(KEYINPUT0), .B(n1078), .Z(n1239) );
XNOR2_X1 U905 ( .A(n1212), .B(KEYINPUT34), .ZN(n1238) );
AND2_X1 U906 ( .A1(n1230), .A2(n1092), .ZN(n1212) );
AND3_X1 U907 ( .A1(n1088), .A2(n1240), .A3(n1241), .ZN(n1230) );
XNOR2_X1 U908 ( .A(n1242), .B(KEYINPUT33), .ZN(n1088) );
XOR2_X1 U909 ( .A(n1210), .B(n1243), .Z(G30) );
NAND2_X1 U910 ( .A1(n1244), .A2(G128), .ZN(n1243) );
XNOR2_X1 U911 ( .A(KEYINPUT60), .B(KEYINPUT27), .ZN(n1244) );
NAND4_X1 U912 ( .A1(n1228), .A2(n1200), .A3(n1245), .A4(n1229), .ZN(n1210) );
AND3_X1 U913 ( .A1(n1246), .A2(n1240), .A3(n1105), .ZN(n1228) );
NAND2_X1 U914 ( .A1(n1247), .A2(n1248), .ZN(G3) );
NAND2_X1 U915 ( .A1(n1189), .A2(n1249), .ZN(n1248) );
XOR2_X1 U916 ( .A(KEYINPUT11), .B(n1250), .Z(n1247) );
NOR2_X1 U917 ( .A1(n1189), .A2(n1249), .ZN(n1250) );
INV_X1 U918 ( .A(G101), .ZN(n1249) );
NOR3_X1 U919 ( .A1(n1206), .A2(n1205), .A3(n1072), .ZN(n1189) );
NAND3_X1 U920 ( .A1(n1245), .A2(n1195), .A3(n1229), .ZN(n1205) );
XNOR2_X1 U921 ( .A(G125), .B(n1211), .ZN(G27) );
NAND3_X1 U922 ( .A1(n1066), .A2(n1229), .A3(n1217), .ZN(n1211) );
AND3_X1 U923 ( .A1(n1092), .A2(n1240), .A3(n1207), .ZN(n1217) );
NAND2_X1 U924 ( .A1(n1251), .A2(n1094), .ZN(n1240) );
NAND4_X1 U925 ( .A1(G902), .A2(G953), .A3(n1252), .A4(n1253), .ZN(n1251) );
INV_X1 U926 ( .A(G900), .ZN(n1253) );
INV_X1 U927 ( .A(n1196), .ZN(n1066) );
XNOR2_X1 U928 ( .A(n1202), .B(n1254), .ZN(G24) );
XOR2_X1 U929 ( .A(KEYINPUT57), .B(G122), .Z(n1254) );
AND4_X1 U930 ( .A1(n1197), .A2(n1073), .A3(n1231), .A4(n1106), .ZN(n1202) );
NOR2_X1 U931 ( .A1(n1246), .A2(n1105), .ZN(n1073) );
XOR2_X1 U932 ( .A(n1201), .B(n1255), .Z(G21) );
NOR2_X1 U933 ( .A1(KEYINPUT16), .A2(n1256), .ZN(n1255) );
AND4_X1 U934 ( .A1(n1197), .A2(n1064), .A3(n1105), .A4(n1246), .ZN(n1201) );
XNOR2_X1 U935 ( .A(n1257), .B(n1191), .ZN(G18) );
AND3_X1 U936 ( .A1(n1241), .A2(n1200), .A3(n1197), .ZN(n1191) );
INV_X1 U937 ( .A(n1090), .ZN(n1200) );
NAND2_X1 U938 ( .A1(n1258), .A2(n1231), .ZN(n1090) );
XOR2_X1 U939 ( .A(n1259), .B(KEYINPUT14), .Z(n1231) );
XNOR2_X1 U940 ( .A(G113), .B(n1260), .ZN(G15) );
NAND4_X1 U941 ( .A1(KEYINPUT49), .A2(n1197), .A3(n1092), .A4(n1241), .ZN(n1260) );
INV_X1 U942 ( .A(n1072), .ZN(n1241) );
NAND2_X1 U943 ( .A1(n1261), .A2(n1105), .ZN(n1072) );
INV_X1 U944 ( .A(n1093), .ZN(n1092) );
NAND2_X1 U945 ( .A1(n1259), .A2(n1106), .ZN(n1093) );
NOR3_X1 U946 ( .A1(n1075), .A2(n1262), .A3(n1196), .ZN(n1197) );
NAND2_X1 U947 ( .A1(n1086), .A2(n1263), .ZN(n1196) );
XOR2_X1 U948 ( .A(n1264), .B(KEYINPUT46), .Z(n1086) );
INV_X1 U949 ( .A(n1229), .ZN(n1075) );
XNOR2_X1 U950 ( .A(G110), .B(n1265), .ZN(G12) );
NAND4_X1 U951 ( .A1(n1207), .A2(n1064), .A3(n1266), .A4(n1245), .ZN(n1265) );
XOR2_X1 U952 ( .A(n1242), .B(KEYINPUT37), .Z(n1245) );
NAND2_X1 U953 ( .A1(n1263), .A2(n1264), .ZN(n1242) );
NAND3_X1 U954 ( .A1(n1267), .A2(n1268), .A3(n1103), .ZN(n1264) );
NAND2_X1 U955 ( .A1(n1269), .A2(n1180), .ZN(n1103) );
NAND2_X1 U956 ( .A1(KEYINPUT29), .A2(n1180), .ZN(n1268) );
OR2_X1 U957 ( .A1(n1104), .A2(KEYINPUT29), .ZN(n1267) );
OR2_X1 U958 ( .A1(n1180), .A2(n1269), .ZN(n1104) );
AND3_X1 U959 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1269) );
NAND2_X1 U960 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
INV_X1 U961 ( .A(KEYINPUT21), .ZN(n1274) );
XNOR2_X1 U962 ( .A(n1176), .B(n1177), .ZN(n1273) );
INV_X1 U963 ( .A(n1275), .ZN(n1177) );
NAND3_X1 U964 ( .A1(n1275), .A2(n1176), .A3(KEYINPUT21), .ZN(n1270) );
XNOR2_X1 U965 ( .A(n1276), .B(n1277), .ZN(n1176) );
NAND2_X1 U966 ( .A1(G227), .A2(n1057), .ZN(n1276) );
XNOR2_X1 U967 ( .A(n1278), .B(n1279), .ZN(n1275) );
XNOR2_X1 U968 ( .A(KEYINPUT15), .B(n1049), .ZN(n1279) );
XNOR2_X1 U969 ( .A(n1280), .B(n1281), .ZN(n1278) );
INV_X1 U970 ( .A(G469), .ZN(n1180) );
XNOR2_X1 U971 ( .A(n1087), .B(KEYINPUT3), .ZN(n1263) );
AND2_X1 U972 ( .A1(n1282), .A2(G221), .ZN(n1087) );
XOR2_X1 U973 ( .A(n1283), .B(KEYINPUT12), .Z(n1282) );
NOR2_X1 U974 ( .A1(n1262), .A2(n1284), .ZN(n1266) );
XNOR2_X1 U975 ( .A(n1229), .B(KEYINPUT24), .ZN(n1284) );
NOR2_X1 U976 ( .A1(n1285), .A2(n1077), .ZN(n1229) );
XNOR2_X1 U977 ( .A(n1286), .B(n1186), .ZN(n1077) );
NAND2_X1 U978 ( .A1(G210), .A2(n1287), .ZN(n1186) );
NAND2_X1 U979 ( .A1(n1288), .A2(n1272), .ZN(n1286) );
XOR2_X1 U980 ( .A(n1289), .B(n1140), .Z(n1288) );
XNOR2_X1 U981 ( .A(n1290), .B(n1291), .ZN(n1140) );
XOR2_X1 U982 ( .A(G122), .B(G110), .Z(n1291) );
XOR2_X1 U983 ( .A(n1292), .B(n1293), .Z(n1290) );
NOR2_X1 U984 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NOR2_X1 U985 ( .A1(G107), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U986 ( .A(KEYINPUT7), .B(n1281), .ZN(n1296) );
NOR2_X1 U987 ( .A1(n1049), .A2(n1281), .ZN(n1294) );
XNOR2_X1 U988 ( .A(G104), .B(G101), .ZN(n1281) );
INV_X1 U989 ( .A(G107), .ZN(n1049) );
NAND3_X1 U990 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1292) );
INV_X1 U991 ( .A(n1300), .ZN(n1299) );
NAND2_X1 U992 ( .A1(KEYINPUT36), .A2(n1301), .ZN(n1298) );
XOR2_X1 U993 ( .A(n1302), .B(n1303), .Z(n1301) );
NAND2_X1 U994 ( .A1(G119), .A2(n1257), .ZN(n1302) );
NAND2_X1 U995 ( .A1(n1304), .A2(n1305), .ZN(n1297) );
INV_X1 U996 ( .A(KEYINPUT36), .ZN(n1305) );
NAND3_X1 U997 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1289) );
NAND2_X1 U998 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND3_X1 U999 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1310) );
NAND2_X1 U1000 ( .A1(KEYINPUT4), .A2(n1314), .ZN(n1313) );
NAND2_X1 U1001 ( .A1(KEYINPUT50), .A2(n1220), .ZN(n1312) );
NAND2_X1 U1002 ( .A1(n1315), .A2(n1316), .ZN(n1311) );
INV_X1 U1003 ( .A(KEYINPUT50), .ZN(n1316) );
NAND2_X1 U1004 ( .A1(n1220), .A2(n1317), .ZN(n1315) );
NAND2_X1 U1005 ( .A1(KEYINPUT39), .A2(n1318), .ZN(n1317) );
INV_X1 U1006 ( .A(n1319), .ZN(n1309) );
NAND4_X1 U1007 ( .A1(n1319), .A2(n1314), .A3(n1220), .A4(n1318), .ZN(n1307) );
INV_X1 U1008 ( .A(KEYINPUT4), .ZN(n1318) );
INV_X1 U1009 ( .A(KEYINPUT39), .ZN(n1314) );
NAND2_X1 U1010 ( .A1(KEYINPUT4), .A2(n1320), .ZN(n1306) );
NAND2_X1 U1011 ( .A1(n1220), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1012 ( .A1(KEYINPUT39), .A2(n1319), .ZN(n1321) );
NAND3_X1 U1013 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1319) );
NAND2_X1 U1014 ( .A1(n1222), .A2(n1325), .ZN(n1324) );
INV_X1 U1015 ( .A(KEYINPUT35), .ZN(n1325) );
NAND3_X1 U1016 ( .A1(KEYINPUT35), .A2(n1326), .A3(n1185), .ZN(n1323) );
OR2_X1 U1017 ( .A1(n1185), .A2(n1326), .ZN(n1322) );
NOR2_X1 U1018 ( .A1(KEYINPUT38), .A2(n1222), .ZN(n1326) );
XOR2_X1 U1019 ( .A(G125), .B(KEYINPUT28), .Z(n1185) );
AND2_X1 U1020 ( .A1(G224), .A2(n1057), .ZN(n1220) );
XNOR2_X1 U1021 ( .A(KEYINPUT0), .B(n1078), .ZN(n1285) );
AND2_X1 U1022 ( .A1(G214), .A2(n1287), .ZN(n1078) );
NAND2_X1 U1023 ( .A1(n1327), .A2(n1272), .ZN(n1287) );
INV_X1 U1024 ( .A(n1195), .ZN(n1262) );
NAND2_X1 U1025 ( .A1(n1094), .A2(n1328), .ZN(n1195) );
NAND3_X1 U1026 ( .A1(n1141), .A2(n1252), .A3(G902), .ZN(n1328) );
NOR2_X1 U1027 ( .A1(n1057), .A2(G898), .ZN(n1141) );
NAND3_X1 U1028 ( .A1(n1252), .A2(n1057), .A3(G952), .ZN(n1094) );
NAND2_X1 U1029 ( .A1(G237), .A2(G234), .ZN(n1252) );
INV_X1 U1030 ( .A(n1206), .ZN(n1064) );
NAND2_X1 U1031 ( .A1(n1258), .A2(n1259), .ZN(n1206) );
XNOR2_X1 U1032 ( .A(n1329), .B(n1110), .ZN(n1259) );
NOR2_X1 U1033 ( .A1(n1155), .A2(G902), .ZN(n1110) );
INV_X1 U1034 ( .A(n1152), .ZN(n1155) );
XNOR2_X1 U1035 ( .A(n1330), .B(n1331), .ZN(n1152) );
XOR2_X1 U1036 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1037 ( .A(G122), .B(n1257), .ZN(n1333) );
XNOR2_X1 U1038 ( .A(n1334), .B(G128), .ZN(n1332) );
XOR2_X1 U1039 ( .A(n1335), .B(n1336), .Z(n1330) );
NOR2_X1 U1040 ( .A1(G107), .A2(KEYINPUT40), .ZN(n1336) );
XOR2_X1 U1041 ( .A(n1337), .B(n1338), .Z(n1335) );
NOR2_X1 U1042 ( .A1(G134), .A2(KEYINPUT32), .ZN(n1338) );
OR2_X1 U1043 ( .A1(n1147), .A2(n1339), .ZN(n1337) );
INV_X1 U1044 ( .A(G217), .ZN(n1147) );
NAND2_X1 U1045 ( .A1(KEYINPUT1), .A2(n1153), .ZN(n1329) );
INV_X1 U1046 ( .A(G478), .ZN(n1153) );
INV_X1 U1047 ( .A(n1106), .ZN(n1258) );
XOR2_X1 U1048 ( .A(n1340), .B(n1159), .Z(n1106) );
INV_X1 U1049 ( .A(G475), .ZN(n1159) );
NAND2_X1 U1050 ( .A1(n1157), .A2(n1272), .ZN(n1340) );
XNOR2_X1 U1051 ( .A(n1341), .B(n1342), .ZN(n1157) );
XOR2_X1 U1052 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1053 ( .A(n1134), .B(G122), .ZN(n1344) );
INV_X1 U1054 ( .A(G125), .ZN(n1134) );
XNOR2_X1 U1055 ( .A(n1226), .B(G140), .ZN(n1343) );
INV_X1 U1056 ( .A(G146), .ZN(n1226) );
XOR2_X1 U1057 ( .A(n1345), .B(n1346), .Z(n1341) );
XNOR2_X1 U1058 ( .A(n1347), .B(G104), .ZN(n1346) );
INV_X1 U1059 ( .A(G113), .ZN(n1347) );
NAND2_X1 U1060 ( .A1(KEYINPUT56), .A2(n1348), .ZN(n1345) );
XNOR2_X1 U1061 ( .A(G131), .B(n1349), .ZN(n1348) );
NAND2_X1 U1062 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NAND2_X1 U1063 ( .A1(n1352), .A2(n1334), .ZN(n1351) );
XOR2_X1 U1064 ( .A(n1353), .B(KEYINPUT19), .Z(n1350) );
OR2_X1 U1065 ( .A1(n1334), .A2(n1352), .ZN(n1353) );
NAND3_X1 U1066 ( .A1(n1327), .A2(n1057), .A3(G214), .ZN(n1352) );
NOR2_X1 U1067 ( .A1(n1105), .A2(n1261), .ZN(n1207) );
INV_X1 U1068 ( .A(n1246), .ZN(n1261) );
NAND2_X1 U1069 ( .A1(n1354), .A2(n1102), .ZN(n1246) );
NAND3_X1 U1070 ( .A1(n1355), .A2(n1356), .A3(G217), .ZN(n1102) );
NAND2_X1 U1071 ( .A1(n1145), .A2(n1272), .ZN(n1356) );
XOR2_X1 U1072 ( .A(KEYINPUT61), .B(n1101), .Z(n1354) );
AND3_X1 U1073 ( .A1(n1357), .A2(n1272), .A3(n1145), .ZN(n1101) );
XNOR2_X1 U1074 ( .A(n1358), .B(n1359), .ZN(n1145) );
XOR2_X1 U1075 ( .A(n1277), .B(n1360), .Z(n1359) );
XOR2_X1 U1076 ( .A(G110), .B(G140), .Z(n1277) );
XOR2_X1 U1077 ( .A(n1361), .B(n1362), .Z(n1358) );
NOR2_X1 U1078 ( .A1(G125), .A2(KEYINPUT55), .ZN(n1362) );
XNOR2_X1 U1079 ( .A(G119), .B(n1363), .ZN(n1361) );
NOR3_X1 U1080 ( .A1(n1364), .A2(KEYINPUT18), .A3(n1365), .ZN(n1363) );
NOR3_X1 U1081 ( .A1(n1366), .A2(n1339), .A3(n1367), .ZN(n1365) );
XNOR2_X1 U1082 ( .A(G137), .B(n1368), .ZN(n1366) );
XNOR2_X1 U1083 ( .A(KEYINPUT5), .B(KEYINPUT41), .ZN(n1368) );
NOR2_X1 U1084 ( .A1(n1369), .A2(n1127), .ZN(n1364) );
NOR2_X1 U1085 ( .A1(n1339), .A2(n1367), .ZN(n1369) );
INV_X1 U1086 ( .A(G221), .ZN(n1367) );
NAND2_X1 U1087 ( .A1(G234), .A2(n1057), .ZN(n1339) );
NAND2_X1 U1088 ( .A1(G217), .A2(n1355), .ZN(n1357) );
XNOR2_X1 U1089 ( .A(KEYINPUT45), .B(n1283), .ZN(n1355) );
NAND2_X1 U1090 ( .A1(G234), .A2(n1272), .ZN(n1283) );
XOR2_X1 U1091 ( .A(n1370), .B(n1171), .Z(n1105) );
INV_X1 U1092 ( .A(G472), .ZN(n1171) );
NAND2_X1 U1093 ( .A1(n1371), .A2(n1272), .ZN(n1370) );
INV_X1 U1094 ( .A(G902), .ZN(n1272) );
XOR2_X1 U1095 ( .A(n1372), .B(n1373), .Z(n1371) );
XOR2_X1 U1096 ( .A(KEYINPUT63), .B(KEYINPUT13), .Z(n1373) );
XOR2_X1 U1097 ( .A(n1169), .B(n1168), .Z(n1372) );
XNOR2_X1 U1098 ( .A(n1374), .B(G101), .ZN(n1168) );
NAND3_X1 U1099 ( .A1(n1327), .A2(n1057), .A3(G210), .ZN(n1374) );
INV_X1 U1100 ( .A(G953), .ZN(n1057) );
INV_X1 U1101 ( .A(G237), .ZN(n1327) );
XOR2_X1 U1102 ( .A(n1280), .B(n1375), .Z(n1169) );
NOR2_X1 U1103 ( .A1(n1300), .A2(n1304), .ZN(n1375) );
NAND2_X1 U1104 ( .A1(n1376), .A2(n1377), .ZN(n1304) );
NAND2_X1 U1105 ( .A1(n1378), .A2(G119), .ZN(n1377) );
XNOR2_X1 U1106 ( .A(G116), .B(n1303), .ZN(n1378) );
NAND3_X1 U1107 ( .A1(n1303), .A2(n1257), .A3(n1256), .ZN(n1376) );
INV_X1 U1108 ( .A(G119), .ZN(n1256) );
NOR3_X1 U1109 ( .A1(n1257), .A2(G119), .A3(n1303), .ZN(n1300) );
XOR2_X1 U1110 ( .A(G113), .B(KEYINPUT47), .Z(n1303) );
INV_X1 U1111 ( .A(G116), .ZN(n1257) );
XOR2_X1 U1112 ( .A(n1379), .B(n1380), .Z(n1280) );
XNOR2_X1 U1113 ( .A(KEYINPUT58), .B(n1127), .ZN(n1380) );
INV_X1 U1114 ( .A(G137), .ZN(n1127) );
XNOR2_X1 U1115 ( .A(n1126), .B(n1130), .ZN(n1379) );
INV_X1 U1116 ( .A(G131), .ZN(n1130) );
XNOR2_X1 U1117 ( .A(G134), .B(n1222), .ZN(n1126) );
XNOR2_X1 U1118 ( .A(n1334), .B(n1360), .ZN(n1222) );
XOR2_X1 U1119 ( .A(G128), .B(G146), .Z(n1360) );
INV_X1 U1120 ( .A(G143), .ZN(n1334) );
endmodule


