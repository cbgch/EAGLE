//Key = 1101011010111000000010100110100101010000100000100011100000111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;

XNOR2_X1 U710 ( .A(G107), .B(n980), .ZN(G9) );
NOR2_X1 U711 ( .A1(n981), .A2(n982), .ZN(G75) );
NOR4_X1 U712 ( .A1(G953), .A2(n983), .A3(n984), .A4(n985), .ZN(n982) );
NOR2_X1 U713 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U714 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR2_X1 U715 ( .A1(n990), .A2(n991), .ZN(n989) );
INV_X1 U716 ( .A(n992), .ZN(n991) );
NOR2_X1 U717 ( .A1(n993), .A2(n994), .ZN(n990) );
NOR2_X1 U718 ( .A1(n995), .A2(n996), .ZN(n994) );
NOR2_X1 U719 ( .A1(n997), .A2(n998), .ZN(n995) );
NOR2_X1 U720 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR2_X1 U721 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U722 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U723 ( .A1(n1005), .A2(n1006), .ZN(n997) );
NOR2_X1 U724 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
AND2_X1 U725 ( .A1(n1009), .A2(n1010), .ZN(n1007) );
NOR3_X1 U726 ( .A1(n1006), .A2(n1011), .A3(n1000), .ZN(n993) );
NOR2_X1 U727 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U728 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NOR4_X1 U729 ( .A1(n1016), .A2(n1000), .A3(n1006), .A4(n996), .ZN(n988) );
INV_X1 U730 ( .A(n1017), .ZN(n996) );
INV_X1 U731 ( .A(n1018), .ZN(n1000) );
NOR2_X1 U732 ( .A1(n1019), .A2(n1020), .ZN(n1016) );
NOR3_X1 U733 ( .A1(n983), .A2(G953), .A3(G952), .ZN(n981) );
AND4_X1 U734 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n1024), .ZN(n983) );
NOR3_X1 U735 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
XNOR2_X1 U736 ( .A(KEYINPUT45), .B(n1028), .ZN(n1027) );
NAND4_X1 U737 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1025) );
NAND2_X1 U738 ( .A1(KEYINPUT19), .A2(n1033), .ZN(n1032) );
NAND2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1031) );
INV_X1 U740 ( .A(KEYINPUT19), .ZN(n1035) );
NAND2_X1 U741 ( .A1(n1036), .A2(n1004), .ZN(n1034) );
NAND2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1030) );
NAND2_X1 U743 ( .A1(n1039), .A2(n1040), .ZN(n1029) );
INV_X1 U744 ( .A(n1038), .ZN(n1040) );
XOR2_X1 U745 ( .A(KEYINPUT26), .B(n1037), .Z(n1039) );
AND3_X1 U746 ( .A1(n1041), .A2(n1042), .A3(n1015), .ZN(n1023) );
NAND2_X1 U747 ( .A1(G475), .A2(n1043), .ZN(n1022) );
XOR2_X1 U748 ( .A(n1044), .B(n1045), .Z(G72) );
NOR2_X1 U749 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U750 ( .A1(G227), .A2(n1048), .ZN(n1046) );
NOR3_X1 U751 ( .A1(KEYINPUT4), .A2(n1049), .A3(n1050), .ZN(n1044) );
AND2_X1 U752 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR3_X1 U753 ( .A1(n1052), .A2(n1047), .A3(n1051), .ZN(n1049) );
NAND2_X1 U754 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
OR2_X1 U755 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U756 ( .A(n1057), .B(KEYINPUT48), .Z(n1053) );
NAND2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1057) );
XNOR2_X1 U758 ( .A(n1058), .B(n1059), .ZN(n1055) );
XOR2_X1 U759 ( .A(n1060), .B(n1061), .Z(n1059) );
XNOR2_X1 U760 ( .A(KEYINPUT14), .B(n1062), .ZN(n1058) );
NOR2_X1 U761 ( .A1(KEYINPUT36), .A2(n1063), .ZN(n1062) );
XOR2_X1 U762 ( .A(G134), .B(n1064), .Z(n1063) );
NOR2_X1 U763 ( .A1(G953), .A2(n1065), .ZN(n1052) );
XOR2_X1 U764 ( .A(n1066), .B(n1067), .Z(G69) );
XOR2_X1 U765 ( .A(n1068), .B(n1069), .Z(n1067) );
NAND2_X1 U766 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U767 ( .A(n1072), .B(n1073), .Z(n1070) );
XNOR2_X1 U768 ( .A(KEYINPUT28), .B(n1074), .ZN(n1072) );
NOR2_X1 U769 ( .A1(n1075), .A2(KEYINPUT13), .ZN(n1074) );
NAND2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1068) );
NAND3_X1 U771 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
XOR2_X1 U772 ( .A(n1081), .B(KEYINPUT37), .Z(n1080) );
XOR2_X1 U773 ( .A(KEYINPUT5), .B(G953), .Z(n1076) );
NAND3_X1 U774 ( .A1(n1082), .A2(n1071), .A3(KEYINPUT31), .ZN(n1066) );
INV_X1 U775 ( .A(n1083), .ZN(n1071) );
OR2_X1 U776 ( .A1(n1048), .A2(G224), .ZN(n1082) );
NOR2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(G66) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
XOR2_X1 U779 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U780 ( .A1(KEYINPUT9), .A2(n1090), .ZN(n1089) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1037), .ZN(n1088) );
AND2_X1 U782 ( .A1(n1090), .A2(KEYINPUT9), .ZN(n1086) );
NOR2_X1 U783 ( .A1(n1084), .A2(n1092), .ZN(G63) );
XOR2_X1 U784 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND3_X1 U785 ( .A1(n1091), .A2(G478), .A3(KEYINPUT58), .ZN(n1093) );
NOR2_X1 U786 ( .A1(n1084), .A2(n1095), .ZN(G60) );
XOR2_X1 U787 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U788 ( .A1(n1091), .A2(G475), .ZN(n1096) );
XNOR2_X1 U789 ( .A(G104), .B(n1098), .ZN(G6) );
NOR2_X1 U790 ( .A1(n1084), .A2(n1099), .ZN(G57) );
XOR2_X1 U791 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U792 ( .A(n1102), .B(n1103), .Z(n1101) );
XNOR2_X1 U793 ( .A(n1104), .B(n1105), .ZN(n1103) );
NOR2_X1 U794 ( .A1(KEYINPUT2), .A2(n1106), .ZN(n1105) );
NOR2_X1 U795 ( .A1(KEYINPUT29), .A2(n1107), .ZN(n1104) );
XOR2_X1 U796 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U797 ( .A(n1110), .B(KEYINPUT30), .Z(n1109) );
NAND2_X1 U798 ( .A1(n1091), .A2(G472), .ZN(n1102) );
XOR2_X1 U799 ( .A(n1111), .B(n1112), .Z(n1100) );
NOR2_X1 U800 ( .A1(n1084), .A2(n1113), .ZN(G54) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U802 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U803 ( .A(G110), .B(G140), .ZN(n1117) );
NAND2_X1 U804 ( .A1(n1091), .A2(G469), .ZN(n1116) );
INV_X1 U805 ( .A(n1118), .ZN(n1091) );
XNOR2_X1 U806 ( .A(n1119), .B(n1120), .ZN(n1114) );
NOR2_X1 U807 ( .A1(n1084), .A2(n1121), .ZN(G51) );
XOR2_X1 U808 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U810 ( .A1(n1126), .A2(KEYINPUT53), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1118), .ZN(n1126) );
NAND2_X1 U812 ( .A1(G902), .A2(n985), .ZN(n1118) );
NAND3_X1 U813 ( .A1(n1078), .A2(n1128), .A3(n1065), .ZN(n985) );
AND4_X1 U814 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1065) );
NOR3_X1 U815 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
INV_X1 U816 ( .A(n1136), .ZN(n1135) );
NOR2_X1 U817 ( .A1(n1137), .A2(n1033), .ZN(n1133) );
NOR3_X1 U818 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1137) );
XOR2_X1 U819 ( .A(KEYINPUT15), .B(n1141), .Z(n1138) );
XOR2_X1 U820 ( .A(KEYINPUT43), .B(n1142), .Z(n1128) );
AND2_X1 U821 ( .A1(n1081), .A2(n1079), .ZN(n1142) );
AND3_X1 U822 ( .A1(n1143), .A2(n980), .A3(n1098), .ZN(n1079) );
NAND3_X1 U823 ( .A1(n1018), .A2(n1144), .A3(n1020), .ZN(n1098) );
NAND3_X1 U824 ( .A1(n1018), .A2(n1144), .A3(n1019), .ZN(n980) );
AND4_X1 U825 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1078) );
XOR2_X1 U826 ( .A(n1149), .B(n1150), .Z(n1122) );
NOR2_X1 U827 ( .A1(KEYINPUT18), .A2(n1151), .ZN(n1150) );
XOR2_X1 U828 ( .A(G125), .B(n1152), .Z(n1151) );
NOR2_X1 U829 ( .A1(KEYINPUT41), .A2(n1111), .ZN(n1152) );
NOR2_X1 U830 ( .A1(n1048), .A2(G952), .ZN(n1084) );
XOR2_X1 U831 ( .A(G146), .B(n1153), .Z(G48) );
NOR2_X1 U832 ( .A1(n1033), .A2(n1154), .ZN(n1153) );
XOR2_X1 U833 ( .A(KEYINPUT12), .B(n1141), .Z(n1154) );
AND2_X1 U834 ( .A1(n1155), .A2(n1020), .ZN(n1141) );
XOR2_X1 U835 ( .A(n1156), .B(n1136), .Z(G45) );
NAND4_X1 U836 ( .A1(n1157), .A2(n1002), .A3(n1026), .A4(n1158), .ZN(n1136) );
XNOR2_X1 U837 ( .A(G140), .B(n1129), .ZN(G42) );
NAND3_X1 U838 ( .A1(n1159), .A2(n1013), .A3(n1160), .ZN(n1129) );
XOR2_X1 U839 ( .A(G137), .B(n1134), .Z(G39) );
AND3_X1 U840 ( .A1(n1155), .A2(n1159), .A3(n992), .ZN(n1134) );
XNOR2_X1 U841 ( .A(G134), .B(n1131), .ZN(G36) );
NAND3_X1 U842 ( .A1(n1157), .A2(n1019), .A3(n1159), .ZN(n1131) );
XNOR2_X1 U843 ( .A(G131), .B(n1130), .ZN(G33) );
NAND3_X1 U844 ( .A1(n1159), .A2(n1157), .A3(n1020), .ZN(n1130) );
AND3_X1 U845 ( .A1(n1013), .A2(n1161), .A3(n1008), .ZN(n1157) );
INV_X1 U846 ( .A(n1006), .ZN(n1159) );
NAND2_X1 U847 ( .A1(n1162), .A2(n1036), .ZN(n1006) );
XOR2_X1 U848 ( .A(n1004), .B(KEYINPUT16), .Z(n1162) );
NAND3_X1 U849 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(G30) );
NAND2_X1 U850 ( .A1(KEYINPUT63), .A2(n1166), .ZN(n1165) );
OR3_X1 U851 ( .A1(n1166), .A2(KEYINPUT63), .A3(G128), .ZN(n1164) );
NAND2_X1 U852 ( .A1(G128), .A2(n1167), .ZN(n1163) );
NAND2_X1 U853 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
INV_X1 U854 ( .A(KEYINPUT63), .ZN(n1169) );
XNOR2_X1 U855 ( .A(KEYINPUT24), .B(n1166), .ZN(n1168) );
NAND2_X1 U856 ( .A1(n1139), .A2(n1170), .ZN(n1166) );
XOR2_X1 U857 ( .A(KEYINPUT44), .B(n1002), .Z(n1170) );
AND2_X1 U858 ( .A1(n1155), .A2(n1019), .ZN(n1139) );
AND4_X1 U859 ( .A1(n1171), .A2(n1013), .A3(n1009), .A4(n1161), .ZN(n1155) );
XOR2_X1 U860 ( .A(n1110), .B(n1143), .Z(G3) );
NAND3_X1 U861 ( .A1(n1008), .A2(n1144), .A3(n992), .ZN(n1143) );
XOR2_X1 U862 ( .A(n1172), .B(n1173), .Z(G27) );
NAND2_X1 U863 ( .A1(n1140), .A2(n1174), .ZN(n1173) );
XOR2_X1 U864 ( .A(KEYINPUT39), .B(n1002), .Z(n1174) );
AND2_X1 U865 ( .A1(n1017), .A2(n1160), .ZN(n1140) );
AND4_X1 U866 ( .A1(n1020), .A2(n1010), .A3(n1009), .A4(n1161), .ZN(n1160) );
NAND2_X1 U867 ( .A1(n1175), .A2(n1176), .ZN(n1161) );
NAND3_X1 U868 ( .A1(G902), .A2(n1177), .A3(n1047), .ZN(n1176) );
NOR2_X1 U869 ( .A1(G900), .A2(n1048), .ZN(n1047) );
XNOR2_X1 U870 ( .A(KEYINPUT22), .B(n987), .ZN(n1175) );
XNOR2_X1 U871 ( .A(G122), .B(n1178), .ZN(G24) );
NAND2_X1 U872 ( .A1(KEYINPUT6), .A2(n1179), .ZN(n1178) );
INV_X1 U873 ( .A(n1145), .ZN(n1179) );
NAND4_X1 U874 ( .A1(n1180), .A2(n1018), .A3(n1026), .A4(n1158), .ZN(n1145) );
NOR2_X1 U875 ( .A1(n1009), .A2(n1171), .ZN(n1018) );
XOR2_X1 U876 ( .A(n1146), .B(n1181), .Z(G21) );
XOR2_X1 U877 ( .A(KEYINPUT25), .B(G119), .Z(n1181) );
NAND4_X1 U878 ( .A1(n1180), .A2(n992), .A3(n1171), .A4(n1009), .ZN(n1146) );
XOR2_X1 U879 ( .A(n1182), .B(n1147), .Z(G18) );
NAND3_X1 U880 ( .A1(n1008), .A2(n1019), .A3(n1180), .ZN(n1147) );
NOR2_X1 U881 ( .A1(n1158), .A2(n1183), .ZN(n1019) );
XNOR2_X1 U882 ( .A(G113), .B(n1148), .ZN(G15) );
NAND3_X1 U883 ( .A1(n1020), .A2(n1008), .A3(n1180), .ZN(n1148) );
AND2_X1 U884 ( .A1(n1017), .A2(n1184), .ZN(n1180) );
NOR2_X1 U885 ( .A1(n1014), .A2(n1185), .ZN(n1017) );
INV_X1 U886 ( .A(n1015), .ZN(n1185) );
NOR2_X1 U887 ( .A1(n1010), .A2(n1009), .ZN(n1008) );
AND2_X1 U888 ( .A1(n1183), .A2(n1158), .ZN(n1020) );
XNOR2_X1 U889 ( .A(G110), .B(n1081), .ZN(G12) );
NAND4_X1 U890 ( .A1(n992), .A2(n1144), .A3(n1010), .A4(n1009), .ZN(n1081) );
XNOR2_X1 U891 ( .A(n1038), .B(n1037), .ZN(n1009) );
AND2_X1 U892 ( .A1(G217), .A2(n1186), .ZN(n1037) );
NAND2_X1 U893 ( .A1(n1090), .A2(n1187), .ZN(n1038) );
XNOR2_X1 U894 ( .A(n1188), .B(n1189), .ZN(n1090) );
XOR2_X1 U895 ( .A(G110), .B(n1190), .Z(n1189) );
XOR2_X1 U896 ( .A(G137), .B(G119), .Z(n1190) );
XOR2_X1 U897 ( .A(n1191), .B(n1056), .Z(n1188) );
XOR2_X1 U898 ( .A(n1192), .B(n1193), .Z(n1191) );
NAND2_X1 U899 ( .A1(G221), .A2(n1194), .ZN(n1192) );
INV_X1 U900 ( .A(n1171), .ZN(n1010) );
XOR2_X1 U901 ( .A(n1021), .B(KEYINPUT33), .Z(n1171) );
XNOR2_X1 U902 ( .A(G472), .B(n1195), .ZN(n1021) );
NOR2_X1 U903 ( .A1(G902), .A2(n1196), .ZN(n1195) );
XOR2_X1 U904 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U905 ( .A(n1112), .B(n1108), .Z(n1198) );
NAND3_X1 U906 ( .A1(n1199), .A2(n1048), .A3(n1200), .ZN(n1108) );
XOR2_X1 U907 ( .A(KEYINPUT32), .B(G210), .Z(n1200) );
XNOR2_X1 U908 ( .A(n1201), .B(n1202), .ZN(n1112) );
XOR2_X1 U909 ( .A(G116), .B(G113), .Z(n1202) );
NAND2_X1 U910 ( .A1(KEYINPUT35), .A2(G119), .ZN(n1201) );
XOR2_X1 U911 ( .A(n1203), .B(n1204), .Z(n1197) );
NOR2_X1 U912 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U913 ( .A(n1207), .B(KEYINPUT8), .Z(n1206) );
NAND2_X1 U914 ( .A1(n1106), .A2(n1208), .ZN(n1207) );
NOR2_X1 U915 ( .A1(n1106), .A2(n1208), .ZN(n1205) );
XNOR2_X1 U916 ( .A(KEYINPUT10), .B(n1209), .ZN(n1203) );
NOR2_X1 U917 ( .A1(KEYINPUT61), .A2(n1110), .ZN(n1209) );
AND2_X1 U918 ( .A1(n1184), .A2(n1013), .ZN(n1144) );
AND2_X1 U919 ( .A1(n1015), .A2(n1014), .ZN(n1013) );
NAND2_X1 U920 ( .A1(n1041), .A2(n1028), .ZN(n1014) );
NAND3_X1 U921 ( .A1(n1210), .A2(n1187), .A3(n1211), .ZN(n1028) );
XOR2_X1 U922 ( .A(KEYINPUT59), .B(G469), .Z(n1210) );
NAND2_X1 U923 ( .A1(n1212), .A2(n1213), .ZN(n1041) );
NAND2_X1 U924 ( .A1(n1211), .A2(n1187), .ZN(n1213) );
XOR2_X1 U925 ( .A(n1214), .B(n1215), .Z(n1211) );
XNOR2_X1 U926 ( .A(n1216), .B(n1217), .ZN(n1215) );
NOR2_X1 U927 ( .A1(KEYINPUT49), .A2(n1119), .ZN(n1217) );
XOR2_X1 U928 ( .A(n1218), .B(n1061), .Z(n1119) );
XNOR2_X1 U929 ( .A(n1193), .B(n1219), .ZN(n1061) );
NOR2_X1 U930 ( .A1(KEYINPUT56), .A2(n1220), .ZN(n1219) );
XOR2_X1 U931 ( .A(n1221), .B(n1110), .Z(n1218) );
INV_X1 U932 ( .A(G101), .ZN(n1110) );
XNOR2_X1 U933 ( .A(G110), .B(KEYINPUT54), .ZN(n1216) );
XOR2_X1 U934 ( .A(n1222), .B(n1120), .Z(n1214) );
XNOR2_X1 U935 ( .A(n1106), .B(n1223), .ZN(n1120) );
AND2_X1 U936 ( .A1(n1048), .A2(G227), .ZN(n1223) );
NAND2_X1 U937 ( .A1(n1224), .A2(n1225), .ZN(n1106) );
NAND2_X1 U938 ( .A1(n1226), .A2(n1064), .ZN(n1225) );
INV_X1 U939 ( .A(G137), .ZN(n1064) );
XOR2_X1 U940 ( .A(n1227), .B(KEYINPUT1), .Z(n1226) );
NAND2_X1 U941 ( .A1(n1228), .A2(G137), .ZN(n1224) );
XOR2_X1 U942 ( .A(KEYINPUT20), .B(n1229), .Z(n1228) );
INV_X1 U943 ( .A(n1227), .ZN(n1229) );
XOR2_X1 U944 ( .A(n1230), .B(n1231), .Z(n1227) );
INV_X1 U945 ( .A(n1060), .ZN(n1231) );
XNOR2_X1 U946 ( .A(G131), .B(KEYINPUT52), .ZN(n1060) );
XNOR2_X1 U947 ( .A(G134), .B(KEYINPUT21), .ZN(n1230) );
NAND2_X1 U948 ( .A1(KEYINPUT51), .A2(G140), .ZN(n1222) );
XNOR2_X1 U949 ( .A(G469), .B(KEYINPUT59), .ZN(n1212) );
NAND2_X1 U950 ( .A1(n1232), .A2(G221), .ZN(n1015) );
XOR2_X1 U951 ( .A(n1186), .B(KEYINPUT34), .Z(n1232) );
NAND2_X1 U952 ( .A1(G234), .A2(n1187), .ZN(n1186) );
AND2_X1 U953 ( .A1(n1002), .A2(n1233), .ZN(n1184) );
NAND2_X1 U954 ( .A1(n987), .A2(n1234), .ZN(n1233) );
NAND3_X1 U955 ( .A1(n1083), .A2(n1177), .A3(G902), .ZN(n1234) );
NOR2_X1 U956 ( .A1(G898), .A2(n1048), .ZN(n1083) );
NAND3_X1 U957 ( .A1(n1177), .A2(n1048), .A3(G952), .ZN(n987) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1177) );
INV_X1 U959 ( .A(n1033), .ZN(n1002) );
NAND2_X1 U960 ( .A1(n1003), .A2(n1004), .ZN(n1033) );
NAND2_X1 U961 ( .A1(G214), .A2(n1235), .ZN(n1004) );
INV_X1 U962 ( .A(n1036), .ZN(n1003) );
XNOR2_X1 U963 ( .A(n1236), .B(n1127), .ZN(n1036) );
NAND2_X1 U964 ( .A1(G210), .A2(n1235), .ZN(n1127) );
NAND2_X1 U965 ( .A1(n1199), .A2(n1187), .ZN(n1235) );
NAND2_X1 U966 ( .A1(n1237), .A2(n1187), .ZN(n1236) );
XOR2_X1 U967 ( .A(n1124), .B(n1238), .Z(n1237) );
XOR2_X1 U968 ( .A(n1149), .B(n1239), .Z(n1238) );
NAND3_X1 U969 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
NAND2_X1 U970 ( .A1(KEYINPUT17), .A2(G125), .ZN(n1242) );
NAND3_X1 U971 ( .A1(n1172), .A2(n1243), .A3(n1111), .ZN(n1241) );
INV_X1 U972 ( .A(G125), .ZN(n1172) );
NAND2_X1 U973 ( .A1(n1208), .A2(n1244), .ZN(n1240) );
NAND2_X1 U974 ( .A1(n1245), .A2(n1243), .ZN(n1244) );
INV_X1 U975 ( .A(KEYINPUT17), .ZN(n1243) );
XOR2_X1 U976 ( .A(KEYINPUT46), .B(G125), .Z(n1245) );
INV_X1 U977 ( .A(n1111), .ZN(n1208) );
XNOR2_X1 U978 ( .A(n1220), .B(n1246), .ZN(n1111) );
XOR2_X1 U979 ( .A(KEYINPUT38), .B(n1193), .Z(n1246) );
XOR2_X1 U980 ( .A(G146), .B(G128), .Z(n1193) );
XNOR2_X1 U981 ( .A(n1156), .B(KEYINPUT40), .ZN(n1220) );
NAND2_X1 U982 ( .A1(G224), .A2(n1048), .ZN(n1149) );
XNOR2_X1 U983 ( .A(n1075), .B(n1073), .ZN(n1124) );
XOR2_X1 U984 ( .A(G110), .B(G122), .Z(n1073) );
AND3_X1 U985 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1075) );
OR3_X1 U986 ( .A1(n1250), .A2(G119), .A3(n1182), .ZN(n1249) );
NAND3_X1 U987 ( .A1(n1250), .A2(n1182), .A3(n1251), .ZN(n1248) );
INV_X1 U988 ( .A(G119), .ZN(n1251) );
NAND2_X1 U989 ( .A1(n1252), .A2(G119), .ZN(n1247) );
XOR2_X1 U990 ( .A(n1182), .B(n1250), .Z(n1252) );
XOR2_X1 U991 ( .A(n1253), .B(n1254), .Z(n1250) );
XOR2_X1 U992 ( .A(KEYINPUT23), .B(G113), .Z(n1254) );
XOR2_X1 U993 ( .A(n1255), .B(G101), .Z(n1253) );
NAND2_X1 U994 ( .A1(KEYINPUT62), .A2(n1221), .ZN(n1255) );
XOR2_X1 U995 ( .A(G107), .B(n1256), .Z(n1221) );
INV_X1 U996 ( .A(G116), .ZN(n1182) );
NOR2_X1 U997 ( .A1(n1026), .A2(n1158), .ZN(n992) );
NAND3_X1 U998 ( .A1(n1257), .A2(n1258), .A3(n1042), .ZN(n1158) );
OR2_X1 U999 ( .A1(n1043), .A2(G475), .ZN(n1042) );
OR2_X1 U1000 ( .A1(n1259), .A2(G475), .ZN(n1258) );
NAND3_X1 U1001 ( .A1(n1043), .A2(n1259), .A3(G475), .ZN(n1257) );
INV_X1 U1002 ( .A(KEYINPUT27), .ZN(n1259) );
NAND2_X1 U1003 ( .A1(n1097), .A2(n1187), .ZN(n1043) );
XNOR2_X1 U1004 ( .A(n1260), .B(n1261), .ZN(n1097) );
XNOR2_X1 U1005 ( .A(n1056), .B(n1262), .ZN(n1261) );
XNOR2_X1 U1006 ( .A(n1263), .B(n1264), .ZN(n1262) );
NAND2_X1 U1007 ( .A1(n1265), .A2(KEYINPUT0), .ZN(n1264) );
XOR2_X1 U1008 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U1009 ( .A(KEYINPUT42), .B(G122), .Z(n1267) );
XNOR2_X1 U1010 ( .A(G113), .B(n1256), .ZN(n1266) );
XOR2_X1 U1011 ( .A(G104), .B(KEYINPUT57), .Z(n1256) );
NAND2_X1 U1012 ( .A1(KEYINPUT11), .A2(n1268), .ZN(n1263) );
XOR2_X1 U1013 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U1014 ( .A(n1156), .B(KEYINPUT3), .Z(n1270) );
INV_X1 U1015 ( .A(G143), .ZN(n1156) );
NAND4_X1 U1016 ( .A1(KEYINPUT50), .A2(G214), .A3(n1199), .A4(n1048), .ZN(n1269) );
INV_X1 U1017 ( .A(G237), .ZN(n1199) );
XOR2_X1 U1018 ( .A(G140), .B(G125), .Z(n1056) );
XNOR2_X1 U1019 ( .A(G131), .B(n1271), .ZN(n1260) );
XOR2_X1 U1020 ( .A(KEYINPUT7), .B(G146), .Z(n1271) );
INV_X1 U1021 ( .A(n1183), .ZN(n1026) );
XOR2_X1 U1022 ( .A(n1272), .B(G478), .Z(n1183) );
NAND2_X1 U1023 ( .A1(n1094), .A2(n1187), .ZN(n1272) );
INV_X1 U1024 ( .A(G902), .ZN(n1187) );
XNOR2_X1 U1025 ( .A(n1273), .B(n1274), .ZN(n1094) );
XOR2_X1 U1026 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U1027 ( .A(G128), .B(n1277), .Z(n1276) );
NOR2_X1 U1028 ( .A1(KEYINPUT55), .A2(n1278), .ZN(n1277) );
XOR2_X1 U1029 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U1030 ( .A(G116), .B(G107), .Z(n1280) );
XOR2_X1 U1031 ( .A(KEYINPUT47), .B(G122), .Z(n1279) );
AND2_X1 U1032 ( .A1(n1194), .A2(G217), .ZN(n1275) );
AND2_X1 U1033 ( .A1(G234), .A2(n1048), .ZN(n1194) );
INV_X1 U1034 ( .A(G953), .ZN(n1048) );
XNOR2_X1 U1035 ( .A(G134), .B(n1281), .ZN(n1273) );
XOR2_X1 U1036 ( .A(KEYINPUT60), .B(G143), .Z(n1281) );
endmodule


