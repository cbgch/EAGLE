//Key = 0111110110101011100011010110100000011110100111100010100010001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;

XNOR2_X1 U766 ( .A(G107), .B(n1064), .ZN(G9) );
NAND3_X1 U767 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
XNOR2_X1 U768 ( .A(KEYINPUT62), .B(n1068), .ZN(n1066) );
NOR2_X1 U769 ( .A1(n1069), .A2(n1070), .ZN(G75) );
NOR4_X1 U770 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NOR2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
NOR2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NOR3_X1 U773 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NOR3_X1 U774 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1080) );
NOR2_X1 U775 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U776 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
INV_X1 U778 ( .A(n1091), .ZN(n1083) );
NOR2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1082) );
NOR3_X1 U780 ( .A1(n1092), .A2(n1094), .A3(n1086), .ZN(n1077) );
NOR3_X1 U781 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
NOR2_X1 U782 ( .A1(n1098), .A2(n1081), .ZN(n1097) );
INV_X1 U783 ( .A(n1099), .ZN(n1081) );
NOR2_X1 U784 ( .A1(n1067), .A2(n1100), .ZN(n1098) );
NOR3_X1 U785 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1096) );
XNOR2_X1 U786 ( .A(KEYINPUT40), .B(n1079), .ZN(n1101) );
NOR2_X1 U787 ( .A1(n1104), .A2(n1079), .ZN(n1095) );
NAND3_X1 U788 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1071) );
NOR3_X1 U789 ( .A1(n1108), .A2(G952), .A3(n1073), .ZN(n1069) );
AND4_X1 U790 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1073) );
NOR4_X1 U791 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1112) );
NOR2_X1 U792 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XOR2_X1 U793 ( .A(KEYINPUT44), .B(G475), .Z(n1118) );
INV_X1 U794 ( .A(n1119), .ZN(n1117) );
NOR2_X1 U795 ( .A1(n1120), .A2(n1121), .ZN(n1111) );
XNOR2_X1 U796 ( .A(G469), .B(n1122), .ZN(n1121) );
XNOR2_X1 U797 ( .A(n1123), .B(n1124), .ZN(n1120) );
XOR2_X1 U798 ( .A(n1125), .B(n1126), .Z(G72) );
NOR3_X1 U799 ( .A1(n1127), .A2(KEYINPUT53), .A3(n1128), .ZN(n1126) );
NOR2_X1 U800 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U801 ( .A1(n1131), .A2(n1132), .ZN(n1125) );
NAND2_X1 U802 ( .A1(n1133), .A2(n1127), .ZN(n1132) );
XNOR2_X1 U803 ( .A(n1134), .B(n1107), .ZN(n1133) );
NAND3_X1 U804 ( .A1(G900), .A2(n1134), .A3(G953), .ZN(n1131) );
XNOR2_X1 U805 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U806 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U807 ( .A1(KEYINPUT63), .A2(n1139), .ZN(n1137) );
INV_X1 U808 ( .A(n1140), .ZN(n1139) );
XNOR2_X1 U809 ( .A(n1141), .B(n1142), .ZN(n1135) );
NAND2_X1 U810 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
INV_X1 U811 ( .A(n1145), .ZN(n1144) );
XOR2_X1 U812 ( .A(n1146), .B(KEYINPUT18), .Z(n1143) );
NAND2_X1 U813 ( .A1(G140), .A2(n1147), .ZN(n1146) );
XNOR2_X1 U814 ( .A(KEYINPUT3), .B(n1148), .ZN(n1147) );
XOR2_X1 U815 ( .A(n1149), .B(n1150), .Z(G69) );
NOR2_X1 U816 ( .A1(n1151), .A2(n1127), .ZN(n1150) );
NOR2_X1 U817 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U818 ( .A1(n1154), .A2(n1155), .ZN(n1149) );
NAND2_X1 U819 ( .A1(n1156), .A2(n1127), .ZN(n1155) );
XOR2_X1 U820 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U821 ( .A1(n1159), .A2(n1106), .ZN(n1157) );
XNOR2_X1 U822 ( .A(n1074), .B(KEYINPUT30), .ZN(n1159) );
INV_X1 U823 ( .A(n1160), .ZN(n1074) );
NAND3_X1 U824 ( .A1(n1158), .A2(G898), .A3(G953), .ZN(n1154) );
AND2_X1 U825 ( .A1(KEYINPUT36), .A2(n1161), .ZN(n1158) );
NOR2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(G66) );
XNOR2_X1 U827 ( .A(n1164), .B(n1165), .ZN(n1163) );
NOR2_X1 U828 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NOR2_X1 U829 ( .A1(n1168), .A2(n1169), .ZN(G63) );
XOR2_X1 U830 ( .A(KEYINPUT49), .B(n1162), .Z(n1169) );
XOR2_X1 U831 ( .A(n1170), .B(n1171), .Z(n1168) );
NOR2_X1 U832 ( .A1(KEYINPUT39), .A2(n1172), .ZN(n1171) );
XOR2_X1 U833 ( .A(n1173), .B(n1174), .Z(n1172) );
NAND2_X1 U834 ( .A1(n1175), .A2(G478), .ZN(n1170) );
NOR2_X1 U835 ( .A1(n1162), .A2(n1176), .ZN(G60) );
XOR2_X1 U836 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND3_X1 U837 ( .A1(n1175), .A2(G475), .A3(KEYINPUT37), .ZN(n1177) );
XNOR2_X1 U838 ( .A(n1179), .B(n1180), .ZN(G6) );
NAND2_X1 U839 ( .A1(KEYINPUT35), .A2(G104), .ZN(n1180) );
NOR2_X1 U840 ( .A1(n1162), .A2(n1181), .ZN(G57) );
XOR2_X1 U841 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U842 ( .A(n1184), .B(n1185), .ZN(n1183) );
NAND3_X1 U843 ( .A1(n1175), .A2(G472), .A3(KEYINPUT1), .ZN(n1184) );
INV_X1 U844 ( .A(n1167), .ZN(n1175) );
NOR2_X1 U845 ( .A1(n1162), .A2(n1186), .ZN(G54) );
XOR2_X1 U846 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U847 ( .A(n1189), .B(n1190), .ZN(n1188) );
XNOR2_X1 U848 ( .A(n1138), .B(n1191), .ZN(n1187) );
XOR2_X1 U849 ( .A(KEYINPUT57), .B(n1192), .Z(n1191) );
NOR2_X1 U850 ( .A1(n1193), .A2(n1167), .ZN(n1192) );
NOR2_X1 U851 ( .A1(n1162), .A2(n1194), .ZN(G51) );
XOR2_X1 U852 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U853 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U854 ( .A1(n1123), .A2(n1167), .ZN(n1198) );
NAND2_X1 U855 ( .A1(G902), .A2(n1199), .ZN(n1167) );
NAND3_X1 U856 ( .A1(n1106), .A2(n1160), .A3(n1107), .ZN(n1199) );
AND4_X1 U857 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1107) );
NOR4_X1 U858 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
INV_X1 U859 ( .A(n1208), .ZN(n1207) );
INV_X1 U860 ( .A(n1209), .ZN(n1206) );
NAND2_X1 U861 ( .A1(n1099), .A2(n1210), .ZN(n1202) );
NAND2_X1 U862 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND4_X1 U863 ( .A1(n1213), .A2(n1100), .A3(n1088), .A4(n1214), .ZN(n1212) );
NAND2_X1 U864 ( .A1(n1215), .A2(n1216), .ZN(n1211) );
NAND3_X1 U865 ( .A1(n1065), .A2(n1088), .A3(n1067), .ZN(n1160) );
AND4_X1 U866 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1106) );
NOR4_X1 U867 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
NOR2_X1 U868 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
INV_X1 U869 ( .A(KEYINPUT8), .ZN(n1226) );
NOR2_X1 U870 ( .A1(KEYINPUT17), .A2(n1227), .ZN(n1223) );
NOR2_X1 U871 ( .A1(n1228), .A2(n1229), .ZN(n1222) );
INV_X1 U872 ( .A(n1230), .ZN(n1229) );
XNOR2_X1 U873 ( .A(n1213), .B(KEYINPUT31), .ZN(n1228) );
NOR3_X1 U874 ( .A1(n1091), .A2(n1231), .A3(n1232), .ZN(n1221) );
NOR2_X1 U875 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NOR3_X1 U876 ( .A1(n1235), .A2(KEYINPUT8), .A3(n1236), .ZN(n1234) );
NOR2_X1 U877 ( .A1(n1237), .A2(n1238), .ZN(n1231) );
AND3_X1 U878 ( .A1(KEYINPUT17), .A2(n1236), .A3(n1067), .ZN(n1237) );
NAND3_X1 U879 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1091) );
NOR2_X1 U880 ( .A1(n1179), .A2(n1242), .ZN(n1219) );
AND3_X1 U881 ( .A1(n1065), .A2(n1088), .A3(n1100), .ZN(n1179) );
INV_X1 U882 ( .A(n1068), .ZN(n1088) );
NOR4_X1 U883 ( .A1(n1243), .A2(n1244), .A3(KEYINPUT41), .A4(n1245), .ZN(n1197) );
INV_X1 U884 ( .A(n1246), .ZN(n1245) );
NOR3_X1 U885 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1244) );
AND2_X1 U886 ( .A1(n1247), .A2(n1249), .ZN(n1243) );
INV_X1 U887 ( .A(KEYINPUT45), .ZN(n1247) );
NOR2_X1 U888 ( .A1(n1127), .A2(G952), .ZN(n1162) );
XNOR2_X1 U889 ( .A(n1250), .B(n1200), .ZN(G48) );
NAND3_X1 U890 ( .A1(n1100), .A2(n1236), .A3(n1216), .ZN(n1200) );
XNOR2_X1 U891 ( .A(G146), .B(KEYINPUT38), .ZN(n1250) );
XNOR2_X1 U892 ( .A(G143), .B(n1201), .ZN(G45) );
NAND4_X1 U893 ( .A1(n1251), .A2(n1236), .A3(n1252), .A4(n1253), .ZN(n1201) );
XNOR2_X1 U894 ( .A(G140), .B(n1254), .ZN(G42) );
NAND3_X1 U895 ( .A1(n1099), .A2(n1213), .A3(n1255), .ZN(n1254) );
NOR3_X1 U896 ( .A1(n1235), .A2(n1256), .A3(n1068), .ZN(n1255) );
XNOR2_X1 U897 ( .A(n1257), .B(KEYINPUT15), .ZN(n1256) );
INV_X1 U898 ( .A(n1100), .ZN(n1235) );
NAND2_X1 U899 ( .A1(n1258), .A2(n1259), .ZN(G39) );
NAND2_X1 U900 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND2_X1 U901 ( .A1(n1262), .A2(n1263), .ZN(n1258) );
NAND2_X1 U902 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U903 ( .A1(G137), .A2(n1266), .ZN(n1265) );
OR2_X1 U904 ( .A1(n1266), .A2(n1260), .ZN(n1264) );
NOR2_X1 U905 ( .A1(KEYINPUT9), .A2(n1267), .ZN(n1260) );
INV_X1 U906 ( .A(KEYINPUT10), .ZN(n1266) );
INV_X1 U907 ( .A(n1261), .ZN(n1262) );
NAND2_X1 U908 ( .A1(n1099), .A2(n1268), .ZN(n1261) );
XOR2_X1 U909 ( .A(KEYINPUT34), .B(n1269), .Z(n1268) );
NOR2_X1 U910 ( .A1(n1270), .A2(n1079), .ZN(n1269) );
XNOR2_X1 U911 ( .A(G134), .B(n1208), .ZN(G36) );
NAND3_X1 U912 ( .A1(n1251), .A2(n1067), .A3(n1099), .ZN(n1208) );
XNOR2_X1 U913 ( .A(G131), .B(n1209), .ZN(G33) );
NAND3_X1 U914 ( .A1(n1251), .A2(n1100), .A3(n1099), .ZN(n1209) );
NOR2_X1 U915 ( .A1(n1271), .A2(n1102), .ZN(n1099) );
XOR2_X1 U916 ( .A(n1272), .B(KEYINPUT51), .Z(n1102) );
XNOR2_X1 U917 ( .A(KEYINPUT58), .B(n1103), .ZN(n1271) );
AND2_X1 U918 ( .A1(n1273), .A2(n1239), .ZN(n1251) );
XNOR2_X1 U919 ( .A(n1274), .B(n1205), .ZN(G30) );
AND3_X1 U920 ( .A1(n1067), .A2(n1236), .A3(n1216), .ZN(n1205) );
INV_X1 U921 ( .A(n1270), .ZN(n1216) );
NAND2_X1 U922 ( .A1(n1273), .A2(n1275), .ZN(n1270) );
NOR3_X1 U923 ( .A1(n1276), .A2(n1257), .A3(n1068), .ZN(n1273) );
INV_X1 U924 ( .A(n1104), .ZN(n1236) );
XOR2_X1 U925 ( .A(n1217), .B(n1277), .Z(G3) );
XOR2_X1 U926 ( .A(KEYINPUT20), .B(G101), .Z(n1277) );
NAND3_X1 U927 ( .A1(n1239), .A2(n1240), .A3(n1230), .ZN(n1217) );
XOR2_X1 U928 ( .A(n1204), .B(n1278), .Z(G27) );
NOR2_X1 U929 ( .A1(KEYINPUT47), .A2(n1148), .ZN(n1278) );
AND4_X1 U930 ( .A1(n1213), .A2(n1241), .A3(n1279), .A4(n1100), .ZN(n1204) );
NOR2_X1 U931 ( .A1(n1257), .A2(n1104), .ZN(n1279) );
INV_X1 U932 ( .A(n1214), .ZN(n1257) );
NAND2_X1 U933 ( .A1(n1076), .A2(n1280), .ZN(n1214) );
NAND4_X1 U934 ( .A1(G902), .A2(G953), .A3(n1281), .A4(n1130), .ZN(n1280) );
INV_X1 U935 ( .A(G900), .ZN(n1130) );
XNOR2_X1 U936 ( .A(G122), .B(n1218), .ZN(G24) );
NAND4_X1 U937 ( .A1(n1241), .A2(n1065), .A3(n1252), .A4(n1253), .ZN(n1218) );
NOR3_X1 U938 ( .A1(n1104), .A2(n1233), .A3(n1086), .ZN(n1065) );
INV_X1 U939 ( .A(n1110), .ZN(n1086) );
NOR2_X1 U940 ( .A1(n1240), .A2(n1275), .ZN(n1110) );
XOR2_X1 U941 ( .A(n1282), .B(n1242), .Z(G21) );
AND3_X1 U942 ( .A1(n1215), .A2(n1275), .A3(n1283), .ZN(n1242) );
NAND2_X1 U943 ( .A1(KEYINPUT21), .A2(n1284), .ZN(n1282) );
XNOR2_X1 U944 ( .A(G116), .B(n1227), .ZN(G18) );
NAND3_X1 U945 ( .A1(n1067), .A2(n1239), .A3(n1283), .ZN(n1227) );
NOR2_X1 U946 ( .A1(n1253), .A2(n1109), .ZN(n1067) );
INV_X1 U947 ( .A(n1252), .ZN(n1109) );
XOR2_X1 U948 ( .A(n1225), .B(n1285), .Z(G15) );
NOR2_X1 U949 ( .A1(G113), .A2(KEYINPUT13), .ZN(n1285) );
NAND3_X1 U950 ( .A1(n1100), .A2(n1239), .A3(n1283), .ZN(n1225) );
NOR4_X1 U951 ( .A1(n1092), .A2(n1104), .A3(n1276), .A4(n1233), .ZN(n1283) );
INV_X1 U952 ( .A(n1241), .ZN(n1092) );
NOR2_X1 U953 ( .A1(n1090), .A2(n1115), .ZN(n1241) );
XOR2_X1 U954 ( .A(n1286), .B(KEYINPUT55), .Z(n1090) );
XOR2_X1 U955 ( .A(n1275), .B(KEYINPUT46), .Z(n1239) );
NOR2_X1 U956 ( .A1(n1252), .A2(n1287), .ZN(n1100) );
XNOR2_X1 U957 ( .A(G110), .B(n1288), .ZN(G12) );
NAND2_X1 U958 ( .A1(n1230), .A2(n1213), .ZN(n1288) );
INV_X1 U959 ( .A(n1093), .ZN(n1213) );
NAND2_X1 U960 ( .A1(n1276), .A2(n1275), .ZN(n1093) );
XOR2_X1 U961 ( .A(n1289), .B(n1166), .Z(n1275) );
NAND2_X1 U962 ( .A1(G217), .A2(n1290), .ZN(n1166) );
NAND2_X1 U963 ( .A1(n1164), .A2(n1291), .ZN(n1289) );
XNOR2_X1 U964 ( .A(n1292), .B(n1293), .ZN(n1164) );
XNOR2_X1 U965 ( .A(n1284), .B(n1294), .ZN(n1293) );
XNOR2_X1 U966 ( .A(n1267), .B(G128), .ZN(n1294) );
XOR2_X1 U967 ( .A(n1295), .B(n1296), .Z(n1292) );
XNOR2_X1 U968 ( .A(n1297), .B(n1298), .ZN(n1296) );
NOR2_X1 U969 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U970 ( .A(n1301), .B(KEYINPUT26), .Z(n1300) );
NAND2_X1 U971 ( .A1(G146), .A2(n1302), .ZN(n1301) );
NOR2_X1 U972 ( .A1(G146), .A2(n1302), .ZN(n1299) );
NAND2_X1 U973 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U974 ( .A1(n1305), .A2(n1145), .ZN(n1304) );
NAND2_X1 U975 ( .A1(n1306), .A2(n1148), .ZN(n1303) );
NAND2_X1 U976 ( .A1(n1305), .A2(n1307), .ZN(n1306) );
XNOR2_X1 U977 ( .A(KEYINPUT14), .B(KEYINPUT2), .ZN(n1305) );
NAND2_X1 U978 ( .A1(G221), .A2(n1308), .ZN(n1295) );
INV_X1 U979 ( .A(n1240), .ZN(n1276) );
XNOR2_X1 U980 ( .A(n1309), .B(G472), .ZN(n1240) );
NAND3_X1 U981 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1309) );
XNOR2_X1 U982 ( .A(KEYINPUT43), .B(n1291), .ZN(n1312) );
NAND2_X1 U983 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
INV_X1 U984 ( .A(KEYINPUT59), .ZN(n1314) );
XNOR2_X1 U985 ( .A(n1182), .B(n1315), .ZN(n1313) );
INV_X1 U986 ( .A(n1185), .ZN(n1315) );
NAND3_X1 U987 ( .A1(n1185), .A2(n1182), .A3(KEYINPUT59), .ZN(n1310) );
XOR2_X1 U988 ( .A(n1316), .B(n1317), .Z(n1182) );
XOR2_X1 U989 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U990 ( .A(G113), .B(G116), .ZN(n1319) );
NAND2_X1 U991 ( .A1(KEYINPUT4), .A2(G119), .ZN(n1318) );
XOR2_X1 U992 ( .A(n1320), .B(n1321), .Z(n1316) );
XNOR2_X1 U993 ( .A(n1322), .B(n1323), .ZN(n1185) );
NAND3_X1 U994 ( .A1(n1324), .A2(n1127), .A3(G210), .ZN(n1322) );
NOR4_X1 U995 ( .A1(n1079), .A2(n1068), .A3(n1104), .A4(n1233), .ZN(n1230) );
INV_X1 U996 ( .A(n1238), .ZN(n1233) );
NAND2_X1 U997 ( .A1(n1325), .A2(n1076), .ZN(n1238) );
NAND3_X1 U998 ( .A1(n1105), .A2(n1281), .A3(n1326), .ZN(n1076) );
XNOR2_X1 U999 ( .A(G952), .B(KEYINPUT52), .ZN(n1326) );
INV_X1 U1000 ( .A(n1108), .ZN(n1105) );
XOR2_X1 U1001 ( .A(G953), .B(KEYINPUT42), .Z(n1108) );
NAND4_X1 U1002 ( .A1(G902), .A2(G953), .A3(n1281), .A4(n1153), .ZN(n1325) );
INV_X1 U1003 ( .A(G898), .ZN(n1153) );
NAND2_X1 U1004 ( .A1(G234), .A2(G237), .ZN(n1281) );
NAND2_X1 U1005 ( .A1(n1327), .A2(n1272), .ZN(n1104) );
NAND3_X1 U1006 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1272) );
NAND2_X1 U1007 ( .A1(KEYINPUT6), .A2(n1124), .ZN(n1330) );
OR3_X1 U1008 ( .A1(n1124), .A2(KEYINPUT6), .A3(n1123), .ZN(n1329) );
NAND2_X1 U1009 ( .A1(n1331), .A2(n1123), .ZN(n1328) );
NAND2_X1 U1010 ( .A1(G210), .A2(n1332), .ZN(n1123) );
NAND2_X1 U1011 ( .A1(n1333), .A2(n1334), .ZN(n1331) );
INV_X1 U1012 ( .A(KEYINPUT6), .ZN(n1334) );
XNOR2_X1 U1013 ( .A(n1124), .B(KEYINPUT61), .ZN(n1333) );
AND2_X1 U1014 ( .A1(n1335), .A2(n1291), .ZN(n1124) );
XNOR2_X1 U1015 ( .A(n1336), .B(n1195), .ZN(n1335) );
XNOR2_X1 U1016 ( .A(n1161), .B(KEYINPUT27), .ZN(n1195) );
XOR2_X1 U1017 ( .A(n1337), .B(n1338), .Z(n1161) );
XOR2_X1 U1018 ( .A(n1339), .B(n1340), .Z(n1338) );
XNOR2_X1 U1019 ( .A(n1284), .B(G116), .ZN(n1340) );
INV_X1 U1020 ( .A(G119), .ZN(n1284) );
XOR2_X1 U1021 ( .A(KEYINPUT56), .B(G122), .Z(n1339) );
XNOR2_X1 U1022 ( .A(n1341), .B(n1342), .ZN(n1337) );
INV_X1 U1023 ( .A(n1190), .ZN(n1342) );
XOR2_X1 U1024 ( .A(G110), .B(n1323), .Z(n1190) );
XOR2_X1 U1025 ( .A(n1343), .B(G113), .Z(n1341) );
NAND3_X1 U1026 ( .A1(n1344), .A2(n1345), .A3(n1346), .ZN(n1343) );
NAND2_X1 U1027 ( .A1(G107), .A2(n1347), .ZN(n1346) );
NAND2_X1 U1028 ( .A1(KEYINPUT32), .A2(n1348), .ZN(n1345) );
NAND2_X1 U1029 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
XNOR2_X1 U1030 ( .A(KEYINPUT0), .B(n1347), .ZN(n1349) );
NAND2_X1 U1031 ( .A1(n1351), .A2(n1352), .ZN(n1344) );
INV_X1 U1032 ( .A(KEYINPUT32), .ZN(n1352) );
NAND2_X1 U1033 ( .A1(n1353), .A2(n1354), .ZN(n1351) );
NAND2_X1 U1034 ( .A1(KEYINPUT0), .A2(n1347), .ZN(n1354) );
OR3_X1 U1035 ( .A1(G107), .A2(KEYINPUT0), .A3(n1347), .ZN(n1353) );
NAND2_X1 U1036 ( .A1(KEYINPUT5), .A2(n1355), .ZN(n1336) );
NAND2_X1 U1037 ( .A1(n1356), .A2(n1246), .ZN(n1355) );
NAND2_X1 U1038 ( .A1(n1248), .A2(n1249), .ZN(n1246) );
OR2_X1 U1039 ( .A1(n1249), .A2(n1248), .ZN(n1356) );
NOR2_X1 U1040 ( .A1(n1152), .A2(G953), .ZN(n1248) );
INV_X1 U1041 ( .A(G224), .ZN(n1152) );
XNOR2_X1 U1042 ( .A(n1321), .B(n1357), .ZN(n1249) );
XNOR2_X1 U1043 ( .A(KEYINPUT19), .B(n1148), .ZN(n1357) );
XNOR2_X1 U1044 ( .A(n1358), .B(n1359), .ZN(n1321) );
XNOR2_X1 U1045 ( .A(G143), .B(n1360), .ZN(n1359) );
NAND2_X1 U1046 ( .A1(KEYINPUT60), .A2(n1361), .ZN(n1360) );
XNOR2_X1 U1047 ( .A(KEYINPUT16), .B(n1274), .ZN(n1361) );
INV_X1 U1048 ( .A(G128), .ZN(n1274) );
NAND2_X1 U1049 ( .A1(KEYINPUT25), .A2(n1362), .ZN(n1358) );
XNOR2_X1 U1050 ( .A(KEYINPUT58), .B(n1113), .ZN(n1327) );
INV_X1 U1051 ( .A(n1103), .ZN(n1113) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1332), .ZN(n1103) );
NAND2_X1 U1053 ( .A1(n1363), .A2(n1291), .ZN(n1332) );
NAND2_X1 U1054 ( .A1(n1364), .A2(n1286), .ZN(n1068) );
XNOR2_X1 U1055 ( .A(n1122), .B(n1365), .ZN(n1286) );
NOR2_X1 U1056 ( .A1(KEYINPUT54), .A2(n1193), .ZN(n1365) );
INV_X1 U1057 ( .A(G469), .ZN(n1193) );
NAND2_X1 U1058 ( .A1(n1366), .A2(n1291), .ZN(n1122) );
XOR2_X1 U1059 ( .A(n1367), .B(n1368), .Z(n1366) );
XOR2_X1 U1060 ( .A(n1189), .B(n1323), .Z(n1368) );
XOR2_X1 U1061 ( .A(G101), .B(KEYINPUT29), .Z(n1323) );
XOR2_X1 U1062 ( .A(n1369), .B(n1370), .Z(n1189) );
XNOR2_X1 U1063 ( .A(n1347), .B(n1371), .ZN(n1370) );
XNOR2_X1 U1064 ( .A(n1307), .B(G107), .ZN(n1371) );
INV_X1 U1065 ( .A(G104), .ZN(n1347) );
XOR2_X1 U1066 ( .A(n1320), .B(n1372), .Z(n1369) );
NOR2_X1 U1067 ( .A1(G953), .A2(n1129), .ZN(n1372) );
INV_X1 U1068 ( .A(G227), .ZN(n1129) );
XNOR2_X1 U1069 ( .A(G131), .B(n1140), .ZN(n1320) );
XNOR2_X1 U1070 ( .A(G134), .B(n1267), .ZN(n1140) );
INV_X1 U1071 ( .A(G137), .ZN(n1267) );
XOR2_X1 U1072 ( .A(n1373), .B(n1374), .Z(n1367) );
XNOR2_X1 U1073 ( .A(n1375), .B(KEYINPUT7), .ZN(n1374) );
NAND2_X1 U1074 ( .A1(KEYINPUT28), .A2(n1297), .ZN(n1375) );
INV_X1 U1075 ( .A(G110), .ZN(n1297) );
NAND2_X1 U1076 ( .A1(KEYINPUT50), .A2(n1138), .ZN(n1373) );
XOR2_X1 U1077 ( .A(G128), .B(n1376), .Z(n1138) );
XNOR2_X1 U1078 ( .A(n1115), .B(KEYINPUT11), .ZN(n1364) );
INV_X1 U1079 ( .A(n1089), .ZN(n1115) );
NAND2_X1 U1080 ( .A1(G221), .A2(n1290), .ZN(n1089) );
NAND2_X1 U1081 ( .A1(G234), .A2(n1291), .ZN(n1290) );
INV_X1 U1082 ( .A(n1215), .ZN(n1079) );
NOR2_X1 U1083 ( .A1(n1252), .A2(n1253), .ZN(n1215) );
INV_X1 U1084 ( .A(n1287), .ZN(n1253) );
NOR2_X1 U1085 ( .A1(n1377), .A2(n1114), .ZN(n1287) );
NOR2_X1 U1086 ( .A1(n1119), .A2(G475), .ZN(n1114) );
AND2_X1 U1087 ( .A1(n1378), .A2(n1119), .ZN(n1377) );
NAND2_X1 U1088 ( .A1(n1178), .A2(n1291), .ZN(n1119) );
XOR2_X1 U1089 ( .A(n1379), .B(n1380), .Z(n1178) );
XNOR2_X1 U1090 ( .A(n1381), .B(n1376), .ZN(n1380) );
XNOR2_X1 U1091 ( .A(G143), .B(n1362), .ZN(n1376) );
INV_X1 U1092 ( .A(G146), .ZN(n1362) );
NAND3_X1 U1093 ( .A1(n1382), .A2(n1383), .A3(n1384), .ZN(n1381) );
NAND2_X1 U1094 ( .A1(n1145), .A2(n1142), .ZN(n1384) );
INV_X1 U1095 ( .A(G131), .ZN(n1142) );
NOR2_X1 U1096 ( .A1(n1148), .A2(G140), .ZN(n1145) );
NAND3_X1 U1097 ( .A1(G131), .A2(n1148), .A3(n1307), .ZN(n1383) );
INV_X1 U1098 ( .A(G140), .ZN(n1307) );
INV_X1 U1099 ( .A(G125), .ZN(n1148) );
NAND2_X1 U1100 ( .A1(n1385), .A2(G140), .ZN(n1382) );
XNOR2_X1 U1101 ( .A(G125), .B(G131), .ZN(n1385) );
XOR2_X1 U1102 ( .A(n1386), .B(n1387), .Z(n1379) );
AND3_X1 U1103 ( .A1(G214), .A2(n1127), .A3(n1324), .ZN(n1387) );
XOR2_X1 U1104 ( .A(n1363), .B(KEYINPUT22), .Z(n1324) );
INV_X1 U1105 ( .A(G237), .ZN(n1363) );
NAND2_X1 U1106 ( .A1(n1388), .A2(n1389), .ZN(n1386) );
OR2_X1 U1107 ( .A1(n1390), .A2(G104), .ZN(n1389) );
XOR2_X1 U1108 ( .A(n1391), .B(KEYINPUT48), .Z(n1388) );
NAND2_X1 U1109 ( .A1(G104), .A2(n1390), .ZN(n1391) );
XOR2_X1 U1110 ( .A(G113), .B(G122), .Z(n1390) );
XOR2_X1 U1111 ( .A(KEYINPUT33), .B(G475), .Z(n1378) );
XNOR2_X1 U1112 ( .A(n1392), .B(G478), .ZN(n1252) );
NAND2_X1 U1113 ( .A1(n1393), .A2(n1291), .ZN(n1392) );
INV_X1 U1114 ( .A(G902), .ZN(n1291) );
XNOR2_X1 U1115 ( .A(n1173), .B(n1174), .ZN(n1393) );
XNOR2_X1 U1116 ( .A(n1394), .B(n1395), .ZN(n1174) );
NOR2_X1 U1117 ( .A1(KEYINPUT24), .A2(n1396), .ZN(n1395) );
INV_X1 U1118 ( .A(G134), .ZN(n1396) );
NAND2_X1 U1119 ( .A1(G217), .A2(n1308), .ZN(n1394) );
AND2_X1 U1120 ( .A1(G234), .A2(n1127), .ZN(n1308) );
INV_X1 U1121 ( .A(G953), .ZN(n1127) );
XOR2_X1 U1122 ( .A(n1397), .B(n1398), .Z(n1173) );
NOR2_X1 U1123 ( .A1(n1399), .A2(n1400), .ZN(n1398) );
XOR2_X1 U1124 ( .A(n1401), .B(KEYINPUT23), .Z(n1400) );
NAND2_X1 U1125 ( .A1(n1402), .A2(n1350), .ZN(n1401) );
INV_X1 U1126 ( .A(G107), .ZN(n1350) );
XOR2_X1 U1127 ( .A(KEYINPUT12), .B(n1403), .Z(n1402) );
AND2_X1 U1128 ( .A1(n1403), .A2(G107), .ZN(n1399) );
XOR2_X1 U1129 ( .A(G116), .B(G122), .Z(n1403) );
XNOR2_X1 U1130 ( .A(G128), .B(G143), .ZN(n1397) );
endmodule


