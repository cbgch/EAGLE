//Key = 0110100111101010111111111110000010001011000001001101011001010110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311;

XNOR2_X1 U720 ( .A(G107), .B(n1000), .ZN(G9) );
NOR2_X1 U721 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR3_X1 U722 ( .A1(n1003), .A2(G953), .A3(n1004), .ZN(n1002) );
INV_X1 U723 ( .A(n1005), .ZN(n1004) );
XNOR2_X1 U724 ( .A(KEYINPUT63), .B(n1006), .ZN(n1003) );
NOR4_X1 U725 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1006), .ZN(n1001) );
INV_X1 U726 ( .A(G952), .ZN(n1006) );
NOR2_X1 U727 ( .A1(n1010), .A2(KEYINPUT26), .ZN(n1009) );
AND4_X1 U728 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
NAND4_X1 U729 ( .A1(n1015), .A2(n1005), .A3(n1016), .A4(n1017), .ZN(n1007) );
NAND4_X1 U730 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1016) );
NOR2_X1 U731 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U732 ( .A1(n1024), .A2(n1025), .ZN(n1019) );
NAND2_X1 U733 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NAND3_X1 U734 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1027) );
NAND2_X1 U735 ( .A1(n1031), .A2(n1032), .ZN(n1018) );
NAND4_X1 U736 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1005) );
NOR3_X1 U737 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR2_X1 U738 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND3_X1 U739 ( .A1(n1042), .A2(n1043), .A3(n1028), .ZN(n1037) );
NOR3_X1 U740 ( .A1(n1022), .A2(n1044), .A3(n1045), .ZN(n1035) );
NOR3_X1 U741 ( .A1(n1046), .A2(KEYINPUT58), .A3(n1047), .ZN(n1045) );
AND2_X1 U742 ( .A1(n1046), .A2(KEYINPUT58), .ZN(n1044) );
NAND4_X1 U743 ( .A1(n1014), .A2(n1013), .A3(n1011), .A4(n1048), .ZN(n1015) );
NAND3_X1 U744 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND2_X1 U745 ( .A1(KEYINPUT26), .A2(n1012), .ZN(n1051) );
NAND2_X1 U746 ( .A1(n1020), .A2(n1052), .ZN(n1050) );
NAND2_X1 U747 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
OR2_X1 U748 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U749 ( .A1(n1057), .A2(n1058), .ZN(n1049) );
INV_X1 U750 ( .A(n1023), .ZN(n1014) );
XOR2_X1 U751 ( .A(n1059), .B(n1060), .Z(G72) );
NOR2_X1 U752 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
XNOR2_X1 U753 ( .A(n1063), .B(n1064), .ZN(n1062) );
NAND4_X1 U754 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1059) );
INV_X1 U755 ( .A(n1061), .ZN(n1068) );
NAND2_X1 U756 ( .A1(G953), .A2(n1069), .ZN(n1066) );
XOR2_X1 U757 ( .A(n1070), .B(n1071), .Z(G69) );
NAND2_X1 U758 ( .A1(G953), .A2(n1072), .ZN(n1071) );
NAND2_X1 U759 ( .A1(G898), .A2(G224), .ZN(n1072) );
NAND3_X1 U760 ( .A1(n1073), .A2(n1074), .A3(KEYINPUT38), .ZN(n1070) );
NAND2_X1 U761 ( .A1(KEYINPUT8), .A2(n1075), .ZN(n1074) );
XOR2_X1 U762 ( .A(n1076), .B(n1077), .Z(n1075) );
OR3_X1 U763 ( .A1(n1076), .A2(n1077), .A3(KEYINPUT8), .ZN(n1073) );
NOR2_X1 U764 ( .A1(G953), .A2(n1078), .ZN(n1077) );
NAND2_X1 U765 ( .A1(n1079), .A2(n1080), .ZN(n1076) );
NAND2_X1 U766 ( .A1(G953), .A2(n1081), .ZN(n1080) );
XNOR2_X1 U767 ( .A(n1082), .B(n1083), .ZN(n1079) );
XNOR2_X1 U768 ( .A(n1084), .B(n1085), .ZN(n1083) );
NAND2_X1 U769 ( .A1(KEYINPUT62), .A2(n1086), .ZN(n1084) );
NOR2_X1 U770 ( .A1(n1087), .A2(n1088), .ZN(G66) );
XOR2_X1 U771 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U772 ( .A1(n1046), .A2(n1091), .ZN(n1090) );
NOR2_X1 U773 ( .A1(n1087), .A2(n1092), .ZN(G63) );
XOR2_X1 U774 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR3_X1 U775 ( .A1(n1091), .A2(KEYINPUT3), .A3(n1041), .ZN(n1093) );
NOR2_X1 U776 ( .A1(n1087), .A2(n1095), .ZN(G60) );
XNOR2_X1 U777 ( .A(n1096), .B(n1097), .ZN(n1095) );
NOR3_X1 U778 ( .A1(n1091), .A2(KEYINPUT0), .A3(n1098), .ZN(n1097) );
XOR2_X1 U779 ( .A(n1099), .B(n1100), .Z(G6) );
NAND2_X1 U780 ( .A1(KEYINPUT51), .A2(G104), .ZN(n1100) );
NOR2_X1 U781 ( .A1(n1087), .A2(n1101), .ZN(G57) );
XOR2_X1 U782 ( .A(n1102), .B(n1103), .Z(n1101) );
XNOR2_X1 U783 ( .A(G101), .B(n1104), .ZN(n1103) );
XNOR2_X1 U784 ( .A(KEYINPUT61), .B(KEYINPUT29), .ZN(n1104) );
XOR2_X1 U785 ( .A(n1105), .B(n1106), .Z(n1102) );
NOR2_X1 U786 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U787 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U788 ( .A(KEYINPUT33), .B(n1111), .Z(n1109) );
AND2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NOR2_X1 U790 ( .A1(n1091), .A2(n1112), .ZN(n1111) );
INV_X1 U791 ( .A(G472), .ZN(n1112) );
XOR2_X1 U792 ( .A(n1113), .B(n1114), .Z(n1110) );
XNOR2_X1 U793 ( .A(n1115), .B(n1116), .ZN(n1113) );
NOR2_X1 U794 ( .A1(KEYINPUT56), .A2(n1117), .ZN(n1116) );
NOR2_X1 U795 ( .A1(n1087), .A2(n1118), .ZN(G54) );
XOR2_X1 U796 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U797 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U798 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XOR2_X1 U799 ( .A(KEYINPUT27), .B(n1125), .Z(n1124) );
AND2_X1 U800 ( .A1(n1115), .A2(n1126), .ZN(n1125) );
NOR2_X1 U801 ( .A1(n1115), .A2(n1126), .ZN(n1123) );
XOR2_X1 U802 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U803 ( .A1(KEYINPUT42), .A2(n1129), .ZN(n1128) );
XOR2_X1 U804 ( .A(n1130), .B(KEYINPUT32), .Z(n1129) );
NOR2_X1 U805 ( .A1(KEYINPUT28), .A2(n1131), .ZN(n1121) );
XNOR2_X1 U806 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR2_X1 U807 ( .A1(KEYINPUT13), .A2(n1134), .ZN(n1133) );
XNOR2_X1 U808 ( .A(G110), .B(KEYINPUT4), .ZN(n1134) );
NOR2_X1 U809 ( .A1(n1135), .A2(n1091), .ZN(n1119) );
NOR2_X1 U810 ( .A1(n1087), .A2(n1136), .ZN(G51) );
XOR2_X1 U811 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U812 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U813 ( .A1(n1141), .A2(n1091), .ZN(n1140) );
NAND2_X1 U814 ( .A1(G902), .A2(n1008), .ZN(n1091) );
NAND3_X1 U815 ( .A1(n1065), .A2(n1142), .A3(n1078), .ZN(n1008) );
AND4_X1 U816 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1078) );
AND4_X1 U817 ( .A1(n1000), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1146) );
NAND2_X1 U818 ( .A1(n1058), .A2(n1150), .ZN(n1000) );
NOR4_X1 U819 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1145) );
NOR2_X1 U820 ( .A1(KEYINPUT9), .A2(n1155), .ZN(n1154) );
NAND4_X1 U821 ( .A1(n1012), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1155) );
NOR2_X1 U822 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
INV_X1 U823 ( .A(KEYINPUT9), .ZN(n1159) );
NOR2_X1 U824 ( .A1(n1161), .A2(n1099), .ZN(n1152) );
NAND2_X1 U825 ( .A1(n1162), .A2(n1150), .ZN(n1099) );
AND3_X1 U826 ( .A1(n1163), .A2(n1164), .A3(n1011), .ZN(n1150) );
INV_X1 U827 ( .A(KEYINPUT21), .ZN(n1161) );
NOR4_X1 U828 ( .A1(KEYINPUT21), .A2(n1165), .A3(n1032), .A4(n1166), .ZN(n1151) );
INV_X1 U829 ( .A(n1011), .ZN(n1032) );
NAND3_X1 U830 ( .A1(n1167), .A2(n1025), .A3(n1164), .ZN(n1165) );
NAND3_X1 U831 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(n1143) );
XNOR2_X1 U832 ( .A(n1057), .B(KEYINPUT39), .ZN(n1170) );
XNOR2_X1 U833 ( .A(KEYINPUT14), .B(n1067), .ZN(n1142) );
AND4_X1 U834 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1065) );
AND3_X1 U835 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1174) );
NAND3_X1 U836 ( .A1(n1178), .A2(n1179), .A3(n1012), .ZN(n1177) );
NAND2_X1 U837 ( .A1(n1157), .A2(n1180), .ZN(n1173) );
NAND2_X1 U838 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U839 ( .A1(n1183), .A2(n1162), .ZN(n1181) );
NAND2_X1 U840 ( .A1(KEYINPUT59), .A2(n1184), .ZN(n1139) );
XOR2_X1 U841 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U842 ( .A1(KEYINPUT5), .A2(n1187), .ZN(n1185) );
NOR2_X1 U843 ( .A1(n1017), .A2(G952), .ZN(n1087) );
XOR2_X1 U844 ( .A(n1176), .B(n1188), .Z(G48) );
NOR2_X1 U845 ( .A1(G146), .A2(KEYINPUT15), .ZN(n1188) );
NAND4_X1 U846 ( .A1(n1189), .A2(n1178), .A3(n1162), .A4(n1168), .ZN(n1176) );
XOR2_X1 U847 ( .A(n1190), .B(n1191), .Z(G45) );
NAND2_X1 U848 ( .A1(n1192), .A2(KEYINPUT48), .ZN(n1191) );
XNOR2_X1 U849 ( .A(G143), .B(KEYINPUT19), .ZN(n1192) );
NAND2_X1 U850 ( .A1(n1193), .A2(n1194), .ZN(n1190) );
XNOR2_X1 U851 ( .A(KEYINPUT31), .B(n1029), .ZN(n1194) );
INV_X1 U852 ( .A(n1182), .ZN(n1193) );
NAND4_X1 U853 ( .A1(n1189), .A2(n1178), .A3(n1039), .A4(n1195), .ZN(n1182) );
XOR2_X1 U854 ( .A(n1172), .B(n1196), .Z(G42) );
NAND2_X1 U855 ( .A1(KEYINPUT16), .A2(G140), .ZN(n1196) );
NAND3_X1 U856 ( .A1(n1162), .A2(n1179), .A3(n1183), .ZN(n1172) );
NAND2_X1 U857 ( .A1(n1197), .A2(n1198), .ZN(G39) );
NAND2_X1 U858 ( .A1(G137), .A2(n1171), .ZN(n1198) );
XOR2_X1 U859 ( .A(n1199), .B(KEYINPUT60), .Z(n1197) );
OR2_X1 U860 ( .A1(n1171), .A2(G137), .ZN(n1199) );
NAND3_X1 U861 ( .A1(n1168), .A2(n1020), .A3(n1183), .ZN(n1171) );
XNOR2_X1 U862 ( .A(G134), .B(n1067), .ZN(G36) );
NAND3_X1 U863 ( .A1(n1157), .A2(n1058), .A3(n1183), .ZN(n1067) );
INV_X1 U864 ( .A(n1200), .ZN(n1183) );
XNOR2_X1 U865 ( .A(n1201), .B(n1202), .ZN(G33) );
NOR4_X1 U866 ( .A1(KEYINPUT40), .A2(n1029), .A3(n1166), .A4(n1200), .ZN(n1202) );
NAND3_X1 U867 ( .A1(n1189), .A2(n1203), .A3(n1013), .ZN(n1200) );
INV_X1 U868 ( .A(n1031), .ZN(n1013) );
NAND2_X1 U869 ( .A1(n1026), .A2(n1028), .ZN(n1031) );
INV_X1 U870 ( .A(n1053), .ZN(n1189) );
XNOR2_X1 U871 ( .A(n1204), .B(KEYINPUT2), .ZN(n1053) );
INV_X1 U872 ( .A(n1157), .ZN(n1029) );
XNOR2_X1 U873 ( .A(G128), .B(n1175), .ZN(G30) );
NAND4_X1 U874 ( .A1(n1178), .A2(n1168), .A3(n1058), .A4(n1164), .ZN(n1175) );
NAND2_X1 U875 ( .A1(n1205), .A2(n1206), .ZN(G3) );
NAND2_X1 U876 ( .A1(G101), .A2(n1144), .ZN(n1206) );
XOR2_X1 U877 ( .A(KEYINPUT22), .B(n1207), .Z(n1205) );
NOR2_X1 U878 ( .A1(G101), .A2(n1144), .ZN(n1207) );
NAND3_X1 U879 ( .A1(n1169), .A2(n1164), .A3(n1157), .ZN(n1144) );
XNOR2_X1 U880 ( .A(G125), .B(n1208), .ZN(G27) );
NAND4_X1 U881 ( .A1(n1209), .A2(n1178), .A3(n1162), .A4(n1179), .ZN(n1208) );
AND2_X1 U882 ( .A1(n1158), .A2(n1203), .ZN(n1178) );
NAND2_X1 U883 ( .A1(n1023), .A2(n1210), .ZN(n1203) );
NAND3_X1 U884 ( .A1(G902), .A2(n1211), .A3(n1061), .ZN(n1210) );
NOR2_X1 U885 ( .A1(G900), .A2(n1017), .ZN(n1061) );
XNOR2_X1 U886 ( .A(n1057), .B(KEYINPUT10), .ZN(n1209) );
XNOR2_X1 U887 ( .A(G122), .B(n1149), .ZN(G24) );
NAND4_X1 U888 ( .A1(n1057), .A2(n1011), .A3(n1212), .A4(n1163), .ZN(n1149) );
NOR2_X1 U889 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
NOR2_X1 U890 ( .A1(n1215), .A2(n1216), .ZN(n1011) );
XNOR2_X1 U891 ( .A(G119), .B(n1217), .ZN(G21) );
NAND3_X1 U892 ( .A1(n1057), .A2(n1169), .A3(n1168), .ZN(n1217) );
AND2_X1 U893 ( .A1(n1216), .A2(n1215), .ZN(n1168) );
INV_X1 U894 ( .A(n1033), .ZN(n1216) );
XNOR2_X1 U895 ( .A(G116), .B(n1148), .ZN(G18) );
NAND4_X1 U896 ( .A1(n1057), .A2(n1157), .A3(n1058), .A4(n1163), .ZN(n1148) );
NOR2_X1 U897 ( .A1(n1039), .A2(n1213), .ZN(n1058) );
INV_X1 U898 ( .A(n1195), .ZN(n1213) );
XNOR2_X1 U899 ( .A(G113), .B(n1160), .ZN(G15) );
NAND3_X1 U900 ( .A1(n1157), .A2(n1163), .A3(n1012), .ZN(n1160) );
NOR2_X1 U901 ( .A1(n1166), .A2(n1022), .ZN(n1012) );
INV_X1 U902 ( .A(n1057), .ZN(n1022) );
NOR2_X1 U903 ( .A1(n1056), .A2(n1218), .ZN(n1057) );
INV_X1 U904 ( .A(n1055), .ZN(n1218) );
INV_X1 U905 ( .A(n1162), .ZN(n1166) );
NOR2_X1 U906 ( .A1(n1195), .A2(n1214), .ZN(n1162) );
INV_X1 U907 ( .A(n1039), .ZN(n1214) );
NOR2_X1 U908 ( .A1(n1215), .A2(n1033), .ZN(n1157) );
XNOR2_X1 U909 ( .A(G110), .B(n1147), .ZN(G12) );
NAND3_X1 U910 ( .A1(n1169), .A2(n1164), .A3(n1179), .ZN(n1147) );
INV_X1 U911 ( .A(n1030), .ZN(n1179) );
NAND2_X1 U912 ( .A1(n1033), .A2(n1215), .ZN(n1030) );
NAND2_X1 U913 ( .A1(n1043), .A2(n1219), .ZN(n1215) );
OR2_X1 U914 ( .A1(n1046), .A2(n1047), .ZN(n1219) );
NAND2_X1 U915 ( .A1(n1047), .A2(n1046), .ZN(n1043) );
NAND2_X1 U916 ( .A1(G217), .A2(n1220), .ZN(n1046) );
NOR2_X1 U917 ( .A1(n1089), .A2(G902), .ZN(n1047) );
XOR2_X1 U918 ( .A(n1221), .B(n1222), .Z(n1089) );
XNOR2_X1 U919 ( .A(n1223), .B(n1224), .ZN(n1222) );
NAND2_X1 U920 ( .A1(KEYINPUT54), .A2(n1225), .ZN(n1223) );
XOR2_X1 U921 ( .A(n1226), .B(n1227), .Z(n1221) );
NOR2_X1 U922 ( .A1(KEYINPUT30), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U923 ( .A(G128), .B(n1229), .ZN(n1228) );
XNOR2_X1 U924 ( .A(n1230), .B(n1231), .ZN(n1226) );
NAND3_X1 U925 ( .A1(n1232), .A2(n1017), .A3(G234), .ZN(n1230) );
XOR2_X1 U926 ( .A(KEYINPUT47), .B(G221), .Z(n1232) );
XOR2_X1 U927 ( .A(n1233), .B(G472), .Z(n1033) );
NAND2_X1 U928 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U929 ( .A(n1236), .B(n1237), .Z(n1234) );
XNOR2_X1 U930 ( .A(n1238), .B(n1239), .ZN(n1237) );
NOR2_X1 U931 ( .A1(KEYINPUT52), .A2(n1240), .ZN(n1239) );
INV_X1 U932 ( .A(n1115), .ZN(n1240) );
NAND2_X1 U933 ( .A1(n1241), .A2(KEYINPUT24), .ZN(n1238) );
XOR2_X1 U934 ( .A(n1242), .B(n1243), .Z(n1241) );
XNOR2_X1 U935 ( .A(KEYINPUT49), .B(n1105), .ZN(n1243) );
NAND3_X1 U936 ( .A1(G210), .A2(n1017), .A3(n1244), .ZN(n1105) );
XNOR2_X1 U937 ( .A(G237), .B(KEYINPUT41), .ZN(n1244) );
NAND2_X1 U938 ( .A1(KEYINPUT25), .A2(n1245), .ZN(n1242) );
INV_X1 U939 ( .A(G101), .ZN(n1245) );
XOR2_X1 U940 ( .A(n1117), .B(n1114), .Z(n1236) );
XOR2_X1 U941 ( .A(n1246), .B(G113), .Z(n1114) );
XOR2_X1 U942 ( .A(n1247), .B(KEYINPUT57), .Z(n1117) );
XNOR2_X1 U943 ( .A(n1204), .B(KEYINPUT44), .ZN(n1164) );
NAND2_X1 U944 ( .A1(n1056), .A2(n1055), .ZN(n1204) );
NAND2_X1 U945 ( .A1(G221), .A2(n1220), .ZN(n1055) );
NAND2_X1 U946 ( .A1(G234), .A2(n1235), .ZN(n1220) );
XOR2_X1 U947 ( .A(n1248), .B(n1135), .Z(n1056) );
INV_X1 U948 ( .A(G469), .ZN(n1135) );
NAND3_X1 U949 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1248) );
XNOR2_X1 U950 ( .A(KEYINPUT20), .B(n1235), .ZN(n1251) );
NAND2_X1 U951 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
NAND2_X1 U952 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U953 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
XNOR2_X1 U954 ( .A(n1258), .B(n1259), .ZN(n1256) );
XNOR2_X1 U955 ( .A(G110), .B(n1260), .ZN(n1252) );
INV_X1 U956 ( .A(n1132), .ZN(n1260) );
NAND2_X1 U957 ( .A1(n1261), .A2(n1262), .ZN(n1249) );
NAND2_X1 U958 ( .A1(n1263), .A2(n1257), .ZN(n1262) );
INV_X1 U959 ( .A(KEYINPUT11), .ZN(n1257) );
NAND2_X1 U960 ( .A1(n1264), .A2(n1255), .ZN(n1263) );
INV_X1 U961 ( .A(KEYINPUT46), .ZN(n1255) );
XNOR2_X1 U962 ( .A(G110), .B(n1132), .ZN(n1264) );
XOR2_X1 U963 ( .A(G140), .B(n1265), .Z(n1132) );
NOR2_X1 U964 ( .A1(G953), .A2(n1069), .ZN(n1265) );
INV_X1 U965 ( .A(G227), .ZN(n1069) );
XNOR2_X1 U966 ( .A(n1259), .B(n1063), .ZN(n1261) );
INV_X1 U967 ( .A(n1258), .ZN(n1063) );
XNOR2_X1 U968 ( .A(n1115), .B(n1266), .ZN(n1258) );
INV_X1 U969 ( .A(n1127), .ZN(n1266) );
XOR2_X1 U970 ( .A(G131), .B(n1267), .Z(n1115) );
XNOR2_X1 U971 ( .A(n1225), .B(G134), .ZN(n1267) );
INV_X1 U972 ( .A(G137), .ZN(n1225) );
NOR2_X1 U973 ( .A1(KEYINPUT43), .A2(n1130), .ZN(n1259) );
XNOR2_X1 U974 ( .A(n1085), .B(KEYINPUT36), .ZN(n1130) );
AND2_X1 U975 ( .A1(n1020), .A2(n1163), .ZN(n1169) );
NOR2_X1 U976 ( .A1(n1025), .A2(n1156), .ZN(n1163) );
INV_X1 U977 ( .A(n1167), .ZN(n1156) );
NAND2_X1 U978 ( .A1(n1023), .A2(n1268), .ZN(n1167) );
NAND4_X1 U979 ( .A1(G953), .A2(G902), .A3(n1211), .A4(n1081), .ZN(n1268) );
INV_X1 U980 ( .A(G898), .ZN(n1081) );
NAND3_X1 U981 ( .A1(n1211), .A2(n1017), .A3(G952), .ZN(n1023) );
NAND2_X1 U982 ( .A1(G237), .A2(G234), .ZN(n1211) );
INV_X1 U983 ( .A(n1158), .ZN(n1025) );
NOR2_X1 U984 ( .A1(n1026), .A2(n1269), .ZN(n1158) );
INV_X1 U985 ( .A(n1028), .ZN(n1269) );
NAND2_X1 U986 ( .A1(G214), .A2(n1270), .ZN(n1028) );
XOR2_X1 U987 ( .A(n1034), .B(KEYINPUT50), .Z(n1026) );
XNOR2_X1 U988 ( .A(n1271), .B(n1141), .ZN(n1034) );
NAND2_X1 U989 ( .A1(G210), .A2(n1270), .ZN(n1141) );
NAND2_X1 U990 ( .A1(n1272), .A2(n1235), .ZN(n1270) );
NAND2_X1 U991 ( .A1(n1273), .A2(n1235), .ZN(n1271) );
XOR2_X1 U992 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U993 ( .A(n1137), .B(n1186), .ZN(n1275) );
XNOR2_X1 U994 ( .A(n1247), .B(G125), .ZN(n1186) );
XNOR2_X1 U995 ( .A(n1127), .B(KEYINPUT55), .ZN(n1247) );
XOR2_X1 U996 ( .A(G146), .B(n1276), .Z(n1127) );
XNOR2_X1 U997 ( .A(n1277), .B(n1086), .ZN(n1137) );
XNOR2_X1 U998 ( .A(n1278), .B(n1231), .ZN(n1086) );
INV_X1 U999 ( .A(G110), .ZN(n1231) );
XNOR2_X1 U1000 ( .A(n1279), .B(n1280), .ZN(n1277) );
INV_X1 U1001 ( .A(n1085), .ZN(n1280) );
XOR2_X1 U1002 ( .A(G101), .B(n1281), .Z(n1085) );
XOR2_X1 U1003 ( .A(G107), .B(G104), .Z(n1281) );
NAND2_X1 U1004 ( .A1(KEYINPUT17), .A2(n1082), .ZN(n1279) );
XOR2_X1 U1005 ( .A(n1282), .B(n1283), .Z(n1082) );
NAND2_X1 U1006 ( .A1(KEYINPUT18), .A2(n1246), .ZN(n1282) );
XOR2_X1 U1007 ( .A(G116), .B(n1229), .Z(n1246) );
XOR2_X1 U1008 ( .A(G119), .B(KEYINPUT23), .Z(n1229) );
XOR2_X1 U1009 ( .A(n1187), .B(n1284), .Z(n1274) );
XNOR2_X1 U1010 ( .A(KEYINPUT6), .B(KEYINPUT45), .ZN(n1284) );
NAND2_X1 U1011 ( .A1(G224), .A2(n1017), .ZN(n1187) );
NOR2_X1 U1012 ( .A1(n1195), .A2(n1039), .ZN(n1020) );
XOR2_X1 U1013 ( .A(n1285), .B(n1098), .Z(n1039) );
INV_X1 U1014 ( .A(G475), .ZN(n1098) );
NAND2_X1 U1015 ( .A1(n1096), .A2(n1235), .ZN(n1285) );
INV_X1 U1016 ( .A(G902), .ZN(n1235) );
XNOR2_X1 U1017 ( .A(n1286), .B(n1287), .ZN(n1096) );
XNOR2_X1 U1018 ( .A(n1288), .B(n1289), .ZN(n1287) );
XOR2_X1 U1019 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U1020 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
OR2_X1 U1021 ( .A1(n1201), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1022 ( .A(n1295), .B(KEYINPUT34), .Z(n1292) );
NAND2_X1 U1023 ( .A1(n1294), .A2(n1201), .ZN(n1295) );
INV_X1 U1024 ( .A(G131), .ZN(n1201) );
XNOR2_X1 U1025 ( .A(n1296), .B(G143), .ZN(n1294) );
NAND3_X1 U1026 ( .A1(n1272), .A2(n1017), .A3(G214), .ZN(n1296) );
INV_X1 U1027 ( .A(G237), .ZN(n1272) );
NAND2_X1 U1028 ( .A1(n1297), .A2(n1298), .ZN(n1290) );
NAND4_X1 U1029 ( .A1(KEYINPUT7), .A2(KEYINPUT1), .A3(n1283), .A4(n1278), .ZN(n1298) );
NAND2_X1 U1030 ( .A1(n1299), .A2(n1300), .ZN(n1297) );
NAND2_X1 U1031 ( .A1(n1301), .A2(n1278), .ZN(n1300) );
OR2_X1 U1032 ( .A1(n1283), .A2(KEYINPUT1), .ZN(n1301) );
NAND2_X1 U1033 ( .A1(KEYINPUT7), .A2(n1283), .ZN(n1299) );
INV_X1 U1034 ( .A(G113), .ZN(n1283) );
INV_X1 U1035 ( .A(n1224), .ZN(n1288) );
XOR2_X1 U1036 ( .A(G146), .B(n1064), .Z(n1224) );
XOR2_X1 U1037 ( .A(G125), .B(G140), .Z(n1064) );
XOR2_X1 U1038 ( .A(n1302), .B(G104), .Z(n1286) );
XNOR2_X1 U1039 ( .A(KEYINPUT53), .B(KEYINPUT37), .ZN(n1302) );
NAND3_X1 U1040 ( .A1(n1303), .A2(n1304), .A3(n1042), .ZN(n1195) );
NAND2_X1 U1041 ( .A1(n1040), .A2(n1041), .ZN(n1042) );
NAND2_X1 U1042 ( .A1(n1041), .A2(n1305), .ZN(n1304) );
OR3_X1 U1043 ( .A1(n1041), .A2(n1040), .A3(n1305), .ZN(n1303) );
INV_X1 U1044 ( .A(KEYINPUT12), .ZN(n1305) );
NOR2_X1 U1045 ( .A1(n1094), .A2(G902), .ZN(n1040) );
XNOR2_X1 U1046 ( .A(n1306), .B(n1307), .ZN(n1094) );
XOR2_X1 U1047 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1048 ( .A(G107), .B(n1310), .Z(n1309) );
NOR2_X1 U1049 ( .A1(KEYINPUT35), .A2(n1276), .ZN(n1310) );
XOR2_X1 U1050 ( .A(G128), .B(G143), .Z(n1276) );
AND3_X1 U1051 ( .A1(G234), .A2(n1017), .A3(G217), .ZN(n1308) );
INV_X1 U1052 ( .A(G953), .ZN(n1017) );
XNOR2_X1 U1053 ( .A(G116), .B(n1311), .ZN(n1306) );
XNOR2_X1 U1054 ( .A(G134), .B(n1278), .ZN(n1311) );
INV_X1 U1055 ( .A(G122), .ZN(n1278) );
INV_X1 U1056 ( .A(G478), .ZN(n1041) );
endmodule


