//Key = 1001010001001011111000100100110000101011111101000100101000001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U741 ( .A(G107), .B(n1024), .ZN(G9) );
NAND4_X1 U742 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
XNOR2_X1 U743 ( .A(n1029), .B(KEYINPUT22), .ZN(n1025) );
NOR2_X1 U744 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U745 ( .A1(n1032), .A2(n1033), .A3(G953), .A4(n1034), .ZN(n1031) );
NOR2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U748 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U751 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
XOR2_X1 U753 ( .A(n1050), .B(KEYINPUT1), .Z(n1048) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR3_X1 U757 ( .A1(n1052), .A2(n1057), .A3(n1045), .ZN(n1037) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U759 ( .A1(n1060), .A2(n1041), .ZN(n1059) );
NOR2_X1 U760 ( .A1(n1061), .A2(n1029), .ZN(n1060) );
AND2_X1 U761 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1039), .ZN(n1058) );
NOR2_X1 U763 ( .A1(n1027), .A2(n1065), .ZN(n1064) );
NAND3_X1 U764 ( .A1(n1066), .A2(G952), .A3(n1067), .ZN(n1032) );
NOR3_X1 U765 ( .A1(n1068), .A2(G953), .A3(n1034), .ZN(n1030) );
AND4_X1 U766 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1072), .ZN(n1034) );
NOR4_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1072) );
XNOR2_X1 U768 ( .A(n1077), .B(n1078), .ZN(n1076) );
XOR2_X1 U769 ( .A(KEYINPUT33), .B(n1055), .Z(n1075) );
NOR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
INV_X1 U771 ( .A(KEYINPUT35), .ZN(n1080) );
NOR3_X1 U772 ( .A1(n1081), .A2(n1063), .A3(n1082), .ZN(n1079) );
AND2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U774 ( .A1(KEYINPUT35), .A2(n1085), .ZN(n1073) );
NOR2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1071) );
INV_X1 U776 ( .A(n1049), .ZN(n1086) );
XNOR2_X1 U777 ( .A(n1088), .B(n1089), .ZN(n1070) );
NAND2_X1 U778 ( .A1(KEYINPUT14), .A2(G478), .ZN(n1088) );
XOR2_X1 U779 ( .A(n1090), .B(n1091), .Z(n1069) );
NAND2_X1 U780 ( .A1(KEYINPUT49), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U781 ( .A(G952), .B(KEYINPUT41), .ZN(n1068) );
NAND2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(G72) );
NAND3_X1 U783 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
XOR2_X1 U784 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U785 ( .A1(KEYINPUT24), .A2(n1100), .ZN(n1099) );
XOR2_X1 U786 ( .A(n1101), .B(KEYINPUT30), .Z(n1100) );
NAND2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1093) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1103) );
XOR2_X1 U789 ( .A(KEYINPUT0), .B(G953), .Z(n1095) );
XNOR2_X1 U790 ( .A(n1104), .B(n1098), .ZN(n1102) );
NAND2_X1 U791 ( .A1(G953), .A2(n1105), .ZN(n1098) );
NAND2_X1 U792 ( .A1(G900), .A2(G227), .ZN(n1105) );
NAND2_X1 U793 ( .A1(n1106), .A2(n1101), .ZN(n1104) );
NAND2_X1 U794 ( .A1(n1107), .A2(n1108), .ZN(n1101) );
NAND2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XOR2_X1 U796 ( .A(n1111), .B(n1112), .Z(n1107) );
XOR2_X1 U797 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U798 ( .A1(KEYINPUT60), .A2(n1115), .ZN(n1113) );
INV_X1 U799 ( .A(KEYINPUT24), .ZN(n1106) );
XOR2_X1 U800 ( .A(n1116), .B(n1117), .Z(G69) );
XOR2_X1 U801 ( .A(n1118), .B(n1119), .Z(n1117) );
NAND2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U803 ( .A(KEYINPUT45), .B(G953), .Z(n1120) );
NAND2_X1 U804 ( .A1(n1122), .A2(n1123), .ZN(n1118) );
XOR2_X1 U805 ( .A(n1124), .B(n1125), .Z(n1122) );
NOR3_X1 U806 ( .A1(n1126), .A2(KEYINPUT58), .A3(n1127), .ZN(n1116) );
AND2_X1 U807 ( .A1(G224), .A2(G898), .ZN(n1127) );
NOR2_X1 U808 ( .A1(n1128), .A2(n1129), .ZN(G66) );
XOR2_X1 U809 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U810 ( .A1(KEYINPUT2), .A2(n1132), .ZN(n1131) );
XOR2_X1 U811 ( .A(n1133), .B(n1134), .Z(n1132) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
NOR3_X1 U813 ( .A1(n1128), .A2(n1137), .A3(n1138), .ZN(G63) );
NOR4_X1 U814 ( .A1(n1139), .A2(n1140), .A3(KEYINPUT56), .A4(n1141), .ZN(n1138) );
INV_X1 U815 ( .A(n1142), .ZN(n1139) );
NOR2_X1 U816 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
NOR3_X1 U817 ( .A1(n1140), .A2(n1144), .A3(n1141), .ZN(n1143) );
INV_X1 U818 ( .A(G478), .ZN(n1141) );
AND2_X1 U819 ( .A1(n1145), .A2(KEYINPUT56), .ZN(n1144) );
NOR2_X1 U820 ( .A1(KEYINPUT46), .A2(n1145), .ZN(n1142) );
XNOR2_X1 U821 ( .A(n1146), .B(KEYINPUT19), .ZN(n1145) );
NOR2_X1 U822 ( .A1(n1128), .A2(n1147), .ZN(G60) );
XNOR2_X1 U823 ( .A(n1148), .B(n1149), .ZN(n1147) );
AND2_X1 U824 ( .A1(G475), .A2(n1135), .ZN(n1149) );
XOR2_X1 U825 ( .A(n1150), .B(n1151), .Z(G6) );
XOR2_X1 U826 ( .A(KEYINPUT44), .B(G104), .Z(n1151) );
NOR2_X1 U827 ( .A1(n1128), .A2(n1152), .ZN(G57) );
XOR2_X1 U828 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U829 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U830 ( .A(n1157), .B(n1158), .ZN(n1156) );
AND2_X1 U831 ( .A1(G472), .A2(n1135), .ZN(n1158) );
INV_X1 U832 ( .A(n1140), .ZN(n1135) );
XOR2_X1 U833 ( .A(KEYINPUT39), .B(n1159), .Z(n1155) );
XOR2_X1 U834 ( .A(n1160), .B(n1161), .Z(n1153) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1160) );
NOR2_X1 U836 ( .A1(n1128), .A2(n1164), .ZN(G54) );
XOR2_X1 U837 ( .A(n1165), .B(n1166), .Z(n1164) );
XNOR2_X1 U838 ( .A(n1167), .B(n1168), .ZN(n1166) );
NOR2_X1 U839 ( .A1(n1081), .A2(n1140), .ZN(n1168) );
INV_X1 U840 ( .A(G469), .ZN(n1081) );
XOR2_X1 U841 ( .A(n1169), .B(n1170), .Z(n1165) );
NOR2_X1 U842 ( .A1(KEYINPUT20), .A2(G140), .ZN(n1170) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1169) );
NOR2_X1 U844 ( .A1(n1128), .A2(n1173), .ZN(G51) );
NOR2_X1 U845 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
XOR2_X1 U846 ( .A(n1176), .B(n1177), .Z(n1175) );
AND2_X1 U847 ( .A1(n1178), .A2(KEYINPUT54), .ZN(n1177) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1140), .ZN(n1176) );
NAND2_X1 U849 ( .A1(G902), .A2(n1180), .ZN(n1140) );
NAND2_X1 U850 ( .A1(n1067), .A2(n1181), .ZN(n1180) );
XOR2_X1 U851 ( .A(KEYINPUT55), .B(n1066), .Z(n1181) );
INV_X1 U852 ( .A(n1096), .ZN(n1066) );
NAND4_X1 U853 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1096) );
NOR4_X1 U854 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
NOR2_X1 U855 ( .A1(n1052), .A2(n1190), .ZN(n1189) );
NOR2_X1 U856 ( .A1(n1191), .A2(n1192), .ZN(n1188) );
XOR2_X1 U857 ( .A(n1193), .B(KEYINPUT32), .Z(n1191) );
NAND2_X1 U858 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
INV_X1 U859 ( .A(n1196), .ZN(n1187) );
AND2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1184) );
INV_X1 U861 ( .A(n1121), .ZN(n1067) );
NAND4_X1 U862 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1121) );
NOR4_X1 U863 ( .A1(n1203), .A2(n1204), .A3(n1150), .A4(n1205), .ZN(n1202) );
NOR3_X1 U864 ( .A1(n1206), .A2(n1045), .A3(n1207), .ZN(n1205) );
AND3_X1 U865 ( .A1(n1208), .A2(n1028), .A3(n1065), .ZN(n1150) );
NOR2_X1 U866 ( .A1(n1209), .A2(n1210), .ZN(n1201) );
NOR2_X1 U867 ( .A1(KEYINPUT54), .A2(n1178), .ZN(n1174) );
XNOR2_X1 U868 ( .A(n1211), .B(n1212), .ZN(n1178) );
XOR2_X1 U869 ( .A(n1213), .B(G125), .Z(n1211) );
NOR2_X1 U870 ( .A1(n1126), .A2(G952), .ZN(n1128) );
XOR2_X1 U871 ( .A(n1214), .B(n1196), .Z(G48) );
NAND3_X1 U872 ( .A1(n1195), .A2(n1055), .A3(n1215), .ZN(n1196) );
INV_X1 U873 ( .A(n1216), .ZN(n1055) );
XNOR2_X1 U874 ( .A(n1186), .B(n1217), .ZN(G45) );
XOR2_X1 U875 ( .A(KEYINPUT36), .B(G143), .Z(n1217) );
AND3_X1 U876 ( .A1(n1047), .A2(n1218), .A3(n1219), .ZN(n1186) );
XOR2_X1 U877 ( .A(G140), .B(n1220), .Z(G42) );
NOR2_X1 U878 ( .A1(n1221), .A2(n1052), .ZN(n1220) );
XOR2_X1 U879 ( .A(n1190), .B(KEYINPUT8), .Z(n1221) );
NAND4_X1 U880 ( .A1(n1195), .A2(n1065), .A3(n1216), .A4(n1222), .ZN(n1190) );
NAND2_X1 U881 ( .A1(n1223), .A2(n1224), .ZN(G39) );
NAND2_X1 U882 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
XOR2_X1 U883 ( .A(KEYINPUT28), .B(n1227), .Z(n1223) );
NOR2_X1 U884 ( .A1(n1225), .A2(n1226), .ZN(n1227) );
INV_X1 U885 ( .A(G137), .ZN(n1226) );
INV_X1 U886 ( .A(n1183), .ZN(n1225) );
NAND3_X1 U887 ( .A1(n1228), .A2(n1229), .A3(n1195), .ZN(n1183) );
XOR2_X1 U888 ( .A(n1115), .B(n1198), .Z(G36) );
NAND3_X1 U889 ( .A1(n1228), .A2(n1027), .A3(n1219), .ZN(n1198) );
INV_X1 U890 ( .A(G134), .ZN(n1115) );
XOR2_X1 U891 ( .A(n1230), .B(n1197), .Z(G33) );
NAND3_X1 U892 ( .A1(n1228), .A2(n1065), .A3(n1219), .ZN(n1197) );
AND2_X1 U893 ( .A1(n1195), .A2(n1054), .ZN(n1219) );
AND2_X1 U894 ( .A1(n1029), .A2(n1231), .ZN(n1195) );
INV_X1 U895 ( .A(n1052), .ZN(n1228) );
NAND2_X1 U896 ( .A1(n1232), .A2(n1049), .ZN(n1052) );
INV_X1 U897 ( .A(n1050), .ZN(n1232) );
XNOR2_X1 U898 ( .A(G128), .B(n1233), .ZN(G30) );
NAND4_X1 U899 ( .A1(n1194), .A2(n1047), .A3(n1234), .A4(n1231), .ZN(n1233) );
XOR2_X1 U900 ( .A(KEYINPUT57), .B(n1029), .Z(n1234) );
NOR3_X1 U901 ( .A1(n1207), .A2(n1216), .A3(n1056), .ZN(n1194) );
XOR2_X1 U902 ( .A(G101), .B(n1204), .Z(G3) );
AND3_X1 U903 ( .A1(n1235), .A2(n1208), .A3(n1054), .ZN(n1204) );
XOR2_X1 U904 ( .A(n1236), .B(n1182), .Z(G27) );
NAND4_X1 U905 ( .A1(n1215), .A2(n1085), .A3(n1216), .A4(n1231), .ZN(n1182) );
NAND2_X1 U906 ( .A1(n1036), .A2(n1237), .ZN(n1231) );
NAND4_X1 U907 ( .A1(n1109), .A2(G902), .A3(n1238), .A4(n1110), .ZN(n1237) );
INV_X1 U908 ( .A(G900), .ZN(n1110) );
AND3_X1 U909 ( .A1(n1222), .A2(n1047), .A3(n1065), .ZN(n1215) );
XOR2_X1 U910 ( .A(G122), .B(n1203), .Z(G24) );
AND3_X1 U911 ( .A1(n1028), .A2(n1218), .A3(n1239), .ZN(n1203) );
NAND2_X1 U912 ( .A1(n1240), .A2(n1241), .ZN(n1218) );
OR2_X1 U913 ( .A1(n1207), .A2(KEYINPUT62), .ZN(n1241) );
NAND3_X1 U914 ( .A1(n1242), .A2(n1243), .A3(KEYINPUT62), .ZN(n1240) );
INV_X1 U915 ( .A(n1244), .ZN(n1243) );
INV_X1 U916 ( .A(n1045), .ZN(n1028) );
NAND2_X1 U917 ( .A1(n1216), .A2(n1056), .ZN(n1045) );
XNOR2_X1 U918 ( .A(G119), .B(n1245), .ZN(G21) );
NAND2_X1 U919 ( .A1(KEYINPUT3), .A2(n1210), .ZN(n1245) );
AND2_X1 U920 ( .A1(n1229), .A2(n1239), .ZN(n1210) );
NOR3_X1 U921 ( .A1(n1056), .A2(n1216), .A3(n1041), .ZN(n1229) );
INV_X1 U922 ( .A(n1222), .ZN(n1056) );
XOR2_X1 U923 ( .A(G116), .B(n1209), .Z(G18) );
AND3_X1 U924 ( .A1(n1239), .A2(n1027), .A3(n1054), .ZN(n1209) );
INV_X1 U925 ( .A(n1207), .ZN(n1027) );
NAND2_X1 U926 ( .A1(n1244), .A2(n1242), .ZN(n1207) );
XNOR2_X1 U927 ( .A(n1199), .B(n1246), .ZN(G15) );
XOR2_X1 U928 ( .A(KEYINPUT7), .B(G113), .Z(n1246) );
NAND3_X1 U929 ( .A1(n1065), .A2(n1239), .A3(n1054), .ZN(n1199) );
NOR2_X1 U930 ( .A1(n1222), .A2(n1216), .ZN(n1054) );
AND2_X1 U931 ( .A1(n1085), .A2(n1026), .ZN(n1239) );
INV_X1 U932 ( .A(n1039), .ZN(n1085) );
NAND2_X1 U933 ( .A1(n1062), .A2(n1247), .ZN(n1039) );
NOR2_X1 U934 ( .A1(n1242), .A2(n1244), .ZN(n1065) );
INV_X1 U935 ( .A(n1248), .ZN(n1242) );
XOR2_X1 U936 ( .A(n1171), .B(n1200), .Z(G12) );
NAND4_X1 U937 ( .A1(n1235), .A2(n1208), .A3(n1216), .A4(n1222), .ZN(n1200) );
XNOR2_X1 U938 ( .A(n1087), .B(KEYINPUT17), .ZN(n1222) );
XNOR2_X1 U939 ( .A(n1249), .B(n1136), .ZN(n1087) );
AND2_X1 U940 ( .A1(G217), .A2(n1250), .ZN(n1136) );
NAND2_X1 U941 ( .A1(n1251), .A2(n1083), .ZN(n1249) );
XOR2_X1 U942 ( .A(n1133), .B(n1252), .Z(n1251) );
INV_X1 U943 ( .A(n1134), .ZN(n1252) );
XOR2_X1 U944 ( .A(n1253), .B(n1254), .Z(n1134) );
XOR2_X1 U945 ( .A(KEYINPUT61), .B(G146), .Z(n1254) );
XOR2_X1 U946 ( .A(n1255), .B(G110), .Z(n1253) );
NAND2_X1 U947 ( .A1(G221), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U948 ( .A(n1257), .B(n1258), .ZN(n1133) );
XOR2_X1 U949 ( .A(n1163), .B(n1259), .Z(n1258) );
XOR2_X1 U950 ( .A(n1260), .B(G472), .Z(n1216) );
NAND2_X1 U951 ( .A1(n1261), .A2(n1083), .ZN(n1260) );
XOR2_X1 U952 ( .A(n1262), .B(n1161), .Z(n1261) );
XNOR2_X1 U953 ( .A(n1263), .B(n1264), .ZN(n1161) );
NAND2_X1 U954 ( .A1(KEYINPUT12), .A2(n1265), .ZN(n1263) );
XNOR2_X1 U955 ( .A(n1266), .B(n1267), .ZN(n1262) );
NOR2_X1 U956 ( .A1(KEYINPUT47), .A2(n1268), .ZN(n1267) );
XOR2_X1 U957 ( .A(G101), .B(n1269), .Z(n1268) );
NOR2_X1 U958 ( .A1(n1159), .A2(KEYINPUT37), .ZN(n1269) );
AND3_X1 U959 ( .A1(n1270), .A2(n1126), .A3(G210), .ZN(n1159) );
NOR2_X1 U960 ( .A1(KEYINPUT26), .A2(n1271), .ZN(n1266) );
XNOR2_X1 U961 ( .A(n1272), .B(n1273), .ZN(n1271) );
NOR2_X1 U962 ( .A1(KEYINPUT50), .A2(n1274), .ZN(n1273) );
XOR2_X1 U963 ( .A(n1275), .B(G137), .Z(n1274) );
INV_X1 U964 ( .A(n1206), .ZN(n1208) );
NAND2_X1 U965 ( .A1(n1026), .A2(n1029), .ZN(n1206) );
NOR2_X1 U966 ( .A1(n1062), .A2(n1063), .ZN(n1029) );
INV_X1 U967 ( .A(n1247), .ZN(n1063) );
NAND2_X1 U968 ( .A1(G221), .A2(n1250), .ZN(n1247) );
NAND2_X1 U969 ( .A1(G234), .A2(n1276), .ZN(n1250) );
XOR2_X1 U970 ( .A(KEYINPUT9), .B(G902), .Z(n1276) );
XOR2_X1 U971 ( .A(n1277), .B(G469), .Z(n1062) );
NAND2_X1 U972 ( .A1(n1083), .A2(n1084), .ZN(n1277) );
NAND3_X1 U973 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1084) );
NAND2_X1 U974 ( .A1(n1281), .A2(n1167), .ZN(n1280) );
NAND2_X1 U975 ( .A1(n1282), .A2(n1283), .ZN(n1279) );
INV_X1 U976 ( .A(KEYINPUT34), .ZN(n1283) );
NAND2_X1 U977 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
XNOR2_X1 U978 ( .A(n1167), .B(KEYINPUT4), .ZN(n1284) );
NAND2_X1 U979 ( .A1(KEYINPUT34), .A2(n1286), .ZN(n1278) );
NAND2_X1 U980 ( .A1(n1287), .A2(n1288), .ZN(n1286) );
OR3_X1 U981 ( .A1(n1281), .A2(n1167), .A3(KEYINPUT4), .ZN(n1288) );
INV_X1 U982 ( .A(n1285), .ZN(n1281) );
XOR2_X1 U983 ( .A(n1289), .B(n1172), .Z(n1285) );
AND2_X1 U984 ( .A1(G227), .A2(n1126), .ZN(n1172) );
NAND2_X1 U985 ( .A1(n1290), .A2(KEYINPUT5), .ZN(n1289) );
XOR2_X1 U986 ( .A(n1171), .B(G140), .Z(n1290) );
NAND2_X1 U987 ( .A1(KEYINPUT4), .A2(n1167), .ZN(n1287) );
XNOR2_X1 U988 ( .A(n1291), .B(n1292), .ZN(n1167) );
INV_X1 U989 ( .A(n1114), .ZN(n1292) );
XOR2_X1 U990 ( .A(n1293), .B(n1163), .Z(n1114) );
XOR2_X1 U991 ( .A(G128), .B(G137), .Z(n1163) );
NAND2_X1 U992 ( .A1(KEYINPUT40), .A2(n1294), .ZN(n1293) );
INV_X1 U993 ( .A(n1295), .ZN(n1294) );
XOR2_X1 U994 ( .A(n1162), .B(n1296), .Z(n1291) );
XOR2_X1 U995 ( .A(n1275), .B(G101), .Z(n1162) );
XOR2_X1 U996 ( .A(n1230), .B(n1297), .Z(n1275) );
XOR2_X1 U997 ( .A(KEYINPUT27), .B(G134), .Z(n1297) );
INV_X1 U998 ( .A(G131), .ZN(n1230) );
AND2_X1 U999 ( .A1(n1047), .A2(n1298), .ZN(n1026) );
NAND2_X1 U1000 ( .A1(n1036), .A2(n1299), .ZN(n1298) );
NAND3_X1 U1001 ( .A1(n1300), .A2(n1238), .A3(G902), .ZN(n1299) );
INV_X1 U1002 ( .A(n1123), .ZN(n1300) );
NAND2_X1 U1003 ( .A1(n1109), .A2(n1301), .ZN(n1123) );
INV_X1 U1004 ( .A(G898), .ZN(n1301) );
XOR2_X1 U1005 ( .A(n1126), .B(KEYINPUT18), .Z(n1109) );
NAND3_X1 U1006 ( .A1(n1238), .A2(n1126), .A3(G952), .ZN(n1036) );
NAND2_X1 U1007 ( .A1(G234), .A2(G237), .ZN(n1238) );
INV_X1 U1008 ( .A(n1192), .ZN(n1047) );
NAND2_X1 U1009 ( .A1(n1050), .A2(n1049), .ZN(n1192) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1302), .ZN(n1049) );
XNOR2_X1 U1011 ( .A(n1092), .B(n1303), .ZN(n1050) );
NOR2_X1 U1012 ( .A1(n1091), .A2(KEYINPUT6), .ZN(n1303) );
INV_X1 U1013 ( .A(n1179), .ZN(n1091) );
NAND2_X1 U1014 ( .A1(G210), .A2(n1302), .ZN(n1179) );
NAND2_X1 U1015 ( .A1(n1304), .A2(n1083), .ZN(n1302) );
XOR2_X1 U1016 ( .A(KEYINPUT43), .B(G237), .Z(n1304) );
AND3_X1 U1017 ( .A1(n1305), .A2(n1306), .A3(n1083), .ZN(n1092) );
NAND2_X1 U1018 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XNOR2_X1 U1019 ( .A(n1212), .B(KEYINPUT59), .ZN(n1308) );
NAND2_X1 U1020 ( .A1(n1212), .A2(n1309), .ZN(n1305) );
INV_X1 U1021 ( .A(n1307), .ZN(n1309) );
XOR2_X1 U1022 ( .A(n1310), .B(KEYINPUT13), .Z(n1307) );
NAND2_X1 U1023 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND2_X1 U1024 ( .A1(n1213), .A2(n1236), .ZN(n1312) );
INV_X1 U1025 ( .A(G125), .ZN(n1236) );
NAND2_X1 U1026 ( .A1(n1313), .A2(G125), .ZN(n1311) );
XOR2_X1 U1027 ( .A(KEYINPUT48), .B(n1314), .Z(n1313) );
INV_X1 U1028 ( .A(n1213), .ZN(n1314) );
XOR2_X1 U1029 ( .A(n1315), .B(n1272), .Z(n1213) );
XNOR2_X1 U1030 ( .A(n1157), .B(G128), .ZN(n1272) );
NAND2_X1 U1031 ( .A1(KEYINPUT38), .A2(n1295), .ZN(n1157) );
NAND2_X1 U1032 ( .A1(G224), .A2(n1126), .ZN(n1315) );
XNOR2_X1 U1033 ( .A(n1316), .B(n1125), .ZN(n1212) );
XNOR2_X1 U1034 ( .A(n1317), .B(n1318), .ZN(n1125) );
XOR2_X1 U1035 ( .A(G122), .B(G101), .Z(n1318) );
XNOR2_X1 U1036 ( .A(n1319), .B(n1320), .ZN(n1317) );
NOR2_X1 U1037 ( .A1(G110), .A2(KEYINPUT23), .ZN(n1320) );
NOR2_X1 U1038 ( .A1(KEYINPUT11), .A2(n1296), .ZN(n1319) );
XOR2_X1 U1039 ( .A(G104), .B(n1321), .Z(n1296) );
NAND2_X1 U1040 ( .A1(KEYINPUT29), .A2(n1124), .ZN(n1316) );
NAND2_X1 U1041 ( .A1(n1322), .A2(n1323), .ZN(n1124) );
NAND2_X1 U1042 ( .A1(n1265), .A2(n1264), .ZN(n1323) );
XOR2_X1 U1043 ( .A(KEYINPUT25), .B(n1324), .Z(n1322) );
NOR2_X1 U1044 ( .A1(n1265), .A2(n1264), .ZN(n1324) );
XOR2_X1 U1045 ( .A(G116), .B(n1257), .Z(n1265) );
XOR2_X1 U1046 ( .A(G119), .B(KEYINPUT53), .Z(n1257) );
INV_X1 U1047 ( .A(n1041), .ZN(n1235) );
NAND2_X1 U1048 ( .A1(n1248), .A2(n1244), .ZN(n1041) );
XNOR2_X1 U1049 ( .A(n1325), .B(n1078), .ZN(n1244) );
XNOR2_X1 U1050 ( .A(G475), .B(KEYINPUT10), .ZN(n1078) );
NAND2_X1 U1051 ( .A1(KEYINPUT42), .A2(n1077), .ZN(n1325) );
AND2_X1 U1052 ( .A1(n1326), .A2(n1148), .ZN(n1077) );
XNOR2_X1 U1053 ( .A(n1327), .B(n1328), .ZN(n1148) );
XOR2_X1 U1054 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1055 ( .A(n1331), .B(G122), .Z(n1330) );
INV_X1 U1056 ( .A(G104), .ZN(n1331) );
NAND4_X1 U1057 ( .A1(KEYINPUT52), .A2(G214), .A3(n1270), .A4(n1126), .ZN(n1329) );
INV_X1 U1058 ( .A(G237), .ZN(n1270) );
XOR2_X1 U1059 ( .A(n1332), .B(n1111), .Z(n1327) );
XOR2_X1 U1060 ( .A(G131), .B(n1259), .Z(n1111) );
XOR2_X1 U1061 ( .A(G125), .B(G140), .Z(n1259) );
XOR2_X1 U1062 ( .A(n1295), .B(n1264), .Z(n1332) );
XOR2_X1 U1063 ( .A(G113), .B(KEYINPUT51), .Z(n1264) );
XOR2_X1 U1064 ( .A(n1214), .B(n1333), .Z(n1295) );
INV_X1 U1065 ( .A(G146), .ZN(n1214) );
XOR2_X1 U1066 ( .A(KEYINPUT16), .B(G902), .Z(n1326) );
XOR2_X1 U1067 ( .A(n1089), .B(n1334), .Z(n1248) );
XOR2_X1 U1068 ( .A(KEYINPUT31), .B(G478), .Z(n1334) );
NAND2_X1 U1069 ( .A1(n1146), .A2(n1083), .ZN(n1089) );
INV_X1 U1070 ( .A(G902), .ZN(n1083) );
XOR2_X1 U1071 ( .A(n1335), .B(n1336), .Z(n1146) );
XOR2_X1 U1072 ( .A(G116), .B(n1337), .Z(n1336) );
XOR2_X1 U1073 ( .A(G134), .B(G122), .Z(n1337) );
XOR2_X1 U1074 ( .A(n1338), .B(n1321), .Z(n1335) );
XOR2_X1 U1075 ( .A(G107), .B(KEYINPUT63), .Z(n1321) );
XOR2_X1 U1076 ( .A(n1339), .B(n1340), .Z(n1338) );
AND2_X1 U1077 ( .A1(n1256), .A2(G217), .ZN(n1340) );
AND2_X1 U1078 ( .A1(G234), .A2(n1126), .ZN(n1256) );
INV_X1 U1079 ( .A(G953), .ZN(n1126) );
NAND2_X1 U1080 ( .A1(n1341), .A2(KEYINPUT15), .ZN(n1339) );
XNOR2_X1 U1081 ( .A(G128), .B(n1333), .ZN(n1341) );
XOR2_X1 U1082 ( .A(G143), .B(KEYINPUT21), .Z(n1333) );
INV_X1 U1083 ( .A(G110), .ZN(n1171) );
endmodule


