//Key = 1001111101011001100001010000100011110100111100000010010100000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459;

XNOR2_X1 U781 ( .A(G107), .B(n1102), .ZN(G9) );
NOR2_X1 U782 ( .A1(n1103), .A2(n1104), .ZN(G75) );
NOR4_X1 U783 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1104) );
NOR2_X1 U784 ( .A1(KEYINPUT23), .A2(n1109), .ZN(n1108) );
AND3_X1 U785 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NOR3_X1 U786 ( .A1(n1111), .A2(n1113), .A3(n1114), .ZN(n1107) );
NOR2_X1 U787 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U788 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NOR2_X1 U789 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NOR3_X1 U790 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
XNOR2_X1 U791 ( .A(KEYINPUT34), .B(n1124), .ZN(n1121) );
NOR4_X1 U792 ( .A1(KEYINPUT50), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1119) );
INV_X1 U793 ( .A(n1128), .ZN(n1126) );
INV_X1 U794 ( .A(n1124), .ZN(n1125) );
NOR3_X1 U795 ( .A1(n1124), .A2(n1129), .A3(n1127), .ZN(n1115) );
NOR2_X1 U796 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U797 ( .A1(n1132), .A2(n1123), .ZN(n1131) );
NOR2_X1 U798 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U799 ( .A1(n1135), .A2(n1118), .ZN(n1130) );
NOR2_X1 U800 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
AND2_X1 U801 ( .A1(n1128), .A2(KEYINPUT50), .ZN(n1136) );
NAND3_X1 U802 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1105) );
NAND4_X1 U803 ( .A1(n1110), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1140) );
NAND3_X1 U804 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1143) );
NAND2_X1 U805 ( .A1(n1147), .A2(n1148), .ZN(n1144) );
NAND2_X1 U806 ( .A1(n1149), .A2(n1111), .ZN(n1142) );
NAND2_X1 U807 ( .A1(KEYINPUT23), .A2(n1112), .ZN(n1149) );
NAND2_X1 U808 ( .A1(n1113), .A2(n1127), .ZN(n1141) );
NOR3_X1 U809 ( .A1(n1123), .A2(n1118), .A3(n1124), .ZN(n1110) );
INV_X1 U810 ( .A(n1150), .ZN(n1123) );
AND3_X1 U811 ( .A1(n1138), .A2(n1139), .A3(n1151), .ZN(n1103) );
NAND4_X1 U812 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1138) );
NOR4_X1 U813 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
XOR2_X1 U814 ( .A(KEYINPUT0), .B(n1160), .Z(n1159) );
NOR2_X1 U815 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U816 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U817 ( .A1(G902), .A2(n1165), .ZN(n1163) );
AND2_X1 U818 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
INV_X1 U819 ( .A(n1112), .ZN(n1158) );
XOR2_X1 U820 ( .A(n1168), .B(KEYINPUT12), .Z(n1157) );
NAND2_X1 U821 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U822 ( .A1(n1170), .A2(n1169), .ZN(n1156) );
XNOR2_X1 U823 ( .A(n1171), .B(KEYINPUT58), .ZN(n1169) );
INV_X1 U824 ( .A(n1172), .ZN(n1170) );
XNOR2_X1 U825 ( .A(n1173), .B(n1174), .ZN(n1154) );
XNOR2_X1 U826 ( .A(n1175), .B(G478), .ZN(n1153) );
XNOR2_X1 U827 ( .A(n1176), .B(G472), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1177), .B(n1178), .Z(G72) );
XOR2_X1 U829 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U830 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U831 ( .A(n1183), .B(n1184), .Z(n1182) );
XNOR2_X1 U832 ( .A(n1185), .B(n1186), .ZN(n1184) );
XOR2_X1 U833 ( .A(n1187), .B(n1188), .Z(n1183) );
XNOR2_X1 U834 ( .A(KEYINPUT44), .B(KEYINPUT39), .ZN(n1187) );
NOR2_X1 U835 ( .A1(G953), .A2(n1189), .ZN(n1179) );
NOR2_X1 U836 ( .A1(n1190), .A2(n1191), .ZN(n1177) );
AND2_X1 U837 ( .A1(G227), .A2(G900), .ZN(n1190) );
XOR2_X1 U838 ( .A(n1192), .B(n1193), .Z(G69) );
XOR2_X1 U839 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U840 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
XOR2_X1 U841 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U842 ( .A(G113), .B(n1200), .ZN(n1199) );
NAND2_X1 U843 ( .A1(n1201), .A2(KEYINPUT55), .ZN(n1200) );
XOR2_X1 U844 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U845 ( .A1(G898), .A2(n1139), .ZN(n1196) );
NAND2_X1 U846 ( .A1(n1204), .A2(n1139), .ZN(n1194) );
NAND2_X1 U847 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XNOR2_X1 U848 ( .A(n1207), .B(KEYINPUT17), .ZN(n1205) );
NAND2_X1 U849 ( .A1(n1208), .A2(n1209), .ZN(n1192) );
NAND2_X1 U850 ( .A1(G898), .A2(G224), .ZN(n1209) );
INV_X1 U851 ( .A(n1191), .ZN(n1208) );
XOR2_X1 U852 ( .A(G953), .B(KEYINPUT35), .Z(n1191) );
NOR2_X1 U853 ( .A1(n1210), .A2(n1211), .ZN(G66) );
XOR2_X1 U854 ( .A(n1212), .B(n1167), .Z(n1211) );
NOR2_X1 U855 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
XNOR2_X1 U856 ( .A(KEYINPUT6), .B(n1164), .ZN(n1214) );
NOR2_X1 U857 ( .A1(n1210), .A2(n1215), .ZN(G63) );
NOR3_X1 U858 ( .A1(n1175), .A2(n1216), .A3(n1217), .ZN(n1215) );
NOR3_X1 U859 ( .A1(n1218), .A2(n1219), .A3(n1213), .ZN(n1217) );
NOR2_X1 U860 ( .A1(n1220), .A2(n1221), .ZN(n1216) );
NOR2_X1 U861 ( .A1(n1222), .A2(n1219), .ZN(n1220) );
NOR2_X1 U862 ( .A1(n1210), .A2(n1223), .ZN(G60) );
NOR3_X1 U863 ( .A1(n1172), .A2(n1224), .A3(n1225), .ZN(n1223) );
NOR3_X1 U864 ( .A1(n1226), .A2(n1171), .A3(n1213), .ZN(n1225) );
NOR2_X1 U865 ( .A1(n1227), .A2(n1228), .ZN(n1224) );
NOR2_X1 U866 ( .A1(n1222), .A2(n1171), .ZN(n1227) );
INV_X1 U867 ( .A(n1106), .ZN(n1222) );
XNOR2_X1 U868 ( .A(G104), .B(n1229), .ZN(G6) );
NAND2_X1 U869 ( .A1(n1137), .A2(n1230), .ZN(n1229) );
NOR3_X1 U870 ( .A1(n1210), .A2(n1231), .A3(n1232), .ZN(G57) );
NOR2_X1 U871 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XNOR2_X1 U872 ( .A(n1235), .B(KEYINPUT63), .ZN(n1234) );
INV_X1 U873 ( .A(n1236), .ZN(n1233) );
NOR2_X1 U874 ( .A1(n1236), .A2(n1237), .ZN(n1231) );
XNOR2_X1 U875 ( .A(KEYINPUT47), .B(n1238), .ZN(n1237) );
INV_X1 U876 ( .A(n1235), .ZN(n1238) );
XNOR2_X1 U877 ( .A(n1239), .B(n1240), .ZN(n1235) );
NOR2_X1 U878 ( .A1(n1241), .A2(n1213), .ZN(n1240) );
XNOR2_X1 U879 ( .A(n1242), .B(n1243), .ZN(n1239) );
NAND2_X1 U880 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
XOR2_X1 U881 ( .A(n1246), .B(KEYINPUT25), .Z(n1244) );
NOR2_X1 U882 ( .A1(n1210), .A2(n1247), .ZN(G54) );
XOR2_X1 U883 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U884 ( .A(n1250), .B(n1251), .ZN(n1249) );
NAND2_X1 U885 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
OR2_X1 U886 ( .A1(n1254), .A2(KEYINPUT31), .ZN(n1253) );
NAND3_X1 U887 ( .A1(G140), .A2(n1255), .A3(KEYINPUT31), .ZN(n1252) );
XNOR2_X1 U888 ( .A(n1256), .B(n1257), .ZN(n1248) );
XOR2_X1 U889 ( .A(n1258), .B(n1259), .Z(n1256) );
NOR2_X1 U890 ( .A1(n1174), .A2(n1213), .ZN(n1259) );
INV_X1 U891 ( .A(G469), .ZN(n1174) );
NOR3_X1 U892 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(G51) );
NOR3_X1 U893 ( .A1(n1263), .A2(n1139), .A3(n1151), .ZN(n1262) );
INV_X1 U894 ( .A(G952), .ZN(n1151) );
AND2_X1 U895 ( .A1(n1263), .A2(n1210), .ZN(n1261) );
NOR2_X1 U896 ( .A1(n1139), .A2(G952), .ZN(n1210) );
INV_X1 U897 ( .A(KEYINPUT46), .ZN(n1263) );
XOR2_X1 U898 ( .A(n1264), .B(n1265), .Z(n1260) );
XOR2_X1 U899 ( .A(n1266), .B(n1267), .Z(n1265) );
NOR2_X1 U900 ( .A1(n1268), .A2(n1213), .ZN(n1267) );
NAND2_X1 U901 ( .A1(G902), .A2(n1106), .ZN(n1213) );
NAND3_X1 U902 ( .A1(n1206), .A2(n1269), .A3(n1189), .ZN(n1106) );
AND4_X1 U903 ( .A1(n1270), .A2(n1271), .A3(n1272), .A4(n1273), .ZN(n1189) );
AND4_X1 U904 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1273) );
NOR3_X1 U905 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1272) );
AND2_X1 U906 ( .A1(KEYINPUT43), .A2(n1281), .ZN(n1280) );
NOR3_X1 U907 ( .A1(KEYINPUT43), .A2(n1134), .A3(n1282), .ZN(n1279) );
AND4_X1 U908 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1206) );
AND4_X1 U909 ( .A1(n1102), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n1286) );
NAND2_X1 U910 ( .A1(n1128), .A2(n1230), .ZN(n1102) );
NOR2_X1 U911 ( .A1(n1290), .A2(n1118), .ZN(n1230) );
NAND4_X1 U912 ( .A1(n1137), .A2(n1291), .A3(n1292), .A4(n1293), .ZN(n1285) );
NAND2_X1 U913 ( .A1(KEYINPUT53), .A2(n1290), .ZN(n1293) );
NAND2_X1 U914 ( .A1(n1294), .A2(n1295), .ZN(n1292) );
INV_X1 U915 ( .A(KEYINPUT53), .ZN(n1295) );
NAND2_X1 U916 ( .A1(n1296), .A2(n1297), .ZN(n1294) );
INV_X1 U917 ( .A(n1298), .ZN(n1296) );
NOR2_X1 U918 ( .A1(KEYINPUT26), .A2(n1299), .ZN(n1266) );
XOR2_X1 U919 ( .A(n1300), .B(n1301), .Z(n1264) );
NOR2_X1 U920 ( .A1(KEYINPUT60), .A2(n1302), .ZN(n1301) );
XNOR2_X1 U921 ( .A(n1303), .B(n1304), .ZN(n1302) );
XNOR2_X1 U922 ( .A(G125), .B(KEYINPUT42), .ZN(n1303) );
XNOR2_X1 U923 ( .A(G146), .B(n1270), .ZN(G48) );
NAND3_X1 U924 ( .A1(n1305), .A2(n1306), .A3(n1137), .ZN(n1270) );
XNOR2_X1 U925 ( .A(G143), .B(n1307), .ZN(G45) );
NAND2_X1 U926 ( .A1(KEYINPUT21), .A2(n1278), .ZN(n1307) );
AND4_X1 U927 ( .A1(n1305), .A2(n1133), .A3(n1308), .A4(n1309), .ZN(n1278) );
XNOR2_X1 U928 ( .A(G140), .B(n1271), .ZN(G42) );
NAND3_X1 U929 ( .A1(n1310), .A2(n1134), .A3(n1137), .ZN(n1271) );
XOR2_X1 U930 ( .A(G137), .B(n1311), .Z(G39) );
NOR2_X1 U931 ( .A1(KEYINPUT22), .A2(n1277), .ZN(n1311) );
NAND3_X1 U932 ( .A1(n1150), .A2(n1306), .A3(n1310), .ZN(n1277) );
XOR2_X1 U933 ( .A(n1312), .B(G134), .Z(G36) );
NAND2_X1 U934 ( .A1(KEYINPUT5), .A2(n1276), .ZN(n1312) );
NAND3_X1 U935 ( .A1(n1133), .A2(n1128), .A3(n1310), .ZN(n1276) );
XNOR2_X1 U936 ( .A(G131), .B(n1275), .ZN(G33) );
NAND3_X1 U937 ( .A1(n1310), .A2(n1133), .A3(n1137), .ZN(n1275) );
AND3_X1 U938 ( .A1(n1313), .A2(n1111), .A3(n1112), .ZN(n1310) );
NOR2_X1 U939 ( .A1(n1127), .A2(n1113), .ZN(n1112) );
NAND2_X1 U940 ( .A1(n1148), .A2(n1314), .ZN(n1127) );
INV_X1 U941 ( .A(n1147), .ZN(n1314) );
XOR2_X1 U942 ( .A(n1274), .B(n1315), .Z(G30) );
XNOR2_X1 U943 ( .A(G128), .B(KEYINPUT57), .ZN(n1315) );
NAND3_X1 U944 ( .A1(n1128), .A2(n1306), .A3(n1305), .ZN(n1274) );
AND2_X1 U945 ( .A1(n1297), .A2(n1313), .ZN(n1305) );
XNOR2_X1 U946 ( .A(G101), .B(n1316), .ZN(G3) );
NAND2_X1 U947 ( .A1(KEYINPUT40), .A2(n1207), .ZN(n1316) );
INV_X1 U948 ( .A(n1269), .ZN(n1207) );
NAND3_X1 U949 ( .A1(n1133), .A2(n1317), .A3(n1150), .ZN(n1269) );
XNOR2_X1 U950 ( .A(n1318), .B(n1281), .ZN(G27) );
NOR2_X1 U951 ( .A1(n1282), .A2(n1319), .ZN(n1281) );
NAND4_X1 U952 ( .A1(n1146), .A2(n1137), .A3(n1320), .A4(n1313), .ZN(n1282) );
NAND2_X1 U953 ( .A1(n1124), .A2(n1321), .ZN(n1313) );
NAND3_X1 U954 ( .A1(G902), .A2(n1322), .A3(n1181), .ZN(n1321) );
NOR2_X1 U955 ( .A1(n1139), .A2(G900), .ZN(n1181) );
XNOR2_X1 U956 ( .A(G122), .B(n1283), .ZN(G24) );
NAND4_X1 U957 ( .A1(n1323), .A2(n1291), .A3(n1308), .A4(n1309), .ZN(n1283) );
INV_X1 U958 ( .A(n1118), .ZN(n1291) );
NAND2_X1 U959 ( .A1(n1324), .A2(n1325), .ZN(n1118) );
XNOR2_X1 U960 ( .A(G119), .B(n1284), .ZN(G21) );
NAND3_X1 U961 ( .A1(n1150), .A2(n1306), .A3(n1323), .ZN(n1284) );
NAND2_X1 U962 ( .A1(n1326), .A2(n1327), .ZN(n1306) );
OR3_X1 U963 ( .A1(n1325), .A2(n1324), .A3(KEYINPUT19), .ZN(n1327) );
NAND2_X1 U964 ( .A1(KEYINPUT19), .A2(n1134), .ZN(n1326) );
XNOR2_X1 U965 ( .A(G116), .B(n1289), .ZN(G18) );
NAND3_X1 U966 ( .A1(n1133), .A2(n1128), .A3(n1323), .ZN(n1289) );
NOR2_X1 U967 ( .A1(n1328), .A2(n1309), .ZN(n1128) );
XOR2_X1 U968 ( .A(n1288), .B(n1329), .Z(G15) );
NAND2_X1 U969 ( .A1(KEYINPUT62), .A2(G113), .ZN(n1329) );
NAND3_X1 U970 ( .A1(n1137), .A2(n1133), .A3(n1323), .ZN(n1288) );
AND3_X1 U971 ( .A1(n1320), .A2(n1298), .A3(n1146), .ZN(n1323) );
INV_X1 U972 ( .A(n1111), .ZN(n1146) );
AND2_X1 U973 ( .A1(n1324), .A2(n1330), .ZN(n1133) );
XNOR2_X1 U974 ( .A(KEYINPUT19), .B(n1325), .ZN(n1330) );
INV_X1 U975 ( .A(n1331), .ZN(n1324) );
AND2_X1 U976 ( .A1(n1309), .A2(n1328), .ZN(n1137) );
XNOR2_X1 U977 ( .A(G110), .B(n1287), .ZN(G12) );
NAND3_X1 U978 ( .A1(n1150), .A2(n1317), .A3(n1134), .ZN(n1287) );
INV_X1 U979 ( .A(n1319), .ZN(n1134) );
NAND2_X1 U980 ( .A1(n1325), .A2(n1331), .ZN(n1319) );
NAND3_X1 U981 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1331) );
XOR2_X1 U982 ( .A(KEYINPUT3), .B(n1161), .Z(n1334) );
NOR3_X1 U983 ( .A1(n1335), .A2(G902), .A3(n1167), .ZN(n1161) );
NAND2_X1 U984 ( .A1(n1335), .A2(n1167), .ZN(n1333) );
XNOR2_X1 U985 ( .A(n1336), .B(n1337), .ZN(n1167) );
XOR2_X1 U986 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U987 ( .A(n1340), .B(n1341), .Z(n1339) );
NAND3_X1 U988 ( .A1(G234), .A2(n1139), .A3(G221), .ZN(n1341) );
NAND2_X1 U989 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
OR2_X1 U990 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
XOR2_X1 U991 ( .A(n1346), .B(KEYINPUT10), .Z(n1342) );
NAND2_X1 U992 ( .A1(n1345), .A2(n1344), .ZN(n1346) );
NOR2_X1 U993 ( .A1(G137), .A2(KEYINPUT56), .ZN(n1338) );
XOR2_X1 U994 ( .A(n1347), .B(n1348), .Z(n1336) );
XNOR2_X1 U995 ( .A(G110), .B(n1349), .ZN(n1348) );
NAND2_X1 U996 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NAND2_X1 U997 ( .A1(G140), .A2(n1318), .ZN(n1351) );
XOR2_X1 U998 ( .A(n1352), .B(KEYINPUT1), .Z(n1350) );
NAND2_X1 U999 ( .A1(G125), .A2(n1353), .ZN(n1352) );
INV_X1 U1000 ( .A(G140), .ZN(n1353) );
XNOR2_X1 U1001 ( .A(G146), .B(KEYINPUT54), .ZN(n1347) );
NOR2_X1 U1002 ( .A1(n1164), .A2(G234), .ZN(n1335) );
NAND2_X1 U1003 ( .A1(G902), .A2(G217), .ZN(n1332) );
NAND2_X1 U1004 ( .A1(n1354), .A2(n1355), .ZN(n1325) );
NAND2_X1 U1005 ( .A1(n1176), .A2(n1356), .ZN(n1355) );
NAND2_X1 U1006 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
NAND2_X1 U1007 ( .A1(G472), .A2(n1359), .ZN(n1358) );
INV_X1 U1008 ( .A(n1360), .ZN(n1176) );
NAND2_X1 U1009 ( .A1(n1361), .A2(n1241), .ZN(n1354) );
INV_X1 U1010 ( .A(G472), .ZN(n1241) );
NAND2_X1 U1011 ( .A1(n1359), .A2(n1362), .ZN(n1361) );
NAND2_X1 U1012 ( .A1(n1360), .A2(n1357), .ZN(n1362) );
INV_X1 U1013 ( .A(KEYINPUT59), .ZN(n1357) );
NAND2_X1 U1014 ( .A1(n1363), .A2(n1364), .ZN(n1360) );
XOR2_X1 U1015 ( .A(n1365), .B(n1366), .Z(n1363) );
XNOR2_X1 U1016 ( .A(n1236), .B(G101), .ZN(n1366) );
NOR3_X1 U1017 ( .A1(G237), .A2(G953), .A3(n1268), .ZN(n1236) );
INV_X1 U1018 ( .A(G210), .ZN(n1268) );
NAND3_X1 U1019 ( .A1(n1246), .A2(n1245), .A3(KEYINPUT32), .ZN(n1365) );
NAND2_X1 U1020 ( .A1(n1367), .A2(n1368), .ZN(n1245) );
XNOR2_X1 U1021 ( .A(n1369), .B(n1370), .ZN(n1368) );
XNOR2_X1 U1022 ( .A(n1304), .B(n1371), .ZN(n1367) );
NAND2_X1 U1023 ( .A1(n1372), .A2(n1373), .ZN(n1246) );
XOR2_X1 U1024 ( .A(n1369), .B(n1370), .Z(n1373) );
NAND2_X1 U1025 ( .A1(KEYINPUT41), .A2(n1374), .ZN(n1369) );
INV_X1 U1026 ( .A(G113), .ZN(n1374) );
XNOR2_X1 U1027 ( .A(n1375), .B(n1371), .ZN(n1372) );
INV_X1 U1028 ( .A(KEYINPUT20), .ZN(n1359) );
INV_X1 U1029 ( .A(n1290), .ZN(n1317) );
NAND2_X1 U1030 ( .A1(n1297), .A2(n1298), .ZN(n1290) );
NAND2_X1 U1031 ( .A1(n1124), .A2(n1376), .ZN(n1298) );
NAND4_X1 U1032 ( .A1(G953), .A2(G902), .A3(n1322), .A4(n1377), .ZN(n1376) );
INV_X1 U1033 ( .A(G898), .ZN(n1377) );
NAND3_X1 U1034 ( .A1(n1322), .A2(n1139), .A3(G952), .ZN(n1124) );
NAND2_X1 U1035 ( .A1(G237), .A2(G234), .ZN(n1322) );
AND2_X1 U1036 ( .A1(n1320), .A2(n1111), .ZN(n1297) );
NAND2_X1 U1037 ( .A1(n1378), .A2(n1379), .ZN(n1111) );
NAND2_X1 U1038 ( .A1(G469), .A2(n1173), .ZN(n1379) );
XOR2_X1 U1039 ( .A(n1380), .B(KEYINPUT36), .Z(n1378) );
OR2_X1 U1040 ( .A1(n1173), .A2(G469), .ZN(n1380) );
NAND2_X1 U1041 ( .A1(n1381), .A2(n1364), .ZN(n1173) );
XOR2_X1 U1042 ( .A(n1254), .B(n1382), .Z(n1381) );
XNOR2_X1 U1043 ( .A(n1258), .B(n1383), .ZN(n1382) );
NOR3_X1 U1044 ( .A1(n1384), .A2(KEYINPUT24), .A3(n1385), .ZN(n1383) );
NOR3_X1 U1045 ( .A1(n1251), .A2(n1386), .A3(n1387), .ZN(n1385) );
NOR2_X1 U1046 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NOR2_X1 U1047 ( .A1(KEYINPUT61), .A2(n1257), .ZN(n1386) );
XOR2_X1 U1048 ( .A(n1390), .B(KEYINPUT4), .Z(n1384) );
NAND3_X1 U1049 ( .A1(n1391), .A2(n1392), .A3(n1251), .ZN(n1390) );
INV_X1 U1050 ( .A(n1371), .ZN(n1251) );
XOR2_X1 U1051 ( .A(n1188), .B(KEYINPUT9), .Z(n1371) );
XNOR2_X1 U1052 ( .A(n1393), .B(n1394), .ZN(n1188) );
XNOR2_X1 U1053 ( .A(G134), .B(G137), .ZN(n1393) );
NAND2_X1 U1054 ( .A1(KEYINPUT61), .A2(n1388), .ZN(n1392) );
NAND2_X1 U1055 ( .A1(n1257), .A2(n1389), .ZN(n1391) );
INV_X1 U1056 ( .A(KEYINPUT61), .ZN(n1389) );
NAND2_X1 U1057 ( .A1(n1388), .A2(n1395), .ZN(n1257) );
NAND2_X1 U1058 ( .A1(n1396), .A2(n1186), .ZN(n1395) );
OR2_X1 U1059 ( .A1(n1186), .A2(n1396), .ZN(n1388) );
XOR2_X1 U1060 ( .A(G101), .B(n1397), .Z(n1396) );
NOR2_X1 U1061 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
NOR2_X1 U1062 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
INV_X1 U1063 ( .A(KEYINPUT14), .ZN(n1400) );
NOR2_X1 U1064 ( .A1(KEYINPUT14), .A2(n1402), .ZN(n1398) );
XNOR2_X1 U1065 ( .A(n1403), .B(n1404), .ZN(n1186) );
NOR3_X1 U1066 ( .A1(KEYINPUT27), .A2(n1405), .A3(n1406), .ZN(n1404) );
AND2_X1 U1067 ( .A1(KEYINPUT16), .A2(n1407), .ZN(n1406) );
NOR2_X1 U1068 ( .A1(KEYINPUT16), .A2(n1408), .ZN(n1405) );
NOR2_X1 U1069 ( .A1(G146), .A2(n1409), .ZN(n1408) );
NAND2_X1 U1070 ( .A1(G227), .A2(n1139), .ZN(n1258) );
XOR2_X1 U1071 ( .A(G110), .B(G140), .Z(n1254) );
NOR2_X1 U1072 ( .A1(n1122), .A2(n1113), .ZN(n1320) );
INV_X1 U1073 ( .A(n1145), .ZN(n1113) );
NAND2_X1 U1074 ( .A1(G221), .A2(n1410), .ZN(n1145) );
NAND2_X1 U1075 ( .A1(G234), .A2(n1364), .ZN(n1410) );
OR2_X1 U1076 ( .A1(n1148), .A2(n1147), .ZN(n1122) );
NOR2_X1 U1077 ( .A1(n1411), .A2(n1412), .ZN(n1147) );
XOR2_X1 U1078 ( .A(n1413), .B(n1414), .Z(n1148) );
NOR2_X1 U1079 ( .A1(n1412), .A2(n1415), .ZN(n1414) );
XNOR2_X1 U1080 ( .A(G210), .B(KEYINPUT38), .ZN(n1415) );
NOR2_X1 U1081 ( .A1(G902), .A2(G237), .ZN(n1412) );
NAND2_X1 U1082 ( .A1(n1416), .A2(n1364), .ZN(n1413) );
INV_X1 U1083 ( .A(G902), .ZN(n1364) );
XNOR2_X1 U1084 ( .A(n1299), .B(n1417), .ZN(n1416) );
XOR2_X1 U1085 ( .A(n1418), .B(n1300), .Z(n1417) );
NAND2_X1 U1086 ( .A1(G224), .A2(n1139), .ZN(n1300) );
INV_X1 U1087 ( .A(G953), .ZN(n1139) );
NAND4_X1 U1088 ( .A1(KEYINPUT7), .A2(n1419), .A3(n1420), .A4(n1421), .ZN(n1418) );
NAND3_X1 U1089 ( .A1(KEYINPUT8), .A2(n1422), .A3(n1304), .ZN(n1421) );
INV_X1 U1090 ( .A(n1375), .ZN(n1304) );
NAND2_X1 U1091 ( .A1(KEYINPUT45), .A2(n1423), .ZN(n1422) );
NAND3_X1 U1092 ( .A1(n1424), .A2(n1425), .A3(n1375), .ZN(n1420) );
INV_X1 U1093 ( .A(KEYINPUT8), .ZN(n1425) );
NAND2_X1 U1094 ( .A1(n1426), .A2(n1423), .ZN(n1424) );
NAND2_X1 U1095 ( .A1(n1318), .A2(n1427), .ZN(n1423) );
INV_X1 U1096 ( .A(G125), .ZN(n1318) );
NAND2_X1 U1097 ( .A1(G125), .A2(n1428), .ZN(n1419) );
NAND2_X1 U1098 ( .A1(n1429), .A2(n1427), .ZN(n1428) );
INV_X1 U1099 ( .A(KEYINPUT2), .ZN(n1427) );
XNOR2_X1 U1100 ( .A(n1426), .B(n1375), .ZN(n1429) );
XNOR2_X1 U1101 ( .A(n1403), .B(n1407), .ZN(n1375) );
XOR2_X1 U1102 ( .A(G143), .B(G146), .Z(n1407) );
XNOR2_X1 U1103 ( .A(G128), .B(KEYINPUT37), .ZN(n1403) );
INV_X1 U1104 ( .A(KEYINPUT45), .ZN(n1426) );
XOR2_X1 U1105 ( .A(n1430), .B(n1431), .Z(n1299) );
XNOR2_X1 U1106 ( .A(n1202), .B(n1198), .ZN(n1431) );
XNOR2_X1 U1107 ( .A(n1432), .B(n1433), .ZN(n1198) );
XNOR2_X1 U1108 ( .A(KEYINPUT48), .B(n1243), .ZN(n1433) );
INV_X1 U1109 ( .A(G101), .ZN(n1243) );
XNOR2_X1 U1110 ( .A(n1370), .B(n1434), .ZN(n1432) );
NOR2_X1 U1111 ( .A1(n1435), .A2(KEYINPUT13), .ZN(n1434) );
INV_X1 U1112 ( .A(n1402), .ZN(n1435) );
NAND2_X1 U1113 ( .A1(n1436), .A2(n1401), .ZN(n1402) );
NAND2_X1 U1114 ( .A1(n1437), .A2(G107), .ZN(n1401) );
XNOR2_X1 U1115 ( .A(KEYINPUT52), .B(G104), .ZN(n1437) );
NAND2_X1 U1116 ( .A1(n1438), .A2(n1439), .ZN(n1436) );
INV_X1 U1117 ( .A(G107), .ZN(n1439) );
XOR2_X1 U1118 ( .A(KEYINPUT52), .B(G104), .Z(n1438) );
XNOR2_X1 U1119 ( .A(n1440), .B(n1345), .ZN(n1370) );
XNOR2_X1 U1120 ( .A(G119), .B(KEYINPUT11), .ZN(n1345) );
OR2_X1 U1121 ( .A1(KEYINPUT49), .A2(n1255), .ZN(n1202) );
INV_X1 U1122 ( .A(G110), .ZN(n1255) );
NOR2_X1 U1123 ( .A1(n1309), .A2(n1308), .ZN(n1150) );
INV_X1 U1124 ( .A(n1328), .ZN(n1308) );
XOR2_X1 U1125 ( .A(n1441), .B(n1442), .Z(n1328) );
INV_X1 U1126 ( .A(n1175), .ZN(n1442) );
NOR2_X1 U1127 ( .A1(n1221), .A2(G902), .ZN(n1175) );
INV_X1 U1128 ( .A(n1218), .ZN(n1221) );
XNOR2_X1 U1129 ( .A(n1443), .B(n1444), .ZN(n1218) );
XOR2_X1 U1130 ( .A(n1445), .B(n1446), .Z(n1444) );
XNOR2_X1 U1131 ( .A(n1344), .B(G107), .ZN(n1446) );
INV_X1 U1132 ( .A(G128), .ZN(n1344) );
XNOR2_X1 U1133 ( .A(n1409), .B(G134), .ZN(n1445) );
XNOR2_X1 U1134 ( .A(n1447), .B(n1448), .ZN(n1443) );
INV_X1 U1135 ( .A(n1440), .ZN(n1448) );
XOR2_X1 U1136 ( .A(G116), .B(KEYINPUT51), .Z(n1440) );
XOR2_X1 U1137 ( .A(n1449), .B(n1450), .Z(n1447) );
NOR3_X1 U1138 ( .A1(n1166), .A2(G953), .A3(n1164), .ZN(n1450) );
INV_X1 U1139 ( .A(G217), .ZN(n1164) );
INV_X1 U1140 ( .A(G234), .ZN(n1166) );
NAND2_X1 U1141 ( .A1(KEYINPUT15), .A2(n1203), .ZN(n1449) );
NAND2_X1 U1142 ( .A1(KEYINPUT28), .A2(n1219), .ZN(n1441) );
INV_X1 U1143 ( .A(G478), .ZN(n1219) );
XNOR2_X1 U1144 ( .A(n1172), .B(n1171), .ZN(n1309) );
INV_X1 U1145 ( .A(G475), .ZN(n1171) );
NOR2_X1 U1146 ( .A1(n1228), .A2(G902), .ZN(n1172) );
INV_X1 U1147 ( .A(n1226), .ZN(n1228) );
XNOR2_X1 U1148 ( .A(n1451), .B(n1452), .ZN(n1226) );
XOR2_X1 U1149 ( .A(n1453), .B(n1454), .Z(n1452) );
XNOR2_X1 U1150 ( .A(n1409), .B(n1455), .ZN(n1454) );
NOR2_X1 U1151 ( .A1(KEYINPUT18), .A2(n1456), .ZN(n1455) );
XOR2_X1 U1152 ( .A(G104), .B(n1430), .Z(n1456) );
XOR2_X1 U1153 ( .A(G113), .B(n1203), .Z(n1430) );
XOR2_X1 U1154 ( .A(G122), .B(KEYINPUT29), .Z(n1203) );
INV_X1 U1155 ( .A(G143), .ZN(n1409) );
NOR3_X1 U1156 ( .A1(n1411), .A2(G953), .A3(G237), .ZN(n1453) );
INV_X1 U1157 ( .A(G214), .ZN(n1411) );
XOR2_X1 U1158 ( .A(n1457), .B(n1185), .Z(n1451) );
XOR2_X1 U1159 ( .A(G140), .B(G125), .Z(n1185) );
XOR2_X1 U1160 ( .A(n1458), .B(n1394), .Z(n1457) );
XOR2_X1 U1161 ( .A(G131), .B(KEYINPUT30), .Z(n1394) );
NAND2_X1 U1162 ( .A1(KEYINPUT33), .A2(n1459), .ZN(n1458) );
INV_X1 U1163 ( .A(G146), .ZN(n1459) );
endmodule


