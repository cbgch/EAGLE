//Key = 0010000101010011110100011001000101111111011110100010101001101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
n1426;

XOR2_X1 U771 ( .A(n1086), .B(n1087), .Z(G9) );
NAND2_X1 U772 ( .A1(KEYINPUT44), .A2(n1088), .ZN(n1087) );
NOR2_X1 U773 ( .A1(n1089), .A2(n1090), .ZN(G75) );
NOR4_X1 U774 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
NOR3_X1 U775 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
NOR2_X1 U776 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NOR2_X1 U777 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U778 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U779 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U780 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U781 ( .A1(n1108), .A2(n1109), .ZN(n1102) );
NOR2_X1 U782 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR2_X1 U783 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NOR3_X1 U784 ( .A1(n1105), .A2(n1114), .A3(n1109), .ZN(n1098) );
NOR2_X1 U785 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR3_X1 U786 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1092) );
XOR2_X1 U787 ( .A(KEYINPUT21), .B(n1120), .Z(n1117) );
NAND3_X1 U788 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1091) );
NAND2_X1 U789 ( .A1(n1124), .A2(n1125), .ZN(n1122) );
XNOR2_X1 U790 ( .A(KEYINPUT28), .B(n1118), .ZN(n1124) );
OR4_X1 U791 ( .A1(n1095), .A2(n1101), .A3(n1105), .A4(n1109), .ZN(n1118) );
INV_X1 U792 ( .A(n1126), .ZN(n1105) );
NOR3_X1 U793 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1089) );
AND4_X1 U794 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1093) );
NOR4_X1 U795 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1130) );
NOR2_X1 U796 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NOR2_X1 U797 ( .A1(G469), .A2(n1137), .ZN(n1133) );
NOR2_X1 U798 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
AND2_X1 U799 ( .A1(n1136), .A2(KEYINPUT62), .ZN(n1139) );
NAND2_X1 U800 ( .A1(KEYINPUT50), .A2(n1140), .ZN(n1136) );
NOR2_X1 U801 ( .A1(KEYINPUT62), .A2(n1141), .ZN(n1138) );
INV_X1 U802 ( .A(n1140), .ZN(n1141) );
XOR2_X1 U803 ( .A(n1142), .B(n1143), .Z(n1132) );
NAND3_X1 U804 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1131) );
XOR2_X1 U805 ( .A(n1147), .B(KEYINPUT5), .Z(n1146) );
XOR2_X1 U806 ( .A(n1148), .B(n1149), .Z(n1144) );
XOR2_X1 U807 ( .A(KEYINPUT8), .B(G472), .Z(n1149) );
NOR3_X1 U808 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1129) );
INV_X1 U809 ( .A(n1119), .ZN(n1151) );
NAND2_X1 U810 ( .A1(G478), .A2(n1153), .ZN(n1127) );
NAND2_X1 U811 ( .A1(n1154), .A2(n1155), .ZN(G72) );
NAND2_X1 U812 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U813 ( .A1(G953), .A2(n1158), .ZN(n1157) );
NAND2_X1 U814 ( .A1(G900), .A2(G227), .ZN(n1158) );
INV_X1 U815 ( .A(n1159), .ZN(n1156) );
NAND2_X1 U816 ( .A1(n1159), .A2(n1160), .ZN(n1154) );
NAND2_X1 U817 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U818 ( .A1(G953), .A2(n1163), .ZN(n1162) );
INV_X1 U819 ( .A(n1164), .ZN(n1161) );
XOR2_X1 U820 ( .A(n1165), .B(n1166), .Z(n1159) );
NOR4_X1 U821 ( .A1(KEYINPUT10), .A2(n1164), .A3(n1167), .A4(n1168), .ZN(n1166) );
XOR2_X1 U822 ( .A(n1169), .B(KEYINPUT11), .Z(n1168) );
NAND2_X1 U823 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
NOR2_X1 U824 ( .A1(n1170), .A2(n1171), .ZN(n1167) );
XOR2_X1 U825 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U826 ( .A(n1174), .B(G134), .Z(n1172) );
XNOR2_X1 U827 ( .A(G125), .B(n1175), .ZN(n1170) );
XOR2_X1 U828 ( .A(KEYINPUT31), .B(G140), .Z(n1175) );
NAND2_X1 U829 ( .A1(n1176), .A2(n1177), .ZN(n1165) );
XOR2_X1 U830 ( .A(n1178), .B(KEYINPUT55), .Z(n1176) );
XOR2_X1 U831 ( .A(n1179), .B(n1180), .Z(G69) );
NOR2_X1 U832 ( .A1(n1181), .A2(n1121), .ZN(n1180) );
AND2_X1 U833 ( .A1(n1182), .A2(n1178), .ZN(n1121) );
AND3_X1 U834 ( .A1(G898), .A2(G953), .A3(G224), .ZN(n1181) );
NAND2_X1 U835 ( .A1(KEYINPUT17), .A2(n1183), .ZN(n1179) );
NAND2_X1 U836 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
INV_X1 U837 ( .A(n1186), .ZN(n1185) );
XOR2_X1 U838 ( .A(n1187), .B(n1188), .Z(n1184) );
NAND3_X1 U839 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1187) );
NAND2_X1 U840 ( .A1(n1192), .A2(n1193), .ZN(n1190) );
INV_X1 U841 ( .A(KEYINPUT57), .ZN(n1193) );
NAND2_X1 U842 ( .A1(n1194), .A2(KEYINPUT57), .ZN(n1189) );
NOR2_X1 U843 ( .A1(n1195), .A2(n1196), .ZN(G66) );
NOR2_X1 U844 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XOR2_X1 U845 ( .A(n1199), .B(KEYINPUT52), .Z(n1198) );
NAND2_X1 U846 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
OR2_X1 U847 ( .A1(n1128), .A2(n1202), .ZN(n1201) );
NOR4_X1 U848 ( .A1(n1200), .A2(n1203), .A3(n1204), .A4(n1202), .ZN(n1197) );
XNOR2_X1 U849 ( .A(n1205), .B(KEYINPUT26), .ZN(n1202) );
NOR2_X1 U850 ( .A1(n1195), .A2(n1206), .ZN(G63) );
XOR2_X1 U851 ( .A(n1207), .B(n1208), .Z(n1206) );
AND2_X1 U852 ( .A1(G478), .A2(n1209), .ZN(n1208) );
NOR2_X1 U853 ( .A1(n1195), .A2(n1210), .ZN(G60) );
XOR2_X1 U854 ( .A(n1211), .B(n1212), .Z(n1210) );
AND2_X1 U855 ( .A1(G475), .A2(n1209), .ZN(n1212) );
XNOR2_X1 U856 ( .A(G104), .B(n1213), .ZN(G6) );
NAND2_X1 U857 ( .A1(KEYINPUT36), .A2(n1214), .ZN(n1213) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1215), .ZN(G57) );
XOR2_X1 U859 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U860 ( .A(n1218), .B(n1219), .Z(n1217) );
AND2_X1 U861 ( .A1(G472), .A2(n1209), .ZN(n1219) );
NOR2_X1 U862 ( .A1(KEYINPUT20), .A2(n1220), .ZN(n1218) );
NOR2_X1 U863 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND3_X1 U864 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1216) );
NAND2_X1 U865 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
INV_X1 U866 ( .A(KEYINPUT60), .ZN(n1227) );
NAND3_X1 U867 ( .A1(KEYINPUT60), .A2(n1228), .A3(n1229), .ZN(n1224) );
OR2_X1 U868 ( .A1(n1229), .A2(n1228), .ZN(n1223) );
NOR2_X1 U869 ( .A1(n1230), .A2(n1226), .ZN(n1228) );
XNOR2_X1 U870 ( .A(n1231), .B(n1232), .ZN(n1226) );
NAND2_X1 U871 ( .A1(KEYINPUT61), .A2(n1233), .ZN(n1231) );
INV_X1 U872 ( .A(KEYINPUT27), .ZN(n1230) );
NOR2_X1 U873 ( .A1(n1195), .A2(n1234), .ZN(G54) );
XOR2_X1 U874 ( .A(n1235), .B(n1236), .Z(n1234) );
XOR2_X1 U875 ( .A(n1237), .B(n1238), .Z(n1235) );
NOR2_X1 U876 ( .A1(n1135), .A2(n1239), .ZN(n1238) );
INV_X1 U877 ( .A(G469), .ZN(n1135) );
NAND2_X1 U878 ( .A1(KEYINPUT2), .A2(n1240), .ZN(n1237) );
NOR2_X1 U879 ( .A1(n1195), .A2(n1241), .ZN(G51) );
NOR2_X1 U880 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U881 ( .A(KEYINPUT13), .B(n1244), .Z(n1243) );
NOR2_X1 U882 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
AND2_X1 U883 ( .A1(n1246), .A2(n1245), .ZN(n1242) );
XNOR2_X1 U884 ( .A(n1247), .B(n1248), .ZN(n1245) );
NOR2_X1 U885 ( .A1(KEYINPUT4), .A2(n1249), .ZN(n1248) );
NAND2_X1 U886 ( .A1(n1209), .A2(n1250), .ZN(n1246) );
INV_X1 U887 ( .A(n1239), .ZN(n1209) );
NAND2_X1 U888 ( .A1(G902), .A2(n1205), .ZN(n1239) );
NAND2_X1 U889 ( .A1(n1123), .A2(n1182), .ZN(n1205) );
AND4_X1 U890 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1182) );
NOR4_X1 U891 ( .A1(n1255), .A2(n1088), .A3(n1214), .A4(n1256), .ZN(n1254) );
INV_X1 U892 ( .A(n1257), .ZN(n1256) );
AND3_X1 U893 ( .A1(n1258), .A2(n1259), .A3(n1116), .ZN(n1214) );
AND3_X1 U894 ( .A1(n1258), .A2(n1259), .A3(n1115), .ZN(n1088) );
NOR2_X1 U895 ( .A1(n1260), .A2(n1261), .ZN(n1253) );
NOR2_X1 U896 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XOR2_X1 U897 ( .A(n1264), .B(KEYINPUT25), .Z(n1263) );
NOR3_X1 U898 ( .A1(n1101), .A2(n1265), .A3(n1266), .ZN(n1260) );
INV_X1 U899 ( .A(n1177), .ZN(n1123) );
NAND4_X1 U900 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1177) );
AND4_X1 U901 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1270) );
OR2_X1 U902 ( .A1(KEYINPUT29), .A2(n1275), .ZN(n1274) );
AND2_X1 U903 ( .A1(n1276), .A2(n1277), .ZN(n1269) );
NAND2_X1 U904 ( .A1(n1116), .A2(n1278), .ZN(n1267) );
NAND2_X1 U905 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND4_X1 U906 ( .A1(KEYINPUT29), .A2(n1281), .A3(n1282), .A4(n1111), .ZN(n1280) );
NAND2_X1 U907 ( .A1(n1283), .A2(n1284), .ZN(n1279) );
NOR2_X1 U908 ( .A1(n1178), .A2(G952), .ZN(n1195) );
XOR2_X1 U909 ( .A(n1275), .B(n1285), .Z(G48) );
NAND2_X1 U910 ( .A1(KEYINPUT46), .A2(G146), .ZN(n1285) );
NAND2_X1 U911 ( .A1(n1286), .A2(n1282), .ZN(n1275) );
XOR2_X1 U912 ( .A(n1287), .B(n1273), .Z(G45) );
NAND4_X1 U913 ( .A1(n1283), .A2(n1125), .A3(n1288), .A4(n1289), .ZN(n1273) );
NAND2_X1 U914 ( .A1(n1290), .A2(n1291), .ZN(G42) );
NAND2_X1 U915 ( .A1(G140), .A2(n1272), .ZN(n1291) );
XOR2_X1 U916 ( .A(KEYINPUT23), .B(n1292), .Z(n1290) );
NOR2_X1 U917 ( .A1(G140), .A2(n1272), .ZN(n1292) );
NAND3_X1 U918 ( .A1(n1284), .A2(n1106), .A3(n1286), .ZN(n1272) );
AND3_X1 U919 ( .A1(n1111), .A2(n1293), .A3(n1116), .ZN(n1286) );
NAND2_X1 U920 ( .A1(n1294), .A2(n1295), .ZN(G39) );
NAND2_X1 U921 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U922 ( .A(KEYINPUT63), .B(n1298), .Z(n1294) );
NOR2_X1 U923 ( .A1(n1296), .A2(n1297), .ZN(n1298) );
INV_X1 U924 ( .A(G137), .ZN(n1297) );
INV_X1 U925 ( .A(n1268), .ZN(n1296) );
NAND4_X1 U926 ( .A1(n1284), .A2(n1111), .A3(n1299), .A4(n1300), .ZN(n1268) );
NOR3_X1 U927 ( .A1(n1301), .A2(n1281), .A3(n1302), .ZN(n1300) );
XOR2_X1 U928 ( .A(n1303), .B(n1271), .Z(G36) );
NAND3_X1 U929 ( .A1(n1284), .A2(n1115), .A3(n1283), .ZN(n1271) );
INV_X1 U930 ( .A(n1097), .ZN(n1284) );
XNOR2_X1 U931 ( .A(G131), .B(n1304), .ZN(G33) );
NAND3_X1 U932 ( .A1(n1283), .A2(n1116), .A3(n1305), .ZN(n1304) );
XOR2_X1 U933 ( .A(n1097), .B(KEYINPUT38), .Z(n1305) );
NAND2_X1 U934 ( .A1(n1306), .A2(n1119), .ZN(n1097) );
AND3_X1 U935 ( .A1(n1111), .A2(n1293), .A3(n1107), .ZN(n1283) );
XOR2_X1 U936 ( .A(n1307), .B(KEYINPUT53), .Z(n1111) );
XOR2_X1 U937 ( .A(n1277), .B(n1308), .Z(G30) );
XOR2_X1 U938 ( .A(n1309), .B(KEYINPUT12), .Z(n1308) );
NAND4_X1 U939 ( .A1(n1282), .A2(n1115), .A3(n1307), .A4(n1293), .ZN(n1277) );
XOR2_X1 U940 ( .A(n1255), .B(n1310), .Z(G3) );
NOR2_X1 U941 ( .A1(KEYINPUT59), .A2(n1311), .ZN(n1310) );
AND3_X1 U942 ( .A1(n1299), .A2(n1259), .A3(n1107), .ZN(n1255) );
INV_X1 U943 ( .A(n1265), .ZN(n1259) );
NAND3_X1 U944 ( .A1(n1307), .A2(n1312), .A3(n1313), .ZN(n1265) );
XNOR2_X1 U945 ( .A(G125), .B(n1276), .ZN(G27) );
NAND4_X1 U946 ( .A1(n1126), .A2(n1106), .A3(n1314), .A4(n1116), .ZN(n1276) );
NOR2_X1 U947 ( .A1(n1281), .A2(n1262), .ZN(n1314) );
INV_X1 U948 ( .A(n1293), .ZN(n1281) );
NAND2_X1 U949 ( .A1(n1095), .A2(n1315), .ZN(n1293) );
NAND3_X1 U950 ( .A1(G902), .A2(n1316), .A3(n1164), .ZN(n1315) );
NOR2_X1 U951 ( .A1(n1178), .A2(G900), .ZN(n1164) );
INV_X1 U952 ( .A(n1266), .ZN(n1106) );
XOR2_X1 U953 ( .A(G122), .B(n1317), .Z(G24) );
NOR2_X1 U954 ( .A1(n1262), .A2(n1264), .ZN(n1317) );
NAND4_X1 U955 ( .A1(n1318), .A2(n1258), .A3(n1288), .A4(n1289), .ZN(n1264) );
INV_X1 U956 ( .A(n1109), .ZN(n1258) );
NAND2_X1 U957 ( .A1(n1302), .A2(n1301), .ZN(n1109) );
XOR2_X1 U958 ( .A(n1319), .B(n1251), .Z(G21) );
NAND3_X1 U959 ( .A1(n1299), .A2(n1282), .A3(n1318), .ZN(n1251) );
NOR3_X1 U960 ( .A1(n1301), .A2(n1302), .A3(n1262), .ZN(n1282) );
INV_X1 U961 ( .A(n1320), .ZN(n1301) );
INV_X1 U962 ( .A(n1101), .ZN(n1299) );
XNOR2_X1 U963 ( .A(G116), .B(n1252), .ZN(G18) );
NAND4_X1 U964 ( .A1(n1318), .A2(n1107), .A3(n1115), .A4(n1125), .ZN(n1252) );
INV_X1 U965 ( .A(n1262), .ZN(n1125) );
XOR2_X1 U966 ( .A(n1321), .B(KEYINPUT3), .Z(n1262) );
NOR2_X1 U967 ( .A1(n1288), .A2(n1322), .ZN(n1115) );
INV_X1 U968 ( .A(n1145), .ZN(n1288) );
XOR2_X1 U969 ( .A(n1323), .B(n1257), .Z(G15) );
NAND4_X1 U970 ( .A1(n1318), .A2(n1107), .A3(n1116), .A4(n1313), .ZN(n1257) );
INV_X1 U971 ( .A(n1321), .ZN(n1313) );
NOR2_X1 U972 ( .A1(n1289), .A2(n1145), .ZN(n1116) );
INV_X1 U973 ( .A(n1322), .ZN(n1289) );
NOR2_X1 U974 ( .A1(n1320), .A2(n1302), .ZN(n1107) );
AND2_X1 U975 ( .A1(n1126), .A2(n1312), .ZN(n1318) );
NOR2_X1 U976 ( .A1(n1112), .A2(n1150), .ZN(n1126) );
INV_X1 U977 ( .A(n1113), .ZN(n1150) );
XOR2_X1 U978 ( .A(G110), .B(n1324), .Z(G12) );
NOR4_X1 U979 ( .A1(n1321), .A2(n1325), .A3(n1266), .A4(n1101), .ZN(n1324) );
NAND2_X1 U980 ( .A1(n1322), .A2(n1145), .ZN(n1101) );
XNOR2_X1 U981 ( .A(G475), .B(n1326), .ZN(n1145) );
NOR2_X1 U982 ( .A1(G902), .A2(n1211), .ZN(n1326) );
NAND2_X1 U983 ( .A1(n1327), .A2(n1328), .ZN(n1211) );
NAND2_X1 U984 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
NAND2_X1 U985 ( .A1(KEYINPUT35), .A2(n1331), .ZN(n1330) );
OR2_X1 U986 ( .A1(n1332), .A2(KEYINPUT47), .ZN(n1331) );
INV_X1 U987 ( .A(n1333), .ZN(n1329) );
NAND2_X1 U988 ( .A1(n1332), .A2(n1334), .ZN(n1327) );
NAND2_X1 U989 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND2_X1 U990 ( .A1(n1333), .A2(KEYINPUT35), .ZN(n1336) );
XNOR2_X1 U991 ( .A(G104), .B(n1337), .ZN(n1333) );
XOR2_X1 U992 ( .A(G122), .B(G113), .Z(n1337) );
INV_X1 U993 ( .A(KEYINPUT47), .ZN(n1335) );
XNOR2_X1 U994 ( .A(n1338), .B(n1339), .ZN(n1332) );
XOR2_X1 U995 ( .A(n1340), .B(n1341), .Z(n1339) );
NAND2_X1 U996 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
OR2_X1 U997 ( .A1(n1344), .A2(G125), .ZN(n1343) );
XOR2_X1 U998 ( .A(n1345), .B(KEYINPUT48), .Z(n1342) );
NAND2_X1 U999 ( .A1(G125), .A2(n1344), .ZN(n1345) );
XNOR2_X1 U1000 ( .A(G131), .B(n1346), .ZN(n1338) );
AND3_X1 U1001 ( .A1(G214), .A2(n1178), .A3(n1347), .ZN(n1346) );
NOR2_X1 U1002 ( .A1(n1348), .A2(n1152), .ZN(n1322) );
NOR3_X1 U1003 ( .A1(G478), .A2(G902), .A3(n1207), .ZN(n1152) );
AND2_X1 U1004 ( .A1(n1349), .A2(n1153), .ZN(n1348) );
NAND2_X1 U1005 ( .A1(n1350), .A2(n1204), .ZN(n1153) );
INV_X1 U1006 ( .A(n1207), .ZN(n1350) );
XOR2_X1 U1007 ( .A(n1351), .B(n1352), .Z(n1207) );
NOR2_X1 U1008 ( .A1(KEYINPUT22), .A2(n1353), .ZN(n1352) );
XOR2_X1 U1009 ( .A(n1354), .B(n1355), .Z(n1353) );
XOR2_X1 U1010 ( .A(G128), .B(n1356), .Z(n1355) );
XOR2_X1 U1011 ( .A(G143), .B(G134), .Z(n1356) );
XOR2_X1 U1012 ( .A(n1086), .B(n1357), .Z(n1354) );
XOR2_X1 U1013 ( .A(G122), .B(G116), .Z(n1357) );
NAND3_X1 U1014 ( .A1(G234), .A2(G217), .A3(n1358), .ZN(n1351) );
XOR2_X1 U1015 ( .A(n1178), .B(KEYINPUT51), .Z(n1358) );
XOR2_X1 U1016 ( .A(KEYINPUT30), .B(G478), .Z(n1349) );
NAND2_X1 U1017 ( .A1(n1302), .A2(n1320), .ZN(n1266) );
NAND2_X1 U1018 ( .A1(n1359), .A2(n1360), .ZN(n1320) );
NAND2_X1 U1019 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
INV_X1 U1020 ( .A(KEYINPUT32), .ZN(n1362) );
NAND2_X1 U1021 ( .A1(n1128), .A2(n1147), .ZN(n1361) );
NAND2_X1 U1022 ( .A1(n1363), .A2(n1203), .ZN(n1147) );
OR2_X1 U1023 ( .A1(n1203), .A2(n1363), .ZN(n1128) );
NAND2_X1 U1024 ( .A1(KEYINPUT32), .A2(n1364), .ZN(n1359) );
XOR2_X1 U1025 ( .A(n1363), .B(n1203), .Z(n1364) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1365), .ZN(n1203) );
AND2_X1 U1027 ( .A1(n1200), .A2(n1204), .ZN(n1363) );
XOR2_X1 U1028 ( .A(n1366), .B(n1367), .Z(n1200) );
XOR2_X1 U1029 ( .A(n1368), .B(n1369), .Z(n1367) );
XOR2_X1 U1030 ( .A(G140), .B(G137), .Z(n1369) );
XOR2_X1 U1031 ( .A(KEYINPUT19), .B(G146), .Z(n1368) );
XOR2_X1 U1032 ( .A(n1370), .B(n1371), .Z(n1366) );
XOR2_X1 U1033 ( .A(n1372), .B(n1373), .Z(n1371) );
NAND3_X1 U1034 ( .A1(G234), .A2(n1178), .A3(G221), .ZN(n1373) );
NAND2_X1 U1035 ( .A1(n1374), .A2(n1375), .ZN(n1372) );
NAND2_X1 U1036 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
XOR2_X1 U1037 ( .A(KEYINPUT54), .B(n1378), .Z(n1374) );
NOR2_X1 U1038 ( .A1(n1376), .A2(n1377), .ZN(n1378) );
XOR2_X1 U1039 ( .A(G128), .B(G119), .Z(n1377) );
NAND2_X1 U1040 ( .A1(KEYINPUT15), .A2(G125), .ZN(n1370) );
XOR2_X1 U1041 ( .A(n1379), .B(G472), .Z(n1302) );
NAND2_X1 U1042 ( .A1(KEYINPUT7), .A2(n1380), .ZN(n1379) );
XNOR2_X1 U1043 ( .A(KEYINPUT1), .B(n1148), .ZN(n1380) );
NAND2_X1 U1044 ( .A1(n1381), .A2(n1204), .ZN(n1148) );
XOR2_X1 U1045 ( .A(n1382), .B(n1383), .Z(n1381) );
XOR2_X1 U1046 ( .A(n1233), .B(n1229), .Z(n1383) );
XOR2_X1 U1047 ( .A(n1384), .B(n1385), .Z(n1229) );
XOR2_X1 U1048 ( .A(KEYINPUT24), .B(G113), .Z(n1385) );
NAND3_X1 U1049 ( .A1(n1386), .A2(n1387), .A3(n1388), .ZN(n1384) );
NAND2_X1 U1050 ( .A1(KEYINPUT0), .A2(G116), .ZN(n1388) );
NAND3_X1 U1051 ( .A1(n1389), .A2(n1390), .A3(n1319), .ZN(n1387) );
INV_X1 U1052 ( .A(KEYINPUT0), .ZN(n1390) );
OR2_X1 U1053 ( .A1(n1319), .A2(n1389), .ZN(n1386) );
NOR2_X1 U1054 ( .A1(n1391), .A2(G116), .ZN(n1389) );
INV_X1 U1055 ( .A(KEYINPUT33), .ZN(n1391) );
INV_X1 U1056 ( .A(G119), .ZN(n1319) );
XOR2_X1 U1057 ( .A(n1232), .B(n1392), .Z(n1382) );
XOR2_X1 U1058 ( .A(KEYINPUT6), .B(n1393), .Z(n1392) );
NOR2_X1 U1059 ( .A1(n1221), .A2(n1394), .ZN(n1393) );
XOR2_X1 U1060 ( .A(KEYINPUT56), .B(n1222), .Z(n1394) );
NOR2_X1 U1061 ( .A1(n1311), .A2(n1395), .ZN(n1222) );
AND2_X1 U1062 ( .A1(n1311), .A2(n1395), .ZN(n1221) );
NAND3_X1 U1063 ( .A1(n1347), .A2(n1178), .A3(n1396), .ZN(n1395) );
XOR2_X1 U1064 ( .A(KEYINPUT40), .B(G210), .Z(n1396) );
NAND2_X1 U1065 ( .A1(n1397), .A2(n1312), .ZN(n1325) );
NAND2_X1 U1066 ( .A1(n1095), .A2(n1398), .ZN(n1312) );
NAND3_X1 U1067 ( .A1(n1186), .A2(n1316), .A3(G902), .ZN(n1398) );
NOR2_X1 U1068 ( .A1(n1178), .A2(G898), .ZN(n1186) );
NAND3_X1 U1069 ( .A1(n1316), .A2(n1178), .A3(G952), .ZN(n1095) );
NAND2_X1 U1070 ( .A1(G237), .A2(G234), .ZN(n1316) );
XOR2_X1 U1071 ( .A(KEYINPUT45), .B(n1307), .Z(n1397) );
AND2_X1 U1072 ( .A1(n1112), .A2(n1113), .ZN(n1307) );
NAND2_X1 U1073 ( .A1(G221), .A2(n1365), .ZN(n1113) );
NAND2_X1 U1074 ( .A1(G234), .A2(n1204), .ZN(n1365) );
XNOR2_X1 U1075 ( .A(n1140), .B(G469), .ZN(n1112) );
NAND2_X1 U1076 ( .A1(n1399), .A2(n1204), .ZN(n1140) );
XOR2_X1 U1077 ( .A(n1236), .B(n1240), .Z(n1399) );
XOR2_X1 U1078 ( .A(n1344), .B(n1376), .Z(n1240) );
INV_X1 U1079 ( .A(G140), .ZN(n1344) );
XNOR2_X1 U1080 ( .A(n1400), .B(n1401), .ZN(n1236) );
XOR2_X1 U1081 ( .A(n1402), .B(n1403), .Z(n1401) );
XOR2_X1 U1082 ( .A(G104), .B(G101), .Z(n1403) );
XOR2_X1 U1083 ( .A(KEYINPUT49), .B(G107), .Z(n1402) );
XOR2_X1 U1084 ( .A(n1404), .B(n1232), .Z(n1400) );
XNOR2_X1 U1085 ( .A(n1405), .B(n1173), .ZN(n1232) );
XOR2_X1 U1086 ( .A(G131), .B(G137), .Z(n1173) );
NAND2_X1 U1087 ( .A1(KEYINPUT14), .A2(n1303), .ZN(n1405) );
INV_X1 U1088 ( .A(G134), .ZN(n1303) );
XOR2_X1 U1089 ( .A(n1174), .B(n1406), .Z(n1404) );
NOR2_X1 U1090 ( .A1(G953), .A2(n1163), .ZN(n1406) );
INV_X1 U1091 ( .A(G227), .ZN(n1163) );
NAND2_X1 U1092 ( .A1(n1407), .A2(n1408), .ZN(n1174) );
NAND2_X1 U1093 ( .A1(n1341), .A2(n1309), .ZN(n1408) );
XOR2_X1 U1094 ( .A(KEYINPUT41), .B(n1409), .Z(n1407) );
NOR2_X1 U1095 ( .A1(n1341), .A2(n1309), .ZN(n1409) );
INV_X1 U1096 ( .A(G128), .ZN(n1309) );
XOR2_X1 U1097 ( .A(n1287), .B(G146), .Z(n1341) );
INV_X1 U1098 ( .A(G143), .ZN(n1287) );
NAND2_X1 U1099 ( .A1(n1120), .A2(n1119), .ZN(n1321) );
NAND2_X1 U1100 ( .A1(G214), .A2(n1410), .ZN(n1119) );
INV_X1 U1101 ( .A(n1306), .ZN(n1120) );
XOR2_X1 U1102 ( .A(n1411), .B(n1250), .Z(n1306) );
INV_X1 U1103 ( .A(n1143), .ZN(n1250) );
NAND2_X1 U1104 ( .A1(G210), .A2(n1410), .ZN(n1143) );
NAND2_X1 U1105 ( .A1(n1204), .A2(n1347), .ZN(n1410) );
INV_X1 U1106 ( .A(G237), .ZN(n1347) );
NAND2_X1 U1107 ( .A1(n1412), .A2(KEYINPUT39), .ZN(n1411) );
XOR2_X1 U1108 ( .A(n1142), .B(KEYINPUT43), .Z(n1412) );
NAND2_X1 U1109 ( .A1(n1413), .A2(n1204), .ZN(n1142) );
INV_X1 U1110 ( .A(G902), .ZN(n1204) );
XNOR2_X1 U1111 ( .A(n1249), .B(n1414), .ZN(n1413) );
XOR2_X1 U1112 ( .A(n1247), .B(KEYINPUT9), .Z(n1414) );
XOR2_X1 U1113 ( .A(n1188), .B(n1415), .Z(n1247) );
XOR2_X1 U1114 ( .A(n1416), .B(n1417), .Z(n1415) );
AND2_X1 U1115 ( .A1(n1178), .A2(G224), .ZN(n1417) );
INV_X1 U1116 ( .A(G953), .ZN(n1178) );
NOR3_X1 U1117 ( .A1(n1194), .A2(KEYINPUT18), .A3(n1418), .ZN(n1416) );
INV_X1 U1118 ( .A(n1191), .ZN(n1418) );
NAND2_X1 U1119 ( .A1(n1419), .A2(n1192), .ZN(n1191) );
NOR2_X1 U1120 ( .A1(n1192), .A2(n1419), .ZN(n1194) );
XOR2_X1 U1121 ( .A(n1420), .B(n1421), .Z(n1419) );
XNOR2_X1 U1122 ( .A(G104), .B(n1422), .ZN(n1421) );
NAND2_X1 U1123 ( .A1(KEYINPUT58), .A2(n1086), .ZN(n1422) );
INV_X1 U1124 ( .A(G107), .ZN(n1086) );
NAND2_X1 U1125 ( .A1(KEYINPUT16), .A2(n1311), .ZN(n1420) );
INV_X1 U1126 ( .A(G101), .ZN(n1311) );
XNOR2_X1 U1127 ( .A(n1423), .B(n1424), .ZN(n1192) );
XOR2_X1 U1128 ( .A(KEYINPUT37), .B(G119), .Z(n1424) );
XOR2_X1 U1129 ( .A(n1323), .B(G116), .Z(n1423) );
INV_X1 U1130 ( .A(G113), .ZN(n1323) );
XOR2_X1 U1131 ( .A(G122), .B(n1376), .Z(n1188) );
XNOR2_X1 U1132 ( .A(G110), .B(KEYINPUT42), .ZN(n1376) );
XNOR2_X1 U1133 ( .A(n1233), .B(G125), .ZN(n1249) );
XOR2_X1 U1134 ( .A(n1425), .B(n1426), .Z(n1233) );
XOR2_X1 U1135 ( .A(G146), .B(G128), .Z(n1426) );
NAND2_X1 U1136 ( .A1(KEYINPUT34), .A2(G143), .ZN(n1425) );
endmodule


