//Key = 0000101000000010010111101110000000001101010111110111001101000101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328;

XNOR2_X1 U733 ( .A(G107), .B(n1006), .ZN(G9) );
NOR2_X1 U734 ( .A1(n1007), .A2(n1008), .ZN(G75) );
NOR4_X1 U735 ( .A1(n1009), .A2(n1010), .A3(G953), .A4(n1011), .ZN(n1008) );
NOR2_X1 U736 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NOR2_X1 U737 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR3_X1 U738 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
NOR3_X1 U739 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1017) );
AND3_X1 U740 ( .A1(n1022), .A2(n1023), .A3(KEYINPUT35), .ZN(n1021) );
NOR2_X1 U741 ( .A1(n1024), .A2(n1022), .ZN(n1020) );
NOR2_X1 U742 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NOR2_X1 U743 ( .A1(KEYINPUT35), .A2(n1027), .ZN(n1026) );
NOR3_X1 U744 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1025) );
NOR2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1019) );
NOR2_X1 U746 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR3_X1 U747 ( .A1(n1022), .A2(n1035), .A3(n1032), .ZN(n1014) );
NOR2_X1 U748 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NOR2_X1 U749 ( .A1(n1038), .A2(n1018), .ZN(n1037) );
NOR2_X1 U750 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR3_X1 U751 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1039) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1016), .ZN(n1036) );
NOR2_X1 U753 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
INV_X1 U755 ( .A(n1049), .ZN(n1012) );
NOR3_X1 U756 ( .A1(n1011), .A2(G953), .A3(G952), .ZN(n1007) );
AND4_X1 U757 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1011) );
NOR2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
XNOR2_X1 U759 ( .A(G472), .B(n1056), .ZN(n1055) );
NOR2_X1 U760 ( .A1(n1057), .A2(KEYINPUT10), .ZN(n1056) );
XOR2_X1 U761 ( .A(n1058), .B(n1059), .Z(n1054) );
NOR2_X1 U762 ( .A1(n1060), .A2(KEYINPUT0), .ZN(n1059) );
XOR2_X1 U763 ( .A(n1061), .B(n1062), .Z(G72) );
NOR2_X1 U764 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
XNOR2_X1 U765 ( .A(n1065), .B(n1066), .ZN(n1064) );
XOR2_X1 U766 ( .A(n1067), .B(n1068), .Z(n1066) );
NOR2_X1 U767 ( .A1(KEYINPUT2), .A2(n1069), .ZN(n1068) );
NAND2_X1 U768 ( .A1(n1070), .A2(n1071), .ZN(n1061) );
NAND2_X1 U769 ( .A1(KEYINPUT47), .A2(n1072), .ZN(n1071) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U771 ( .A1(G953), .A2(n1075), .ZN(n1074) );
INV_X1 U772 ( .A(n1063), .ZN(n1073) );
NAND2_X1 U773 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
NAND2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
XOR2_X1 U775 ( .A(KEYINPUT60), .B(n1080), .Z(n1079) );
XOR2_X1 U776 ( .A(n1081), .B(n1082), .Z(G69) );
NOR2_X1 U777 ( .A1(n1083), .A2(n1077), .ZN(n1082) );
NOR2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U779 ( .A1(n1086), .A2(n1087), .ZN(n1081) );
NAND2_X1 U780 ( .A1(n1088), .A2(n1077), .ZN(n1087) );
XOR2_X1 U781 ( .A(n1089), .B(n1090), .Z(n1088) );
OR3_X1 U782 ( .A1(n1085), .A2(n1090), .A3(n1077), .ZN(n1086) );
XNOR2_X1 U783 ( .A(n1091), .B(n1092), .ZN(n1090) );
XNOR2_X1 U784 ( .A(n1093), .B(n1094), .ZN(n1092) );
XOR2_X1 U785 ( .A(n1095), .B(KEYINPUT19), .Z(n1091) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XOR2_X1 U787 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U788 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NOR2_X1 U789 ( .A1(n1096), .A2(n1102), .ZN(G63) );
XOR2_X1 U790 ( .A(n1103), .B(n1104), .Z(n1102) );
AND2_X1 U791 ( .A1(G478), .A2(n1105), .ZN(n1103) );
NOR3_X1 U792 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(G60) );
NOR3_X1 U793 ( .A1(n1109), .A2(G953), .A3(G952), .ZN(n1108) );
AND2_X1 U794 ( .A1(n1109), .A2(n1096), .ZN(n1107) );
INV_X1 U795 ( .A(KEYINPUT48), .ZN(n1109) );
XNOR2_X1 U796 ( .A(n1110), .B(n1111), .ZN(n1106) );
AND2_X1 U797 ( .A1(G475), .A2(n1105), .ZN(n1111) );
XNOR2_X1 U798 ( .A(G104), .B(n1112), .ZN(G6) );
NOR2_X1 U799 ( .A1(n1096), .A2(n1113), .ZN(G57) );
XNOR2_X1 U800 ( .A(n1114), .B(n1115), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1116), .B(n1117), .Z(n1115) );
AND2_X1 U802 ( .A1(G472), .A2(n1105), .ZN(n1117) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
XOR2_X1 U804 ( .A(n1120), .B(KEYINPUT43), .Z(n1119) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U806 ( .A(n1123), .B(KEYINPUT32), .Z(n1121) );
NOR2_X1 U807 ( .A1(n1096), .A2(n1124), .ZN(G54) );
XOR2_X1 U808 ( .A(n1125), .B(n1126), .Z(n1124) );
XOR2_X1 U809 ( .A(n1127), .B(n1128), .Z(n1126) );
NOR2_X1 U810 ( .A1(KEYINPUT33), .A2(n1129), .ZN(n1127) );
XOR2_X1 U811 ( .A(n1130), .B(n1131), .Z(n1125) );
XOR2_X1 U812 ( .A(KEYINPUT46), .B(G110), .Z(n1131) );
NAND3_X1 U813 ( .A1(n1105), .A2(G469), .A3(KEYINPUT20), .ZN(n1130) );
INV_X1 U814 ( .A(n1101), .ZN(n1105) );
NOR2_X1 U815 ( .A1(n1096), .A2(n1132), .ZN(G51) );
XOR2_X1 U816 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U817 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U818 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR3_X1 U819 ( .A1(n1084), .A2(KEYINPUT56), .A3(G953), .ZN(n1137) );
NOR3_X1 U820 ( .A1(n1101), .A2(n1042), .A3(n1139), .ZN(n1135) );
NAND2_X1 U821 ( .A1(n1140), .A2(n1009), .ZN(n1101) );
NAND3_X1 U822 ( .A1(n1089), .A2(n1080), .A3(n1078), .ZN(n1009) );
AND3_X1 U823 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1078) );
NAND2_X1 U824 ( .A1(n1040), .A2(n1144), .ZN(n1143) );
NAND2_X1 U825 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U826 ( .A1(n1147), .A2(n1034), .ZN(n1146) );
XOR2_X1 U827 ( .A(n1148), .B(KEYINPUT13), .Z(n1145) );
AND3_X1 U828 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1080) );
NAND2_X1 U829 ( .A1(n1034), .A2(n1152), .ZN(n1151) );
NAND2_X1 U830 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND4_X1 U831 ( .A1(n1046), .A2(n1051), .A3(n1040), .A4(n1155), .ZN(n1154) );
NAND3_X1 U832 ( .A1(n1156), .A2(n1157), .A3(n1053), .ZN(n1153) );
OR2_X1 U833 ( .A1(n1158), .A2(KEYINPUT58), .ZN(n1157) );
NAND2_X1 U834 ( .A1(KEYINPUT58), .A2(n1159), .ZN(n1156) );
NAND2_X1 U835 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
AND4_X1 U836 ( .A1(n1162), .A2(n1112), .A3(n1163), .A4(n1164), .ZN(n1089) );
NOR4_X1 U837 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
NOR2_X1 U838 ( .A1(KEYINPUT3), .A2(n1169), .ZN(n1168) );
NOR2_X1 U839 ( .A1(KEYINPUT9), .A2(n1170), .ZN(n1167) );
NOR2_X1 U840 ( .A1(n1171), .A2(n1172), .ZN(n1166) );
NOR3_X1 U841 ( .A1(n1173), .A2(n1174), .A3(n1022), .ZN(n1165) );
AND3_X1 U842 ( .A1(n1175), .A2(n1006), .A3(n1176), .ZN(n1163) );
NAND3_X1 U843 ( .A1(n1177), .A2(n1178), .A3(n1033), .ZN(n1006) );
NAND3_X1 U844 ( .A1(n1177), .A2(n1178), .A3(n1034), .ZN(n1112) );
NAND3_X1 U845 ( .A1(n1179), .A2(n1032), .A3(n1180), .ZN(n1162) );
INV_X1 U846 ( .A(n1051), .ZN(n1032) );
NAND2_X1 U847 ( .A1(n1181), .A2(n1182), .ZN(n1179) );
NAND4_X1 U848 ( .A1(KEYINPUT9), .A2(n1177), .A3(n1183), .A4(n1184), .ZN(n1182) );
NAND4_X1 U849 ( .A1(KEYINPUT3), .A2(n1033), .A3(n1174), .A4(n1185), .ZN(n1181) );
XOR2_X1 U850 ( .A(n1186), .B(KEYINPUT44), .Z(n1140) );
XOR2_X1 U851 ( .A(n1187), .B(n1188), .Z(n1133) );
NOR2_X1 U852 ( .A1(G125), .A2(KEYINPUT7), .ZN(n1188) );
NOR2_X1 U853 ( .A1(n1077), .A2(G952), .ZN(n1096) );
XNOR2_X1 U854 ( .A(G146), .B(n1189), .ZN(G48) );
NAND4_X1 U855 ( .A1(KEYINPUT39), .A2(n1147), .A3(n1034), .A4(n1040), .ZN(n1189) );
XOR2_X1 U856 ( .A(G143), .B(n1190), .Z(G45) );
NOR2_X1 U857 ( .A1(n1171), .A2(n1148), .ZN(n1190) );
NAND3_X1 U858 ( .A1(n1183), .A2(n1184), .A3(n1158), .ZN(n1148) );
XOR2_X1 U859 ( .A(G140), .B(n1191), .Z(G42) );
NOR2_X1 U860 ( .A1(KEYINPUT1), .A2(n1142), .ZN(n1191) );
NAND4_X1 U861 ( .A1(n1034), .A2(n1046), .A3(n1192), .A4(n1053), .ZN(n1142) );
NOR2_X1 U862 ( .A1(n1160), .A2(n1027), .ZN(n1192) );
XNOR2_X1 U863 ( .A(G137), .B(n1141), .ZN(G39) );
NAND3_X1 U864 ( .A1(n1050), .A2(n1053), .A3(n1147), .ZN(n1141) );
XOR2_X1 U865 ( .A(n1193), .B(n1149), .Z(G36) );
NAND3_X1 U866 ( .A1(n1053), .A2(n1033), .A3(n1158), .ZN(n1149) );
INV_X1 U867 ( .A(n1194), .ZN(n1158) );
XOR2_X1 U868 ( .A(G131), .B(n1195), .Z(G33) );
NOR4_X1 U869 ( .A1(KEYINPUT23), .A2(n1016), .A3(n1196), .A4(n1194), .ZN(n1195) );
NAND2_X1 U870 ( .A1(n1161), .A2(n1155), .ZN(n1194) );
INV_X1 U871 ( .A(n1053), .ZN(n1016) );
NOR2_X1 U872 ( .A1(n1041), .A2(n1197), .ZN(n1053) );
NOR2_X1 U873 ( .A1(n1043), .A2(n1042), .ZN(n1197) );
INV_X1 U874 ( .A(G214), .ZN(n1043) );
XOR2_X1 U875 ( .A(n1198), .B(n1150), .Z(G30) );
NAND3_X1 U876 ( .A1(n1033), .A2(n1040), .A3(n1147), .ZN(n1150) );
NOR4_X1 U877 ( .A1(n1027), .A2(n1047), .A3(n1174), .A4(n1160), .ZN(n1147) );
INV_X1 U878 ( .A(n1155), .ZN(n1160) );
XOR2_X1 U879 ( .A(n1199), .B(n1200), .Z(G3) );
XOR2_X1 U880 ( .A(n1122), .B(KEYINPUT12), .Z(n1200) );
NAND2_X1 U881 ( .A1(n1201), .A2(n1040), .ZN(n1199) );
XOR2_X1 U882 ( .A(n1172), .B(KEYINPUT21), .Z(n1201) );
NAND3_X1 U883 ( .A1(n1050), .A2(n1202), .A3(n1161), .ZN(n1172) );
NOR3_X1 U884 ( .A1(n1048), .A2(n1047), .A3(n1027), .ZN(n1161) );
XNOR2_X1 U885 ( .A(G125), .B(n1203), .ZN(G27) );
NAND4_X1 U886 ( .A1(n1204), .A2(n1155), .A3(n1051), .A4(n1205), .ZN(n1203) );
NOR2_X1 U887 ( .A1(n1206), .A2(n1196), .ZN(n1205) );
NAND2_X1 U888 ( .A1(n1207), .A2(n1208), .ZN(n1155) );
NAND3_X1 U889 ( .A1(G902), .A2(n1049), .A3(n1063), .ZN(n1208) );
NOR2_X1 U890 ( .A1(G900), .A2(n1077), .ZN(n1063) );
XOR2_X1 U891 ( .A(KEYINPUT16), .B(n1040), .Z(n1204) );
XOR2_X1 U892 ( .A(n1209), .B(n1170), .Z(G24) );
NAND4_X1 U893 ( .A1(n1051), .A2(n1177), .A3(n1210), .A4(n1180), .ZN(n1170) );
NOR2_X1 U894 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
INV_X1 U895 ( .A(n1018), .ZN(n1177) );
NAND2_X1 U896 ( .A1(n1174), .A2(n1213), .ZN(n1018) );
XNOR2_X1 U897 ( .A(G119), .B(n1214), .ZN(G21) );
NAND4_X1 U898 ( .A1(KEYINPUT51), .A2(n1215), .A3(n1050), .A4(n1048), .ZN(n1214) );
NAND2_X1 U899 ( .A1(n1216), .A2(n1217), .ZN(G18) );
NAND2_X1 U900 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U901 ( .A(KEYINPUT49), .B(n1220), .Z(n1216) );
NOR2_X1 U902 ( .A1(n1218), .A2(n1219), .ZN(n1220) );
INV_X1 U903 ( .A(n1169), .ZN(n1218) );
NAND3_X1 U904 ( .A1(n1174), .A2(n1033), .A3(n1215), .ZN(n1169) );
NOR2_X1 U905 ( .A1(n1184), .A2(n1212), .ZN(n1033) );
INV_X1 U906 ( .A(n1183), .ZN(n1212) );
XOR2_X1 U907 ( .A(n1221), .B(KEYINPUT50), .Z(n1183) );
XOR2_X1 U908 ( .A(n1222), .B(n1175), .Z(G15) );
NAND3_X1 U909 ( .A1(n1174), .A2(n1034), .A3(n1215), .ZN(n1175) );
INV_X1 U910 ( .A(n1173), .ZN(n1215) );
NAND3_X1 U911 ( .A1(n1180), .A2(n1185), .A3(n1051), .ZN(n1173) );
NOR2_X1 U912 ( .A1(n1028), .A2(n1223), .ZN(n1051) );
NOR2_X1 U913 ( .A1(n1030), .A2(n1029), .ZN(n1223) );
INV_X1 U914 ( .A(n1224), .ZN(n1029) );
INV_X1 U915 ( .A(G221), .ZN(n1030) );
INV_X1 U916 ( .A(n1047), .ZN(n1185) );
XOR2_X1 U917 ( .A(n1225), .B(KEYINPUT27), .Z(n1047) );
INV_X1 U918 ( .A(n1196), .ZN(n1034) );
NAND2_X1 U919 ( .A1(n1221), .A2(n1184), .ZN(n1196) );
INV_X1 U920 ( .A(n1211), .ZN(n1184) );
XNOR2_X1 U921 ( .A(G110), .B(n1176), .ZN(G12) );
NAND3_X1 U922 ( .A1(n1050), .A2(n1178), .A3(n1046), .ZN(n1176) );
INV_X1 U923 ( .A(n1206), .ZN(n1046) );
NAND2_X1 U924 ( .A1(n1048), .A2(n1213), .ZN(n1206) );
XNOR2_X1 U925 ( .A(n1225), .B(KEYINPUT45), .ZN(n1213) );
XNOR2_X1 U926 ( .A(n1057), .B(G472), .ZN(n1225) );
AND2_X1 U927 ( .A1(n1226), .A2(n1186), .ZN(n1057) );
NAND3_X1 U928 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1226) );
NAND2_X1 U929 ( .A1(n1118), .A2(n1114), .ZN(n1229) );
NOR2_X1 U930 ( .A1(n1122), .A2(n1123), .ZN(n1118) );
OR3_X1 U931 ( .A1(n1114), .A2(n1230), .A3(n1122), .ZN(n1228) );
NAND2_X1 U932 ( .A1(n1231), .A2(n1122), .ZN(n1227) );
XOR2_X1 U933 ( .A(n1114), .B(n1230), .Z(n1231) );
INV_X1 U934 ( .A(n1123), .ZN(n1230) );
NAND3_X1 U935 ( .A1(n1232), .A2(n1077), .A3(G210), .ZN(n1123) );
XOR2_X1 U936 ( .A(n1233), .B(n1234), .Z(n1114) );
XOR2_X1 U937 ( .A(n1235), .B(n1236), .Z(n1234) );
XOR2_X1 U938 ( .A(n1222), .B(n1237), .Z(n1233) );
INV_X1 U939 ( .A(n1174), .ZN(n1048) );
XOR2_X1 U940 ( .A(n1058), .B(n1060), .Z(n1174) );
INV_X1 U941 ( .A(n1100), .ZN(n1060) );
NAND2_X1 U942 ( .A1(G217), .A2(n1224), .ZN(n1100) );
NAND2_X1 U943 ( .A1(n1238), .A2(n1186), .ZN(n1058) );
XOR2_X1 U944 ( .A(KEYINPUT18), .B(n1239), .Z(n1238) );
INV_X1 U945 ( .A(n1098), .ZN(n1239) );
XOR2_X1 U946 ( .A(n1240), .B(n1241), .Z(n1098) );
XNOR2_X1 U947 ( .A(n1242), .B(n1243), .ZN(n1241) );
XOR2_X1 U948 ( .A(n1244), .B(n1245), .Z(n1243) );
NOR2_X1 U949 ( .A1(KEYINPUT11), .A2(n1246), .ZN(n1245) );
XOR2_X1 U950 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U951 ( .A(G119), .B(G110), .Z(n1248) );
XOR2_X1 U952 ( .A(KEYINPUT63), .B(G128), .Z(n1247) );
NAND3_X1 U953 ( .A1(n1249), .A2(n1077), .A3(G221), .ZN(n1244) );
XOR2_X1 U954 ( .A(KEYINPUT62), .B(G234), .Z(n1249) );
XNOR2_X1 U955 ( .A(n1250), .B(n1065), .ZN(n1240) );
XOR2_X1 U956 ( .A(G125), .B(G140), .Z(n1065) );
AND2_X1 U957 ( .A1(n1180), .A2(n1023), .ZN(n1178) );
INV_X1 U958 ( .A(n1027), .ZN(n1023) );
NAND2_X1 U959 ( .A1(n1028), .A2(n1251), .ZN(n1027) );
NAND2_X1 U960 ( .A1(G221), .A2(n1224), .ZN(n1251) );
NAND2_X1 U961 ( .A1(n1252), .A2(G234), .ZN(n1224) );
XNOR2_X1 U962 ( .A(n1253), .B(G469), .ZN(n1028) );
NAND2_X1 U963 ( .A1(n1254), .A2(n1186), .ZN(n1253) );
XNOR2_X1 U964 ( .A(n1128), .B(n1255), .ZN(n1254) );
XOR2_X1 U965 ( .A(G140), .B(G110), .Z(n1255) );
XNOR2_X1 U966 ( .A(n1256), .B(n1257), .ZN(n1128) );
XOR2_X1 U967 ( .A(n1237), .B(n1258), .Z(n1257) );
XOR2_X1 U968 ( .A(n1069), .B(KEYINPUT36), .Z(n1237) );
XNOR2_X1 U969 ( .A(n1259), .B(n1242), .ZN(n1069) );
XOR2_X1 U970 ( .A(G137), .B(KEYINPUT15), .Z(n1242) );
XOR2_X1 U971 ( .A(G131), .B(n1193), .Z(n1259) );
INV_X1 U972 ( .A(G134), .ZN(n1193) );
XOR2_X1 U973 ( .A(n1067), .B(n1260), .Z(n1256) );
XOR2_X1 U974 ( .A(KEYINPUT54), .B(n1261), .Z(n1260) );
NOR2_X1 U975 ( .A1(G953), .A2(n1075), .ZN(n1261) );
INV_X1 U976 ( .A(G227), .ZN(n1075) );
XOR2_X1 U977 ( .A(n1262), .B(G128), .Z(n1067) );
NAND3_X1 U978 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1262) );
XOR2_X1 U979 ( .A(n1266), .B(KEYINPUT41), .Z(n1265) );
NAND2_X1 U980 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
OR3_X1 U981 ( .A1(n1269), .A2(G146), .A3(KEYINPUT42), .ZN(n1268) );
NAND2_X1 U982 ( .A1(n1270), .A2(KEYINPUT42), .ZN(n1267) );
OR2_X1 U983 ( .A1(n1271), .A2(KEYINPUT6), .ZN(n1264) );
NAND3_X1 U984 ( .A1(G146), .A2(n1269), .A3(KEYINPUT6), .ZN(n1263) );
INV_X1 U985 ( .A(n1272), .ZN(n1269) );
AND2_X1 U986 ( .A1(n1040), .A2(n1202), .ZN(n1180) );
NAND2_X1 U987 ( .A1(n1207), .A2(n1273), .ZN(n1202) );
NAND4_X1 U988 ( .A1(G953), .A2(G902), .A3(n1049), .A4(n1085), .ZN(n1273) );
INV_X1 U989 ( .A(G898), .ZN(n1085) );
NAND3_X1 U990 ( .A1(n1049), .A2(n1077), .A3(n1274), .ZN(n1207) );
XNOR2_X1 U991 ( .A(G952), .B(KEYINPUT55), .ZN(n1274) );
NAND2_X1 U992 ( .A1(G237), .A2(G234), .ZN(n1049) );
INV_X1 U993 ( .A(n1171), .ZN(n1040) );
NAND2_X1 U994 ( .A1(n1041), .A2(n1275), .ZN(n1171) );
NAND2_X1 U995 ( .A1(G214), .A2(n1276), .ZN(n1275) );
XNOR2_X1 U996 ( .A(n1277), .B(n1278), .ZN(n1041) );
NOR2_X1 U997 ( .A1(n1042), .A2(n1279), .ZN(n1278) );
XOR2_X1 U998 ( .A(n1139), .B(KEYINPUT38), .Z(n1279) );
INV_X1 U999 ( .A(G210), .ZN(n1139) );
INV_X1 U1000 ( .A(n1276), .ZN(n1042) );
NAND2_X1 U1001 ( .A1(n1252), .A2(n1232), .ZN(n1276) );
XOR2_X1 U1002 ( .A(KEYINPUT28), .B(n1186), .Z(n1252) );
NAND2_X1 U1003 ( .A1(n1280), .A2(n1186), .ZN(n1277) );
XOR2_X1 U1004 ( .A(n1138), .B(n1281), .Z(n1280) );
NAND2_X1 U1005 ( .A1(n1282), .A2(KEYINPUT25), .ZN(n1281) );
XOR2_X1 U1006 ( .A(n1283), .B(n1235), .Z(n1282) );
INV_X1 U1007 ( .A(n1187), .ZN(n1235) );
XOR2_X1 U1008 ( .A(n1284), .B(G128), .Z(n1187) );
NAND3_X1 U1009 ( .A1(n1285), .A2(n1271), .A3(KEYINPUT57), .ZN(n1284) );
INV_X1 U1010 ( .A(n1270), .ZN(n1271) );
NOR2_X1 U1011 ( .A1(n1272), .A2(G146), .ZN(n1270) );
NAND2_X1 U1012 ( .A1(n1272), .A2(G146), .ZN(n1285) );
XNOR2_X1 U1013 ( .A(G143), .B(KEYINPUT4), .ZN(n1272) );
XNOR2_X1 U1014 ( .A(G125), .B(n1286), .ZN(n1283) );
NOR2_X1 U1015 ( .A1(G953), .A2(n1084), .ZN(n1286) );
INV_X1 U1016 ( .A(G224), .ZN(n1084) );
NAND2_X1 U1017 ( .A1(n1287), .A2(n1288), .ZN(n1138) );
NAND2_X1 U1018 ( .A1(n1289), .A2(n1093), .ZN(n1288) );
XOR2_X1 U1019 ( .A(KEYINPUT26), .B(n1290), .Z(n1287) );
NOR2_X1 U1020 ( .A1(n1093), .A2(n1289), .ZN(n1290) );
XOR2_X1 U1021 ( .A(n1291), .B(n1258), .Z(n1289) );
INV_X1 U1022 ( .A(n1095), .ZN(n1258) );
XOR2_X1 U1023 ( .A(n1122), .B(n1292), .Z(n1095) );
XOR2_X1 U1024 ( .A(G107), .B(G104), .Z(n1292) );
INV_X1 U1025 ( .A(G101), .ZN(n1122) );
NOR2_X1 U1026 ( .A1(KEYINPUT31), .A2(n1094), .ZN(n1291) );
XNOR2_X1 U1027 ( .A(G113), .B(n1293), .ZN(n1094) );
NOR2_X1 U1028 ( .A1(KEYINPUT5), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1029 ( .A(KEYINPUT17), .B(n1236), .Z(n1294) );
XOR2_X1 U1030 ( .A(G119), .B(n1295), .Z(n1236) );
XOR2_X1 U1031 ( .A(G122), .B(n1296), .Z(n1093) );
NOR2_X1 U1032 ( .A1(G110), .A2(KEYINPUT53), .ZN(n1296) );
INV_X1 U1033 ( .A(n1022), .ZN(n1050) );
NAND2_X1 U1034 ( .A1(n1211), .A2(n1221), .ZN(n1022) );
XOR2_X1 U1035 ( .A(n1297), .B(G478), .Z(n1221) );
OR2_X1 U1036 ( .A1(n1104), .A2(G902), .ZN(n1297) );
XNOR2_X1 U1037 ( .A(n1298), .B(n1299), .ZN(n1104) );
XOR2_X1 U1038 ( .A(G107), .B(n1300), .Z(n1299) );
XOR2_X1 U1039 ( .A(G143), .B(G134), .Z(n1300) );
XOR2_X1 U1040 ( .A(n1301), .B(n1302), .Z(n1298) );
XOR2_X1 U1041 ( .A(n1303), .B(n1304), .Z(n1302) );
AND3_X1 U1042 ( .A1(G234), .A2(n1077), .A3(G217), .ZN(n1304) );
NOR2_X1 U1043 ( .A1(KEYINPUT40), .A2(n1305), .ZN(n1303) );
XNOR2_X1 U1044 ( .A(n1295), .B(n1306), .ZN(n1305) );
NOR2_X1 U1045 ( .A1(KEYINPUT52), .A2(n1209), .ZN(n1306) );
XNOR2_X1 U1046 ( .A(n1219), .B(KEYINPUT59), .ZN(n1295) );
INV_X1 U1047 ( .A(G116), .ZN(n1219) );
NAND2_X1 U1048 ( .A1(KEYINPUT22), .A2(n1198), .ZN(n1301) );
INV_X1 U1049 ( .A(G128), .ZN(n1198) );
XOR2_X1 U1050 ( .A(n1307), .B(G475), .Z(n1211) );
NAND2_X1 U1051 ( .A1(n1110), .A2(n1186), .ZN(n1307) );
INV_X1 U1052 ( .A(G902), .ZN(n1186) );
XNOR2_X1 U1053 ( .A(n1308), .B(n1309), .ZN(n1110) );
XOR2_X1 U1054 ( .A(n1310), .B(n1311), .Z(n1309) );
NAND2_X1 U1055 ( .A1(KEYINPUT61), .A2(n1222), .ZN(n1311) );
INV_X1 U1056 ( .A(G113), .ZN(n1222) );
NAND3_X1 U1057 ( .A1(n1312), .A2(n1313), .A3(n1314), .ZN(n1310) );
NAND2_X1 U1058 ( .A1(KEYINPUT34), .A2(n1315), .ZN(n1314) );
NAND3_X1 U1059 ( .A1(n1316), .A2(n1317), .A3(n1318), .ZN(n1313) );
INV_X1 U1060 ( .A(KEYINPUT34), .ZN(n1317) );
OR2_X1 U1061 ( .A1(n1318), .A2(n1316), .ZN(n1312) );
NOR2_X1 U1062 ( .A1(n1319), .A2(n1315), .ZN(n1316) );
XNOR2_X1 U1063 ( .A(n1320), .B(n1250), .ZN(n1315) );
XOR2_X1 U1064 ( .A(G146), .B(KEYINPUT30), .Z(n1250) );
XOR2_X1 U1065 ( .A(n1321), .B(KEYINPUT14), .Z(n1320) );
NAND2_X1 U1066 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NAND2_X1 U1067 ( .A1(G125), .A2(n1129), .ZN(n1323) );
XOR2_X1 U1068 ( .A(KEYINPUT37), .B(n1324), .Z(n1322) );
NOR2_X1 U1069 ( .A1(G125), .A2(n1129), .ZN(n1324) );
INV_X1 U1070 ( .A(G140), .ZN(n1129) );
INV_X1 U1071 ( .A(KEYINPUT24), .ZN(n1319) );
XOR2_X1 U1072 ( .A(n1325), .B(n1326), .Z(n1318) );
XOR2_X1 U1073 ( .A(G143), .B(n1327), .Z(n1326) );
NOR2_X1 U1074 ( .A1(KEYINPUT8), .A2(G131), .ZN(n1327) );
NAND3_X1 U1075 ( .A1(n1232), .A2(n1077), .A3(n1328), .ZN(n1325) );
XOR2_X1 U1076 ( .A(KEYINPUT29), .B(G214), .Z(n1328) );
INV_X1 U1077 ( .A(G953), .ZN(n1077) );
INV_X1 U1078 ( .A(G237), .ZN(n1232) );
XOR2_X1 U1079 ( .A(G104), .B(n1209), .Z(n1308) );
INV_X1 U1080 ( .A(G122), .ZN(n1209) );
endmodule


