//Key = 1010100111000011100000100010000001111101110101111110000010101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339;

XOR2_X1 U735 ( .A(n1013), .B(n1014), .Z(G9) );
XNOR2_X1 U736 ( .A(KEYINPUT50), .B(n1015), .ZN(n1014) );
NOR2_X1 U737 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U738 ( .A1(G953), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1017) );
NOR3_X1 U739 ( .A1(n1021), .A2(KEYINPUT38), .A3(n1022), .ZN(n1019) );
INV_X1 U740 ( .A(n1023), .ZN(n1022) );
NOR2_X1 U741 ( .A1(n1024), .A2(n1025), .ZN(n1021) );
NOR3_X1 U742 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
NOR3_X1 U743 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1027) );
NOR2_X1 U744 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U745 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U746 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR3_X1 U747 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1030) );
NOR2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1029) );
XNOR2_X1 U749 ( .A(n1043), .B(KEYINPUT5), .ZN(n1041) );
NOR3_X1 U750 ( .A1(n1039), .A2(n1044), .A3(n1033), .ZN(n1024) );
NOR3_X1 U751 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
AND2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U753 ( .A1(n1050), .A2(n1028), .ZN(n1046) );
INV_X1 U754 ( .A(n1051), .ZN(n1028) );
NOR3_X1 U755 ( .A1(n1018), .A2(G953), .A3(G952), .ZN(n1016) );
AND4_X1 U756 ( .A1(n1043), .A2(n1052), .A3(n1053), .A4(n1054), .ZN(n1018) );
NOR3_X1 U757 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
XNOR2_X1 U758 ( .A(n1058), .B(KEYINPUT35), .ZN(n1057) );
XNOR2_X1 U759 ( .A(n1059), .B(n1060), .ZN(n1056) );
NOR2_X1 U760 ( .A1(KEYINPUT53), .A2(n1061), .ZN(n1060) );
XNOR2_X1 U761 ( .A(G475), .B(KEYINPUT37), .ZN(n1061) );
XNOR2_X1 U762 ( .A(n1062), .B(G478), .ZN(n1053) );
XOR2_X1 U763 ( .A(n1063), .B(n1064), .Z(G72) );
NOR3_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NOR2_X1 U765 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NOR2_X1 U766 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U767 ( .A1(G140), .A2(n1072), .ZN(n1071) );
XNOR2_X1 U768 ( .A(KEYINPUT42), .B(G125), .ZN(n1072) );
XOR2_X1 U769 ( .A(n1073), .B(KEYINPUT39), .Z(n1065) );
NAND4_X1 U770 ( .A1(n1069), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1073) );
OR3_X1 U771 ( .A1(n1077), .A2(G140), .A3(KEYINPUT42), .ZN(n1076) );
NAND2_X1 U772 ( .A1(KEYINPUT42), .A2(n1077), .ZN(n1075) );
XOR2_X1 U773 ( .A(n1078), .B(n1079), .Z(n1069) );
NOR2_X1 U774 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U776 ( .A(G131), .B(KEYINPUT6), .ZN(n1083) );
AND2_X1 U777 ( .A1(n1084), .A2(n1082), .ZN(n1080) );
XOR2_X1 U778 ( .A(G137), .B(n1085), .Z(n1082) );
NOR2_X1 U779 ( .A1(G134), .A2(KEYINPUT52), .ZN(n1085) );
NAND2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1063) );
NAND2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U782 ( .A(n1090), .B(KEYINPUT22), .Z(n1086) );
NAND2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U784 ( .A1(G953), .A2(n1093), .ZN(n1092) );
NAND2_X1 U785 ( .A1(G227), .A2(n1094), .ZN(n1093) );
NAND2_X1 U786 ( .A1(G900), .A2(n1095), .ZN(n1094) );
INV_X1 U787 ( .A(KEYINPUT0), .ZN(n1095) );
NAND2_X1 U788 ( .A1(KEYINPUT0), .A2(n1066), .ZN(n1091) );
XOR2_X1 U789 ( .A(n1096), .B(n1097), .Z(G69) );
XOR2_X1 U790 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U791 ( .A1(G953), .A2(n1100), .ZN(n1099) );
NAND2_X1 U792 ( .A1(G898), .A2(G224), .ZN(n1100) );
NAND2_X1 U793 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U794 ( .A1(G953), .A2(n1103), .ZN(n1102) );
XOR2_X1 U795 ( .A(n1104), .B(n1105), .Z(n1101) );
XNOR2_X1 U796 ( .A(n1106), .B(KEYINPUT60), .ZN(n1105) );
NAND2_X1 U797 ( .A1(n1107), .A2(KEYINPUT46), .ZN(n1106) );
XNOR2_X1 U798 ( .A(n1108), .B(KEYINPUT3), .ZN(n1107) );
AND2_X1 U799 ( .A1(n1109), .A2(n1089), .ZN(n1096) );
NOR2_X1 U800 ( .A1(n1110), .A2(n1111), .ZN(G66) );
NOR2_X1 U801 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U803 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
AND2_X1 U805 ( .A1(n1117), .A2(n1116), .ZN(n1112) );
INV_X1 U806 ( .A(KEYINPUT14), .ZN(n1117) );
NOR2_X1 U807 ( .A1(n1110), .A2(n1120), .ZN(G63) );
NOR3_X1 U808 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
NOR2_X1 U809 ( .A1(KEYINPUT58), .A2(n1124), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1062), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n1130), .A2(n1131), .ZN(n1128) );
NOR3_X1 U814 ( .A1(n1132), .A2(n1133), .A3(n1131), .ZN(n1121) );
NOR2_X1 U815 ( .A1(n1126), .A2(n1134), .ZN(n1133) );
XNOR2_X1 U816 ( .A(n1124), .B(n1135), .ZN(n1134) );
XOR2_X1 U817 ( .A(KEYINPUT4), .B(KEYINPUT2), .Z(n1135) );
INV_X1 U818 ( .A(n1129), .ZN(n1124) );
INV_X1 U819 ( .A(KEYINPUT58), .ZN(n1126) );
NOR2_X1 U820 ( .A1(n1110), .A2(n1136), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1059), .A2(n1137), .A3(n1138), .ZN(n1136) );
AND3_X1 U822 ( .A1(n1139), .A2(G475), .A3(n1118), .ZN(n1138) );
NOR2_X1 U823 ( .A1(n1140), .A2(n1139), .ZN(n1137) );
AND2_X1 U824 ( .A1(n1020), .A2(G475), .ZN(n1140) );
INV_X1 U825 ( .A(n1130), .ZN(n1020) );
NAND2_X1 U826 ( .A1(n1141), .A2(n1142), .ZN(G6) );
NAND3_X1 U827 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1142) );
NAND2_X1 U828 ( .A1(G104), .A2(n1146), .ZN(n1141) );
NAND2_X1 U829 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U830 ( .A1(KEYINPUT23), .A2(n1143), .ZN(n1148) );
NAND2_X1 U831 ( .A1(n1149), .A2(n1150), .ZN(n1147) );
INV_X1 U832 ( .A(KEYINPUT23), .ZN(n1150) );
NAND2_X1 U833 ( .A1(n1143), .A2(n1144), .ZN(n1149) );
INV_X1 U834 ( .A(KEYINPUT21), .ZN(n1144) );
AND4_X1 U835 ( .A1(n1151), .A2(n1051), .A3(n1152), .A4(n1153), .ZN(n1143) );
XNOR2_X1 U836 ( .A(KEYINPUT31), .B(n1154), .ZN(n1153) );
NOR3_X1 U837 ( .A1(n1110), .A2(n1155), .A3(n1156), .ZN(G57) );
NOR3_X1 U838 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
NOR2_X1 U839 ( .A1(n1160), .A2(n1161), .ZN(n1155) );
NOR2_X1 U840 ( .A1(n1158), .A2(n1159), .ZN(n1161) );
XOR2_X1 U841 ( .A(n1162), .B(KEYINPUT7), .Z(n1159) );
NAND2_X1 U842 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U843 ( .A1(n1164), .A2(n1163), .ZN(n1158) );
AND2_X1 U844 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
NAND2_X1 U845 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1170), .ZN(n1165) );
XNOR2_X1 U847 ( .A(n1167), .B(KEYINPUT57), .ZN(n1170) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(n1167) );
NAND2_X1 U849 ( .A1(n1118), .A2(G472), .ZN(n1164) );
INV_X1 U850 ( .A(n1157), .ZN(n1160) );
NAND2_X1 U851 ( .A1(n1173), .A2(n1174), .ZN(n1157) );
OR2_X1 U852 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U853 ( .A(n1177), .B(KEYINPUT19), .Z(n1173) );
NAND2_X1 U854 ( .A1(n1176), .A2(n1175), .ZN(n1177) );
INV_X1 U855 ( .A(G101), .ZN(n1176) );
NOR2_X1 U856 ( .A1(n1110), .A2(n1178), .ZN(G54) );
XOR2_X1 U857 ( .A(n1179), .B(n1180), .Z(n1178) );
XNOR2_X1 U858 ( .A(n1181), .B(n1182), .ZN(n1180) );
XNOR2_X1 U859 ( .A(n1183), .B(G110), .ZN(n1182) );
XNOR2_X1 U860 ( .A(n1184), .B(n1185), .ZN(n1179) );
XNOR2_X1 U861 ( .A(n1186), .B(n1187), .ZN(n1185) );
NOR2_X1 U862 ( .A1(KEYINPUT20), .A2(n1171), .ZN(n1187) );
NAND3_X1 U863 ( .A1(n1118), .A2(G469), .A3(KEYINPUT16), .ZN(n1186) );
NOR3_X1 U864 ( .A1(n1110), .A2(n1188), .A3(n1189), .ZN(G51) );
NOR4_X1 U865 ( .A1(n1190), .A2(n1132), .A3(KEYINPUT55), .A4(n1191), .ZN(n1189) );
NOR2_X1 U866 ( .A1(n1192), .A2(n1193), .ZN(n1188) );
NOR3_X1 U867 ( .A1(n1132), .A2(n1194), .A3(n1191), .ZN(n1193) );
NOR2_X1 U868 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
INV_X1 U869 ( .A(KEYINPUT55), .ZN(n1196) );
INV_X1 U870 ( .A(n1118), .ZN(n1132) );
NOR2_X1 U871 ( .A1(n1197), .A2(n1130), .ZN(n1118) );
NOR2_X1 U872 ( .A1(n1109), .A2(n1088), .ZN(n1130) );
NAND4_X1 U873 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1088) );
NOR3_X1 U874 ( .A1(n1202), .A2(n1203), .A3(n1204), .ZN(n1201) );
NAND2_X1 U875 ( .A1(n1052), .A2(n1205), .ZN(n1200) );
NAND3_X1 U876 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1205) );
XOR2_X1 U877 ( .A(KEYINPUT36), .B(n1209), .Z(n1208) );
NOR2_X1 U878 ( .A1(n1154), .A2(n1210), .ZN(n1209) );
NAND3_X1 U879 ( .A1(n1151), .A2(n1048), .A3(n1211), .ZN(n1207) );
XOR2_X1 U880 ( .A(KEYINPUT8), .B(n1212), .Z(n1206) );
NAND4_X1 U881 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1109) );
AND4_X1 U882 ( .A1(n1013), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1216) );
NAND3_X1 U883 ( .A1(n1220), .A2(n1221), .A3(n1051), .ZN(n1013) );
NAND2_X1 U884 ( .A1(n1221), .A2(n1045), .ZN(n1215) );
NAND2_X1 U885 ( .A1(n1222), .A2(n1223), .ZN(n1045) );
NAND3_X1 U886 ( .A1(n1224), .A2(n1225), .A3(n1049), .ZN(n1223) );
NAND2_X1 U887 ( .A1(n1151), .A2(n1051), .ZN(n1222) );
INV_X1 U888 ( .A(n1190), .ZN(n1192) );
NAND2_X1 U889 ( .A1(n1195), .A2(KEYINPUT48), .ZN(n1190) );
XOR2_X1 U890 ( .A(n1226), .B(n1227), .Z(n1195) );
XOR2_X1 U891 ( .A(n1228), .B(KEYINPUT34), .Z(n1227) );
AND2_X1 U892 ( .A1(n1229), .A2(G953), .ZN(n1110) );
XNOR2_X1 U893 ( .A(G952), .B(KEYINPUT61), .ZN(n1229) );
XNOR2_X1 U894 ( .A(G146), .B(n1198), .ZN(G48) );
NAND3_X1 U895 ( .A1(n1151), .A2(n1230), .A3(n1231), .ZN(n1198) );
XNOR2_X1 U896 ( .A(G143), .B(n1199), .ZN(G45) );
NAND3_X1 U897 ( .A1(n1211), .A2(n1048), .A3(n1232), .ZN(n1199) );
NOR3_X1 U898 ( .A1(n1042), .A2(n1233), .A3(n1234), .ZN(n1232) );
XNOR2_X1 U899 ( .A(G140), .B(n1235), .ZN(G42) );
NAND3_X1 U900 ( .A1(n1236), .A2(n1052), .A3(n1237), .ZN(n1235) );
XNOR2_X1 U901 ( .A(n1035), .B(KEYINPUT49), .ZN(n1237) );
INV_X1 U902 ( .A(n1210), .ZN(n1236) );
XNOR2_X1 U903 ( .A(G137), .B(n1238), .ZN(G39) );
NAND2_X1 U904 ( .A1(n1212), .A2(n1052), .ZN(n1238) );
AND2_X1 U905 ( .A1(n1231), .A2(n1049), .ZN(n1212) );
XNOR2_X1 U906 ( .A(n1202), .B(n1239), .ZN(G36) );
NAND2_X1 U907 ( .A1(KEYINPUT9), .A2(G134), .ZN(n1239) );
AND4_X1 U908 ( .A1(n1211), .A2(n1048), .A3(n1052), .A4(n1220), .ZN(n1202) );
XNOR2_X1 U909 ( .A(G131), .B(n1240), .ZN(G33) );
NAND4_X1 U910 ( .A1(n1211), .A2(n1151), .A3(n1052), .A4(n1241), .ZN(n1240) );
XOR2_X1 U911 ( .A(KEYINPUT59), .B(n1048), .Z(n1241) );
INV_X1 U912 ( .A(n1033), .ZN(n1052) );
NAND2_X1 U913 ( .A1(n1242), .A2(n1038), .ZN(n1033) );
INV_X1 U914 ( .A(n1040), .ZN(n1242) );
XOR2_X1 U915 ( .A(G128), .B(n1204), .Z(G30) );
AND3_X1 U916 ( .A1(n1220), .A2(n1230), .A3(n1231), .ZN(n1204) );
AND3_X1 U917 ( .A1(n1243), .A2(n1225), .A3(n1211), .ZN(n1231) );
AND2_X1 U918 ( .A1(n1244), .A2(n1035), .ZN(n1211) );
XNOR2_X1 U919 ( .A(G101), .B(n1213), .ZN(G3) );
NAND3_X1 U920 ( .A1(n1048), .A2(n1221), .A3(n1049), .ZN(n1213) );
XNOR2_X1 U921 ( .A(n1077), .B(n1203), .ZN(G27) );
NOR3_X1 U922 ( .A1(n1039), .A2(n1042), .A3(n1210), .ZN(n1203) );
NAND4_X1 U923 ( .A1(n1244), .A2(n1151), .A3(n1224), .A4(n1225), .ZN(n1210) );
AND2_X1 U924 ( .A1(n1245), .A2(n1023), .ZN(n1244) );
NAND2_X1 U925 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U926 ( .A1(n1066), .A2(G902), .ZN(n1247) );
NOR2_X1 U927 ( .A1(n1089), .A2(G900), .ZN(n1066) );
NAND2_X1 U928 ( .A1(G952), .A2(n1089), .ZN(n1246) );
XNOR2_X1 U929 ( .A(G122), .B(n1214), .ZN(G24) );
NAND4_X1 U930 ( .A1(n1248), .A2(n1051), .A3(n1249), .A4(n1250), .ZN(n1214) );
NOR2_X1 U931 ( .A1(n1058), .A2(n1225), .ZN(n1051) );
XNOR2_X1 U932 ( .A(G119), .B(n1219), .ZN(G21) );
NAND4_X1 U933 ( .A1(n1049), .A2(n1248), .A3(n1243), .A4(n1225), .ZN(n1219) );
XNOR2_X1 U934 ( .A(n1224), .B(KEYINPUT54), .ZN(n1243) );
INV_X1 U935 ( .A(n1026), .ZN(n1049) );
XNOR2_X1 U936 ( .A(G116), .B(n1218), .ZN(G18) );
NAND3_X1 U937 ( .A1(n1248), .A2(n1220), .A3(n1048), .ZN(n1218) );
INV_X1 U938 ( .A(n1050), .ZN(n1220) );
NAND2_X1 U939 ( .A1(n1251), .A2(n1250), .ZN(n1050) );
XNOR2_X1 U940 ( .A(G113), .B(n1217), .ZN(G15) );
NAND3_X1 U941 ( .A1(n1048), .A2(n1248), .A3(n1151), .ZN(n1217) );
NOR2_X1 U942 ( .A1(n1250), .A2(n1234), .ZN(n1151) );
INV_X1 U943 ( .A(n1249), .ZN(n1234) );
XNOR2_X1 U944 ( .A(n1251), .B(KEYINPUT13), .ZN(n1249) );
AND2_X1 U945 ( .A1(n1043), .A2(n1152), .ZN(n1248) );
INV_X1 U946 ( .A(n1039), .ZN(n1043) );
NAND2_X1 U947 ( .A1(n1252), .A2(n1037), .ZN(n1039) );
INV_X1 U948 ( .A(n1036), .ZN(n1252) );
NOR2_X1 U949 ( .A1(n1225), .A2(n1224), .ZN(n1048) );
XNOR2_X1 U950 ( .A(G110), .B(n1253), .ZN(G12) );
NAND4_X1 U951 ( .A1(n1224), .A2(n1221), .A3(n1254), .A4(n1225), .ZN(n1253) );
XOR2_X1 U952 ( .A(n1055), .B(KEYINPUT1), .Z(n1225) );
XNOR2_X1 U953 ( .A(n1255), .B(n1119), .ZN(n1055) );
AND2_X1 U954 ( .A1(G217), .A2(n1256), .ZN(n1119) );
NAND2_X1 U955 ( .A1(n1197), .A2(n1116), .ZN(n1255) );
NAND2_X1 U956 ( .A1(n1257), .A2(n1258), .ZN(n1116) );
NAND2_X1 U957 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U958 ( .A(n1261), .B(KEYINPUT10), .Z(n1257) );
OR2_X1 U959 ( .A1(n1260), .A2(n1259), .ZN(n1261) );
XOR2_X1 U960 ( .A(n1262), .B(G137), .Z(n1259) );
NAND2_X1 U961 ( .A1(G221), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U962 ( .A(n1264), .B(n1265), .ZN(n1260) );
XOR2_X1 U963 ( .A(G119), .B(G110), .Z(n1265) );
XOR2_X1 U964 ( .A(n1266), .B(n1267), .Z(n1264) );
NAND2_X1 U965 ( .A1(KEYINPUT63), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U966 ( .A(KEYINPUT11), .B(n1026), .ZN(n1254) );
NAND2_X1 U967 ( .A1(n1233), .A2(n1251), .ZN(n1026) );
XNOR2_X1 U968 ( .A(n1059), .B(G475), .ZN(n1251) );
NOR2_X1 U969 ( .A1(n1139), .A2(G902), .ZN(n1059) );
XOR2_X1 U970 ( .A(n1269), .B(n1270), .Z(n1139) );
XOR2_X1 U971 ( .A(n1271), .B(n1272), .Z(n1270) );
XNOR2_X1 U972 ( .A(n1273), .B(n1274), .ZN(n1272) );
NOR2_X1 U973 ( .A1(KEYINPUT28), .A2(n1275), .ZN(n1274) );
XNOR2_X1 U974 ( .A(KEYINPUT62), .B(n1268), .ZN(n1275) );
NAND2_X1 U975 ( .A1(n1074), .A2(n1276), .ZN(n1268) );
NAND2_X1 U976 ( .A1(G125), .A2(n1183), .ZN(n1276) );
INV_X1 U977 ( .A(n1070), .ZN(n1074) );
NOR2_X1 U978 ( .A1(n1183), .A2(G125), .ZN(n1070) );
NAND4_X1 U979 ( .A1(KEYINPUT33), .A2(G214), .A3(n1277), .A4(n1089), .ZN(n1273) );
XNOR2_X1 U980 ( .A(G113), .B(n1145), .ZN(n1271) );
INV_X1 U981 ( .A(G104), .ZN(n1145) );
XOR2_X1 U982 ( .A(n1278), .B(n1279), .Z(n1269) );
XNOR2_X1 U983 ( .A(n1084), .B(G122), .ZN(n1279) );
INV_X1 U984 ( .A(G131), .ZN(n1084) );
XNOR2_X1 U985 ( .A(G146), .B(G143), .ZN(n1278) );
INV_X1 U986 ( .A(n1250), .ZN(n1233) );
XNOR2_X1 U987 ( .A(n1280), .B(n1281), .ZN(n1250) );
XNOR2_X1 U988 ( .A(KEYINPUT41), .B(n1131), .ZN(n1281) );
INV_X1 U989 ( .A(G478), .ZN(n1131) );
NAND2_X1 U990 ( .A1(KEYINPUT15), .A2(n1282), .ZN(n1280) );
INV_X1 U991 ( .A(n1062), .ZN(n1282) );
NOR2_X1 U992 ( .A1(n1129), .A2(G902), .ZN(n1062) );
XNOR2_X1 U993 ( .A(n1283), .B(n1284), .ZN(n1129) );
XOR2_X1 U994 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U995 ( .A(G128), .B(n1287), .ZN(n1286) );
NAND2_X1 U996 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U997 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U998 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
NAND2_X1 U999 ( .A1(KEYINPUT45), .A2(n1015), .ZN(n1293) );
INV_X1 U1000 ( .A(KEYINPUT30), .ZN(n1292) );
NAND2_X1 U1001 ( .A1(G107), .A2(n1294), .ZN(n1288) );
NAND2_X1 U1002 ( .A1(KEYINPUT45), .A2(n1295), .ZN(n1294) );
OR2_X1 U1003 ( .A1(n1290), .A2(KEYINPUT30), .ZN(n1295) );
XOR2_X1 U1004 ( .A(G116), .B(G122), .Z(n1290) );
AND2_X1 U1005 ( .A1(G217), .A2(n1263), .ZN(n1285) );
AND2_X1 U1006 ( .A1(G234), .A2(n1089), .ZN(n1263) );
XNOR2_X1 U1007 ( .A(G134), .B(n1296), .ZN(n1283) );
XNOR2_X1 U1008 ( .A(KEYINPUT18), .B(n1297), .ZN(n1296) );
INV_X1 U1009 ( .A(G143), .ZN(n1297) );
AND2_X1 U1010 ( .A1(n1152), .A2(n1035), .ZN(n1221) );
INV_X1 U1011 ( .A(n1154), .ZN(n1035) );
NAND2_X1 U1012 ( .A1(n1036), .A2(n1037), .ZN(n1154) );
NAND2_X1 U1013 ( .A1(G221), .A2(n1298), .ZN(n1037) );
XNOR2_X1 U1014 ( .A(KEYINPUT40), .B(n1256), .ZN(n1298) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1197), .ZN(n1256) );
XNOR2_X1 U1016 ( .A(n1299), .B(G469), .ZN(n1036) );
NAND2_X1 U1017 ( .A1(n1300), .A2(n1197), .ZN(n1299) );
XOR2_X1 U1018 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1019 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1020 ( .A(n1181), .B(n1305), .Z(n1304) );
NOR2_X1 U1021 ( .A1(KEYINPUT25), .A2(n1306), .ZN(n1305) );
XNOR2_X1 U1022 ( .A(n1307), .B(n1308), .ZN(n1306) );
INV_X1 U1023 ( .A(n1184), .ZN(n1308) );
XOR2_X1 U1024 ( .A(n1078), .B(n1309), .Z(n1184) );
INV_X1 U1025 ( .A(n1108), .ZN(n1309) );
XOR2_X1 U1026 ( .A(n1310), .B(n1267), .Z(n1078) );
NAND2_X1 U1027 ( .A1(n1311), .A2(KEYINPUT43), .ZN(n1310) );
XNOR2_X1 U1028 ( .A(G143), .B(KEYINPUT29), .ZN(n1311) );
NOR2_X1 U1029 ( .A1(KEYINPUT27), .A2(n1312), .ZN(n1307) );
NAND2_X1 U1030 ( .A1(G227), .A2(n1089), .ZN(n1181) );
NAND2_X1 U1031 ( .A1(KEYINPUT26), .A2(n1183), .ZN(n1303) );
INV_X1 U1032 ( .A(G140), .ZN(n1183) );
XNOR2_X1 U1033 ( .A(G110), .B(n1313), .ZN(n1301) );
XNOR2_X1 U1034 ( .A(KEYINPUT51), .B(KEYINPUT47), .ZN(n1313) );
AND2_X1 U1035 ( .A1(n1230), .A2(n1314), .ZN(n1152) );
NAND2_X1 U1036 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND3_X1 U1037 ( .A1(n1317), .A2(n1318), .A3(n1023), .ZN(n1316) );
OR2_X1 U1038 ( .A1(G952), .A2(G953), .ZN(n1318) );
NAND2_X1 U1039 ( .A1(G953), .A2(n1319), .ZN(n1317) );
OR3_X1 U1040 ( .A1(G898), .A2(KEYINPUT32), .A3(n1197), .ZN(n1319) );
NAND2_X1 U1041 ( .A1(KEYINPUT32), .A2(n1320), .ZN(n1315) );
NAND4_X1 U1042 ( .A1(G953), .A2(G902), .A3(n1023), .A4(n1103), .ZN(n1320) );
INV_X1 U1043 ( .A(G898), .ZN(n1103) );
NAND2_X1 U1044 ( .A1(G237), .A2(G234), .ZN(n1023) );
INV_X1 U1045 ( .A(n1042), .ZN(n1230) );
NAND2_X1 U1046 ( .A1(n1040), .A2(n1038), .ZN(n1042) );
NAND2_X1 U1047 ( .A1(G214), .A2(n1321), .ZN(n1038) );
XOR2_X1 U1048 ( .A(n1322), .B(n1191), .Z(n1040) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1321), .ZN(n1191) );
NAND2_X1 U1050 ( .A1(n1277), .A2(n1197), .ZN(n1321) );
NAND2_X1 U1051 ( .A1(n1323), .A2(n1197), .ZN(n1322) );
XOR2_X1 U1052 ( .A(n1226), .B(n1324), .Z(n1323) );
XOR2_X1 U1053 ( .A(n1325), .B(KEYINPUT12), .Z(n1324) );
NAND2_X1 U1054 ( .A1(KEYINPUT56), .A2(n1228), .ZN(n1325) );
AND2_X1 U1055 ( .A1(G224), .A2(n1089), .ZN(n1228) );
XOR2_X1 U1056 ( .A(n1326), .B(n1327), .Z(n1226) );
XNOR2_X1 U1057 ( .A(n1077), .B(n1108), .ZN(n1327) );
XOR2_X1 U1058 ( .A(G101), .B(n1328), .Z(n1108) );
XNOR2_X1 U1059 ( .A(n1015), .B(G104), .ZN(n1328) );
INV_X1 U1060 ( .A(G107), .ZN(n1015) );
INV_X1 U1061 ( .A(G125), .ZN(n1077) );
XNOR2_X1 U1062 ( .A(n1104), .B(n1168), .ZN(n1326) );
INV_X1 U1063 ( .A(n1169), .ZN(n1168) );
XOR2_X1 U1064 ( .A(n1329), .B(n1172), .Z(n1104) );
XNOR2_X1 U1065 ( .A(G110), .B(G122), .ZN(n1329) );
INV_X1 U1066 ( .A(n1058), .ZN(n1224) );
XNOR2_X1 U1067 ( .A(n1330), .B(G472), .ZN(n1058) );
NAND2_X1 U1068 ( .A1(n1331), .A2(n1197), .ZN(n1330) );
INV_X1 U1069 ( .A(G902), .ZN(n1197) );
XOR2_X1 U1070 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1071 ( .A(n1175), .B(n1172), .ZN(n1333) );
XNOR2_X1 U1072 ( .A(n1334), .B(n1335), .ZN(n1172) );
XOR2_X1 U1073 ( .A(KEYINPUT44), .B(G119), .Z(n1335) );
XNOR2_X1 U1074 ( .A(G113), .B(G116), .ZN(n1334) );
NAND3_X1 U1075 ( .A1(n1277), .A2(n1089), .A3(G210), .ZN(n1175) );
INV_X1 U1076 ( .A(G953), .ZN(n1089) );
INV_X1 U1077 ( .A(G237), .ZN(n1277) );
XOR2_X1 U1078 ( .A(n1336), .B(n1337), .Z(n1332) );
NOR2_X1 U1079 ( .A1(KEYINPUT24), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1080 ( .A(n1312), .B(n1169), .ZN(n1338) );
XOR2_X1 U1081 ( .A(G143), .B(n1267), .Z(n1169) );
XOR2_X1 U1082 ( .A(G128), .B(G146), .Z(n1267) );
INV_X1 U1083 ( .A(n1171), .ZN(n1312) );
XOR2_X1 U1084 ( .A(G131), .B(n1339), .Z(n1171) );
XOR2_X1 U1085 ( .A(G137), .B(G134), .Z(n1339) );
XNOR2_X1 U1086 ( .A(G101), .B(KEYINPUT17), .ZN(n1336) );
endmodule


