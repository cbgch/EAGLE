//Key = 1101011000100000010101000000110011000100000010010101000000100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347;

XOR2_X1 U727 ( .A(n1021), .B(n1022), .Z(G9) );
NOR2_X1 U728 ( .A1(KEYINPUT24), .A2(n1023), .ZN(n1022) );
INV_X1 U729 ( .A(G107), .ZN(n1023) );
NOR3_X1 U730 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1021) );
INV_X1 U731 ( .A(n1027), .ZN(n1025) );
NOR2_X1 U732 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U733 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
XOR2_X1 U734 ( .A(n1034), .B(KEYINPUT8), .Z(n1033) );
NOR2_X1 U735 ( .A1(n1035), .A2(n1036), .ZN(n1032) );
NOR2_X1 U736 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U737 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
INV_X1 U738 ( .A(KEYINPUT54), .ZN(n1040) );
NOR4_X1 U739 ( .A1(n1024), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NOR2_X1 U740 ( .A1(n1044), .A2(n1043), .ZN(n1037) );
NOR2_X1 U741 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U742 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U743 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
AND2_X1 U744 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U745 ( .A1(n1053), .A2(n1041), .ZN(n1049) );
NOR4_X1 U746 ( .A1(KEYINPUT54), .A2(n1024), .A3(n1041), .A4(n1042), .ZN(n1045) );
NAND3_X1 U747 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1030) );
NAND3_X1 U748 ( .A1(n1052), .A2(n1057), .A3(n1058), .ZN(n1056) );
INV_X1 U749 ( .A(n1043), .ZN(n1058) );
NAND2_X1 U750 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND3_X1 U751 ( .A1(n1061), .A2(n1027), .A3(n1062), .ZN(n1060) );
NAND2_X1 U752 ( .A1(n1063), .A2(n1064), .ZN(n1059) );
NAND3_X1 U753 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
NAND3_X1 U754 ( .A1(n1068), .A2(n1061), .A3(n1069), .ZN(n1067) );
NAND3_X1 U755 ( .A1(n1070), .A2(n1062), .A3(n1071), .ZN(n1065) );
NOR3_X1 U756 ( .A1(n1072), .A2(G953), .A3(G952), .ZN(n1028) );
INV_X1 U757 ( .A(n1054), .ZN(n1072) );
NAND4_X1 U758 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1054) );
NOR4_X1 U759 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
XOR2_X1 U760 ( .A(KEYINPUT38), .B(n1081), .Z(n1080) );
XOR2_X1 U761 ( .A(n1070), .B(KEYINPUT29), .Z(n1077) );
NOR3_X1 U762 ( .A1(n1071), .A2(n1082), .A3(n1069), .ZN(n1075) );
XOR2_X1 U763 ( .A(n1083), .B(n1084), .Z(n1074) );
NOR2_X1 U764 ( .A1(n1085), .A2(KEYINPUT61), .ZN(n1084) );
XOR2_X1 U765 ( .A(G472), .B(n1086), .Z(n1073) );
NOR2_X1 U766 ( .A1(n1087), .A2(KEYINPUT48), .ZN(n1086) );
XOR2_X1 U767 ( .A(n1088), .B(n1089), .Z(G72) );
XOR2_X1 U768 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U769 ( .A1(G953), .A2(n1092), .ZN(n1091) );
NAND2_X1 U770 ( .A1(G900), .A2(G227), .ZN(n1092) );
NAND2_X1 U771 ( .A1(n1093), .A2(n1094), .ZN(n1090) );
NAND2_X1 U772 ( .A1(G953), .A2(n1095), .ZN(n1094) );
XOR2_X1 U773 ( .A(n1096), .B(n1097), .Z(n1093) );
XOR2_X1 U774 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U775 ( .A(n1100), .B(n1101), .Z(n1096) );
XNOR2_X1 U776 ( .A(G125), .B(KEYINPUT9), .ZN(n1101) );
NAND2_X1 U777 ( .A1(KEYINPUT1), .A2(n1102), .ZN(n1100) );
AND2_X1 U778 ( .A1(n1034), .A2(n1055), .ZN(n1088) );
XOR2_X1 U779 ( .A(n1103), .B(n1104), .Z(G69) );
NOR2_X1 U780 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U781 ( .A(n1107), .B(KEYINPUT10), .Z(n1106) );
NAND3_X1 U782 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
XOR2_X1 U783 ( .A(n1111), .B(KEYINPUT39), .Z(n1110) );
NAND2_X1 U784 ( .A1(G953), .A2(n1112), .ZN(n1109) );
NOR2_X1 U785 ( .A1(n1108), .A2(n1111), .ZN(n1105) );
NAND2_X1 U786 ( .A1(n1055), .A2(n1031), .ZN(n1111) );
XOR2_X1 U787 ( .A(n1113), .B(n1114), .Z(n1108) );
XNOR2_X1 U788 ( .A(n1115), .B(KEYINPUT26), .ZN(n1114) );
NAND2_X1 U789 ( .A1(KEYINPUT37), .A2(n1116), .ZN(n1115) );
XOR2_X1 U790 ( .A(n1117), .B(n1118), .Z(n1113) );
NAND2_X1 U791 ( .A1(G953), .A2(n1119), .ZN(n1103) );
NAND2_X1 U792 ( .A1(G898), .A2(G224), .ZN(n1119) );
NOR2_X1 U793 ( .A1(n1120), .A2(n1121), .ZN(G66) );
XNOR2_X1 U794 ( .A(n1122), .B(n1123), .ZN(n1121) );
NAND2_X1 U795 ( .A1(n1124), .A2(G217), .ZN(n1123) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1125), .ZN(G63) );
XNOR2_X1 U797 ( .A(n1126), .B(n1127), .ZN(n1125) );
NAND2_X1 U798 ( .A1(n1124), .A2(G478), .ZN(n1126) );
NOR2_X1 U799 ( .A1(n1120), .A2(n1128), .ZN(G60) );
NOR2_X1 U800 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
XOR2_X1 U801 ( .A(KEYINPUT55), .B(n1131), .Z(n1130) );
NOR2_X1 U802 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U803 ( .A(n1134), .B(KEYINPUT45), .Z(n1132) );
AND2_X1 U804 ( .A1(n1134), .A2(n1133), .ZN(n1129) );
NAND2_X1 U805 ( .A1(n1124), .A2(G475), .ZN(n1134) );
XOR2_X1 U806 ( .A(G104), .B(n1135), .Z(G6) );
NOR2_X1 U807 ( .A1(n1120), .A2(n1136), .ZN(G57) );
XOR2_X1 U808 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U809 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U810 ( .A1(KEYINPUT25), .A2(n1141), .ZN(n1140) );
XOR2_X1 U811 ( .A(n1142), .B(n1143), .Z(n1141) );
XNOR2_X1 U812 ( .A(G101), .B(KEYINPUT23), .ZN(n1143) );
NAND2_X1 U813 ( .A1(n1124), .A2(G472), .ZN(n1139) );
NOR2_X1 U814 ( .A1(n1120), .A2(n1144), .ZN(G54) );
XOR2_X1 U815 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U816 ( .A1(n1124), .A2(G469), .ZN(n1146) );
NAND2_X1 U817 ( .A1(n1147), .A2(KEYINPUT21), .ZN(n1145) );
XOR2_X1 U818 ( .A(n1148), .B(n1149), .Z(n1147) );
XOR2_X1 U819 ( .A(KEYINPUT43), .B(n1150), .Z(n1149) );
XOR2_X1 U820 ( .A(n1151), .B(n1152), .Z(n1148) );
NAND2_X1 U821 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
NAND2_X1 U822 ( .A1(n1098), .A2(n1155), .ZN(n1154) );
NAND2_X1 U823 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U824 ( .A1(KEYINPUT27), .A2(n1158), .ZN(n1157) );
NAND3_X1 U825 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1153) );
INV_X1 U826 ( .A(KEYINPUT27), .ZN(n1161) );
OR2_X1 U827 ( .A1(n1156), .A2(KEYINPUT12), .ZN(n1160) );
NAND2_X1 U828 ( .A1(n1156), .A2(n1162), .ZN(n1159) );
NAND2_X1 U829 ( .A1(n1163), .A2(n1158), .ZN(n1162) );
INV_X1 U830 ( .A(KEYINPUT12), .ZN(n1158) );
NOR3_X1 U831 ( .A1(n1120), .A2(n1164), .A3(n1165), .ZN(G51) );
NOR2_X1 U832 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U833 ( .A(n1168), .B(n1169), .Z(n1167) );
NOR2_X1 U834 ( .A1(KEYINPUT46), .A2(n1170), .ZN(n1168) );
NOR2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(n1164) );
XOR2_X1 U836 ( .A(n1173), .B(n1169), .Z(n1172) );
XNOR2_X1 U837 ( .A(n1174), .B(n1175), .ZN(n1169) );
NAND2_X1 U838 ( .A1(n1124), .A2(n1083), .ZN(n1174) );
AND2_X1 U839 ( .A1(G902), .A2(n1176), .ZN(n1124) );
OR2_X1 U840 ( .A1(n1031), .A2(n1034), .ZN(n1176) );
NAND4_X1 U841 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1034) );
NOR4_X1 U842 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
NOR2_X1 U843 ( .A1(n1185), .A2(n1186), .ZN(n1179) );
NAND4_X1 U844 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1031) );
AND3_X1 U845 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
OR3_X1 U846 ( .A1(n1048), .A2(n1053), .A3(n1026), .ZN(n1191) );
AND2_X1 U847 ( .A1(n1194), .A2(n1195), .ZN(n1053) );
NAND2_X1 U848 ( .A1(n1196), .A2(n1078), .ZN(n1195) );
NAND2_X1 U849 ( .A1(n1135), .A2(n1197), .ZN(n1189) );
NOR3_X1 U850 ( .A1(n1024), .A2(n1026), .A3(n1042), .ZN(n1135) );
NAND3_X1 U851 ( .A1(n1027), .A2(n1198), .A3(n1199), .ZN(n1188) );
XOR2_X1 U852 ( .A(KEYINPUT20), .B(n1200), .Z(n1198) );
NAND2_X1 U853 ( .A1(n1201), .A2(n1202), .ZN(n1187) );
NAND3_X1 U854 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1202) );
XOR2_X1 U855 ( .A(n1206), .B(KEYINPUT4), .Z(n1205) );
NAND4_X1 U856 ( .A1(n1207), .A2(n1052), .A3(n1027), .A4(n1051), .ZN(n1206) );
XOR2_X1 U857 ( .A(n1208), .B(KEYINPUT15), .Z(n1207) );
NAND4_X1 U858 ( .A1(n1208), .A2(n1024), .A3(n1051), .A4(n1209), .ZN(n1204) );
NOR2_X1 U859 ( .A1(n1042), .A2(n1197), .ZN(n1209) );
INV_X1 U860 ( .A(KEYINPUT63), .ZN(n1197) );
INV_X1 U861 ( .A(n1052), .ZN(n1024) );
XOR2_X1 U862 ( .A(n1210), .B(KEYINPUT40), .Z(n1203) );
NOR2_X1 U863 ( .A1(KEYINPUT46), .A2(n1211), .ZN(n1173) );
INV_X1 U864 ( .A(n1170), .ZN(n1211) );
XOR2_X1 U865 ( .A(n1212), .B(n1213), .Z(n1170) );
NOR2_X1 U866 ( .A1(G125), .A2(KEYINPUT22), .ZN(n1213) );
NOR2_X1 U867 ( .A1(n1055), .A2(G952), .ZN(n1120) );
XOR2_X1 U868 ( .A(G146), .B(n1186), .Z(G48) );
AND3_X1 U869 ( .A1(n1214), .A2(n1201), .A3(n1215), .ZN(n1186) );
XOR2_X1 U870 ( .A(n1216), .B(n1177), .Z(G45) );
NAND4_X1 U871 ( .A1(n1201), .A2(n1051), .A3(n1200), .A4(n1217), .ZN(n1177) );
AND3_X1 U872 ( .A1(n1079), .A2(n1218), .A3(n1219), .ZN(n1217) );
XOR2_X1 U873 ( .A(n1102), .B(n1178), .Z(G42) );
NAND4_X1 U874 ( .A1(n1220), .A2(n1062), .A3(n1214), .A4(n1219), .ZN(n1178) );
INV_X1 U875 ( .A(G140), .ZN(n1102) );
XOR2_X1 U876 ( .A(G137), .B(n1185), .Z(G39) );
AND3_X1 U877 ( .A1(n1062), .A2(n1063), .A3(n1215), .ZN(n1185) );
XNOR2_X1 U878 ( .A(G134), .B(n1221), .ZN(G36) );
NAND2_X1 U879 ( .A1(KEYINPUT58), .A2(n1184), .ZN(n1221) );
AND2_X1 U880 ( .A1(n1222), .A2(n1027), .ZN(n1184) );
XOR2_X1 U881 ( .A(n1183), .B(n1223), .Z(G33) );
NOR2_X1 U882 ( .A1(KEYINPUT13), .A2(n1224), .ZN(n1223) );
INV_X1 U883 ( .A(G131), .ZN(n1224) );
AND2_X1 U884 ( .A1(n1222), .A2(n1214), .ZN(n1183) );
AND4_X1 U885 ( .A1(n1062), .A2(n1200), .A3(n1051), .A4(n1219), .ZN(n1222) );
INV_X1 U886 ( .A(n1036), .ZN(n1062) );
NAND2_X1 U887 ( .A1(n1068), .A2(n1225), .ZN(n1036) );
XOR2_X1 U888 ( .A(G128), .B(n1182), .Z(G30) );
AND3_X1 U889 ( .A1(n1027), .A2(n1201), .A3(n1215), .ZN(n1182) );
AND4_X1 U890 ( .A1(n1051), .A2(n1226), .A3(n1219), .A4(n1078), .ZN(n1215) );
XOR2_X1 U891 ( .A(G101), .B(n1227), .Z(G3) );
NOR4_X1 U892 ( .A1(KEYINPUT57), .A2(n1026), .A3(n1048), .A4(n1194), .ZN(n1227) );
INV_X1 U893 ( .A(n1200), .ZN(n1194) );
INV_X1 U894 ( .A(n1063), .ZN(n1048) );
NAND3_X1 U895 ( .A1(n1051), .A2(n1208), .A3(n1201), .ZN(n1026) );
XOR2_X1 U896 ( .A(G125), .B(n1181), .Z(G27) );
AND4_X1 U897 ( .A1(n1214), .A2(n1228), .A3(n1229), .A4(n1196), .ZN(n1181) );
AND2_X1 U898 ( .A1(n1078), .A2(n1219), .ZN(n1229) );
NAND2_X1 U899 ( .A1(n1043), .A2(n1230), .ZN(n1219) );
NAND4_X1 U900 ( .A1(G953), .A2(G902), .A3(n1231), .A4(n1095), .ZN(n1230) );
INV_X1 U901 ( .A(G900), .ZN(n1095) );
XNOR2_X1 U902 ( .A(G122), .B(n1193), .ZN(G24) );
NAND4_X1 U903 ( .A1(n1199), .A2(n1052), .A3(n1079), .A4(n1218), .ZN(n1193) );
NOR2_X1 U904 ( .A1(n1078), .A2(n1226), .ZN(n1052) );
XOR2_X1 U905 ( .A(n1232), .B(n1192), .Z(G21) );
NAND4_X1 U906 ( .A1(n1063), .A2(n1199), .A3(n1226), .A4(n1078), .ZN(n1192) );
INV_X1 U907 ( .A(n1196), .ZN(n1226) );
NAND2_X1 U908 ( .A1(n1233), .A2(n1234), .ZN(G18) );
NAND2_X1 U909 ( .A1(G116), .A2(n1235), .ZN(n1234) );
XOR2_X1 U910 ( .A(n1236), .B(KEYINPUT56), .Z(n1233) );
OR2_X1 U911 ( .A1(n1235), .A2(G116), .ZN(n1236) );
NAND3_X1 U912 ( .A1(n1199), .A2(n1027), .A3(n1200), .ZN(n1235) );
NOR2_X1 U913 ( .A1(n1079), .A2(n1237), .ZN(n1027) );
AND2_X1 U914 ( .A1(n1228), .A2(n1208), .ZN(n1199) );
INV_X1 U915 ( .A(n1066), .ZN(n1228) );
NAND2_X1 U916 ( .A1(n1061), .A2(n1201), .ZN(n1066) );
XOR2_X1 U917 ( .A(G113), .B(n1238), .Z(G15) );
NOR2_X1 U918 ( .A1(n1239), .A2(n1210), .ZN(n1238) );
NAND4_X1 U919 ( .A1(n1214), .A2(n1200), .A3(n1061), .A4(n1208), .ZN(n1210) );
INV_X1 U920 ( .A(n1041), .ZN(n1061) );
NAND2_X1 U921 ( .A1(n1070), .A2(n1240), .ZN(n1041) );
NOR2_X1 U922 ( .A1(n1078), .A2(n1196), .ZN(n1200) );
INV_X1 U923 ( .A(n1042), .ZN(n1214) );
NAND2_X1 U924 ( .A1(n1241), .A2(n1079), .ZN(n1042) );
XOR2_X1 U925 ( .A(KEYINPUT62), .B(n1237), .Z(n1241) );
XOR2_X1 U926 ( .A(n1242), .B(n1243), .Z(G12) );
NAND2_X1 U927 ( .A1(KEYINPUT49), .A2(G110), .ZN(n1243) );
NAND4_X1 U928 ( .A1(n1244), .A2(n1220), .A3(n1063), .A4(n1208), .ZN(n1242) );
NAND2_X1 U929 ( .A1(n1043), .A2(n1245), .ZN(n1208) );
NAND4_X1 U930 ( .A1(G953), .A2(G902), .A3(n1231), .A4(n1112), .ZN(n1245) );
INV_X1 U931 ( .A(G898), .ZN(n1112) );
NAND3_X1 U932 ( .A1(n1231), .A2(n1055), .A3(G952), .ZN(n1043) );
NAND2_X1 U933 ( .A1(G237), .A2(G234), .ZN(n1231) );
NOR2_X1 U934 ( .A1(n1218), .A2(n1079), .ZN(n1063) );
XNOR2_X1 U935 ( .A(n1246), .B(G475), .ZN(n1079) );
NAND2_X1 U936 ( .A1(n1133), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U937 ( .A(n1248), .B(n1249), .ZN(n1133) );
XOR2_X1 U938 ( .A(n1250), .B(n1251), .Z(n1248) );
XOR2_X1 U939 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U940 ( .A(G122), .B(G113), .Z(n1253) );
XOR2_X1 U941 ( .A(KEYINPUT50), .B(KEYINPUT35), .Z(n1252) );
XOR2_X1 U942 ( .A(n1254), .B(n1255), .Z(n1250) );
XNOR2_X1 U943 ( .A(n1256), .B(n1257), .ZN(n1255) );
XNOR2_X1 U944 ( .A(G104), .B(n1258), .ZN(n1254) );
NOR2_X1 U945 ( .A1(KEYINPUT30), .A2(n1259), .ZN(n1258) );
XOR2_X1 U946 ( .A(G143), .B(n1260), .Z(n1259) );
AND3_X1 U947 ( .A1(G214), .A2(n1055), .A3(n1261), .ZN(n1260) );
INV_X1 U948 ( .A(n1237), .ZN(n1218) );
NOR2_X1 U949 ( .A1(n1081), .A2(n1082), .ZN(n1237) );
NOR3_X1 U950 ( .A1(G478), .A2(G902), .A3(n1127), .ZN(n1082) );
AND2_X1 U951 ( .A1(G478), .A2(n1262), .ZN(n1081) );
OR2_X1 U952 ( .A1(n1127), .A2(G902), .ZN(n1262) );
XNOR2_X1 U953 ( .A(n1263), .B(n1264), .ZN(n1127) );
XOR2_X1 U954 ( .A(G107), .B(n1265), .Z(n1264) );
XOR2_X1 U955 ( .A(G122), .B(G116), .Z(n1265) );
XOR2_X1 U956 ( .A(n1266), .B(n1267), .Z(n1263) );
NOR3_X1 U957 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1267) );
INV_X1 U958 ( .A(G234), .ZN(n1270) );
XOR2_X1 U959 ( .A(KEYINPUT34), .B(G953), .Z(n1268) );
NAND2_X1 U960 ( .A1(KEYINPUT17), .A2(n1271), .ZN(n1266) );
XNOR2_X1 U961 ( .A(G134), .B(n1272), .ZN(n1271) );
NAND2_X1 U962 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NAND2_X1 U963 ( .A1(G143), .A2(n1275), .ZN(n1274) );
XOR2_X1 U964 ( .A(n1276), .B(KEYINPUT11), .Z(n1273) );
NAND2_X1 U965 ( .A1(G128), .A2(n1216), .ZN(n1276) );
AND3_X1 U966 ( .A1(n1196), .A2(n1078), .A3(n1051), .ZN(n1220) );
NOR2_X1 U967 ( .A1(n1070), .A2(n1071), .ZN(n1051) );
INV_X1 U968 ( .A(n1240), .ZN(n1071) );
NAND2_X1 U969 ( .A1(G221), .A2(n1277), .ZN(n1240) );
NAND2_X1 U970 ( .A1(G234), .A2(n1247), .ZN(n1277) );
XOR2_X1 U971 ( .A(n1278), .B(G469), .Z(n1070) );
NAND2_X1 U972 ( .A1(n1279), .A2(n1247), .ZN(n1278) );
XOR2_X1 U973 ( .A(n1280), .B(n1281), .Z(n1279) );
XNOR2_X1 U974 ( .A(n1156), .B(n1152), .ZN(n1281) );
XOR2_X1 U975 ( .A(G110), .B(G140), .Z(n1152) );
XNOR2_X1 U976 ( .A(n1099), .B(n1282), .ZN(n1156) );
XNOR2_X1 U977 ( .A(n1216), .B(n1283), .ZN(n1099) );
XOR2_X1 U978 ( .A(n1150), .B(n1098), .Z(n1280) );
AND2_X1 U979 ( .A1(G227), .A2(n1055), .ZN(n1150) );
NAND3_X1 U980 ( .A1(n1284), .A2(n1285), .A3(n1286), .ZN(n1078) );
NAND2_X1 U981 ( .A1(n1122), .A2(n1287), .ZN(n1286) );
OR3_X1 U982 ( .A1(n1287), .A2(n1122), .A3(G902), .ZN(n1285) );
AND2_X1 U983 ( .A1(n1288), .A2(n1289), .ZN(n1122) );
NAND2_X1 U984 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U985 ( .A(KEYINPUT3), .B(n1292), .Z(n1288) );
NOR2_X1 U986 ( .A1(n1290), .A2(n1291), .ZN(n1292) );
XOR2_X1 U987 ( .A(n1293), .B(G137), .Z(n1291) );
NAND3_X1 U988 ( .A1(G221), .A2(n1055), .A3(G234), .ZN(n1293) );
AND2_X1 U989 ( .A1(n1294), .A2(n1295), .ZN(n1290) );
NAND2_X1 U990 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
NAND2_X1 U991 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
OR2_X1 U992 ( .A1(n1300), .A2(KEYINPUT18), .ZN(n1298) );
XOR2_X1 U993 ( .A(n1301), .B(n1302), .Z(n1296) );
INV_X1 U994 ( .A(n1249), .ZN(n1301) );
NAND2_X1 U995 ( .A1(n1300), .A2(n1303), .ZN(n1294) );
NAND2_X1 U996 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
INV_X1 U997 ( .A(KEYINPUT18), .ZN(n1305) );
NAND2_X1 U998 ( .A1(n1306), .A2(n1299), .ZN(n1304) );
INV_X1 U999 ( .A(KEYINPUT42), .ZN(n1299) );
XOR2_X1 U1000 ( .A(n1302), .B(n1249), .Z(n1306) );
XOR2_X1 U1001 ( .A(G146), .B(G125), .Z(n1249) );
XNOR2_X1 U1002 ( .A(KEYINPUT2), .B(n1307), .ZN(n1302) );
NOR2_X1 U1003 ( .A1(KEYINPUT31), .A2(n1257), .ZN(n1307) );
XNOR2_X1 U1004 ( .A(G140), .B(KEYINPUT33), .ZN(n1257) );
XOR2_X1 U1005 ( .A(G110), .B(n1308), .Z(n1300) );
XOR2_X1 U1006 ( .A(G128), .B(G119), .Z(n1308) );
NOR2_X1 U1007 ( .A1(n1269), .A2(G234), .ZN(n1287) );
INV_X1 U1008 ( .A(G217), .ZN(n1269) );
NAND2_X1 U1009 ( .A1(G902), .A2(G217), .ZN(n1284) );
XNOR2_X1 U1010 ( .A(n1087), .B(G472), .ZN(n1196) );
AND3_X1 U1011 ( .A1(n1309), .A2(n1310), .A3(n1247), .ZN(n1087) );
NAND3_X1 U1012 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1310) );
INV_X1 U1013 ( .A(KEYINPUT19), .ZN(n1313) );
XOR2_X1 U1014 ( .A(n1314), .B(n1315), .Z(n1311) );
NAND2_X1 U1015 ( .A1(n1316), .A2(KEYINPUT19), .ZN(n1309) );
XOR2_X1 U1016 ( .A(n1317), .B(n1315), .Z(n1316) );
XOR2_X1 U1017 ( .A(n1142), .B(n1318), .Z(n1315) );
NOR2_X1 U1018 ( .A1(G101), .A2(KEYINPUT14), .ZN(n1318) );
NAND3_X1 U1019 ( .A1(n1261), .A2(n1055), .A3(G210), .ZN(n1142) );
INV_X1 U1020 ( .A(G237), .ZN(n1261) );
NAND2_X1 U1021 ( .A1(n1312), .A2(n1314), .ZN(n1317) );
INV_X1 U1022 ( .A(KEYINPUT7), .ZN(n1314) );
XOR2_X1 U1023 ( .A(n1137), .B(KEYINPUT6), .Z(n1312) );
XOR2_X1 U1024 ( .A(n1319), .B(n1320), .Z(n1137) );
XNOR2_X1 U1025 ( .A(G113), .B(n1321), .ZN(n1320) );
NAND2_X1 U1026 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
NAND2_X1 U1027 ( .A1(G116), .A2(n1232), .ZN(n1323) );
XOR2_X1 U1028 ( .A(n1324), .B(KEYINPUT36), .Z(n1322) );
OR2_X1 U1029 ( .A1(n1232), .A2(G116), .ZN(n1324) );
INV_X1 U1030 ( .A(G119), .ZN(n1232) );
XOR2_X1 U1031 ( .A(n1212), .B(n1098), .Z(n1319) );
INV_X1 U1032 ( .A(n1163), .ZN(n1098) );
XOR2_X1 U1033 ( .A(n1325), .B(n1256), .Z(n1163) );
XOR2_X1 U1034 ( .A(G131), .B(KEYINPUT41), .Z(n1256) );
XNOR2_X1 U1035 ( .A(G134), .B(G137), .ZN(n1325) );
XOR2_X1 U1036 ( .A(n1239), .B(KEYINPUT51), .Z(n1244) );
INV_X1 U1037 ( .A(n1201), .ZN(n1239) );
NOR2_X1 U1038 ( .A1(n1068), .A2(n1069), .ZN(n1201) );
INV_X1 U1039 ( .A(n1225), .ZN(n1069) );
NAND2_X1 U1040 ( .A1(G214), .A2(n1326), .ZN(n1225) );
XOR2_X1 U1041 ( .A(KEYINPUT5), .B(n1327), .Z(n1326) );
XNOR2_X1 U1042 ( .A(n1085), .B(n1083), .ZN(n1068) );
NOR2_X1 U1043 ( .A1(n1328), .A2(n1327), .ZN(n1083) );
NOR2_X1 U1044 ( .A1(G902), .A2(G237), .ZN(n1327) );
INV_X1 U1045 ( .A(G210), .ZN(n1328) );
AND3_X1 U1046 ( .A1(n1329), .A2(n1247), .A3(n1330), .ZN(n1085) );
XOR2_X1 U1047 ( .A(n1331), .B(KEYINPUT16), .Z(n1330) );
OR2_X1 U1048 ( .A1(n1332), .A2(n1175), .ZN(n1331) );
INV_X1 U1049 ( .A(G902), .ZN(n1247) );
NAND2_X1 U1050 ( .A1(n1175), .A2(n1332), .ZN(n1329) );
XNOR2_X1 U1051 ( .A(n1212), .B(n1333), .ZN(n1332) );
XOR2_X1 U1052 ( .A(G125), .B(n1171), .Z(n1333) );
INV_X1 U1053 ( .A(n1166), .ZN(n1171) );
NAND2_X1 U1054 ( .A1(G224), .A2(n1055), .ZN(n1166) );
INV_X1 U1055 ( .A(G953), .ZN(n1055) );
XOR2_X1 U1056 ( .A(n1334), .B(n1283), .Z(n1212) );
XNOR2_X1 U1057 ( .A(G146), .B(n1275), .ZN(n1283) );
INV_X1 U1058 ( .A(G128), .ZN(n1275) );
NAND2_X1 U1059 ( .A1(n1335), .A2(KEYINPUT28), .ZN(n1334) );
XOR2_X1 U1060 ( .A(n1216), .B(KEYINPUT59), .Z(n1335) );
INV_X1 U1061 ( .A(G143), .ZN(n1216) );
AND2_X1 U1062 ( .A1(n1336), .A2(n1337), .ZN(n1175) );
NAND2_X1 U1063 ( .A1(n1338), .A2(n1118), .ZN(n1337) );
NAND2_X1 U1064 ( .A1(n1282), .A2(n1339), .ZN(n1336) );
XNOR2_X1 U1065 ( .A(n1340), .B(n1338), .ZN(n1339) );
XNOR2_X1 U1066 ( .A(n1341), .B(n1116), .ZN(n1338) );
XOR2_X1 U1067 ( .A(n1342), .B(n1343), .Z(n1116) );
XOR2_X1 U1068 ( .A(G119), .B(G113), .Z(n1343) );
NAND2_X1 U1069 ( .A1(KEYINPUT0), .A2(G116), .ZN(n1342) );
NAND2_X1 U1070 ( .A1(KEYINPUT32), .A2(n1117), .ZN(n1341) );
XNOR2_X1 U1071 ( .A(n1344), .B(n1345), .ZN(n1117) );
XOR2_X1 U1072 ( .A(G122), .B(G110), .Z(n1345) );
XNOR2_X1 U1073 ( .A(KEYINPUT60), .B(KEYINPUT44), .ZN(n1344) );
XNOR2_X1 U1074 ( .A(KEYINPUT53), .B(KEYINPUT47), .ZN(n1340) );
INV_X1 U1075 ( .A(n1118), .ZN(n1282) );
XOR2_X1 U1076 ( .A(n1346), .B(n1347), .Z(n1118) );
XOR2_X1 U1077 ( .A(KEYINPUT52), .B(G107), .Z(n1347) );
XNOR2_X1 U1078 ( .A(G104), .B(G101), .ZN(n1346) );
endmodule


