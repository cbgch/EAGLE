//Key = 0001111000000011111010000011111010010000000001100111110010101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365;

XNOR2_X1 U753 ( .A(G107), .B(n1042), .ZN(G9) );
NOR2_X1 U754 ( .A1(n1043), .A2(n1044), .ZN(G75) );
NOR3_X1 U755 ( .A1(n1045), .A2(G953), .A3(n1046), .ZN(n1044) );
XOR2_X1 U756 ( .A(n1047), .B(KEYINPUT19), .Z(n1045) );
NAND3_X1 U757 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NAND2_X1 U759 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND3_X1 U760 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
NAND2_X1 U765 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U767 ( .A1(n1064), .A2(n1070), .A3(n1060), .ZN(n1053) );
NAND2_X1 U768 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U769 ( .A1(n1057), .A2(n1073), .ZN(n1072) );
OR2_X1 U770 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND2_X1 U771 ( .A1(n1055), .A2(n1076), .ZN(n1071) );
NAND2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U774 ( .A(n1081), .ZN(n1051) );
NOR3_X1 U775 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1043) );
AND4_X1 U776 ( .A1(n1082), .A2(n1055), .A3(n1060), .A4(n1083), .ZN(n1046) );
NOR3_X1 U777 ( .A1(n1084), .A2(n1079), .A3(n1085), .ZN(n1083) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U780 ( .A1(KEYINPUT21), .A2(n1090), .ZN(n1088) );
NOR2_X1 U781 ( .A1(n1091), .A2(KEYINPUT39), .ZN(n1090) );
NOR2_X1 U782 ( .A1(n1092), .A2(n1093), .ZN(n1086) );
NOR2_X1 U783 ( .A1(n1094), .A2(KEYINPUT39), .ZN(n1092) );
NOR2_X1 U784 ( .A1(KEYINPUT21), .A2(n1095), .ZN(n1094) );
XOR2_X1 U785 ( .A(n1096), .B(KEYINPUT33), .Z(n1084) );
NAND3_X1 U786 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NAND2_X1 U787 ( .A1(KEYINPUT7), .A2(n1100), .ZN(n1098) );
OR2_X1 U788 ( .A1(n1101), .A2(KEYINPUT7), .ZN(n1097) );
XOR2_X1 U789 ( .A(n1102), .B(n1103), .Z(G72) );
NOR2_X1 U790 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NAND2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1102) );
OR3_X1 U793 ( .A1(n1048), .A2(G953), .A3(n1110), .ZN(n1109) );
NAND3_X1 U794 ( .A1(n1111), .A2(n1112), .A3(n1110), .ZN(n1108) );
XNOR2_X1 U795 ( .A(n1113), .B(n1114), .ZN(n1110) );
XOR2_X1 U796 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND3_X1 U797 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1115) );
NAND2_X1 U798 ( .A1(G140), .A2(n1120), .ZN(n1119) );
OR3_X1 U799 ( .A1(n1120), .A2(G140), .A3(n1121), .ZN(n1118) );
NAND2_X1 U800 ( .A1(KEYINPUT60), .A2(n1122), .ZN(n1120) );
NAND2_X1 U801 ( .A1(G125), .A2(n1121), .ZN(n1117) );
INV_X1 U802 ( .A(KEYINPUT14), .ZN(n1121) );
XNOR2_X1 U803 ( .A(G131), .B(n1123), .ZN(n1113) );
NOR2_X1 U804 ( .A1(KEYINPUT1), .A2(n1124), .ZN(n1123) );
NAND2_X1 U805 ( .A1(G953), .A2(n1107), .ZN(n1112) );
XOR2_X1 U806 ( .A(KEYINPUT36), .B(n1048), .Z(n1111) );
XOR2_X1 U807 ( .A(n1125), .B(n1126), .Z(G69) );
NOR2_X1 U808 ( .A1(n1050), .A2(G953), .ZN(n1126) );
NAND2_X1 U809 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
NAND2_X1 U810 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
OR2_X1 U811 ( .A1(n1105), .A2(G224), .ZN(n1130) );
NAND2_X1 U812 ( .A1(G953), .A2(n1131), .ZN(n1127) );
NAND2_X1 U813 ( .A1(G898), .A2(n1132), .ZN(n1131) );
OR2_X1 U814 ( .A1(n1129), .A2(G224), .ZN(n1132) );
XNOR2_X1 U815 ( .A(n1133), .B(n1134), .ZN(n1129) );
XNOR2_X1 U816 ( .A(n1135), .B(KEYINPUT30), .ZN(n1134) );
NAND2_X1 U817 ( .A1(KEYINPUT26), .A2(n1136), .ZN(n1135) );
XNOR2_X1 U818 ( .A(n1137), .B(G110), .ZN(n1136) );
XOR2_X1 U819 ( .A(n1138), .B(n1139), .Z(n1133) );
NAND2_X1 U820 ( .A1(KEYINPUT3), .A2(n1140), .ZN(n1138) );
NOR2_X1 U821 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XOR2_X1 U822 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U823 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U824 ( .A1(KEYINPUT29), .A2(n1147), .ZN(n1143) );
NOR2_X1 U825 ( .A1(n1141), .A2(n1148), .ZN(G63) );
XNOR2_X1 U826 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U827 ( .A1(n1100), .A2(n1146), .ZN(n1150) );
NOR2_X1 U828 ( .A1(n1141), .A2(n1151), .ZN(G60) );
XNOR2_X1 U829 ( .A(n1152), .B(n1153), .ZN(n1151) );
AND2_X1 U830 ( .A1(G475), .A2(n1154), .ZN(n1153) );
XNOR2_X1 U831 ( .A(G104), .B(n1155), .ZN(G6) );
NOR2_X1 U832 ( .A1(n1141), .A2(n1156), .ZN(G57) );
XOR2_X1 U833 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U834 ( .A(n1159), .B(n1160), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1161), .B(n1162), .Z(n1157) );
XOR2_X1 U836 ( .A(KEYINPUT49), .B(n1163), .Z(n1162) );
AND2_X1 U837 ( .A1(G472), .A2(n1154), .ZN(n1163) );
NAND2_X1 U838 ( .A1(KEYINPUT27), .A2(n1164), .ZN(n1161) );
NOR2_X1 U839 ( .A1(n1141), .A2(n1165), .ZN(G54) );
XOR2_X1 U840 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(n1167) );
XNOR2_X1 U842 ( .A(n1170), .B(n1116), .ZN(n1169) );
XOR2_X1 U843 ( .A(n1171), .B(n1172), .Z(n1166) );
XOR2_X1 U844 ( .A(KEYINPUT52), .B(n1173), .Z(n1172) );
AND2_X1 U845 ( .A1(G469), .A2(n1154), .ZN(n1173) );
NAND2_X1 U846 ( .A1(n1174), .A2(KEYINPUT63), .ZN(n1171) );
XOR2_X1 U847 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR3_X1 U848 ( .A1(n1106), .A2(KEYINPUT57), .A3(G953), .ZN(n1176) );
XNOR2_X1 U849 ( .A(G110), .B(G140), .ZN(n1175) );
NOR2_X1 U850 ( .A1(n1141), .A2(n1177), .ZN(G51) );
XNOR2_X1 U851 ( .A(n1178), .B(n1179), .ZN(n1177) );
XNOR2_X1 U852 ( .A(n1180), .B(n1181), .ZN(n1179) );
NAND3_X1 U853 ( .A1(n1154), .A2(n1089), .A3(KEYINPUT18), .ZN(n1181) );
INV_X1 U854 ( .A(n1095), .ZN(n1089) );
INV_X1 U855 ( .A(n1146), .ZN(n1154) );
NAND2_X1 U856 ( .A1(G902), .A2(n1182), .ZN(n1146) );
NAND2_X1 U857 ( .A1(n1050), .A2(n1048), .ZN(n1182) );
AND4_X1 U858 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1048) );
AND4_X1 U859 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1186) );
AND2_X1 U860 ( .A1(n1191), .A2(n1192), .ZN(n1185) );
NAND2_X1 U861 ( .A1(n1193), .A2(n1194), .ZN(n1183) );
XNOR2_X1 U862 ( .A(KEYINPUT61), .B(n1063), .ZN(n1194) );
AND4_X1 U863 ( .A1(n1042), .A2(n1155), .A3(n1195), .A4(n1196), .ZN(n1050) );
AND4_X1 U864 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1196) );
NOR3_X1 U865 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1195) );
NOR3_X1 U866 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
AND2_X1 U867 ( .A1(n1204), .A2(n1207), .ZN(n1202) );
INV_X1 U868 ( .A(KEYINPUT48), .ZN(n1204) );
AND3_X1 U869 ( .A1(n1208), .A2(n1209), .A3(n1074), .ZN(n1201) );
NAND3_X1 U870 ( .A1(n1210), .A2(n1055), .A3(n1211), .ZN(n1155) );
NAND3_X1 U871 ( .A1(n1212), .A2(n1055), .A3(n1210), .ZN(n1042) );
NAND2_X1 U872 ( .A1(n1213), .A2(KEYINPUT15), .ZN(n1180) );
XNOR2_X1 U873 ( .A(G125), .B(n1214), .ZN(n1213) );
NOR2_X1 U874 ( .A1(n1105), .A2(G952), .ZN(n1141) );
XOR2_X1 U875 ( .A(G146), .B(n1215), .Z(G48) );
NOR2_X1 U876 ( .A1(KEYINPUT11), .A2(n1192), .ZN(n1215) );
NAND3_X1 U877 ( .A1(n1211), .A2(n1205), .A3(n1216), .ZN(n1192) );
XNOR2_X1 U878 ( .A(G143), .B(n1191), .ZN(G45) );
NAND3_X1 U879 ( .A1(n1217), .A2(n1074), .A3(n1218), .ZN(n1191) );
NOR3_X1 U880 ( .A1(n1077), .A2(n1219), .A3(n1082), .ZN(n1218) );
XNOR2_X1 U881 ( .A(G140), .B(n1190), .ZN(G42) );
NAND4_X1 U882 ( .A1(n1057), .A2(n1217), .A3(n1211), .A4(n1075), .ZN(n1190) );
NAND2_X1 U883 ( .A1(n1220), .A2(n1221), .ZN(G39) );
NAND2_X1 U884 ( .A1(n1222), .A2(G137), .ZN(n1221) );
XOR2_X1 U885 ( .A(KEYINPUT46), .B(n1223), .Z(n1220) );
NOR2_X1 U886 ( .A1(G137), .A2(n1222), .ZN(n1223) );
AND2_X1 U887 ( .A1(n1224), .A2(n1225), .ZN(n1222) );
OR2_X1 U888 ( .A1(n1184), .A2(KEYINPUT13), .ZN(n1225) );
NAND3_X1 U889 ( .A1(n1216), .A2(n1064), .A3(n1057), .ZN(n1184) );
NAND4_X1 U890 ( .A1(n1064), .A2(n1226), .A3(n1216), .A4(KEYINPUT13), .ZN(n1224) );
INV_X1 U891 ( .A(n1057), .ZN(n1226) );
XOR2_X1 U892 ( .A(G134), .B(n1227), .Z(G36) );
NOR2_X1 U893 ( .A1(n1063), .A2(n1228), .ZN(n1227) );
XOR2_X1 U894 ( .A(n1229), .B(n1230), .Z(G33) );
XOR2_X1 U895 ( .A(KEYINPUT9), .B(G131), .Z(n1230) );
NOR2_X1 U896 ( .A1(KEYINPUT47), .A2(n1189), .ZN(n1229) );
NAND2_X1 U897 ( .A1(n1193), .A2(n1211), .ZN(n1189) );
INV_X1 U898 ( .A(n1062), .ZN(n1211) );
INV_X1 U899 ( .A(n1228), .ZN(n1193) );
NAND3_X1 U900 ( .A1(n1217), .A2(n1074), .A3(n1057), .ZN(n1228) );
NOR2_X1 U901 ( .A1(n1231), .A2(n1079), .ZN(n1057) );
XNOR2_X1 U902 ( .A(G128), .B(n1188), .ZN(G30) );
NAND3_X1 U903 ( .A1(n1212), .A2(n1205), .A3(n1216), .ZN(n1188) );
AND3_X1 U904 ( .A1(n1232), .A2(n1233), .A3(n1217), .ZN(n1216) );
AND2_X1 U905 ( .A1(n1234), .A2(n1235), .ZN(n1217) );
XNOR2_X1 U906 ( .A(G101), .B(n1200), .ZN(G3) );
NAND3_X1 U907 ( .A1(n1210), .A2(n1064), .A3(n1074), .ZN(n1200) );
XOR2_X1 U908 ( .A(n1187), .B(n1236), .Z(G27) );
NAND2_X1 U909 ( .A1(KEYINPUT62), .A2(G125), .ZN(n1236) );
NAND3_X1 U910 ( .A1(n1075), .A2(n1235), .A3(n1208), .ZN(n1187) );
NOR3_X1 U911 ( .A1(n1237), .A2(n1077), .A3(n1062), .ZN(n1208) );
NAND2_X1 U912 ( .A1(n1081), .A2(n1238), .ZN(n1235) );
NAND4_X1 U913 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1107), .ZN(n1238) );
INV_X1 U914 ( .A(G900), .ZN(n1107) );
XNOR2_X1 U915 ( .A(G122), .B(n1199), .ZN(G24) );
NAND3_X1 U916 ( .A1(n1060), .A2(n1055), .A3(n1240), .ZN(n1199) );
NOR3_X1 U917 ( .A1(n1241), .A2(n1219), .A3(n1082), .ZN(n1240) );
INV_X1 U918 ( .A(n1242), .ZN(n1082) );
NOR2_X1 U919 ( .A1(n1233), .A2(n1232), .ZN(n1055) );
XNOR2_X1 U920 ( .A(n1243), .B(n1207), .ZN(G21) );
NOR2_X1 U921 ( .A1(n1206), .A2(n1077), .ZN(n1207) );
NAND3_X1 U922 ( .A1(n1060), .A2(n1064), .A3(n1244), .ZN(n1206) );
NOR3_X1 U923 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
INV_X1 U924 ( .A(n1237), .ZN(n1060) );
XNOR2_X1 U925 ( .A(G116), .B(n1198), .ZN(G18) );
OR4_X1 U926 ( .A1(n1248), .A2(n1237), .A3(n1063), .A4(n1241), .ZN(n1198) );
INV_X1 U927 ( .A(n1212), .ZN(n1063) );
INV_X1 U928 ( .A(n1074), .ZN(n1248) );
XNOR2_X1 U929 ( .A(n1249), .B(n1250), .ZN(G15) );
NOR3_X1 U930 ( .A1(n1251), .A2(KEYINPUT24), .A3(n1077), .ZN(n1250) );
INV_X1 U931 ( .A(n1205), .ZN(n1077) );
XOR2_X1 U932 ( .A(KEYINPUT45), .B(n1252), .Z(n1251) );
NOR4_X1 U933 ( .A1(n1246), .A2(n1253), .A3(n1237), .A4(n1062), .ZN(n1252) );
NAND2_X1 U934 ( .A1(n1254), .A2(n1242), .ZN(n1062) );
XNOR2_X1 U935 ( .A(KEYINPUT34), .B(n1255), .ZN(n1254) );
NAND2_X1 U936 ( .A1(n1069), .A2(n1256), .ZN(n1237) );
XNOR2_X1 U937 ( .A(n1074), .B(KEYINPUT44), .ZN(n1253) );
NOR2_X1 U938 ( .A1(n1232), .A2(n1247), .ZN(n1074) );
INV_X1 U939 ( .A(n1233), .ZN(n1247) );
INV_X1 U940 ( .A(n1209), .ZN(n1246) );
XNOR2_X1 U941 ( .A(n1197), .B(n1257), .ZN(G12) );
NOR2_X1 U942 ( .A1(KEYINPUT8), .A2(n1258), .ZN(n1257) );
INV_X1 U943 ( .A(G110), .ZN(n1258) );
NAND3_X1 U944 ( .A1(n1210), .A2(n1064), .A3(n1075), .ZN(n1197) );
NOR2_X1 U945 ( .A1(n1233), .A2(n1245), .ZN(n1075) );
INV_X1 U946 ( .A(n1232), .ZN(n1245) );
XOR2_X1 U947 ( .A(n1259), .B(n1145), .Z(n1232) );
NAND2_X1 U948 ( .A1(G217), .A2(n1260), .ZN(n1145) );
NAND2_X1 U949 ( .A1(n1147), .A2(n1261), .ZN(n1259) );
XOR2_X1 U950 ( .A(n1262), .B(n1263), .Z(n1147) );
XNOR2_X1 U951 ( .A(n1264), .B(n1265), .ZN(n1263) );
NOR2_X1 U952 ( .A1(KEYINPUT10), .A2(n1266), .ZN(n1265) );
NAND2_X1 U953 ( .A1(KEYINPUT17), .A2(G110), .ZN(n1264) );
XOR2_X1 U954 ( .A(n1267), .B(n1268), .Z(n1262) );
NOR2_X1 U955 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
INV_X1 U956 ( .A(G221), .ZN(n1269) );
XOR2_X1 U957 ( .A(n1271), .B(n1272), .Z(n1267) );
XNOR2_X1 U958 ( .A(G128), .B(n1273), .ZN(n1272) );
XNOR2_X1 U959 ( .A(KEYINPUT59), .B(KEYINPUT4), .ZN(n1273) );
XOR2_X1 U960 ( .A(n1274), .B(n1275), .Z(n1271) );
XNOR2_X1 U961 ( .A(G119), .B(n1276), .ZN(n1274) );
XNOR2_X1 U962 ( .A(n1277), .B(G472), .ZN(n1233) );
NAND2_X1 U963 ( .A1(n1278), .A2(n1261), .ZN(n1277) );
XNOR2_X1 U964 ( .A(n1164), .B(n1279), .ZN(n1278) );
XOR2_X1 U965 ( .A(n1280), .B(n1160), .Z(n1279) );
XNOR2_X1 U966 ( .A(n1281), .B(n1282), .ZN(n1160) );
XNOR2_X1 U967 ( .A(G101), .B(n1283), .ZN(n1282) );
NAND2_X1 U968 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U969 ( .A1(n1286), .A2(n1249), .ZN(n1285) );
XOR2_X1 U970 ( .A(n1287), .B(KEYINPUT42), .Z(n1284) );
OR2_X1 U971 ( .A1(n1286), .A2(n1249), .ZN(n1287) );
XOR2_X1 U972 ( .A(n1288), .B(KEYINPUT32), .Z(n1286) );
NAND2_X1 U973 ( .A1(n1289), .A2(G210), .ZN(n1281) );
NOR2_X1 U974 ( .A1(n1159), .A2(n1290), .ZN(n1280) );
XOR2_X1 U975 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n1290) );
INV_X1 U976 ( .A(n1170), .ZN(n1164) );
NAND2_X1 U977 ( .A1(n1291), .A2(n1292), .ZN(n1064) );
OR3_X1 U978 ( .A1(n1255), .A2(n1242), .A3(KEYINPUT34), .ZN(n1292) );
NAND2_X1 U979 ( .A1(KEYINPUT34), .A2(n1212), .ZN(n1291) );
NOR2_X1 U980 ( .A1(n1242), .A2(n1219), .ZN(n1212) );
INV_X1 U981 ( .A(n1255), .ZN(n1219) );
NAND2_X1 U982 ( .A1(n1099), .A2(n1101), .ZN(n1255) );
NAND2_X1 U983 ( .A1(G478), .A2(n1293), .ZN(n1101) );
NAND2_X1 U984 ( .A1(n1149), .A2(n1261), .ZN(n1293) );
NAND3_X1 U985 ( .A1(n1100), .A2(n1261), .A3(n1149), .ZN(n1099) );
XNOR2_X1 U986 ( .A(n1294), .B(n1295), .ZN(n1149) );
NOR2_X1 U987 ( .A1(n1270), .A2(n1296), .ZN(n1295) );
INV_X1 U988 ( .A(G217), .ZN(n1296) );
NAND2_X1 U989 ( .A1(G234), .A2(n1105), .ZN(n1270) );
NAND2_X1 U990 ( .A1(KEYINPUT28), .A2(n1297), .ZN(n1294) );
XOR2_X1 U991 ( .A(n1298), .B(n1299), .Z(n1297) );
XOR2_X1 U992 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U993 ( .A(n1302), .B(n1303), .Z(n1298) );
NOR2_X1 U994 ( .A1(KEYINPUT0), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U995 ( .A(G116), .B(G122), .ZN(n1304) );
XNOR2_X1 U996 ( .A(G107), .B(KEYINPUT41), .ZN(n1302) );
INV_X1 U997 ( .A(G478), .ZN(n1100) );
XNOR2_X1 U998 ( .A(n1305), .B(G475), .ZN(n1242) );
NAND2_X1 U999 ( .A1(n1261), .A2(n1152), .ZN(n1305) );
NAND2_X1 U1000 ( .A1(n1306), .A2(n1307), .ZN(n1152) );
NAND2_X1 U1001 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XOR2_X1 U1002 ( .A(KEYINPUT20), .B(n1310), .Z(n1306) );
NOR2_X1 U1003 ( .A1(n1308), .A2(n1309), .ZN(n1310) );
XNOR2_X1 U1004 ( .A(n1311), .B(n1312), .ZN(n1309) );
XNOR2_X1 U1005 ( .A(n1249), .B(G104), .ZN(n1312) );
XNOR2_X1 U1006 ( .A(n1313), .B(n1137), .ZN(n1311) );
INV_X1 U1007 ( .A(G122), .ZN(n1137) );
XNOR2_X1 U1008 ( .A(KEYINPUT54), .B(KEYINPUT43), .ZN(n1313) );
XOR2_X1 U1009 ( .A(n1314), .B(n1315), .Z(n1308) );
XOR2_X1 U1010 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1011 ( .A(KEYINPUT35), .B(n1318), .ZN(n1317) );
NOR2_X1 U1012 ( .A1(G131), .A2(KEYINPUT22), .ZN(n1316) );
XOR2_X1 U1013 ( .A(n1319), .B(n1275), .Z(n1314) );
XNOR2_X1 U1014 ( .A(n1122), .B(n1320), .ZN(n1275) );
XOR2_X1 U1015 ( .A(KEYINPUT37), .B(G140), .Z(n1320) );
XNOR2_X1 U1016 ( .A(n1321), .B(n1322), .ZN(n1319) );
NAND2_X1 U1017 ( .A1(n1289), .A2(G214), .ZN(n1321) );
NOR2_X1 U1018 ( .A1(G953), .A2(G237), .ZN(n1289) );
NOR2_X1 U1019 ( .A1(n1066), .A2(n1241), .ZN(n1210) );
NAND2_X1 U1020 ( .A1(n1205), .A2(n1209), .ZN(n1241) );
NAND2_X1 U1021 ( .A1(n1323), .A2(n1081), .ZN(n1209) );
NAND3_X1 U1022 ( .A1(n1239), .A2(n1105), .A3(G952), .ZN(n1081) );
NAND4_X1 U1023 ( .A1(G953), .A2(G902), .A3(n1239), .A4(n1324), .ZN(n1323) );
INV_X1 U1024 ( .A(G898), .ZN(n1324) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1239) );
NOR2_X1 U1026 ( .A1(n1080), .A2(n1079), .ZN(n1205) );
AND2_X1 U1027 ( .A1(G214), .A2(n1325), .ZN(n1079) );
INV_X1 U1028 ( .A(n1231), .ZN(n1080) );
XNOR2_X1 U1029 ( .A(n1091), .B(n1095), .ZN(n1231) );
NAND2_X1 U1030 ( .A1(G210), .A2(n1325), .ZN(n1095) );
NAND2_X1 U1031 ( .A1(n1261), .A2(n1326), .ZN(n1325) );
INV_X1 U1032 ( .A(G237), .ZN(n1326) );
INV_X1 U1033 ( .A(n1093), .ZN(n1091) );
NAND2_X1 U1034 ( .A1(n1327), .A2(n1261), .ZN(n1093) );
XNOR2_X1 U1035 ( .A(n1159), .B(n1328), .ZN(n1327) );
XNOR2_X1 U1036 ( .A(n1329), .B(n1330), .ZN(n1328) );
INV_X1 U1037 ( .A(n1178), .ZN(n1330) );
XNOR2_X1 U1038 ( .A(n1331), .B(n1332), .ZN(n1178) );
XOR2_X1 U1039 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1040 ( .A(KEYINPUT56), .B(n1335), .ZN(n1334) );
NOR2_X1 U1041 ( .A1(KEYINPUT55), .A2(n1336), .ZN(n1335) );
XNOR2_X1 U1042 ( .A(G122), .B(G110), .ZN(n1336) );
NAND2_X1 U1043 ( .A1(G224), .A2(n1105), .ZN(n1333) );
INV_X1 U1044 ( .A(G953), .ZN(n1105) );
XNOR2_X1 U1045 ( .A(n1140), .B(n1139), .ZN(n1331) );
XNOR2_X1 U1046 ( .A(n1249), .B(n1288), .ZN(n1139) );
XNOR2_X1 U1047 ( .A(G116), .B(n1243), .ZN(n1288) );
INV_X1 U1048 ( .A(G119), .ZN(n1243) );
INV_X1 U1049 ( .A(G113), .ZN(n1249) );
AND2_X1 U1050 ( .A1(n1337), .A2(n1338), .ZN(n1140) );
NAND2_X1 U1051 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
INV_X1 U1052 ( .A(G101), .ZN(n1340) );
XNOR2_X1 U1053 ( .A(n1341), .B(n1342), .ZN(n1339) );
NAND2_X1 U1054 ( .A1(G101), .A2(n1343), .ZN(n1337) );
XNOR2_X1 U1055 ( .A(G104), .B(n1342), .ZN(n1343) );
NOR2_X1 U1056 ( .A1(G107), .A2(KEYINPUT2), .ZN(n1342) );
NAND2_X1 U1057 ( .A1(KEYINPUT58), .A2(n1122), .ZN(n1329) );
INV_X1 U1058 ( .A(G125), .ZN(n1122) );
INV_X1 U1059 ( .A(n1214), .ZN(n1159) );
NAND2_X1 U1060 ( .A1(n1344), .A2(n1345), .ZN(n1214) );
NAND2_X1 U1061 ( .A1(n1301), .A2(n1266), .ZN(n1345) );
NAND2_X1 U1062 ( .A1(n1346), .A2(n1322), .ZN(n1344) );
INV_X1 U1063 ( .A(n1266), .ZN(n1322) );
XNOR2_X1 U1064 ( .A(n1301), .B(KEYINPUT25), .ZN(n1346) );
XOR2_X1 U1065 ( .A(G128), .B(G143), .Z(n1301) );
INV_X1 U1066 ( .A(n1234), .ZN(n1066) );
NOR2_X1 U1067 ( .A1(n1069), .A2(n1068), .ZN(n1234) );
INV_X1 U1068 ( .A(n1256), .ZN(n1068) );
NAND2_X1 U1069 ( .A1(G221), .A2(n1260), .ZN(n1256) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1261), .ZN(n1260) );
XOR2_X1 U1071 ( .A(n1347), .B(G469), .Z(n1069) );
NAND2_X1 U1072 ( .A1(n1348), .A2(n1261), .ZN(n1347) );
INV_X1 U1073 ( .A(G902), .ZN(n1261) );
XOR2_X1 U1074 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1075 ( .A(n1351), .B(n1352), .Z(n1350) );
XNOR2_X1 U1076 ( .A(n1106), .B(G140), .ZN(n1352) );
INV_X1 U1077 ( .A(G227), .ZN(n1106) );
NOR2_X1 U1078 ( .A1(n1353), .A2(KEYINPUT38), .ZN(n1351) );
NOR2_X1 U1079 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1080 ( .A(n1356), .B(KEYINPUT50), .Z(n1355) );
NAND2_X1 U1081 ( .A1(n1357), .A2(n1116), .ZN(n1356) );
NOR2_X1 U1082 ( .A1(n1116), .A2(n1357), .ZN(n1354) );
XNOR2_X1 U1083 ( .A(n1168), .B(KEYINPUT51), .ZN(n1357) );
XOR2_X1 U1084 ( .A(G101), .B(n1358), .Z(n1168) );
XNOR2_X1 U1085 ( .A(G107), .B(n1341), .ZN(n1358) );
INV_X1 U1086 ( .A(G104), .ZN(n1341) );
XOR2_X1 U1087 ( .A(n1359), .B(n1360), .Z(n1116) );
XNOR2_X1 U1088 ( .A(KEYINPUT40), .B(n1361), .ZN(n1360) );
INV_X1 U1089 ( .A(G128), .ZN(n1361) );
NAND2_X1 U1090 ( .A1(n1362), .A2(n1363), .ZN(n1359) );
NAND2_X1 U1091 ( .A1(n1266), .A2(n1318), .ZN(n1363) );
XOR2_X1 U1092 ( .A(KEYINPUT53), .B(n1364), .Z(n1362) );
NOR2_X1 U1093 ( .A1(n1266), .A2(n1318), .ZN(n1364) );
INV_X1 U1094 ( .A(G143), .ZN(n1318) );
XOR2_X1 U1095 ( .A(G146), .B(KEYINPUT23), .Z(n1266) );
XNOR2_X1 U1096 ( .A(n1170), .B(n1365), .ZN(n1349) );
NOR2_X1 U1097 ( .A1(G110), .A2(KEYINPUT12), .ZN(n1365) );
XOR2_X1 U1098 ( .A(G131), .B(n1124), .Z(n1170) );
XNOR2_X1 U1099 ( .A(n1300), .B(n1276), .ZN(n1124) );
XOR2_X1 U1100 ( .A(G137), .B(KEYINPUT16), .Z(n1276) );
XNOR2_X1 U1101 ( .A(G134), .B(KEYINPUT31), .ZN(n1300) );
endmodule


