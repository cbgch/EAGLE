//Key = 1001100010000001011110000000101010001101111111100001100001000011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281;

XOR2_X1 U707 ( .A(n975), .B(n976), .Z(G9) );
NOR2_X1 U708 ( .A1(n977), .A2(n978), .ZN(G75) );
NOR2_X1 U709 ( .A1(n979), .A2(n980), .ZN(n978) );
INV_X1 U710 ( .A(n981), .ZN(n979) );
NOR3_X1 U711 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n977) );
NOR4_X1 U712 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n983) );
NOR2_X1 U713 ( .A1(n989), .A2(n990), .ZN(n986) );
NOR2_X1 U714 ( .A1(n991), .A2(n992), .ZN(n990) );
NOR2_X1 U715 ( .A1(n993), .A2(n994), .ZN(n991) );
NOR2_X1 U716 ( .A1(n995), .A2(n996), .ZN(n993) );
NOR2_X1 U717 ( .A1(n997), .A2(n998), .ZN(n989) );
NOR2_X1 U718 ( .A1(n999), .A2(n1000), .ZN(n997) );
NOR2_X1 U719 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NAND3_X1 U720 ( .A1(n981), .A2(n1003), .A3(n1004), .ZN(n982) );
NAND4_X1 U721 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n1004) );
NAND2_X1 U722 ( .A1(n985), .A2(n1009), .ZN(n1008) );
NAND3_X1 U723 ( .A1(n1010), .A2(n1011), .A3(KEYINPUT47), .ZN(n1009) );
INV_X1 U724 ( .A(n1012), .ZN(n985) );
NAND3_X1 U725 ( .A1(n1013), .A2(n1014), .A3(n1012), .ZN(n1007) );
NAND2_X1 U726 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U727 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U728 ( .A1(n1011), .A2(n1019), .ZN(n1013) );
NAND2_X1 U729 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
OR2_X1 U730 ( .A1(n1022), .A2(KEYINPUT47), .ZN(n1021) );
NAND4_X1 U731 ( .A1(n1023), .A2(n1005), .A3(n1024), .A4(n1025), .ZN(n981) );
NOR4_X1 U732 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1025) );
XNOR2_X1 U733 ( .A(n1030), .B(KEYINPUT42), .ZN(n1028) );
XOR2_X1 U734 ( .A(n1031), .B(n1032), .Z(n1027) );
NOR2_X1 U735 ( .A1(G472), .A2(KEYINPUT6), .ZN(n1032) );
INV_X1 U736 ( .A(n1002), .ZN(n1026) );
XOR2_X1 U737 ( .A(n1033), .B(n1034), .Z(n1024) );
XOR2_X1 U738 ( .A(KEYINPUT31), .B(G469), .Z(n1034) );
NAND2_X1 U739 ( .A1(KEYINPUT40), .A2(n1035), .ZN(n1033) );
XNOR2_X1 U740 ( .A(n1036), .B(n1037), .ZN(n1023) );
XOR2_X1 U741 ( .A(n1038), .B(n1039), .Z(G72) );
XOR2_X1 U742 ( .A(n1040), .B(n1041), .Z(n1039) );
NOR2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
XOR2_X1 U744 ( .A(n1003), .B(KEYINPUT41), .Z(n1043) );
NOR2_X1 U745 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
XOR2_X1 U746 ( .A(KEYINPUT35), .B(n1046), .Z(n1045) );
NOR2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1040) );
XOR2_X1 U748 ( .A(n1049), .B(n1050), .Z(n1048) );
XOR2_X1 U749 ( .A(G134), .B(n1051), .Z(n1050) );
XOR2_X1 U750 ( .A(KEYINPUT27), .B(G140), .Z(n1051) );
XOR2_X1 U751 ( .A(n1052), .B(n1053), .Z(n1049) );
XNOR2_X1 U752 ( .A(G125), .B(n1054), .ZN(n1052) );
NOR2_X1 U753 ( .A1(n1055), .A2(n1003), .ZN(n1038) );
NOR2_X1 U754 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XOR2_X1 U755 ( .A(n1058), .B(n1059), .Z(G69) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1003), .ZN(n1059) );
AND2_X1 U757 ( .A1(G224), .A2(G898), .ZN(n1060) );
NAND2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(n1058) );
NAND2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U760 ( .A1(n1065), .A2(n1066), .ZN(n1061) );
XNOR2_X1 U761 ( .A(n1063), .B(KEYINPUT33), .ZN(n1066) );
AND2_X1 U762 ( .A1(n1003), .A2(n1067), .ZN(n1063) );
INV_X1 U763 ( .A(n1064), .ZN(n1065) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U766 ( .A(n1072), .B(n1073), .Z(n1068) );
XOR2_X1 U767 ( .A(KEYINPUT26), .B(n1074), .Z(n1073) );
NOR3_X1 U768 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(G66) );
NOR2_X1 U769 ( .A1(n980), .A2(n1078), .ZN(n1077) );
INV_X1 U770 ( .A(KEYINPUT11), .ZN(n1078) );
NOR2_X1 U771 ( .A1(KEYINPUT11), .A2(n1079), .ZN(n1076) );
XOR2_X1 U772 ( .A(n1080), .B(n1081), .Z(n1075) );
NOR2_X1 U773 ( .A1(n1037), .A2(n1082), .ZN(n1081) );
NAND2_X1 U774 ( .A1(KEYINPUT3), .A2(n1083), .ZN(n1080) );
NOR2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(G63) );
XOR2_X1 U776 ( .A(n1086), .B(n1087), .Z(n1085) );
NAND3_X1 U777 ( .A1(G478), .A2(n1088), .A3(n1089), .ZN(n1086) );
XNOR2_X1 U778 ( .A(KEYINPUT43), .B(n984), .ZN(n1088) );
NOR3_X1 U779 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(G60) );
NOR2_X1 U780 ( .A1(n980), .A2(n1093), .ZN(n1092) );
INV_X1 U781 ( .A(KEYINPUT2), .ZN(n1093) );
OR2_X1 U782 ( .A1(G952), .A2(G953), .ZN(n980) );
NOR2_X1 U783 ( .A1(KEYINPUT2), .A2(n1079), .ZN(n1091) );
INV_X1 U784 ( .A(n1084), .ZN(n1079) );
XOR2_X1 U785 ( .A(n1094), .B(n1095), .Z(n1090) );
NAND2_X1 U786 ( .A1(n1096), .A2(G475), .ZN(n1094) );
NAND3_X1 U787 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(G6) );
NAND3_X1 U788 ( .A1(n994), .A2(n1100), .A3(n1101), .ZN(n1099) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND2_X1 U790 ( .A1(KEYINPUT18), .A2(n1104), .ZN(n1103) );
NAND3_X1 U791 ( .A1(G104), .A2(n1105), .A3(n1102), .ZN(n1098) );
INV_X1 U792 ( .A(KEYINPUT13), .ZN(n1102) );
NAND3_X1 U793 ( .A1(n1101), .A2(n994), .A3(KEYINPUT18), .ZN(n1105) );
NAND2_X1 U794 ( .A1(KEYINPUT13), .A2(n1104), .ZN(n1097) );
NOR2_X1 U795 ( .A1(n1084), .A2(n1106), .ZN(G57) );
XOR2_X1 U796 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U798 ( .A1(n1096), .A2(G472), .ZN(n1109) );
XOR2_X1 U799 ( .A(n1111), .B(n1112), .Z(n1107) );
NOR2_X1 U800 ( .A1(n1084), .A2(n1113), .ZN(G54) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U802 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U803 ( .A(KEYINPUT58), .B(KEYINPUT39), .Z(n1117) );
NOR2_X1 U804 ( .A1(KEYINPUT16), .A2(n1118), .ZN(n1116) );
XOR2_X1 U805 ( .A(n1119), .B(n1120), .Z(n1118) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1114) );
XOR2_X1 U807 ( .A(n1123), .B(n1053), .Z(n1121) );
NAND2_X1 U808 ( .A1(n1096), .A2(G469), .ZN(n1123) );
INV_X1 U809 ( .A(n1082), .ZN(n1096) );
NOR2_X1 U810 ( .A1(n1084), .A2(n1124), .ZN(G51) );
XNOR2_X1 U811 ( .A(n1125), .B(n1126), .ZN(n1124) );
XNOR2_X1 U812 ( .A(n1127), .B(n1128), .ZN(n1125) );
NOR3_X1 U813 ( .A1(n1082), .A2(KEYINPUT50), .A3(n1129), .ZN(n1128) );
NAND2_X1 U814 ( .A1(n1089), .A2(n984), .ZN(n1082) );
OR3_X1 U815 ( .A1(n1044), .A2(n1046), .A3(n1067), .ZN(n984) );
NAND4_X1 U816 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1067) );
AND4_X1 U817 ( .A1(n976), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1133) );
NAND4_X1 U818 ( .A1(n1000), .A2(n1137), .A3(n1015), .A4(n1138), .ZN(n976) );
NAND2_X1 U819 ( .A1(n994), .A2(n1139), .ZN(n1132) );
NAND2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U821 ( .A(KEYINPUT17), .B(n1101), .Z(n1140) );
NOR4_X1 U822 ( .A1(n1017), .A2(n1142), .A3(n987), .A4(n1143), .ZN(n1101) );
NAND3_X1 U823 ( .A1(n1137), .A2(n1138), .A3(n1144), .ZN(n1130) );
INV_X1 U824 ( .A(n1145), .ZN(n1046) );
NAND4_X1 U825 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1044) );
NOR4_X1 U826 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1149) );
XOR2_X1 U827 ( .A(n1154), .B(KEYINPUT28), .Z(n1089) );
NOR2_X1 U828 ( .A1(KEYINPUT9), .A2(n1155), .ZN(n1127) );
XOR2_X1 U829 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U830 ( .A1(KEYINPUT63), .A2(n1158), .ZN(n1157) );
NOR2_X1 U831 ( .A1(n1003), .A2(G952), .ZN(n1084) );
XNOR2_X1 U832 ( .A(n1148), .B(n1159), .ZN(G48) );
NOR2_X1 U833 ( .A1(KEYINPUT14), .A2(n1160), .ZN(n1159) );
NAND3_X1 U834 ( .A1(n1161), .A2(n994), .A3(n1162), .ZN(n1148) );
XOR2_X1 U835 ( .A(G143), .B(n1163), .Z(G45) );
NOR2_X1 U836 ( .A1(KEYINPUT38), .A2(n1146), .ZN(n1163) );
NAND4_X1 U837 ( .A1(n1164), .A2(n994), .A3(n1029), .A4(n1165), .ZN(n1146) );
XNOR2_X1 U838 ( .A(G140), .B(n1147), .ZN(G42) );
NAND3_X1 U839 ( .A1(n1005), .A2(n1161), .A3(n1166), .ZN(n1147) );
NOR3_X1 U840 ( .A1(n1022), .A2(n1167), .A3(n1142), .ZN(n1166) );
XOR2_X1 U841 ( .A(n1168), .B(n1169), .Z(G39) );
XOR2_X1 U842 ( .A(KEYINPUT51), .B(G137), .Z(n1169) );
NAND2_X1 U843 ( .A1(KEYINPUT37), .A2(n1152), .ZN(n1168) );
AND3_X1 U844 ( .A1(n1162), .A2(n1011), .A3(n1005), .ZN(n1152) );
XOR2_X1 U845 ( .A(G134), .B(n1153), .Z(G36) );
AND3_X1 U846 ( .A1(n1005), .A2(n1137), .A3(n1164), .ZN(n1153) );
XOR2_X1 U847 ( .A(n1170), .B(G131), .Z(G33) );
NAND2_X1 U848 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
OR2_X1 U849 ( .A1(n1145), .A2(KEYINPUT54), .ZN(n1172) );
NAND3_X1 U850 ( .A1(n1005), .A2(n1161), .A3(n1164), .ZN(n1145) );
NOR3_X1 U851 ( .A1(n1142), .A2(n1167), .A3(n1020), .ZN(n1164) );
NAND4_X1 U852 ( .A1(n1167), .A2(n1005), .A3(n1173), .A4(KEYINPUT54), .ZN(n1171) );
NOR3_X1 U853 ( .A1(n1017), .A2(n1142), .A3(n1020), .ZN(n1173) );
INV_X1 U854 ( .A(n998), .ZN(n1005) );
NAND2_X1 U855 ( .A1(n1174), .A2(n996), .ZN(n998) );
INV_X1 U856 ( .A(n1175), .ZN(n1167) );
XOR2_X1 U857 ( .A(n1151), .B(n1176), .Z(G30) );
XOR2_X1 U858 ( .A(KEYINPUT10), .B(G128), .Z(n1176) );
AND3_X1 U859 ( .A1(n1137), .A2(n994), .A3(n1162), .ZN(n1151) );
AND4_X1 U860 ( .A1(n1177), .A2(n1178), .A3(n1000), .A4(n1175), .ZN(n1162) );
XOR2_X1 U861 ( .A(n1131), .B(n1179), .Z(G3) );
NAND2_X1 U862 ( .A1(KEYINPUT20), .A2(G101), .ZN(n1179) );
NAND2_X1 U863 ( .A1(n1180), .A2(n1181), .ZN(n1131) );
INV_X1 U864 ( .A(n1020), .ZN(n1180) );
XOR2_X1 U865 ( .A(G125), .B(n1150), .Z(G27) );
AND4_X1 U866 ( .A1(n994), .A2(n1175), .A3(n1010), .A4(n1182), .ZN(n1150) );
NOR2_X1 U867 ( .A1(n992), .A2(n1017), .ZN(n1182) );
NAND2_X1 U868 ( .A1(n1183), .A2(n1184), .ZN(n1175) );
NAND3_X1 U869 ( .A1(n1185), .A2(n1012), .A3(n1047), .ZN(n1184) );
AND2_X1 U870 ( .A1(n1070), .A2(n1057), .ZN(n1047) );
INV_X1 U871 ( .A(G900), .ZN(n1057) );
INV_X1 U872 ( .A(n1186), .ZN(n994) );
XOR2_X1 U873 ( .A(n1187), .B(n1136), .Z(G24) );
NAND4_X1 U874 ( .A1(n1006), .A2(n1015), .A3(n1188), .A4(n1138), .ZN(n1136) );
AND2_X1 U875 ( .A1(n1165), .A2(n1029), .ZN(n1188) );
INV_X1 U876 ( .A(n987), .ZN(n1015) );
NAND2_X1 U877 ( .A1(n1189), .A2(n1190), .ZN(n987) );
XOR2_X1 U878 ( .A(G119), .B(n1191), .Z(G21) );
NOR2_X1 U879 ( .A1(n1192), .A2(n1186), .ZN(n1191) );
XOR2_X1 U880 ( .A(n1141), .B(KEYINPUT21), .Z(n1192) );
NAND3_X1 U881 ( .A1(n1177), .A2(n1006), .A3(n1193), .ZN(n1141) );
NOR3_X1 U882 ( .A1(n988), .A2(n1143), .A3(n1190), .ZN(n1193) );
INV_X1 U883 ( .A(n1011), .ZN(n988) );
INV_X1 U884 ( .A(n992), .ZN(n1006) );
XOR2_X1 U885 ( .A(n1194), .B(n1195), .Z(G18) );
NAND2_X1 U886 ( .A1(KEYINPUT62), .A2(G116), .ZN(n1195) );
NAND4_X1 U887 ( .A1(n1196), .A2(n1144), .A3(n1137), .A4(n1197), .ZN(n1194) );
INV_X1 U888 ( .A(n1018), .ZN(n1137) );
NAND2_X1 U889 ( .A1(n1198), .A2(n1165), .ZN(n1018) );
XOR2_X1 U890 ( .A(n1030), .B(KEYINPUT23), .Z(n1165) );
XNOR2_X1 U891 ( .A(n1029), .B(KEYINPUT25), .ZN(n1198) );
XOR2_X1 U892 ( .A(n1186), .B(KEYINPUT8), .Z(n1196) );
XNOR2_X1 U893 ( .A(G113), .B(n1135), .ZN(G15) );
NAND3_X1 U894 ( .A1(n1144), .A2(n1138), .A3(n1161), .ZN(n1135) );
INV_X1 U895 ( .A(n1017), .ZN(n1161) );
NAND2_X1 U896 ( .A1(n1199), .A2(n1029), .ZN(n1017) );
INV_X1 U897 ( .A(n1030), .ZN(n1199) );
NOR2_X1 U898 ( .A1(n992), .A2(n1020), .ZN(n1144) );
NAND2_X1 U899 ( .A1(n1177), .A2(n1190), .ZN(n1020) );
INV_X1 U900 ( .A(n1178), .ZN(n1190) );
XOR2_X1 U901 ( .A(n1189), .B(KEYINPUT36), .Z(n1177) );
NAND2_X1 U902 ( .A1(n1200), .A2(n1002), .ZN(n992) );
XNOR2_X1 U903 ( .A(G110), .B(n1134), .ZN(G12) );
NAND2_X1 U904 ( .A1(n1010), .A2(n1181), .ZN(n1134) );
AND3_X1 U905 ( .A1(n1000), .A2(n1138), .A3(n1011), .ZN(n1181) );
NOR2_X1 U906 ( .A1(n1029), .A2(n1030), .ZN(n1011) );
XNOR2_X1 U907 ( .A(n1201), .B(G478), .ZN(n1030) );
NAND2_X1 U908 ( .A1(n1087), .A2(n1154), .ZN(n1201) );
XNOR2_X1 U909 ( .A(n1202), .B(n1203), .ZN(n1087) );
XOR2_X1 U910 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U911 ( .A(G134), .B(G116), .Z(n1205) );
XOR2_X1 U912 ( .A(KEYINPUT55), .B(G143), .Z(n1204) );
XOR2_X1 U913 ( .A(n1206), .B(n1207), .Z(n1202) );
XNOR2_X1 U914 ( .A(n1208), .B(n1209), .ZN(n1207) );
NOR2_X1 U915 ( .A1(G128), .A2(KEYINPUT59), .ZN(n1209) );
NAND2_X1 U916 ( .A1(KEYINPUT44), .A2(n1187), .ZN(n1208) );
XOR2_X1 U917 ( .A(n1210), .B(G107), .Z(n1206) );
NAND3_X1 U918 ( .A1(G234), .A2(n1003), .A3(G217), .ZN(n1210) );
XNOR2_X1 U919 ( .A(n1211), .B(G475), .ZN(n1029) );
NAND2_X1 U920 ( .A1(n1095), .A2(n1154), .ZN(n1211) );
XNOR2_X1 U921 ( .A(n1212), .B(n1213), .ZN(n1095) );
XOR2_X1 U922 ( .A(n1214), .B(n1215), .Z(n1213) );
XNOR2_X1 U923 ( .A(n1216), .B(n1217), .ZN(n1215) );
NOR2_X1 U924 ( .A1(KEYINPUT48), .A2(n1218), .ZN(n1217) );
XOR2_X1 U925 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U926 ( .A(G143), .B(G131), .Z(n1220) );
AND3_X1 U927 ( .A1(G214), .A2(n1003), .A3(n1221), .ZN(n1219) );
NAND2_X1 U928 ( .A1(KEYINPUT57), .A2(n1104), .ZN(n1216) );
XNOR2_X1 U929 ( .A(G113), .B(n1222), .ZN(n1212) );
XOR2_X1 U930 ( .A(G140), .B(G122), .Z(n1222) );
NOR2_X1 U931 ( .A1(n1186), .A2(n1143), .ZN(n1138) );
INV_X1 U932 ( .A(n1197), .ZN(n1143) );
NAND2_X1 U933 ( .A1(n1223), .A2(n1183), .ZN(n1197) );
NAND3_X1 U934 ( .A1(n1224), .A2(n1012), .A3(G952), .ZN(n1183) );
XOR2_X1 U935 ( .A(KEYINPUT32), .B(G953), .Z(n1224) );
NAND4_X1 U936 ( .A1(n1070), .A2(n1185), .A3(n1012), .A4(n1071), .ZN(n1223) );
INV_X1 U937 ( .A(G898), .ZN(n1071) );
NAND2_X1 U938 ( .A1(G237), .A2(G234), .ZN(n1012) );
XOR2_X1 U939 ( .A(G902), .B(KEYINPUT29), .Z(n1185) );
XOR2_X1 U940 ( .A(G953), .B(KEYINPUT53), .Z(n1070) );
NAND2_X1 U941 ( .A1(n995), .A2(n996), .ZN(n1186) );
NAND2_X1 U942 ( .A1(G214), .A2(n1225), .ZN(n996) );
INV_X1 U943 ( .A(n1174), .ZN(n995) );
XNOR2_X1 U944 ( .A(n1226), .B(n1129), .ZN(n1174) );
NAND2_X1 U945 ( .A1(G210), .A2(n1225), .ZN(n1129) );
NAND2_X1 U946 ( .A1(n1221), .A2(n1154), .ZN(n1225) );
NAND2_X1 U947 ( .A1(n1227), .A2(n1154), .ZN(n1226) );
XOR2_X1 U948 ( .A(n1228), .B(n1229), .Z(n1227) );
XNOR2_X1 U949 ( .A(n1126), .B(n1158), .ZN(n1229) );
XNOR2_X1 U950 ( .A(n1214), .B(n1230), .ZN(n1158) );
NAND2_X1 U951 ( .A1(n1231), .A2(n1232), .ZN(n1126) );
NAND2_X1 U952 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XOR2_X1 U953 ( .A(n1072), .B(KEYINPUT56), .Z(n1233) );
NAND2_X1 U954 ( .A1(n1235), .A2(n1074), .ZN(n1231) );
INV_X1 U955 ( .A(n1234), .ZN(n1074) );
XOR2_X1 U956 ( .A(KEYINPUT24), .B(n1236), .Z(n1235) );
INV_X1 U957 ( .A(n1072), .ZN(n1236) );
XOR2_X1 U958 ( .A(n1237), .B(n1238), .Z(n1072) );
XNOR2_X1 U959 ( .A(n1239), .B(n1240), .ZN(n1238) );
XOR2_X1 U960 ( .A(n1104), .B(n1241), .Z(n1240) );
NAND2_X1 U961 ( .A1(KEYINPUT4), .A2(n1111), .ZN(n1241) );
INV_X1 U962 ( .A(G104), .ZN(n1104) );
NAND2_X1 U963 ( .A1(KEYINPUT46), .A2(n975), .ZN(n1239) );
INV_X1 U964 ( .A(G107), .ZN(n975) );
XOR2_X1 U965 ( .A(G110), .B(n1187), .Z(n1237) );
INV_X1 U966 ( .A(G122), .ZN(n1187) );
XOR2_X1 U967 ( .A(n1156), .B(KEYINPUT7), .Z(n1228) );
NAND2_X1 U968 ( .A1(G224), .A2(n1003), .ZN(n1156) );
INV_X1 U969 ( .A(n1142), .ZN(n1000) );
NAND2_X1 U970 ( .A1(n1001), .A2(n1002), .ZN(n1142) );
NAND2_X1 U971 ( .A1(G221), .A2(n1242), .ZN(n1002) );
INV_X1 U972 ( .A(n1200), .ZN(n1001) );
XNOR2_X1 U973 ( .A(n1035), .B(G469), .ZN(n1200) );
AND2_X1 U974 ( .A1(n1243), .A2(n1154), .ZN(n1035) );
XOR2_X1 U975 ( .A(n1244), .B(n1245), .Z(n1243) );
XNOR2_X1 U976 ( .A(n1246), .B(n1247), .ZN(n1245) );
NOR2_X1 U977 ( .A1(KEYINPUT5), .A2(n1053), .ZN(n1247) );
XNOR2_X1 U978 ( .A(n1248), .B(n1249), .ZN(n1053) );
NAND3_X1 U979 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1248) );
NAND2_X1 U980 ( .A1(G146), .A2(n1253), .ZN(n1252) );
NAND2_X1 U981 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
INV_X1 U982 ( .A(KEYINPUT45), .ZN(n1255) );
NAND2_X1 U983 ( .A1(G143), .A2(n1256), .ZN(n1254) );
XOR2_X1 U984 ( .A(KEYINPUT15), .B(G146), .Z(n1256) );
NAND2_X1 U985 ( .A1(KEYINPUT45), .A2(n1257), .ZN(n1250) );
NAND2_X1 U986 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NAND3_X1 U987 ( .A1(KEYINPUT15), .A2(G143), .A3(n1160), .ZN(n1259) );
OR2_X1 U988 ( .A1(n1160), .A2(KEYINPUT15), .ZN(n1258) );
INV_X1 U989 ( .A(G146), .ZN(n1160) );
NAND2_X1 U990 ( .A1(KEYINPUT30), .A2(n1119), .ZN(n1246) );
NOR2_X1 U991 ( .A1(n1056), .A2(G953), .ZN(n1119) );
INV_X1 U992 ( .A(G227), .ZN(n1056) );
XNOR2_X1 U993 ( .A(n1122), .B(n1120), .ZN(n1244) );
XNOR2_X1 U994 ( .A(n1260), .B(n1261), .ZN(n1122) );
XOR2_X1 U995 ( .A(G107), .B(G104), .Z(n1261) );
XOR2_X1 U996 ( .A(n1111), .B(n1262), .Z(n1260) );
INV_X1 U997 ( .A(G101), .ZN(n1111) );
INV_X1 U998 ( .A(n1022), .ZN(n1010) );
NAND2_X1 U999 ( .A1(n1178), .A2(n1189), .ZN(n1022) );
XOR2_X1 U1000 ( .A(n1031), .B(G472), .Z(n1189) );
NAND2_X1 U1001 ( .A1(n1263), .A2(n1264), .ZN(n1031) );
XOR2_X1 U1002 ( .A(n1110), .B(n1265), .Z(n1264) );
XOR2_X1 U1003 ( .A(n1112), .B(n1266), .Z(n1265) );
NOR2_X1 U1004 ( .A1(G101), .A2(KEYINPUT60), .ZN(n1266) );
NAND3_X1 U1005 ( .A1(n1221), .A2(n1003), .A3(G210), .ZN(n1112) );
INV_X1 U1006 ( .A(G237), .ZN(n1221) );
XOR2_X1 U1007 ( .A(n1267), .B(n1268), .Z(n1110) );
XOR2_X1 U1008 ( .A(n1230), .B(n1269), .Z(n1268) );
XOR2_X1 U1009 ( .A(KEYINPUT12), .B(G146), .Z(n1269) );
XNOR2_X1 U1010 ( .A(n1270), .B(n1271), .ZN(n1230) );
NOR2_X1 U1011 ( .A1(KEYINPUT34), .A2(n1249), .ZN(n1271) );
XOR2_X1 U1012 ( .A(G128), .B(KEYINPUT1), .Z(n1249) );
NAND2_X1 U1013 ( .A1(KEYINPUT19), .A2(n1253), .ZN(n1270) );
INV_X1 U1014 ( .A(G143), .ZN(n1253) );
XOR2_X1 U1015 ( .A(n1234), .B(n1262), .Z(n1267) );
XOR2_X1 U1016 ( .A(n1054), .B(n1272), .Z(n1262) );
NOR2_X1 U1017 ( .A1(G134), .A2(KEYINPUT22), .ZN(n1272) );
XOR2_X1 U1018 ( .A(G131), .B(G137), .Z(n1054) );
XNOR2_X1 U1019 ( .A(G113), .B(n1273), .ZN(n1234) );
XOR2_X1 U1020 ( .A(G119), .B(G116), .Z(n1273) );
XOR2_X1 U1021 ( .A(KEYINPUT52), .B(G902), .Z(n1263) );
XNOR2_X1 U1022 ( .A(n1274), .B(n1037), .ZN(n1178) );
NAND2_X1 U1023 ( .A1(G217), .A2(n1242), .ZN(n1037) );
NAND2_X1 U1024 ( .A1(G234), .A2(n1154), .ZN(n1242) );
NAND2_X1 U1025 ( .A1(KEYINPUT0), .A2(n1036), .ZN(n1274) );
NAND2_X1 U1026 ( .A1(n1083), .A2(n1154), .ZN(n1036) );
INV_X1 U1027 ( .A(G902), .ZN(n1154) );
XNOR2_X1 U1028 ( .A(n1275), .B(n1276), .ZN(n1083) );
XOR2_X1 U1029 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1030 ( .A(G137), .B(G128), .Z(n1278) );
XOR2_X1 U1031 ( .A(KEYINPUT61), .B(KEYINPUT49), .Z(n1277) );
XOR2_X1 U1032 ( .A(n1279), .B(n1280), .Z(n1275) );
XOR2_X1 U1033 ( .A(n1214), .B(n1120), .Z(n1280) );
XOR2_X1 U1034 ( .A(G110), .B(G140), .Z(n1120) );
XOR2_X1 U1035 ( .A(G125), .B(G146), .Z(n1214) );
XOR2_X1 U1036 ( .A(n1281), .B(G119), .Z(n1279) );
NAND3_X1 U1037 ( .A1(G234), .A2(n1003), .A3(G221), .ZN(n1281) );
INV_X1 U1038 ( .A(G953), .ZN(n1003) );
endmodule


