//Key = 0100011010001001101011111110010000101010001010100000011011110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336;

XNOR2_X1 U747 ( .A(n1022), .B(n1023), .ZN(G9) );
NOR2_X1 U748 ( .A1(KEYINPUT0), .A2(n1024), .ZN(n1023) );
NAND4_X1 U749 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(G75) );
NOR3_X1 U750 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND2_X1 U751 ( .A1(n1032), .A2(n1033), .ZN(n1027) );
NAND2_X1 U752 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND4_X1 U753 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND2_X1 U754 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND2_X1 U755 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
OR2_X1 U757 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1048), .A2(n1049), .ZN(n1040) );
NAND3_X1 U759 ( .A1(n1042), .A2(n1050), .A3(n1048), .ZN(n1034) );
NAND2_X1 U760 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U761 ( .A1(n1053), .A2(n1054), .A3(n1036), .ZN(n1052) );
NAND2_X1 U762 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XNOR2_X1 U763 ( .A(n1037), .B(KEYINPUT61), .ZN(n1056) );
INV_X1 U764 ( .A(n1039), .ZN(n1055) );
NAND3_X1 U765 ( .A1(n1057), .A2(n1058), .A3(n1039), .ZN(n1053) );
NAND2_X1 U766 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND2_X1 U767 ( .A1(n1061), .A2(n1037), .ZN(n1051) );
INV_X1 U768 ( .A(n1062), .ZN(n1032) );
NAND4_X1 U769 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1025) );
NOR3_X1 U770 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1066) );
XOR2_X1 U771 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U772 ( .A1(n1072), .A2(KEYINPUT3), .ZN(n1071) );
XOR2_X1 U773 ( .A(n1073), .B(n1074), .Z(n1068) );
NOR2_X1 U774 ( .A1(G475), .A2(KEYINPUT4), .ZN(n1074) );
NAND3_X1 U775 ( .A1(n1039), .A2(n1046), .A3(n1075), .ZN(n1067) );
NAND2_X1 U776 ( .A1(G478), .A2(n1076), .ZN(n1075) );
NOR3_X1 U777 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1065) );
NOR3_X1 U778 ( .A1(n1080), .A2(KEYINPUT27), .A3(n1081), .ZN(n1079) );
INV_X1 U779 ( .A(G469), .ZN(n1080) );
NOR2_X1 U780 ( .A1(G469), .A2(n1082), .ZN(n1078) );
NOR2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U782 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U783 ( .A1(KEYINPUT27), .A2(n1081), .ZN(n1085) );
INV_X1 U784 ( .A(n1087), .ZN(n1081) );
AND2_X1 U785 ( .A1(n1087), .A2(n1086), .ZN(n1083) );
XOR2_X1 U786 ( .A(KEYINPUT33), .B(KEYINPUT14), .Z(n1086) );
XOR2_X1 U787 ( .A(KEYINPUT15), .B(n1088), .Z(n1064) );
XOR2_X1 U788 ( .A(n1089), .B(n1090), .Z(G72) );
NOR2_X1 U789 ( .A1(n1091), .A2(n1026), .ZN(n1090) );
AND2_X1 U790 ( .A1(G227), .A2(G900), .ZN(n1091) );
NOR2_X1 U791 ( .A1(KEYINPUT51), .A2(n1092), .ZN(n1089) );
XOR2_X1 U792 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR3_X1 U793 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1094) );
NOR2_X1 U794 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
XOR2_X1 U796 ( .A(n1099), .B(KEYINPUT57), .Z(n1101) );
XOR2_X1 U797 ( .A(n1102), .B(n1103), .Z(n1099) );
XNOR2_X1 U798 ( .A(n1104), .B(n1105), .ZN(n1103) );
NAND2_X1 U799 ( .A1(KEYINPUT5), .A2(n1106), .ZN(n1104) );
XOR2_X1 U800 ( .A(n1107), .B(n1108), .Z(n1102) );
NOR2_X1 U801 ( .A1(KEYINPUT48), .A2(n1109), .ZN(n1108) );
XNOR2_X1 U802 ( .A(G134), .B(G140), .ZN(n1107) );
INV_X1 U803 ( .A(n1098), .ZN(n1100) );
XOR2_X1 U804 ( .A(n1110), .B(n1111), .Z(n1098) );
NAND2_X1 U805 ( .A1(n1026), .A2(n1031), .ZN(n1093) );
NAND2_X1 U806 ( .A1(n1112), .A2(n1113), .ZN(G69) );
NAND3_X1 U807 ( .A1(n1114), .A2(n1115), .A3(G953), .ZN(n1113) );
NAND2_X1 U808 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U809 ( .A1(G898), .A2(G224), .ZN(n1114) );
NAND3_X1 U810 ( .A1(n1118), .A2(n1117), .A3(n1119), .ZN(n1112) );
XNOR2_X1 U811 ( .A(n1116), .B(n1120), .ZN(n1119) );
NAND2_X1 U812 ( .A1(n1026), .A2(n1121), .ZN(n1120) );
NAND2_X1 U813 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
INV_X1 U814 ( .A(n1029), .ZN(n1123) );
XOR2_X1 U815 ( .A(n1030), .B(KEYINPUT24), .Z(n1122) );
AND3_X1 U816 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1116) );
INV_X1 U817 ( .A(n1127), .ZN(n1126) );
NAND2_X1 U818 ( .A1(n1128), .A2(n1129), .ZN(n1125) );
NAND2_X1 U819 ( .A1(n1130), .A2(n1131), .ZN(n1124) );
XNOR2_X1 U820 ( .A(n1128), .B(KEYINPUT19), .ZN(n1131) );
AND3_X1 U821 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1128) );
NAND2_X1 U822 ( .A1(KEYINPUT47), .A2(n1135), .ZN(n1134) );
NAND3_X1 U823 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1133) );
INV_X1 U824 ( .A(KEYINPUT47), .ZN(n1137) );
OR2_X1 U825 ( .A1(n1138), .A2(n1136), .ZN(n1132) );
NOR2_X1 U826 ( .A1(n1139), .A2(n1135), .ZN(n1136) );
INV_X1 U827 ( .A(KEYINPUT54), .ZN(n1139) );
INV_X1 U828 ( .A(n1129), .ZN(n1130) );
INV_X1 U829 ( .A(KEYINPUT41), .ZN(n1117) );
NAND2_X1 U830 ( .A1(G953), .A2(n1140), .ZN(n1118) );
NOR2_X1 U831 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XOR2_X1 U832 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U833 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U834 ( .A1(KEYINPUT1), .A2(n1147), .ZN(n1143) );
NOR2_X1 U835 ( .A1(n1141), .A2(n1148), .ZN(G63) );
XOR2_X1 U836 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND2_X1 U837 ( .A1(n1151), .A2(G478), .ZN(n1149) );
NOR2_X1 U838 ( .A1(n1141), .A2(n1152), .ZN(G60) );
XOR2_X1 U839 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U840 ( .A1(n1151), .A2(G475), .ZN(n1153) );
XOR2_X1 U841 ( .A(G104), .B(n1155), .Z(G6) );
NOR2_X1 U842 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NOR2_X1 U843 ( .A1(n1141), .A2(n1158), .ZN(G57) );
NOR2_X1 U844 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U845 ( .A(KEYINPUT40), .B(n1161), .Z(n1160) );
NOR2_X1 U846 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U847 ( .A(G101), .B(n1164), .ZN(n1163) );
NOR2_X1 U848 ( .A1(n1165), .A2(n1166), .ZN(n1159) );
INV_X1 U849 ( .A(n1162), .ZN(n1166) );
XOR2_X1 U850 ( .A(n1167), .B(n1168), .Z(n1162) );
NOR2_X1 U851 ( .A1(KEYINPUT55), .A2(n1169), .ZN(n1168) );
NAND2_X1 U852 ( .A1(n1151), .A2(G472), .ZN(n1167) );
XOR2_X1 U853 ( .A(n1164), .B(G101), .Z(n1165) );
NAND2_X1 U854 ( .A1(KEYINPUT25), .A2(n1170), .ZN(n1164) );
NOR2_X1 U855 ( .A1(n1141), .A2(n1171), .ZN(G54) );
XOR2_X1 U856 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U857 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U858 ( .A(G110), .B(KEYINPUT16), .ZN(n1175) );
NAND2_X1 U859 ( .A1(n1151), .A2(G469), .ZN(n1174) );
XOR2_X1 U860 ( .A(n1176), .B(n1177), .Z(n1172) );
NOR2_X1 U861 ( .A1(n1141), .A2(n1178), .ZN(G51) );
XOR2_X1 U862 ( .A(n1179), .B(n1180), .Z(n1178) );
NAND2_X1 U863 ( .A1(n1151), .A2(n1181), .ZN(n1179) );
INV_X1 U864 ( .A(n1145), .ZN(n1151) );
NAND2_X1 U865 ( .A1(G902), .A2(n1182), .ZN(n1145) );
OR3_X1 U866 ( .A1(n1031), .A2(n1030), .A3(n1029), .ZN(n1182) );
NAND2_X1 U867 ( .A1(n1183), .A2(n1184), .ZN(n1029) );
NAND2_X1 U868 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U869 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U870 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
NAND2_X1 U871 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND2_X1 U872 ( .A1(n1061), .A2(n1193), .ZN(n1192) );
NAND2_X1 U873 ( .A1(n1194), .A2(n1195), .ZN(n1191) );
NAND2_X1 U874 ( .A1(n1196), .A2(n1061), .ZN(n1187) );
NAND4_X1 U875 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1022), .ZN(n1030) );
OR2_X1 U876 ( .A1(n1200), .A2(n1156), .ZN(n1022) );
NAND2_X1 U877 ( .A1(n1201), .A2(n1037), .ZN(n1156) );
NAND3_X1 U878 ( .A1(n1194), .A2(n1201), .A3(n1202), .ZN(n1197) );
XNOR2_X1 U879 ( .A(n1037), .B(KEYINPUT22), .ZN(n1202) );
NAND4_X1 U880 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1031) );
NOR4_X1 U881 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
INV_X1 U882 ( .A(n1211), .ZN(n1210) );
NAND2_X1 U883 ( .A1(n1212), .A2(n1049), .ZN(n1205) );
NAND2_X1 U884 ( .A1(n1157), .A2(n1200), .ZN(n1049) );
INV_X1 U885 ( .A(n1193), .ZN(n1200) );
INV_X1 U886 ( .A(n1213), .ZN(n1212) );
NOR2_X1 U887 ( .A1(n1026), .A2(G952), .ZN(n1141) );
XOR2_X1 U888 ( .A(G146), .B(n1214), .Z(G48) );
NOR2_X1 U889 ( .A1(n1157), .A2(n1213), .ZN(n1214) );
XOR2_X1 U890 ( .A(n1215), .B(n1203), .Z(G45) );
NAND4_X1 U891 ( .A1(n1216), .A2(n1189), .A3(n1217), .A4(n1218), .ZN(n1203) );
XOR2_X1 U892 ( .A(G140), .B(n1209), .Z(G42) );
AND4_X1 U893 ( .A1(n1059), .A2(n1219), .A3(n1194), .A4(n1060), .ZN(n1209) );
XOR2_X1 U894 ( .A(G137), .B(n1208), .Z(G39) );
AND2_X1 U895 ( .A1(n1219), .A2(n1196), .ZN(n1208) );
INV_X1 U896 ( .A(n1220), .ZN(n1196) );
XNOR2_X1 U897 ( .A(G134), .B(n1204), .ZN(G36) );
NAND3_X1 U898 ( .A1(n1189), .A2(n1193), .A3(n1219), .ZN(n1204) );
XNOR2_X1 U899 ( .A(n1207), .B(n1221), .ZN(G33) );
XNOR2_X1 U900 ( .A(G131), .B(KEYINPUT49), .ZN(n1221) );
AND3_X1 U901 ( .A1(n1189), .A2(n1194), .A3(n1219), .ZN(n1207) );
AND4_X1 U902 ( .A1(n1036), .A2(n1217), .A3(n1218), .A4(n1039), .ZN(n1219) );
XOR2_X1 U903 ( .A(G128), .B(n1222), .Z(G30) );
NOR2_X1 U904 ( .A1(n1213), .A2(n1223), .ZN(n1222) );
XOR2_X1 U905 ( .A(KEYINPUT8), .B(n1193), .Z(n1223) );
NAND3_X1 U906 ( .A1(n1224), .A2(n1217), .A3(n1225), .ZN(n1213) );
XNOR2_X1 U907 ( .A(G101), .B(n1198), .ZN(G3) );
NAND3_X1 U908 ( .A1(n1189), .A2(n1201), .A3(n1042), .ZN(n1198) );
XOR2_X1 U909 ( .A(n1106), .B(n1211), .Z(G27) );
NAND4_X1 U910 ( .A1(n1225), .A2(n1048), .A3(n1194), .A4(n1060), .ZN(n1211) );
AND3_X1 U911 ( .A1(n1061), .A2(n1218), .A3(n1059), .ZN(n1225) );
NAND2_X1 U912 ( .A1(n1062), .A2(n1226), .ZN(n1218) );
NAND3_X1 U913 ( .A1(n1227), .A2(n1228), .A3(n1095), .ZN(n1226) );
NOR2_X1 U914 ( .A1(n1026), .A2(G900), .ZN(n1095) );
NAND2_X1 U915 ( .A1(n1229), .A2(n1230), .ZN(G24) );
NAND2_X1 U916 ( .A1(n1231), .A2(n1183), .ZN(n1230) );
XOR2_X1 U917 ( .A(n1232), .B(KEYINPUT37), .Z(n1229) );
OR2_X1 U918 ( .A1(n1183), .A2(n1231), .ZN(n1232) );
XNOR2_X1 U919 ( .A(G122), .B(KEYINPUT38), .ZN(n1231) );
NAND3_X1 U920 ( .A1(n1185), .A2(n1037), .A3(n1216), .ZN(n1183) );
AND3_X1 U921 ( .A1(n1233), .A2(n1234), .A3(n1061), .ZN(n1216) );
NOR2_X1 U922 ( .A1(n1224), .A2(n1059), .ZN(n1037) );
XOR2_X1 U923 ( .A(G119), .B(n1235), .Z(G21) );
NOR4_X1 U924 ( .A1(KEYINPUT63), .A2(n1236), .A3(n1220), .A4(n1237), .ZN(n1235) );
NAND3_X1 U925 ( .A1(n1224), .A2(n1059), .A3(n1042), .ZN(n1220) );
INV_X1 U926 ( .A(n1061), .ZN(n1236) );
XOR2_X1 U927 ( .A(G116), .B(n1238), .Z(G18) );
NOR3_X1 U928 ( .A1(n1239), .A2(n1058), .A3(n1240), .ZN(n1238) );
XOR2_X1 U929 ( .A(KEYINPUT44), .B(n1048), .Z(n1240) );
INV_X1 U930 ( .A(n1189), .ZN(n1058) );
NAND3_X1 U931 ( .A1(n1193), .A2(n1241), .A3(n1061), .ZN(n1239) );
XNOR2_X1 U932 ( .A(n1195), .B(KEYINPUT42), .ZN(n1061) );
NOR2_X1 U933 ( .A1(n1233), .A2(n1242), .ZN(n1193) );
XNOR2_X1 U934 ( .A(G113), .B(n1243), .ZN(G15) );
NAND4_X1 U935 ( .A1(n1185), .A2(n1189), .A3(n1195), .A4(n1244), .ZN(n1243) );
XOR2_X1 U936 ( .A(KEYINPUT9), .B(n1194), .Z(n1244) );
INV_X1 U937 ( .A(n1157), .ZN(n1194) );
NAND2_X1 U938 ( .A1(n1242), .A2(n1233), .ZN(n1157) );
NOR2_X1 U939 ( .A1(n1060), .A2(n1059), .ZN(n1189) );
INV_X1 U940 ( .A(n1237), .ZN(n1185) );
NAND2_X1 U941 ( .A1(n1048), .A2(n1241), .ZN(n1237) );
NOR2_X1 U942 ( .A1(n1047), .A2(n1245), .ZN(n1048) );
INV_X1 U943 ( .A(n1046), .ZN(n1245) );
XNOR2_X1 U944 ( .A(G110), .B(n1199), .ZN(G12) );
NAND4_X1 U945 ( .A1(n1059), .A2(n1042), .A3(n1201), .A4(n1060), .ZN(n1199) );
INV_X1 U946 ( .A(n1224), .ZN(n1060) );
XOR2_X1 U947 ( .A(n1063), .B(KEYINPUT59), .Z(n1224) );
XOR2_X1 U948 ( .A(n1246), .B(G472), .Z(n1063) );
NAND2_X1 U949 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
XNOR2_X1 U950 ( .A(n1170), .B(n1249), .ZN(n1247) );
XOR2_X1 U951 ( .A(G101), .B(n1250), .Z(n1249) );
NOR3_X1 U952 ( .A1(KEYINPUT13), .A2(n1251), .A3(n1252), .ZN(n1250) );
NOR2_X1 U953 ( .A1(n1169), .A2(n1253), .ZN(n1252) );
INV_X1 U954 ( .A(KEYINPUT12), .ZN(n1253) );
XOR2_X1 U955 ( .A(n1254), .B(n1255), .Z(n1169) );
NOR2_X1 U956 ( .A1(KEYINPUT12), .A2(n1256), .ZN(n1251) );
NOR2_X1 U957 ( .A1(n1255), .A2(n1254), .ZN(n1256) );
XOR2_X1 U958 ( .A(n1257), .B(n1258), .Z(n1254) );
NOR2_X1 U959 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U960 ( .A(n1261), .B(KEYINPUT23), .Z(n1260) );
NAND2_X1 U961 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NOR2_X1 U962 ( .A1(n1263), .A2(n1262), .ZN(n1259) );
XOR2_X1 U963 ( .A(KEYINPUT60), .B(G116), .Z(n1262) );
INV_X1 U964 ( .A(G119), .ZN(n1263) );
XNOR2_X1 U965 ( .A(n1264), .B(n1215), .ZN(n1255) );
NAND2_X1 U966 ( .A1(G210), .A2(n1265), .ZN(n1170) );
AND3_X1 U967 ( .A1(n1195), .A2(n1241), .A3(n1217), .ZN(n1201) );
INV_X1 U968 ( .A(n1044), .ZN(n1217) );
NAND2_X1 U969 ( .A1(n1047), .A2(n1046), .ZN(n1044) );
NAND2_X1 U970 ( .A1(G221), .A2(n1266), .ZN(n1046) );
XNOR2_X1 U971 ( .A(n1087), .B(G469), .ZN(n1047) );
NAND2_X1 U972 ( .A1(n1267), .A2(n1248), .ZN(n1087) );
XOR2_X1 U973 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U974 ( .A(n1270), .B(n1271), .Z(n1269) );
XNOR2_X1 U975 ( .A(KEYINPUT31), .B(KEYINPUT30), .ZN(n1271) );
NAND2_X1 U976 ( .A1(KEYINPUT29), .A2(G110), .ZN(n1270) );
XOR2_X1 U977 ( .A(n1272), .B(n1273), .Z(n1268) );
INV_X1 U978 ( .A(n1176), .ZN(n1273) );
XOR2_X1 U979 ( .A(n1274), .B(n1275), .Z(n1176) );
XNOR2_X1 U980 ( .A(n1110), .B(n1276), .ZN(n1275) );
XOR2_X1 U981 ( .A(KEYINPUT53), .B(G140), .Z(n1276) );
NAND2_X1 U982 ( .A1(KEYINPUT21), .A2(n1215), .ZN(n1110) );
INV_X1 U983 ( .A(G143), .ZN(n1215) );
XNOR2_X1 U984 ( .A(n1277), .B(n1264), .ZN(n1274) );
XOR2_X1 U985 ( .A(n1278), .B(n1279), .Z(n1264) );
XNOR2_X1 U986 ( .A(n1280), .B(KEYINPUT20), .ZN(n1279) );
NAND2_X1 U987 ( .A1(n1281), .A2(KEYINPUT6), .ZN(n1280) );
XNOR2_X1 U988 ( .A(G134), .B(n1282), .ZN(n1281) );
NOR2_X1 U989 ( .A1(KEYINPUT10), .A2(n1105), .ZN(n1282) );
XNOR2_X1 U990 ( .A(n1109), .B(n1111), .ZN(n1278) );
XOR2_X1 U991 ( .A(G131), .B(KEYINPUT32), .Z(n1109) );
NAND2_X1 U992 ( .A1(G227), .A2(n1026), .ZN(n1277) );
NAND2_X1 U993 ( .A1(KEYINPUT56), .A2(n1177), .ZN(n1272) );
XOR2_X1 U994 ( .A(G101), .B(n1283), .Z(n1177) );
NAND2_X1 U995 ( .A1(n1284), .A2(n1062), .ZN(n1241) );
NAND3_X1 U996 ( .A1(n1228), .A2(n1026), .A3(G952), .ZN(n1062) );
NAND3_X1 U997 ( .A1(n1227), .A2(n1228), .A3(n1127), .ZN(n1284) );
NOR2_X1 U998 ( .A1(n1026), .A2(G898), .ZN(n1127) );
NAND2_X1 U999 ( .A1(G237), .A2(n1285), .ZN(n1228) );
XOR2_X1 U1000 ( .A(G902), .B(KEYINPUT43), .Z(n1227) );
AND2_X1 U1001 ( .A1(n1286), .A2(n1077), .ZN(n1195) );
INV_X1 U1002 ( .A(n1036), .ZN(n1077) );
XOR2_X1 U1003 ( .A(n1287), .B(n1181), .Z(n1036) );
AND2_X1 U1004 ( .A1(G210), .A2(n1288), .ZN(n1181) );
NAND2_X1 U1005 ( .A1(n1180), .A2(n1248), .ZN(n1287) );
XOR2_X1 U1006 ( .A(n1289), .B(n1290), .Z(n1180) );
XNOR2_X1 U1007 ( .A(n1111), .B(n1291), .ZN(n1290) );
XOR2_X1 U1008 ( .A(n1129), .B(n1292), .Z(n1291) );
NOR2_X1 U1009 ( .A1(G953), .A2(n1140), .ZN(n1292) );
INV_X1 U1010 ( .A(G224), .ZN(n1140) );
NAND2_X1 U1011 ( .A1(n1293), .A2(n1294), .ZN(n1129) );
OR2_X1 U1012 ( .A1(n1295), .A2(G110), .ZN(n1294) );
XOR2_X1 U1013 ( .A(n1296), .B(KEYINPUT52), .Z(n1293) );
NAND2_X1 U1014 ( .A1(G110), .A2(n1295), .ZN(n1296) );
XOR2_X1 U1015 ( .A(G146), .B(G128), .Z(n1111) );
XOR2_X1 U1016 ( .A(n1297), .B(n1138), .Z(n1289) );
XNOR2_X1 U1017 ( .A(n1298), .B(n1283), .ZN(n1138) );
XNOR2_X1 U1018 ( .A(G104), .B(n1024), .ZN(n1283) );
INV_X1 U1019 ( .A(G107), .ZN(n1024) );
NAND2_X1 U1020 ( .A1(KEYINPUT34), .A2(G101), .ZN(n1298) );
XNOR2_X1 U1021 ( .A(n1299), .B(n1135), .ZN(n1297) );
XNOR2_X1 U1022 ( .A(n1300), .B(n1301), .ZN(n1135) );
INV_X1 U1023 ( .A(n1257), .ZN(n1301) );
XNOR2_X1 U1024 ( .A(G113), .B(KEYINPUT50), .ZN(n1257) );
XOR2_X1 U1025 ( .A(n1302), .B(G119), .Z(n1300) );
INV_X1 U1026 ( .A(G116), .ZN(n1302) );
XOR2_X1 U1027 ( .A(n1039), .B(KEYINPUT45), .Z(n1286) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1303), .ZN(n1039) );
XNOR2_X1 U1029 ( .A(KEYINPUT36), .B(n1288), .ZN(n1303) );
OR2_X1 U1030 ( .A1(G902), .A2(G237), .ZN(n1288) );
NOR2_X1 U1031 ( .A1(n1234), .A2(n1233), .ZN(n1042) );
XNOR2_X1 U1032 ( .A(n1073), .B(G475), .ZN(n1233) );
NAND2_X1 U1033 ( .A1(n1304), .A2(n1248), .ZN(n1073) );
XNOR2_X1 U1034 ( .A(n1154), .B(KEYINPUT58), .ZN(n1304) );
XNOR2_X1 U1035 ( .A(n1305), .B(G131), .ZN(n1154) );
XOR2_X1 U1036 ( .A(n1306), .B(n1307), .Z(n1305) );
XOR2_X1 U1037 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1038 ( .A(G113), .B(G104), .Z(n1309) );
XOR2_X1 U1039 ( .A(KEYINPUT46), .B(KEYINPUT11), .Z(n1308) );
XOR2_X1 U1040 ( .A(n1310), .B(n1311), .Z(n1306) );
XOR2_X1 U1041 ( .A(n1312), .B(n1313), .Z(n1311) );
NAND2_X1 U1042 ( .A1(KEYINPUT26), .A2(n1295), .ZN(n1313) );
INV_X1 U1043 ( .A(G122), .ZN(n1295) );
NAND2_X1 U1044 ( .A1(G214), .A2(n1265), .ZN(n1312) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1265) );
XOR2_X1 U1046 ( .A(n1314), .B(n1299), .Z(n1310) );
XNOR2_X1 U1047 ( .A(n1106), .B(G143), .ZN(n1299) );
INV_X1 U1048 ( .A(G125), .ZN(n1106) );
INV_X1 U1049 ( .A(n1242), .ZN(n1234) );
NOR2_X1 U1050 ( .A1(n1088), .A2(n1315), .ZN(n1242) );
AND2_X1 U1051 ( .A1(G478), .A2(n1076), .ZN(n1315) );
NOR2_X1 U1052 ( .A1(n1076), .A2(G478), .ZN(n1088) );
NAND2_X1 U1053 ( .A1(n1150), .A2(n1248), .ZN(n1076) );
XNOR2_X1 U1054 ( .A(n1316), .B(n1317), .ZN(n1150) );
XOR2_X1 U1055 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1056 ( .A(G128), .B(G122), .Z(n1319) );
XOR2_X1 U1057 ( .A(G143), .B(G134), .Z(n1318) );
XOR2_X1 U1058 ( .A(n1320), .B(n1321), .Z(n1316) );
XOR2_X1 U1059 ( .A(G116), .B(G107), .Z(n1321) );
NAND2_X1 U1060 ( .A1(G217), .A2(n1322), .ZN(n1320) );
XOR2_X1 U1061 ( .A(n1070), .B(n1323), .Z(n1059) );
NOR2_X1 U1062 ( .A1(n1072), .A2(KEYINPUT17), .ZN(n1323) );
INV_X1 U1063 ( .A(n1146), .ZN(n1072) );
NAND2_X1 U1064 ( .A1(G217), .A2(n1266), .ZN(n1146) );
NAND2_X1 U1065 ( .A1(n1324), .A2(n1285), .ZN(n1266) );
XOR2_X1 U1066 ( .A(G234), .B(KEYINPUT2), .Z(n1285) );
XOR2_X1 U1067 ( .A(KEYINPUT62), .B(G902), .Z(n1324) );
NAND2_X1 U1068 ( .A1(n1248), .A2(n1147), .ZN(n1070) );
NAND2_X1 U1069 ( .A1(n1325), .A2(n1326), .ZN(n1147) );
OR2_X1 U1070 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
XOR2_X1 U1071 ( .A(n1329), .B(KEYINPUT39), .Z(n1325) );
NAND2_X1 U1072 ( .A1(n1328), .A2(n1327), .ZN(n1329) );
XNOR2_X1 U1073 ( .A(n1330), .B(n1331), .ZN(n1327) );
NOR2_X1 U1074 ( .A1(KEYINPUT35), .A2(n1105), .ZN(n1331) );
XOR2_X1 U1075 ( .A(G137), .B(KEYINPUT28), .Z(n1105) );
NAND2_X1 U1076 ( .A1(G221), .A2(n1322), .ZN(n1330) );
AND2_X1 U1077 ( .A1(G234), .A2(n1026), .ZN(n1322) );
INV_X1 U1078 ( .A(G953), .ZN(n1026) );
XNOR2_X1 U1079 ( .A(n1314), .B(n1332), .ZN(n1328) );
XOR2_X1 U1080 ( .A(G125), .B(n1333), .Z(n1332) );
NOR2_X1 U1081 ( .A1(KEYINPUT7), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1082 ( .A(n1335), .B(n1336), .Z(n1334) );
XOR2_X1 U1083 ( .A(G119), .B(G110), .Z(n1336) );
NAND2_X1 U1084 ( .A1(KEYINPUT18), .A2(G128), .ZN(n1335) );
XNOR2_X1 U1085 ( .A(G146), .B(G140), .ZN(n1314) );
INV_X1 U1086 ( .A(G902), .ZN(n1248) );
endmodule


