//Key = 0111110011011001011101000011111101010100111001000010110111011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368;

NAND2_X1 U756 ( .A1(n1043), .A2(n1044), .ZN(G9) );
NAND3_X1 U757 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
XNOR2_X1 U758 ( .A(n1048), .B(KEYINPUT41), .ZN(n1047) );
NAND2_X1 U759 ( .A1(n1049), .A2(n1050), .ZN(n1043) );
NAND2_X1 U760 ( .A1(n1045), .A2(n1046), .ZN(n1050) );
XNOR2_X1 U761 ( .A(KEYINPUT24), .B(n1051), .ZN(n1046) );
XNOR2_X1 U762 ( .A(KEYINPUT18), .B(n1052), .ZN(n1049) );
INV_X1 U763 ( .A(n1048), .ZN(n1052) );
XOR2_X1 U764 ( .A(G107), .B(KEYINPUT56), .Z(n1048) );
NOR2_X1 U765 ( .A1(n1053), .A2(n1054), .ZN(G75) );
NOR3_X1 U766 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NAND3_X1 U767 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1055) );
NAND2_X1 U768 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U769 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND4_X1 U770 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
NAND2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND3_X1 U772 ( .A1(n1071), .A2(n1072), .A3(KEYINPUT6), .ZN(n1069) );
NAND3_X1 U773 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1067) );
NAND2_X1 U774 ( .A1(n1071), .A2(n1076), .ZN(n1074) );
NAND2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
OR2_X1 U776 ( .A1(n1079), .A2(KEYINPUT6), .ZN(n1078) );
NAND2_X1 U777 ( .A1(n1080), .A2(n1081), .ZN(n1073) );
NAND2_X1 U778 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND3_X1 U779 ( .A1(G221), .A2(n1084), .A3(n1085), .ZN(n1083) );
NAND3_X1 U780 ( .A1(n1071), .A2(n1086), .A3(n1080), .ZN(n1063) );
NAND2_X1 U781 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND3_X1 U782 ( .A1(n1089), .A2(n1090), .A3(n1065), .ZN(n1088) );
NAND2_X1 U783 ( .A1(n1091), .A2(n1070), .ZN(n1090) );
OR3_X1 U784 ( .A1(n1092), .A2(n1093), .A3(n1091), .ZN(n1089) );
NAND2_X1 U785 ( .A1(n1045), .A2(n1075), .ZN(n1087) );
INV_X1 U786 ( .A(n1094), .ZN(n1061) );
AND3_X1 U787 ( .A1(n1058), .A2(n1059), .A3(n1095), .ZN(n1053) );
NAND4_X1 U788 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1058) );
NOR4_X1 U789 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
XNOR2_X1 U790 ( .A(KEYINPUT62), .B(n1104), .ZN(n1103) );
XOR2_X1 U791 ( .A(n1105), .B(n1106), .Z(n1100) );
XOR2_X1 U792 ( .A(KEYINPUT51), .B(KEYINPUT25), .Z(n1106) );
XOR2_X1 U793 ( .A(n1107), .B(G472), .Z(n1105) );
NAND2_X1 U794 ( .A1(KEYINPUT1), .A2(n1108), .ZN(n1107) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1091), .ZN(n1098) );
NAND2_X1 U796 ( .A1(G475), .A2(n1110), .ZN(n1097) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1096) );
NAND2_X1 U798 ( .A1(KEYINPUT60), .A2(n1113), .ZN(n1112) );
XOR2_X1 U799 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U800 ( .A1(KEYINPUT22), .A2(n1116), .ZN(n1115) );
NOR2_X1 U801 ( .A1(n1117), .A2(n1059), .ZN(n1116) );
AND2_X1 U802 ( .A1(G227), .A2(G900), .ZN(n1117) );
NOR2_X1 U803 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
NOR2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1118) );
XNOR2_X1 U806 ( .A(KEYINPUT58), .B(n1121), .ZN(n1123) );
NAND2_X1 U807 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
NAND2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U809 ( .A(n1128), .B(n1129), .Z(n1124) );
XOR2_X1 U810 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR3_X1 U811 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR2_X1 U812 ( .A1(KEYINPUT29), .A2(n1135), .ZN(n1134) );
NOR3_X1 U813 ( .A1(n1136), .A2(G131), .A3(n1137), .ZN(n1133) );
INV_X1 U814 ( .A(KEYINPUT29), .ZN(n1136) );
AND2_X1 U815 ( .A1(n1137), .A2(G131), .ZN(n1132) );
NAND2_X1 U816 ( .A1(KEYINPUT52), .A2(n1135), .ZN(n1137) );
XNOR2_X1 U817 ( .A(G125), .B(G140), .ZN(n1128) );
XNOR2_X1 U818 ( .A(n1120), .B(KEYINPUT10), .ZN(n1122) );
AND2_X1 U819 ( .A1(n1138), .A2(n1057), .ZN(n1120) );
XNOR2_X1 U820 ( .A(KEYINPUT59), .B(n1059), .ZN(n1138) );
XOR2_X1 U821 ( .A(n1139), .B(n1140), .Z(G69) );
NOR2_X1 U822 ( .A1(n1141), .A2(n1059), .ZN(n1140) );
NOR2_X1 U823 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U824 ( .A1(n1144), .A2(n1145), .ZN(n1139) );
NAND3_X1 U825 ( .A1(n1056), .A2(n1059), .A3(n1146), .ZN(n1145) );
NAND2_X1 U826 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U827 ( .A1(KEYINPUT46), .A2(n1143), .ZN(n1148) );
XOR2_X1 U828 ( .A(n1149), .B(KEYINPUT7), .Z(n1144) );
NAND3_X1 U829 ( .A1(n1147), .A2(n1150), .A3(n1151), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1056), .B(KEYINPUT30), .Z(n1151) );
NAND2_X1 U831 ( .A1(n1126), .A2(n1143), .ZN(n1150) );
XNOR2_X1 U832 ( .A(n1152), .B(n1153), .ZN(n1147) );
NOR2_X1 U833 ( .A1(KEYINPUT38), .A2(n1154), .ZN(n1153) );
NOR2_X1 U834 ( .A1(n1155), .A2(n1156), .ZN(G66) );
XOR2_X1 U835 ( .A(n1157), .B(n1158), .Z(n1156) );
NAND2_X1 U836 ( .A1(KEYINPUT50), .A2(n1159), .ZN(n1158) );
NAND2_X1 U837 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1155), .A2(n1162), .ZN(G63) );
XOR2_X1 U839 ( .A(n1163), .B(n1164), .Z(n1162) );
AND2_X1 U840 ( .A1(G478), .A2(n1160), .ZN(n1163) );
NOR2_X1 U841 ( .A1(n1155), .A2(n1165), .ZN(G60) );
XNOR2_X1 U842 ( .A(n1166), .B(n1167), .ZN(n1165) );
AND2_X1 U843 ( .A1(G475), .A2(n1160), .ZN(n1167) );
XNOR2_X1 U844 ( .A(G104), .B(n1168), .ZN(G6) );
NAND4_X1 U845 ( .A1(n1169), .A2(n1170), .A3(n1075), .A4(n1171), .ZN(n1168) );
NOR2_X1 U846 ( .A1(n1155), .A2(n1172), .ZN(G57) );
XOR2_X1 U847 ( .A(n1173), .B(n1174), .Z(n1172) );
AND2_X1 U848 ( .A1(G472), .A2(n1160), .ZN(n1173) );
NOR2_X1 U849 ( .A1(n1155), .A2(n1175), .ZN(G54) );
XOR2_X1 U850 ( .A(n1176), .B(n1177), .Z(n1175) );
XNOR2_X1 U851 ( .A(n1178), .B(n1179), .ZN(n1177) );
XNOR2_X1 U852 ( .A(n1180), .B(n1181), .ZN(n1176) );
NOR2_X1 U853 ( .A1(n1182), .A2(KEYINPUT36), .ZN(n1181) );
NOR3_X1 U854 ( .A1(n1183), .A2(KEYINPUT39), .A3(n1184), .ZN(n1180) );
NOR3_X1 U855 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(G51) );
AND2_X1 U856 ( .A1(KEYINPUT57), .A2(n1155), .ZN(n1187) );
NOR2_X1 U857 ( .A1(n1059), .A2(G952), .ZN(n1155) );
NOR3_X1 U858 ( .A1(KEYINPUT57), .A2(n1059), .A3(n1095), .ZN(n1186) );
INV_X1 U859 ( .A(G952), .ZN(n1095) );
XOR2_X1 U860 ( .A(n1188), .B(n1189), .Z(n1185) );
NAND3_X1 U861 ( .A1(G210), .A2(n1190), .A3(n1160), .ZN(n1189) );
INV_X1 U862 ( .A(n1183), .ZN(n1160) );
NAND2_X1 U863 ( .A1(G902), .A2(n1191), .ZN(n1183) );
OR2_X1 U864 ( .A1(n1057), .A2(n1056), .ZN(n1191) );
NAND4_X1 U865 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1056) );
NOR3_X1 U866 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1195) );
NOR2_X1 U867 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
INV_X1 U868 ( .A(n1201), .ZN(n1200) );
NOR2_X1 U869 ( .A1(n1202), .A2(n1203), .ZN(n1199) );
AND2_X1 U870 ( .A1(n1075), .A2(n1204), .ZN(n1202) );
NOR2_X1 U871 ( .A1(n1051), .A2(n1205), .ZN(n1197) );
XNOR2_X1 U872 ( .A(KEYINPUT33), .B(n1206), .ZN(n1205) );
NAND4_X1 U873 ( .A1(n1207), .A2(n1075), .A3(n1072), .A4(n1171), .ZN(n1051) );
NOR2_X1 U874 ( .A1(n1208), .A2(n1209), .ZN(n1196) );
NOR2_X1 U875 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
AND3_X1 U876 ( .A1(n1080), .A2(n1093), .A3(n1169), .ZN(n1211) );
NOR4_X1 U877 ( .A1(n1212), .A2(n1213), .A3(n1070), .A4(n1077), .ZN(n1210) );
INV_X1 U878 ( .A(n1075), .ZN(n1070) );
NOR2_X1 U879 ( .A1(KEYINPUT9), .A2(n1214), .ZN(n1213) );
NOR2_X1 U880 ( .A1(n1045), .A2(n1082), .ZN(n1214) );
NOR2_X1 U881 ( .A1(n1169), .A2(n1215), .ZN(n1212) );
INV_X1 U882 ( .A(KEYINPUT9), .ZN(n1215) );
NAND4_X1 U883 ( .A1(n1216), .A2(n1217), .A3(n1218), .A4(n1219), .ZN(n1057) );
NOR4_X1 U884 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1219) );
NOR3_X1 U885 ( .A1(n1224), .A2(n1225), .A3(n1226), .ZN(n1223) );
NOR2_X1 U886 ( .A1(KEYINPUT2), .A2(n1227), .ZN(n1226) );
NOR4_X1 U887 ( .A1(n1091), .A2(n1228), .A3(n1082), .A4(n1229), .ZN(n1227) );
INV_X1 U888 ( .A(n1065), .ZN(n1228) );
AND2_X1 U889 ( .A1(n1230), .A2(KEYINPUT2), .ZN(n1225) );
OR2_X1 U890 ( .A1(n1231), .A2(n1232), .ZN(n1218) );
NAND2_X1 U891 ( .A1(n1072), .A2(n1233), .ZN(n1217) );
NAND2_X1 U892 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U893 ( .A1(n1236), .A2(n1092), .ZN(n1235) );
NAND2_X1 U894 ( .A1(n1170), .A2(n1237), .ZN(n1216) );
NAND2_X1 U895 ( .A1(n1234), .A2(n1238), .ZN(n1237) );
NAND4_X1 U896 ( .A1(n1206), .A2(n1231), .A3(n1229), .A4(n1239), .ZN(n1238) );
NOR2_X1 U897 ( .A1(n1102), .A2(n1240), .ZN(n1239) );
INV_X1 U898 ( .A(KEYINPUT3), .ZN(n1231) );
NAND2_X1 U899 ( .A1(KEYINPUT26), .A2(n1241), .ZN(n1188) );
XOR2_X1 U900 ( .A(G146), .B(n1242), .Z(G48) );
NOR2_X1 U901 ( .A1(n1077), .A2(n1234), .ZN(n1242) );
XOR2_X1 U902 ( .A(G143), .B(n1222), .Z(G45) );
AND4_X1 U903 ( .A1(n1169), .A2(n1204), .A3(n1092), .A4(n1229), .ZN(n1222) );
XOR2_X1 U904 ( .A(G140), .B(n1221), .Z(G42) );
NOR3_X1 U905 ( .A1(n1077), .A2(n1230), .A3(n1240), .ZN(n1221) );
INV_X1 U906 ( .A(n1170), .ZN(n1077) );
XOR2_X1 U907 ( .A(G137), .B(n1243), .Z(G39) );
NOR2_X1 U908 ( .A1(n1230), .A2(n1224), .ZN(n1243) );
XNOR2_X1 U909 ( .A(G134), .B(n1244), .ZN(G36) );
NAND4_X1 U910 ( .A1(KEYINPUT35), .A2(n1236), .A3(n1072), .A4(n1092), .ZN(n1244) );
XOR2_X1 U911 ( .A(G131), .B(n1220), .Z(G33) );
AND3_X1 U912 ( .A1(n1236), .A2(n1092), .A3(n1170), .ZN(n1220) );
INV_X1 U913 ( .A(n1230), .ZN(n1236) );
NAND4_X1 U914 ( .A1(n1207), .A2(n1065), .A3(n1229), .A4(n1066), .ZN(n1230) );
XNOR2_X1 U915 ( .A(n1245), .B(n1246), .ZN(G30) );
NOR2_X1 U916 ( .A1(n1079), .A2(n1234), .ZN(n1246) );
NAND3_X1 U917 ( .A1(n1169), .A2(n1229), .A3(n1247), .ZN(n1234) );
XNOR2_X1 U918 ( .A(G101), .B(n1194), .ZN(G3) );
NAND4_X1 U919 ( .A1(n1080), .A2(n1169), .A3(n1092), .A4(n1171), .ZN(n1194) );
XNOR2_X1 U920 ( .A(G125), .B(n1232), .ZN(G27) );
NAND4_X1 U921 ( .A1(n1093), .A2(n1170), .A3(n1248), .A4(n1071), .ZN(n1232) );
INV_X1 U922 ( .A(n1102), .ZN(n1071) );
AND2_X1 U923 ( .A1(n1229), .A2(n1045), .ZN(n1248) );
NAND2_X1 U924 ( .A1(n1094), .A2(n1249), .ZN(n1229) );
NAND4_X1 U925 ( .A1(G902), .A2(n1126), .A3(n1250), .A4(n1127), .ZN(n1249) );
INV_X1 U926 ( .A(G900), .ZN(n1127) );
XNOR2_X1 U927 ( .A(G122), .B(n1251), .ZN(G24) );
NAND3_X1 U928 ( .A1(n1201), .A2(n1075), .A3(n1252), .ZN(n1251) );
XNOR2_X1 U929 ( .A(n1204), .B(KEYINPUT17), .ZN(n1252) );
NOR2_X1 U930 ( .A1(n1104), .A2(n1253), .ZN(n1204) );
XNOR2_X1 U931 ( .A(G119), .B(n1254), .ZN(G21) );
NAND2_X1 U932 ( .A1(n1201), .A2(n1203), .ZN(n1254) );
INV_X1 U933 ( .A(n1224), .ZN(n1203) );
NAND2_X1 U934 ( .A1(n1080), .A2(n1247), .ZN(n1224) );
AND2_X1 U935 ( .A1(n1255), .A2(n1101), .ZN(n1247) );
XNOR2_X1 U936 ( .A(n1256), .B(n1257), .ZN(n1255) );
XNOR2_X1 U937 ( .A(G116), .B(n1192), .ZN(G18) );
NAND3_X1 U938 ( .A1(n1072), .A2(n1092), .A3(n1201), .ZN(n1192) );
INV_X1 U939 ( .A(n1079), .ZN(n1072) );
NAND2_X1 U940 ( .A1(n1253), .A2(n1258), .ZN(n1079) );
XNOR2_X1 U941 ( .A(G113), .B(n1193), .ZN(G15) );
NAND3_X1 U942 ( .A1(n1170), .A2(n1092), .A3(n1201), .ZN(n1193) );
NOR3_X1 U943 ( .A1(n1206), .A2(n1208), .A3(n1102), .ZN(n1201) );
NAND2_X1 U944 ( .A1(n1085), .A2(n1259), .ZN(n1102) );
NAND2_X1 U945 ( .A1(G221), .A2(n1084), .ZN(n1259) );
NAND2_X1 U946 ( .A1(n1260), .A2(n1261), .ZN(n1092) );
NAND2_X1 U947 ( .A1(n1075), .A2(n1256), .ZN(n1261) );
NOR2_X1 U948 ( .A1(n1101), .A2(n1262), .ZN(n1075) );
INV_X1 U949 ( .A(n1257), .ZN(n1262) );
OR3_X1 U950 ( .A1(n1101), .A2(n1257), .A3(n1256), .ZN(n1260) );
INV_X1 U951 ( .A(KEYINPUT53), .ZN(n1256) );
NOR2_X1 U952 ( .A1(n1258), .A2(n1253), .ZN(n1170) );
XNOR2_X1 U953 ( .A(G110), .B(n1263), .ZN(G12) );
NAND4_X1 U954 ( .A1(n1264), .A2(n1080), .A3(n1169), .A4(n1093), .ZN(n1263) );
INV_X1 U955 ( .A(n1240), .ZN(n1093) );
NAND2_X1 U956 ( .A1(n1257), .A2(n1101), .ZN(n1240) );
XNOR2_X1 U957 ( .A(n1265), .B(n1161), .ZN(n1101) );
AND2_X1 U958 ( .A1(G217), .A2(n1084), .ZN(n1161) );
OR2_X1 U959 ( .A1(n1159), .A2(G902), .ZN(n1265) );
XOR2_X1 U960 ( .A(n1266), .B(n1267), .Z(n1159) );
XOR2_X1 U961 ( .A(G137), .B(n1268), .Z(n1267) );
AND3_X1 U962 ( .A1(G221), .A2(n1059), .A3(G234), .ZN(n1268) );
NAND3_X1 U963 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1266) );
OR2_X1 U964 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND3_X1 U965 ( .A1(n1273), .A2(n1272), .A3(KEYINPUT40), .ZN(n1270) );
XNOR2_X1 U966 ( .A(n1274), .B(n1275), .ZN(n1272) );
XOR2_X1 U967 ( .A(KEYINPUT55), .B(G146), .Z(n1275) );
NAND2_X1 U968 ( .A1(n1276), .A2(n1277), .ZN(n1274) );
NAND2_X1 U969 ( .A1(G140), .A2(n1278), .ZN(n1277) );
XOR2_X1 U970 ( .A(KEYINPUT12), .B(n1279), .Z(n1276) );
NOR2_X1 U971 ( .A1(G140), .A2(n1278), .ZN(n1279) );
AND2_X1 U972 ( .A1(KEYINPUT28), .A2(n1280), .ZN(n1273) );
OR2_X1 U973 ( .A1(n1280), .A2(KEYINPUT40), .ZN(n1269) );
XOR2_X1 U974 ( .A(n1281), .B(n1282), .Z(n1280) );
XNOR2_X1 U975 ( .A(KEYINPUT5), .B(n1245), .ZN(n1282) );
XNOR2_X1 U976 ( .A(G110), .B(G119), .ZN(n1281) );
XNOR2_X1 U977 ( .A(n1283), .B(G472), .ZN(n1257) );
NAND2_X1 U978 ( .A1(KEYINPUT45), .A2(n1108), .ZN(n1283) );
OR2_X1 U979 ( .A1(n1174), .A2(G902), .ZN(n1108) );
XNOR2_X1 U980 ( .A(n1284), .B(n1285), .ZN(n1174) );
XOR2_X1 U981 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U982 ( .A(G101), .B(n1288), .ZN(n1287) );
AND3_X1 U983 ( .A1(G210), .A2(n1059), .A3(n1289), .ZN(n1288) );
NAND2_X1 U984 ( .A1(n1290), .A2(n1291), .ZN(n1286) );
NAND2_X1 U985 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U986 ( .A(KEYINPUT16), .B(n1294), .ZN(n1292) );
XOR2_X1 U987 ( .A(n1295), .B(KEYINPUT23), .Z(n1290) );
OR2_X1 U988 ( .A1(n1293), .A2(G113), .ZN(n1295) );
XNOR2_X1 U989 ( .A(G116), .B(n1296), .ZN(n1293) );
INV_X1 U990 ( .A(G119), .ZN(n1296) );
XNOR2_X1 U991 ( .A(n1178), .B(n1297), .ZN(n1284) );
NOR2_X1 U992 ( .A1(n1206), .A2(n1082), .ZN(n1169) );
INV_X1 U993 ( .A(n1207), .ZN(n1082) );
NOR2_X1 U994 ( .A1(n1085), .A2(n1298), .ZN(n1207) );
AND2_X1 U995 ( .A1(G221), .A2(n1084), .ZN(n1298) );
NAND2_X1 U996 ( .A1(G234), .A2(n1299), .ZN(n1084) );
XNOR2_X1 U997 ( .A(n1300), .B(n1184), .ZN(n1085) );
INV_X1 U998 ( .A(G469), .ZN(n1184) );
NAND2_X1 U999 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XNOR2_X1 U1000 ( .A(n1179), .B(n1303), .ZN(n1301) );
XOR2_X1 U1001 ( .A(n1182), .B(n1304), .Z(n1303) );
NOR2_X1 U1002 ( .A1(KEYINPUT13), .A2(n1178), .ZN(n1304) );
XNOR2_X1 U1003 ( .A(n1305), .B(KEYINPUT61), .ZN(n1178) );
NAND2_X1 U1004 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1005 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
INV_X1 U1006 ( .A(n1310), .ZN(n1309) );
NAND2_X1 U1007 ( .A1(n1311), .A2(n1310), .ZN(n1306) );
XOR2_X1 U1008 ( .A(G131), .B(KEYINPUT37), .Z(n1310) );
XOR2_X1 U1009 ( .A(n1308), .B(n1312), .Z(n1311) );
XOR2_X1 U1010 ( .A(KEYINPUT49), .B(KEYINPUT4), .Z(n1312) );
XOR2_X1 U1011 ( .A(n1135), .B(KEYINPUT43), .Z(n1308) );
XOR2_X1 U1012 ( .A(G134), .B(G137), .Z(n1135) );
AND2_X1 U1013 ( .A1(n1313), .A2(n1314), .ZN(n1182) );
NAND3_X1 U1014 ( .A1(G227), .A2(n1059), .A3(n1315), .ZN(n1314) );
XNOR2_X1 U1015 ( .A(G110), .B(G140), .ZN(n1315) );
NAND2_X1 U1016 ( .A1(n1316), .A2(n1317), .ZN(n1313) );
NAND2_X1 U1017 ( .A1(G227), .A2(n1059), .ZN(n1317) );
XOR2_X1 U1018 ( .A(G140), .B(G110), .Z(n1316) );
XOR2_X1 U1019 ( .A(n1318), .B(n1319), .Z(n1179) );
XOR2_X1 U1020 ( .A(n1130), .B(KEYINPUT8), .Z(n1318) );
NAND3_X1 U1021 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1130) );
NAND2_X1 U1022 ( .A1(G128), .A2(n1323), .ZN(n1322) );
NAND2_X1 U1023 ( .A1(KEYINPUT44), .A2(n1324), .ZN(n1321) );
NAND2_X1 U1024 ( .A1(n1325), .A2(n1245), .ZN(n1324) );
XNOR2_X1 U1025 ( .A(KEYINPUT42), .B(n1326), .ZN(n1325) );
NAND2_X1 U1026 ( .A1(n1327), .A2(n1328), .ZN(n1320) );
INV_X1 U1027 ( .A(KEYINPUT44), .ZN(n1328) );
NAND2_X1 U1028 ( .A1(n1329), .A2(n1330), .ZN(n1327) );
NAND3_X1 U1029 ( .A1(KEYINPUT42), .A2(n1245), .A3(n1326), .ZN(n1330) );
INV_X1 U1030 ( .A(G128), .ZN(n1245) );
OR2_X1 U1031 ( .A1(n1326), .A2(KEYINPUT42), .ZN(n1329) );
INV_X1 U1032 ( .A(n1045), .ZN(n1206) );
NOR2_X1 U1033 ( .A1(n1065), .A2(n1091), .ZN(n1045) );
INV_X1 U1034 ( .A(n1066), .ZN(n1091) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1190), .ZN(n1066) );
XOR2_X1 U1036 ( .A(n1331), .B(n1113), .Z(n1065) );
NAND2_X1 U1037 ( .A1(n1332), .A2(G210), .ZN(n1113) );
XOR2_X1 U1038 ( .A(n1190), .B(KEYINPUT63), .Z(n1332) );
NAND2_X1 U1039 ( .A1(n1299), .A2(n1289), .ZN(n1190) );
XNOR2_X1 U1040 ( .A(G902), .B(KEYINPUT14), .ZN(n1299) );
XOR2_X1 U1041 ( .A(n1111), .B(KEYINPUT19), .Z(n1331) );
OR2_X1 U1042 ( .A1(n1241), .A2(G902), .ZN(n1111) );
XNOR2_X1 U1043 ( .A(n1333), .B(n1334), .ZN(n1241) );
XOR2_X1 U1044 ( .A(n1335), .B(n1336), .Z(n1334) );
XNOR2_X1 U1045 ( .A(n1278), .B(n1337), .ZN(n1336) );
NOR2_X1 U1046 ( .A1(KEYINPUT47), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1047 ( .A(KEYINPUT21), .B(n1152), .ZN(n1338) );
XOR2_X1 U1048 ( .A(n1339), .B(n1319), .Z(n1152) );
XOR2_X1 U1049 ( .A(G101), .B(n1340), .Z(n1319) );
XNOR2_X1 U1050 ( .A(n1341), .B(G104), .ZN(n1340) );
INV_X1 U1051 ( .A(G107), .ZN(n1341) );
XNOR2_X1 U1052 ( .A(G113), .B(n1342), .ZN(n1339) );
NOR2_X1 U1053 ( .A1(KEYINPUT54), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1054 ( .A(G116), .B(n1344), .Z(n1343) );
NOR2_X1 U1055 ( .A1(G119), .A2(KEYINPUT20), .ZN(n1344) );
NOR2_X1 U1056 ( .A1(G953), .A2(n1142), .ZN(n1335) );
INV_X1 U1057 ( .A(G224), .ZN(n1142) );
XOR2_X1 U1058 ( .A(n1154), .B(n1297), .Z(n1333) );
XNOR2_X1 U1059 ( .A(n1345), .B(n1323), .ZN(n1297) );
XNOR2_X1 U1060 ( .A(G128), .B(KEYINPUT0), .ZN(n1345) );
XOR2_X1 U1061 ( .A(n1346), .B(G110), .Z(n1154) );
NAND2_X1 U1062 ( .A1(KEYINPUT15), .A2(n1347), .ZN(n1346) );
AND2_X1 U1063 ( .A1(n1104), .A2(n1253), .ZN(n1080) );
NOR2_X1 U1064 ( .A1(n1348), .A2(n1109), .ZN(n1253) );
NOR3_X1 U1065 ( .A1(G475), .A2(G902), .A3(n1349), .ZN(n1109) );
INV_X1 U1066 ( .A(n1166), .ZN(n1349) );
AND2_X1 U1067 ( .A1(n1350), .A2(n1110), .ZN(n1348) );
NAND2_X1 U1068 ( .A1(n1166), .A2(n1302), .ZN(n1110) );
INV_X1 U1069 ( .A(G902), .ZN(n1302) );
XNOR2_X1 U1070 ( .A(n1351), .B(n1352), .ZN(n1166) );
XOR2_X1 U1071 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1072 ( .A(n1347), .B(G104), .ZN(n1354) );
XNOR2_X1 U1073 ( .A(G131), .B(n1278), .ZN(n1353) );
INV_X1 U1074 ( .A(G125), .ZN(n1278) );
XOR2_X1 U1075 ( .A(n1355), .B(n1356), .Z(n1351) );
XNOR2_X1 U1076 ( .A(n1357), .B(n1326), .ZN(n1356) );
INV_X1 U1077 ( .A(n1323), .ZN(n1326) );
XOR2_X1 U1078 ( .A(G143), .B(G146), .Z(n1323) );
NOR2_X1 U1079 ( .A1(G140), .A2(KEYINPUT34), .ZN(n1357) );
XNOR2_X1 U1080 ( .A(n1358), .B(n1359), .ZN(n1355) );
NAND2_X1 U1081 ( .A1(KEYINPUT27), .A2(n1294), .ZN(n1359) );
INV_X1 U1082 ( .A(G113), .ZN(n1294) );
NAND4_X1 U1083 ( .A1(KEYINPUT31), .A2(G214), .A3(n1289), .A4(n1059), .ZN(n1358) );
INV_X1 U1084 ( .A(G237), .ZN(n1289) );
XNOR2_X1 U1085 ( .A(G475), .B(KEYINPUT11), .ZN(n1350) );
INV_X1 U1086 ( .A(n1258), .ZN(n1104) );
XNOR2_X1 U1087 ( .A(n1360), .B(G478), .ZN(n1258) );
OR2_X1 U1088 ( .A1(n1164), .A2(G902), .ZN(n1360) );
XNOR2_X1 U1089 ( .A(n1361), .B(n1362), .ZN(n1164) );
XOR2_X1 U1090 ( .A(n1363), .B(n1364), .Z(n1362) );
XNOR2_X1 U1091 ( .A(G107), .B(n1365), .ZN(n1364) );
NOR2_X1 U1092 ( .A1(G134), .A2(KEYINPUT32), .ZN(n1365) );
NAND3_X1 U1093 ( .A1(G234), .A2(n1059), .A3(G217), .ZN(n1363) );
XOR2_X1 U1094 ( .A(n1366), .B(n1367), .Z(n1361) );
XNOR2_X1 U1095 ( .A(n1347), .B(G116), .ZN(n1367) );
INV_X1 U1096 ( .A(G122), .ZN(n1347) );
XNOR2_X1 U1097 ( .A(G143), .B(G128), .ZN(n1366) );
XNOR2_X1 U1098 ( .A(n1208), .B(KEYINPUT48), .ZN(n1264) );
INV_X1 U1099 ( .A(n1171), .ZN(n1208) );
NAND2_X1 U1100 ( .A1(n1094), .A2(n1368), .ZN(n1171) );
NAND4_X1 U1101 ( .A1(G902), .A2(n1126), .A3(n1250), .A4(n1143), .ZN(n1368) );
INV_X1 U1102 ( .A(G898), .ZN(n1143) );
XOR2_X1 U1103 ( .A(KEYINPUT46), .B(G953), .Z(n1126) );
NAND3_X1 U1104 ( .A1(n1250), .A2(n1059), .A3(G952), .ZN(n1094) );
INV_X1 U1105 ( .A(G953), .ZN(n1059) );
NAND2_X1 U1106 ( .A1(G237), .A2(G234), .ZN(n1250) );
endmodule


