//Key = 1000001011010010111001011000100010110100100101001001110001001100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318;

XNOR2_X1 U723 ( .A(G107), .B(n985), .ZN(G9) );
NAND4_X1 U724 ( .A1(n986), .A2(n987), .A3(n988), .A4(n989), .ZN(n985) );
OR2_X1 U725 ( .A1(n990), .A2(KEYINPUT20), .ZN(n989) );
NAND2_X1 U726 ( .A1(KEYINPUT20), .A2(n991), .ZN(n988) );
NAND2_X1 U727 ( .A1(n992), .A2(n993), .ZN(n991) );
NAND4_X1 U728 ( .A1(n994), .A2(n995), .A3(n996), .A4(n997), .ZN(G75) );
NAND4_X1 U729 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(n996) );
NOR4_X1 U730 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1001) );
INV_X1 U731 ( .A(n1006), .ZN(n1003) );
NAND2_X1 U732 ( .A1(n1007), .A2(n1008), .ZN(n1002) );
XNOR2_X1 U733 ( .A(n1009), .B(n1010), .ZN(n1007) );
NAND2_X1 U734 ( .A1(KEYINPUT37), .A2(n1011), .ZN(n1010) );
NOR3_X1 U735 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1000) );
NOR3_X1 U736 ( .A1(n1015), .A2(KEYINPUT38), .A3(n1016), .ZN(n1014) );
AND2_X1 U737 ( .A1(n1015), .A2(KEYINPUT38), .ZN(n1013) );
XOR2_X1 U738 ( .A(n1017), .B(n1018), .Z(n1012) );
XNOR2_X1 U739 ( .A(n1019), .B(KEYINPUT2), .ZN(n998) );
NAND2_X1 U740 ( .A1(n1020), .A2(n1021), .ZN(n995) );
NAND2_X1 U741 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND3_X1 U742 ( .A1(n987), .A2(n1024), .A3(n1025), .ZN(n1023) );
NAND2_X1 U743 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NAND2_X1 U744 ( .A1(n999), .A2(n1028), .ZN(n1027) );
NAND2_X1 U745 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND2_X1 U746 ( .A1(n1031), .A2(n1032), .ZN(n1026) );
NAND2_X1 U747 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
INV_X1 U749 ( .A(n1037), .ZN(n1033) );
NAND3_X1 U750 ( .A1(n1031), .A2(n1038), .A3(n999), .ZN(n1022) );
NAND2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U752 ( .A1(n1025), .A2(n1041), .ZN(n1040) );
NAND2_X1 U753 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U754 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U755 ( .A1(n987), .A2(n1046), .ZN(n1039) );
NAND2_X1 U756 ( .A1(n993), .A2(n1047), .ZN(n1046) );
NAND2_X1 U757 ( .A1(n1005), .A2(n1048), .ZN(n1047) );
INV_X1 U758 ( .A(n1049), .ZN(n1020) );
XOR2_X1 U759 ( .A(n1050), .B(n1051), .Z(G72) );
XOR2_X1 U760 ( .A(n1052), .B(n1053), .Z(n1051) );
NOR2_X1 U761 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U762 ( .A(n1056), .B(KEYINPUT57), .Z(n1055) );
NAND2_X1 U763 ( .A1(G900), .A2(G227), .ZN(n1056) );
NAND2_X1 U764 ( .A1(n1057), .A2(n1058), .ZN(n1052) );
NAND2_X1 U765 ( .A1(G953), .A2(n1059), .ZN(n1058) );
XOR2_X1 U766 ( .A(n1060), .B(n1061), .Z(n1057) );
XOR2_X1 U767 ( .A(n1062), .B(n1063), .Z(n1061) );
XOR2_X1 U768 ( .A(n1064), .B(n1065), .Z(n1062) );
NAND2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NAND2_X1 U770 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U771 ( .A1(KEYINPUT52), .A2(G140), .ZN(n1069) );
NAND2_X1 U772 ( .A1(KEYINPUT52), .A2(n1070), .ZN(n1066) );
XOR2_X1 U773 ( .A(n1071), .B(n1072), .Z(n1060) );
XOR2_X1 U774 ( .A(KEYINPUT63), .B(n1073), .Z(n1072) );
NOR2_X1 U775 ( .A1(KEYINPUT26), .A2(n1074), .ZN(n1073) );
XNOR2_X1 U776 ( .A(KEYINPUT46), .B(n1075), .ZN(n1074) );
INV_X1 U777 ( .A(G134), .ZN(n1075) );
NAND2_X1 U778 ( .A1(KEYINPUT0), .A2(n1076), .ZN(n1071) );
NAND2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1050) );
NAND2_X1 U780 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U781 ( .A(KEYINPUT41), .B(n1081), .Z(n1080) );
XNOR2_X1 U782 ( .A(G953), .B(KEYINPUT30), .ZN(n1077) );
XOR2_X1 U783 ( .A(n1082), .B(n1083), .Z(G69) );
NOR2_X1 U784 ( .A1(n1084), .A2(n1054), .ZN(n1083) );
XNOR2_X1 U785 ( .A(G953), .B(KEYINPUT27), .ZN(n1054) );
NOR2_X1 U786 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR3_X1 U787 ( .A1(n1087), .A2(KEYINPUT3), .A3(n1088), .ZN(n1082) );
NOR3_X1 U788 ( .A1(n1089), .A2(G953), .A3(n1090), .ZN(n1088) );
NOR2_X1 U789 ( .A1(n1091), .A2(n1092), .ZN(n1087) );
XOR2_X1 U790 ( .A(n1093), .B(KEYINPUT61), .Z(n1092) );
NAND2_X1 U791 ( .A1(n997), .A2(n1094), .ZN(n1093) );
NOR2_X1 U792 ( .A1(n1095), .A2(n1089), .ZN(n1091) );
NOR2_X1 U793 ( .A1(G898), .A2(n997), .ZN(n1095) );
NOR2_X1 U794 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XOR2_X1 U795 ( .A(KEYINPUT42), .B(n1098), .Z(n1097) );
XOR2_X1 U796 ( .A(n1099), .B(n1100), .Z(n1096) );
NOR2_X1 U797 ( .A1(n1015), .A2(n1101), .ZN(n1099) );
NOR2_X1 U798 ( .A1(n1098), .A2(n1102), .ZN(G63) );
NOR3_X1 U799 ( .A1(n1009), .A2(n1103), .A3(n1104), .ZN(n1102) );
NOR4_X1 U800 ( .A1(n1105), .A2(n1101), .A3(KEYINPUT55), .A4(n1011), .ZN(n1104) );
NOR2_X1 U801 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NOR3_X1 U802 ( .A1(n1011), .A2(KEYINPUT55), .A3(n994), .ZN(n1107) );
INV_X1 U803 ( .A(G478), .ZN(n1011) );
NOR2_X1 U804 ( .A1(n1098), .A2(n1108), .ZN(G60) );
XOR2_X1 U805 ( .A(n1109), .B(n1110), .Z(n1108) );
XNOR2_X1 U806 ( .A(KEYINPUT5), .B(n1111), .ZN(n1110) );
AND2_X1 U807 ( .A1(G475), .A2(n1112), .ZN(n1109) );
XOR2_X1 U808 ( .A(G104), .B(n1113), .Z(G6) );
NOR3_X1 U809 ( .A1(n1098), .A2(n1114), .A3(n1115), .ZN(G57) );
NOR2_X1 U810 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U811 ( .A(n1118), .B(KEYINPUT59), .Z(n1117) );
INV_X1 U812 ( .A(n1119), .ZN(n1116) );
NOR2_X1 U813 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
XNOR2_X1 U814 ( .A(KEYINPUT58), .B(n1118), .ZN(n1120) );
NAND3_X1 U815 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1118) );
NAND2_X1 U816 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND3_X1 U817 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1122) );
NAND2_X1 U818 ( .A1(n1129), .A2(G101), .ZN(n1121) );
XNOR2_X1 U819 ( .A(n1126), .B(n1125), .ZN(n1129) );
INV_X1 U820 ( .A(n1127), .ZN(n1125) );
NAND2_X1 U821 ( .A1(n1112), .A2(G472), .ZN(n1127) );
NOR3_X1 U822 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(G54) );
NOR3_X1 U823 ( .A1(n1133), .A2(G953), .A3(G952), .ZN(n1132) );
AND2_X1 U824 ( .A1(n1133), .A2(n1098), .ZN(n1131) );
INV_X1 U825 ( .A(KEYINPUT19), .ZN(n1133) );
XOR2_X1 U826 ( .A(n1134), .B(n1135), .Z(n1130) );
XOR2_X1 U827 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U828 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U829 ( .A1(KEYINPUT60), .A2(n1140), .ZN(n1138) );
XOR2_X1 U830 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U831 ( .A(KEYINPUT31), .B(n1143), .ZN(n1142) );
XNOR2_X1 U832 ( .A(n1144), .B(n1145), .ZN(n1136) );
NAND3_X1 U833 ( .A1(n1112), .A2(G469), .A3(KEYINPUT21), .ZN(n1144) );
XOR2_X1 U834 ( .A(n1146), .B(n1147), .Z(n1134) );
XNOR2_X1 U835 ( .A(n1148), .B(G110), .ZN(n1147) );
XOR2_X1 U836 ( .A(KEYINPUT53), .B(KEYINPUT24), .Z(n1146) );
NOR2_X1 U837 ( .A1(n1098), .A2(n1149), .ZN(G51) );
XNOR2_X1 U838 ( .A(n1150), .B(n1151), .ZN(n1149) );
XNOR2_X1 U839 ( .A(n1152), .B(n1153), .ZN(n1151) );
NOR2_X1 U840 ( .A1(KEYINPUT47), .A2(n1154), .ZN(n1153) );
XNOR2_X1 U841 ( .A(n1155), .B(n1156), .ZN(n1154) );
NOR2_X1 U842 ( .A1(KEYINPUT1), .A2(n1157), .ZN(n1156) );
NAND2_X1 U843 ( .A1(KEYINPUT9), .A2(n1158), .ZN(n1152) );
OR2_X1 U844 ( .A1(n1101), .A2(n1018), .ZN(n1158) );
INV_X1 U845 ( .A(n1112), .ZN(n1101) );
NOR2_X1 U846 ( .A1(n1159), .A2(n994), .ZN(n1112) );
AND3_X1 U847 ( .A1(n1079), .A2(n1090), .A3(n1081), .ZN(n994) );
AND4_X1 U848 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1081) );
INV_X1 U849 ( .A(n1094), .ZN(n1090) );
NAND2_X1 U850 ( .A1(n1164), .A2(n1165), .ZN(n1094) );
NOR4_X1 U851 ( .A1(n1166), .A2(n1167), .A3(n1113), .A4(n1168), .ZN(n1165) );
INV_X1 U852 ( .A(n1169), .ZN(n1168) );
NOR3_X1 U853 ( .A1(n1029), .A2(n1170), .A3(n1171), .ZN(n1113) );
NOR4_X1 U854 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1164) );
NOR2_X1 U855 ( .A1(n993), .A2(n1176), .ZN(n1175) );
INV_X1 U856 ( .A(n1177), .ZN(n993) );
NOR3_X1 U857 ( .A1(n1171), .A2(n1170), .A3(n1030), .ZN(n1174) );
NOR4_X1 U858 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1173) );
XNOR2_X1 U859 ( .A(KEYINPUT23), .B(n1170), .ZN(n1181) );
INV_X1 U860 ( .A(n1182), .ZN(n1172) );
AND4_X1 U861 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1079) );
NOR2_X1 U862 ( .A1(n997), .A2(G952), .ZN(n1098) );
XNOR2_X1 U863 ( .A(G146), .B(n1183), .ZN(G48) );
NAND3_X1 U864 ( .A1(n1187), .A2(n1177), .A3(n1188), .ZN(n1183) );
XNOR2_X1 U865 ( .A(G143), .B(n1184), .ZN(G45) );
NAND4_X1 U866 ( .A1(n1189), .A2(n1177), .A3(n1019), .A4(n1190), .ZN(n1184) );
XNOR2_X1 U867 ( .A(n1148), .B(n1191), .ZN(G42) );
NOR2_X1 U868 ( .A1(KEYINPUT13), .A2(n1185), .ZN(n1191) );
NAND3_X1 U869 ( .A1(n1192), .A2(n1037), .A3(n1025), .ZN(n1185) );
XNOR2_X1 U870 ( .A(G137), .B(n1186), .ZN(G39) );
NAND3_X1 U871 ( .A1(n1188), .A2(n1031), .A3(n1025), .ZN(n1186) );
XNOR2_X1 U872 ( .A(G134), .B(n1160), .ZN(G36) );
NAND3_X1 U873 ( .A1(n1189), .A2(n986), .A3(n1025), .ZN(n1160) );
XNOR2_X1 U874 ( .A(G131), .B(n1161), .ZN(G33) );
NAND3_X1 U875 ( .A1(n1189), .A2(n1187), .A3(n1025), .ZN(n1161) );
AND2_X1 U876 ( .A1(n1048), .A2(n1193), .ZN(n1025) );
AND3_X1 U877 ( .A1(n1037), .A2(n1194), .A3(n1195), .ZN(n1189) );
XNOR2_X1 U878 ( .A(G128), .B(n1162), .ZN(G30) );
NAND3_X1 U879 ( .A1(n986), .A2(n1177), .A3(n1188), .ZN(n1162) );
AND4_X1 U880 ( .A1(n1196), .A2(n1037), .A3(n1194), .A4(n1045), .ZN(n1188) );
XNOR2_X1 U881 ( .A(G101), .B(n1197), .ZN(G3) );
NAND2_X1 U882 ( .A1(n1198), .A2(n1177), .ZN(n1197) );
XOR2_X1 U883 ( .A(n1176), .B(KEYINPUT51), .Z(n1198) );
NAND3_X1 U884 ( .A1(n992), .A2(n1031), .A3(n1195), .ZN(n1176) );
INV_X1 U885 ( .A(n1042), .ZN(n1195) );
XNOR2_X1 U886 ( .A(G125), .B(n1163), .ZN(G27) );
NAND3_X1 U887 ( .A1(n1192), .A2(n1177), .A3(n999), .ZN(n1163) );
AND4_X1 U888 ( .A1(n1187), .A2(n1044), .A3(n1194), .A4(n1045), .ZN(n1192) );
NAND2_X1 U889 ( .A1(n1049), .A2(n1199), .ZN(n1194) );
NAND4_X1 U890 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1059), .ZN(n1199) );
INV_X1 U891 ( .A(G900), .ZN(n1059) );
XOR2_X1 U892 ( .A(G122), .B(n1201), .Z(G24) );
NOR4_X1 U893 ( .A1(n1178), .A2(n1179), .A3(n1170), .A4(n1180), .ZN(n1201) );
INV_X1 U894 ( .A(n987), .ZN(n1170) );
NOR2_X1 U895 ( .A1(n1202), .A2(n1045), .ZN(n987) );
XNOR2_X1 U896 ( .A(G119), .B(n1182), .ZN(G21) );
NAND4_X1 U897 ( .A1(n1196), .A2(n1203), .A3(n1031), .A4(n1045), .ZN(n1182) );
INV_X1 U898 ( .A(n1180), .ZN(n1203) );
XNOR2_X1 U899 ( .A(n1204), .B(n1167), .ZN(G18) );
NOR3_X1 U900 ( .A1(n1042), .A2(n1030), .A3(n1180), .ZN(n1167) );
INV_X1 U901 ( .A(n986), .ZN(n1030) );
NOR2_X1 U902 ( .A1(n1019), .A2(n1178), .ZN(n986) );
XNOR2_X1 U903 ( .A(n1205), .B(n1166), .ZN(G15) );
NOR3_X1 U904 ( .A1(n1042), .A2(n1029), .A3(n1180), .ZN(n1166) );
NAND3_X1 U905 ( .A1(n1177), .A2(n1206), .A3(n999), .ZN(n1180) );
NOR2_X1 U906 ( .A1(n1207), .A2(n1035), .ZN(n999) );
NAND2_X1 U907 ( .A1(n1196), .A2(n1208), .ZN(n1042) );
XNOR2_X1 U908 ( .A(n1044), .B(KEYINPUT44), .ZN(n1196) );
XNOR2_X1 U909 ( .A(G110), .B(n1169), .ZN(G12) );
NAND4_X1 U910 ( .A1(n990), .A2(n1044), .A3(n1031), .A4(n1045), .ZN(n1169) );
INV_X1 U911 ( .A(n1208), .ZN(n1045) );
NOR2_X1 U912 ( .A1(n1004), .A2(n1209), .ZN(n1208) );
NOR2_X1 U913 ( .A1(n1015), .A2(n1016), .ZN(n1209) );
AND2_X1 U914 ( .A1(n1016), .A2(n1015), .ZN(n1004) );
NAND2_X1 U915 ( .A1(G217), .A2(n1210), .ZN(n1015) );
NOR2_X1 U916 ( .A1(n1100), .A2(G902), .ZN(n1016) );
XNOR2_X1 U917 ( .A(n1211), .B(n1212), .ZN(n1100) );
XOR2_X1 U918 ( .A(n1213), .B(n1214), .Z(n1212) );
XNOR2_X1 U919 ( .A(n1215), .B(G110), .ZN(n1214) );
XOR2_X1 U920 ( .A(KEYINPUT39), .B(G128), .Z(n1213) );
XOR2_X1 U921 ( .A(n1216), .B(n1063), .Z(n1211) );
XOR2_X1 U922 ( .A(n1217), .B(n1218), .Z(n1216) );
AND2_X1 U923 ( .A1(n1219), .A2(G221), .ZN(n1218) );
NAND3_X1 U924 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1217) );
NAND2_X1 U925 ( .A1(KEYINPUT50), .A2(n1068), .ZN(n1221) );
OR2_X1 U926 ( .A1(n1223), .A2(KEYINPUT50), .ZN(n1220) );
NAND2_X1 U927 ( .A1(n1224), .A2(n1225), .ZN(n1031) );
OR2_X1 U928 ( .A1(n1029), .A2(KEYINPUT48), .ZN(n1225) );
INV_X1 U929 ( .A(n1187), .ZN(n1029) );
NOR2_X1 U930 ( .A1(n1190), .A2(n1179), .ZN(n1187) );
NAND3_X1 U931 ( .A1(n1178), .A2(n1179), .A3(KEYINPUT48), .ZN(n1224) );
INV_X1 U932 ( .A(n1019), .ZN(n1179) );
XNOR2_X1 U933 ( .A(n1226), .B(G475), .ZN(n1019) );
NAND2_X1 U934 ( .A1(n1159), .A2(n1111), .ZN(n1226) );
NAND2_X1 U935 ( .A1(n1227), .A2(n1228), .ZN(n1111) );
NAND2_X1 U936 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
XOR2_X1 U937 ( .A(KEYINPUT32), .B(n1231), .Z(n1227) );
NOR2_X1 U938 ( .A1(n1229), .A2(n1230), .ZN(n1231) );
XNOR2_X1 U939 ( .A(G104), .B(n1232), .ZN(n1230) );
XNOR2_X1 U940 ( .A(G122), .B(n1205), .ZN(n1232) );
XNOR2_X1 U941 ( .A(n1233), .B(n1234), .ZN(n1229) );
XOR2_X1 U942 ( .A(n1076), .B(n1235), .Z(n1234) );
NAND2_X1 U943 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U944 ( .A1(G143), .A2(n1238), .ZN(n1237) );
NAND2_X1 U945 ( .A1(n1223), .A2(n1222), .ZN(n1238) );
NAND2_X1 U946 ( .A1(n1068), .A2(n1148), .ZN(n1222) );
INV_X1 U947 ( .A(n1070), .ZN(n1223) );
NOR2_X1 U948 ( .A1(n1148), .A2(n1068), .ZN(n1070) );
INV_X1 U949 ( .A(G140), .ZN(n1148) );
NAND2_X1 U950 ( .A1(n1239), .A2(n1240), .ZN(n1236) );
XNOR2_X1 U951 ( .A(G140), .B(n1068), .ZN(n1239) );
XOR2_X1 U952 ( .A(n1143), .B(n1241), .Z(n1233) );
NOR3_X1 U953 ( .A1(n1242), .A2(G237), .A3(n1243), .ZN(n1241) );
INV_X1 U954 ( .A(G214), .ZN(n1243) );
XNOR2_X1 U955 ( .A(KEYINPUT25), .B(n997), .ZN(n1242) );
INV_X1 U956 ( .A(n1190), .ZN(n1178) );
NAND2_X1 U957 ( .A1(n1244), .A2(n1245), .ZN(n1190) );
NAND2_X1 U958 ( .A1(G478), .A2(n1246), .ZN(n1245) );
XOR2_X1 U959 ( .A(KEYINPUT34), .B(n1247), .Z(n1244) );
NOR2_X1 U960 ( .A1(G478), .A2(n1246), .ZN(n1247) );
INV_X1 U961 ( .A(n1009), .ZN(n1246) );
NOR2_X1 U962 ( .A1(G902), .A2(n1106), .ZN(n1009) );
INV_X1 U963 ( .A(n1105), .ZN(n1106) );
NAND2_X1 U964 ( .A1(n1248), .A2(n1249), .ZN(n1105) );
NAND4_X1 U965 ( .A1(G217), .A2(n1219), .A3(n1250), .A4(n1251), .ZN(n1249) );
NAND2_X1 U966 ( .A1(n1252), .A2(n1253), .ZN(n1248) );
NAND2_X1 U967 ( .A1(n1250), .A2(n1251), .ZN(n1253) );
NAND2_X1 U968 ( .A1(n1254), .A2(n1255), .ZN(n1251) );
INV_X1 U969 ( .A(n1256), .ZN(n1255) );
XNOR2_X1 U970 ( .A(n1257), .B(n1258), .ZN(n1254) );
XOR2_X1 U971 ( .A(n1259), .B(KEYINPUT54), .Z(n1250) );
NAND2_X1 U972 ( .A1(n1260), .A2(n1256), .ZN(n1259) );
NAND3_X1 U973 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1256) );
OR2_X1 U974 ( .A1(n1264), .A2(G134), .ZN(n1263) );
NAND2_X1 U975 ( .A1(n1265), .A2(n1266), .ZN(n1262) );
INV_X1 U976 ( .A(KEYINPUT43), .ZN(n1266) );
NAND2_X1 U977 ( .A1(n1267), .A2(n1264), .ZN(n1265) );
XNOR2_X1 U978 ( .A(KEYINPUT40), .B(G134), .ZN(n1267) );
NAND2_X1 U979 ( .A1(KEYINPUT43), .A2(n1268), .ZN(n1261) );
NAND2_X1 U980 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
OR2_X1 U981 ( .A1(G134), .A2(KEYINPUT40), .ZN(n1270) );
NAND3_X1 U982 ( .A1(G134), .A2(n1264), .A3(KEYINPUT40), .ZN(n1269) );
XOR2_X1 U983 ( .A(n1065), .B(KEYINPUT4), .Z(n1264) );
XNOR2_X1 U984 ( .A(n1258), .B(n1271), .ZN(n1260) );
INV_X1 U985 ( .A(n1257), .ZN(n1271) );
NAND2_X1 U986 ( .A1(G217), .A2(n1219), .ZN(n1252) );
AND2_X1 U987 ( .A1(n1272), .A2(n997), .ZN(n1219) );
XNOR2_X1 U988 ( .A(G234), .B(KEYINPUT14), .ZN(n1272) );
INV_X1 U989 ( .A(n1202), .ZN(n1044) );
NAND2_X1 U990 ( .A1(n1273), .A2(n1006), .ZN(n1202) );
NAND2_X1 U991 ( .A1(G472), .A2(n1274), .ZN(n1006) );
XNOR2_X1 U992 ( .A(KEYINPUT45), .B(n1008), .ZN(n1273) );
OR2_X1 U993 ( .A1(n1274), .A2(G472), .ZN(n1008) );
NAND2_X1 U994 ( .A1(n1275), .A2(n1159), .ZN(n1274) );
XNOR2_X1 U995 ( .A(n1119), .B(n1276), .ZN(n1275) );
NOR2_X1 U996 ( .A1(n1124), .A2(n1277), .ZN(n1276) );
XOR2_X1 U997 ( .A(KEYINPUT7), .B(n1278), .Z(n1277) );
NOR2_X1 U998 ( .A1(n1128), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U999 ( .A(KEYINPUT8), .B(n1280), .ZN(n1279) );
NOR2_X1 U1000 ( .A1(G101), .A2(n1126), .ZN(n1124) );
INV_X1 U1001 ( .A(n1280), .ZN(n1126) );
NAND3_X1 U1002 ( .A1(n1281), .A2(n997), .A3(G210), .ZN(n1280) );
XNOR2_X1 U1003 ( .A(n1282), .B(n1283), .ZN(n1119) );
XNOR2_X1 U1004 ( .A(n1205), .B(n1284), .ZN(n1283) );
NOR2_X1 U1005 ( .A1(KEYINPUT15), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U1006 ( .A(G119), .B(n1286), .ZN(n1285) );
NOR2_X1 U1007 ( .A1(KEYINPUT29), .A2(n1204), .ZN(n1286) );
INV_X1 U1008 ( .A(G113), .ZN(n1205) );
XNOR2_X1 U1009 ( .A(n1139), .B(n1287), .ZN(n1282) );
XOR2_X1 U1010 ( .A(G137), .B(n1288), .Z(n1139) );
INV_X1 U1011 ( .A(n1171), .ZN(n990) );
NAND2_X1 U1012 ( .A1(n1177), .A2(n992), .ZN(n1171) );
AND2_X1 U1013 ( .A1(n1037), .A2(n1206), .ZN(n992) );
NAND2_X1 U1014 ( .A1(n1049), .A2(n1289), .ZN(n1206) );
NAND4_X1 U1015 ( .A1(G902), .A2(G953), .A3(n1200), .A4(n1086), .ZN(n1289) );
INV_X1 U1016 ( .A(G898), .ZN(n1086) );
NAND3_X1 U1017 ( .A1(n1200), .A2(n997), .A3(G952), .ZN(n1049) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1200) );
NOR2_X1 U1019 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
AND2_X1 U1020 ( .A1(G221), .A2(n1210), .ZN(n1035) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1159), .ZN(n1210) );
INV_X1 U1022 ( .A(n1207), .ZN(n1036) );
XNOR2_X1 U1023 ( .A(n1290), .B(G469), .ZN(n1207) );
NAND2_X1 U1024 ( .A1(n1291), .A2(n1159), .ZN(n1290) );
XOR2_X1 U1025 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U1026 ( .A(n1288), .B(n1294), .Z(n1293) );
XOR2_X1 U1027 ( .A(n1141), .B(n1063), .Z(n1294) );
XNOR2_X1 U1028 ( .A(G137), .B(n1143), .ZN(n1063) );
XOR2_X1 U1029 ( .A(n1065), .B(n1295), .Z(n1141) );
XNOR2_X1 U1030 ( .A(n1128), .B(n1296), .ZN(n1295) );
NOR2_X1 U1031 ( .A1(KEYINPUT49), .A2(n1297), .ZN(n1296) );
INV_X1 U1032 ( .A(G101), .ZN(n1128) );
XOR2_X1 U1033 ( .A(n1298), .B(n1076), .Z(n1288) );
XNOR2_X1 U1034 ( .A(G131), .B(KEYINPUT56), .ZN(n1076) );
XNOR2_X1 U1035 ( .A(G134), .B(KEYINPUT33), .ZN(n1298) );
XOR2_X1 U1036 ( .A(n1299), .B(n1300), .Z(n1292) );
XOR2_X1 U1037 ( .A(n1145), .B(KEYINPUT10), .Z(n1300) );
NAND2_X1 U1038 ( .A1(G227), .A2(n997), .ZN(n1145) );
INV_X1 U1039 ( .A(G953), .ZN(n997) );
NAND2_X1 U1040 ( .A1(KEYINPUT11), .A2(n1301), .ZN(n1299) );
XNOR2_X1 U1041 ( .A(n1302), .B(n1303), .ZN(n1301) );
NOR2_X1 U1042 ( .A1(G140), .A2(KEYINPUT22), .ZN(n1303) );
NOR2_X1 U1043 ( .A1(n1048), .A2(n1005), .ZN(n1177) );
INV_X1 U1044 ( .A(n1193), .ZN(n1005) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1304), .ZN(n1193) );
XOR2_X1 U1046 ( .A(n1305), .B(n1017), .Z(n1048) );
NAND2_X1 U1047 ( .A1(n1306), .A2(n1159), .ZN(n1017) );
XNOR2_X1 U1048 ( .A(n1307), .B(n1157), .ZN(n1306) );
INV_X1 U1049 ( .A(n1068), .ZN(n1157) );
XOR2_X1 U1050 ( .A(G125), .B(KEYINPUT18), .Z(n1068) );
XNOR2_X1 U1051 ( .A(n1308), .B(n1309), .ZN(n1307) );
INV_X1 U1052 ( .A(n1155), .ZN(n1309) );
XOR2_X1 U1053 ( .A(n1287), .B(n1310), .Z(n1155) );
NOR2_X1 U1054 ( .A1(G953), .A2(n1085), .ZN(n1310) );
INV_X1 U1055 ( .A(G224), .ZN(n1085) );
XOR2_X1 U1056 ( .A(n1065), .B(n1311), .Z(n1287) );
NOR2_X1 U1057 ( .A1(KEYINPUT62), .A2(n1143), .ZN(n1311) );
XNOR2_X1 U1058 ( .A(G146), .B(KEYINPUT17), .ZN(n1143) );
XNOR2_X1 U1059 ( .A(G128), .B(n1240), .ZN(n1065) );
INV_X1 U1060 ( .A(G143), .ZN(n1240) );
NAND2_X1 U1061 ( .A1(KEYINPUT16), .A2(n1150), .ZN(n1308) );
INV_X1 U1062 ( .A(n1089), .ZN(n1150) );
XNOR2_X1 U1063 ( .A(n1312), .B(n1313), .ZN(n1089) );
XOR2_X1 U1064 ( .A(n1258), .B(n1314), .Z(n1313) );
XNOR2_X1 U1065 ( .A(n1315), .B(n1316), .ZN(n1314) );
NOR2_X1 U1066 ( .A1(KEYINPUT12), .A2(n1297), .ZN(n1316) );
XNOR2_X1 U1067 ( .A(G104), .B(n1257), .ZN(n1297) );
XOR2_X1 U1068 ( .A(G107), .B(KEYINPUT36), .Z(n1257) );
NAND2_X1 U1069 ( .A1(KEYINPUT6), .A2(n1302), .ZN(n1315) );
INV_X1 U1070 ( .A(G110), .ZN(n1302) );
XNOR2_X1 U1071 ( .A(n1204), .B(G122), .ZN(n1258) );
INV_X1 U1072 ( .A(G116), .ZN(n1204) );
XOR2_X1 U1073 ( .A(n1317), .B(n1318), .Z(n1312) );
XNOR2_X1 U1074 ( .A(KEYINPUT28), .B(n1215), .ZN(n1318) );
INV_X1 U1075 ( .A(G119), .ZN(n1215) );
XNOR2_X1 U1076 ( .A(G113), .B(G101), .ZN(n1317) );
NAND2_X1 U1077 ( .A1(KEYINPUT35), .A2(n1018), .ZN(n1305) );
NAND2_X1 U1078 ( .A1(G210), .A2(n1304), .ZN(n1018) );
NAND2_X1 U1079 ( .A1(n1281), .A2(n1159), .ZN(n1304) );
INV_X1 U1080 ( .A(G902), .ZN(n1159) );
INV_X1 U1081 ( .A(G237), .ZN(n1281) );
endmodule


