//Key = 1010011100100110001010000100001001100100011101111011110110101110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282;

XNOR2_X1 U701 ( .A(G107), .B(n980), .ZN(G9) );
NOR2_X1 U702 ( .A1(n981), .A2(n982), .ZN(G75) );
NOR3_X1 U703 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n982) );
NOR2_X1 U704 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U705 ( .A1(n988), .A2(n989), .ZN(n986) );
XOR2_X1 U706 ( .A(n990), .B(KEYINPUT41), .Z(n989) );
NAND4_X1 U707 ( .A1(n991), .A2(n992), .A3(n993), .A4(n994), .ZN(n990) );
NOR3_X1 U708 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n988) );
NOR2_X1 U709 ( .A1(n998), .A2(n999), .ZN(n997) );
AND2_X1 U710 ( .A1(n1000), .A2(n992), .ZN(n998) );
NOR2_X1 U711 ( .A1(n991), .A2(n1001), .ZN(n996) );
NOR4_X1 U712 ( .A1(KEYINPUT48), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1001) );
INV_X1 U713 ( .A(n1005), .ZN(n1002) );
INV_X1 U714 ( .A(n994), .ZN(n995) );
NAND3_X1 U715 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n983) );
NAND3_X1 U716 ( .A1(n1005), .A2(n1009), .A3(n991), .ZN(n1008) );
NAND2_X1 U717 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND3_X1 U718 ( .A1(n994), .A2(n1012), .A3(n1013), .ZN(n1011) );
NAND2_X1 U719 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NAND3_X1 U720 ( .A1(n1016), .A2(n1017), .A3(KEYINPUT48), .ZN(n1015) );
INV_X1 U721 ( .A(n1018), .ZN(n1014) );
NAND2_X1 U722 ( .A1(n992), .A2(n1019), .ZN(n1010) );
NAND3_X1 U723 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1019) );
NAND2_X1 U724 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
XNOR2_X1 U725 ( .A(KEYINPUT16), .B(n987), .ZN(n1024) );
NAND3_X1 U726 ( .A1(n1025), .A2(n1026), .A3(n1013), .ZN(n1021) );
NAND2_X1 U727 ( .A1(n994), .A2(n1027), .ZN(n1020) );
NAND2_X1 U728 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U729 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
AND3_X1 U730 ( .A1(n1006), .A2(n1007), .A3(n1032), .ZN(n981) );
NAND4_X1 U731 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1006) );
NOR4_X1 U732 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
XNOR2_X1 U733 ( .A(n1041), .B(n1042), .ZN(n1040) );
XOR2_X1 U734 ( .A(n1043), .B(n1044), .Z(n1039) );
NOR3_X1 U735 ( .A1(n1017), .A2(n1045), .A3(n1030), .ZN(n1035) );
NAND2_X1 U736 ( .A1(n1046), .A2(n1047), .ZN(G72) );
NAND2_X1 U737 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XOR2_X1 U738 ( .A(KEYINPUT37), .B(n1050), .Z(n1046) );
NOR2_X1 U739 ( .A1(n1048), .A2(n1049), .ZN(n1050) );
NAND2_X1 U740 ( .A1(G953), .A2(n1051), .ZN(n1049) );
NAND2_X1 U741 ( .A1(G900), .A2(G227), .ZN(n1051) );
NAND2_X1 U742 ( .A1(n1052), .A2(n1053), .ZN(n1048) );
NAND2_X1 U743 ( .A1(n1054), .A2(n1007), .ZN(n1053) );
XNOR2_X1 U744 ( .A(n1055), .B(n1056), .ZN(n1054) );
NAND3_X1 U745 ( .A1(G900), .A2(n1056), .A3(G953), .ZN(n1052) );
XOR2_X1 U746 ( .A(n1057), .B(n1058), .Z(n1056) );
XNOR2_X1 U747 ( .A(n1059), .B(n1060), .ZN(n1058) );
INV_X1 U748 ( .A(G140), .ZN(n1059) );
XOR2_X1 U749 ( .A(n1061), .B(n1062), .Z(G69) );
XOR2_X1 U750 ( .A(n1063), .B(n1064), .Z(n1062) );
NAND2_X1 U751 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
OR2_X1 U752 ( .A1(n1007), .A2(G898), .ZN(n1066) );
XOR2_X1 U753 ( .A(n1067), .B(n1068), .Z(n1065) );
XOR2_X1 U754 ( .A(n1069), .B(n1070), .Z(n1068) );
NAND2_X1 U755 ( .A1(KEYINPUT34), .A2(n1071), .ZN(n1069) );
XNOR2_X1 U756 ( .A(n1072), .B(KEYINPUT38), .ZN(n1067) );
NAND2_X1 U757 ( .A1(KEYINPUT61), .A2(n1073), .ZN(n1072) );
NAND2_X1 U758 ( .A1(G953), .A2(n1074), .ZN(n1063) );
NAND2_X1 U759 ( .A1(n1075), .A2(G224), .ZN(n1074) );
XNOR2_X1 U760 ( .A(G898), .B(KEYINPUT6), .ZN(n1075) );
NOR2_X1 U761 ( .A1(n1076), .A2(G953), .ZN(n1061) );
NOR2_X1 U762 ( .A1(n1077), .A2(n1078), .ZN(G66) );
NOR3_X1 U763 ( .A1(n1041), .A2(n1079), .A3(n1080), .ZN(n1078) );
NOR3_X1 U764 ( .A1(n1081), .A2(n1042), .A3(n1082), .ZN(n1080) );
INV_X1 U765 ( .A(n1083), .ZN(n1081) );
NOR2_X1 U766 ( .A1(n1084), .A2(n1083), .ZN(n1079) );
NOR2_X1 U767 ( .A1(n1085), .A2(n1042), .ZN(n1084) );
NOR2_X1 U768 ( .A1(n1077), .A2(n1086), .ZN(G63) );
XOR2_X1 U769 ( .A(n1087), .B(n1088), .Z(n1086) );
AND2_X1 U770 ( .A1(G478), .A2(n1089), .ZN(n1088) );
NOR2_X1 U771 ( .A1(n1077), .A2(n1090), .ZN(G60) );
XOR2_X1 U772 ( .A(n1091), .B(n1092), .Z(n1090) );
NOR2_X1 U773 ( .A1(KEYINPUT59), .A2(n1093), .ZN(n1092) );
XNOR2_X1 U774 ( .A(n1094), .B(n1095), .ZN(n1093) );
NAND2_X1 U775 ( .A1(n1089), .A2(G475), .ZN(n1091) );
XNOR2_X1 U776 ( .A(G104), .B(n1096), .ZN(G6) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1097), .ZN(G57) );
XOR2_X1 U778 ( .A(n1098), .B(n1099), .Z(n1097) );
XOR2_X1 U779 ( .A(n1100), .B(n1101), .Z(n1099) );
AND2_X1 U780 ( .A1(G472), .A2(n1089), .ZN(n1101) );
NAND2_X1 U781 ( .A1(n1102), .A2(KEYINPUT0), .ZN(n1100) );
XOR2_X1 U782 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U783 ( .A(KEYINPUT20), .B(n1105), .Z(n1104) );
NOR2_X1 U784 ( .A1(KEYINPUT22), .A2(n1106), .ZN(n1105) );
INV_X1 U785 ( .A(n1107), .ZN(n1106) );
XOR2_X1 U786 ( .A(n1108), .B(n1109), .Z(n1103) );
XNOR2_X1 U787 ( .A(n1110), .B(n1111), .ZN(n1098) );
NOR2_X1 U788 ( .A1(n1077), .A2(n1112), .ZN(G54) );
XOR2_X1 U789 ( .A(n1113), .B(n1114), .Z(n1112) );
XNOR2_X1 U790 ( .A(n1108), .B(n1115), .ZN(n1114) );
XOR2_X1 U791 ( .A(n1116), .B(n1117), .Z(n1113) );
AND2_X1 U792 ( .A1(G469), .A2(n1089), .ZN(n1117) );
NOR2_X1 U793 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
XOR2_X1 U794 ( .A(KEYINPUT17), .B(n1120), .Z(n1119) );
AND2_X1 U795 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U796 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
XNOR2_X1 U797 ( .A(n1123), .B(KEYINPUT52), .ZN(n1122) );
NOR2_X1 U798 ( .A1(n1077), .A2(n1124), .ZN(G51) );
XOR2_X1 U799 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR3_X1 U800 ( .A1(n1082), .A2(KEYINPUT19), .A3(n1044), .ZN(n1125) );
INV_X1 U801 ( .A(n1089), .ZN(n1082) );
NOR2_X1 U802 ( .A1(n1127), .A2(n1085), .ZN(n1089) );
INV_X1 U803 ( .A(n985), .ZN(n1085) );
NAND2_X1 U804 ( .A1(n1055), .A2(n1076), .ZN(n985) );
AND4_X1 U805 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1076) );
AND4_X1 U806 ( .A1(n1096), .A2(n980), .A3(n1132), .A4(n1133), .ZN(n1131) );
NAND3_X1 U807 ( .A1(n993), .A2(n994), .A3(n1134), .ZN(n980) );
NAND3_X1 U808 ( .A1(n1134), .A2(n994), .A3(n1000), .ZN(n1096) );
NOR3_X1 U809 ( .A1(n1135), .A2(n1136), .A3(n1137), .ZN(n1130) );
NOR3_X1 U810 ( .A1(n1138), .A2(n1139), .A3(n1028), .ZN(n1137) );
INV_X1 U811 ( .A(KEYINPUT21), .ZN(n1138) );
NOR2_X1 U812 ( .A1(KEYINPUT21), .A2(n1140), .ZN(n1136) );
INV_X1 U813 ( .A(n1141), .ZN(n1135) );
AND4_X1 U814 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1055) );
NOR4_X1 U815 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
AND2_X1 U816 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
NAND2_X1 U817 ( .A1(n1152), .A2(n1153), .ZN(n1142) );
XNOR2_X1 U818 ( .A(KEYINPUT54), .B(n1028), .ZN(n1153) );
INV_X1 U819 ( .A(n1154), .ZN(n1028) );
NOR2_X1 U820 ( .A1(n1007), .A2(G952), .ZN(n1077) );
XNOR2_X1 U821 ( .A(G146), .B(n1155), .ZN(G48) );
NAND2_X1 U822 ( .A1(n1152), .A2(n1154), .ZN(n1155) );
AND2_X1 U823 ( .A1(n1000), .A2(n1156), .ZN(n1152) );
XNOR2_X1 U824 ( .A(G143), .B(n1151), .ZN(G45) );
NAND4_X1 U825 ( .A1(n1157), .A2(n1158), .A3(n1154), .A4(n1159), .ZN(n1151) );
AND3_X1 U826 ( .A1(n1023), .A2(n1018), .A3(n1160), .ZN(n1159) );
XNOR2_X1 U827 ( .A(G140), .B(n1161), .ZN(G42) );
NOR2_X1 U828 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NOR2_X1 U829 ( .A1(n1164), .A2(n1143), .ZN(n1163) );
NAND2_X1 U830 ( .A1(n1165), .A2(n1013), .ZN(n1143) );
INV_X1 U831 ( .A(KEYINPUT45), .ZN(n1164) );
NOR3_X1 U832 ( .A1(KEYINPUT45), .A2(n1165), .A3(n987), .ZN(n1162) );
AND2_X1 U833 ( .A1(n1166), .A2(n1018), .ZN(n1165) );
XOR2_X1 U834 ( .A(n1167), .B(n1149), .Z(G39) );
AND3_X1 U835 ( .A1(n1013), .A2(n1156), .A3(n1005), .ZN(n1149) );
XNOR2_X1 U836 ( .A(G137), .B(KEYINPUT10), .ZN(n1167) );
XOR2_X1 U837 ( .A(G134), .B(n1148), .Z(G36) );
AND2_X1 U838 ( .A1(n1168), .A2(n993), .ZN(n1148) );
XNOR2_X1 U839 ( .A(n1169), .B(n1147), .ZN(G33) );
AND2_X1 U840 ( .A1(n1168), .A2(n1000), .ZN(n1147) );
AND4_X1 U841 ( .A1(n1023), .A2(n1013), .A3(n1018), .A4(n1157), .ZN(n1168) );
INV_X1 U842 ( .A(n987), .ZN(n1013) );
NAND2_X1 U843 ( .A1(n1031), .A2(n1170), .ZN(n987) );
XOR2_X1 U844 ( .A(G128), .B(n1146), .Z(G30) );
AND3_X1 U845 ( .A1(n993), .A2(n1154), .A3(n1156), .ZN(n1146) );
AND4_X1 U846 ( .A1(n1026), .A2(n1018), .A3(n1037), .A4(n1157), .ZN(n1156) );
XNOR2_X1 U847 ( .A(G101), .B(n1141), .ZN(G3) );
NAND3_X1 U848 ( .A1(n1023), .A2(n1134), .A3(n1005), .ZN(n1141) );
XNOR2_X1 U849 ( .A(G125), .B(n1150), .ZN(G27) );
NAND3_X1 U850 ( .A1(n1166), .A2(n1154), .A3(n992), .ZN(n1150) );
AND4_X1 U851 ( .A1(n1026), .A2(n1000), .A3(n1025), .A4(n1157), .ZN(n1166) );
NAND2_X1 U852 ( .A1(n999), .A2(n1171), .ZN(n1157) );
OR4_X1 U853 ( .A1(n1007), .A2(n1127), .A3(n1172), .A4(G900), .ZN(n1171) );
XOR2_X1 U854 ( .A(G122), .B(n1173), .Z(G24) );
NOR2_X1 U855 ( .A1(KEYINPUT12), .A2(n1128), .ZN(n1173) );
NAND4_X1 U856 ( .A1(n1174), .A2(n994), .A3(n1160), .A4(n1158), .ZN(n1128) );
NOR2_X1 U857 ( .A1(n1037), .A2(n1026), .ZN(n994) );
XNOR2_X1 U858 ( .A(G119), .B(n1129), .ZN(G21) );
NAND4_X1 U859 ( .A1(n1174), .A2(n1005), .A3(n1026), .A4(n1037), .ZN(n1129) );
XNOR2_X1 U860 ( .A(G116), .B(n1133), .ZN(G18) );
NAND3_X1 U861 ( .A1(n1023), .A2(n993), .A3(n1174), .ZN(n1133) );
AND3_X1 U862 ( .A1(n1154), .A2(n1175), .A3(n992), .ZN(n1174) );
NOR2_X1 U863 ( .A1(n1158), .A2(n1176), .ZN(n993) );
XNOR2_X1 U864 ( .A(n1140), .B(n1177), .ZN(G15) );
NOR2_X1 U865 ( .A1(KEYINPUT23), .A2(n1178), .ZN(n1177) );
NAND2_X1 U866 ( .A1(n1139), .A2(n1154), .ZN(n1140) );
AND4_X1 U867 ( .A1(n992), .A2(n1000), .A3(n1023), .A4(n1175), .ZN(n1139) );
NOR2_X1 U868 ( .A1(n1026), .A2(n1025), .ZN(n1023) );
AND2_X1 U869 ( .A1(n1176), .A2(n1158), .ZN(n1000) );
NOR2_X1 U870 ( .A1(n1004), .A2(n1017), .ZN(n992) );
XNOR2_X1 U871 ( .A(G110), .B(n1132), .ZN(G12) );
NAND4_X1 U872 ( .A1(n1026), .A2(n1005), .A3(n1025), .A4(n1134), .ZN(n1132) );
AND3_X1 U873 ( .A1(n1154), .A2(n1175), .A3(n1018), .ZN(n1134) );
NOR2_X1 U874 ( .A1(n1016), .A2(n1017), .ZN(n1018) );
INV_X1 U875 ( .A(n1003), .ZN(n1017) );
NAND2_X1 U876 ( .A1(G221), .A2(n1179), .ZN(n1003) );
INV_X1 U877 ( .A(n1004), .ZN(n1016) );
XNOR2_X1 U878 ( .A(n1033), .B(KEYINPUT57), .ZN(n1004) );
XOR2_X1 U879 ( .A(n1180), .B(G469), .Z(n1033) );
NAND2_X1 U880 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U881 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U882 ( .A(n1115), .B(n1185), .Z(n1184) );
XNOR2_X1 U883 ( .A(n1186), .B(n1187), .ZN(n1185) );
NOR2_X1 U884 ( .A1(G140), .A2(KEYINPUT49), .ZN(n1187) );
NAND2_X1 U885 ( .A1(KEYINPUT58), .A2(n1108), .ZN(n1186) );
XNOR2_X1 U886 ( .A(n1188), .B(n1189), .ZN(n1115) );
NAND2_X1 U887 ( .A1(n1190), .A2(KEYINPUT25), .ZN(n1188) );
XNOR2_X1 U888 ( .A(n1191), .B(KEYINPUT39), .ZN(n1190) );
XOR2_X1 U889 ( .A(n1192), .B(n1193), .Z(n1183) );
XNOR2_X1 U890 ( .A(G110), .B(n1123), .ZN(n1193) );
NAND2_X1 U891 ( .A1(G227), .A2(n1007), .ZN(n1123) );
XOR2_X1 U892 ( .A(KEYINPUT60), .B(KEYINPUT55), .Z(n1192) );
XNOR2_X1 U893 ( .A(KEYINPUT18), .B(n1127), .ZN(n1181) );
NAND2_X1 U894 ( .A1(n1194), .A2(n999), .ZN(n1175) );
INV_X1 U895 ( .A(n991), .ZN(n999) );
NOR3_X1 U896 ( .A1(n1172), .A2(G953), .A3(n1032), .ZN(n991) );
INV_X1 U897 ( .A(G952), .ZN(n1032) );
XOR2_X1 U898 ( .A(KEYINPUT47), .B(n1195), .Z(n1194) );
NOR4_X1 U899 ( .A1(G898), .A2(n1172), .A3(n1127), .A4(n1196), .ZN(n1195) );
XNOR2_X1 U900 ( .A(KEYINPUT30), .B(n1007), .ZN(n1196) );
AND2_X1 U901 ( .A1(G237), .A2(G234), .ZN(n1172) );
NOR2_X1 U902 ( .A1(n1031), .A2(n1030), .ZN(n1154) );
INV_X1 U903 ( .A(n1170), .ZN(n1030) );
NAND2_X1 U904 ( .A1(G214), .A2(n1197), .ZN(n1170) );
XNOR2_X1 U905 ( .A(KEYINPUT50), .B(n1198), .ZN(n1197) );
XOR2_X1 U906 ( .A(n1199), .B(n1043), .Z(n1031) );
NAND2_X1 U907 ( .A1(n1200), .A2(n1127), .ZN(n1043) );
XNOR2_X1 U908 ( .A(n1126), .B(KEYINPUT27), .ZN(n1200) );
XNOR2_X1 U909 ( .A(n1201), .B(n1202), .ZN(n1126) );
XOR2_X1 U910 ( .A(n1203), .B(n1204), .Z(n1202) );
NAND2_X1 U911 ( .A1(G224), .A2(n1007), .ZN(n1204) );
NAND2_X1 U912 ( .A1(n1205), .A2(KEYINPUT53), .ZN(n1203) );
XOR2_X1 U913 ( .A(n1206), .B(n1070), .Z(n1205) );
NAND2_X1 U914 ( .A1(n1207), .A2(n1208), .ZN(n1070) );
NAND2_X1 U915 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XNOR2_X1 U916 ( .A(G101), .B(KEYINPUT40), .ZN(n1209) );
NAND2_X1 U917 ( .A1(n1191), .A2(n1211), .ZN(n1207) );
XNOR2_X1 U918 ( .A(G101), .B(KEYINPUT42), .ZN(n1211) );
INV_X1 U919 ( .A(n1210), .ZN(n1191) );
XOR2_X1 U920 ( .A(G104), .B(n1212), .Z(n1210) );
INV_X1 U921 ( .A(G107), .ZN(n1212) );
NAND2_X1 U922 ( .A1(KEYINPUT43), .A2(n1073), .ZN(n1206) );
XNOR2_X1 U923 ( .A(n1178), .B(n1213), .ZN(n1073) );
NOR2_X1 U924 ( .A1(KEYINPUT9), .A2(n1214), .ZN(n1213) );
XOR2_X1 U925 ( .A(n1215), .B(G119), .Z(n1214) );
NAND2_X1 U926 ( .A1(KEYINPUT7), .A2(n1216), .ZN(n1215) );
XOR2_X1 U927 ( .A(n1057), .B(n1071), .Z(n1201) );
XNOR2_X1 U928 ( .A(n1217), .B(n1218), .ZN(n1071) );
XOR2_X1 U929 ( .A(KEYINPUT28), .B(G122), .Z(n1218) );
INV_X1 U930 ( .A(G110), .ZN(n1217) );
XNOR2_X1 U931 ( .A(G125), .B(n1107), .ZN(n1057) );
NAND2_X1 U932 ( .A1(KEYINPUT33), .A2(n1044), .ZN(n1199) );
NAND2_X1 U933 ( .A1(G210), .A2(n1198), .ZN(n1044) );
NAND2_X1 U934 ( .A1(n1219), .A2(n1127), .ZN(n1198) );
XOR2_X1 U935 ( .A(KEYINPUT62), .B(G237), .Z(n1219) );
INV_X1 U936 ( .A(n1037), .ZN(n1025) );
XNOR2_X1 U937 ( .A(n1220), .B(G472), .ZN(n1037) );
NAND2_X1 U938 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XNOR2_X1 U939 ( .A(KEYINPUT51), .B(n1127), .ZN(n1222) );
XOR2_X1 U940 ( .A(n1223), .B(n1224), .Z(n1221) );
XNOR2_X1 U941 ( .A(n1110), .B(n1189), .ZN(n1224) );
XNOR2_X1 U942 ( .A(n1111), .B(n1107), .ZN(n1189) );
XOR2_X1 U943 ( .A(n1225), .B(n1226), .Z(n1107) );
INV_X1 U944 ( .A(G101), .ZN(n1111) );
NAND2_X1 U945 ( .A1(n1227), .A2(G210), .ZN(n1110) );
XOR2_X1 U946 ( .A(n1228), .B(n1229), .Z(n1223) );
NOR2_X1 U947 ( .A1(KEYINPUT11), .A2(n1109), .ZN(n1229) );
XNOR2_X1 U948 ( .A(n1230), .B(n1231), .ZN(n1109) );
XOR2_X1 U949 ( .A(KEYINPUT15), .B(G119), .Z(n1231) );
XNOR2_X1 U950 ( .A(G113), .B(G116), .ZN(n1230) );
NAND2_X1 U951 ( .A1(n1232), .A2(n1108), .ZN(n1228) );
XNOR2_X1 U952 ( .A(n1060), .B(KEYINPUT5), .ZN(n1108) );
XOR2_X1 U953 ( .A(G131), .B(n1233), .Z(n1060) );
XNOR2_X1 U954 ( .A(n1234), .B(G134), .ZN(n1233) );
XNOR2_X1 U955 ( .A(KEYINPUT26), .B(KEYINPUT24), .ZN(n1232) );
NOR2_X1 U956 ( .A1(n1158), .A2(n1160), .ZN(n1005) );
INV_X1 U957 ( .A(n1176), .ZN(n1160) );
XOR2_X1 U958 ( .A(n1038), .B(KEYINPUT56), .Z(n1176) );
XOR2_X1 U959 ( .A(G478), .B(n1235), .Z(n1038) );
NOR2_X1 U960 ( .A1(n1087), .A2(G902), .ZN(n1235) );
AND2_X1 U961 ( .A1(n1236), .A2(n1237), .ZN(n1087) );
NAND2_X1 U962 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
XOR2_X1 U963 ( .A(KEYINPUT13), .B(n1240), .Z(n1236) );
NOR2_X1 U964 ( .A1(n1238), .A2(n1239), .ZN(n1240) );
NAND2_X1 U965 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
XNOR2_X1 U966 ( .A(G217), .B(KEYINPUT46), .ZN(n1241) );
XNOR2_X1 U967 ( .A(n1243), .B(n1244), .ZN(n1238) );
XNOR2_X1 U968 ( .A(n1216), .B(n1245), .ZN(n1244) );
XOR2_X1 U969 ( .A(G134), .B(G122), .Z(n1245) );
INV_X1 U970 ( .A(G116), .ZN(n1216) );
XNOR2_X1 U971 ( .A(G107), .B(n1225), .ZN(n1243) );
XOR2_X1 U972 ( .A(G128), .B(G143), .Z(n1225) );
NAND2_X1 U973 ( .A1(n1246), .A2(n1034), .ZN(n1158) );
NAND2_X1 U974 ( .A1(n1247), .A2(n1248), .ZN(n1034) );
XNOR2_X1 U975 ( .A(n1045), .B(KEYINPUT63), .ZN(n1246) );
NOR2_X1 U976 ( .A1(n1248), .A2(n1247), .ZN(n1045) );
AND2_X1 U977 ( .A1(n1249), .A2(n1127), .ZN(n1247) );
XNOR2_X1 U978 ( .A(n1095), .B(n1250), .ZN(n1249) );
INV_X1 U979 ( .A(n1094), .ZN(n1250) );
XNOR2_X1 U980 ( .A(n1251), .B(n1252), .ZN(n1094) );
XOR2_X1 U981 ( .A(G104), .B(n1253), .Z(n1252) );
NOR2_X1 U982 ( .A1(KEYINPUT3), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U983 ( .A(G140), .B(KEYINPUT4), .ZN(n1251) );
XNOR2_X1 U984 ( .A(n1255), .B(n1226), .ZN(n1095) );
XOR2_X1 U985 ( .A(n1256), .B(n1257), .Z(n1255) );
NOR2_X1 U986 ( .A1(KEYINPUT31), .A2(n1258), .ZN(n1257) );
NOR2_X1 U987 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U988 ( .A(KEYINPUT29), .B(n1261), .Z(n1260) );
AND2_X1 U989 ( .A1(n1169), .A2(n1262), .ZN(n1261) );
NOR2_X1 U990 ( .A1(n1169), .A2(n1262), .ZN(n1259) );
XNOR2_X1 U991 ( .A(n1263), .B(G143), .ZN(n1262) );
NAND2_X1 U992 ( .A1(n1227), .A2(G214), .ZN(n1263) );
NOR2_X1 U993 ( .A1(G953), .A2(G237), .ZN(n1227) );
INV_X1 U994 ( .A(G131), .ZN(n1169) );
NAND2_X1 U995 ( .A1(n1264), .A2(n1265), .ZN(n1256) );
NAND2_X1 U996 ( .A1(n1266), .A2(n1178), .ZN(n1265) );
INV_X1 U997 ( .A(G113), .ZN(n1178) );
NAND2_X1 U998 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
OR2_X1 U999 ( .A1(G122), .A2(KEYINPUT32), .ZN(n1268) );
NAND2_X1 U1000 ( .A1(G122), .A2(n1269), .ZN(n1264) );
NAND2_X1 U1001 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U1002 ( .A1(G113), .A2(n1267), .ZN(n1271) );
INV_X1 U1003 ( .A(KEYINPUT35), .ZN(n1267) );
INV_X1 U1004 ( .A(KEYINPUT32), .ZN(n1270) );
INV_X1 U1005 ( .A(G475), .ZN(n1248) );
XOR2_X1 U1006 ( .A(n1272), .B(n1041), .Z(n1026) );
NOR2_X1 U1007 ( .A1(n1083), .A2(G902), .ZN(n1041) );
XNOR2_X1 U1008 ( .A(n1273), .B(n1274), .ZN(n1083) );
XNOR2_X1 U1009 ( .A(G128), .B(n1254), .ZN(n1274) );
INV_X1 U1010 ( .A(G125), .ZN(n1254) );
XOR2_X1 U1011 ( .A(n1275), .B(n1276), .Z(n1273) );
XOR2_X1 U1012 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U1013 ( .A(KEYINPUT14), .B(G119), .Z(n1278) );
XOR2_X1 U1014 ( .A(KEYINPUT8), .B(KEYINPUT36), .Z(n1277) );
XOR2_X1 U1015 ( .A(n1279), .B(n1280), .Z(n1275) );
XOR2_X1 U1016 ( .A(n1226), .B(n1121), .Z(n1280) );
XOR2_X1 U1017 ( .A(G110), .B(G140), .Z(n1121) );
XOR2_X1 U1018 ( .A(G146), .B(KEYINPUT1), .Z(n1226) );
XOR2_X1 U1019 ( .A(n1281), .B(n1282), .Z(n1279) );
NOR2_X1 U1020 ( .A1(KEYINPUT44), .A2(n1234), .ZN(n1282) );
INV_X1 U1021 ( .A(G137), .ZN(n1234) );
NAND2_X1 U1022 ( .A1(n1242), .A2(G221), .ZN(n1281) );
AND2_X1 U1023 ( .A1(G234), .A2(n1007), .ZN(n1242) );
INV_X1 U1024 ( .A(G953), .ZN(n1007) );
NAND2_X1 U1025 ( .A1(KEYINPUT2), .A2(n1042), .ZN(n1272) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1179), .ZN(n1042) );
NAND2_X1 U1027 ( .A1(G234), .A2(n1127), .ZN(n1179) );
INV_X1 U1028 ( .A(G902), .ZN(n1127) );
endmodule


