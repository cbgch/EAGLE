//Key = 0010101110011100101101011111110111100111110101100101000000000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381;

XNOR2_X1 U763 ( .A(G107), .B(n1058), .ZN(G9) );
NOR2_X1 U764 ( .A1(n1059), .A2(n1060), .ZN(G75) );
NOR4_X1 U765 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
XOR2_X1 U766 ( .A(n1065), .B(KEYINPUT3), .Z(n1064) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U768 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
NAND2_X1 U769 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NAND3_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NAND2_X1 U771 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
NAND2_X1 U772 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND3_X1 U773 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NAND3_X1 U774 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1078) );
OR2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1066) );
NOR2_X1 U776 ( .A1(n1088), .A2(n1086), .ZN(n1063) );
NAND3_X1 U777 ( .A1(n1074), .A2(n1076), .A3(n1070), .ZN(n1086) );
NAND3_X1 U778 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1061) );
NAND3_X1 U779 ( .A1(n1068), .A2(n1092), .A3(n1070), .ZN(n1091) );
INV_X1 U780 ( .A(n1093), .ZN(n1070) );
NAND2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NAND2_X1 U782 ( .A1(n1076), .A2(n1096), .ZN(n1095) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U784 ( .A1(n1082), .A2(n1099), .ZN(n1098) );
NAND2_X1 U785 ( .A1(n1084), .A2(n1100), .ZN(n1097) );
NAND2_X1 U786 ( .A1(n1074), .A2(n1101), .ZN(n1094) );
AND2_X1 U787 ( .A1(n1082), .A2(n1084), .ZN(n1074) );
NOR3_X1 U788 ( .A1(n1102), .A2(G953), .A3(G952), .ZN(n1059) );
INV_X1 U789 ( .A(n1089), .ZN(n1102) );
NAND4_X1 U790 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1089) );
NOR4_X1 U791 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1106) );
NOR2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U793 ( .A(KEYINPUT56), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR3_X1 U795 ( .A1(KEYINPUT56), .A2(n1113), .A3(n1115), .ZN(n1109) );
XOR2_X1 U796 ( .A(KEYINPUT5), .B(n1116), .Z(n1108) );
NAND3_X1 U797 ( .A1(n1117), .A2(n1118), .A3(n1119), .ZN(n1107) );
XOR2_X1 U798 ( .A(n1120), .B(KEYINPUT35), .Z(n1119) );
NAND2_X1 U799 ( .A1(n1115), .A2(n1113), .ZN(n1118) );
NOR2_X1 U800 ( .A1(n1121), .A2(KEYINPUT53), .ZN(n1115) );
NOR3_X1 U801 ( .A1(n1122), .A2(n1085), .A3(n1075), .ZN(n1105) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(n1104) );
XOR2_X1 U803 ( .A(n1125), .B(KEYINPUT14), .Z(n1124) );
NAND2_X1 U804 ( .A1(KEYINPUT39), .A2(n1126), .ZN(n1123) );
NOR2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1103) );
AND2_X1 U806 ( .A1(n1129), .A2(G469), .ZN(n1128) );
XOR2_X1 U807 ( .A(n1130), .B(n1131), .Z(G72) );
XOR2_X1 U808 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U809 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND2_X1 U810 ( .A1(G900), .A2(G227), .ZN(n1135) );
INV_X1 U811 ( .A(n1136), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NAND2_X1 U813 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U814 ( .A(G953), .B(KEYINPUT32), .ZN(n1139) );
XOR2_X1 U815 ( .A(n1141), .B(n1142), .Z(n1137) );
NOR2_X1 U816 ( .A1(KEYINPUT54), .A2(n1143), .ZN(n1141) );
NOR2_X1 U817 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U818 ( .A(KEYINPUT52), .B(n1146), .Z(n1145) );
NOR2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XNOR2_X1 U820 ( .A(G128), .B(n1149), .ZN(n1147) );
NOR2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
XOR2_X1 U822 ( .A(G128), .B(n1149), .Z(n1151) );
NOR2_X1 U823 ( .A1(n1152), .A2(G953), .ZN(n1130) );
NOR2_X1 U824 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XOR2_X1 U825 ( .A(KEYINPUT51), .B(n1155), .Z(n1154) );
XOR2_X1 U826 ( .A(n1156), .B(n1157), .Z(G69) );
NOR2_X1 U827 ( .A1(n1158), .A2(n1136), .ZN(n1157) );
XOR2_X1 U828 ( .A(G953), .B(KEYINPUT4), .Z(n1136) );
AND2_X1 U829 ( .A1(G224), .A2(G898), .ZN(n1158) );
NAND2_X1 U830 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
NAND2_X1 U831 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U832 ( .A(KEYINPUT19), .B(n1163), .Z(n1159) );
NOR3_X1 U833 ( .A1(n1162), .A2(n1164), .A3(n1161), .ZN(n1163) );
AND2_X1 U834 ( .A1(n1090), .A2(n1165), .ZN(n1161) );
NAND2_X1 U835 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U836 ( .A(n1168), .B(KEYINPUT41), .Z(n1166) );
NAND2_X1 U837 ( .A1(n1169), .A2(n1058), .ZN(n1168) );
INV_X1 U838 ( .A(n1170), .ZN(n1169) );
XNOR2_X1 U839 ( .A(n1171), .B(n1172), .ZN(n1162) );
XNOR2_X1 U840 ( .A(n1173), .B(KEYINPUT58), .ZN(n1172) );
NAND2_X1 U841 ( .A1(KEYINPUT26), .A2(n1174), .ZN(n1173) );
XOR2_X1 U842 ( .A(n1175), .B(n1176), .Z(n1171) );
NOR2_X1 U843 ( .A1(n1177), .A2(n1178), .ZN(G66) );
XNOR2_X1 U844 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U845 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U846 ( .A1(n1177), .A2(n1183), .ZN(G63) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND3_X1 U848 ( .A1(G902), .A2(G478), .A3(n1186), .ZN(n1184) );
XOR2_X1 U849 ( .A(n1062), .B(KEYINPUT63), .Z(n1186) );
NOR2_X1 U850 ( .A1(n1177), .A2(n1187), .ZN(G60) );
XNOR2_X1 U851 ( .A(n1188), .B(n1189), .ZN(n1187) );
NOR2_X1 U852 ( .A1(n1190), .A2(n1182), .ZN(n1189) );
XOR2_X1 U853 ( .A(G104), .B(n1191), .Z(G6) );
NOR2_X1 U854 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NOR2_X1 U855 ( .A1(n1177), .A2(n1194), .ZN(G57) );
NOR2_X1 U856 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U857 ( .A(KEYINPUT10), .B(n1197), .Z(n1196) );
NOR2_X1 U858 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
AND2_X1 U859 ( .A1(n1199), .A2(n1198), .ZN(n1195) );
XOR2_X1 U860 ( .A(n1200), .B(G101), .Z(n1198) );
NAND2_X1 U861 ( .A1(KEYINPUT34), .A2(n1201), .ZN(n1200) );
XNOR2_X1 U862 ( .A(n1202), .B(n1203), .ZN(n1199) );
XNOR2_X1 U863 ( .A(n1204), .B(n1150), .ZN(n1203) );
INV_X1 U864 ( .A(n1148), .ZN(n1150) );
XNOR2_X1 U865 ( .A(n1205), .B(n1206), .ZN(n1202) );
NOR2_X1 U866 ( .A1(KEYINPUT48), .A2(n1207), .ZN(n1206) );
NOR3_X1 U867 ( .A1(n1182), .A2(KEYINPUT30), .A3(n1208), .ZN(n1205) );
NOR3_X1 U868 ( .A1(n1209), .A2(n1177), .A3(n1210), .ZN(G54) );
NOR3_X1 U869 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
XOR2_X1 U870 ( .A(n1214), .B(n1215), .Z(n1211) );
NOR2_X1 U871 ( .A1(KEYINPUT42), .A2(n1216), .ZN(n1215) );
NOR2_X1 U872 ( .A1(n1217), .A2(n1218), .ZN(n1209) );
XOR2_X1 U873 ( .A(n1214), .B(n1219), .Z(n1218) );
NOR2_X1 U874 ( .A1(KEYINPUT42), .A2(n1220), .ZN(n1219) );
NOR2_X1 U875 ( .A1(n1182), .A2(n1221), .ZN(n1214) );
INV_X1 U876 ( .A(G469), .ZN(n1221) );
NOR2_X1 U877 ( .A1(n1212), .A2(n1213), .ZN(n1217) );
INV_X1 U878 ( .A(KEYINPUT46), .ZN(n1213) );
NOR2_X1 U879 ( .A1(n1177), .A2(n1222), .ZN(G51) );
XOR2_X1 U880 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U881 ( .A(n1225), .B(n1226), .Z(n1224) );
NOR2_X1 U882 ( .A1(n1126), .A2(n1182), .ZN(n1226) );
NAND2_X1 U883 ( .A1(G902), .A2(n1062), .ZN(n1182) );
NAND3_X1 U884 ( .A1(n1167), .A2(n1155), .A3(n1227), .ZN(n1062) );
NOR3_X1 U885 ( .A1(n1170), .A2(n1228), .A3(n1153), .ZN(n1227) );
NAND4_X1 U886 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1153) );
XOR2_X1 U887 ( .A(n1058), .B(KEYINPUT23), .Z(n1228) );
NAND3_X1 U888 ( .A1(n1233), .A2(n1234), .A3(n1084), .ZN(n1058) );
NAND3_X1 U889 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1170) );
NAND2_X1 U890 ( .A1(n1238), .A2(n1101), .ZN(n1237) );
XOR2_X1 U891 ( .A(n1193), .B(KEYINPUT29), .Z(n1238) );
NAND4_X1 U892 ( .A1(n1239), .A2(n1084), .A3(n1100), .A4(n1240), .ZN(n1193) );
AND3_X1 U893 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1155) );
NAND3_X1 U894 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
INV_X1 U895 ( .A(n1247), .ZN(n1246) );
NAND2_X1 U896 ( .A1(n1248), .A2(n1249), .ZN(n1245) );
OR2_X1 U897 ( .A1(n1087), .A2(KEYINPUT13), .ZN(n1248) );
NAND3_X1 U898 ( .A1(n1250), .A2(n1088), .A3(n1100), .ZN(n1244) );
NAND2_X1 U899 ( .A1(KEYINPUT13), .A2(n1233), .ZN(n1250) );
AND4_X1 U900 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1167) );
NAND3_X1 U901 ( .A1(n1233), .A2(n1099), .A3(n1255), .ZN(n1251) );
NAND3_X1 U902 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1225) );
NAND2_X1 U903 ( .A1(KEYINPUT55), .A2(n1259), .ZN(n1258) );
OR3_X1 U904 ( .A1(n1260), .A2(KEYINPUT55), .A3(G125), .ZN(n1257) );
NAND2_X1 U905 ( .A1(G125), .A2(n1260), .ZN(n1256) );
NAND2_X1 U906 ( .A1(KEYINPUT8), .A2(n1204), .ZN(n1260) );
NOR2_X1 U907 ( .A1(n1090), .A2(G952), .ZN(n1177) );
XOR2_X1 U908 ( .A(n1229), .B(n1261), .Z(G48) );
XOR2_X1 U909 ( .A(KEYINPUT45), .B(G146), .Z(n1261) );
NAND3_X1 U910 ( .A1(n1239), .A2(n1101), .A3(n1262), .ZN(n1229) );
XNOR2_X1 U911 ( .A(G143), .B(n1230), .ZN(G45) );
NAND4_X1 U912 ( .A1(n1263), .A2(n1264), .A3(n1099), .A4(n1265), .ZN(n1230) );
NOR3_X1 U913 ( .A1(n1266), .A2(n1192), .A3(n1249), .ZN(n1265) );
INV_X1 U914 ( .A(n1101), .ZN(n1192) );
XNOR2_X1 U915 ( .A(G140), .B(n1231), .ZN(G42) );
NAND4_X1 U916 ( .A1(n1076), .A2(n1267), .A3(n1080), .A4(n1239), .ZN(n1231) );
XNOR2_X1 U917 ( .A(G137), .B(n1232), .ZN(G39) );
NAND3_X1 U918 ( .A1(n1262), .A2(n1068), .A3(n1076), .ZN(n1232) );
XOR2_X1 U919 ( .A(G134), .B(n1268), .Z(G36) );
NOR3_X1 U920 ( .A1(n1247), .A2(n1269), .A3(n1087), .ZN(n1268) );
INV_X1 U921 ( .A(n1233), .ZN(n1087) );
XNOR2_X1 U922 ( .A(n1100), .B(KEYINPUT0), .ZN(n1269) );
XOR2_X1 U923 ( .A(G131), .B(n1270), .Z(G33) );
NOR4_X1 U924 ( .A1(KEYINPUT1), .A2(n1249), .A3(n1088), .A4(n1247), .ZN(n1270) );
NAND3_X1 U925 ( .A1(n1099), .A2(n1263), .A3(n1076), .ZN(n1247) );
NOR2_X1 U926 ( .A1(n1271), .A2(n1075), .ZN(n1076) );
INV_X1 U927 ( .A(n1239), .ZN(n1088) );
XNOR2_X1 U928 ( .A(G128), .B(n1241), .ZN(G30) );
NAND3_X1 U929 ( .A1(n1233), .A2(n1101), .A3(n1262), .ZN(n1241) );
AND2_X1 U930 ( .A1(n1267), .A2(n1272), .ZN(n1262) );
NOR3_X1 U931 ( .A1(n1273), .A2(n1274), .A3(n1249), .ZN(n1267) );
INV_X1 U932 ( .A(n1100), .ZN(n1249) );
XNOR2_X1 U933 ( .A(G101), .B(n1275), .ZN(G3) );
NAND2_X1 U934 ( .A1(KEYINPUT37), .A2(n1276), .ZN(n1275) );
INV_X1 U935 ( .A(n1235), .ZN(n1276) );
NAND3_X1 U936 ( .A1(n1234), .A2(n1099), .A3(n1068), .ZN(n1235) );
NAND2_X1 U937 ( .A1(n1277), .A2(n1278), .ZN(G27) );
NAND2_X1 U938 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XOR2_X1 U939 ( .A(n1242), .B(KEYINPUT24), .Z(n1279) );
NAND2_X1 U940 ( .A1(n1281), .A2(G125), .ZN(n1277) );
XNOR2_X1 U941 ( .A(KEYINPUT11), .B(n1242), .ZN(n1281) );
NAND4_X1 U942 ( .A1(n1082), .A2(n1101), .A3(n1239), .A4(n1282), .ZN(n1242) );
NOR3_X1 U943 ( .A1(n1272), .A2(n1274), .A3(n1273), .ZN(n1282) );
INV_X1 U944 ( .A(n1263), .ZN(n1273) );
NAND2_X1 U945 ( .A1(n1093), .A2(n1283), .ZN(n1263) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1284), .A4(n1140), .ZN(n1283) );
INV_X1 U947 ( .A(G900), .ZN(n1140) );
INV_X1 U948 ( .A(n1081), .ZN(n1274) );
XNOR2_X1 U949 ( .A(G122), .B(n1252), .ZN(G24) );
NAND4_X1 U950 ( .A1(n1285), .A2(n1255), .A3(n1084), .A4(n1264), .ZN(n1252) );
XNOR2_X1 U951 ( .A(G119), .B(n1253), .ZN(G21) );
NAND4_X1 U952 ( .A1(n1068), .A2(n1255), .A3(n1272), .A4(n1081), .ZN(n1253) );
XNOR2_X1 U953 ( .A(G116), .B(n1286), .ZN(G18) );
NAND3_X1 U954 ( .A1(n1287), .A2(n1233), .A3(n1255), .ZN(n1286) );
NOR2_X1 U955 ( .A1(n1285), .A2(n1288), .ZN(n1233) );
XOR2_X1 U956 ( .A(n1099), .B(KEYINPUT9), .Z(n1287) );
XNOR2_X1 U957 ( .A(G113), .B(n1254), .ZN(G15) );
NAND3_X1 U958 ( .A1(n1255), .A2(n1099), .A3(n1239), .ZN(n1254) );
NOR2_X1 U959 ( .A1(n1264), .A2(n1266), .ZN(n1239) );
NAND2_X1 U960 ( .A1(n1289), .A2(n1290), .ZN(n1099) );
OR3_X1 U961 ( .A1(n1081), .A2(n1080), .A3(KEYINPUT20), .ZN(n1290) );
NAND2_X1 U962 ( .A1(KEYINPUT20), .A2(n1084), .ZN(n1289) );
NOR2_X1 U963 ( .A1(n1081), .A2(n1272), .ZN(n1084) );
AND3_X1 U964 ( .A1(n1101), .A2(n1240), .A3(n1082), .ZN(n1255) );
AND2_X1 U965 ( .A1(n1083), .A2(n1291), .ZN(n1082) );
NAND2_X1 U966 ( .A1(n1292), .A2(n1293), .ZN(G12) );
NAND2_X1 U967 ( .A1(G110), .A2(n1236), .ZN(n1293) );
XOR2_X1 U968 ( .A(KEYINPUT49), .B(n1294), .Z(n1292) );
NOR2_X1 U969 ( .A1(G110), .A2(n1236), .ZN(n1294) );
NAND4_X1 U970 ( .A1(n1068), .A2(n1234), .A3(n1080), .A4(n1081), .ZN(n1236) );
NAND2_X1 U971 ( .A1(n1295), .A2(n1296), .ZN(n1081) );
NAND2_X1 U972 ( .A1(n1121), .A2(n1181), .ZN(n1296) );
XOR2_X1 U973 ( .A(n1297), .B(KEYINPUT59), .Z(n1295) );
NAND2_X1 U974 ( .A1(n1113), .A2(n1114), .ZN(n1297) );
INV_X1 U975 ( .A(n1121), .ZN(n1114) );
NOR2_X1 U976 ( .A1(n1298), .A2(G902), .ZN(n1121) );
INV_X1 U977 ( .A(n1179), .ZN(n1298) );
XNOR2_X1 U978 ( .A(n1299), .B(n1300), .ZN(n1179) );
NOR2_X1 U979 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
AND2_X1 U980 ( .A1(KEYINPUT60), .A2(n1303), .ZN(n1302) );
NOR2_X1 U981 ( .A1(KEYINPUT15), .A2(n1303), .ZN(n1301) );
XOR2_X1 U982 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U983 ( .A(G128), .B(G110), .Z(n1305) );
XNOR2_X1 U984 ( .A(n1306), .B(n1307), .ZN(n1304) );
NAND2_X1 U985 ( .A1(KEYINPUT40), .A2(n1308), .ZN(n1307) );
NAND2_X1 U986 ( .A1(KEYINPUT27), .A2(n1309), .ZN(n1306) );
XOR2_X1 U987 ( .A(G146), .B(n1142), .Z(n1309) );
XNOR2_X1 U988 ( .A(n1310), .B(n1311), .ZN(n1299) );
INV_X1 U989 ( .A(G137), .ZN(n1311) );
NAND2_X1 U990 ( .A1(G221), .A2(n1312), .ZN(n1310) );
INV_X1 U991 ( .A(n1181), .ZN(n1113) );
NAND2_X1 U992 ( .A1(G217), .A2(n1313), .ZN(n1181) );
INV_X1 U993 ( .A(n1272), .ZN(n1080) );
XNOR2_X1 U994 ( .A(n1117), .B(KEYINPUT57), .ZN(n1272) );
XNOR2_X1 U995 ( .A(n1314), .B(n1208), .ZN(n1117) );
INV_X1 U996 ( .A(G472), .ZN(n1208) );
NAND2_X1 U997 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U998 ( .A(n1317), .B(n1318), .Z(n1315) );
XNOR2_X1 U999 ( .A(n1319), .B(n1207), .ZN(n1318) );
XNOR2_X1 U1000 ( .A(G113), .B(n1320), .ZN(n1207) );
XNOR2_X1 U1001 ( .A(n1308), .B(G116), .ZN(n1320) );
INV_X1 U1002 ( .A(G119), .ZN(n1308) );
XOR2_X1 U1003 ( .A(n1321), .B(n1201), .Z(n1317) );
AND3_X1 U1004 ( .A1(n1322), .A2(n1090), .A3(G210), .ZN(n1201) );
NAND2_X1 U1005 ( .A1(KEYINPUT43), .A2(n1204), .ZN(n1321) );
AND3_X1 U1006 ( .A1(n1101), .A2(n1240), .A3(n1100), .ZN(n1234) );
NOR2_X1 U1007 ( .A1(n1083), .A2(n1085), .ZN(n1100) );
INV_X1 U1008 ( .A(n1291), .ZN(n1085) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1313), .ZN(n1291) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1316), .ZN(n1313) );
NOR2_X1 U1011 ( .A1(n1122), .A2(n1323), .ZN(n1083) );
AND2_X1 U1012 ( .A1(n1324), .A2(n1129), .ZN(n1323) );
XNOR2_X1 U1013 ( .A(G469), .B(KEYINPUT61), .ZN(n1324) );
NOR2_X1 U1014 ( .A1(n1129), .A2(G469), .ZN(n1122) );
NAND2_X1 U1015 ( .A1(n1325), .A2(n1316), .ZN(n1129) );
XNOR2_X1 U1016 ( .A(n1212), .B(n1216), .ZN(n1325) );
INV_X1 U1017 ( .A(n1220), .ZN(n1216) );
XNOR2_X1 U1018 ( .A(n1326), .B(n1327), .ZN(n1220) );
XOR2_X1 U1019 ( .A(G140), .B(G110), .Z(n1327) );
NAND2_X1 U1020 ( .A1(G227), .A2(n1090), .ZN(n1326) );
XOR2_X1 U1021 ( .A(n1328), .B(n1329), .Z(n1212) );
XOR2_X1 U1022 ( .A(G104), .B(n1330), .Z(n1329) );
XOR2_X1 U1023 ( .A(n1319), .B(n1149), .Z(n1328) );
XNOR2_X1 U1024 ( .A(G101), .B(n1148), .ZN(n1319) );
XNOR2_X1 U1025 ( .A(n1331), .B(n1332), .ZN(n1148) );
XNOR2_X1 U1026 ( .A(G134), .B(G137), .ZN(n1331) );
NAND2_X1 U1027 ( .A1(n1093), .A2(n1333), .ZN(n1240) );
NAND3_X1 U1028 ( .A1(G902), .A2(n1284), .A3(n1164), .ZN(n1333) );
NOR2_X1 U1029 ( .A1(n1090), .A2(G898), .ZN(n1164) );
NAND3_X1 U1030 ( .A1(n1284), .A2(n1090), .A3(G952), .ZN(n1093) );
NAND2_X1 U1031 ( .A1(G237), .A2(G234), .ZN(n1284) );
NOR2_X1 U1032 ( .A1(n1073), .A2(n1075), .ZN(n1101) );
AND2_X1 U1033 ( .A1(G214), .A2(n1334), .ZN(n1075) );
INV_X1 U1034 ( .A(n1271), .ZN(n1073) );
XOR2_X1 U1035 ( .A(n1125), .B(n1126), .Z(n1271) );
NAND2_X1 U1036 ( .A1(G210), .A2(n1334), .ZN(n1126) );
NAND2_X1 U1037 ( .A1(n1335), .A2(n1316), .ZN(n1334) );
XNOR2_X1 U1038 ( .A(KEYINPUT21), .B(n1322), .ZN(n1335) );
NAND2_X1 U1039 ( .A1(n1336), .A2(n1316), .ZN(n1125) );
XOR2_X1 U1040 ( .A(n1223), .B(n1337), .Z(n1336) );
XOR2_X1 U1041 ( .A(KEYINPUT22), .B(n1338), .Z(n1337) );
NOR2_X1 U1042 ( .A1(KEYINPUT44), .A2(n1339), .ZN(n1338) );
XNOR2_X1 U1043 ( .A(G125), .B(n1259), .ZN(n1339) );
INV_X1 U1044 ( .A(n1204), .ZN(n1259) );
XNOR2_X1 U1045 ( .A(n1340), .B(G128), .ZN(n1204) );
NAND2_X1 U1046 ( .A1(n1341), .A2(KEYINPUT12), .ZN(n1340) );
XOR2_X1 U1047 ( .A(n1342), .B(G143), .Z(n1341) );
NAND2_X1 U1048 ( .A1(KEYINPUT2), .A2(n1343), .ZN(n1342) );
XOR2_X1 U1049 ( .A(KEYINPUT36), .B(G146), .Z(n1343) );
XOR2_X1 U1050 ( .A(n1344), .B(n1345), .Z(n1223) );
AND2_X1 U1051 ( .A1(n1090), .A2(G224), .ZN(n1345) );
NAND2_X1 U1052 ( .A1(n1346), .A2(n1347), .ZN(n1344) );
NAND2_X1 U1053 ( .A1(n1348), .A2(n1176), .ZN(n1347) );
XOR2_X1 U1054 ( .A(n1349), .B(KEYINPUT50), .Z(n1346) );
OR2_X1 U1055 ( .A1(n1176), .A2(n1348), .ZN(n1349) );
XOR2_X1 U1056 ( .A(n1175), .B(n1174), .Z(n1348) );
XOR2_X1 U1057 ( .A(n1350), .B(n1351), .Z(n1174) );
XNOR2_X1 U1058 ( .A(G119), .B(n1352), .ZN(n1351) );
NAND2_X1 U1059 ( .A1(KEYINPUT28), .A2(G113), .ZN(n1352) );
NAND2_X1 U1060 ( .A1(KEYINPUT33), .A2(G116), .ZN(n1350) );
XNOR2_X1 U1061 ( .A(G101), .B(n1353), .ZN(n1175) );
NOR2_X1 U1062 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NOR3_X1 U1063 ( .A1(KEYINPUT7), .A2(G107), .A3(n1356), .ZN(n1355) );
NOR2_X1 U1064 ( .A1(n1357), .A2(n1358), .ZN(n1354) );
INV_X1 U1065 ( .A(KEYINPUT7), .ZN(n1358) );
XNOR2_X1 U1066 ( .A(G107), .B(n1356), .ZN(n1357) );
XNOR2_X1 U1067 ( .A(n1359), .B(G110), .ZN(n1176) );
NAND2_X1 U1068 ( .A1(KEYINPUT6), .A2(n1360), .ZN(n1359) );
NOR2_X1 U1069 ( .A1(n1264), .A2(n1285), .ZN(n1068) );
INV_X1 U1070 ( .A(n1266), .ZN(n1285) );
XNOR2_X1 U1071 ( .A(n1120), .B(KEYINPUT38), .ZN(n1266) );
XNOR2_X1 U1072 ( .A(n1361), .B(n1190), .ZN(n1120) );
INV_X1 U1073 ( .A(G475), .ZN(n1190) );
NAND2_X1 U1074 ( .A1(n1362), .A2(n1188), .ZN(n1361) );
NAND2_X1 U1075 ( .A1(n1363), .A2(n1364), .ZN(n1188) );
NAND2_X1 U1076 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XOR2_X1 U1077 ( .A(n1367), .B(KEYINPUT47), .Z(n1363) );
OR2_X1 U1078 ( .A1(n1366), .A2(n1365), .ZN(n1367) );
XNOR2_X1 U1079 ( .A(n1368), .B(n1369), .ZN(n1365) );
XNOR2_X1 U1080 ( .A(G113), .B(n1356), .ZN(n1369) );
INV_X1 U1081 ( .A(G104), .ZN(n1356) );
NAND2_X1 U1082 ( .A1(KEYINPUT31), .A2(n1360), .ZN(n1368) );
XNOR2_X1 U1083 ( .A(n1370), .B(n1371), .ZN(n1366) );
XOR2_X1 U1084 ( .A(n1149), .B(n1142), .Z(n1371) );
XNOR2_X1 U1085 ( .A(G140), .B(n1280), .ZN(n1142) );
INV_X1 U1086 ( .A(G125), .ZN(n1280) );
XOR2_X1 U1087 ( .A(G143), .B(G146), .Z(n1149) );
XOR2_X1 U1088 ( .A(n1372), .B(n1373), .Z(n1370) );
NOR2_X1 U1089 ( .A1(KEYINPUT17), .A2(n1332), .ZN(n1373) );
XOR2_X1 U1090 ( .A(G131), .B(KEYINPUT16), .Z(n1332) );
NAND3_X1 U1091 ( .A1(n1322), .A2(n1090), .A3(G214), .ZN(n1372) );
INV_X1 U1092 ( .A(G237), .ZN(n1322) );
XNOR2_X1 U1093 ( .A(KEYINPUT62), .B(n1316), .ZN(n1362) );
INV_X1 U1094 ( .A(n1288), .ZN(n1264) );
NOR2_X1 U1095 ( .A1(n1116), .A2(n1127), .ZN(n1288) );
AND2_X1 U1096 ( .A1(n1374), .A2(G478), .ZN(n1127) );
NOR2_X1 U1097 ( .A1(n1374), .A2(G478), .ZN(n1116) );
NAND2_X1 U1098 ( .A1(n1185), .A2(n1316), .ZN(n1374) );
INV_X1 U1099 ( .A(G902), .ZN(n1316) );
XOR2_X1 U1100 ( .A(n1375), .B(n1376), .Z(n1185) );
XNOR2_X1 U1101 ( .A(n1360), .B(n1377), .ZN(n1376) );
XOR2_X1 U1102 ( .A(G143), .B(G134), .Z(n1377) );
INV_X1 U1103 ( .A(G122), .ZN(n1360) );
XOR2_X1 U1104 ( .A(n1378), .B(n1330), .Z(n1375) );
XOR2_X1 U1105 ( .A(G107), .B(G128), .Z(n1330) );
XNOR2_X1 U1106 ( .A(n1379), .B(n1380), .ZN(n1378) );
NAND2_X1 U1107 ( .A1(KEYINPUT25), .A2(n1381), .ZN(n1380) );
INV_X1 U1108 ( .A(G116), .ZN(n1381) );
NAND3_X1 U1109 ( .A1(G217), .A2(n1312), .A3(KEYINPUT18), .ZN(n1379) );
AND2_X1 U1110 ( .A1(G234), .A2(n1090), .ZN(n1312) );
INV_X1 U1111 ( .A(G953), .ZN(n1090) );
endmodule


