//Key = 0010000111011100000001010011111010011101001001000011010110010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287;

XNOR2_X1 U712 ( .A(G107), .B(n985), .ZN(G9) );
NOR2_X1 U713 ( .A1(n986), .A2(n987), .ZN(G75) );
NOR4_X1 U714 ( .A1(n988), .A2(n989), .A3(G953), .A4(n990), .ZN(n987) );
NOR3_X1 U715 ( .A1(n991), .A2(n992), .A3(n993), .ZN(n989) );
NOR2_X1 U716 ( .A1(n994), .A2(n995), .ZN(n992) );
NAND3_X1 U717 ( .A1(n996), .A2(n997), .A3(n998), .ZN(n988) );
NAND2_X1 U718 ( .A1(n999), .A2(n1000), .ZN(n997) );
NAND2_X1 U719 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NAND3_X1 U720 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
NAND2_X1 U721 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NAND2_X1 U722 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
OR2_X1 U723 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NAND2_X1 U724 ( .A1(n1012), .A2(n1013), .ZN(n1006) );
NAND2_X1 U725 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND2_X1 U726 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U727 ( .A1(n1018), .A2(n1019), .ZN(n1001) );
NAND2_X1 U728 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
OR2_X1 U729 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
INV_X1 U730 ( .A(n991), .ZN(n1018) );
NAND3_X1 U731 ( .A1(n1008), .A2(n1012), .A3(n1005), .ZN(n991) );
INV_X1 U732 ( .A(n1024), .ZN(n1005) );
XOR2_X1 U733 ( .A(KEYINPUT22), .B(G952), .Z(n996) );
NOR3_X1 U734 ( .A1(n1025), .A2(G953), .A3(n990), .ZN(n986) );
AND4_X1 U735 ( .A1(n1026), .A2(n1012), .A3(n1027), .A4(n1028), .ZN(n990) );
NOR4_X1 U736 ( .A1(n1029), .A2(n1030), .A3(n1016), .A4(n1031), .ZN(n1028) );
XNOR2_X1 U737 ( .A(n1032), .B(KEYINPUT26), .ZN(n1031) );
INV_X1 U738 ( .A(n1033), .ZN(n1030) );
NOR2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1029) );
NOR2_X1 U740 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
AND2_X1 U741 ( .A1(n1038), .A2(KEYINPUT37), .ZN(n1037) );
NOR2_X1 U742 ( .A1(n1039), .A2(n1040), .ZN(n1036) );
NOR2_X1 U743 ( .A1(n1038), .A2(KEYINPUT2), .ZN(n1039) );
AND4_X1 U744 ( .A1(G475), .A2(n1038), .A3(KEYINPUT2), .A4(KEYINPUT37), .ZN(n1034) );
NOR2_X1 U745 ( .A1(n1041), .A2(n1042), .ZN(n1027) );
XOR2_X1 U746 ( .A(KEYINPUT1), .B(n1043), .Z(n1042) );
XNOR2_X1 U747 ( .A(G478), .B(n1044), .ZN(n1041) );
XOR2_X1 U748 ( .A(n1045), .B(KEYINPUT17), .Z(n1026) );
XOR2_X1 U749 ( .A(KEYINPUT4), .B(G952), .Z(n1025) );
XOR2_X1 U750 ( .A(n1046), .B(n1047), .Z(G72) );
NOR2_X1 U751 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1046) );
NAND2_X1 U754 ( .A1(n1054), .A2(n1049), .ZN(n1053) );
XNOR2_X1 U755 ( .A(n1055), .B(n1056), .ZN(n1054) );
NOR2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND3_X1 U757 ( .A1(G900), .A2(n1055), .A3(G953), .ZN(n1052) );
NAND3_X1 U758 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1055) );
NAND2_X1 U759 ( .A1(KEYINPUT25), .A2(n1062), .ZN(n1061) );
NAND3_X1 U760 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1060) );
INV_X1 U761 ( .A(KEYINPUT25), .ZN(n1064) );
OR2_X1 U762 ( .A1(n1065), .A2(n1063), .ZN(n1059) );
NOR2_X1 U763 ( .A1(KEYINPUT6), .A2(n1062), .ZN(n1063) );
XNOR2_X1 U764 ( .A(n1066), .B(n1067), .ZN(n1062) );
NAND2_X1 U765 ( .A1(KEYINPUT23), .A2(n1068), .ZN(n1066) );
XOR2_X1 U766 ( .A(G134), .B(n1069), .Z(n1068) );
NAND2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(G69) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1049), .ZN(n1071) );
XNOR2_X1 U769 ( .A(n1073), .B(n1074), .ZN(n1072) );
NOR2_X1 U770 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
XOR2_X1 U771 ( .A(n1077), .B(KEYINPUT16), .Z(n1075) );
NAND2_X1 U772 ( .A1(n1078), .A2(G953), .ZN(n1070) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U774 ( .A1(n1073), .A2(G224), .ZN(n1080) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1079) );
INV_X1 U776 ( .A(n1073), .ZN(n1082) );
NOR3_X1 U777 ( .A1(KEYINPUT49), .A2(n1083), .A3(n1084), .ZN(n1073) );
XNOR2_X1 U778 ( .A(n1085), .B(n1086), .ZN(n1084) );
NAND2_X1 U779 ( .A1(KEYINPUT8), .A2(n1087), .ZN(n1085) );
NAND2_X1 U780 ( .A1(G898), .A2(G224), .ZN(n1081) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(G66) );
XOR2_X1 U782 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR2_X1 U784 ( .A1(n1088), .A2(n1094), .ZN(G63) );
XOR2_X1 U785 ( .A(n1095), .B(n1096), .Z(n1094) );
XOR2_X1 U786 ( .A(n1097), .B(KEYINPUT7), .Z(n1095) );
NAND2_X1 U787 ( .A1(n1092), .A2(G478), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1088), .A2(n1098), .ZN(G60) );
NOR3_X1 U789 ( .A1(n1038), .A2(n1099), .A3(n1100), .ZN(n1098) );
AND3_X1 U790 ( .A1(n1101), .A2(G475), .A3(n1092), .ZN(n1100) );
NOR2_X1 U791 ( .A1(n1102), .A2(n1101), .ZN(n1099) );
NOR2_X1 U792 ( .A1(n998), .A2(n1040), .ZN(n1102) );
NAND2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(G6) );
OR2_X1 U794 ( .A1(n1105), .A2(G104), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1106), .B(KEYINPUT44), .Z(n1103) );
NAND2_X1 U796 ( .A1(G104), .A2(n1105), .ZN(n1106) );
NOR3_X1 U797 ( .A1(n1088), .A2(n1107), .A3(n1108), .ZN(G57) );
NOR2_X1 U798 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
XNOR2_X1 U799 ( .A(n1111), .B(KEYINPUT29), .ZN(n1110) );
NOR2_X1 U800 ( .A1(G101), .A2(n1112), .ZN(n1107) );
XNOR2_X1 U801 ( .A(n1113), .B(n1114), .ZN(n1112) );
XOR2_X1 U802 ( .A(KEYINPUT30), .B(KEYINPUT19), .Z(n1114) );
INV_X1 U803 ( .A(n1111), .ZN(n1113) );
XNOR2_X1 U804 ( .A(n1115), .B(n1116), .ZN(n1111) );
XNOR2_X1 U805 ( .A(n1117), .B(n1118), .ZN(n1116) );
NAND2_X1 U806 ( .A1(n1092), .A2(G472), .ZN(n1117) );
XNOR2_X1 U807 ( .A(n1119), .B(n1120), .ZN(n1115) );
NAND2_X1 U808 ( .A1(n1121), .A2(KEYINPUT12), .ZN(n1119) );
XNOR2_X1 U809 ( .A(n1122), .B(KEYINPUT54), .ZN(n1121) );
NOR2_X1 U810 ( .A1(n1088), .A2(n1123), .ZN(G54) );
XNOR2_X1 U811 ( .A(n1124), .B(n1125), .ZN(n1123) );
XOR2_X1 U812 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U813 ( .A(n1128), .B(n1129), .Z(n1127) );
XNOR2_X1 U814 ( .A(n1130), .B(n1067), .ZN(n1129) );
NAND2_X1 U815 ( .A1(n1092), .A2(G469), .ZN(n1130) );
XNOR2_X1 U816 ( .A(n1131), .B(n1132), .ZN(n1128) );
NOR2_X1 U817 ( .A1(G110), .A2(KEYINPUT24), .ZN(n1132) );
XOR2_X1 U818 ( .A(n1133), .B(n1134), .Z(n1126) );
XNOR2_X1 U819 ( .A(KEYINPUT3), .B(n1135), .ZN(n1134) );
INV_X1 U820 ( .A(G140), .ZN(n1135) );
XOR2_X1 U821 ( .A(KEYINPUT47), .B(KEYINPUT40), .Z(n1133) );
NOR2_X1 U822 ( .A1(n1088), .A2(n1136), .ZN(G51) );
XOR2_X1 U823 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U824 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U825 ( .A1(n1092), .A2(n1141), .ZN(n1139) );
NOR2_X1 U826 ( .A1(n1142), .A2(n998), .ZN(n1092) );
NOR4_X1 U827 ( .A1(n1143), .A2(n1077), .A3(n1058), .A4(n1076), .ZN(n998) );
NAND4_X1 U828 ( .A1(n1144), .A2(n1105), .A3(n1145), .A4(n985), .ZN(n1076) );
NAND3_X1 U829 ( .A1(n1012), .A2(n1146), .A3(n994), .ZN(n985) );
NAND3_X1 U830 ( .A1(n1012), .A2(n1146), .A3(n995), .ZN(n1105) );
NAND3_X1 U831 ( .A1(n999), .A2(n1146), .A3(n1010), .ZN(n1144) );
NAND4_X1 U832 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1058) );
AND3_X1 U833 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NAND2_X1 U834 ( .A1(n1154), .A2(n1155), .ZN(n1149) );
NAND2_X1 U835 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U836 ( .A1(n1158), .A2(n994), .ZN(n1157) );
XOR2_X1 U837 ( .A(n1159), .B(KEYINPUT43), .Z(n1156) );
NAND3_X1 U838 ( .A1(n1158), .A2(n999), .A3(n1160), .ZN(n1147) );
XNOR2_X1 U839 ( .A(n1008), .B(KEYINPUT59), .ZN(n1160) );
NAND4_X1 U840 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1077) );
XOR2_X1 U841 ( .A(n1057), .B(KEYINPUT38), .Z(n1143) );
XNOR2_X1 U842 ( .A(G125), .B(KEYINPUT18), .ZN(n1137) );
NOR2_X1 U843 ( .A1(n1049), .A2(G952), .ZN(n1088) );
XNOR2_X1 U844 ( .A(G146), .B(n1151), .ZN(G48) );
NAND3_X1 U845 ( .A1(n995), .A2(n1154), .A3(n1158), .ZN(n1151) );
XOR2_X1 U846 ( .A(n1153), .B(n1165), .Z(G45) );
NAND2_X1 U847 ( .A1(KEYINPUT21), .A2(G143), .ZN(n1165) );
NAND3_X1 U848 ( .A1(n1166), .A2(n1011), .A3(n1167), .ZN(n1153) );
NOR3_X1 U849 ( .A1(n1014), .A2(n1168), .A3(n1169), .ZN(n1167) );
XNOR2_X1 U850 ( .A(G140), .B(n1170), .ZN(G42) );
NAND2_X1 U851 ( .A1(KEYINPUT11), .A2(n1057), .ZN(n1170) );
AND2_X1 U852 ( .A1(n1010), .A2(n1171), .ZN(n1057) );
XOR2_X1 U853 ( .A(G137), .B(n1172), .Z(G39) );
NOR3_X1 U854 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
XNOR2_X1 U855 ( .A(G134), .B(n1148), .ZN(G36) );
NAND4_X1 U856 ( .A1(n1166), .A2(n1008), .A3(n1011), .A4(n994), .ZN(n1148) );
XNOR2_X1 U857 ( .A(n1152), .B(n1176), .ZN(G33) );
NOR2_X1 U858 ( .A1(KEYINPUT57), .A2(n1177), .ZN(n1176) );
NAND2_X1 U859 ( .A1(n1171), .A2(n1011), .ZN(n1152) );
AND3_X1 U860 ( .A1(n1008), .A2(n995), .A3(n1166), .ZN(n1171) );
INV_X1 U861 ( .A(n1175), .ZN(n1008) );
NAND2_X1 U862 ( .A1(n1017), .A2(n1178), .ZN(n1175) );
XNOR2_X1 U863 ( .A(KEYINPUT36), .B(n1179), .ZN(n1178) );
XNOR2_X1 U864 ( .A(G128), .B(n1180), .ZN(G30) );
NAND3_X1 U865 ( .A1(n1158), .A2(n994), .A3(n1181), .ZN(n1180) );
XNOR2_X1 U866 ( .A(n1154), .B(KEYINPUT39), .ZN(n1181) );
INV_X1 U867 ( .A(n1173), .ZN(n1158) );
NAND3_X1 U868 ( .A1(n1182), .A2(n1183), .A3(n1166), .ZN(n1173) );
NOR2_X1 U869 ( .A1(n1020), .A2(n1184), .ZN(n1166) );
INV_X1 U870 ( .A(n1185), .ZN(n1184) );
XOR2_X1 U871 ( .A(n1145), .B(n1186), .Z(G3) );
NAND2_X1 U872 ( .A1(KEYINPUT32), .A2(G101), .ZN(n1186) );
NAND3_X1 U873 ( .A1(n1011), .A2(n1146), .A3(n999), .ZN(n1145) );
NOR3_X1 U874 ( .A1(n1014), .A2(n1187), .A3(n1020), .ZN(n1146) );
XOR2_X1 U875 ( .A(n1188), .B(n1189), .Z(G27) );
NOR2_X1 U876 ( .A1(KEYINPUT61), .A2(n1190), .ZN(n1189) );
INV_X1 U877 ( .A(G125), .ZN(n1190) );
NOR2_X1 U878 ( .A1(n1014), .A2(n1159), .ZN(n1188) );
NAND4_X1 U879 ( .A1(n1010), .A2(n995), .A3(n1003), .A4(n1185), .ZN(n1159) );
NAND2_X1 U880 ( .A1(n1024), .A2(n1191), .ZN(n1185) );
NAND4_X1 U881 ( .A1(G953), .A2(G902), .A3(n1192), .A4(n1051), .ZN(n1191) );
INV_X1 U882 ( .A(G900), .ZN(n1051) );
XNOR2_X1 U883 ( .A(G122), .B(n1161), .ZN(G24) );
NAND4_X1 U884 ( .A1(n1193), .A2(n1012), .A3(n1194), .A4(n1195), .ZN(n1161) );
NOR2_X1 U885 ( .A1(n1183), .A2(n1182), .ZN(n1012) );
XNOR2_X1 U886 ( .A(G119), .B(n1162), .ZN(G21) );
NAND4_X1 U887 ( .A1(n999), .A2(n1193), .A3(n1182), .A4(n1183), .ZN(n1162) );
XOR2_X1 U888 ( .A(n1163), .B(n1196), .Z(G18) );
NAND2_X1 U889 ( .A1(KEYINPUT51), .A2(G116), .ZN(n1196) );
NAND3_X1 U890 ( .A1(n1193), .A2(n994), .A3(n1011), .ZN(n1163) );
AND2_X1 U891 ( .A1(n1197), .A2(n1194), .ZN(n994) );
XNOR2_X1 U892 ( .A(G113), .B(n1164), .ZN(G15) );
NAND3_X1 U893 ( .A1(n1011), .A2(n1193), .A3(n995), .ZN(n1164) );
NOR2_X1 U894 ( .A1(n1194), .A2(n1168), .ZN(n995) );
INV_X1 U895 ( .A(n1169), .ZN(n1194) );
NOR3_X1 U896 ( .A1(n1014), .A2(n1187), .A3(n993), .ZN(n1193) );
INV_X1 U897 ( .A(n1003), .ZN(n993) );
NOR2_X1 U898 ( .A1(n1022), .A2(n1043), .ZN(n1003) );
INV_X1 U899 ( .A(n1023), .ZN(n1043) );
INV_X1 U900 ( .A(n1154), .ZN(n1014) );
NOR2_X1 U901 ( .A1(n1183), .A2(n1198), .ZN(n1011) );
INV_X1 U902 ( .A(n1182), .ZN(n1198) );
XOR2_X1 U903 ( .A(G110), .B(n1199), .Z(G12) );
NOR2_X1 U904 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NOR2_X1 U905 ( .A1(KEYINPUT58), .A2(n1202), .ZN(n1201) );
INV_X1 U906 ( .A(n1203), .ZN(n1202) );
NOR2_X1 U907 ( .A1(KEYINPUT45), .A2(n1203), .ZN(n1200) );
NAND3_X1 U908 ( .A1(n1010), .A2(n999), .A3(n1204), .ZN(n1203) );
NOR3_X1 U909 ( .A1(n1020), .A2(n1187), .A3(n1205), .ZN(n1204) );
XNOR2_X1 U910 ( .A(n1154), .B(KEYINPUT31), .ZN(n1205) );
NOR2_X1 U911 ( .A1(n1017), .A2(n1016), .ZN(n1154) );
INV_X1 U912 ( .A(n1179), .ZN(n1016) );
NAND2_X1 U913 ( .A1(G214), .A2(n1206), .ZN(n1179) );
INV_X1 U914 ( .A(n1032), .ZN(n1017) );
XNOR2_X1 U915 ( .A(n1207), .B(n1141), .ZN(n1032) );
AND2_X1 U916 ( .A1(G210), .A2(n1206), .ZN(n1141) );
NAND2_X1 U917 ( .A1(n1208), .A2(n1142), .ZN(n1206) );
INV_X1 U918 ( .A(G237), .ZN(n1208) );
NAND2_X1 U919 ( .A1(n1209), .A2(n1142), .ZN(n1207) );
XOR2_X1 U920 ( .A(n1140), .B(n1210), .Z(n1209) );
XOR2_X1 U921 ( .A(KEYINPUT48), .B(n1211), .Z(n1210) );
NOR2_X1 U922 ( .A1(G125), .A2(n1212), .ZN(n1211) );
XNOR2_X1 U923 ( .A(KEYINPUT42), .B(KEYINPUT34), .ZN(n1212) );
XOR2_X1 U924 ( .A(n1213), .B(n1214), .Z(n1140) );
XOR2_X1 U925 ( .A(n1086), .B(n1215), .Z(n1214) );
XNOR2_X1 U926 ( .A(G110), .B(n1216), .ZN(n1086) );
XNOR2_X1 U927 ( .A(n1087), .B(n1217), .ZN(n1213) );
AND2_X1 U928 ( .A1(n1049), .A2(G224), .ZN(n1217) );
XOR2_X1 U929 ( .A(n1118), .B(n1218), .Z(n1087) );
AND2_X1 U930 ( .A1(n1024), .A2(n1219), .ZN(n1187) );
NAND3_X1 U931 ( .A1(G902), .A2(n1192), .A3(n1083), .ZN(n1219) );
NOR2_X1 U932 ( .A1(n1049), .A2(G898), .ZN(n1083) );
NAND3_X1 U933 ( .A1(n1192), .A2(n1049), .A3(G952), .ZN(n1024) );
NAND2_X1 U934 ( .A1(G237), .A2(G234), .ZN(n1192) );
NAND2_X1 U935 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NAND2_X1 U936 ( .A1(G221), .A2(n1220), .ZN(n1023) );
NAND2_X1 U937 ( .A1(n1045), .A2(n1033), .ZN(n1022) );
NAND2_X1 U938 ( .A1(G469), .A2(n1221), .ZN(n1033) );
OR2_X1 U939 ( .A1(n1221), .A2(G469), .ZN(n1045) );
NAND3_X1 U940 ( .A1(n1222), .A2(n1223), .A3(n1142), .ZN(n1221) );
OR3_X1 U941 ( .A1(n1224), .A2(n1225), .A3(KEYINPUT9), .ZN(n1223) );
NAND2_X1 U942 ( .A1(n1226), .A2(KEYINPUT9), .ZN(n1222) );
XOR2_X1 U943 ( .A(n1225), .B(n1224), .Z(n1226) );
XNOR2_X1 U944 ( .A(n1227), .B(n1228), .ZN(n1224) );
NOR2_X1 U945 ( .A1(KEYINPUT41), .A2(n1131), .ZN(n1228) );
NOR2_X1 U946 ( .A1(n1050), .A2(G953), .ZN(n1131) );
INV_X1 U947 ( .A(G227), .ZN(n1050) );
XNOR2_X1 U948 ( .A(G110), .B(G140), .ZN(n1227) );
XNOR2_X1 U949 ( .A(n1229), .B(n1124), .ZN(n1225) );
XNOR2_X1 U950 ( .A(n1230), .B(n1218), .ZN(n1124) );
XNOR2_X1 U951 ( .A(n1109), .B(n1231), .ZN(n1218) );
XOR2_X1 U952 ( .A(G107), .B(G104), .Z(n1231) );
NAND2_X1 U953 ( .A1(KEYINPUT35), .A2(n1067), .ZN(n1229) );
XNOR2_X1 U954 ( .A(n1232), .B(n1233), .ZN(n1067) );
NOR2_X1 U955 ( .A1(G128), .A2(KEYINPUT10), .ZN(n1233) );
INV_X1 U956 ( .A(n1174), .ZN(n999) );
NAND2_X1 U957 ( .A1(n1197), .A2(n1169), .ZN(n1174) );
XNOR2_X1 U958 ( .A(n1044), .B(n1234), .ZN(n1169) );
NOR2_X1 U959 ( .A1(G478), .A2(KEYINPUT60), .ZN(n1234) );
OR2_X1 U960 ( .A1(n1096), .A2(G902), .ZN(n1044) );
XNOR2_X1 U961 ( .A(n1235), .B(n1236), .ZN(n1096) );
XOR2_X1 U962 ( .A(G107), .B(n1237), .Z(n1236) );
NOR2_X1 U963 ( .A1(KEYINPUT63), .A2(n1238), .ZN(n1237) );
XOR2_X1 U964 ( .A(n1239), .B(n1240), .Z(n1238) );
NOR2_X1 U965 ( .A1(KEYINPUT52), .A2(G134), .ZN(n1240) );
XNOR2_X1 U966 ( .A(G128), .B(G143), .ZN(n1239) );
XOR2_X1 U967 ( .A(n1241), .B(n1242), .Z(n1235) );
NOR2_X1 U968 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
INV_X1 U969 ( .A(G217), .ZN(n1244) );
NAND2_X1 U970 ( .A1(KEYINPUT53), .A2(n1245), .ZN(n1241) );
XNOR2_X1 U971 ( .A(n1216), .B(G116), .ZN(n1245) );
INV_X1 U972 ( .A(G122), .ZN(n1216) );
XNOR2_X1 U973 ( .A(n1195), .B(KEYINPUT33), .ZN(n1197) );
INV_X1 U974 ( .A(n1168), .ZN(n1195) );
XOR2_X1 U975 ( .A(n1038), .B(n1040), .Z(n1168) );
INV_X1 U976 ( .A(G475), .ZN(n1040) );
NOR2_X1 U977 ( .A1(n1101), .A2(G902), .ZN(n1038) );
NAND2_X1 U978 ( .A1(n1246), .A2(n1247), .ZN(n1101) );
NAND2_X1 U979 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
INV_X1 U980 ( .A(n1250), .ZN(n1249) );
XOR2_X1 U981 ( .A(KEYINPUT28), .B(n1251), .Z(n1248) );
NAND2_X1 U982 ( .A1(n1250), .A2(n1252), .ZN(n1246) );
XNOR2_X1 U983 ( .A(n1251), .B(KEYINPUT27), .ZN(n1252) );
XNOR2_X1 U984 ( .A(n1253), .B(n1254), .ZN(n1251) );
XOR2_X1 U985 ( .A(G104), .B(n1255), .Z(n1254) );
XOR2_X1 U986 ( .A(KEYINPUT46), .B(G146), .Z(n1255) );
XOR2_X1 U987 ( .A(n1256), .B(n1065), .Z(n1253) );
NAND2_X1 U988 ( .A1(n1257), .A2(KEYINPUT13), .ZN(n1256) );
XNOR2_X1 U989 ( .A(G122), .B(n1258), .ZN(n1257) );
NOR2_X1 U990 ( .A1(G113), .A2(KEYINPUT14), .ZN(n1258) );
XNOR2_X1 U991 ( .A(n1259), .B(n1260), .ZN(n1250) );
XNOR2_X1 U992 ( .A(G143), .B(n1177), .ZN(n1260) );
INV_X1 U993 ( .A(G131), .ZN(n1177) );
NAND2_X1 U994 ( .A1(G214), .A2(n1261), .ZN(n1259) );
AND2_X1 U995 ( .A1(n1262), .A2(n1183), .ZN(n1010) );
XNOR2_X1 U996 ( .A(n1263), .B(n1093), .ZN(n1183) );
AND2_X1 U997 ( .A1(G217), .A2(n1220), .ZN(n1093) );
NAND2_X1 U998 ( .A1(G234), .A2(n1142), .ZN(n1220) );
NAND2_X1 U999 ( .A1(n1091), .A2(n1142), .ZN(n1263) );
INV_X1 U1000 ( .A(G902), .ZN(n1142) );
XOR2_X1 U1001 ( .A(n1264), .B(n1265), .Z(n1091) );
XOR2_X1 U1002 ( .A(n1266), .B(n1267), .Z(n1265) );
XNOR2_X1 U1003 ( .A(n1268), .B(n1269), .ZN(n1267) );
NOR2_X1 U1004 ( .A1(G110), .A2(KEYINPUT15), .ZN(n1269) );
NAND2_X1 U1005 ( .A1(KEYINPUT50), .A2(n1270), .ZN(n1268) );
XOR2_X1 U1006 ( .A(n1271), .B(n1272), .Z(n1264) );
NOR2_X1 U1007 ( .A1(n1243), .A2(n1273), .ZN(n1272) );
INV_X1 U1008 ( .A(G221), .ZN(n1273) );
NAND2_X1 U1009 ( .A1(G234), .A2(n1049), .ZN(n1243) );
INV_X1 U1010 ( .A(G953), .ZN(n1049) );
XOR2_X1 U1011 ( .A(n1274), .B(G128), .Z(n1271) );
NAND2_X1 U1012 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND2_X1 U1013 ( .A1(G146), .A2(n1065), .ZN(n1276) );
XOR2_X1 U1014 ( .A(KEYINPUT55), .B(n1277), .Z(n1275) );
NOR2_X1 U1015 ( .A1(G146), .A2(n1065), .ZN(n1277) );
XOR2_X1 U1016 ( .A(G125), .B(G140), .Z(n1065) );
XNOR2_X1 U1017 ( .A(n1182), .B(KEYINPUT20), .ZN(n1262) );
XNOR2_X1 U1018 ( .A(n1278), .B(G472), .ZN(n1182) );
NAND2_X1 U1019 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XOR2_X1 U1020 ( .A(n1120), .B(n1281), .Z(n1280) );
XNOR2_X1 U1021 ( .A(n1282), .B(n1109), .ZN(n1281) );
INV_X1 U1022 ( .A(G101), .ZN(n1109) );
NAND2_X1 U1023 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U1024 ( .A1(n1122), .A2(n1118), .ZN(n1284) );
XOR2_X1 U1025 ( .A(KEYINPUT56), .B(n1285), .Z(n1283) );
NOR2_X1 U1026 ( .A1(n1122), .A2(n1118), .ZN(n1285) );
XOR2_X1 U1027 ( .A(G113), .B(n1286), .Z(n1118) );
XNOR2_X1 U1028 ( .A(n1270), .B(G116), .ZN(n1286) );
INV_X1 U1029 ( .A(G119), .ZN(n1270) );
XNOR2_X1 U1030 ( .A(n1230), .B(n1215), .ZN(n1122) );
XOR2_X1 U1031 ( .A(G128), .B(n1232), .Z(n1215) );
XOR2_X1 U1032 ( .A(G143), .B(G146), .Z(n1232) );
XNOR2_X1 U1033 ( .A(n1069), .B(n1287), .ZN(n1230) );
NOR2_X1 U1034 ( .A1(G134), .A2(KEYINPUT0), .ZN(n1287) );
XOR2_X1 U1035 ( .A(G131), .B(n1266), .Z(n1069) );
XOR2_X1 U1036 ( .A(G137), .B(KEYINPUT62), .Z(n1266) );
NAND2_X1 U1037 ( .A1(G210), .A2(n1261), .ZN(n1120) );
NOR2_X1 U1038 ( .A1(G953), .A2(G237), .ZN(n1261) );
XNOR2_X1 U1039 ( .A(G902), .B(KEYINPUT5), .ZN(n1279) );
endmodule


