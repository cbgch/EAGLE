//Key = 0011000101000100010110011101101001100100001001010011010010111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;

XOR2_X1 U780 ( .A(n1087), .B(n1088), .Z(G9) );
NOR2_X1 U781 ( .A1(KEYINPUT41), .A2(n1089), .ZN(n1088) );
INV_X1 U782 ( .A(G107), .ZN(n1089) );
NOR2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(G75) );
NOR4_X1 U784 ( .A1(n1092), .A2(n1093), .A3(G953), .A4(n1094), .ZN(n1091) );
NOR2_X1 U785 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NOR2_X1 U786 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U789 ( .A1(KEYINPUT23), .A2(n1103), .ZN(n1102) );
NOR4_X1 U790 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1103) );
NOR3_X1 U791 ( .A1(n1108), .A2(n1104), .A3(n1109), .ZN(n1101) );
NOR3_X1 U792 ( .A1(n1110), .A2(n1111), .A3(n1112), .ZN(n1109) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1107), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U795 ( .A1(n1106), .A2(n1116), .ZN(n1110) );
NOR3_X1 U796 ( .A1(n1107), .A2(n1104), .A3(n1117), .ZN(n1097) );
NOR2_X1 U797 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR3_X1 U798 ( .A1(n1108), .A2(n1120), .A3(n1121), .ZN(n1119) );
XNOR2_X1 U799 ( .A(n1122), .B(KEYINPUT52), .ZN(n1120) );
NOR3_X1 U800 ( .A1(n1106), .A2(n1123), .A3(n1100), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U802 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
AND2_X1 U803 ( .A1(n1128), .A2(KEYINPUT23), .ZN(n1124) );
NAND2_X1 U804 ( .A1(n1129), .A2(n1130), .ZN(n1092) );
NAND3_X1 U805 ( .A1(n1131), .A2(n1132), .A3(n1133), .ZN(n1130) );
NOR3_X1 U806 ( .A1(n1108), .A2(n1106), .A3(n1107), .ZN(n1133) );
XNOR2_X1 U807 ( .A(n1104), .B(KEYINPUT10), .ZN(n1132) );
INV_X1 U808 ( .A(n1134), .ZN(n1104) );
XNOR2_X1 U809 ( .A(n1135), .B(KEYINPUT20), .ZN(n1131) );
NOR3_X1 U810 ( .A1(n1094), .A2(G953), .A3(G952), .ZN(n1090) );
AND4_X1 U811 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1094) );
NOR4_X1 U812 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
AND2_X1 U813 ( .A1(n1144), .A2(G469), .ZN(n1143) );
INV_X1 U814 ( .A(n1121), .ZN(n1141) );
NOR2_X1 U815 ( .A1(n1145), .A2(n1146), .ZN(n1138) );
XNOR2_X1 U816 ( .A(G472), .B(n1147), .ZN(n1146) );
XOR2_X1 U817 ( .A(n1148), .B(n1149), .Z(n1145) );
NOR2_X1 U818 ( .A1(KEYINPUT40), .A2(n1150), .ZN(n1149) );
XNOR2_X1 U819 ( .A(n1151), .B(n1152), .ZN(n1136) );
XOR2_X1 U820 ( .A(n1153), .B(n1154), .Z(G72) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR3_X1 U822 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1156) );
NOR2_X1 U823 ( .A1(G953), .A2(n1160), .ZN(n1155) );
XNOR2_X1 U824 ( .A(n1161), .B(n1159), .ZN(n1160) );
NAND2_X1 U825 ( .A1(n1162), .A2(KEYINPUT30), .ZN(n1159) );
XOR2_X1 U826 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U827 ( .A(n1165), .B(n1166), .ZN(n1164) );
NOR2_X1 U828 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
AND3_X1 U829 ( .A1(KEYINPUT5), .A2(n1169), .A3(G125), .ZN(n1168) );
NOR2_X1 U830 ( .A1(KEYINPUT5), .A2(n1170), .ZN(n1167) );
XOR2_X1 U831 ( .A(n1171), .B(n1172), .Z(n1163) );
XNOR2_X1 U832 ( .A(KEYINPUT25), .B(n1173), .ZN(n1171) );
NOR2_X1 U833 ( .A1(G131), .A2(KEYINPUT46), .ZN(n1173) );
NAND3_X1 U834 ( .A1(G953), .A2(n1174), .A3(KEYINPUT47), .ZN(n1153) );
NAND2_X1 U835 ( .A1(G900), .A2(G227), .ZN(n1174) );
NAND2_X1 U836 ( .A1(n1175), .A2(n1176), .ZN(G69) );
NAND2_X1 U837 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND3_X1 U838 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1177) );
XNOR2_X1 U839 ( .A(n1182), .B(n1183), .ZN(n1181) );
NAND2_X1 U840 ( .A1(n1157), .A2(n1184), .ZN(n1182) );
OR2_X1 U841 ( .A1(n1157), .A2(G224), .ZN(n1179) );
NAND2_X1 U842 ( .A1(n1185), .A2(n1186), .ZN(n1175) );
NAND2_X1 U843 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U844 ( .A1(n1189), .A2(n1183), .ZN(n1188) );
INV_X1 U845 ( .A(KEYINPUT44), .ZN(n1183) );
NAND2_X1 U846 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NAND2_X1 U847 ( .A1(n1192), .A2(n1157), .ZN(n1191) );
NAND2_X1 U848 ( .A1(G224), .A2(G953), .ZN(n1190) );
NAND3_X1 U849 ( .A1(n1184), .A2(n1157), .A3(KEYINPUT44), .ZN(n1187) );
INV_X1 U850 ( .A(n1178), .ZN(n1185) );
NAND2_X1 U851 ( .A1(n1193), .A2(n1180), .ZN(n1178) );
INV_X1 U852 ( .A(n1194), .ZN(n1180) );
XOR2_X1 U853 ( .A(n1195), .B(n1196), .Z(n1193) );
XOR2_X1 U854 ( .A(n1197), .B(n1198), .Z(n1196) );
NAND2_X1 U855 ( .A1(KEYINPUT59), .A2(n1199), .ZN(n1197) );
NOR2_X1 U856 ( .A1(n1200), .A2(n1201), .ZN(G66) );
NOR3_X1 U857 ( .A1(n1148), .A2(n1202), .A3(n1203), .ZN(n1201) );
NOR2_X1 U858 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NOR2_X1 U859 ( .A1(n1129), .A2(n1150), .ZN(n1204) );
NOR3_X1 U860 ( .A1(n1206), .A2(n1150), .A3(n1207), .ZN(n1202) );
INV_X1 U861 ( .A(n1205), .ZN(n1206) );
NOR2_X1 U862 ( .A1(n1200), .A2(n1208), .ZN(G63) );
XOR2_X1 U863 ( .A(n1209), .B(n1210), .Z(n1208) );
NAND2_X1 U864 ( .A1(n1211), .A2(G478), .ZN(n1209) );
NOR2_X1 U865 ( .A1(n1200), .A2(n1212), .ZN(G60) );
XOR2_X1 U866 ( .A(n1213), .B(n1214), .Z(n1212) );
NAND2_X1 U867 ( .A1(n1211), .A2(G475), .ZN(n1213) );
XNOR2_X1 U868 ( .A(G104), .B(n1215), .ZN(G6) );
NAND4_X1 U869 ( .A1(n1216), .A2(n1217), .A3(n1122), .A4(n1218), .ZN(n1215) );
XNOR2_X1 U870 ( .A(n1219), .B(KEYINPUT27), .ZN(n1216) );
NOR2_X1 U871 ( .A1(n1200), .A2(n1220), .ZN(G57) );
XOR2_X1 U872 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U873 ( .A(n1223), .B(n1224), .Z(n1222) );
XNOR2_X1 U874 ( .A(n1225), .B(n1226), .ZN(n1224) );
NAND3_X1 U875 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1223) );
NAND2_X1 U876 ( .A1(KEYINPUT21), .A2(n1230), .ZN(n1229) );
NAND2_X1 U877 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U878 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND4_X1 U879 ( .A1(n1231), .A2(n1235), .A3(KEYINPUT51), .A4(n1233), .ZN(n1228) );
NAND2_X1 U880 ( .A1(n1236), .A2(n1237), .ZN(n1227) );
NAND3_X1 U881 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1237) );
NAND2_X1 U882 ( .A1(KEYINPUT51), .A2(KEYINPUT21), .ZN(n1240) );
NAND2_X1 U883 ( .A1(KEYINPUT37), .A2(n1241), .ZN(n1239) );
NAND2_X1 U884 ( .A1(n1231), .A2(n1242), .ZN(n1241) );
NAND2_X1 U885 ( .A1(n1235), .A2(n1234), .ZN(n1242) );
INV_X1 U886 ( .A(KEYINPUT51), .ZN(n1234) );
INV_X1 U887 ( .A(KEYINPUT21), .ZN(n1235) );
OR2_X1 U888 ( .A1(n1243), .A2(KEYINPUT37), .ZN(n1238) );
INV_X1 U889 ( .A(n1233), .ZN(n1236) );
XNOR2_X1 U890 ( .A(n1244), .B(KEYINPUT12), .ZN(n1233) );
XNOR2_X1 U891 ( .A(n1245), .B(n1246), .ZN(n1221) );
NOR3_X1 U892 ( .A1(n1207), .A2(KEYINPUT38), .A3(n1247), .ZN(n1246) );
INV_X1 U893 ( .A(G472), .ZN(n1247) );
INV_X1 U894 ( .A(n1211), .ZN(n1207) );
NOR2_X1 U895 ( .A1(n1200), .A2(n1248), .ZN(G54) );
XOR2_X1 U896 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U897 ( .A(n1251), .B(n1252), .Z(n1250) );
NOR3_X1 U898 ( .A1(n1253), .A2(n1254), .A3(n1255), .ZN(n1251) );
XNOR2_X1 U899 ( .A(KEYINPUT16), .B(n1256), .ZN(n1253) );
XOR2_X1 U900 ( .A(n1257), .B(KEYINPUT48), .Z(n1249) );
NAND2_X1 U901 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
NOR2_X1 U902 ( .A1(n1200), .A2(n1260), .ZN(G51) );
XOR2_X1 U903 ( .A(n1261), .B(n1262), .Z(n1260) );
XNOR2_X1 U904 ( .A(n1231), .B(n1263), .ZN(n1262) );
XOR2_X1 U905 ( .A(n1264), .B(n1265), .Z(n1261) );
XNOR2_X1 U906 ( .A(n1266), .B(n1267), .ZN(n1265) );
NAND2_X1 U907 ( .A1(n1211), .A2(n1152), .ZN(n1266) );
NOR2_X1 U908 ( .A1(n1254), .A2(n1129), .ZN(n1211) );
INV_X1 U909 ( .A(n1256), .ZN(n1129) );
NAND2_X1 U910 ( .A1(n1161), .A2(n1192), .ZN(n1256) );
INV_X1 U911 ( .A(n1184), .ZN(n1192) );
NAND4_X1 U912 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1184) );
NOR2_X1 U913 ( .A1(n1272), .A2(n1087), .ZN(n1270) );
NOR4_X1 U914 ( .A1(n1116), .A2(n1273), .A3(n1106), .A4(n1274), .ZN(n1087) );
INV_X1 U915 ( .A(n1275), .ZN(n1116) );
NAND2_X1 U916 ( .A1(n1276), .A2(n1277), .ZN(n1268) );
NAND3_X1 U917 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
NAND3_X1 U918 ( .A1(n1281), .A2(n1137), .A3(n1282), .ZN(n1280) );
NAND2_X1 U919 ( .A1(n1218), .A2(n1283), .ZN(n1279) );
NAND2_X1 U920 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
NAND2_X1 U921 ( .A1(n1111), .A2(n1286), .ZN(n1285) );
INV_X1 U922 ( .A(KEYINPUT43), .ZN(n1286) );
NAND2_X1 U923 ( .A1(n1137), .A2(n1287), .ZN(n1284) );
NAND2_X1 U924 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XNOR2_X1 U925 ( .A(n1115), .B(KEYINPUT35), .ZN(n1288) );
NAND3_X1 U926 ( .A1(KEYINPUT43), .A2(n1111), .A3(n1274), .ZN(n1278) );
AND2_X1 U927 ( .A1(n1290), .A2(n1122), .ZN(n1111) );
AND4_X1 U928 ( .A1(n1291), .A2(n1292), .A3(n1293), .A4(n1294), .ZN(n1161) );
NOR4_X1 U929 ( .A1(n1295), .A2(n1296), .A3(n1297), .A4(n1298), .ZN(n1294) );
AND2_X1 U930 ( .A1(n1299), .A2(n1300), .ZN(n1293) );
NAND3_X1 U931 ( .A1(n1114), .A2(n1275), .A3(n1301), .ZN(n1291) );
NAND2_X1 U932 ( .A1(KEYINPUT45), .A2(n1302), .ZN(n1264) );
NOR2_X1 U933 ( .A1(n1157), .A2(G952), .ZN(n1200) );
NAND2_X1 U934 ( .A1(n1303), .A2(n1304), .ZN(G48) );
NAND2_X1 U935 ( .A1(G146), .A2(n1292), .ZN(n1304) );
XOR2_X1 U936 ( .A(KEYINPUT2), .B(n1305), .Z(n1303) );
NOR2_X1 U937 ( .A1(G146), .A2(n1292), .ZN(n1305) );
NAND4_X1 U938 ( .A1(n1217), .A2(n1281), .A3(n1306), .A4(n1128), .ZN(n1292) );
XOR2_X1 U939 ( .A(G143), .B(n1298), .Z(G45) );
AND4_X1 U940 ( .A1(n1307), .A2(n1308), .A3(n1135), .A4(n1309), .ZN(n1298) );
NOR3_X1 U941 ( .A1(n1289), .A2(n1105), .A3(n1310), .ZN(n1309) );
XOR2_X1 U942 ( .A(n1311), .B(n1297), .Z(G42) );
AND3_X1 U943 ( .A1(n1301), .A2(n1290), .A3(n1115), .ZN(n1297) );
NAND2_X1 U944 ( .A1(KEYINPUT9), .A2(n1169), .ZN(n1311) );
XOR2_X1 U945 ( .A(G137), .B(n1296), .Z(G39) );
AND3_X1 U946 ( .A1(n1301), .A2(n1137), .A3(n1281), .ZN(n1296) );
NAND2_X1 U947 ( .A1(n1312), .A2(n1313), .ZN(G36) );
NAND2_X1 U948 ( .A1(G134), .A2(n1314), .ZN(n1313) );
XOR2_X1 U949 ( .A(n1315), .B(KEYINPUT4), .Z(n1312) );
OR2_X1 U950 ( .A1(n1314), .A2(G134), .ZN(n1315) );
NAND3_X1 U951 ( .A1(n1301), .A2(n1275), .A3(n1316), .ZN(n1314) );
XNOR2_X1 U952 ( .A(n1114), .B(KEYINPUT42), .ZN(n1316) );
XOR2_X1 U953 ( .A(n1295), .B(n1317), .Z(G33) );
NOR2_X1 U954 ( .A1(KEYINPUT18), .A2(n1318), .ZN(n1317) );
AND3_X1 U955 ( .A1(n1114), .A2(n1290), .A3(n1301), .ZN(n1295) );
NOR4_X1 U956 ( .A1(n1310), .A2(n1105), .A3(n1100), .A4(n1095), .ZN(n1301) );
INV_X1 U957 ( .A(n1319), .ZN(n1095) );
INV_X1 U958 ( .A(n1128), .ZN(n1105) );
NAND2_X1 U959 ( .A1(n1320), .A2(n1321), .ZN(G30) );
NAND2_X1 U960 ( .A1(G128), .A2(n1300), .ZN(n1321) );
XOR2_X1 U961 ( .A(n1322), .B(KEYINPUT26), .Z(n1320) );
OR2_X1 U962 ( .A1(n1300), .A2(G128), .ZN(n1322) );
NAND4_X1 U963 ( .A1(n1135), .A2(n1218), .A3(n1275), .A4(n1323), .ZN(n1300) );
NOR2_X1 U964 ( .A1(n1310), .A2(n1324), .ZN(n1323) );
XOR2_X1 U965 ( .A(n1325), .B(n1326), .Z(G3) );
NOR3_X1 U966 ( .A1(n1327), .A2(n1274), .A3(n1107), .ZN(n1326) );
INV_X1 U967 ( .A(n1137), .ZN(n1107) );
INV_X1 U968 ( .A(n1218), .ZN(n1274) );
NAND3_X1 U969 ( .A1(n1328), .A2(n1329), .A3(n1114), .ZN(n1327) );
INV_X1 U970 ( .A(n1289), .ZN(n1114) );
OR2_X1 U971 ( .A1(n1276), .A2(KEYINPUT57), .ZN(n1329) );
NAND2_X1 U972 ( .A1(KEYINPUT57), .A2(n1330), .ZN(n1328) );
NAND2_X1 U973 ( .A1(n1219), .A2(n1331), .ZN(n1330) );
NAND2_X1 U974 ( .A1(KEYINPUT62), .A2(n1226), .ZN(n1325) );
XNOR2_X1 U975 ( .A(G125), .B(n1299), .ZN(G27) );
NAND4_X1 U976 ( .A1(n1282), .A2(n1217), .A3(n1115), .A4(n1306), .ZN(n1299) );
INV_X1 U977 ( .A(n1310), .ZN(n1306) );
NAND2_X1 U978 ( .A1(n1134), .A2(n1332), .ZN(n1310) );
NAND2_X1 U979 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NAND3_X1 U980 ( .A1(G953), .A2(n1158), .A3(G902), .ZN(n1333) );
INV_X1 U981 ( .A(G900), .ZN(n1158) );
AND2_X1 U982 ( .A1(n1290), .A2(n1135), .ZN(n1217) );
XOR2_X1 U983 ( .A(G122), .B(n1272), .Z(G24) );
AND4_X1 U984 ( .A1(n1307), .A2(n1308), .A3(n1122), .A4(n1335), .ZN(n1272) );
NOR2_X1 U985 ( .A1(n1273), .A2(n1108), .ZN(n1335) );
INV_X1 U986 ( .A(n1106), .ZN(n1122) );
NAND2_X1 U987 ( .A1(n1336), .A2(n1337), .ZN(n1106) );
XNOR2_X1 U988 ( .A(n1338), .B(KEYINPUT11), .ZN(n1336) );
XNOR2_X1 U989 ( .A(G119), .B(n1339), .ZN(G21) );
NAND4_X1 U990 ( .A1(n1219), .A2(n1340), .A3(n1137), .A4(n1341), .ZN(n1339) );
NOR2_X1 U991 ( .A1(n1324), .A2(n1108), .ZN(n1341) );
INV_X1 U992 ( .A(n1281), .ZN(n1324) );
NOR2_X1 U993 ( .A1(n1342), .A2(n1337), .ZN(n1281) );
INV_X1 U994 ( .A(n1338), .ZN(n1342) );
XNOR2_X1 U995 ( .A(KEYINPUT36), .B(n1331), .ZN(n1340) );
INV_X1 U996 ( .A(n1343), .ZN(n1219) );
XNOR2_X1 U997 ( .A(G116), .B(n1269), .ZN(G18) );
NAND2_X1 U998 ( .A1(n1344), .A2(n1275), .ZN(n1269) );
NOR2_X1 U999 ( .A1(n1307), .A2(n1345), .ZN(n1275) );
XNOR2_X1 U1000 ( .A(G113), .B(n1271), .ZN(G15) );
NAND2_X1 U1001 ( .A1(n1344), .A2(n1290), .ZN(n1271) );
AND2_X1 U1002 ( .A1(n1345), .A2(n1307), .ZN(n1290) );
INV_X1 U1003 ( .A(n1308), .ZN(n1345) );
NOR3_X1 U1004 ( .A1(n1289), .A2(n1273), .A3(n1108), .ZN(n1344) );
INV_X1 U1005 ( .A(n1282), .ZN(n1108) );
NOR2_X1 U1006 ( .A1(n1126), .A2(n1142), .ZN(n1282) );
INV_X1 U1007 ( .A(n1346), .ZN(n1126) );
INV_X1 U1008 ( .A(n1276), .ZN(n1273) );
NAND2_X1 U1009 ( .A1(n1337), .A2(n1338), .ZN(n1289) );
XNOR2_X1 U1010 ( .A(G110), .B(n1347), .ZN(G12) );
NAND4_X1 U1011 ( .A1(n1115), .A2(n1137), .A3(n1276), .A4(n1218), .ZN(n1347) );
XOR2_X1 U1012 ( .A(n1128), .B(KEYINPUT32), .Z(n1218) );
NOR2_X1 U1013 ( .A1(n1142), .A2(n1346), .ZN(n1128) );
NOR2_X1 U1014 ( .A1(n1348), .A2(n1140), .ZN(n1346) );
NOR2_X1 U1015 ( .A1(n1144), .A2(G469), .ZN(n1140) );
AND2_X1 U1016 ( .A1(n1349), .A2(n1144), .ZN(n1348) );
NAND2_X1 U1017 ( .A1(n1350), .A2(n1351), .ZN(n1144) );
XNOR2_X1 U1018 ( .A(KEYINPUT53), .B(n1254), .ZN(n1351) );
XOR2_X1 U1019 ( .A(n1352), .B(n1252), .Z(n1350) );
XNOR2_X1 U1020 ( .A(n1353), .B(n1354), .ZN(n1252) );
XNOR2_X1 U1021 ( .A(n1355), .B(n1172), .ZN(n1354) );
XOR2_X1 U1022 ( .A(G128), .B(n1356), .Z(n1172) );
NOR2_X1 U1023 ( .A1(KEYINPUT54), .A2(n1357), .ZN(n1356) );
NAND2_X1 U1024 ( .A1(KEYINPUT63), .A2(n1358), .ZN(n1355) );
XNOR2_X1 U1025 ( .A(n1359), .B(n1360), .ZN(n1358) );
NOR2_X1 U1026 ( .A1(n1361), .A2(n1362), .ZN(n1352) );
XOR2_X1 U1027 ( .A(n1259), .B(KEYINPUT17), .Z(n1362) );
NAND3_X1 U1028 ( .A1(G227), .A2(n1157), .A3(n1363), .ZN(n1259) );
INV_X1 U1029 ( .A(n1364), .ZN(n1363) );
INV_X1 U1030 ( .A(n1258), .ZN(n1361) );
NAND2_X1 U1031 ( .A1(n1364), .A2(n1365), .ZN(n1258) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1157), .ZN(n1365) );
XNOR2_X1 U1033 ( .A(G110), .B(n1169), .ZN(n1364) );
XNOR2_X1 U1034 ( .A(KEYINPUT55), .B(n1255), .ZN(n1349) );
INV_X1 U1035 ( .A(G469), .ZN(n1255) );
INV_X1 U1036 ( .A(n1127), .ZN(n1142) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1366), .ZN(n1127) );
NOR2_X1 U1038 ( .A1(n1343), .A2(n1331), .ZN(n1276) );
INV_X1 U1039 ( .A(n1135), .ZN(n1331) );
NOR2_X1 U1040 ( .A1(n1319), .A2(n1100), .ZN(n1135) );
XOR2_X1 U1041 ( .A(n1121), .B(KEYINPUT60), .Z(n1100) );
NAND2_X1 U1042 ( .A1(G214), .A2(n1367), .ZN(n1121) );
NAND2_X1 U1043 ( .A1(n1368), .A2(n1369), .ZN(n1319) );
NAND2_X1 U1044 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1045 ( .A1(n1372), .A2(n1373), .ZN(n1370) );
NAND2_X1 U1046 ( .A1(KEYINPUT13), .A2(n1374), .ZN(n1373) );
NAND2_X1 U1047 ( .A1(n1151), .A2(n1375), .ZN(n1368) );
NAND2_X1 U1048 ( .A1(KEYINPUT13), .A2(n1376), .ZN(n1375) );
NAND2_X1 U1049 ( .A1(n1152), .A2(n1372), .ZN(n1376) );
INV_X1 U1050 ( .A(KEYINPUT1), .ZN(n1372) );
INV_X1 U1051 ( .A(n1371), .ZN(n1152) );
NAND2_X1 U1052 ( .A1(G210), .A2(n1367), .ZN(n1371) );
NAND2_X1 U1053 ( .A1(n1377), .A2(n1254), .ZN(n1367) );
XOR2_X1 U1054 ( .A(KEYINPUT24), .B(G237), .Z(n1377) );
INV_X1 U1055 ( .A(n1374), .ZN(n1151) );
NAND2_X1 U1056 ( .A1(n1378), .A2(n1254), .ZN(n1374) );
XOR2_X1 U1057 ( .A(n1263), .B(n1379), .Z(n1378) );
NOR2_X1 U1058 ( .A1(n1380), .A2(n1381), .ZN(n1379) );
XOR2_X1 U1059 ( .A(n1382), .B(KEYINPUT28), .Z(n1381) );
NAND2_X1 U1060 ( .A1(n1383), .A2(n1267), .ZN(n1382) );
NOR2_X1 U1061 ( .A1(n1267), .A2(n1383), .ZN(n1380) );
XNOR2_X1 U1062 ( .A(G125), .B(n1243), .ZN(n1383) );
INV_X1 U1063 ( .A(n1231), .ZN(n1243) );
NAND2_X1 U1064 ( .A1(G224), .A2(n1157), .ZN(n1267) );
XOR2_X1 U1065 ( .A(n1198), .B(n1384), .Z(n1263) );
NOR2_X1 U1066 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
XOR2_X1 U1067 ( .A(n1387), .B(KEYINPUT33), .Z(n1386) );
NAND2_X1 U1068 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
XNOR2_X1 U1069 ( .A(KEYINPUT7), .B(n1390), .ZN(n1389) );
XOR2_X1 U1070 ( .A(n1195), .B(KEYINPUT22), .Z(n1388) );
NOR2_X1 U1071 ( .A1(n1390), .A2(n1195), .ZN(n1385) );
XOR2_X1 U1072 ( .A(n1391), .B(n1392), .Z(n1195) );
XNOR2_X1 U1073 ( .A(n1359), .B(n1393), .ZN(n1392) );
NOR2_X1 U1074 ( .A1(G101), .A2(KEYINPUT49), .ZN(n1393) );
INV_X1 U1075 ( .A(G104), .ZN(n1359) );
NAND2_X1 U1076 ( .A1(KEYINPUT3), .A2(n1394), .ZN(n1391) );
INV_X1 U1077 ( .A(n1360), .ZN(n1394) );
INV_X1 U1078 ( .A(n1199), .ZN(n1390) );
XNOR2_X1 U1079 ( .A(n1395), .B(n1396), .ZN(n1199) );
NOR2_X1 U1080 ( .A1(KEYINPUT15), .A2(n1397), .ZN(n1396) );
XNOR2_X1 U1081 ( .A(G113), .B(G119), .ZN(n1395) );
XNOR2_X1 U1082 ( .A(G110), .B(G122), .ZN(n1198) );
NAND2_X1 U1083 ( .A1(n1398), .A2(n1134), .ZN(n1343) );
NAND2_X1 U1084 ( .A1(G237), .A2(G234), .ZN(n1134) );
NAND2_X1 U1085 ( .A1(n1334), .A2(n1399), .ZN(n1398) );
NAND2_X1 U1086 ( .A1(G902), .A2(n1194), .ZN(n1399) );
NOR2_X1 U1087 ( .A1(G898), .A2(n1157), .ZN(n1194) );
NAND2_X1 U1088 ( .A1(G952), .A2(n1400), .ZN(n1334) );
XNOR2_X1 U1089 ( .A(KEYINPUT19), .B(n1157), .ZN(n1400) );
NOR2_X1 U1090 ( .A1(n1308), .A2(n1307), .ZN(n1137) );
XNOR2_X1 U1091 ( .A(n1401), .B(G475), .ZN(n1307) );
NAND2_X1 U1092 ( .A1(n1214), .A2(n1254), .ZN(n1401) );
XNOR2_X1 U1093 ( .A(n1402), .B(n1403), .ZN(n1214) );
XNOR2_X1 U1094 ( .A(n1404), .B(n1405), .ZN(n1403) );
NOR2_X1 U1095 ( .A1(G113), .A2(KEYINPUT0), .ZN(n1405) );
NAND2_X1 U1096 ( .A1(n1406), .A2(KEYINPUT34), .ZN(n1404) );
XOR2_X1 U1097 ( .A(n1407), .B(n1408), .Z(n1406) );
XOR2_X1 U1098 ( .A(n1357), .B(n1170), .Z(n1408) );
XNOR2_X1 U1099 ( .A(n1409), .B(n1318), .ZN(n1407) );
INV_X1 U1100 ( .A(G131), .ZN(n1318) );
NAND2_X1 U1101 ( .A1(G214), .A2(n1410), .ZN(n1409) );
XNOR2_X1 U1102 ( .A(G104), .B(G122), .ZN(n1402) );
XNOR2_X1 U1103 ( .A(n1411), .B(G478), .ZN(n1308) );
NAND2_X1 U1104 ( .A1(n1210), .A2(n1254), .ZN(n1411) );
XNOR2_X1 U1105 ( .A(n1412), .B(n1413), .ZN(n1210) );
XNOR2_X1 U1106 ( .A(n1414), .B(n1415), .ZN(n1413) );
XOR2_X1 U1107 ( .A(G143), .B(G134), .Z(n1415) );
XOR2_X1 U1108 ( .A(n1416), .B(n1417), .Z(n1412) );
AND2_X1 U1109 ( .A1(n1418), .A2(G217), .ZN(n1417) );
NAND2_X1 U1110 ( .A1(n1419), .A2(n1420), .ZN(n1416) );
NAND2_X1 U1111 ( .A1(n1421), .A2(n1360), .ZN(n1420) );
XOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1422), .Z(n1419) );
NOR2_X1 U1113 ( .A1(n1360), .A2(n1421), .ZN(n1422) );
XNOR2_X1 U1114 ( .A(G122), .B(n1397), .ZN(n1421) );
INV_X1 U1115 ( .A(G116), .ZN(n1397) );
XOR2_X1 U1116 ( .A(G107), .B(KEYINPUT31), .Z(n1360) );
NOR2_X1 U1117 ( .A1(n1338), .A2(n1337), .ZN(n1115) );
XNOR2_X1 U1118 ( .A(n1423), .B(n1150), .ZN(n1337) );
NAND2_X1 U1119 ( .A1(G217), .A2(n1366), .ZN(n1150) );
NAND2_X1 U1120 ( .A1(G234), .A2(n1254), .ZN(n1366) );
XNOR2_X1 U1121 ( .A(n1148), .B(KEYINPUT8), .ZN(n1423) );
NOR2_X1 U1122 ( .A1(n1205), .A2(G902), .ZN(n1148) );
XNOR2_X1 U1123 ( .A(n1424), .B(n1425), .ZN(n1205) );
XOR2_X1 U1124 ( .A(KEYINPUT56), .B(KEYINPUT39), .Z(n1425) );
XNOR2_X1 U1125 ( .A(n1426), .B(n1427), .ZN(n1424) );
INV_X1 U1126 ( .A(G110), .ZN(n1427) );
XOR2_X1 U1127 ( .A(n1428), .B(n1429), .Z(n1426) );
XNOR2_X1 U1128 ( .A(n1414), .B(n1430), .ZN(n1429) );
XOR2_X1 U1129 ( .A(G146), .B(G137), .Z(n1430) );
INV_X1 U1130 ( .A(G128), .ZN(n1414) );
XOR2_X1 U1131 ( .A(n1431), .B(n1432), .Z(n1428) );
NOR2_X1 U1132 ( .A1(n1433), .A2(n1434), .ZN(n1432) );
AND3_X1 U1133 ( .A1(KEYINPUT6), .A2(n1302), .A3(G140), .ZN(n1434) );
INV_X1 U1134 ( .A(G125), .ZN(n1302) );
NOR2_X1 U1135 ( .A1(KEYINPUT6), .A2(n1170), .ZN(n1433) );
XNOR2_X1 U1136 ( .A(n1169), .B(G125), .ZN(n1170) );
INV_X1 U1137 ( .A(G140), .ZN(n1169) );
XNOR2_X1 U1138 ( .A(n1435), .B(n1436), .ZN(n1431) );
INV_X1 U1139 ( .A(G119), .ZN(n1436) );
NAND2_X1 U1140 ( .A1(G221), .A2(n1418), .ZN(n1435) );
AND2_X1 U1141 ( .A1(G234), .A2(n1157), .ZN(n1418) );
INV_X1 U1142 ( .A(G953), .ZN(n1157) );
XOR2_X1 U1143 ( .A(G472), .B(n1437), .Z(n1338) );
NOR2_X1 U1144 ( .A1(KEYINPUT14), .A2(n1147), .ZN(n1437) );
NAND2_X1 U1145 ( .A1(n1438), .A2(n1254), .ZN(n1147) );
INV_X1 U1146 ( .A(G902), .ZN(n1254) );
XOR2_X1 U1147 ( .A(n1439), .B(n1440), .Z(n1438) );
XNOR2_X1 U1148 ( .A(n1231), .B(n1245), .ZN(n1440) );
XNOR2_X1 U1149 ( .A(n1441), .B(n1442), .ZN(n1245) );
NOR2_X1 U1150 ( .A1(G113), .A2(KEYINPUT61), .ZN(n1442) );
XNOR2_X1 U1151 ( .A(G116), .B(n1443), .ZN(n1441) );
NOR2_X1 U1152 ( .A1(G119), .A2(KEYINPUT29), .ZN(n1443) );
XOR2_X1 U1153 ( .A(G128), .B(n1357), .Z(n1231) );
XOR2_X1 U1154 ( .A(G143), .B(G146), .Z(n1357) );
XNOR2_X1 U1155 ( .A(n1353), .B(n1225), .ZN(n1439) );
NAND2_X1 U1156 ( .A1(G210), .A2(n1410), .ZN(n1225) );
NOR2_X1 U1157 ( .A1(G953), .A2(G237), .ZN(n1410) );
XNOR2_X1 U1158 ( .A(n1244), .B(n1226), .ZN(n1353) );
INV_X1 U1159 ( .A(G101), .ZN(n1226) );
NAND2_X1 U1160 ( .A1(n1444), .A2(n1445), .ZN(n1244) );
NAND2_X1 U1161 ( .A1(G131), .A2(n1165), .ZN(n1445) );
XOR2_X1 U1162 ( .A(KEYINPUT50), .B(n1446), .Z(n1444) );
NOR2_X1 U1163 ( .A1(G131), .A2(n1165), .ZN(n1446) );
XOR2_X1 U1164 ( .A(G137), .B(G134), .Z(n1165) );
endmodule


