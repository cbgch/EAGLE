//Key = 1100101011111000001011110100001100010011100010100100000111110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;

XOR2_X1 U771 ( .A(n1069), .B(n1070), .Z(G9) );
NOR2_X1 U772 ( .A1(G107), .A2(KEYINPUT51), .ZN(n1070) );
NAND3_X1 U773 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1069) );
XNOR2_X1 U774 ( .A(n1074), .B(KEYINPUT49), .ZN(n1073) );
NOR2_X1 U775 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR4_X1 U776 ( .A1(G953), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1076) );
NOR2_X1 U777 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR3_X1 U779 ( .A1(n1084), .A2(n1085), .A3(n1086), .ZN(n1083) );
NOR2_X1 U780 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
NOR2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NOR3_X1 U782 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1089) );
AND2_X1 U783 ( .A1(n1094), .A2(KEYINPUT54), .ZN(n1093) );
NOR4_X1 U784 ( .A1(KEYINPUT54), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1092) );
INV_X1 U785 ( .A(n1098), .ZN(n1096) );
NOR2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1087) );
NOR2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
AND2_X1 U788 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR3_X1 U789 ( .A1(n1100), .A2(n1105), .A3(n1090), .ZN(n1082) );
NOR2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U791 ( .A1(n1108), .A2(n1084), .ZN(n1107) );
INV_X1 U792 ( .A(n1109), .ZN(n1084) );
NOR2_X1 U793 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR2_X1 U794 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NOR2_X1 U795 ( .A1(n1114), .A2(n1086), .ZN(n1106) );
INV_X1 U796 ( .A(n1074), .ZN(n1086) );
NOR2_X1 U797 ( .A1(n1071), .A2(n1115), .ZN(n1114) );
NOR3_X1 U798 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1075) );
AND4_X1 U799 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1077) );
NOR4_X1 U800 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1119) );
XNOR2_X1 U801 ( .A(KEYINPUT43), .B(n1098), .ZN(n1123) );
XOR2_X1 U802 ( .A(n1103), .B(KEYINPUT10), .Z(n1120) );
AND3_X1 U803 ( .A1(n1095), .A2(n1124), .A3(n1125), .ZN(n1118) );
XNOR2_X1 U804 ( .A(n1126), .B(n1127), .ZN(n1117) );
NAND2_X1 U805 ( .A1(KEYINPUT8), .A2(n1128), .ZN(n1127) );
XOR2_X1 U806 ( .A(KEYINPUT37), .B(n1129), .Z(n1116) );
NOR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XNOR2_X1 U808 ( .A(KEYINPUT24), .B(n1132), .ZN(n1131) );
INV_X1 U809 ( .A(n1133), .ZN(n1130) );
XOR2_X1 U810 ( .A(n1134), .B(n1135), .Z(G72) );
XOR2_X1 U811 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U812 ( .A1(G953), .A2(n1138), .ZN(n1137) );
NAND2_X1 U813 ( .A1(G900), .A2(G227), .ZN(n1138) );
NAND2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1136) );
NAND2_X1 U815 ( .A1(G953), .A2(n1141), .ZN(n1140) );
XOR2_X1 U816 ( .A(n1142), .B(n1143), .Z(n1139) );
XNOR2_X1 U817 ( .A(n1144), .B(n1145), .ZN(n1143) );
XOR2_X1 U818 ( .A(KEYINPUT47), .B(G140), .Z(n1145) );
XOR2_X1 U819 ( .A(n1146), .B(n1147), .Z(n1142) );
XOR2_X1 U820 ( .A(n1148), .B(n1149), .Z(n1146) );
NAND2_X1 U821 ( .A1(KEYINPUT59), .A2(n1150), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1151), .A2(G953), .ZN(n1134) );
NAND3_X1 U823 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(G69) );
XOR2_X1 U824 ( .A(n1155), .B(KEYINPUT29), .Z(n1154) );
NAND3_X1 U825 ( .A1(G953), .A2(n1156), .A3(n1157), .ZN(n1155) );
INV_X1 U826 ( .A(n1158), .ZN(n1157) );
NAND2_X1 U827 ( .A1(G898), .A2(G224), .ZN(n1156) );
NAND2_X1 U828 ( .A1(n1159), .A2(n1160), .ZN(n1153) );
NAND2_X1 U829 ( .A1(n1161), .A2(n1162), .ZN(n1159) );
NAND2_X1 U830 ( .A1(n1163), .A2(n1158), .ZN(n1162) );
NAND2_X1 U831 ( .A1(n1164), .A2(n1165), .ZN(n1161) );
XOR2_X1 U832 ( .A(n1166), .B(KEYINPUT16), .Z(n1164) );
NAND4_X1 U833 ( .A1(G224), .A2(n1158), .A3(G898), .A4(G953), .ZN(n1152) );
XNOR2_X1 U834 ( .A(n1166), .B(KEYINPUT45), .ZN(n1158) );
NAND2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U836 ( .A1(G953), .A2(n1169), .ZN(n1168) );
XOR2_X1 U837 ( .A(n1170), .B(n1171), .Z(n1167) );
NAND2_X1 U838 ( .A1(KEYINPUT4), .A2(n1172), .ZN(n1170) );
NOR2_X1 U839 ( .A1(n1173), .A2(n1174), .ZN(G66) );
XNOR2_X1 U840 ( .A(n1175), .B(n1176), .ZN(n1174) );
AND3_X1 U841 ( .A1(n1177), .A2(n1178), .A3(G217), .ZN(n1175) );
NOR2_X1 U842 ( .A1(n1173), .A2(n1179), .ZN(G63) );
XOR2_X1 U843 ( .A(n1180), .B(n1181), .Z(n1179) );
AND2_X1 U844 ( .A1(G478), .A2(n1177), .ZN(n1181) );
NOR2_X1 U845 ( .A1(KEYINPUT19), .A2(n1182), .ZN(n1180) );
NOR2_X1 U846 ( .A1(n1173), .A2(n1183), .ZN(G60) );
NOR3_X1 U847 ( .A1(n1126), .A2(n1184), .A3(n1185), .ZN(n1183) );
NOR3_X1 U848 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
AND2_X1 U849 ( .A1(n1186), .A2(n1187), .ZN(n1184) );
NAND3_X1 U850 ( .A1(G475), .A2(n1079), .A3(KEYINPUT55), .ZN(n1186) );
XNOR2_X1 U851 ( .A(G104), .B(n1189), .ZN(G6) );
NOR2_X1 U852 ( .A1(n1173), .A2(n1190), .ZN(G57) );
XOR2_X1 U853 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U854 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U855 ( .A1(n1195), .A2(KEYINPUT2), .ZN(n1194) );
AND2_X1 U856 ( .A1(G472), .A2(n1177), .ZN(n1193) );
XNOR2_X1 U857 ( .A(n1196), .B(n1197), .ZN(n1191) );
NAND3_X1 U858 ( .A1(n1198), .A2(n1199), .A3(KEYINPUT44), .ZN(n1196) );
NAND2_X1 U859 ( .A1(KEYINPUT1), .A2(n1200), .ZN(n1199) );
NAND3_X1 U860 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1198) );
INV_X1 U861 ( .A(KEYINPUT1), .ZN(n1203) );
NOR2_X1 U862 ( .A1(n1173), .A2(n1204), .ZN(G54) );
XOR2_X1 U863 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U864 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U865 ( .A1(KEYINPUT3), .A2(n1209), .ZN(n1208) );
AND2_X1 U866 ( .A1(G469), .A2(n1177), .ZN(n1207) );
XOR2_X1 U867 ( .A(n1210), .B(n1211), .Z(n1205) );
NOR2_X1 U868 ( .A1(n1173), .A2(n1212), .ZN(G51) );
XOR2_X1 U869 ( .A(n1213), .B(n1214), .Z(n1212) );
NOR2_X1 U870 ( .A1(KEYINPUT17), .A2(n1215), .ZN(n1214) );
XOR2_X1 U871 ( .A(n1216), .B(n1217), .Z(n1215) );
XNOR2_X1 U872 ( .A(n1218), .B(KEYINPUT20), .ZN(n1217) );
NAND2_X1 U873 ( .A1(n1219), .A2(KEYINPUT11), .ZN(n1218) );
XNOR2_X1 U874 ( .A(n1220), .B(n1144), .ZN(n1219) );
NAND2_X1 U875 ( .A1(KEYINPUT23), .A2(n1221), .ZN(n1220) );
NAND2_X1 U876 ( .A1(n1177), .A2(n1222), .ZN(n1213) );
AND2_X1 U877 ( .A1(G902), .A2(n1079), .ZN(n1177) );
NAND2_X1 U878 ( .A1(n1163), .A2(n1151), .ZN(n1079) );
AND4_X1 U879 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1151) );
NOR4_X1 U880 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1226) );
NOR3_X1 U881 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1225) );
NOR4_X1 U882 ( .A1(n1234), .A2(n1235), .A3(n1102), .A4(n1100), .ZN(n1233) );
INV_X1 U883 ( .A(KEYINPUT48), .ZN(n1234) );
NOR2_X1 U884 ( .A1(KEYINPUT48), .A2(n1236), .ZN(n1232) );
INV_X1 U885 ( .A(n1165), .ZN(n1163) );
NAND4_X1 U886 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1165) );
AND4_X1 U887 ( .A1(n1189), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1240) );
NAND3_X1 U888 ( .A1(n1072), .A2(n1074), .A3(n1115), .ZN(n1189) );
NOR2_X1 U889 ( .A1(n1244), .A2(n1245), .ZN(n1239) );
AND3_X1 U890 ( .A1(n1071), .A2(n1074), .A3(n1072), .ZN(n1245) );
INV_X1 U891 ( .A(n1246), .ZN(n1244) );
NOR2_X1 U892 ( .A1(n1160), .A2(G952), .ZN(n1173) );
NAND2_X1 U893 ( .A1(n1247), .A2(n1248), .ZN(G48) );
NAND2_X1 U894 ( .A1(G146), .A2(n1249), .ZN(n1248) );
NAND2_X1 U895 ( .A1(n1230), .A2(n1250), .ZN(n1249) );
NAND2_X1 U896 ( .A1(KEYINPUT32), .A2(KEYINPUT18), .ZN(n1250) );
NAND3_X1 U897 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1247) );
INV_X1 U898 ( .A(KEYINPUT32), .ZN(n1253) );
NAND2_X1 U899 ( .A1(n1230), .A2(n1254), .ZN(n1252) );
INV_X1 U900 ( .A(KEYINPUT18), .ZN(n1254) );
NAND2_X1 U901 ( .A1(KEYINPUT18), .A2(n1255), .ZN(n1251) );
NAND2_X1 U902 ( .A1(n1230), .A2(n1256), .ZN(n1255) );
AND3_X1 U903 ( .A1(n1115), .A2(n1091), .A3(n1257), .ZN(n1230) );
XOR2_X1 U904 ( .A(G143), .B(n1229), .Z(G45) );
AND4_X1 U905 ( .A1(n1102), .A2(n1091), .A3(n1111), .A4(n1258), .ZN(n1229) );
AND3_X1 U906 ( .A1(n1122), .A2(n1259), .A3(n1260), .ZN(n1258) );
XNOR2_X1 U907 ( .A(G140), .B(n1236), .ZN(G42) );
NAND3_X1 U908 ( .A1(n1094), .A2(n1102), .A3(n1261), .ZN(n1236) );
XOR2_X1 U909 ( .A(G137), .B(n1228), .Z(G39) );
AND3_X1 U910 ( .A1(n1257), .A2(n1109), .A3(n1094), .ZN(n1228) );
XNOR2_X1 U911 ( .A(n1150), .B(n1231), .ZN(G36) );
AND2_X1 U912 ( .A1(n1262), .A2(n1071), .ZN(n1231) );
XNOR2_X1 U913 ( .A(G131), .B(n1223), .ZN(G33) );
NAND2_X1 U914 ( .A1(n1262), .A2(n1115), .ZN(n1223) );
AND4_X1 U915 ( .A1(n1094), .A2(n1111), .A3(n1102), .A4(n1259), .ZN(n1262) );
INV_X1 U916 ( .A(n1100), .ZN(n1094) );
NAND3_X1 U917 ( .A1(n1125), .A2(n1098), .A3(n1095), .ZN(n1100) );
XNOR2_X1 U918 ( .A(n1263), .B(n1227), .ZN(G30) );
AND3_X1 U919 ( .A1(n1071), .A2(n1091), .A3(n1257), .ZN(n1227) );
AND4_X1 U920 ( .A1(n1102), .A2(n1121), .A3(n1259), .A4(n1264), .ZN(n1257) );
XNOR2_X1 U921 ( .A(G101), .B(n1246), .ZN(G3) );
NAND3_X1 U922 ( .A1(n1109), .A2(n1072), .A3(n1111), .ZN(n1246) );
NAND2_X1 U923 ( .A1(n1265), .A2(n1266), .ZN(G27) );
NAND2_X1 U924 ( .A1(n1267), .A2(n1144), .ZN(n1266) );
XOR2_X1 U925 ( .A(n1224), .B(KEYINPUT0), .Z(n1267) );
NAND2_X1 U926 ( .A1(n1268), .A2(G125), .ZN(n1265) );
XNOR2_X1 U927 ( .A(KEYINPUT12), .B(n1224), .ZN(n1268) );
NAND3_X1 U928 ( .A1(n1269), .A2(n1091), .A3(n1261), .ZN(n1224) );
INV_X1 U929 ( .A(n1235), .ZN(n1261) );
NAND4_X1 U930 ( .A1(n1115), .A2(n1270), .A3(n1259), .A4(n1264), .ZN(n1235) );
NAND2_X1 U931 ( .A1(n1081), .A2(n1271), .ZN(n1259) );
NAND4_X1 U932 ( .A1(G902), .A2(G953), .A3(n1272), .A4(n1141), .ZN(n1271) );
INV_X1 U933 ( .A(G900), .ZN(n1141) );
XNOR2_X1 U934 ( .A(G122), .B(n1237), .ZN(G24) );
NAND4_X1 U935 ( .A1(n1273), .A2(n1074), .A3(n1122), .A4(n1260), .ZN(n1237) );
NOR2_X1 U936 ( .A1(n1264), .A2(n1113), .ZN(n1074) );
INV_X1 U937 ( .A(n1270), .ZN(n1113) );
NAND2_X1 U938 ( .A1(n1274), .A2(n1275), .ZN(G21) );
NAND2_X1 U939 ( .A1(n1276), .A2(n1238), .ZN(n1275) );
NAND2_X1 U940 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U941 ( .A1(KEYINPUT28), .A2(n1279), .ZN(n1278) );
NAND3_X1 U942 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1274) );
INV_X1 U943 ( .A(KEYINPUT28), .ZN(n1282) );
NAND2_X1 U944 ( .A1(G119), .A2(n1279), .ZN(n1281) );
INV_X1 U945 ( .A(KEYINPUT13), .ZN(n1279) );
NAND2_X1 U946 ( .A1(n1283), .A2(n1277), .ZN(n1280) );
OR2_X1 U947 ( .A1(n1238), .A2(KEYINPUT13), .ZN(n1283) );
NAND4_X1 U948 ( .A1(n1273), .A2(n1109), .A3(n1121), .A4(n1264), .ZN(n1238) );
XNOR2_X1 U949 ( .A(G116), .B(n1243), .ZN(G18) );
NAND3_X1 U950 ( .A1(n1111), .A2(n1071), .A3(n1273), .ZN(n1243) );
NOR2_X1 U951 ( .A1(n1260), .A2(n1284), .ZN(n1071) );
INV_X1 U952 ( .A(n1122), .ZN(n1284) );
NAND2_X1 U953 ( .A1(n1285), .A2(n1286), .ZN(G15) );
NAND2_X1 U954 ( .A1(G113), .A2(n1242), .ZN(n1286) );
XOR2_X1 U955 ( .A(KEYINPUT57), .B(n1287), .Z(n1285) );
NOR2_X1 U956 ( .A1(G113), .A2(n1242), .ZN(n1287) );
NAND3_X1 U957 ( .A1(n1111), .A2(n1115), .A3(n1273), .ZN(n1242) );
AND3_X1 U958 ( .A1(n1091), .A2(n1288), .A3(n1269), .ZN(n1273) );
INV_X1 U959 ( .A(n1090), .ZN(n1269) );
NAND2_X1 U960 ( .A1(n1103), .A2(n1124), .ZN(n1090) );
NOR2_X1 U961 ( .A1(n1122), .A2(n1289), .ZN(n1115) );
INV_X1 U962 ( .A(n1260), .ZN(n1289) );
AND2_X1 U963 ( .A1(n1112), .A2(n1121), .ZN(n1111) );
INV_X1 U964 ( .A(n1264), .ZN(n1112) );
XNOR2_X1 U965 ( .A(G110), .B(n1241), .ZN(G12) );
NAND4_X1 U966 ( .A1(n1109), .A2(n1072), .A3(n1270), .A4(n1264), .ZN(n1241) );
NAND2_X1 U967 ( .A1(n1133), .A2(n1132), .ZN(n1264) );
NAND3_X1 U968 ( .A1(n1290), .A2(n1188), .A3(n1176), .ZN(n1132) );
NAND2_X1 U969 ( .A1(G217), .A2(n1178), .ZN(n1290) );
NAND3_X1 U970 ( .A1(n1291), .A2(n1178), .A3(G217), .ZN(n1133) );
NAND2_X1 U971 ( .A1(n1176), .A2(n1188), .ZN(n1291) );
XOR2_X1 U972 ( .A(n1292), .B(n1293), .Z(n1176) );
XOR2_X1 U973 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U974 ( .A(n1296), .B(n1297), .Z(n1295) );
NOR2_X1 U975 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XOR2_X1 U976 ( .A(n1300), .B(KEYINPUT31), .Z(n1299) );
NAND2_X1 U977 ( .A1(G119), .A2(n1263), .ZN(n1300) );
NOR2_X1 U978 ( .A1(G119), .A2(n1263), .ZN(n1298) );
NAND2_X1 U979 ( .A1(G221), .A2(n1301), .ZN(n1296) );
NAND2_X1 U980 ( .A1(KEYINPUT35), .A2(n1302), .ZN(n1294) );
INV_X1 U981 ( .A(G110), .ZN(n1302) );
XOR2_X1 U982 ( .A(n1303), .B(n1304), .Z(n1292) );
XOR2_X1 U983 ( .A(G137), .B(n1305), .Z(n1304) );
XNOR2_X1 U984 ( .A(G146), .B(KEYINPUT60), .ZN(n1303) );
XOR2_X1 U985 ( .A(n1121), .B(KEYINPUT56), .Z(n1270) );
XNOR2_X1 U986 ( .A(n1306), .B(G472), .ZN(n1121) );
NAND2_X1 U987 ( .A1(n1307), .A2(n1188), .ZN(n1306) );
XOR2_X1 U988 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U989 ( .A(n1200), .B(n1195), .Z(n1309) );
AND3_X1 U990 ( .A1(n1310), .A2(n1311), .A3(G210), .ZN(n1195) );
XOR2_X1 U991 ( .A(n1202), .B(n1201), .Z(n1200) );
XNOR2_X1 U992 ( .A(n1312), .B(n1313), .ZN(n1201) );
XOR2_X1 U993 ( .A(G116), .B(G113), .Z(n1313) );
NAND2_X1 U994 ( .A1(KEYINPUT40), .A2(n1277), .ZN(n1312) );
INV_X1 U995 ( .A(G119), .ZN(n1277) );
XNOR2_X1 U996 ( .A(n1210), .B(n1221), .ZN(n1202) );
XNOR2_X1 U997 ( .A(n1314), .B(n1197), .ZN(n1308) );
XNOR2_X1 U998 ( .A(KEYINPUT53), .B(KEYINPUT38), .ZN(n1314) );
AND3_X1 U999 ( .A1(n1091), .A2(n1288), .A3(n1102), .ZN(n1072) );
NOR2_X1 U1000 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
INV_X1 U1001 ( .A(n1124), .ZN(n1104) );
NAND2_X1 U1002 ( .A1(G221), .A2(n1178), .ZN(n1124) );
NAND2_X1 U1003 ( .A1(n1315), .A2(G234), .ZN(n1178) );
XOR2_X1 U1004 ( .A(n1316), .B(G469), .Z(n1103) );
NAND2_X1 U1005 ( .A1(n1317), .A2(n1188), .ZN(n1316) );
XOR2_X1 U1006 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1007 ( .A(n1209), .B(n1320), .Z(n1319) );
NAND2_X1 U1008 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
OR2_X1 U1009 ( .A1(n1211), .A2(KEYINPUT15), .ZN(n1322) );
XNOR2_X1 U1010 ( .A(n1323), .B(n1324), .ZN(n1211) );
NAND2_X1 U1011 ( .A1(n1325), .A2(n1326), .ZN(n1323) );
NAND2_X1 U1012 ( .A1(n1327), .A2(n1147), .ZN(n1326) );
NAND2_X1 U1013 ( .A1(KEYINPUT15), .A2(n1328), .ZN(n1321) );
XOR2_X1 U1014 ( .A(n1325), .B(n1324), .Z(n1328) );
AND2_X1 U1015 ( .A1(G227), .A2(n1310), .ZN(n1324) );
OR2_X1 U1016 ( .A1(n1147), .A2(n1327), .ZN(n1325) );
XOR2_X1 U1017 ( .A(G101), .B(n1329), .Z(n1327) );
NOR2_X1 U1018 ( .A1(KEYINPUT41), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1019 ( .A(n1331), .B(n1263), .Z(n1147) );
NAND2_X1 U1020 ( .A1(KEYINPUT21), .A2(n1332), .ZN(n1331) );
XNOR2_X1 U1021 ( .A(n1256), .B(G143), .ZN(n1332) );
XNOR2_X1 U1022 ( .A(G110), .B(G140), .ZN(n1209) );
XOR2_X1 U1023 ( .A(n1210), .B(KEYINPUT58), .Z(n1318) );
XOR2_X1 U1024 ( .A(n1333), .B(n1149), .Z(n1210) );
XOR2_X1 U1025 ( .A(G131), .B(n1334), .Z(n1149) );
XOR2_X1 U1026 ( .A(KEYINPUT9), .B(G137), .Z(n1334) );
NAND2_X1 U1027 ( .A1(KEYINPUT61), .A2(n1150), .ZN(n1333) );
NAND2_X1 U1028 ( .A1(n1335), .A2(n1081), .ZN(n1288) );
NAND3_X1 U1029 ( .A1(n1272), .A2(n1160), .A3(G952), .ZN(n1081) );
XOR2_X1 U1030 ( .A(KEYINPUT22), .B(n1336), .Z(n1335) );
AND4_X1 U1031 ( .A1(n1169), .A2(n1272), .A3(G953), .A4(G902), .ZN(n1336) );
NAND2_X1 U1032 ( .A1(G237), .A2(G234), .ZN(n1272) );
INV_X1 U1033 ( .A(G898), .ZN(n1169) );
AND2_X1 U1034 ( .A1(n1337), .A2(n1095), .ZN(n1091) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1338), .ZN(n1095) );
NAND2_X1 U1036 ( .A1(n1098), .A2(n1125), .ZN(n1337) );
INV_X1 U1037 ( .A(n1097), .ZN(n1125) );
NOR2_X1 U1038 ( .A1(n1339), .A2(n1222), .ZN(n1097) );
NAND2_X1 U1039 ( .A1(n1222), .A2(n1339), .ZN(n1098) );
NAND2_X1 U1040 ( .A1(n1340), .A2(n1188), .ZN(n1339) );
XOR2_X1 U1041 ( .A(n1216), .B(n1341), .Z(n1340) );
XNOR2_X1 U1042 ( .A(G125), .B(n1221), .ZN(n1341) );
XNOR2_X1 U1043 ( .A(G146), .B(n1342), .ZN(n1221) );
XNOR2_X1 U1044 ( .A(n1171), .B(n1343), .ZN(n1216) );
XOR2_X1 U1045 ( .A(n1172), .B(n1344), .Z(n1343) );
NAND2_X1 U1046 ( .A1(G224), .A2(n1310), .ZN(n1344) );
NAND3_X1 U1047 ( .A1(n1345), .A2(n1346), .A3(n1347), .ZN(n1172) );
NAND2_X1 U1048 ( .A1(KEYINPUT52), .A2(G110), .ZN(n1347) );
NAND3_X1 U1049 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1346) );
INV_X1 U1050 ( .A(KEYINPUT52), .ZN(n1349) );
OR2_X1 U1051 ( .A1(n1350), .A2(n1348), .ZN(n1345) );
NOR2_X1 U1052 ( .A1(G110), .A2(KEYINPUT63), .ZN(n1348) );
XOR2_X1 U1053 ( .A(n1351), .B(n1352), .Z(n1171) );
XOR2_X1 U1054 ( .A(n1353), .B(n1354), .Z(n1352) );
NAND2_X1 U1055 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1056 ( .A1(KEYINPUT30), .A2(n1330), .ZN(n1356) );
XNOR2_X1 U1057 ( .A(G104), .B(G107), .ZN(n1330) );
OR3_X1 U1058 ( .A1(n1357), .A2(G107), .A3(KEYINPUT30), .ZN(n1355) );
NAND2_X1 U1059 ( .A1(KEYINPUT39), .A2(n1197), .ZN(n1353) );
INV_X1 U1060 ( .A(G101), .ZN(n1197) );
XOR2_X1 U1061 ( .A(n1358), .B(n1359), .Z(n1351) );
NOR2_X1 U1062 ( .A1(KEYINPUT42), .A2(n1360), .ZN(n1359) );
XOR2_X1 U1063 ( .A(G116), .B(n1361), .Z(n1360) );
NOR2_X1 U1064 ( .A1(G119), .A2(KEYINPUT50), .ZN(n1361) );
XNOR2_X1 U1065 ( .A(G113), .B(KEYINPUT25), .ZN(n1358) );
AND2_X1 U1066 ( .A1(G210), .A2(n1338), .ZN(n1222) );
NAND2_X1 U1067 ( .A1(n1315), .A2(n1311), .ZN(n1338) );
XNOR2_X1 U1068 ( .A(G902), .B(KEYINPUT27), .ZN(n1315) );
NOR2_X1 U1069 ( .A1(n1122), .A2(n1260), .ZN(n1109) );
XOR2_X1 U1070 ( .A(n1126), .B(n1362), .Z(n1260) );
XNOR2_X1 U1071 ( .A(KEYINPUT5), .B(n1128), .ZN(n1362) );
INV_X1 U1072 ( .A(G475), .ZN(n1128) );
AND2_X1 U1073 ( .A1(n1187), .A2(n1188), .ZN(n1126) );
XNOR2_X1 U1074 ( .A(n1363), .B(n1364), .ZN(n1187) );
XOR2_X1 U1075 ( .A(n1365), .B(n1366), .Z(n1364) );
NAND2_X1 U1076 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
NAND2_X1 U1077 ( .A1(G146), .A2(n1369), .ZN(n1368) );
NAND2_X1 U1078 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
NAND2_X1 U1079 ( .A1(n1372), .A2(n1144), .ZN(n1371) );
XNOR2_X1 U1080 ( .A(n1373), .B(n1374), .ZN(n1370) );
NAND2_X1 U1081 ( .A1(n1375), .A2(n1256), .ZN(n1367) );
INV_X1 U1082 ( .A(G146), .ZN(n1256) );
NAND2_X1 U1083 ( .A1(n1376), .A2(n1377), .ZN(n1375) );
NAND2_X1 U1084 ( .A1(n1374), .A2(n1373), .ZN(n1377) );
INV_X1 U1085 ( .A(KEYINPUT46), .ZN(n1373) );
NAND2_X1 U1086 ( .A1(n1305), .A2(KEYINPUT46), .ZN(n1376) );
NOR2_X1 U1087 ( .A1(n1378), .A2(n1374), .ZN(n1305) );
NOR2_X1 U1088 ( .A1(n1144), .A2(n1372), .ZN(n1374) );
AND2_X1 U1089 ( .A1(n1372), .A2(n1144), .ZN(n1378) );
INV_X1 U1090 ( .A(G125), .ZN(n1144) );
XOR2_X1 U1091 ( .A(G140), .B(KEYINPUT14), .Z(n1372) );
NAND2_X1 U1092 ( .A1(n1379), .A2(n1380), .ZN(n1365) );
NAND2_X1 U1093 ( .A1(n1381), .A2(n1382), .ZN(n1380) );
XOR2_X1 U1094 ( .A(n1383), .B(KEYINPUT34), .Z(n1379) );
OR2_X1 U1095 ( .A1(n1382), .A2(n1381), .ZN(n1383) );
XNOR2_X1 U1096 ( .A(G143), .B(n1384), .ZN(n1381) );
AND3_X1 U1097 ( .A1(G214), .A2(n1311), .A3(n1310), .ZN(n1384) );
INV_X1 U1098 ( .A(G237), .ZN(n1311) );
XOR2_X1 U1099 ( .A(G131), .B(KEYINPUT36), .Z(n1382) );
XNOR2_X1 U1100 ( .A(n1385), .B(n1357), .ZN(n1363) );
INV_X1 U1101 ( .A(G104), .ZN(n1357) );
NAND2_X1 U1102 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
NAND2_X1 U1103 ( .A1(G113), .A2(n1350), .ZN(n1387) );
XOR2_X1 U1104 ( .A(n1388), .B(KEYINPUT33), .Z(n1386) );
OR2_X1 U1105 ( .A1(n1350), .A2(G113), .ZN(n1388) );
INV_X1 U1106 ( .A(G122), .ZN(n1350) );
XNOR2_X1 U1107 ( .A(n1389), .B(G478), .ZN(n1122) );
NAND2_X1 U1108 ( .A1(n1182), .A2(n1188), .ZN(n1389) );
INV_X1 U1109 ( .A(G902), .ZN(n1188) );
XNOR2_X1 U1110 ( .A(n1390), .B(n1391), .ZN(n1182) );
XOR2_X1 U1111 ( .A(n1392), .B(n1393), .Z(n1391) );
NAND2_X1 U1112 ( .A1(G217), .A2(n1301), .ZN(n1393) );
AND2_X1 U1113 ( .A1(G234), .A2(n1310), .ZN(n1301) );
XOR2_X1 U1114 ( .A(n1160), .B(KEYINPUT26), .Z(n1310) );
INV_X1 U1115 ( .A(G953), .ZN(n1160) );
NAND2_X1 U1116 ( .A1(KEYINPUT62), .A2(n1394), .ZN(n1392) );
XOR2_X1 U1117 ( .A(n1342), .B(n1395), .Z(n1394) );
XNOR2_X1 U1118 ( .A(KEYINPUT7), .B(n1150), .ZN(n1395) );
INV_X1 U1119 ( .A(G134), .ZN(n1150) );
XNOR2_X1 U1120 ( .A(n1263), .B(G143), .ZN(n1342) );
INV_X1 U1121 ( .A(G128), .ZN(n1263) );
XOR2_X1 U1122 ( .A(n1396), .B(n1397), .Z(n1390) );
XOR2_X1 U1123 ( .A(G116), .B(G107), .Z(n1397) );
NAND2_X1 U1124 ( .A1(KEYINPUT6), .A2(G122), .ZN(n1396) );
endmodule


