//Key = 0101001010101111110100101111111010110100011011001000000101100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;

XNOR2_X1 U758 ( .A(G107), .B(n1044), .ZN(G9) );
NAND2_X1 U759 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NOR2_X1 U760 ( .A1(n1047), .A2(n1048), .ZN(G75) );
NOR4_X1 U761 ( .A1(n1049), .A2(n1050), .A3(G953), .A4(n1051), .ZN(n1048) );
NOR3_X1 U762 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1050) );
INV_X1 U763 ( .A(n1055), .ZN(n1054) );
NOR2_X1 U764 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
NOR2_X1 U765 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U766 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U767 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
AND3_X1 U768 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1060) );
NOR4_X1 U769 ( .A1(n1067), .A2(n1068), .A3(n1063), .A4(n1069), .ZN(n1056) );
XNOR2_X1 U770 ( .A(n1066), .B(KEYINPUT4), .ZN(n1068) );
NAND3_X1 U771 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1049) );
XOR2_X1 U772 ( .A(n1073), .B(KEYINPUT25), .Z(n1072) );
NAND2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NAND3_X1 U774 ( .A1(n1076), .A2(n1066), .A3(n1077), .ZN(n1075) );
NAND3_X1 U775 ( .A1(n1055), .A2(n1078), .A3(n1079), .ZN(n1074) );
INV_X1 U776 ( .A(n1052), .ZN(n1079) );
NAND2_X1 U777 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NAND3_X1 U778 ( .A1(n1066), .A2(n1082), .A3(n1083), .ZN(n1081) );
NAND2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1080) );
NAND2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U781 ( .A1(n1088), .A2(n1066), .ZN(n1087) );
XNOR2_X1 U782 ( .A(n1089), .B(KEYINPUT44), .ZN(n1088) );
NAND2_X1 U783 ( .A1(n1083), .A2(n1090), .ZN(n1086) );
NAND2_X1 U784 ( .A1(n1077), .A2(n1046), .ZN(n1071) );
INV_X1 U785 ( .A(n1091), .ZN(n1046) );
NOR3_X1 U786 ( .A1(n1063), .A2(n1059), .A3(n1052), .ZN(n1077) );
NOR3_X1 U787 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1047) );
AND4_X1 U788 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1051) );
NOR4_X1 U789 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1095) );
NOR2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
INV_X1 U791 ( .A(KEYINPUT38), .ZN(n1101) );
NOR2_X1 U792 ( .A1(KEYINPUT38), .A2(n1102), .ZN(n1098) );
XNOR2_X1 U793 ( .A(G469), .B(n1103), .ZN(n1097) );
NAND3_X1 U794 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1096) );
XOR2_X1 U795 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U796 ( .A1(KEYINPUT35), .A2(G475), .ZN(n1107) );
AND3_X1 U797 ( .A1(n1109), .A2(n1110), .A3(n1069), .ZN(n1094) );
NAND2_X1 U798 ( .A1(G478), .A2(n1111), .ZN(n1093) );
XOR2_X1 U799 ( .A(KEYINPUT12), .B(n1112), .Z(n1092) );
XOR2_X1 U800 ( .A(n1113), .B(n1114), .Z(G72) );
XOR2_X1 U801 ( .A(n1115), .B(n1116), .Z(n1114) );
NAND2_X1 U802 ( .A1(G953), .A2(n1117), .ZN(n1116) );
NAND2_X1 U803 ( .A1(G900), .A2(G227), .ZN(n1117) );
NAND3_X1 U804 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(n1115) );
NAND2_X1 U805 ( .A1(G953), .A2(n1121), .ZN(n1120) );
XOR2_X1 U806 ( .A(KEYINPUT15), .B(G900), .Z(n1121) );
NAND2_X1 U807 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
XOR2_X1 U808 ( .A(KEYINPUT24), .B(n1124), .Z(n1122) );
NAND2_X1 U809 ( .A1(n1125), .A2(G125), .ZN(n1118) );
XOR2_X1 U810 ( .A(KEYINPUT11), .B(n1124), .Z(n1125) );
XNOR2_X1 U811 ( .A(n1126), .B(G140), .ZN(n1124) );
NAND2_X1 U812 ( .A1(KEYINPUT42), .A2(n1127), .ZN(n1126) );
XOR2_X1 U813 ( .A(n1128), .B(n1129), .Z(n1127) );
XNOR2_X1 U814 ( .A(n1130), .B(n1131), .ZN(n1129) );
NOR2_X1 U815 ( .A1(KEYINPUT39), .A2(n1132), .ZN(n1131) );
XNOR2_X1 U816 ( .A(G134), .B(n1133), .ZN(n1132) );
XNOR2_X1 U817 ( .A(n1134), .B(KEYINPUT56), .ZN(n1128) );
AND2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(n1113) );
XOR2_X1 U819 ( .A(n1137), .B(n1138), .Z(G69) );
NOR2_X1 U820 ( .A1(n1139), .A2(n1136), .ZN(n1138) );
AND2_X1 U821 ( .A1(G224), .A2(G898), .ZN(n1139) );
NAND2_X1 U822 ( .A1(n1140), .A2(n1141), .ZN(n1137) );
NAND3_X1 U823 ( .A1(n1142), .A2(n1136), .A3(n1143), .ZN(n1141) );
XOR2_X1 U824 ( .A(n1144), .B(KEYINPUT60), .Z(n1140) );
NAND3_X1 U825 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
INV_X1 U826 ( .A(n1143), .ZN(n1147) );
XNOR2_X1 U827 ( .A(n1148), .B(n1149), .ZN(n1143) );
XNOR2_X1 U828 ( .A(KEYINPUT2), .B(n1150), .ZN(n1149) );
XOR2_X1 U829 ( .A(n1151), .B(n1152), .Z(n1148) );
NAND2_X1 U830 ( .A1(G953), .A2(n1153), .ZN(n1146) );
NAND2_X1 U831 ( .A1(n1142), .A2(n1136), .ZN(n1145) );
NOR3_X1 U832 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(G66) );
NOR3_X1 U833 ( .A1(n1157), .A2(n1158), .A3(n1136), .ZN(n1156) );
INV_X1 U834 ( .A(KEYINPUT53), .ZN(n1157) );
NOR2_X1 U835 ( .A1(KEYINPUT53), .A2(n1159), .ZN(n1155) );
NOR2_X1 U836 ( .A1(n1160), .A2(n1161), .ZN(n1154) );
XOR2_X1 U837 ( .A(n1162), .B(KEYINPUT6), .Z(n1161) );
NAND2_X1 U838 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NAND2_X1 U839 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NOR3_X1 U840 ( .A1(n1167), .A2(n1163), .A3(n1168), .ZN(n1160) );
NOR2_X1 U841 ( .A1(n1169), .A2(n1170), .ZN(G63) );
XOR2_X1 U842 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1167), .ZN(n1171) );
INV_X1 U844 ( .A(G478), .ZN(n1173) );
NOR2_X1 U845 ( .A1(n1169), .A2(n1174), .ZN(G60) );
XOR2_X1 U846 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U847 ( .A1(n1177), .A2(n1167), .ZN(n1175) );
XOR2_X1 U848 ( .A(n1178), .B(n1179), .Z(G6) );
NAND2_X1 U849 ( .A1(KEYINPUT63), .A2(G104), .ZN(n1179) );
NOR2_X1 U850 ( .A1(n1169), .A2(n1180), .ZN(G57) );
XOR2_X1 U851 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U852 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U853 ( .A1(n1185), .A2(n1167), .ZN(n1183) );
NOR2_X1 U854 ( .A1(n1169), .A2(n1186), .ZN(G54) );
XOR2_X1 U855 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U856 ( .A(KEYINPUT3), .B(n1189), .Z(n1188) );
NOR2_X1 U857 ( .A1(n1190), .A2(n1167), .ZN(n1189) );
XOR2_X1 U858 ( .A(n1191), .B(n1192), .Z(n1187) );
NOR2_X1 U859 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
NOR2_X1 U860 ( .A1(G110), .A2(n1195), .ZN(n1194) );
XOR2_X1 U861 ( .A(KEYINPUT29), .B(n1196), .Z(n1195) );
NOR2_X1 U862 ( .A1(n1196), .A2(n1150), .ZN(n1193) );
NOR2_X1 U863 ( .A1(n1169), .A2(n1197), .ZN(G51) );
XOR2_X1 U864 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U865 ( .A(n1200), .B(n1201), .ZN(n1198) );
NOR2_X1 U866 ( .A1(n1202), .A2(n1167), .ZN(n1201) );
NAND2_X1 U867 ( .A1(G902), .A2(n1166), .ZN(n1167) );
INV_X1 U868 ( .A(n1070), .ZN(n1166) );
NOR2_X1 U869 ( .A1(n1142), .A2(n1135), .ZN(n1070) );
NAND4_X1 U870 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1135) );
NOR4_X1 U871 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
NOR4_X1 U872 ( .A1(n1211), .A2(n1063), .A3(n1212), .A4(n1213), .ZN(n1210) );
NOR2_X1 U873 ( .A1(KEYINPUT26), .A2(n1214), .ZN(n1213) );
NOR2_X1 U874 ( .A1(n1215), .A2(n1082), .ZN(n1214) );
INV_X1 U875 ( .A(n1216), .ZN(n1215) );
NOR2_X1 U876 ( .A1(n1217), .A2(n1218), .ZN(n1212) );
INV_X1 U877 ( .A(KEYINPUT26), .ZN(n1218) );
NAND2_X1 U878 ( .A1(n1090), .A2(n1219), .ZN(n1211) );
NOR3_X1 U879 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1209) );
XNOR2_X1 U880 ( .A(n1089), .B(KEYINPUT31), .ZN(n1221) );
INV_X1 U881 ( .A(n1223), .ZN(n1208) );
AND2_X1 U882 ( .A1(n1224), .A2(n1225), .ZN(n1205) );
NAND4_X1 U883 ( .A1(n1226), .A2(n1178), .A3(n1227), .A4(n1228), .ZN(n1142) );
AND4_X1 U884 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
NOR2_X1 U885 ( .A1(n1233), .A2(n1234), .ZN(n1227) );
NOR4_X1 U886 ( .A1(n1235), .A2(n1059), .A3(n1236), .A4(n1237), .ZN(n1234) );
XNOR2_X1 U887 ( .A(KEYINPUT21), .B(n1238), .ZN(n1237) );
NOR3_X1 U888 ( .A1(n1091), .A2(n1239), .A3(n1240), .ZN(n1233) );
NOR2_X1 U889 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
INV_X1 U890 ( .A(KEYINPUT33), .ZN(n1242) );
NOR2_X1 U891 ( .A1(n1089), .A2(n1243), .ZN(n1241) );
NOR2_X1 U892 ( .A1(KEYINPUT33), .A2(n1045), .ZN(n1239) );
NAND2_X1 U893 ( .A1(n1066), .A2(n1219), .ZN(n1091) );
NAND3_X1 U894 ( .A1(n1045), .A2(n1066), .A3(n1076), .ZN(n1178) );
INV_X1 U895 ( .A(n1159), .ZN(n1169) );
NAND2_X1 U896 ( .A1(n1158), .A2(G953), .ZN(n1159) );
XNOR2_X1 U897 ( .A(G952), .B(KEYINPUT52), .ZN(n1158) );
XNOR2_X1 U898 ( .A(G146), .B(n1244), .ZN(G48) );
NAND2_X1 U899 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XNOR2_X1 U900 ( .A(G143), .B(n1223), .ZN(G45) );
NAND4_X1 U901 ( .A1(n1217), .A2(n1090), .A3(n1247), .A4(n1089), .ZN(n1223) );
NOR2_X1 U902 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XNOR2_X1 U903 ( .A(G140), .B(n1204), .ZN(G42) );
NAND4_X1 U904 ( .A1(n1083), .A2(n1217), .A3(n1076), .A4(n1250), .ZN(n1204) );
XOR2_X1 U905 ( .A(n1225), .B(n1251), .Z(G39) );
NAND2_X1 U906 ( .A1(KEYINPUT45), .A2(G137), .ZN(n1251) );
NAND3_X1 U907 ( .A1(n1083), .A2(n1055), .A3(n1246), .ZN(n1225) );
NAND2_X1 U908 ( .A1(n1252), .A2(n1253), .ZN(G36) );
NAND4_X1 U909 ( .A1(KEYINPUT8), .A2(n1254), .A3(n1219), .A4(n1255), .ZN(n1253) );
XNOR2_X1 U910 ( .A(KEYINPUT1), .B(n1256), .ZN(n1255) );
NAND2_X1 U911 ( .A1(n1257), .A2(n1258), .ZN(n1252) );
NAND2_X1 U912 ( .A1(n1259), .A2(n1256), .ZN(n1258) );
NAND2_X1 U913 ( .A1(KEYINPUT1), .A2(n1260), .ZN(n1259) );
INV_X1 U914 ( .A(KEYINPUT8), .ZN(n1260) );
NAND2_X1 U915 ( .A1(n1254), .A2(n1219), .ZN(n1257) );
XNOR2_X1 U916 ( .A(G131), .B(n1224), .ZN(G33) );
NAND2_X1 U917 ( .A1(n1254), .A2(n1076), .ZN(n1224) );
AND3_X1 U918 ( .A1(n1217), .A2(n1090), .A3(n1083), .ZN(n1254) );
INV_X1 U919 ( .A(n1063), .ZN(n1083) );
NAND2_X1 U920 ( .A1(n1065), .A2(n1110), .ZN(n1063) );
NAND3_X1 U921 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(G30) );
NAND2_X1 U922 ( .A1(n1207), .A2(n1264), .ZN(n1263) );
INV_X1 U923 ( .A(n1265), .ZN(n1207) );
NAND2_X1 U924 ( .A1(n1266), .A2(n1267), .ZN(n1262) );
INV_X1 U925 ( .A(KEYINPUT57), .ZN(n1267) );
NAND2_X1 U926 ( .A1(G128), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U927 ( .A(KEYINPUT58), .B(n1265), .ZN(n1268) );
NAND2_X1 U928 ( .A1(KEYINPUT57), .A2(n1269), .ZN(n1261) );
NAND2_X1 U929 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND3_X1 U930 ( .A1(KEYINPUT58), .A2(G128), .A3(n1265), .ZN(n1271) );
OR2_X1 U931 ( .A1(n1265), .A2(KEYINPUT58), .ZN(n1270) );
NAND3_X1 U932 ( .A1(n1219), .A2(n1089), .A3(n1246), .ZN(n1265) );
INV_X1 U933 ( .A(n1220), .ZN(n1246) );
NAND3_X1 U934 ( .A1(n1272), .A2(n1273), .A3(n1217), .ZN(n1220) );
AND2_X1 U935 ( .A1(n1082), .A2(n1216), .ZN(n1217) );
XNOR2_X1 U936 ( .A(G101), .B(n1232), .ZN(G3) );
NAND3_X1 U937 ( .A1(n1055), .A2(n1045), .A3(n1090), .ZN(n1232) );
XNOR2_X1 U938 ( .A(G125), .B(n1203), .ZN(G27) );
NAND4_X1 U939 ( .A1(n1245), .A2(n1084), .A3(n1250), .A4(n1216), .ZN(n1203) );
NAND2_X1 U940 ( .A1(n1274), .A2(n1052), .ZN(n1216) );
XOR2_X1 U941 ( .A(KEYINPUT22), .B(n1275), .Z(n1274) );
NOR4_X1 U942 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1136), .ZN(n1275) );
XNOR2_X1 U943 ( .A(G900), .B(KEYINPUT15), .ZN(n1277) );
INV_X1 U944 ( .A(n1279), .ZN(n1276) );
NOR2_X1 U945 ( .A1(n1222), .A2(n1235), .ZN(n1245) );
INV_X1 U946 ( .A(n1076), .ZN(n1222) );
XOR2_X1 U947 ( .A(G122), .B(n1280), .Z(G24) );
NOR2_X1 U948 ( .A1(n1226), .A2(n1281), .ZN(n1280) );
XOR2_X1 U949 ( .A(KEYINPUT48), .B(KEYINPUT19), .Z(n1281) );
NAND4_X1 U950 ( .A1(n1282), .A2(n1066), .A3(n1283), .A4(n1284), .ZN(n1226) );
NOR2_X1 U951 ( .A1(n1285), .A2(n1273), .ZN(n1066) );
XNOR2_X1 U952 ( .A(G119), .B(n1286), .ZN(G21) );
NAND3_X1 U953 ( .A1(n1287), .A2(n1282), .A3(KEYINPUT14), .ZN(n1286) );
INV_X1 U954 ( .A(n1236), .ZN(n1287) );
NAND3_X1 U955 ( .A1(n1272), .A2(n1055), .A3(n1273), .ZN(n1236) );
INV_X1 U956 ( .A(n1288), .ZN(n1273) );
NAND2_X1 U957 ( .A1(n1289), .A2(n1290), .ZN(G18) );
NAND2_X1 U958 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U959 ( .A(KEYINPUT17), .B(n1293), .Z(n1289) );
NOR2_X1 U960 ( .A1(n1291), .A2(n1292), .ZN(n1293) );
INV_X1 U961 ( .A(n1231), .ZN(n1291) );
NAND3_X1 U962 ( .A1(n1282), .A2(n1219), .A3(n1090), .ZN(n1231) );
NOR2_X1 U963 ( .A1(n1283), .A2(n1248), .ZN(n1219) );
XNOR2_X1 U964 ( .A(G113), .B(n1230), .ZN(G15) );
NAND3_X1 U965 ( .A1(n1282), .A2(n1076), .A3(n1090), .ZN(n1230) );
NOR2_X1 U966 ( .A1(n1288), .A2(n1285), .ZN(n1090) );
NOR2_X1 U967 ( .A1(n1284), .A2(n1249), .ZN(n1076) );
AND3_X1 U968 ( .A1(n1089), .A2(n1238), .A3(n1084), .ZN(n1282) );
INV_X1 U969 ( .A(n1059), .ZN(n1084) );
NAND2_X1 U970 ( .A1(n1294), .A2(n1069), .ZN(n1059) );
XNOR2_X1 U971 ( .A(KEYINPUT5), .B(n1067), .ZN(n1294) );
XNOR2_X1 U972 ( .A(G110), .B(n1229), .ZN(G12) );
NAND3_X1 U973 ( .A1(n1055), .A2(n1045), .A3(n1250), .ZN(n1229) );
INV_X1 U974 ( .A(n1062), .ZN(n1250) );
NAND2_X1 U975 ( .A1(n1272), .A2(n1288), .ZN(n1062) );
XNOR2_X1 U976 ( .A(n1105), .B(KEYINPUT13), .ZN(n1288) );
XNOR2_X1 U977 ( .A(n1295), .B(n1185), .ZN(n1105) );
INV_X1 U978 ( .A(G472), .ZN(n1185) );
NAND2_X1 U979 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XNOR2_X1 U980 ( .A(n1184), .B(n1298), .ZN(n1297) );
XNOR2_X1 U981 ( .A(KEYINPUT62), .B(n1299), .ZN(n1298) );
NOR2_X1 U982 ( .A1(KEYINPUT9), .A2(n1181), .ZN(n1299) );
XNOR2_X1 U983 ( .A(n1300), .B(n1301), .ZN(n1181) );
NOR2_X1 U984 ( .A1(KEYINPUT51), .A2(G116), .ZN(n1301) );
XNOR2_X1 U985 ( .A(G113), .B(G119), .ZN(n1300) );
XNOR2_X1 U986 ( .A(n1302), .B(n1303), .ZN(n1184) );
XNOR2_X1 U987 ( .A(n1304), .B(n1305), .ZN(n1303) );
INV_X1 U988 ( .A(G101), .ZN(n1304) );
XOR2_X1 U989 ( .A(n1306), .B(n1307), .Z(n1302) );
AND3_X1 U990 ( .A1(G210), .A2(n1136), .A3(n1308), .ZN(n1307) );
XNOR2_X1 U991 ( .A(G902), .B(KEYINPUT46), .ZN(n1296) );
XOR2_X1 U992 ( .A(n1285), .B(KEYINPUT20), .Z(n1272) );
NAND2_X1 U993 ( .A1(n1109), .A2(n1102), .ZN(n1285) );
NAND3_X1 U994 ( .A1(n1168), .A2(n1278), .A3(n1163), .ZN(n1102) );
INV_X1 U995 ( .A(n1309), .ZN(n1163) );
INV_X1 U996 ( .A(n1165), .ZN(n1109) );
NOR2_X1 U997 ( .A1(n1168), .A2(n1100), .ZN(n1165) );
NOR2_X1 U998 ( .A1(G902), .A2(n1309), .ZN(n1100) );
XNOR2_X1 U999 ( .A(n1310), .B(n1311), .ZN(n1309) );
XOR2_X1 U1000 ( .A(n1312), .B(n1313), .Z(n1311) );
XNOR2_X1 U1001 ( .A(n1264), .B(G119), .ZN(n1313) );
INV_X1 U1002 ( .A(G128), .ZN(n1264) );
XNOR2_X1 U1003 ( .A(KEYINPUT43), .B(n1314), .ZN(n1312) );
XOR2_X1 U1004 ( .A(n1315), .B(n1316), .Z(n1310) );
XNOR2_X1 U1005 ( .A(n1317), .B(n1318), .ZN(n1316) );
XOR2_X1 U1006 ( .A(n1319), .B(n1320), .Z(n1315) );
AND3_X1 U1007 ( .A1(G221), .A2(n1136), .A3(G234), .ZN(n1320) );
NAND2_X1 U1008 ( .A1(KEYINPUT28), .A2(n1150), .ZN(n1319) );
NAND2_X1 U1009 ( .A1(G217), .A2(n1321), .ZN(n1168) );
NOR2_X1 U1010 ( .A1(n1235), .A2(n1243), .ZN(n1045) );
NAND2_X1 U1011 ( .A1(n1082), .A2(n1238), .ZN(n1243) );
NAND2_X1 U1012 ( .A1(n1052), .A2(n1322), .ZN(n1238) );
NAND4_X1 U1013 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1153), .ZN(n1322) );
INV_X1 U1014 ( .A(G898), .ZN(n1153) );
NAND3_X1 U1015 ( .A1(n1279), .A2(n1136), .A3(n1323), .ZN(n1052) );
XOR2_X1 U1016 ( .A(KEYINPUT18), .B(G952), .Z(n1323) );
NAND2_X1 U1017 ( .A1(G237), .A2(G234), .ZN(n1279) );
AND2_X1 U1018 ( .A1(n1067), .A2(n1069), .ZN(n1082) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1321), .ZN(n1069) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1278), .ZN(n1321) );
XNOR2_X1 U1021 ( .A(n1324), .B(n1103), .ZN(n1067) );
NAND2_X1 U1022 ( .A1(n1325), .A2(n1278), .ZN(n1103) );
XOR2_X1 U1023 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1024 ( .A(n1191), .B(n1196), .ZN(n1327) );
XOR2_X1 U1025 ( .A(G140), .B(n1328), .Z(n1196) );
AND2_X1 U1026 ( .A1(n1136), .A2(G227), .ZN(n1328) );
XOR2_X1 U1027 ( .A(n1329), .B(n1330), .Z(n1191) );
XNOR2_X1 U1028 ( .A(n1306), .B(n1331), .ZN(n1329) );
INV_X1 U1029 ( .A(n1134), .ZN(n1331) );
NOR2_X1 U1030 ( .A1(n1332), .A2(n1333), .ZN(n1134) );
INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n1332) );
XNOR2_X1 U1032 ( .A(n1334), .B(n1335), .ZN(n1306) );
XNOR2_X1 U1033 ( .A(n1336), .B(n1256), .ZN(n1334) );
INV_X1 U1034 ( .A(G134), .ZN(n1256) );
NAND2_X1 U1035 ( .A1(KEYINPUT16), .A2(n1318), .ZN(n1336) );
INV_X1 U1036 ( .A(n1133), .ZN(n1318) );
XOR2_X1 U1037 ( .A(G137), .B(KEYINPUT50), .Z(n1133) );
XNOR2_X1 U1038 ( .A(KEYINPUT49), .B(n1150), .ZN(n1326) );
INV_X1 U1039 ( .A(G110), .ZN(n1150) );
NAND2_X1 U1040 ( .A1(KEYINPUT41), .A2(n1190), .ZN(n1324) );
INV_X1 U1041 ( .A(G469), .ZN(n1190) );
INV_X1 U1042 ( .A(n1089), .ZN(n1235) );
NOR2_X1 U1043 ( .A1(n1065), .A2(n1064), .ZN(n1089) );
INV_X1 U1044 ( .A(n1110), .ZN(n1064) );
NAND2_X1 U1045 ( .A1(G214), .A2(n1337), .ZN(n1110) );
XNOR2_X1 U1046 ( .A(n1104), .B(KEYINPUT32), .ZN(n1065) );
XNOR2_X1 U1047 ( .A(n1338), .B(n1202), .ZN(n1104) );
NAND2_X1 U1048 ( .A1(G210), .A2(n1337), .ZN(n1202) );
NAND2_X1 U1049 ( .A1(n1308), .A2(n1278), .ZN(n1337) );
INV_X1 U1050 ( .A(G237), .ZN(n1308) );
NAND2_X1 U1051 ( .A1(n1339), .A2(n1278), .ZN(n1338) );
INV_X1 U1052 ( .A(G902), .ZN(n1278) );
XOR2_X1 U1053 ( .A(n1340), .B(n1341), .Z(n1339) );
XOR2_X1 U1054 ( .A(KEYINPUT30), .B(n1342), .Z(n1341) );
XOR2_X1 U1055 ( .A(KEYINPUT7), .B(KEYINPUT61), .Z(n1342) );
XNOR2_X1 U1056 ( .A(n1343), .B(n1344), .ZN(n1340) );
INV_X1 U1057 ( .A(n1200), .ZN(n1344) );
XNOR2_X1 U1058 ( .A(n1345), .B(n1346), .ZN(n1200) );
XOR2_X1 U1059 ( .A(n1347), .B(n1348), .Z(n1346) );
NAND2_X1 U1060 ( .A1(G224), .A2(n1136), .ZN(n1348) );
NAND2_X1 U1061 ( .A1(n1349), .A2(KEYINPUT37), .ZN(n1347) );
XNOR2_X1 U1062 ( .A(n1151), .B(n1292), .ZN(n1349) );
INV_X1 U1063 ( .A(G116), .ZN(n1292) );
XOR2_X1 U1064 ( .A(n1350), .B(n1330), .Z(n1151) );
XNOR2_X1 U1065 ( .A(n1351), .B(n1352), .ZN(n1330) );
XOR2_X1 U1066 ( .A(KEYINPUT23), .B(G107), .Z(n1352) );
XNOR2_X1 U1067 ( .A(G101), .B(G104), .ZN(n1351) );
XOR2_X1 U1068 ( .A(n1353), .B(G113), .Z(n1350) );
NAND2_X1 U1069 ( .A1(KEYINPUT34), .A2(G119), .ZN(n1353) );
XNOR2_X1 U1070 ( .A(G110), .B(n1354), .ZN(n1345) );
XNOR2_X1 U1071 ( .A(n1123), .B(G122), .ZN(n1354) );
NAND2_X1 U1072 ( .A1(KEYINPUT10), .A2(n1199), .ZN(n1343) );
XOR2_X1 U1073 ( .A(n1355), .B(n1305), .Z(n1199) );
NOR2_X1 U1074 ( .A1(KEYINPUT47), .A2(n1333), .ZN(n1305) );
XOR2_X1 U1075 ( .A(G128), .B(KEYINPUT40), .Z(n1333) );
NOR2_X1 U1076 ( .A1(n1284), .A2(n1283), .ZN(n1055) );
INV_X1 U1077 ( .A(n1249), .ZN(n1283) );
XOR2_X1 U1078 ( .A(n1108), .B(n1177), .Z(n1249) );
INV_X1 U1079 ( .A(G475), .ZN(n1177) );
NOR2_X1 U1080 ( .A1(n1176), .A2(G902), .ZN(n1108) );
XNOR2_X1 U1081 ( .A(n1356), .B(n1357), .ZN(n1176) );
XNOR2_X1 U1082 ( .A(n1317), .B(n1335), .ZN(n1357) );
INV_X1 U1083 ( .A(n1130), .ZN(n1335) );
XOR2_X1 U1084 ( .A(G131), .B(n1355), .Z(n1130) );
XNOR2_X1 U1085 ( .A(G143), .B(n1314), .ZN(n1355) );
INV_X1 U1086 ( .A(G146), .ZN(n1314) );
XNOR2_X1 U1087 ( .A(n1123), .B(G140), .ZN(n1317) );
INV_X1 U1088 ( .A(G125), .ZN(n1123) );
XOR2_X1 U1089 ( .A(n1358), .B(n1359), .Z(n1356) );
NOR2_X1 U1090 ( .A1(KEYINPUT36), .A2(n1360), .ZN(n1359) );
XOR2_X1 U1091 ( .A(G104), .B(n1361), .Z(n1360) );
NOR2_X1 U1092 ( .A1(KEYINPUT59), .A2(n1362), .ZN(n1361) );
XNOR2_X1 U1093 ( .A(G113), .B(G122), .ZN(n1362) );
NAND3_X1 U1094 ( .A1(G214), .A2(n1136), .A3(n1363), .ZN(n1358) );
XNOR2_X1 U1095 ( .A(G237), .B(KEYINPUT54), .ZN(n1363) );
INV_X1 U1096 ( .A(n1248), .ZN(n1284) );
NOR2_X1 U1097 ( .A1(n1112), .A2(n1364), .ZN(n1248) );
AND2_X1 U1098 ( .A1(G478), .A2(n1111), .ZN(n1364) );
NOR2_X1 U1099 ( .A1(n1111), .A2(G478), .ZN(n1112) );
OR2_X1 U1100 ( .A1(n1172), .A2(G902), .ZN(n1111) );
XNOR2_X1 U1101 ( .A(n1365), .B(n1366), .ZN(n1172) );
XOR2_X1 U1102 ( .A(G107), .B(n1367), .Z(n1366) );
XNOR2_X1 U1103 ( .A(n1368), .B(G128), .ZN(n1367) );
INV_X1 U1104 ( .A(G143), .ZN(n1368) );
XNOR2_X1 U1105 ( .A(n1152), .B(n1369), .ZN(n1365) );
XNOR2_X1 U1106 ( .A(n1370), .B(n1371), .ZN(n1369) );
NOR2_X1 U1107 ( .A1(KEYINPUT0), .A2(G134), .ZN(n1371) );
NAND4_X1 U1108 ( .A1(KEYINPUT27), .A2(G217), .A3(G234), .A4(n1136), .ZN(n1370) );
INV_X1 U1109 ( .A(G953), .ZN(n1136) );
XOR2_X1 U1110 ( .A(G116), .B(G122), .Z(n1152) );
endmodule


