//Key = 1011001110100110001010111001010010011110001000011000011100110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348;

XNOR2_X1 U739 ( .A(n1018), .B(n1019), .ZN(G9) );
NOR2_X1 U740 ( .A1(KEYINPUT21), .A2(n1020), .ZN(n1019) );
NOR2_X1 U741 ( .A1(n1021), .A2(n1022), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1023), .A2(n1024), .A3(KEYINPUT17), .A4(G953), .ZN(n1022) );
NAND3_X1 U743 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1023) );
NAND2_X1 U744 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NAND2_X1 U745 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND4_X1 U746 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND3_X1 U748 ( .A1(n1038), .A2(n1039), .A3(KEYINPUT23), .ZN(n1037) );
NAND2_X1 U749 ( .A1(n1040), .A2(n1041), .ZN(n1036) );
NAND2_X1 U750 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NAND2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U752 ( .A1(n1039), .A2(n1041), .A3(n1038), .ZN(n1030) );
NAND3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1041), .ZN(n1039) );
NAND2_X1 U754 ( .A1(n1034), .A2(n1048), .ZN(n1047) );
NAND2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1032), .A2(n1051), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U758 ( .A1(KEYINPUT22), .A2(n1054), .ZN(n1053) );
NAND2_X1 U759 ( .A1(n1033), .A2(n1055), .ZN(n1049) );
NAND2_X1 U760 ( .A1(KEYINPUT23), .A2(n1032), .ZN(n1055) );
OR4_X1 U761 ( .A1(n1056), .A2(KEYINPUT22), .A3(n1057), .A4(n1034), .ZN(n1046) );
INV_X1 U762 ( .A(n1058), .ZN(n1028) );
NAND4_X1 U763 ( .A1(n1032), .A2(n1038), .A3(n1033), .A4(n1059), .ZN(n1025) );
NOR3_X1 U764 ( .A1(n1058), .A2(n1060), .A3(n1061), .ZN(n1059) );
NOR2_X1 U765 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR3_X1 U767 ( .A1(n1024), .A2(G953), .A3(G952), .ZN(n1021) );
AND4_X1 U768 ( .A1(n1044), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1024) );
NOR4_X1 U769 ( .A1(n1069), .A2(n1060), .A3(n1070), .A4(n1071), .ZN(n1068) );
XOR2_X1 U770 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U771 ( .A1(n1074), .A2(KEYINPUT16), .ZN(n1073) );
XNOR2_X1 U772 ( .A(G469), .B(KEYINPUT25), .ZN(n1072) );
NOR2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1070) );
XOR2_X1 U774 ( .A(n1077), .B(KEYINPUT2), .Z(n1075) );
INV_X1 U775 ( .A(n1041), .ZN(n1060) );
NOR3_X1 U776 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1067) );
NOR2_X1 U777 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U778 ( .A(KEYINPUT55), .B(n1083), .Z(n1082) );
INV_X1 U779 ( .A(n1084), .ZN(n1081) );
NOR2_X1 U780 ( .A1(n1084), .A2(n1083), .ZN(n1079) );
XNOR2_X1 U781 ( .A(n1085), .B(KEYINPUT46), .ZN(n1083) );
INV_X1 U782 ( .A(n1034), .ZN(n1078) );
XOR2_X1 U783 ( .A(n1086), .B(n1087), .Z(G72) );
XOR2_X1 U784 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U785 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
AND2_X1 U786 ( .A1(G227), .A2(G900), .ZN(n1090) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NAND2_X1 U788 ( .A1(G953), .A2(n1094), .ZN(n1093) );
XOR2_X1 U789 ( .A(n1095), .B(n1096), .Z(n1092) );
XNOR2_X1 U790 ( .A(n1097), .B(n1098), .ZN(n1096) );
NOR2_X1 U791 ( .A1(KEYINPUT60), .A2(n1099), .ZN(n1098) );
NAND2_X1 U792 ( .A1(KEYINPUT6), .A2(n1100), .ZN(n1097) );
NAND2_X1 U793 ( .A1(n1091), .A2(n1101), .ZN(n1086) );
XOR2_X1 U794 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U795 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U796 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U797 ( .A1(G953), .A2(n1108), .ZN(n1107) );
XNOR2_X1 U798 ( .A(KEYINPUT47), .B(n1109), .ZN(n1108) );
NAND2_X1 U799 ( .A1(n1110), .A2(n1091), .ZN(n1104) );
NAND2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XNOR2_X1 U801 ( .A(KEYINPUT38), .B(n1113), .ZN(n1112) );
NOR2_X1 U802 ( .A1(n1114), .A2(n1091), .ZN(n1102) );
NOR2_X1 U803 ( .A1(n1115), .A2(n1109), .ZN(n1114) );
NOR2_X1 U804 ( .A1(n1116), .A2(n1117), .ZN(G66) );
XNOR2_X1 U805 ( .A(n1118), .B(n1119), .ZN(n1117) );
XOR2_X1 U806 ( .A(KEYINPUT4), .B(n1120), .Z(n1119) );
NOR2_X1 U807 ( .A1(n1084), .A2(n1121), .ZN(n1120) );
NOR3_X1 U808 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(G63) );
AND2_X1 U809 ( .A1(KEYINPUT3), .A2(n1116), .ZN(n1124) );
NOR3_X1 U810 ( .A1(KEYINPUT3), .A2(G953), .A3(G952), .ZN(n1123) );
NOR3_X1 U811 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1122) );
NOR2_X1 U812 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U813 ( .A1(KEYINPUT1), .A2(n1130), .ZN(n1128) );
XOR2_X1 U814 ( .A(n1131), .B(KEYINPUT9), .Z(n1130) );
NOR3_X1 U815 ( .A1(n1132), .A2(KEYINPUT1), .A3(n1131), .ZN(n1126) );
AND2_X1 U816 ( .A1(n1131), .A2(KEYINPUT1), .ZN(n1125) );
OR2_X1 U817 ( .A1(n1121), .A2(n1076), .ZN(n1131) );
NOR2_X1 U818 ( .A1(n1116), .A2(n1133), .ZN(G60) );
XOR2_X1 U819 ( .A(n1134), .B(n1135), .Z(n1133) );
NAND3_X1 U820 ( .A1(G475), .A2(n1136), .A3(n1137), .ZN(n1134) );
XNOR2_X1 U821 ( .A(G902), .B(KEYINPUT10), .ZN(n1137) );
XNOR2_X1 U822 ( .A(G104), .B(n1113), .ZN(G6) );
NOR2_X1 U823 ( .A1(n1116), .A2(n1138), .ZN(G57) );
XOR2_X1 U824 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U825 ( .A(n1141), .B(n1142), .Z(n1140) );
NAND2_X1 U826 ( .A1(KEYINPUT59), .A2(n1143), .ZN(n1142) );
NAND3_X1 U827 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1141) );
NAND2_X1 U828 ( .A1(KEYINPUT50), .A2(n1147), .ZN(n1146) );
NAND3_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1145) );
NAND2_X1 U830 ( .A1(n1151), .A2(n1152), .ZN(n1144) );
NAND2_X1 U831 ( .A1(n1153), .A2(n1149), .ZN(n1152) );
INV_X1 U832 ( .A(KEYINPUT50), .ZN(n1149) );
XNOR2_X1 U833 ( .A(n1147), .B(KEYINPUT31), .ZN(n1153) );
XOR2_X1 U834 ( .A(G101), .B(n1154), .Z(n1139) );
NOR2_X1 U835 ( .A1(n1155), .A2(n1121), .ZN(n1154) );
XNOR2_X1 U836 ( .A(G472), .B(KEYINPUT40), .ZN(n1155) );
NOR2_X1 U837 ( .A1(n1116), .A2(n1156), .ZN(G54) );
XOR2_X1 U838 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U839 ( .A(KEYINPUT36), .B(n1159), .Z(n1158) );
NOR2_X1 U840 ( .A1(n1160), .A2(n1121), .ZN(n1159) );
NAND2_X1 U841 ( .A1(G902), .A2(n1136), .ZN(n1121) );
NAND2_X1 U842 ( .A1(n1161), .A2(n1162), .ZN(n1157) );
NAND3_X1 U843 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(n1162) );
NAND2_X1 U844 ( .A1(n1166), .A2(n1167), .ZN(n1163) );
NAND2_X1 U845 ( .A1(KEYINPUT54), .A2(n1168), .ZN(n1167) );
INV_X1 U846 ( .A(n1169), .ZN(n1166) );
XOR2_X1 U847 ( .A(KEYINPUT7), .B(n1170), .Z(n1161) );
NOR3_X1 U848 ( .A1(n1165), .A2(n1169), .A3(n1171), .ZN(n1170) );
NOR2_X1 U849 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
INV_X1 U850 ( .A(KEYINPUT54), .ZN(n1173) );
NOR2_X1 U851 ( .A1(n1168), .A2(KEYINPUT54), .ZN(n1169) );
NOR2_X1 U852 ( .A1(n1116), .A2(n1174), .ZN(G51) );
XOR2_X1 U853 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U854 ( .A(n1177), .B(G125), .Z(n1175) );
NAND4_X1 U855 ( .A1(n1178), .A2(KEYINPUT24), .A3(G902), .A4(G210), .ZN(n1177) );
XNOR2_X1 U856 ( .A(n1027), .B(KEYINPUT5), .ZN(n1178) );
INV_X1 U857 ( .A(n1136), .ZN(n1027) );
NAND3_X1 U858 ( .A1(n1179), .A2(n1113), .A3(n1111), .ZN(n1136) );
AND4_X1 U859 ( .A1(n1180), .A2(n1181), .A3(n1020), .A4(n1182), .ZN(n1111) );
NOR3_X1 U860 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1182) );
INV_X1 U861 ( .A(n1186), .ZN(n1184) );
NOR2_X1 U862 ( .A1(n1187), .A2(n1042), .ZN(n1183) );
NOR2_X1 U863 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U864 ( .A1(n1057), .A2(n1190), .ZN(n1189) );
NOR3_X1 U865 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1188) );
XOR2_X1 U866 ( .A(n1194), .B(KEYINPUT53), .Z(n1192) );
NAND4_X1 U867 ( .A1(n1195), .A2(n1038), .A3(n1054), .A4(n1194), .ZN(n1020) );
NAND4_X1 U868 ( .A1(n1196), .A2(n1195), .A3(n1197), .A4(n1194), .ZN(n1113) );
INV_X1 U869 ( .A(n1101), .ZN(n1179) );
NAND4_X1 U870 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1101) );
NOR4_X1 U871 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
NOR3_X1 U872 ( .A1(n1206), .A2(n1052), .A3(n1042), .ZN(n1205) );
NOR2_X1 U873 ( .A1(n1207), .A2(n1208), .ZN(n1200) );
NOR2_X1 U874 ( .A1(n1091), .A2(G952), .ZN(n1116) );
XOR2_X1 U875 ( .A(G146), .B(n1208), .Z(G48) );
AND2_X1 U876 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XNOR2_X1 U877 ( .A(n1211), .B(n1207), .ZN(G45) );
AND4_X1 U878 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1207) );
NOR2_X1 U879 ( .A1(n1193), .A2(n1042), .ZN(n1215) );
INV_X1 U880 ( .A(n1216), .ZN(n1042) );
XOR2_X1 U881 ( .A(G140), .B(n1204), .Z(G42) );
AND3_X1 U882 ( .A1(n1196), .A2(n1045), .A3(n1217), .ZN(n1204) );
XNOR2_X1 U883 ( .A(G137), .B(n1198), .ZN(G39) );
NAND4_X1 U884 ( .A1(n1217), .A2(n1033), .A3(n1218), .A4(n1045), .ZN(n1198) );
XNOR2_X1 U885 ( .A(G134), .B(n1199), .ZN(G36) );
NAND3_X1 U886 ( .A1(n1216), .A2(n1054), .A3(n1217), .ZN(n1199) );
XNOR2_X1 U887 ( .A(G131), .B(n1219), .ZN(G33) );
NAND4_X1 U888 ( .A1(KEYINPUT13), .A2(n1217), .A3(n1216), .A4(n1210), .ZN(n1219) );
INV_X1 U889 ( .A(n1206), .ZN(n1217) );
NAND4_X1 U890 ( .A1(n1034), .A2(n1056), .A3(n1212), .A4(n1041), .ZN(n1206) );
NOR2_X1 U891 ( .A1(n1064), .A2(n1220), .ZN(n1034) );
INV_X1 U892 ( .A(n1065), .ZN(n1220) );
NAND2_X1 U893 ( .A1(n1221), .A2(n1222), .ZN(G30) );
NAND2_X1 U894 ( .A1(n1203), .A2(n1223), .ZN(n1222) );
INV_X1 U895 ( .A(n1224), .ZN(n1203) );
XOR2_X1 U896 ( .A(n1225), .B(KEYINPUT15), .Z(n1221) );
NAND2_X1 U897 ( .A1(G128), .A2(n1224), .ZN(n1225) );
NAND2_X1 U898 ( .A1(n1209), .A2(n1054), .ZN(n1224) );
INV_X1 U899 ( .A(n1057), .ZN(n1054) );
AND4_X1 U900 ( .A1(n1195), .A2(n1218), .A3(n1045), .A4(n1212), .ZN(n1209) );
NAND2_X1 U901 ( .A1(n1226), .A2(n1227), .ZN(G3) );
NAND2_X1 U902 ( .A1(G101), .A2(n1228), .ZN(n1227) );
XOR2_X1 U903 ( .A(n1229), .B(KEYINPUT52), .Z(n1226) );
OR2_X1 U904 ( .A1(n1228), .A2(G101), .ZN(n1229) );
NAND2_X1 U905 ( .A1(n1230), .A2(n1216), .ZN(n1228) );
XNOR2_X1 U906 ( .A(n1202), .B(n1231), .ZN(G27) );
XNOR2_X1 U907 ( .A(G125), .B(KEYINPUT34), .ZN(n1231) );
AND4_X1 U908 ( .A1(n1196), .A2(n1232), .A3(n1045), .A4(n1212), .ZN(n1202) );
NAND2_X1 U909 ( .A1(n1058), .A2(n1233), .ZN(n1212) );
NAND4_X1 U910 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1094), .ZN(n1233) );
INV_X1 U911 ( .A(G900), .ZN(n1094) );
NOR2_X1 U912 ( .A1(n1052), .A2(n1218), .ZN(n1196) );
XNOR2_X1 U913 ( .A(n1181), .B(n1235), .ZN(G24) );
NOR2_X1 U914 ( .A1(KEYINPUT11), .A2(n1236), .ZN(n1235) );
NAND4_X1 U915 ( .A1(n1237), .A2(n1038), .A3(n1214), .A4(n1213), .ZN(n1181) );
NOR2_X1 U916 ( .A1(n1045), .A2(n1218), .ZN(n1038) );
XNOR2_X1 U917 ( .A(n1238), .B(n1185), .ZN(G21) );
NOR4_X1 U918 ( .A1(n1191), .A2(n1190), .A3(n1044), .A4(n1197), .ZN(n1185) );
INV_X1 U919 ( .A(n1045), .ZN(n1197) );
XNOR2_X1 U920 ( .A(G116), .B(n1239), .ZN(G18) );
NAND4_X1 U921 ( .A1(KEYINPUT58), .A2(n1216), .A3(n1240), .A4(n1232), .ZN(n1239) );
NOR2_X1 U922 ( .A1(n1241), .A2(n1057), .ZN(n1240) );
NAND2_X1 U923 ( .A1(n1066), .A2(n1213), .ZN(n1057) );
INV_X1 U924 ( .A(n1242), .ZN(n1213) );
XOR2_X1 U925 ( .A(n1194), .B(KEYINPUT63), .Z(n1241) );
NAND2_X1 U926 ( .A1(n1243), .A2(n1244), .ZN(G15) );
OR2_X1 U927 ( .A1(n1180), .A2(G113), .ZN(n1244) );
XOR2_X1 U928 ( .A(n1245), .B(KEYINPUT45), .Z(n1243) );
NAND2_X1 U929 ( .A1(G113), .A2(n1180), .ZN(n1245) );
NAND3_X1 U930 ( .A1(n1210), .A2(n1237), .A3(n1216), .ZN(n1180) );
NOR2_X1 U931 ( .A1(n1045), .A2(n1044), .ZN(n1216) );
INV_X1 U932 ( .A(n1190), .ZN(n1237) );
NAND2_X1 U933 ( .A1(n1232), .A2(n1194), .ZN(n1190) );
AND3_X1 U934 ( .A1(n1062), .A2(n1041), .A3(n1032), .ZN(n1232) );
INV_X1 U935 ( .A(n1052), .ZN(n1210) );
NAND2_X1 U936 ( .A1(n1242), .A2(n1214), .ZN(n1052) );
XNOR2_X1 U937 ( .A(n1066), .B(KEYINPUT30), .ZN(n1214) );
XNOR2_X1 U938 ( .A(G110), .B(n1186), .ZN(G12) );
NAND3_X1 U939 ( .A1(n1044), .A2(n1045), .A3(n1230), .ZN(n1186) );
AND3_X1 U940 ( .A1(n1195), .A2(n1194), .A3(n1033), .ZN(n1230) );
INV_X1 U941 ( .A(n1191), .ZN(n1033) );
NAND2_X1 U942 ( .A1(n1242), .A2(n1066), .ZN(n1191) );
XOR2_X1 U943 ( .A(n1246), .B(G475), .Z(n1066) );
NAND2_X1 U944 ( .A1(n1135), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U945 ( .A(n1248), .B(n1249), .ZN(n1135) );
XOR2_X1 U946 ( .A(n1250), .B(n1251), .Z(n1249) );
XNOR2_X1 U947 ( .A(n1252), .B(n1253), .ZN(n1251) );
NOR3_X1 U948 ( .A1(n1254), .A2(G237), .A3(n1255), .ZN(n1253) );
INV_X1 U949 ( .A(G214), .ZN(n1255) );
XNOR2_X1 U950 ( .A(KEYINPUT61), .B(n1091), .ZN(n1254) );
XNOR2_X1 U951 ( .A(n1256), .B(G113), .ZN(n1250) );
INV_X1 U952 ( .A(G131), .ZN(n1256) );
XOR2_X1 U953 ( .A(n1257), .B(n1258), .Z(n1248) );
XOR2_X1 U954 ( .A(n1259), .B(n1099), .Z(n1257) );
NAND2_X1 U955 ( .A1(KEYINPUT0), .A2(n1236), .ZN(n1259) );
NOR2_X1 U956 ( .A1(n1260), .A2(n1069), .ZN(n1242) );
NOR2_X1 U957 ( .A1(n1077), .A2(G478), .ZN(n1069) );
AND2_X1 U958 ( .A1(n1261), .A2(n1077), .ZN(n1260) );
NAND2_X1 U959 ( .A1(n1132), .A2(n1247), .ZN(n1077) );
INV_X1 U960 ( .A(n1129), .ZN(n1132) );
XNOR2_X1 U961 ( .A(n1262), .B(n1263), .ZN(n1129) );
XOR2_X1 U962 ( .A(G134), .B(n1264), .Z(n1263) );
NOR2_X1 U963 ( .A1(KEYINPUT57), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U964 ( .A(G143), .B(G128), .ZN(n1265) );
XOR2_X1 U965 ( .A(n1266), .B(n1267), .Z(n1262) );
NOR2_X1 U966 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
INV_X1 U967 ( .A(G217), .ZN(n1269) );
NAND2_X1 U968 ( .A1(n1270), .A2(n1271), .ZN(n1266) );
NAND2_X1 U969 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NAND2_X1 U970 ( .A1(KEYINPUT32), .A2(n1274), .ZN(n1273) );
NAND2_X1 U971 ( .A1(n1018), .A2(n1275), .ZN(n1274) );
INV_X1 U972 ( .A(n1276), .ZN(n1272) );
NAND2_X1 U973 ( .A1(G107), .A2(n1277), .ZN(n1270) );
NAND2_X1 U974 ( .A1(n1275), .A2(n1278), .ZN(n1277) );
NAND2_X1 U975 ( .A1(KEYINPUT32), .A2(n1276), .ZN(n1278) );
XOR2_X1 U976 ( .A(G116), .B(n1279), .Z(n1276) );
XNOR2_X1 U977 ( .A(KEYINPUT20), .B(n1236), .ZN(n1279) );
INV_X1 U978 ( .A(G122), .ZN(n1236) );
INV_X1 U979 ( .A(KEYINPUT62), .ZN(n1275) );
XNOR2_X1 U980 ( .A(KEYINPUT56), .B(n1076), .ZN(n1261) );
INV_X1 U981 ( .A(G478), .ZN(n1076) );
NAND2_X1 U982 ( .A1(n1280), .A2(n1281), .ZN(n1194) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1234), .A4(n1109), .ZN(n1281) );
INV_X1 U984 ( .A(G898), .ZN(n1109) );
XNOR2_X1 U985 ( .A(KEYINPUT27), .B(n1058), .ZN(n1280) );
NAND3_X1 U986 ( .A1(n1234), .A2(n1091), .A3(n1282), .ZN(n1058) );
XOR2_X1 U987 ( .A(KEYINPUT26), .B(G952), .Z(n1282) );
NAND2_X1 U988 ( .A1(G237), .A2(G234), .ZN(n1234) );
INV_X1 U989 ( .A(n1193), .ZN(n1195) );
NAND3_X1 U990 ( .A1(n1056), .A2(n1041), .A3(n1062), .ZN(n1193) );
AND2_X1 U991 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NAND2_X1 U992 ( .A1(G214), .A2(n1283), .ZN(n1065) );
NAND2_X1 U993 ( .A1(n1284), .A2(n1247), .ZN(n1283) );
NAND2_X1 U994 ( .A1(n1285), .A2(n1286), .ZN(n1064) );
NAND2_X1 U995 ( .A1(G210), .A2(n1287), .ZN(n1286) );
NAND2_X1 U996 ( .A1(n1247), .A2(n1288), .ZN(n1287) );
OR2_X1 U997 ( .A1(n1284), .A2(n1289), .ZN(n1288) );
NAND3_X1 U998 ( .A1(n1290), .A2(n1247), .A3(n1289), .ZN(n1285) );
XNOR2_X1 U999 ( .A(n1176), .B(n1291), .ZN(n1289) );
NOR2_X1 U1000 ( .A1(G125), .A2(KEYINPUT39), .ZN(n1291) );
XOR2_X1 U1001 ( .A(n1292), .B(n1106), .Z(n1176) );
XOR2_X1 U1002 ( .A(n1293), .B(n1294), .Z(n1106) );
XOR2_X1 U1003 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U1004 ( .A(n1297), .B(n1252), .ZN(n1296) );
NAND2_X1 U1005 ( .A1(KEYINPUT42), .A2(n1238), .ZN(n1297) );
INV_X1 U1006 ( .A(G119), .ZN(n1238) );
XNOR2_X1 U1007 ( .A(G110), .B(G122), .ZN(n1295) );
XOR2_X1 U1008 ( .A(n1298), .B(n1299), .Z(n1293) );
XOR2_X1 U1009 ( .A(n1300), .B(n1301), .Z(n1298) );
NAND2_X1 U1010 ( .A1(KEYINPUT8), .A2(n1018), .ZN(n1300) );
XOR2_X1 U1011 ( .A(n1302), .B(n1303), .Z(n1292) );
NOR2_X1 U1012 ( .A1(G953), .A2(n1115), .ZN(n1303) );
INV_X1 U1013 ( .A(G224), .ZN(n1115) );
NAND2_X1 U1014 ( .A1(G210), .A2(G237), .ZN(n1290) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1304), .ZN(n1041) );
INV_X1 U1016 ( .A(n1032), .ZN(n1056) );
XOR2_X1 U1017 ( .A(n1074), .B(n1160), .Z(n1032) );
INV_X1 U1018 ( .A(G469), .ZN(n1160) );
AND2_X1 U1019 ( .A1(n1305), .A2(n1247), .ZN(n1074) );
NAND2_X1 U1020 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND3_X1 U1021 ( .A1(KEYINPUT37), .A2(n1172), .A3(n1308), .ZN(n1307) );
XNOR2_X1 U1022 ( .A(n1309), .B(KEYINPUT18), .ZN(n1308) );
NAND3_X1 U1023 ( .A1(n1310), .A2(n1311), .A3(n1312), .ZN(n1306) );
XNOR2_X1 U1024 ( .A(KEYINPUT18), .B(n1165), .ZN(n1312) );
INV_X1 U1025 ( .A(n1309), .ZN(n1165) );
XNOR2_X1 U1026 ( .A(n1313), .B(n1314), .ZN(n1309) );
XOR2_X1 U1027 ( .A(n1315), .B(n1299), .Z(n1314) );
XOR2_X1 U1028 ( .A(G101), .B(KEYINPUT51), .Z(n1299) );
XOR2_X1 U1029 ( .A(n1100), .B(n1316), .Z(n1313) );
NOR2_X1 U1030 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
XOR2_X1 U1031 ( .A(KEYINPUT43), .B(n1319), .Z(n1318) );
NOR2_X1 U1032 ( .A1(n1018), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1033 ( .A(KEYINPUT33), .B(n1252), .ZN(n1320) );
INV_X1 U1034 ( .A(G107), .ZN(n1018) );
NOR2_X1 U1035 ( .A1(G107), .A2(n1252), .ZN(n1317) );
INV_X1 U1036 ( .A(G104), .ZN(n1252) );
NAND2_X1 U1037 ( .A1(n1321), .A2(n1322), .ZN(n1100) );
NAND2_X1 U1038 ( .A1(n1323), .A2(n1223), .ZN(n1322) );
XOR2_X1 U1039 ( .A(KEYINPUT14), .B(n1324), .Z(n1321) );
NOR2_X1 U1040 ( .A1(n1223), .A2(n1323), .ZN(n1324) );
XNOR2_X1 U1041 ( .A(n1211), .B(n1325), .ZN(n1323) );
NOR2_X1 U1042 ( .A1(KEYINPUT12), .A2(n1326), .ZN(n1325) );
INV_X1 U1043 ( .A(G143), .ZN(n1211) );
NAND3_X1 U1044 ( .A1(KEYINPUT37), .A2(n1172), .A3(n1327), .ZN(n1311) );
OR2_X1 U1045 ( .A1(n1327), .A2(n1172), .ZN(n1310) );
NAND2_X1 U1046 ( .A1(n1168), .A2(n1164), .ZN(n1172) );
NAND3_X1 U1047 ( .A1(G227), .A2(n1091), .A3(n1328), .ZN(n1164) );
XNOR2_X1 U1048 ( .A(G110), .B(G140), .ZN(n1328) );
NAND2_X1 U1049 ( .A1(n1329), .A2(n1330), .ZN(n1168) );
NAND2_X1 U1050 ( .A1(G227), .A2(n1091), .ZN(n1330) );
XNOR2_X1 U1051 ( .A(G140), .B(n1331), .ZN(n1329) );
INV_X1 U1052 ( .A(KEYINPUT44), .ZN(n1327) );
XOR2_X1 U1053 ( .A(n1085), .B(n1084), .Z(n1045) );
NAND2_X1 U1054 ( .A1(G217), .A2(n1304), .ZN(n1084) );
NAND2_X1 U1055 ( .A1(G234), .A2(n1247), .ZN(n1304) );
NAND2_X1 U1056 ( .A1(n1118), .A2(n1247), .ZN(n1085) );
XNOR2_X1 U1057 ( .A(n1332), .B(n1333), .ZN(n1118) );
XOR2_X1 U1058 ( .A(n1334), .B(n1335), .Z(n1333) );
XNOR2_X1 U1059 ( .A(n1331), .B(n1336), .ZN(n1335) );
NOR2_X1 U1060 ( .A1(KEYINPUT49), .A2(n1337), .ZN(n1336) );
XNOR2_X1 U1061 ( .A(n1099), .B(n1326), .ZN(n1337) );
XOR2_X1 U1062 ( .A(G125), .B(G140), .Z(n1099) );
INV_X1 U1063 ( .A(G110), .ZN(n1331) );
NOR2_X1 U1064 ( .A1(n1338), .A2(n1268), .ZN(n1334) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1091), .ZN(n1268) );
INV_X1 U1066 ( .A(G221), .ZN(n1338) );
XNOR2_X1 U1067 ( .A(G119), .B(n1339), .ZN(n1332) );
XNOR2_X1 U1068 ( .A(G137), .B(n1223), .ZN(n1339) );
INV_X1 U1069 ( .A(G128), .ZN(n1223) );
INV_X1 U1070 ( .A(n1218), .ZN(n1044) );
XNOR2_X1 U1071 ( .A(n1340), .B(G472), .ZN(n1218) );
NAND2_X1 U1072 ( .A1(n1341), .A2(n1247), .ZN(n1340) );
INV_X1 U1073 ( .A(G902), .ZN(n1247) );
XOR2_X1 U1074 ( .A(n1342), .B(n1343), .Z(n1341) );
XNOR2_X1 U1075 ( .A(G101), .B(n1344), .ZN(n1343) );
XNOR2_X1 U1076 ( .A(KEYINPUT48), .B(KEYINPUT41), .ZN(n1344) );
XNOR2_X1 U1077 ( .A(n1345), .B(n1148), .ZN(n1342) );
INV_X1 U1078 ( .A(n1147), .ZN(n1148) );
XOR2_X1 U1079 ( .A(G119), .B(n1301), .Z(n1147) );
XOR2_X1 U1080 ( .A(G116), .B(G113), .Z(n1301) );
XNOR2_X1 U1081 ( .A(n1150), .B(n1143), .ZN(n1345) );
NAND3_X1 U1082 ( .A1(n1284), .A2(n1091), .A3(G210), .ZN(n1143) );
INV_X1 U1083 ( .A(G953), .ZN(n1091) );
INV_X1 U1084 ( .A(G237), .ZN(n1284) );
INV_X1 U1085 ( .A(n1151), .ZN(n1150) );
XNOR2_X1 U1086 ( .A(n1302), .B(n1315), .ZN(n1151) );
XNOR2_X1 U1087 ( .A(n1095), .B(KEYINPUT28), .ZN(n1315) );
XNOR2_X1 U1088 ( .A(G131), .B(n1346), .ZN(n1095) );
XOR2_X1 U1089 ( .A(G137), .B(G134), .Z(n1346) );
XOR2_X1 U1090 ( .A(n1347), .B(n1348), .Z(n1302) );
XOR2_X1 U1091 ( .A(KEYINPUT29), .B(KEYINPUT19), .Z(n1348) );
XNOR2_X1 U1092 ( .A(n1258), .B(G128), .ZN(n1347) );
XNOR2_X1 U1093 ( .A(G143), .B(n1326), .ZN(n1258) );
XNOR2_X1 U1094 ( .A(G146), .B(KEYINPUT35), .ZN(n1326) );
endmodule


