//Key = 0011010101010101001111101011110111101000000101101011101001001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327;

XOR2_X1 U730 ( .A(n1002), .B(n1003), .Z(G9) );
NAND2_X1 U731 ( .A1(KEYINPUT22), .A2(G107), .ZN(n1003) );
NOR2_X1 U732 ( .A1(n1004), .A2(n1005), .ZN(G75) );
NOR3_X1 U733 ( .A1(n1006), .A2(G953), .A3(n1007), .ZN(n1005) );
INV_X1 U734 ( .A(n1008), .ZN(n1007) );
XNOR2_X1 U735 ( .A(G952), .B(KEYINPUT15), .ZN(n1006) );
NOR4_X1 U736 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1004) );
NOR3_X1 U737 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR4_X1 U738 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1014) );
INV_X1 U739 ( .A(KEYINPUT6), .ZN(n1013) );
NOR3_X1 U740 ( .A1(n1019), .A2(n1020), .A3(n1018), .ZN(n1011) );
NOR2_X1 U741 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U742 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U743 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U744 ( .A1(n1027), .A2(n1017), .ZN(n1026) );
NOR2_X1 U745 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR3_X1 U746 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1028) );
NOR2_X1 U747 ( .A1(n1016), .A2(n1033), .ZN(n1025) );
XNOR2_X1 U748 ( .A(n1034), .B(n1035), .ZN(n1033) );
NOR3_X1 U749 ( .A1(n1017), .A2(n1036), .A3(n1016), .ZN(n1021) );
NOR2_X1 U750 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
XOR2_X1 U751 ( .A(KEYINPUT42), .B(n1039), .Z(n1038) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U753 ( .A1(KEYINPUT6), .A2(n1015), .ZN(n1037) );
NAND3_X1 U754 ( .A1(n1042), .A2(n1043), .A3(n1008), .ZN(n1010) );
NAND4_X1 U755 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1008) );
NOR4_X1 U756 ( .A1(n1048), .A2(n1049), .A3(n1032), .A4(n1050), .ZN(n1047) );
XOR2_X1 U757 ( .A(n1051), .B(KEYINPUT52), .Z(n1050) );
INV_X1 U758 ( .A(n1052), .ZN(n1049) );
XOR2_X1 U759 ( .A(n1053), .B(n1054), .Z(n1045) );
NAND2_X1 U760 ( .A1(KEYINPUT57), .A2(n1055), .ZN(n1054) );
XOR2_X1 U761 ( .A(KEYINPUT34), .B(n1056), .Z(n1055) );
NAND3_X1 U762 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1042) );
OR2_X1 U763 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND4_X1 U764 ( .A1(n1062), .A2(n1063), .A3(G952), .A4(n1064), .ZN(n1009) );
NAND2_X1 U765 ( .A1(n1030), .A2(n1065), .ZN(n1064) );
NAND2_X1 U766 ( .A1(n1059), .A2(n1066), .ZN(n1065) );
NOR3_X1 U767 ( .A1(n1017), .A2(n1024), .A3(n1019), .ZN(n1059) );
INV_X1 U768 ( .A(KEYINPUT32), .ZN(n1030) );
XOR2_X1 U769 ( .A(n1067), .B(n1068), .Z(G72) );
XOR2_X1 U770 ( .A(n1069), .B(n1070), .Z(n1068) );
NAND2_X1 U771 ( .A1(G953), .A2(n1071), .ZN(n1070) );
NAND2_X1 U772 ( .A1(G900), .A2(G227), .ZN(n1071) );
NAND2_X1 U773 ( .A1(n1072), .A2(n1073), .ZN(n1069) );
OR2_X1 U774 ( .A1(n1043), .A2(G900), .ZN(n1073) );
XOR2_X1 U775 ( .A(n1074), .B(n1075), .Z(n1072) );
XOR2_X1 U776 ( .A(n1076), .B(n1077), .Z(n1075) );
XNOR2_X1 U777 ( .A(G131), .B(n1078), .ZN(n1077) );
XOR2_X1 U778 ( .A(n1079), .B(n1080), .Z(n1074) );
XNOR2_X1 U779 ( .A(n1081), .B(G134), .ZN(n1080) );
INV_X1 U780 ( .A(G137), .ZN(n1081) );
XNOR2_X1 U781 ( .A(KEYINPUT20), .B(n1082), .ZN(n1079) );
NOR2_X1 U782 ( .A1(n1062), .A2(G953), .ZN(n1067) );
XOR2_X1 U783 ( .A(n1083), .B(n1084), .Z(G69) );
NOR2_X1 U784 ( .A1(n1085), .A2(n1043), .ZN(n1084) );
NOR2_X1 U785 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U786 ( .A1(KEYINPUT10), .A2(n1088), .ZN(n1083) );
XOR2_X1 U787 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U788 ( .A1(G953), .A2(n1063), .ZN(n1090) );
NAND2_X1 U789 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NAND2_X1 U790 ( .A1(G953), .A2(n1087), .ZN(n1092) );
NOR2_X1 U791 ( .A1(n1093), .A2(n1094), .ZN(G66) );
XOR2_X1 U792 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U793 ( .A1(n1053), .A2(n1097), .ZN(n1095) );
NOR2_X1 U794 ( .A1(n1093), .A2(n1098), .ZN(G63) );
NOR2_X1 U795 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XOR2_X1 U796 ( .A(n1101), .B(KEYINPUT45), .Z(n1100) );
NAND2_X1 U797 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U798 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
NOR2_X1 U799 ( .A1(n1097), .A2(n1104), .ZN(n1102) );
INV_X1 U800 ( .A(G478), .ZN(n1104) );
NOR2_X1 U801 ( .A1(n1093), .A2(n1105), .ZN(G60) );
XOR2_X1 U802 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U803 ( .A1(n1108), .A2(n1097), .ZN(n1106) );
XOR2_X1 U804 ( .A(n1109), .B(n1110), .Z(G6) );
XNOR2_X1 U805 ( .A(G104), .B(KEYINPUT55), .ZN(n1110) );
NAND3_X1 U806 ( .A1(n1111), .A2(n1057), .A3(n1060), .ZN(n1109) );
NOR2_X1 U807 ( .A1(n1093), .A2(n1112), .ZN(G57) );
XOR2_X1 U808 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U809 ( .A1(n1115), .A2(KEYINPUT33), .ZN(n1114) );
XOR2_X1 U810 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR3_X1 U811 ( .A1(n1097), .A2(KEYINPUT0), .A3(n1118), .ZN(n1116) );
NAND3_X1 U812 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1113) );
OR2_X1 U813 ( .A1(n1122), .A2(KEYINPUT11), .ZN(n1121) );
NAND3_X1 U814 ( .A1(KEYINPUT11), .A2(n1122), .A3(G101), .ZN(n1120) );
NAND2_X1 U815 ( .A1(n1123), .A2(n1124), .ZN(n1119) );
INV_X1 U816 ( .A(G101), .ZN(n1124) );
NAND2_X1 U817 ( .A1(KEYINPUT11), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U818 ( .A(KEYINPUT19), .B(n1122), .ZN(n1125) );
XOR2_X1 U819 ( .A(n1126), .B(KEYINPUT36), .Z(n1122) );
NOR2_X1 U820 ( .A1(n1093), .A2(n1127), .ZN(G54) );
XOR2_X1 U821 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U822 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U823 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U824 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U825 ( .A(n1136), .B(KEYINPUT37), .Z(n1132) );
OR2_X1 U826 ( .A1(n1134), .A2(n1135), .ZN(n1136) );
XNOR2_X1 U827 ( .A(n1137), .B(n1076), .ZN(n1134) );
NAND2_X1 U828 ( .A1(KEYINPUT51), .A2(n1138), .ZN(n1137) );
NAND2_X1 U829 ( .A1(n1139), .A2(n1140), .ZN(n1130) );
XOR2_X1 U830 ( .A(n1141), .B(KEYINPUT16), .Z(n1139) );
NOR2_X1 U831 ( .A1(n1142), .A2(n1097), .ZN(n1128) );
NOR2_X1 U832 ( .A1(n1093), .A2(n1143), .ZN(G51) );
XOR2_X1 U833 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR3_X1 U834 ( .A1(n1097), .A2(KEYINPUT8), .A3(n1146), .ZN(n1145) );
INV_X1 U835 ( .A(G210), .ZN(n1146) );
NAND2_X1 U836 ( .A1(G902), .A2(n1147), .ZN(n1097) );
NAND2_X1 U837 ( .A1(n1062), .A2(n1063), .ZN(n1147) );
AND2_X1 U838 ( .A1(n1148), .A2(n1149), .ZN(n1063) );
NOR4_X1 U839 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1149) );
NOR3_X1 U840 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
XNOR2_X1 U841 ( .A(KEYINPUT7), .B(n1016), .ZN(n1154) );
INV_X1 U842 ( .A(n1057), .ZN(n1016) );
INV_X1 U843 ( .A(n1157), .ZN(n1152) );
AND4_X1 U844 ( .A1(n1002), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1148) );
NAND3_X1 U845 ( .A1(n1057), .A2(n1061), .A3(n1111), .ZN(n1002) );
AND4_X1 U846 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1062) );
NOR4_X1 U847 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1164) );
INV_X1 U848 ( .A(n1169), .ZN(n1166) );
NOR2_X1 U849 ( .A1(n1170), .A2(n1171), .ZN(n1163) );
NOR2_X1 U850 ( .A1(n1043), .A2(G952), .ZN(n1093) );
XOR2_X1 U851 ( .A(G146), .B(n1168), .Z(G48) );
AND3_X1 U852 ( .A1(n1032), .A2(n1172), .A3(n1173), .ZN(n1168) );
XNOR2_X1 U853 ( .A(n1174), .B(n1162), .ZN(G45) );
NAND3_X1 U854 ( .A1(n1029), .A2(n1172), .A3(n1175), .ZN(n1162) );
NOR3_X1 U855 ( .A1(n1015), .A2(n1176), .A3(n1177), .ZN(n1175) );
NAND2_X1 U856 ( .A1(KEYINPUT9), .A2(n1178), .ZN(n1174) );
XNOR2_X1 U857 ( .A(n1082), .B(n1167), .ZN(G42) );
AND3_X1 U858 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1167) );
XNOR2_X1 U859 ( .A(G137), .B(n1169), .ZN(G39) );
NAND3_X1 U860 ( .A1(n1046), .A2(n1182), .A3(n1183), .ZN(n1169) );
NOR3_X1 U861 ( .A1(n1184), .A2(n1031), .A3(n1179), .ZN(n1183) );
XNOR2_X1 U862 ( .A(G134), .B(n1185), .ZN(G36) );
NOR2_X1 U863 ( .A1(n1171), .A2(KEYINPUT35), .ZN(n1185) );
AND3_X1 U864 ( .A1(n1182), .A2(n1172), .A3(n1186), .ZN(n1171) );
XOR2_X1 U865 ( .A(G131), .B(n1165), .Z(G33) );
AND2_X1 U866 ( .A1(n1181), .A2(n1029), .ZN(n1165) );
NOR3_X1 U867 ( .A1(n1024), .A2(n1184), .A3(n1156), .ZN(n1181) );
INV_X1 U868 ( .A(n1182), .ZN(n1024) );
NOR2_X1 U869 ( .A1(n1040), .A2(n1048), .ZN(n1182) );
INV_X1 U870 ( .A(n1041), .ZN(n1048) );
XNOR2_X1 U871 ( .A(n1170), .B(n1187), .ZN(G30) );
NAND2_X1 U872 ( .A1(KEYINPUT3), .A2(G128), .ZN(n1187) );
AND4_X1 U873 ( .A1(n1032), .A2(n1172), .A3(n1188), .A4(n1061), .ZN(n1170) );
NOR2_X1 U874 ( .A1(n1031), .A2(n1015), .ZN(n1188) );
INV_X1 U875 ( .A(n1184), .ZN(n1172) );
NAND3_X1 U876 ( .A1(n1189), .A2(n1034), .A3(n1190), .ZN(n1184) );
XNOR2_X1 U877 ( .A(G101), .B(n1160), .ZN(G3) );
NAND3_X1 U878 ( .A1(n1029), .A2(n1111), .A3(n1046), .ZN(n1160) );
XNOR2_X1 U879 ( .A(n1078), .B(n1191), .ZN(G27) );
NOR2_X1 U880 ( .A1(n1161), .A2(n1192), .ZN(n1191) );
XOR2_X1 U881 ( .A(KEYINPUT26), .B(KEYINPUT13), .Z(n1192) );
NAND4_X1 U882 ( .A1(n1044), .A2(n1173), .A3(n1179), .A4(n1189), .ZN(n1161) );
NAND2_X1 U883 ( .A1(n1193), .A2(n1019), .ZN(n1189) );
NAND2_X1 U884 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
XOR2_X1 U885 ( .A(KEYINPUT48), .B(G900), .Z(n1195) );
NOR3_X1 U886 ( .A1(n1015), .A2(n1031), .A3(n1156), .ZN(n1173) );
INV_X1 U887 ( .A(n1060), .ZN(n1156) );
XNOR2_X1 U888 ( .A(G122), .B(n1159), .ZN(G24) );
NAND4_X1 U889 ( .A1(n1196), .A2(n1057), .A3(n1197), .A4(n1198), .ZN(n1159) );
NOR2_X1 U890 ( .A1(n1180), .A2(n1032), .ZN(n1057) );
XOR2_X1 U891 ( .A(n1151), .B(n1199), .Z(G21) );
NOR2_X1 U892 ( .A1(KEYINPUT47), .A2(n1200), .ZN(n1199) );
INV_X1 U893 ( .A(G119), .ZN(n1200) );
AND4_X1 U894 ( .A1(n1196), .A2(n1046), .A3(n1032), .A4(n1180), .ZN(n1151) );
XOR2_X1 U895 ( .A(n1201), .B(n1202), .Z(G18) );
NOR2_X1 U896 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
NOR2_X1 U897 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND4_X1 U898 ( .A1(n1044), .A2(n1186), .A3(n1015), .A4(n1207), .ZN(n1206) );
INV_X1 U899 ( .A(KEYINPUT4), .ZN(n1205) );
NOR2_X1 U900 ( .A1(KEYINPUT4), .A2(n1157), .ZN(n1203) );
NAND2_X1 U901 ( .A1(n1196), .A2(n1186), .ZN(n1157) );
AND2_X1 U902 ( .A1(n1029), .A2(n1061), .ZN(n1186) );
NOR2_X1 U903 ( .A1(n1197), .A2(n1176), .ZN(n1061) );
XNOR2_X1 U904 ( .A(G116), .B(KEYINPUT44), .ZN(n1201) );
XOR2_X1 U905 ( .A(G113), .B(n1208), .Z(G15) );
NOR2_X1 U906 ( .A1(KEYINPUT58), .A2(n1158), .ZN(n1208) );
NAND3_X1 U907 ( .A1(n1060), .A2(n1029), .A3(n1196), .ZN(n1158) );
AND3_X1 U908 ( .A1(n1209), .A2(n1207), .A3(n1044), .ZN(n1196) );
INV_X1 U909 ( .A(n1017), .ZN(n1044) );
NAND2_X1 U910 ( .A1(n1035), .A2(n1034), .ZN(n1017) );
NOR2_X1 U911 ( .A1(n1179), .A2(n1180), .ZN(n1029) );
NOR2_X1 U912 ( .A1(n1198), .A2(n1177), .ZN(n1060) );
INV_X1 U913 ( .A(n1197), .ZN(n1177) );
XOR2_X1 U914 ( .A(G110), .B(n1150), .Z(G12) );
AND2_X1 U915 ( .A1(n1066), .A2(n1111), .ZN(n1150) );
INV_X1 U916 ( .A(n1155), .ZN(n1111) );
NAND4_X1 U917 ( .A1(n1190), .A2(n1209), .A3(n1034), .A4(n1207), .ZN(n1155) );
NAND2_X1 U918 ( .A1(n1210), .A2(n1019), .ZN(n1207) );
NAND3_X1 U919 ( .A1(n1211), .A2(n1043), .A3(G952), .ZN(n1019) );
NAND2_X1 U920 ( .A1(n1194), .A2(n1087), .ZN(n1210) );
INV_X1 U921 ( .A(G898), .ZN(n1087) );
AND3_X1 U922 ( .A1(G953), .A2(n1211), .A3(n1212), .ZN(n1194) );
XNOR2_X1 U923 ( .A(G902), .B(KEYINPUT50), .ZN(n1212) );
NAND2_X1 U924 ( .A1(G237), .A2(G234), .ZN(n1211) );
NAND2_X1 U925 ( .A1(G221), .A2(n1213), .ZN(n1034) );
INV_X1 U926 ( .A(n1015), .ZN(n1209) );
NAND2_X1 U927 ( .A1(n1041), .A2(n1040), .ZN(n1015) );
NAND2_X1 U928 ( .A1(n1052), .A2(n1051), .ZN(n1040) );
NAND2_X1 U929 ( .A1(n1214), .A2(n1215), .ZN(n1051) );
NAND2_X1 U930 ( .A1(G210), .A2(n1216), .ZN(n1215) );
INV_X1 U931 ( .A(n1217), .ZN(n1214) );
NAND3_X1 U932 ( .A1(n1216), .A2(n1217), .A3(G210), .ZN(n1052) );
NAND2_X1 U933 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U934 ( .A(n1144), .B(n1220), .Z(n1219) );
XOR2_X1 U935 ( .A(KEYINPUT27), .B(KEYINPUT14), .Z(n1220) );
XOR2_X1 U936 ( .A(n1221), .B(n1222), .Z(n1144) );
XOR2_X1 U937 ( .A(n1223), .B(n1224), .Z(n1222) );
XNOR2_X1 U938 ( .A(KEYINPUT54), .B(n1078), .ZN(n1224) );
NOR2_X1 U939 ( .A1(G953), .A2(n1086), .ZN(n1223) );
INV_X1 U940 ( .A(G224), .ZN(n1086) );
XNOR2_X1 U941 ( .A(n1091), .B(n1225), .ZN(n1221) );
XOR2_X1 U942 ( .A(n1226), .B(n1227), .Z(n1091) );
XOR2_X1 U943 ( .A(n1228), .B(n1229), .Z(n1227) );
NOR2_X1 U944 ( .A1(KEYINPUT53), .A2(n1230), .ZN(n1228) );
XOR2_X1 U945 ( .A(n1231), .B(n1232), .Z(n1226) );
XNOR2_X1 U946 ( .A(n1233), .B(G101), .ZN(n1232) );
NAND2_X1 U947 ( .A1(n1234), .A2(n1235), .ZN(n1231) );
OR2_X1 U948 ( .A1(n1236), .A2(G113), .ZN(n1235) );
XOR2_X1 U949 ( .A(n1237), .B(KEYINPUT49), .Z(n1234) );
NAND2_X1 U950 ( .A1(G113), .A2(n1236), .ZN(n1237) );
XNOR2_X1 U951 ( .A(n1238), .B(KEYINPUT25), .ZN(n1236) );
NAND2_X1 U952 ( .A1(G214), .A2(n1216), .ZN(n1041) );
NAND2_X1 U953 ( .A1(n1239), .A2(n1240), .ZN(n1216) );
INV_X1 U954 ( .A(n1035), .ZN(n1190) );
XNOR2_X1 U955 ( .A(n1241), .B(n1242), .ZN(n1035) );
XNOR2_X1 U956 ( .A(KEYINPUT61), .B(n1142), .ZN(n1242) );
INV_X1 U957 ( .A(G469), .ZN(n1142) );
NAND2_X1 U958 ( .A1(n1243), .A2(n1218), .ZN(n1241) );
XOR2_X1 U959 ( .A(n1244), .B(n1245), .Z(n1243) );
XNOR2_X1 U960 ( .A(n1135), .B(n1076), .ZN(n1245) );
XOR2_X1 U961 ( .A(n1246), .B(n1247), .Z(n1244) );
NOR2_X1 U962 ( .A1(KEYINPUT23), .A2(n1138), .ZN(n1247) );
XNOR2_X1 U963 ( .A(G101), .B(n1248), .ZN(n1138) );
NOR2_X1 U964 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
NOR3_X1 U965 ( .A1(KEYINPUT43), .A2(G107), .A3(n1251), .ZN(n1250) );
NOR2_X1 U966 ( .A1(n1229), .A2(n1252), .ZN(n1249) );
INV_X1 U967 ( .A(KEYINPUT43), .ZN(n1252) );
XNOR2_X1 U968 ( .A(n1251), .B(G107), .ZN(n1229) );
INV_X1 U969 ( .A(G104), .ZN(n1251) );
NAND2_X1 U970 ( .A1(n1141), .A2(n1140), .ZN(n1246) );
NAND2_X1 U971 ( .A1(n1253), .A2(n1254), .ZN(n1140) );
NAND2_X1 U972 ( .A1(G227), .A2(n1043), .ZN(n1254) );
XNOR2_X1 U973 ( .A(G140), .B(n1230), .ZN(n1253) );
NAND3_X1 U974 ( .A1(n1255), .A2(n1043), .A3(G227), .ZN(n1141) );
XNOR2_X1 U975 ( .A(n1082), .B(n1230), .ZN(n1255) );
NOR3_X1 U976 ( .A1(n1032), .A2(n1031), .A3(n1018), .ZN(n1066) );
INV_X1 U977 ( .A(n1046), .ZN(n1018) );
NOR2_X1 U978 ( .A1(n1198), .A2(n1197), .ZN(n1046) );
XOR2_X1 U979 ( .A(n1256), .B(n1108), .Z(n1197) );
INV_X1 U980 ( .A(G475), .ZN(n1108) );
OR2_X1 U981 ( .A1(n1107), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U982 ( .A(n1258), .B(n1259), .ZN(n1107) );
XNOR2_X1 U983 ( .A(G104), .B(n1260), .ZN(n1259) );
NAND2_X1 U984 ( .A1(KEYINPUT5), .A2(n1261), .ZN(n1260) );
XNOR2_X1 U985 ( .A(n1233), .B(G113), .ZN(n1261) );
NAND2_X1 U986 ( .A1(n1262), .A2(KEYINPUT21), .ZN(n1258) );
XOR2_X1 U987 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U988 ( .A(G131), .B(n1265), .Z(n1264) );
NOR3_X1 U989 ( .A1(n1266), .A2(KEYINPUT17), .A3(n1267), .ZN(n1265) );
NOR2_X1 U990 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
XNOR2_X1 U991 ( .A(G125), .B(KEYINPUT60), .ZN(n1269) );
NOR2_X1 U992 ( .A1(n1270), .A2(G125), .ZN(n1268) );
NOR2_X1 U993 ( .A1(KEYINPUT59), .A2(G140), .ZN(n1270) );
NOR2_X1 U994 ( .A1(n1271), .A2(n1082), .ZN(n1266) );
NOR2_X1 U995 ( .A1(KEYINPUT59), .A2(G125), .ZN(n1271) );
XOR2_X1 U996 ( .A(n1272), .B(n1273), .Z(n1263) );
NAND3_X1 U997 ( .A1(n1240), .A2(n1043), .A3(G214), .ZN(n1272) );
INV_X1 U998 ( .A(n1176), .ZN(n1198) );
XOR2_X1 U999 ( .A(n1274), .B(G478), .Z(n1176) );
OR2_X1 U1000 ( .A1(n1103), .A2(n1257), .ZN(n1274) );
XNOR2_X1 U1001 ( .A(n1275), .B(n1276), .ZN(n1103) );
NOR2_X1 U1002 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
INV_X1 U1003 ( .A(G217), .ZN(n1277) );
NAND2_X1 U1004 ( .A1(n1279), .A2(n1280), .ZN(n1275) );
NAND2_X1 U1005 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U1006 ( .A(KEYINPUT63), .B(n1283), .Z(n1279) );
NOR2_X1 U1007 ( .A1(n1281), .A2(n1282), .ZN(n1283) );
XOR2_X1 U1008 ( .A(n1284), .B(n1285), .Z(n1282) );
XNOR2_X1 U1009 ( .A(n1286), .B(G128), .ZN(n1285) );
XNOR2_X1 U1010 ( .A(G143), .B(KEYINPUT1), .ZN(n1284) );
XOR2_X1 U1011 ( .A(n1287), .B(n1288), .Z(n1281) );
XNOR2_X1 U1012 ( .A(n1289), .B(G107), .ZN(n1288) );
INV_X1 U1013 ( .A(G116), .ZN(n1289) );
NAND2_X1 U1014 ( .A1(KEYINPUT24), .A2(n1233), .ZN(n1287) );
INV_X1 U1015 ( .A(G122), .ZN(n1233) );
INV_X1 U1016 ( .A(n1180), .ZN(n1031) );
XNOR2_X1 U1017 ( .A(n1053), .B(n1290), .ZN(n1180) );
XOR2_X1 U1018 ( .A(KEYINPUT56), .B(n1056), .Z(n1290) );
NOR2_X1 U1019 ( .A1(n1257), .A2(n1096), .ZN(n1056) );
XNOR2_X1 U1020 ( .A(n1291), .B(n1292), .ZN(n1096) );
XOR2_X1 U1021 ( .A(n1293), .B(n1294), .Z(n1292) );
NOR2_X1 U1022 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
AND2_X1 U1023 ( .A1(G137), .A2(n1297), .ZN(n1296) );
NOR2_X1 U1024 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
XNOR2_X1 U1025 ( .A(G137), .B(KEYINPUT2), .ZN(n1298) );
NOR2_X1 U1026 ( .A1(n1278), .A2(n1299), .ZN(n1297) );
XNOR2_X1 U1027 ( .A(KEYINPUT41), .B(G221), .ZN(n1299) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1043), .ZN(n1278) );
NOR2_X1 U1029 ( .A1(KEYINPUT30), .A2(n1300), .ZN(n1293) );
INV_X1 U1030 ( .A(n1230), .ZN(n1300) );
XOR2_X1 U1031 ( .A(G110), .B(KEYINPUT28), .Z(n1230) );
XOR2_X1 U1032 ( .A(n1301), .B(n1302), .Z(n1291) );
NOR2_X1 U1033 ( .A1(KEYINPUT39), .A2(n1303), .ZN(n1302) );
XNOR2_X1 U1034 ( .A(G146), .B(n1304), .ZN(n1303) );
NAND3_X1 U1035 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1304) );
NAND2_X1 U1036 ( .A1(KEYINPUT62), .A2(G125), .ZN(n1307) );
NAND3_X1 U1037 ( .A1(n1078), .A2(n1308), .A3(G140), .ZN(n1306) );
INV_X1 U1038 ( .A(G125), .ZN(n1078) );
NAND2_X1 U1039 ( .A1(n1309), .A2(n1082), .ZN(n1305) );
INV_X1 U1040 ( .A(G140), .ZN(n1082) );
NAND2_X1 U1041 ( .A1(n1310), .A2(n1308), .ZN(n1309) );
INV_X1 U1042 ( .A(KEYINPUT62), .ZN(n1308) );
XNOR2_X1 U1043 ( .A(G125), .B(KEYINPUT40), .ZN(n1310) );
XNOR2_X1 U1044 ( .A(G119), .B(G128), .ZN(n1301) );
NAND2_X1 U1045 ( .A1(G217), .A2(n1213), .ZN(n1053) );
NAND2_X1 U1046 ( .A1(G234), .A2(n1239), .ZN(n1213) );
INV_X1 U1047 ( .A(G902), .ZN(n1239) );
INV_X1 U1048 ( .A(n1179), .ZN(n1032) );
XNOR2_X1 U1049 ( .A(n1311), .B(n1312), .ZN(n1179) );
XNOR2_X1 U1050 ( .A(KEYINPUT29), .B(n1118), .ZN(n1312) );
INV_X1 U1051 ( .A(G472), .ZN(n1118) );
NAND2_X1 U1052 ( .A1(n1313), .A2(n1218), .ZN(n1311) );
INV_X1 U1053 ( .A(n1257), .ZN(n1218) );
XOR2_X1 U1054 ( .A(G902), .B(KEYINPUT38), .Z(n1257) );
XNOR2_X1 U1055 ( .A(n1117), .B(n1314), .ZN(n1313) );
XOR2_X1 U1056 ( .A(n1126), .B(n1315), .Z(n1314) );
NOR2_X1 U1057 ( .A1(G101), .A2(KEYINPUT12), .ZN(n1315) );
NAND3_X1 U1058 ( .A1(n1240), .A2(n1043), .A3(G210), .ZN(n1126) );
INV_X1 U1059 ( .A(G953), .ZN(n1043) );
INV_X1 U1060 ( .A(G237), .ZN(n1240) );
XNOR2_X1 U1061 ( .A(n1316), .B(n1317), .ZN(n1117) );
XOR2_X1 U1062 ( .A(n1238), .B(n1225), .Z(n1317) );
NAND2_X1 U1063 ( .A1(n1318), .A2(n1319), .ZN(n1225) );
NAND3_X1 U1064 ( .A1(G128), .A2(n1273), .A3(n1320), .ZN(n1319) );
INV_X1 U1065 ( .A(KEYINPUT46), .ZN(n1320) );
NAND2_X1 U1066 ( .A1(n1076), .A2(KEYINPUT46), .ZN(n1318) );
XOR2_X1 U1067 ( .A(G128), .B(n1273), .Z(n1076) );
XNOR2_X1 U1068 ( .A(n1178), .B(G146), .ZN(n1273) );
INV_X1 U1069 ( .A(G143), .ZN(n1178) );
XNOR2_X1 U1070 ( .A(G116), .B(G119), .ZN(n1238) );
XOR2_X1 U1071 ( .A(n1135), .B(G113), .Z(n1316) );
NAND2_X1 U1072 ( .A1(n1321), .A2(n1322), .ZN(n1135) );
NAND3_X1 U1073 ( .A1(KEYINPUT18), .A2(G137), .A3(n1323), .ZN(n1322) );
XOR2_X1 U1074 ( .A(n1324), .B(G131), .Z(n1323) );
NAND2_X1 U1075 ( .A1(KEYINPUT31), .A2(n1286), .ZN(n1324) );
INV_X1 U1076 ( .A(G134), .ZN(n1286) );
NAND2_X1 U1077 ( .A1(n1325), .A2(n1326), .ZN(n1321) );
NAND2_X1 U1078 ( .A1(KEYINPUT18), .A2(G137), .ZN(n1326) );
XOR2_X1 U1079 ( .A(n1327), .B(G131), .Z(n1325) );
NAND2_X1 U1080 ( .A1(G134), .A2(KEYINPUT31), .ZN(n1327) );
endmodule


