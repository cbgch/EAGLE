//Key = 1101110001110011110001100110110010111000101100011000111000110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273;

XOR2_X1 U700 ( .A(G107), .B(n968), .Z(G9) );
NOR2_X1 U701 ( .A1(n969), .A2(n970), .ZN(G75) );
NOR4_X1 U702 ( .A1(G953), .A2(n971), .A3(n972), .A4(n973), .ZN(n970) );
NOR3_X1 U703 ( .A1(n974), .A2(n975), .A3(n976), .ZN(n972) );
NOR2_X1 U704 ( .A1(n977), .A2(n978), .ZN(n976) );
NOR2_X1 U705 ( .A1(n979), .A2(n980), .ZN(n978) );
NOR3_X1 U706 ( .A1(n981), .A2(n982), .A3(n983), .ZN(n979) );
NOR2_X1 U707 ( .A1(n984), .A2(n985), .ZN(n983) );
NOR2_X1 U708 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U709 ( .A1(n988), .A2(n989), .ZN(n987) );
NOR2_X1 U710 ( .A1(n990), .A2(n991), .ZN(n988) );
NOR2_X1 U711 ( .A1(n992), .A2(n993), .ZN(n990) );
NOR2_X1 U712 ( .A1(n994), .A2(n995), .ZN(n986) );
NOR2_X1 U713 ( .A1(n996), .A2(n997), .ZN(n994) );
NOR2_X1 U714 ( .A1(n998), .A2(n999), .ZN(n996) );
NOR3_X1 U715 ( .A1(n995), .A2(n1000), .A3(n1001), .ZN(n982) );
XNOR2_X1 U716 ( .A(n1002), .B(KEYINPUT7), .ZN(n1000) );
NOR2_X1 U717 ( .A1(n989), .A2(n1003), .ZN(n981) );
NOR4_X1 U718 ( .A1(n1004), .A2(n989), .A3(n985), .A4(n995), .ZN(n977) );
NOR2_X1 U719 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NOR2_X1 U720 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR3_X1 U721 ( .A1(n971), .A2(G953), .A3(G952), .ZN(n969) );
AND4_X1 U722 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1007), .ZN(n971) );
INV_X1 U723 ( .A(n1012), .ZN(n1007) );
NOR2_X1 U724 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
XOR2_X1 U725 ( .A(n1015), .B(KEYINPUT18), .Z(n1013) );
NAND4_X1 U726 ( .A1(n1016), .A2(n1017), .A3(n999), .A4(n993), .ZN(n1015) );
XOR2_X1 U727 ( .A(n1018), .B(n1019), .Z(n1017) );
XNOR2_X1 U728 ( .A(G469), .B(KEYINPUT59), .ZN(n1019) );
NAND2_X1 U729 ( .A1(KEYINPUT61), .A2(n1020), .ZN(n1018) );
XNOR2_X1 U730 ( .A(n1021), .B(n1022), .ZN(n1016) );
NOR2_X1 U731 ( .A1(KEYINPUT56), .A2(n1023), .ZN(n1022) );
XNOR2_X1 U732 ( .A(n1024), .B(n1025), .ZN(n1009) );
XNOR2_X1 U733 ( .A(KEYINPUT6), .B(KEYINPUT45), .ZN(n1024) );
XOR2_X1 U734 ( .A(n1026), .B(n1027), .Z(G72) );
NOR2_X1 U735 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
AND2_X1 U736 ( .A1(G227), .A2(G900), .ZN(n1028) );
NAND2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1026) );
NAND3_X1 U738 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
INV_X1 U739 ( .A(n1035), .ZN(n1034) );
XOR2_X1 U740 ( .A(n1036), .B(n1037), .Z(n1033) );
NAND2_X1 U741 ( .A1(G953), .A2(n1038), .ZN(n1032) );
XOR2_X1 U742 ( .A(n1039), .B(KEYINPUT31), .Z(n1030) );
NAND3_X1 U743 ( .A1(n1035), .A2(n1029), .A3(n1040), .ZN(n1039) );
XNOR2_X1 U744 ( .A(n1036), .B(n1037), .ZN(n1040) );
NAND2_X1 U745 ( .A1(KEYINPUT1), .A2(n1041), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1036) );
NAND2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
XOR2_X1 U748 ( .A(n1046), .B(KEYINPUT12), .Z(n1042) );
OR2_X1 U749 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
XNOR2_X1 U750 ( .A(KEYINPUT51), .B(n1047), .ZN(n1044) );
XNOR2_X1 U751 ( .A(n1048), .B(n1049), .ZN(n1045) );
XOR2_X1 U752 ( .A(KEYINPUT4), .B(KEYINPUT2), .Z(n1049) );
XOR2_X1 U753 ( .A(n1050), .B(n1051), .Z(G69) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
XOR2_X1 U755 ( .A(n1054), .B(KEYINPUT35), .Z(n1053) );
NAND2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U757 ( .A1(n1055), .A2(n1056), .ZN(n1052) );
NAND2_X1 U758 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
XNOR2_X1 U759 ( .A(G953), .B(KEYINPUT13), .ZN(n1057) );
AND2_X1 U760 ( .A1(n1059), .A2(n1060), .ZN(n1055) );
NAND2_X1 U761 ( .A1(G953), .A2(n1061), .ZN(n1060) );
XOR2_X1 U762 ( .A(n1062), .B(n1063), .Z(n1059) );
XOR2_X1 U763 ( .A(n1064), .B(KEYINPUT29), .Z(n1062) );
NAND2_X1 U764 ( .A1(G953), .A2(n1065), .ZN(n1050) );
NAND2_X1 U765 ( .A1(G898), .A2(G224), .ZN(n1065) );
NOR2_X1 U766 ( .A1(n1066), .A2(n1067), .ZN(G66) );
XOR2_X1 U767 ( .A(n1068), .B(n1069), .Z(n1067) );
XOR2_X1 U768 ( .A(n1070), .B(KEYINPUT30), .Z(n1068) );
NAND3_X1 U769 ( .A1(n1071), .A2(G902), .A3(n1072), .ZN(n1070) );
XOR2_X1 U770 ( .A(n973), .B(KEYINPUT46), .Z(n1072) );
NOR3_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(G63) );
AND2_X1 U772 ( .A1(KEYINPUT47), .A2(n1066), .ZN(n1075) );
NOR3_X1 U773 ( .A1(KEYINPUT47), .A2(G953), .A3(G952), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1073) );
XOR2_X1 U775 ( .A(n1078), .B(KEYINPUT11), .Z(n1077) );
NAND2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XOR2_X1 U777 ( .A(n1081), .B(KEYINPUT20), .Z(n1079) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1076) );
XNOR2_X1 U779 ( .A(KEYINPUT54), .B(n1080), .ZN(n1082) );
NAND2_X1 U780 ( .A1(n1083), .A2(G478), .ZN(n1081) );
NOR2_X1 U781 ( .A1(n1066), .A2(n1084), .ZN(G60) );
XOR2_X1 U782 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U783 ( .A1(n1083), .A2(G475), .ZN(n1085) );
XOR2_X1 U784 ( .A(G104), .B(n1087), .Z(G6) );
NOR2_X1 U785 ( .A1(n1066), .A2(n1088), .ZN(G57) );
NOR2_X1 U786 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XOR2_X1 U787 ( .A(n1091), .B(KEYINPUT62), .Z(n1090) );
NAND2_X1 U788 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U789 ( .A1(n1092), .A2(n1093), .ZN(n1089) );
XNOR2_X1 U790 ( .A(n1094), .B(n1095), .ZN(n1093) );
NOR2_X1 U791 ( .A1(KEYINPUT38), .A2(n1096), .ZN(n1095) );
NOR3_X1 U792 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NOR2_X1 U793 ( .A1(KEYINPUT24), .A2(n1100), .ZN(n1099) );
NOR2_X1 U794 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U795 ( .A1(KEYINPUT5), .A2(n1103), .ZN(n1102) );
AND3_X1 U796 ( .A1(n1103), .A2(n1104), .A3(KEYINPUT5), .ZN(n1101) );
NOR2_X1 U797 ( .A1(n1105), .A2(n1106), .ZN(n1098) );
INV_X1 U798 ( .A(KEYINPUT24), .ZN(n1106) );
NOR2_X1 U799 ( .A1(n1107), .A2(n1108), .ZN(n1105) );
XOR2_X1 U800 ( .A(n1103), .B(KEYINPUT5), .Z(n1107) );
NOR2_X1 U801 ( .A1(n1104), .A2(n1103), .ZN(n1097) );
NAND2_X1 U802 ( .A1(n1083), .A2(G472), .ZN(n1094) );
INV_X1 U803 ( .A(n1109), .ZN(n1083) );
NOR2_X1 U804 ( .A1(n1066), .A2(n1110), .ZN(G54) );
XOR2_X1 U805 ( .A(n1111), .B(n1112), .Z(n1110) );
NAND3_X1 U806 ( .A1(G469), .A2(G902), .A3(n1113), .ZN(n1112) );
XOR2_X1 U807 ( .A(n973), .B(KEYINPUT27), .Z(n1113) );
NAND2_X1 U808 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U809 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U810 ( .A(KEYINPUT63), .B(n1118), .Z(n1114) );
NOR2_X1 U811 ( .A1(n1117), .A2(n1116), .ZN(n1118) );
XOR2_X1 U812 ( .A(n1119), .B(n1120), .Z(n1116) );
NAND2_X1 U813 ( .A1(n1121), .A2(KEYINPUT53), .ZN(n1119) );
XOR2_X1 U814 ( .A(n1122), .B(KEYINPUT52), .Z(n1121) );
NOR2_X1 U815 ( .A1(n1066), .A2(n1123), .ZN(G51) );
XOR2_X1 U816 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U817 ( .A1(n1126), .A2(n1109), .ZN(n1125) );
NAND2_X1 U818 ( .A1(G902), .A2(n973), .ZN(n1109) );
OR2_X1 U819 ( .A1(n1058), .A2(n1035), .ZN(n973) );
NAND4_X1 U820 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1035) );
NOR4_X1 U821 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1130) );
NOR2_X1 U822 ( .A1(KEYINPUT19), .A2(n1135), .ZN(n1134) );
AND2_X1 U823 ( .A1(n1136), .A2(n1137), .ZN(n1129) );
NAND2_X1 U824 ( .A1(n1138), .A2(n1139), .ZN(n1127) );
NAND2_X1 U825 ( .A1(n1140), .A2(n1003), .ZN(n1139) );
NAND3_X1 U826 ( .A1(n1141), .A2(n1142), .A3(KEYINPUT19), .ZN(n1140) );
NAND2_X1 U827 ( .A1(n1143), .A2(n1144), .ZN(n1058) );
NOR4_X1 U828 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1087), .ZN(n1144) );
AND3_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1087) );
NOR4_X1 U830 ( .A1(n968), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1143) );
INV_X1 U831 ( .A(n1154), .ZN(n1151) );
AND3_X1 U832 ( .A1(n1155), .A2(n1149), .A3(n1148), .ZN(n968) );
NAND2_X1 U833 ( .A1(n1156), .A2(KEYINPUT15), .ZN(n1124) );
XNOR2_X1 U834 ( .A(n1157), .B(n1158), .ZN(n1156) );
NOR2_X1 U835 ( .A1(n1029), .A2(G952), .ZN(n1066) );
XNOR2_X1 U836 ( .A(G146), .B(n1128), .ZN(G48) );
NAND3_X1 U837 ( .A1(n1150), .A2(n991), .A3(n1159), .ZN(n1128) );
XNOR2_X1 U838 ( .A(n1160), .B(n1135), .ZN(G45) );
NAND3_X1 U839 ( .A1(n1141), .A2(n991), .A3(n1138), .ZN(n1135) );
NAND2_X1 U840 ( .A1(KEYINPUT10), .A2(n1161), .ZN(n1160) );
XNOR2_X1 U841 ( .A(n1162), .B(n1163), .ZN(G42) );
NOR2_X1 U842 ( .A1(KEYINPUT50), .A2(n1137), .ZN(n1163) );
NAND3_X1 U843 ( .A1(n1164), .A2(n997), .A3(n1165), .ZN(n1137) );
INV_X1 U844 ( .A(n1003), .ZN(n1165) );
XOR2_X1 U845 ( .A(G137), .B(n1133), .Z(G39) );
AND3_X1 U846 ( .A1(n1159), .A2(n1166), .A3(n1167), .ZN(n1133) );
XOR2_X1 U847 ( .A(n1168), .B(n1132), .Z(G36) );
AND3_X1 U848 ( .A1(n1167), .A2(n1155), .A3(n1138), .ZN(n1132) );
NAND2_X1 U849 ( .A1(KEYINPUT26), .A2(n1169), .ZN(n1168) );
NAND3_X1 U850 ( .A1(n1170), .A2(n1171), .A3(n1172), .ZN(G33) );
NAND2_X1 U851 ( .A1(G131), .A2(n1173), .ZN(n1172) );
NAND2_X1 U852 ( .A1(n1174), .A2(KEYINPUT34), .ZN(n1173) );
XNOR2_X1 U853 ( .A(n1175), .B(KEYINPUT28), .ZN(n1174) );
NAND3_X1 U854 ( .A1(KEYINPUT34), .A2(n1176), .A3(n1175), .ZN(n1171) );
OR2_X1 U855 ( .A1(n1175), .A2(KEYINPUT34), .ZN(n1170) );
AND3_X1 U856 ( .A1(n1177), .A2(n1178), .A3(n1138), .ZN(n1175) );
AND3_X1 U857 ( .A1(n997), .A2(n1179), .A3(n1006), .ZN(n1138) );
NAND2_X1 U858 ( .A1(KEYINPUT14), .A2(n1003), .ZN(n1178) );
NAND2_X1 U859 ( .A1(n1167), .A2(n1150), .ZN(n1003) );
INV_X1 U860 ( .A(n995), .ZN(n1167) );
NAND2_X1 U861 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
INV_X1 U862 ( .A(KEYINPUT14), .ZN(n1181) );
NAND2_X1 U863 ( .A1(n1150), .A2(n995), .ZN(n1180) );
NAND2_X1 U864 ( .A1(n1182), .A2(n993), .ZN(n995) );
INV_X1 U865 ( .A(n992), .ZN(n1182) );
XNOR2_X1 U866 ( .A(G128), .B(n1183), .ZN(G30) );
NOR2_X1 U867 ( .A1(n1131), .A2(KEYINPUT37), .ZN(n1183) );
AND3_X1 U868 ( .A1(n1155), .A2(n991), .A3(n1159), .ZN(n1131) );
AND4_X1 U869 ( .A1(n997), .A2(n1012), .A3(n1008), .A4(n1179), .ZN(n1159) );
XOR2_X1 U870 ( .A(G101), .B(n1147), .Z(G3) );
AND3_X1 U871 ( .A1(n1006), .A2(n1148), .A3(n1166), .ZN(n1147) );
AND2_X1 U872 ( .A1(n1184), .A2(n997), .ZN(n1148) );
XNOR2_X1 U873 ( .A(G125), .B(n1136), .ZN(G27) );
NAND4_X1 U874 ( .A1(n1164), .A2(n1150), .A3(n1002), .A4(n991), .ZN(n1136) );
AND3_X1 U875 ( .A1(n1012), .A2(n1179), .A3(n1025), .ZN(n1164) );
NAND2_X1 U876 ( .A1(n1185), .A2(n1186), .ZN(n1179) );
NAND2_X1 U877 ( .A1(n1187), .A2(n1038), .ZN(n1186) );
INV_X1 U878 ( .A(G900), .ZN(n1038) );
XOR2_X1 U879 ( .A(G122), .B(n1153), .Z(G24) );
AND4_X1 U880 ( .A1(n1141), .A2(n1002), .A3(n1149), .A4(n1184), .ZN(n1153) );
INV_X1 U881 ( .A(n980), .ZN(n1149) );
NAND2_X1 U882 ( .A1(n1188), .A2(n1025), .ZN(n980) );
AND2_X1 U883 ( .A1(n1189), .A2(n1014), .ZN(n1141) );
XOR2_X1 U884 ( .A(G119), .B(n1152), .Z(G21) );
AND3_X1 U885 ( .A1(n1002), .A2(n1008), .A3(n1190), .ZN(n1152) );
XNOR2_X1 U886 ( .A(n1191), .B(n1146), .ZN(G18) );
AND2_X1 U887 ( .A1(n1192), .A2(n1155), .ZN(n1146) );
INV_X1 U888 ( .A(n1001), .ZN(n1155) );
NAND2_X1 U889 ( .A1(n1189), .A2(n1193), .ZN(n1001) );
XNOR2_X1 U890 ( .A(n1194), .B(n1145), .ZN(G15) );
AND2_X1 U891 ( .A1(n1192), .A2(n1150), .ZN(n1145) );
AND2_X1 U892 ( .A1(n1195), .A2(n1014), .ZN(n1150) );
XNOR2_X1 U893 ( .A(KEYINPUT58), .B(n1010), .ZN(n1195) );
AND3_X1 U894 ( .A1(n1002), .A2(n1184), .A3(n1006), .ZN(n1192) );
AND2_X1 U895 ( .A1(n1188), .A2(n1008), .ZN(n1006) );
XNOR2_X1 U896 ( .A(n1012), .B(KEYINPUT33), .ZN(n1188) );
INV_X1 U897 ( .A(n989), .ZN(n1002) );
NAND2_X1 U898 ( .A1(n1196), .A2(n999), .ZN(n989) );
INV_X1 U899 ( .A(n998), .ZN(n1196) );
NAND2_X1 U900 ( .A1(n1197), .A2(n1198), .ZN(G12) );
NAND2_X1 U901 ( .A1(G110), .A2(n1154), .ZN(n1198) );
XOR2_X1 U902 ( .A(KEYINPUT17), .B(n1199), .Z(n1197) );
NOR2_X1 U903 ( .A1(G110), .A2(n1154), .ZN(n1199) );
NAND3_X1 U904 ( .A1(n1025), .A2(n997), .A3(n1190), .ZN(n1154) );
AND3_X1 U905 ( .A1(n1184), .A2(n1012), .A3(n1166), .ZN(n1190) );
INV_X1 U906 ( .A(n985), .ZN(n1166) );
NAND2_X1 U907 ( .A1(n1010), .A2(n1193), .ZN(n985) );
XOR2_X1 U908 ( .A(n1014), .B(KEYINPUT36), .Z(n1193) );
XNOR2_X1 U909 ( .A(n1200), .B(G475), .ZN(n1014) );
NAND2_X1 U910 ( .A1(n1086), .A2(n1201), .ZN(n1200) );
XNOR2_X1 U911 ( .A(n1202), .B(n1203), .ZN(n1086) );
XOR2_X1 U912 ( .A(n1204), .B(n1205), .Z(n1203) );
XNOR2_X1 U913 ( .A(n1176), .B(G122), .ZN(n1205) );
INV_X1 U914 ( .A(G131), .ZN(n1176) );
XNOR2_X1 U915 ( .A(G146), .B(n1161), .ZN(n1204) );
XOR2_X1 U916 ( .A(n1206), .B(n1207), .Z(n1202) );
XNOR2_X1 U917 ( .A(n1194), .B(G104), .ZN(n1207) );
INV_X1 U918 ( .A(G113), .ZN(n1194) );
XNOR2_X1 U919 ( .A(n1208), .B(n1041), .ZN(n1206) );
XNOR2_X1 U920 ( .A(n1209), .B(n1162), .ZN(n1041) );
NAND2_X1 U921 ( .A1(n1210), .A2(G214), .ZN(n1208) );
INV_X1 U922 ( .A(n1189), .ZN(n1010) );
XOR2_X1 U923 ( .A(G478), .B(n1211), .Z(n1189) );
AND2_X1 U924 ( .A1(n1201), .A2(n1080), .ZN(n1211) );
XOR2_X1 U925 ( .A(n1212), .B(n1213), .Z(n1080) );
XOR2_X1 U926 ( .A(G128), .B(n1214), .Z(n1213) );
XNOR2_X1 U927 ( .A(n1161), .B(G134), .ZN(n1214) );
INV_X1 U928 ( .A(G143), .ZN(n1161) );
XOR2_X1 U929 ( .A(n1215), .B(n1216), .Z(n1212) );
NOR2_X1 U930 ( .A1(KEYINPUT44), .A2(n1217), .ZN(n1216) );
XOR2_X1 U931 ( .A(G107), .B(n1218), .Z(n1217) );
XNOR2_X1 U932 ( .A(G122), .B(n1191), .ZN(n1218) );
NAND2_X1 U933 ( .A1(n1219), .A2(n1220), .ZN(n1215) );
XNOR2_X1 U934 ( .A(G217), .B(KEYINPUT22), .ZN(n1219) );
XNOR2_X1 U935 ( .A(n1221), .B(n1071), .ZN(n1012) );
AND2_X1 U936 ( .A1(G217), .A2(n1222), .ZN(n1071) );
NAND2_X1 U937 ( .A1(n1069), .A2(n1201), .ZN(n1221) );
XNOR2_X1 U938 ( .A(n1223), .B(n1224), .ZN(n1069) );
XNOR2_X1 U939 ( .A(n1225), .B(n1226), .ZN(n1224) );
XOR2_X1 U940 ( .A(n1227), .B(n1228), .Z(n1226) );
NOR2_X1 U941 ( .A1(KEYINPUT60), .A2(n1229), .ZN(n1228) );
XNOR2_X1 U942 ( .A(G140), .B(n1230), .ZN(n1229) );
NAND2_X1 U943 ( .A1(KEYINPUT32), .A2(n1209), .ZN(n1230) );
NAND2_X1 U944 ( .A1(n1220), .A2(G221), .ZN(n1227) );
AND2_X1 U945 ( .A1(G234), .A2(n1029), .ZN(n1220) );
XNOR2_X1 U946 ( .A(G110), .B(n1231), .ZN(n1223) );
XOR2_X1 U947 ( .A(G137), .B(G119), .Z(n1231) );
AND2_X1 U948 ( .A1(n991), .A2(n1232), .ZN(n1184) );
NAND2_X1 U949 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U950 ( .A1(n1187), .A2(n1061), .ZN(n1234) );
INV_X1 U951 ( .A(G898), .ZN(n1061) );
NOR3_X1 U952 ( .A1(n1029), .A2(n975), .A3(n1201), .ZN(n1187) );
INV_X1 U953 ( .A(n1235), .ZN(n975) );
XOR2_X1 U954 ( .A(n1185), .B(KEYINPUT41), .Z(n1233) );
NAND3_X1 U955 ( .A1(n1235), .A2(n1029), .A3(n1236), .ZN(n1185) );
XOR2_X1 U956 ( .A(KEYINPUT48), .B(n974), .Z(n1236) );
XOR2_X1 U957 ( .A(G952), .B(KEYINPUT0), .Z(n974) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1235) );
INV_X1 U959 ( .A(n1142), .ZN(n991) );
NAND2_X1 U960 ( .A1(n992), .A2(n993), .ZN(n1142) );
NAND2_X1 U961 ( .A1(G214), .A2(n1237), .ZN(n993) );
XNOR2_X1 U962 ( .A(n1238), .B(n1239), .ZN(n992) );
XNOR2_X1 U963 ( .A(KEYINPUT55), .B(n1023), .ZN(n1239) );
NAND2_X1 U964 ( .A1(n1240), .A2(n1201), .ZN(n1023) );
XOR2_X1 U965 ( .A(n1241), .B(n1158), .Z(n1240) );
AND2_X1 U966 ( .A1(n1242), .A2(n1243), .ZN(n1158) );
NAND3_X1 U967 ( .A1(G224), .A2(n1244), .A3(n1245), .ZN(n1243) );
XNOR2_X1 U968 ( .A(n1047), .B(G125), .ZN(n1245) );
NAND2_X1 U969 ( .A1(n1246), .A2(n1247), .ZN(n1242) );
NAND2_X1 U970 ( .A1(G224), .A2(n1244), .ZN(n1247) );
XNOR2_X1 U971 ( .A(KEYINPUT42), .B(n1029), .ZN(n1244) );
XNOR2_X1 U972 ( .A(n1209), .B(n1047), .ZN(n1246) );
INV_X1 U973 ( .A(G125), .ZN(n1209) );
NAND2_X1 U974 ( .A1(KEYINPUT43), .A2(n1157), .ZN(n1241) );
XNOR2_X1 U975 ( .A(n1064), .B(n1248), .ZN(n1157) );
NOR2_X1 U976 ( .A1(KEYINPUT57), .A2(n1063), .ZN(n1248) );
XNOR2_X1 U977 ( .A(n1249), .B(n1250), .ZN(n1063) );
XOR2_X1 U978 ( .A(KEYINPUT39), .B(G110), .Z(n1250) );
NAND2_X1 U979 ( .A1(n1251), .A2(KEYINPUT3), .ZN(n1249) );
XNOR2_X1 U980 ( .A(G122), .B(KEYINPUT40), .ZN(n1251) );
XOR2_X1 U981 ( .A(n1252), .B(n1253), .Z(n1064) );
XNOR2_X1 U982 ( .A(n1254), .B(KEYINPUT21), .ZN(n1253) );
NAND2_X1 U983 ( .A1(KEYINPUT25), .A2(n1191), .ZN(n1254) );
XNOR2_X1 U984 ( .A(n1255), .B(n1256), .ZN(n1252) );
NAND2_X1 U985 ( .A1(KEYINPUT9), .A2(n1021), .ZN(n1238) );
INV_X1 U986 ( .A(n1126), .ZN(n1021) );
NAND2_X1 U987 ( .A1(G210), .A2(n1237), .ZN(n1126) );
NAND2_X1 U988 ( .A1(n1257), .A2(n1201), .ZN(n1237) );
INV_X1 U989 ( .A(G237), .ZN(n1257) );
AND2_X1 U990 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND2_X1 U991 ( .A1(G221), .A2(n1222), .ZN(n999) );
NAND2_X1 U992 ( .A1(G234), .A2(n1201), .ZN(n1222) );
XOR2_X1 U993 ( .A(n1020), .B(G469), .Z(n998) );
AND2_X1 U994 ( .A1(n1258), .A2(n1201), .ZN(n1020) );
XOR2_X1 U995 ( .A(n1259), .B(n1120), .Z(n1258) );
XNOR2_X1 U996 ( .A(G110), .B(n1162), .ZN(n1120) );
INV_X1 U997 ( .A(G140), .ZN(n1162) );
XOR2_X1 U998 ( .A(n1117), .B(n1260), .Z(n1259) );
NOR2_X1 U999 ( .A1(KEYINPUT49), .A2(n1122), .ZN(n1260) );
NAND2_X1 U1000 ( .A1(G227), .A2(n1029), .ZN(n1122) );
XNOR2_X1 U1001 ( .A(n1256), .B(n1261), .ZN(n1117) );
XNOR2_X1 U1002 ( .A(KEYINPUT51), .B(n1104), .ZN(n1261) );
XNOR2_X1 U1003 ( .A(n1262), .B(n1263), .ZN(n1256) );
XNOR2_X1 U1004 ( .A(G104), .B(G107), .ZN(n1262) );
INV_X1 U1005 ( .A(n1008), .ZN(n1025) );
XNOR2_X1 U1006 ( .A(n1264), .B(G472), .ZN(n1008) );
NAND3_X1 U1007 ( .A1(n1265), .A2(n1266), .A3(n1201), .ZN(n1264) );
INV_X1 U1008 ( .A(G902), .ZN(n1201) );
NAND2_X1 U1009 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
INV_X1 U1010 ( .A(KEYINPUT8), .ZN(n1268) );
XOR2_X1 U1011 ( .A(n1269), .B(n1092), .Z(n1267) );
NAND3_X1 U1012 ( .A1(n1092), .A2(n1269), .A3(KEYINPUT8), .ZN(n1265) );
XNOR2_X1 U1013 ( .A(n1103), .B(n1104), .ZN(n1269) );
INV_X1 U1014 ( .A(n1108), .ZN(n1104) );
XOR2_X1 U1015 ( .A(n1048), .B(n1270), .Z(n1108) );
INV_X1 U1016 ( .A(n1047), .ZN(n1270) );
XOR2_X1 U1017 ( .A(G143), .B(n1225), .Z(n1047) );
XOR2_X1 U1018 ( .A(G128), .B(G146), .Z(n1225) );
XNOR2_X1 U1019 ( .A(G131), .B(n1271), .ZN(n1048) );
XNOR2_X1 U1020 ( .A(G137), .B(n1169), .ZN(n1271) );
INV_X1 U1021 ( .A(G134), .ZN(n1169) );
XOR2_X1 U1022 ( .A(n1191), .B(n1255), .Z(n1103) );
XOR2_X1 U1023 ( .A(G113), .B(G119), .Z(n1255) );
INV_X1 U1024 ( .A(G116), .ZN(n1191) );
XOR2_X1 U1025 ( .A(n1272), .B(n1263), .Z(n1092) );
XOR2_X1 U1026 ( .A(G101), .B(KEYINPUT16), .Z(n1263) );
NAND2_X1 U1027 ( .A1(n1210), .A2(G210), .ZN(n1272) );
AND2_X1 U1028 ( .A1(n1273), .A2(n1029), .ZN(n1210) );
INV_X1 U1029 ( .A(G953), .ZN(n1029) );
XNOR2_X1 U1030 ( .A(G237), .B(KEYINPUT23), .ZN(n1273) );
endmodule


