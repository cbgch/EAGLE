//Key = 1001000100110010110011000111110011011100001101100100000101011110


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
n2164;

OR2_X1 U1224 ( .A1(n1772), .A2(STATO_REG_0__SCAN_IN), .ZN(n1624) );
INV_X2 U1225 ( .A(n1624), .ZN(n1625) );
NOR4_X2 U1226 ( .A1(n1771), .A2(n2080), .A3(n2091), .A4(AVERAGE), .ZN(n1860));
INV_X2 U1227 ( .A(U280), .ZN(n1775) );
XNOR2_X1 U1228 ( .A(KEYINPUT19), .B(n1626), .ZN(U375) );
NAND2_X1 U1229 ( .A1(n1627), .A2(n1628), .ZN(U344) );
NAND2_X1 U1230 ( .A1(n1629), .A2(DATA_IN_7_), .ZN(n1628) );
XOR2_X1 U1231 ( .A(KEYINPUT11), .B(n1630), .Z(n1627) );
NOR2_X1 U1232 ( .A1(n1631), .A2(n1632), .ZN(n1630) );
XNOR2_X1 U1233 ( .A(KEYINPUT12), .B(n1633), .ZN(n1632) );
NAND2_X1 U1234 ( .A1(n1634), .A2(n1635), .ZN(U343) );
NAND2_X1 U1235 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1633), .ZN(n1635) );
NAND2_X1 U1236 ( .A1(n1629), .A2(DATA_IN_6_), .ZN(n1634) );
NAND2_X1 U1237 ( .A1(n1636), .A2(n1637), .ZN(U342) );
NAND2_X1 U1238 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1633), .ZN(n1637) );
NAND2_X1 U1239 ( .A1(n1629), .A2(DATA_IN_5_), .ZN(n1636) );
NAND2_X1 U1240 ( .A1(n1638), .A2(n1639), .ZN(U341) );
NAND2_X1 U1241 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1633), .ZN(n1639) );
NAND2_X1 U1242 ( .A1(n1629), .A2(DATA_IN_4_), .ZN(n1638) );
NAND2_X1 U1243 ( .A1(n1640), .A2(n1641), .ZN(U340) );
NAND2_X1 U1244 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1633), .ZN(n1641) );
NAND2_X1 U1245 ( .A1(n1629), .A2(DATA_IN_3_), .ZN(n1640) );
NAND2_X1 U1246 ( .A1(n1642), .A2(n1643), .ZN(U339) );
NAND2_X1 U1247 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1633), .ZN(n1643) );
NAND2_X1 U1248 ( .A1(n1629), .A2(DATA_IN_2_), .ZN(n1642) );
NAND2_X1 U1249 ( .A1(n1644), .A2(n1645), .ZN(U338) );
NAND2_X1 U1250 ( .A1(n1629), .A2(DATA_IN_1_), .ZN(n1645) );
NAND2_X1 U1251 ( .A1(n1646), .A2(n1633), .ZN(n1644) );
XNOR2_X1 U1252 ( .A(RMAX_REG_1__SCAN_IN), .B(KEYINPUT16), .ZN(n1646) );
NAND2_X1 U1253 ( .A1(n1647), .A2(n1648), .ZN(U337) );
NAND2_X1 U1254 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1633), .ZN(n1648) );
NAND2_X1 U1255 ( .A1(n1629), .A2(DATA_IN_0_), .ZN(n1647) );
INV_X1 U1256 ( .A(n1633), .ZN(n1629) );
NAND2_X1 U1257 ( .A1(n1626), .A2(n1649), .ZN(n1633) );
OR2_X1 U1258 ( .A1(n1650), .A2(STATO_REG_0__SCAN_IN), .ZN(n1649) );
NAND2_X1 U1259 ( .A1(n1651), .A2(n1652), .ZN(U336) );
NAND2_X1 U1260 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1653), .ZN(n1652) );
NAND2_X1 U1261 ( .A1(n1654), .A2(n1655), .ZN(n1651) );
XNOR2_X1 U1262 ( .A(KEYINPUT39), .B(n1656), .ZN(n1654) );
NAND2_X1 U1263 ( .A1(n1657), .A2(n1658), .ZN(U335) );
NAND2_X1 U1264 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1653), .ZN(n1658) );
NAND2_X1 U1265 ( .A1(n1655), .A2(DATA_IN_6_), .ZN(n1657) );
NAND2_X1 U1266 ( .A1(n1659), .A2(n1660), .ZN(U334) );
NAND2_X1 U1267 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1653), .ZN(n1660) );
NAND2_X1 U1268 ( .A1(n1655), .A2(DATA_IN_5_), .ZN(n1659) );
NAND2_X1 U1269 ( .A1(n1661), .A2(n1662), .ZN(U333) );
NAND2_X1 U1270 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1653), .ZN(n1662) );
NAND2_X1 U1271 ( .A1(n1655), .A2(DATA_IN_4_), .ZN(n1661) );
NAND2_X1 U1272 ( .A1(n1663), .A2(n1664), .ZN(U332) );
NAND2_X1 U1273 ( .A1(n1655), .A2(DATA_IN_3_), .ZN(n1664) );
NAND2_X1 U1274 ( .A1(n1665), .A2(n1653), .ZN(n1663) );
XNOR2_X1 U1275 ( .A(RMIN_REG_3__SCAN_IN), .B(KEYINPUT29), .ZN(n1665) );
NAND2_X1 U1276 ( .A1(n1666), .A2(n1667), .ZN(U331) );
NAND2_X1 U1277 ( .A1(n1655), .A2(DATA_IN_2_), .ZN(n1667) );
XOR2_X1 U1278 ( .A(n1668), .B(KEYINPUT47), .Z(n1666) );
NAND2_X1 U1279 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1653), .ZN(n1668) );
NAND2_X1 U1280 ( .A1(n1669), .A2(n1670), .ZN(U330) );
NAND2_X1 U1281 ( .A1(DATA_IN_1_), .A2(n1671), .ZN(n1670) );
XNOR2_X1 U1282 ( .A(KEYINPUT50), .B(n1653), .ZN(n1671) );
NAND2_X1 U1283 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1653), .ZN(n1669) );
NAND2_X1 U1284 ( .A1(n1672), .A2(n1673), .ZN(U329) );
NAND2_X1 U1285 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1653), .ZN(n1673) );
NAND2_X1 U1286 ( .A1(n1655), .A2(DATA_IN_0_), .ZN(n1672) );
INV_X1 U1287 ( .A(n1653), .ZN(n1655) );
NAND2_X1 U1288 ( .A1(n1626), .A2(n1674), .ZN(n1653) );
NAND2_X1 U1289 ( .A1(n1675), .A2(n1676), .ZN(n1674) );
NAND2_X1 U1290 ( .A1(n1677), .A2(n1678), .ZN(n1675) );
NAND2_X1 U1291 ( .A1(n1679), .A2(n1680), .ZN(n1678) );
NAND3_X1 U1292 ( .A1(n1681), .A2(n1682), .A3(n1683), .ZN(n1680) );
NAND2_X1 U1293 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1656), .ZN(n1683) );
NAND3_X1 U1294 ( .A1(n1684), .A2(n1685), .A3(n1686), .ZN(n1682) );
NAND2_X1 U1295 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1687), .ZN(n1686) );
NAND3_X1 U1296 ( .A1(n1688), .A2(n1689), .A3(n1690), .ZN(n1685) );
NAND2_X1 U1297 ( .A1(DATA_IN_5_), .A2(n1691), .ZN(n1690) );
NAND3_X1 U1298 ( .A1(n1692), .A2(n1693), .A3(n1694), .ZN(n1689) );
NAND2_X1 U1299 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1695), .ZN(n1694) );
NAND3_X1 U1300 ( .A1(n1696), .A2(n1697), .A3(n1698), .ZN(n1693) );
NAND2_X1 U1301 ( .A1(DATA_IN_2_), .A2(n1699), .ZN(n1698) );
NAND3_X1 U1302 ( .A1(n1700), .A2(n1701), .A3(n1702), .ZN(n1697) );
NAND2_X1 U1303 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1703), .ZN(n1702) );
NAND3_X1 U1304 ( .A1(n1704), .A2(n1705), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1701) );
NAND2_X1 U1305 ( .A1(n1706), .A2(DATA_IN_1_), .ZN(n1704) );
XOR2_X1 U1306 ( .A(n1707), .B(KEYINPUT33), .Z(n1706) );
XNOR2_X1 U1307 ( .A(RMIN_REG_1__SCAN_IN), .B(KEYINPUT35), .ZN(n1707) );
NAND2_X1 U1308 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1708), .ZN(n1700) );
NAND2_X1 U1309 ( .A1(n1709), .A2(n1710), .ZN(n1696) );
XNOR2_X1 U1310 ( .A(KEYINPUT5), .B(n1711), .ZN(n1709) );
NAND2_X1 U1311 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1711), .ZN(n1692) );
NAND2_X1 U1312 ( .A1(DATA_IN_4_), .A2(n1712), .ZN(n1688) );
NAND2_X1 U1313 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1713), .ZN(n1684) );
XNOR2_X1 U1314 ( .A(KEYINPUT3), .B(n1714), .ZN(n1713) );
NAND2_X1 U1315 ( .A1(DATA_IN_6_), .A2(n1715), .ZN(n1681) );
XOR2_X1 U1316 ( .A(RMIN_REG_6__SCAN_IN), .B(KEYINPUT27), .Z(n1715) );
NAND2_X1 U1317 ( .A1(DATA_IN_7_), .A2(n1716), .ZN(n1679) );
XOR2_X1 U1318 ( .A(n1650), .B(KEYINPUT28), .Z(n1677) );
NAND2_X1 U1319 ( .A1(n1717), .A2(n1718), .ZN(n1650) );
NAND2_X1 U1320 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1656), .ZN(n1718) );
INV_X1 U1321 ( .A(DATA_IN_7_), .ZN(n1656) );
NAND3_X1 U1322 ( .A1(n1719), .A2(n1720), .A3(n1721), .ZN(n1717) );
XOR2_X1 U1323 ( .A(n1722), .B(KEYINPUT18), .Z(n1721) );
NAND3_X1 U1324 ( .A1(n1723), .A2(n1724), .A3(n1725), .ZN(n1722) );
NAND2_X1 U1325 ( .A1(DATA_IN_5_), .A2(n1726), .ZN(n1725) );
NAND3_X1 U1326 ( .A1(n1727), .A2(n1728), .A3(n1729), .ZN(n1724) );
NAND2_X1 U1327 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1687), .ZN(n1729) );
NAND3_X1 U1328 ( .A1(n1730), .A2(n1731), .A3(n1732), .ZN(n1728) );
NAND2_X1 U1329 ( .A1(DATA_IN_3_), .A2(n1733), .ZN(n1732) );
NAND3_X1 U1330 ( .A1(n1734), .A2(n1735), .A3(n1736), .ZN(n1731) );
NAND2_X1 U1331 ( .A1(RMAX_REG_3__SCAN_IN), .A2(n1711), .ZN(n1736) );
NAND3_X1 U1332 ( .A1(n1737), .A2(n1738), .A3(n1739), .ZN(n1735) );
NAND2_X1 U1333 ( .A1(DATA_IN_2_), .A2(n1740), .ZN(n1739) );
NAND3_X1 U1334 ( .A1(n1741), .A2(n1742), .A3(DATA_IN_0_), .ZN(n1738) );
NAND2_X1 U1335 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1708), .ZN(n1741) );
NAND2_X1 U1336 ( .A1(DATA_IN_1_), .A2(n1743), .ZN(n1737) );
NAND2_X1 U1337 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1703), .ZN(n1734) );
NAND2_X1 U1338 ( .A1(DATA_IN_4_), .A2(n1744), .ZN(n1730) );
XNOR2_X1 U1339 ( .A(n1745), .B(KEYINPUT62), .ZN(n1744) );
NAND2_X1 U1340 ( .A1(n1746), .A2(RMAX_REG_4__SCAN_IN), .ZN(n1727) );
XNOR2_X1 U1341 ( .A(DATA_IN_4_), .B(KEYINPUT9), .ZN(n1746) );
NAND2_X1 U1342 ( .A1(n1747), .A2(n1748), .ZN(n1723) );
XNOR2_X1 U1343 ( .A(KEYINPUT48), .B(n1714), .ZN(n1747) );
NAND2_X1 U1344 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1714), .ZN(n1720) );
NAND2_X1 U1345 ( .A1(DATA_IN_7_), .A2(n1631), .ZN(n1719) );
NAND2_X1 U1346 ( .A1(n1749), .A2(n1750), .ZN(U328) );
NAND2_X1 U1347 ( .A1(DATA_IN_7_), .A2(n1751), .ZN(n1750) );
XOR2_X1 U1348 ( .A(KEYINPUT52), .B(n1752), .Z(n1751) );
NAND2_X1 U1349 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1753), .ZN(n1749) );
NAND2_X1 U1350 ( .A1(n1754), .A2(n1755), .ZN(U327) );
NAND2_X1 U1351 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1753), .ZN(n1755) );
XOR2_X1 U1352 ( .A(n1756), .B(KEYINPUT30), .Z(n1754) );
NAND2_X1 U1353 ( .A1(n1752), .A2(DATA_IN_6_), .ZN(n1756) );
NAND2_X1 U1354 ( .A1(n1757), .A2(n1758), .ZN(U326) );
NAND2_X1 U1355 ( .A1(n1752), .A2(DATA_IN_5_), .ZN(n1758) );
NAND2_X1 U1356 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1753), .ZN(n1757) );
NAND2_X1 U1357 ( .A1(n1759), .A2(n1760), .ZN(U325) );
NAND2_X1 U1358 ( .A1(n1752), .A2(DATA_IN_4_), .ZN(n1760) );
NAND2_X1 U1359 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1753), .ZN(n1759) );
NAND2_X1 U1360 ( .A1(n1761), .A2(n1762), .ZN(U324) );
NAND2_X1 U1361 ( .A1(n1752), .A2(DATA_IN_3_), .ZN(n1762) );
NAND2_X1 U1362 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1753), .ZN(n1761) );
NAND2_X1 U1363 ( .A1(n1763), .A2(n1764), .ZN(U323) );
NAND2_X1 U1364 ( .A1(n1752), .A2(DATA_IN_2_), .ZN(n1764) );
XOR2_X1 U1365 ( .A(n1765), .B(KEYINPUT2), .Z(n1763) );
NAND2_X1 U1366 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1753), .ZN(n1765) );
NAND2_X1 U1367 ( .A1(n1766), .A2(n1767), .ZN(U322) );
NAND2_X1 U1368 ( .A1(n1752), .A2(DATA_IN_1_), .ZN(n1767) );
NAND2_X1 U1369 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1753), .ZN(n1766) );
NAND2_X1 U1370 ( .A1(n1768), .A2(n1769), .ZN(U321) );
NAND2_X1 U1371 ( .A1(n1752), .A2(DATA_IN_0_), .ZN(n1769) );
AND2_X1 U1372 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1770), .ZN(n1752) );
NAND2_X1 U1373 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1753), .ZN(n1768) );
NAND2_X1 U1374 ( .A1(n1626), .A2(n1770), .ZN(n1753) );
NAND2_X1 U1375 ( .A1(n1676), .A2(n1771), .ZN(n1770) );
NAND2_X1 U1376 ( .A1(n1772), .A2(n1676), .ZN(n1626) );
INV_X1 U1377 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1676) );
NAND2_X1 U1378 ( .A1(n1773), .A2(n1774), .ZN(U320) );
NAND2_X1 U1379 ( .A1(n1625), .A2(DATA_IN_7_), .ZN(n1774) );
NAND2_X1 U1380 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1775), .ZN(n1773) );
NAND2_X1 U1381 ( .A1(n1776), .A2(n1777), .ZN(U319) );
NAND2_X1 U1382 ( .A1(n1625), .A2(DATA_IN_6_), .ZN(n1777) );
NAND2_X1 U1383 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1775), .ZN(n1776) );
NAND2_X1 U1384 ( .A1(n1778), .A2(n1779), .ZN(U318) );
NAND2_X1 U1385 ( .A1(n1625), .A2(DATA_IN_5_), .ZN(n1779) );
NAND2_X1 U1386 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1775), .ZN(n1778) );
NAND2_X1 U1387 ( .A1(n1780), .A2(n1781), .ZN(U317) );
NAND2_X1 U1388 ( .A1(n1782), .A2(DATA_IN_4_), .ZN(n1781) );
XNOR2_X1 U1389 ( .A(n1625), .B(KEYINPUT45), .ZN(n1782) );
NAND2_X1 U1390 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1775), .ZN(n1780) );
NAND2_X1 U1391 ( .A1(n1783), .A2(n1784), .ZN(U316) );
NAND2_X1 U1392 ( .A1(n1625), .A2(DATA_IN_3_), .ZN(n1784) );
NAND2_X1 U1393 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1775), .ZN(n1783) );
NAND2_X1 U1394 ( .A1(n1785), .A2(n1786), .ZN(U315) );
NAND2_X1 U1395 ( .A1(n1625), .A2(DATA_IN_2_), .ZN(n1786) );
NAND2_X1 U1396 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1775), .ZN(n1785) );
NAND2_X1 U1397 ( .A1(n1787), .A2(n1788), .ZN(U314) );
NAND2_X1 U1398 ( .A1(DATA_IN_1_), .A2(n1789), .ZN(n1788) );
XNOR2_X1 U1399 ( .A(KEYINPUT40), .B(n1624), .ZN(n1789) );
NAND2_X1 U1400 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1775), .ZN(n1787) );
NAND2_X1 U1401 ( .A1(n1790), .A2(n1791), .ZN(U313) );
NAND2_X1 U1402 ( .A1(n1625), .A2(DATA_IN_0_), .ZN(n1791) );
NAND2_X1 U1403 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1775), .ZN(n1790) );
NAND2_X1 U1404 ( .A1(n1792), .A2(n1793), .ZN(U312) );
NAND2_X1 U1405 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1794), .ZN(n1793) );
XNOR2_X1 U1406 ( .A(KEYINPUT8), .B(n1624), .ZN(n1794) );
NAND2_X1 U1407 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1775), .ZN(n1792) );
NAND2_X1 U1408 ( .A1(n1795), .A2(n1796), .ZN(U311) );
NAND2_X1 U1409 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1625), .ZN(n1796) );
NAND2_X1 U1410 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1775), .ZN(n1795) );
NAND2_X1 U1411 ( .A1(n1797), .A2(n1798), .ZN(U310) );
NAND2_X1 U1412 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1625), .ZN(n1798) );
NAND2_X1 U1413 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1775), .ZN(n1797) );
NAND2_X1 U1414 ( .A1(n1799), .A2(n1800), .ZN(U309) );
NAND2_X1 U1415 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1625), .ZN(n1800) );
NAND2_X1 U1416 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1775), .ZN(n1799) );
NAND2_X1 U1417 ( .A1(n1801), .A2(n1802), .ZN(U308) );
NAND2_X1 U1418 ( .A1(n1803), .A2(REG1_REG_3__SCAN_IN), .ZN(n1802) );
XNOR2_X1 U1419 ( .A(n1625), .B(KEYINPUT59), .ZN(n1803) );
NAND2_X1 U1420 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1775), .ZN(n1801) );
NAND2_X1 U1421 ( .A1(n1804), .A2(n1805), .ZN(U307) );
NAND2_X1 U1422 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1625), .ZN(n1805) );
NAND2_X1 U1423 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1775), .ZN(n1804) );
NAND2_X1 U1424 ( .A1(n1806), .A2(n1807), .ZN(U306) );
NAND2_X1 U1425 ( .A1(n1808), .A2(n1775), .ZN(n1807) );
XOR2_X1 U1426 ( .A(REG2_REG_1__SCAN_IN), .B(KEYINPUT15), .Z(n1808) );
NAND2_X1 U1427 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1625), .ZN(n1806) );
NAND2_X1 U1428 ( .A1(n1809), .A2(n1810), .ZN(U305) );
NAND2_X1 U1429 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1625), .ZN(n1810) );
NAND2_X1 U1430 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1775), .ZN(n1809) );
NAND2_X1 U1431 ( .A1(n1811), .A2(n1812), .ZN(U304) );
NAND2_X1 U1432 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1625), .ZN(n1812) );
NAND2_X1 U1433 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1775), .ZN(n1811) );
NAND2_X1 U1434 ( .A1(n1813), .A2(n1814), .ZN(U303) );
NAND2_X1 U1435 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1775), .ZN(n1814) );
XOR2_X1 U1436 ( .A(KEYINPUT60), .B(n1815), .Z(n1813) );
AND2_X1 U1437 ( .A1(n1625), .A2(REG2_REG_6__SCAN_IN), .ZN(n1815) );
NAND2_X1 U1438 ( .A1(n1816), .A2(n1817), .ZN(U302) );
NAND2_X1 U1439 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1625), .ZN(n1817) );
NAND2_X1 U1440 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1775), .ZN(n1816) );
NAND2_X1 U1441 ( .A1(n1818), .A2(n1819), .ZN(U301) );
NAND2_X1 U1442 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1625), .ZN(n1819) );
NAND2_X1 U1443 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1775), .ZN(n1818) );
NAND2_X1 U1444 ( .A1(n1820), .A2(n1821), .ZN(U300) );
NAND2_X1 U1445 ( .A1(n1822), .A2(n1775), .ZN(n1821) );
XOR2_X1 U1446 ( .A(REG3_REG_3__SCAN_IN), .B(KEYINPUT34), .Z(n1822) );
NAND2_X1 U1447 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1625), .ZN(n1820) );
NAND2_X1 U1448 ( .A1(n1823), .A2(n1824), .ZN(U299) );
NAND2_X1 U1449 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1625), .ZN(n1824) );
NAND2_X1 U1450 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1775), .ZN(n1823) );
NAND2_X1 U1451 ( .A1(n1825), .A2(n1826), .ZN(U298) );
NAND2_X1 U1452 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1625), .ZN(n1826) );
NAND2_X1 U1453 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1775), .ZN(n1825) );
NAND2_X1 U1454 ( .A1(n1827), .A2(n1828), .ZN(U297) );
NAND2_X1 U1455 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1625), .ZN(n1828) );
NAND2_X1 U1456 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1775), .ZN(n1827) );
NAND2_X1 U1457 ( .A1(n1829), .A2(n1830), .ZN(U296) );
NAND2_X1 U1458 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1625), .ZN(n1830) );
NAND2_X1 U1459 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1775), .ZN(n1829) );
NAND2_X1 U1460 ( .A1(n1831), .A2(n1832), .ZN(U295) );
NAND2_X1 U1461 ( .A1(n1833), .A2(n1775), .ZN(n1832) );
XNOR2_X1 U1462 ( .A(REG4_REG_6__SCAN_IN), .B(KEYINPUT55), .ZN(n1833) );
NAND2_X1 U1463 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1625), .ZN(n1831) );
NAND2_X1 U1464 ( .A1(n1834), .A2(n1835), .ZN(U294) );
NAND2_X1 U1465 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1625), .ZN(n1835) );
NAND2_X1 U1466 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1775), .ZN(n1834) );
NAND2_X1 U1467 ( .A1(n1836), .A2(n1837), .ZN(U293) );
NAND2_X1 U1468 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1625), .ZN(n1837) );
NAND2_X1 U1469 ( .A1(REG4_REG_4__SCAN_IN), .A2(n1775), .ZN(n1836) );
NAND2_X1 U1470 ( .A1(n1838), .A2(n1839), .ZN(U292) );
NAND2_X1 U1471 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1625), .ZN(n1839) );
XOR2_X1 U1472 ( .A(KEYINPUT32), .B(n1840), .Z(n1838) );
NOR2_X1 U1473 ( .A1(U280), .A2(n1841), .ZN(n1840) );
NAND2_X1 U1474 ( .A1(n1842), .A2(n1843), .ZN(U291) );
NAND2_X1 U1475 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1625), .ZN(n1843) );
NAND2_X1 U1476 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1775), .ZN(n1842) );
NAND2_X1 U1477 ( .A1(n1844), .A2(n1845), .ZN(U290) );
NAND2_X1 U1478 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1625), .ZN(n1845) );
NAND2_X1 U1479 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1775), .ZN(n1844) );
NAND2_X1 U1480 ( .A1(n1846), .A2(n1847), .ZN(U289) );
NAND2_X1 U1481 ( .A1(n1625), .A2(n1848), .ZN(n1847) );
XOR2_X1 U1482 ( .A(REG3_REG_0__SCAN_IN), .B(KEYINPUT41), .Z(n1848) );
NAND2_X1 U1483 ( .A1(n1849), .A2(REG4_REG_0__SCAN_IN), .ZN(n1846) );
XNOR2_X1 U1484 ( .A(n1775), .B(KEYINPUT61), .ZN(n1849) );
NAND4_X1 U1485 ( .A1(n1850), .A2(n1851), .A3(n1852), .A4(n1853), .ZN(U288));
NAND2_X1 U1486 ( .A1(n1854), .A2(n1855), .ZN(n1853) );
NAND2_X1 U1487 ( .A1(n1856), .A2(n1857), .ZN(n1855) );
NAND2_X1 U1488 ( .A1(n1858), .A2(n1859), .ZN(n1857) );
XNOR2_X1 U1489 ( .A(n1860), .B(KEYINPUT36), .ZN(n1858) );
NAND2_X1 U1490 ( .A1(n1861), .A2(RLAST_REG_7__SCAN_IN), .ZN(n1852) );
NAND2_X1 U1491 ( .A1(n1862), .A2(REG4_REG_7__SCAN_IN), .ZN(n1851) );
NAND2_X1 U1492 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1775), .ZN(n1850) );
NAND4_X1 U1493 ( .A1(n1863), .A2(n1864), .A3(n1865), .A4(n1866), .ZN(U287));
NOR3_X1 U1494 ( .A1(n1867), .A2(n1868), .A3(n1869), .ZN(n1866) );
NOR4_X1 U1495 ( .A1(n1870), .A2(n1871), .A3(n1872), .A4(n1873), .ZN(n1869));
AND2_X1 U1496 ( .A1(n1870), .A2(n1874), .ZN(n1868) );
NAND2_X1 U1497 ( .A1(KEYINPUT26), .A2(n1875), .ZN(n1870) );
XOR2_X1 U1498 ( .A(n1876), .B(KEYINPUT7), .Z(n1867) );
NAND2_X1 U1499 ( .A1(n1862), .A2(REG4_REG_6__SCAN_IN), .ZN(n1876) );
NAND2_X1 U1500 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n1775), .ZN(n1865) );
NAND2_X1 U1501 ( .A1(n1860), .A2(n1877), .ZN(n1864) );
XOR2_X1 U1502 ( .A(KEYINPUT10), .B(n1878), .Z(n1877) );
NOR2_X1 U1503 ( .A1(n1879), .A2(n1880), .ZN(n1878) );
XOR2_X1 U1504 ( .A(n1881), .B(n1882), .Z(n1880) );
NOR2_X1 U1505 ( .A1(n1872), .A2(n1859), .ZN(n1882) );
INV_X1 U1506 ( .A(n1883), .ZN(n1859) );
NAND2_X1 U1507 ( .A1(n1884), .A2(n1875), .ZN(n1881) );
NOR2_X1 U1508 ( .A1(n1875), .A2(n1884), .ZN(n1879) );
INV_X1 U1509 ( .A(KEYINPUT56), .ZN(n1884) );
NAND2_X1 U1510 ( .A1(n1861), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1863) );
NAND4_X1 U1511 ( .A1(n1885), .A2(n1886), .A3(n1887), .A4(n1888), .ZN(U286));
NOR3_X1 U1512 ( .A1(n1889), .A2(n1890), .A3(n1891), .ZN(n1888) );
AND2_X1 U1513 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1861), .ZN(n1891) );
NOR2_X1 U1514 ( .A1(n1892), .A2(n1893), .ZN(n1890) );
AND2_X1 U1515 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1862), .ZN(n1889) );
NAND2_X1 U1516 ( .A1(n1894), .A2(DATA_OUT_REG_5__SCAN_IN), .ZN(n1887) );
XNOR2_X1 U1517 ( .A(n1775), .B(KEYINPUT43), .ZN(n1894) );
NAND2_X1 U1518 ( .A1(n1874), .A2(n1895), .ZN(n1886) );
NAND2_X1 U1519 ( .A1(n1872), .A2(n1873), .ZN(n1895) );
INV_X1 U1520 ( .A(n1856), .ZN(n1874) );
NAND2_X1 U1521 ( .A1(n1896), .A2(n1897), .ZN(n1856) );
NAND2_X1 U1522 ( .A1(n1898), .A2(n1899), .ZN(n1897) );
NAND2_X1 U1523 ( .A1(n1900), .A2(n1860), .ZN(n1885) );
XNOR2_X1 U1524 ( .A(n1883), .B(n1872), .ZN(n1900) );
INV_X1 U1525 ( .A(n1899), .ZN(n1872) );
NAND2_X1 U1526 ( .A1(n1875), .A2(n1901), .ZN(n1899) );
NAND2_X1 U1527 ( .A1(n1902), .A2(n1903), .ZN(n1901) );
INV_X1 U1528 ( .A(n1854), .ZN(n1875) );
NOR2_X1 U1529 ( .A1(n1903), .A2(n1902), .ZN(n1854) );
INV_X1 U1530 ( .A(n1892), .ZN(n1902) );
NAND2_X1 U1531 ( .A1(n1904), .A2(n1905), .ZN(n1892) );
NAND4_X1 U1532 ( .A1(n1906), .A2(n1907), .A3(n1908), .A4(n1909), .ZN(n1905));
NAND2_X1 U1533 ( .A1(n1910), .A2(n1911), .ZN(n1909) );
XNOR2_X1 U1534 ( .A(n1912), .B(DATA_IN_6_), .ZN(n1910) );
NAND2_X1 U1535 ( .A1(n1913), .A2(RESTART), .ZN(n1908) );
XNOR2_X1 U1536 ( .A(RMIN_REG_6__SCAN_IN), .B(n1748), .ZN(n1913) );
INV_X1 U1537 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1748) );
NAND2_X1 U1538 ( .A1(n1914), .A2(n1915), .ZN(n1907) );
NAND2_X1 U1539 ( .A1(n1916), .A2(n1917), .ZN(n1915) );
XNOR2_X1 U1540 ( .A(n1918), .B(KEYINPUT38), .ZN(n1916) );
NAND4_X1 U1541 ( .A1(n1919), .A2(n1920), .A3(n1921), .A4(n1922), .ZN(n1904));
NAND2_X1 U1542 ( .A1(n1923), .A2(n1911), .ZN(n1922) );
XNOR2_X1 U1543 ( .A(REG4_REG_6__SCAN_IN), .B(DATA_IN_6_), .ZN(n1923) );
NAND2_X1 U1544 ( .A1(n1924), .A2(RESTART), .ZN(n1921) );
XNOR2_X1 U1545 ( .A(RMAX_REG_6__SCAN_IN), .B(RMIN_REG_6__SCAN_IN), .ZN(n1924) );
NAND2_X1 U1546 ( .A1(n1925), .A2(n1906), .ZN(n1920) );
NAND2_X1 U1547 ( .A1(n1926), .A2(n1918), .ZN(n1906) );
NAND2_X1 U1548 ( .A1(n1927), .A2(n1917), .ZN(n1919) );
NAND4_X1 U1549 ( .A1(n1928), .A2(n1929), .A3(n1930), .A4(n1931), .ZN(U285));
NOR3_X1 U1550 ( .A1(n1932), .A2(n1933), .A3(n1934), .ZN(n1931) );
NOR3_X1 U1551 ( .A1(n1871), .A2(n1898), .A3(n1935), .ZN(n1934) );
NOR2_X1 U1552 ( .A1(n1936), .A2(n1937), .ZN(n1935) );
NOR2_X1 U1553 ( .A1(n1938), .A2(n1939), .ZN(n1936) );
INV_X1 U1554 ( .A(n1873), .ZN(n1898) );
NAND3_X1 U1555 ( .A1(n1940), .A2(n1941), .A3(n1942), .ZN(n1873) );
XOR2_X1 U1556 ( .A(n1937), .B(KEYINPUT24), .Z(n1942) );
NOR3_X1 U1557 ( .A1(n1943), .A2(n1883), .A3(n1944), .ZN(n1933) );
NOR2_X1 U1558 ( .A1(n1945), .A2(n1937), .ZN(n1944) );
NOR2_X1 U1559 ( .A1(n1946), .A2(n1947), .ZN(n1945) );
NOR3_X1 U1560 ( .A1(n1946), .A2(n1948), .A3(n1947), .ZN(n1883) );
INV_X1 U1561 ( .A(n1937), .ZN(n1948) );
NAND2_X1 U1562 ( .A1(n1903), .A2(n1949), .ZN(n1937) );
NAND2_X1 U1563 ( .A1(n1950), .A2(n1951), .ZN(n1949) );
OR2_X1 U1564 ( .A1(n1951), .A2(n1950), .ZN(n1903) );
AND2_X1 U1565 ( .A1(n1950), .A2(n1952), .ZN(n1932) );
NAND2_X1 U1566 ( .A1(n1953), .A2(n1954), .ZN(n1950) );
NAND2_X1 U1567 ( .A1(n1955), .A2(n1917), .ZN(n1954) );
XNOR2_X1 U1568 ( .A(n1956), .B(n1925), .ZN(n1955) );
XNOR2_X1 U1569 ( .A(KEYINPUT6), .B(n1957), .ZN(n1956) );
NOR2_X1 U1570 ( .A1(KEYINPUT31), .A2(n1918), .ZN(n1957) );
INV_X1 U1571 ( .A(n1927), .ZN(n1918) );
NAND2_X1 U1572 ( .A1(n1958), .A2(n1926), .ZN(n1953) );
INV_X1 U1573 ( .A(n1917), .ZN(n1926) );
NAND2_X1 U1574 ( .A1(n1959), .A2(n1960), .ZN(n1917) );
NAND2_X1 U1575 ( .A1(n1961), .A2(n1962), .ZN(n1960) );
OR2_X1 U1576 ( .A1(n1963), .A2(n1964), .ZN(n1961) );
NAND2_X1 U1577 ( .A1(n1964), .A2(n1963), .ZN(n1959) );
XNOR2_X1 U1578 ( .A(n1914), .B(n1965), .ZN(n1958) );
NOR2_X1 U1579 ( .A1(KEYINPUT44), .A2(n1927), .ZN(n1965) );
NAND2_X1 U1580 ( .A1(n1966), .A2(n1967), .ZN(n1927) );
NAND2_X1 U1581 ( .A1(RESTART), .A2(n1726), .ZN(n1967) );
NAND2_X1 U1582 ( .A1(n1687), .A2(n1911), .ZN(n1966) );
INV_X1 U1583 ( .A(n1925), .ZN(n1914) );
NAND2_X1 U1584 ( .A1(n1968), .A2(n1969), .ZN(n1925) );
NAND2_X1 U1585 ( .A1(RESTART), .A2(n1691), .ZN(n1969) );
NAND2_X1 U1586 ( .A1(n1970), .A2(n1911), .ZN(n1968) );
NAND2_X1 U1587 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1775), .ZN(n1930) );
NAND2_X1 U1588 ( .A1(n1861), .A2(RLAST_REG_4__SCAN_IN), .ZN(n1929) );
NAND2_X1 U1589 ( .A1(n1862), .A2(REG4_REG_4__SCAN_IN), .ZN(n1928) );
NAND4_X1 U1590 ( .A1(n1971), .A2(n1972), .A3(n1973), .A4(n1974), .ZN(U284));
AND4_X1 U1591 ( .A1(n1975), .A2(n1976), .A3(n1977), .A4(n1978), .ZN(n1974));
NAND2_X1 U1592 ( .A1(n1979), .A2(n1941), .ZN(n1978) );
NAND3_X1 U1593 ( .A1(n1896), .A2(n1940), .A3(n1938), .ZN(n1977) );
NAND2_X1 U1594 ( .A1(n1862), .A2(REG4_REG_3__SCAN_IN), .ZN(n1976) );
NAND2_X1 U1595 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1775), .ZN(n1975) );
NAND2_X1 U1596 ( .A1(n1861), .A2(RLAST_REG_3__SCAN_IN), .ZN(n1973) );
NAND3_X1 U1597 ( .A1(n1980), .A2(n1946), .A3(n1860), .ZN(n1972) );
XOR2_X1 U1598 ( .A(n1938), .B(KEYINPUT4), .Z(n1946) );
INV_X1 U1599 ( .A(n1941), .ZN(n1938) );
NAND2_X1 U1600 ( .A1(n1981), .A2(n1951), .ZN(n1941) );
OR2_X1 U1601 ( .A1(n1982), .A2(n1983), .ZN(n1951) );
NAND2_X1 U1602 ( .A1(n1983), .A2(n1982), .ZN(n1981) );
INV_X1 U1603 ( .A(n1947), .ZN(n1980) );
NAND2_X1 U1604 ( .A1(n1952), .A2(n1983), .ZN(n1971) );
NAND2_X1 U1605 ( .A1(n1984), .A2(n1985), .ZN(n1983) );
NAND2_X1 U1606 ( .A1(n1986), .A2(n1962), .ZN(n1985) );
XOR2_X1 U1607 ( .A(n1987), .B(KEYINPUT1), .Z(n1984) );
OR2_X1 U1608 ( .A1(n1962), .A2(n1986), .ZN(n1987) );
XOR2_X1 U1609 ( .A(n1988), .B(n1963), .Z(n1986) );
NAND2_X1 U1610 ( .A1(n1989), .A2(n1990), .ZN(n1963) );
NAND2_X1 U1611 ( .A1(RESTART), .A2(n1745), .ZN(n1990) );
NAND2_X1 U1612 ( .A1(n1695), .A2(n1911), .ZN(n1989) );
INV_X1 U1613 ( .A(DATA_IN_4_), .ZN(n1695) );
NAND2_X1 U1614 ( .A1(KEYINPUT25), .A2(n1991), .ZN(n1988) );
INV_X1 U1615 ( .A(n1964), .ZN(n1991) );
NAND2_X1 U1616 ( .A1(n1992), .A2(n1993), .ZN(n1964) );
NAND2_X1 U1617 ( .A1(RESTART), .A2(n1712), .ZN(n1993) );
OR2_X1 U1618 ( .A1(REG4_REG_4__SCAN_IN), .A2(RESTART), .ZN(n1992) );
NAND2_X1 U1619 ( .A1(n1994), .A2(n1995), .ZN(n1962) );
NAND2_X1 U1620 ( .A1(n1996), .A2(n1997), .ZN(n1995) );
NAND2_X1 U1621 ( .A1(n1998), .A2(n1999), .ZN(n1997) );
NAND2_X1 U1622 ( .A1(n2000), .A2(n2001), .ZN(n1994) );
NAND4_X1 U1623 ( .A1(n2002), .A2(n2003), .A3(n2004), .A4(n2005), .ZN(U283));
NOR4_X1 U1624 ( .A1(n2006), .A2(n2007), .A3(n2008), .A4(n2009), .ZN(n2005));
AND2_X1 U1625 ( .A1(n2010), .A2(n1952), .ZN(n2009) );
INV_X1 U1626 ( .A(n1893), .ZN(n1952) );
AND2_X1 U1627 ( .A1(n2011), .A2(n1979), .ZN(n2008) );
NAND2_X1 U1628 ( .A1(n2012), .A2(n2013), .ZN(n1979) );
NAND2_X1 U1629 ( .A1(n1860), .A2(n1947), .ZN(n2013) );
NAND2_X1 U1630 ( .A1(n1896), .A2(n1939), .ZN(n2012) );
AND4_X1 U1631 ( .A1(n2014), .A2(n1947), .A3(n2015), .A4(n1860), .ZN(n2007));
NAND3_X1 U1632 ( .A1(n2015), .A2(n2014), .A3(n2011), .ZN(n1947) );
NOR4_X1 U1633 ( .A1(n2016), .A2(n1940), .A3(n1871), .A4(n2017), .ZN(n2006));
XNOR2_X1 U1634 ( .A(KEYINPUT23), .B(n2015), .ZN(n2017) );
INV_X1 U1635 ( .A(n1939), .ZN(n1940) );
NAND3_X1 U1636 ( .A1(n2011), .A2(n2018), .A3(n2019), .ZN(n1939) );
XNOR2_X1 U1637 ( .A(KEYINPUT37), .B(n2015), .ZN(n2019) );
NAND2_X1 U1638 ( .A1(n1982), .A2(n2020), .ZN(n2011) );
NAND2_X1 U1639 ( .A1(n2021), .A2(n2010), .ZN(n2020) );
OR2_X1 U1640 ( .A1(n2010), .A2(n2021), .ZN(n1982) );
NAND3_X1 U1641 ( .A1(n2022), .A2(n2023), .A3(n2024), .ZN(n2010) );
NAND3_X1 U1642 ( .A1(n2025), .A2(n1999), .A3(n1998), .ZN(n2024) );
NAND2_X1 U1643 ( .A1(KEYINPUT20), .A2(n1996), .ZN(n2025) );
OR4_X1 U1644 ( .A1(n1998), .A2(KEYINPUT51), .A3(n1999), .A4(n1996), .ZN(n2023) );
NAND2_X1 U1645 ( .A1(n2026), .A2(n1996), .ZN(n2022) );
NAND2_X1 U1646 ( .A1(n2027), .A2(n2028), .ZN(n1996) );
NAND2_X1 U1647 ( .A1(RESTART), .A2(n1710), .ZN(n2028) );
NAND2_X1 U1648 ( .A1(n1841), .A2(n1911), .ZN(n2027) );
NAND2_X1 U1649 ( .A1(n2029), .A2(n2030), .ZN(n2026) );
NAND2_X1 U1650 ( .A1(n2031), .A2(n2000), .ZN(n2030) );
INV_X1 U1651 ( .A(n1999), .ZN(n2000) );
OR2_X1 U1652 ( .A1(n1998), .A2(KEYINPUT51), .ZN(n2031) );
INV_X1 U1653 ( .A(n2001), .ZN(n1998) );
NAND3_X1 U1654 ( .A1(KEYINPUT20), .A2(n2001), .A3(n1999), .ZN(n2029) );
NAND2_X1 U1655 ( .A1(n2032), .A2(n2033), .ZN(n1999) );
NAND2_X1 U1656 ( .A1(n2034), .A2(n2035), .ZN(n2033) );
NAND2_X1 U1657 ( .A1(n2036), .A2(n2037), .ZN(n2034) );
XOR2_X1 U1658 ( .A(KEYINPUT42), .B(n2038), .Z(n2032) );
NOR2_X1 U1659 ( .A1(n2036), .A2(n2037), .ZN(n2038) );
NAND2_X1 U1660 ( .A1(n2039), .A2(n2040), .ZN(n2001) );
NAND2_X1 U1661 ( .A1(RESTART), .A2(n1733), .ZN(n2040) );
NAND2_X1 U1662 ( .A1(n1711), .A2(n1911), .ZN(n2039) );
NAND2_X1 U1663 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1775), .ZN(n2004) );
NAND2_X1 U1664 ( .A1(n1861), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2003) );
NAND2_X1 U1665 ( .A1(n1862), .A2(REG4_REG_2__SCAN_IN), .ZN(n2002) );
NAND4_X1 U1666 ( .A1(n2041), .A2(n2042), .A3(n2043), .A4(n2044), .ZN(U282));
NOR3_X1 U1667 ( .A1(n2045), .A2(n2046), .A3(n2047), .ZN(n2044) );
NOR2_X1 U1668 ( .A1(n2048), .A2(n1943), .ZN(n2047) );
INV_X1 U1669 ( .A(n1860), .ZN(n1943) );
XNOR2_X1 U1670 ( .A(n2014), .B(n2015), .ZN(n2048) );
NAND2_X1 U1671 ( .A1(n2049), .A2(n2021), .ZN(n2014) );
NAND2_X1 U1672 ( .A1(n2050), .A2(n2051), .ZN(n2049) );
XNOR2_X1 U1673 ( .A(n2052), .B(KEYINPUT53), .ZN(n2050) );
NOR2_X1 U1674 ( .A1(n2052), .A2(n2053), .ZN(n2046) );
XNOR2_X1 U1675 ( .A(KEYINPUT49), .B(n1893), .ZN(n2053) );
NOR2_X1 U1676 ( .A1(n2054), .A2(n1871), .ZN(n2045) );
INV_X1 U1677 ( .A(n1896), .ZN(n1871) );
NOR2_X1 U1678 ( .A1(n2055), .A2(n2056), .ZN(n2054) );
XOR2_X1 U1679 ( .A(n2057), .B(KEYINPUT0), .Z(n2056) );
NAND2_X1 U1680 ( .A1(n2016), .A2(n2015), .ZN(n2057) );
NOR2_X1 U1681 ( .A1(n2016), .A2(n2015), .ZN(n2055) );
INV_X1 U1682 ( .A(n2018), .ZN(n2016) );
NAND2_X1 U1683 ( .A1(n2021), .A2(n2058), .ZN(n2018) );
NAND2_X1 U1684 ( .A1(n2059), .A2(n2051), .ZN(n2058) );
OR2_X1 U1685 ( .A1(n2051), .A2(n2059), .ZN(n2021) );
INV_X1 U1686 ( .A(n2052), .ZN(n2059) );
XOR2_X1 U1687 ( .A(n2060), .B(n2035), .Z(n2052) );
NAND2_X1 U1688 ( .A1(n2061), .A2(n2062), .ZN(n2035) );
NAND2_X1 U1689 ( .A1(n2063), .A2(n2064), .ZN(n2062) );
NAND2_X1 U1690 ( .A1(n2065), .A2(n2066), .ZN(n2064) );
XOR2_X1 U1691 ( .A(n2067), .B(KEYINPUT63), .Z(n2065) );
OR2_X1 U1692 ( .A1(n2066), .A2(n2067), .ZN(n2061) );
NAND2_X1 U1693 ( .A1(KEYINPUT14), .A2(n2068), .ZN(n2060) );
XOR2_X1 U1694 ( .A(n2037), .B(n2036), .Z(n2068) );
NAND2_X1 U1695 ( .A1(n2069), .A2(n2070), .ZN(n2036) );
NAND2_X1 U1696 ( .A1(RESTART), .A2(n1699), .ZN(n2070) );
NAND2_X1 U1697 ( .A1(n2071), .A2(n1911), .ZN(n2069) );
NAND2_X1 U1698 ( .A1(n2072), .A2(n2073), .ZN(n2037) );
NAND2_X1 U1699 ( .A1(RESTART), .A2(n1740), .ZN(n2073) );
NAND2_X1 U1700 ( .A1(n1703), .A2(n1911), .ZN(n2072) );
NAND2_X1 U1701 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1775), .ZN(n2043) );
NAND2_X1 U1702 ( .A1(n1861), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2042) );
NAND2_X1 U1703 ( .A1(n1862), .A2(REG4_REG_1__SCAN_IN), .ZN(n2041) );
NAND3_X1 U1704 ( .A1(n2074), .A2(n2075), .A3(n2076), .ZN(U281) );
NOR3_X1 U1705 ( .A1(n2077), .A2(n2078), .A3(n2079), .ZN(n2076) );
AND2_X1 U1706 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1861), .ZN(n2079) );
NOR2_X1 U1707 ( .A1(n2080), .A2(ENABLE), .ZN(n1861) );
NOR2_X1 U1708 ( .A1(n2081), .A2(n2015), .ZN(n2078) );
NAND2_X1 U1709 ( .A1(n2051), .A2(n2082), .ZN(n2015) );
NAND3_X1 U1710 ( .A1(n2083), .A2(n2067), .A3(n2084), .ZN(n2082) );
NAND2_X1 U1711 ( .A1(n2085), .A2(n2086), .ZN(n2051) );
NAND2_X1 U1712 ( .A1(n2083), .A2(n2067), .ZN(n2086) );
NAND3_X1 U1713 ( .A1(n2087), .A2(n2088), .A3(n2089), .ZN(n2083) );
NAND2_X1 U1714 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1911), .ZN(n2088) );
NAND2_X1 U1715 ( .A1(RESTART), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2087) );
NOR2_X1 U1716 ( .A1(n1860), .A2(n1896), .ZN(n2081) );
NOR3_X1 U1717 ( .A1(n1772), .A2(n1775), .A3(n2090), .ZN(n1896) );
NOR2_X1 U1718 ( .A1(n2085), .A2(n1893), .ZN(n2077) );
NAND4_X1 U1719 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2092), .A3(n2090), .A4(U280), .ZN(n1893) );
NAND3_X1 U1720 ( .A1(n2093), .A2(n2094), .A3(RESTART), .ZN(n2090) );
NAND2_X1 U1721 ( .A1(n2095), .A2(n2096), .ZN(n2094) );
NAND2_X1 U1722 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2096) );
NAND2_X1 U1723 ( .A1(n2097), .A2(n2098), .ZN(n2095) );
NAND2_X1 U1724 ( .A1(RMIN_REG_6__SCAN_IN), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2098) );
NAND3_X1 U1725 ( .A1(n2099), .A2(n2100), .A3(n2101), .ZN(n2097) );
OR2_X1 U1726 ( .A1(RMAX_REG_6__SCAN_IN), .A2(RMIN_REG_6__SCAN_IN), .ZN(n2101) );
NAND3_X1 U1727 ( .A1(n2102), .A2(n2103), .A3(n2104), .ZN(n2100) );
NAND2_X1 U1728 ( .A1(n2105), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2104) );
XNOR2_X1 U1729 ( .A(RMAX_REG_5__SCAN_IN), .B(KEYINPUT17), .ZN(n2105) );
NAND3_X1 U1730 ( .A1(n2106), .A2(n2107), .A3(n2108), .ZN(n2103) );
NAND2_X1 U1731 ( .A1(n1745), .A2(n1712), .ZN(n2108) );
INV_X1 U1732 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1712) );
NAND3_X1 U1733 ( .A1(n2109), .A2(n2110), .A3(n2111), .ZN(n2107) );
NAND2_X1 U1734 ( .A1(RMIN_REG_2__SCAN_IN), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2111) );
NAND3_X1 U1735 ( .A1(n2112), .A2(n2113), .A3(n2114), .ZN(n2110) );
NAND2_X1 U1736 ( .A1(n1740), .A2(n1699), .ZN(n2114) );
INV_X1 U1737 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1699) );
INV_X1 U1738 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1740) );
NAND2_X1 U1739 ( .A1(n2115), .A2(n2116), .ZN(n2113) );
OR2_X1 U1740 ( .A1(n2117), .A2(n1743), .ZN(n2115) );
NAND2_X1 U1741 ( .A1(n2117), .A2(n1743), .ZN(n2112) );
NAND2_X1 U1742 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2117) );
NAND2_X1 U1743 ( .A1(n2118), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2109) );
XNOR2_X1 U1744 ( .A(RMIN_REG_3__SCAN_IN), .B(KEYINPUT21), .ZN(n2118) );
NAND2_X1 U1745 ( .A1(n1733), .A2(n1710), .ZN(n2106) );
INV_X1 U1746 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1710) );
INV_X1 U1747 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1733) );
NAND2_X1 U1748 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n2119), .ZN(n2102) );
XNOR2_X1 U1749 ( .A(n1745), .B(KEYINPUT58), .ZN(n2119) );
INV_X1 U1750 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1745) );
NAND2_X1 U1751 ( .A1(n1726), .A2(n1691), .ZN(n2099) );
INV_X1 U1752 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1691) );
INV_X1 U1753 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1726) );
NAND2_X1 U1754 ( .A1(n1631), .A2(n1716), .ZN(n2093) );
INV_X1 U1755 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1716) );
INV_X1 U1756 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1631) );
NAND2_X1 U1757 ( .A1(n2120), .A2(n1911), .ZN(n2092) );
NAND3_X1 U1758 ( .A1(n2091), .A2(n2121), .A3(ENABLE), .ZN(n2120) );
NAND2_X1 U1759 ( .A1(n2122), .A2(n2123), .ZN(n2091) );
NAND2_X1 U1760 ( .A1(n2124), .A2(n2125), .ZN(n2123) );
NAND2_X1 U1761 ( .A1(REG4_REG_7__SCAN_IN), .A2(DATA_IN_7_), .ZN(n2125) );
NAND2_X1 U1762 ( .A1(n2126), .A2(n2127), .ZN(n2124) );
NAND2_X1 U1763 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2127) );
NAND3_X1 U1764 ( .A1(n2128), .A2(n2129), .A3(n2130), .ZN(n2126) );
NAND2_X1 U1765 ( .A1(n1714), .A2(n1912), .ZN(n2130) );
INV_X1 U1766 ( .A(REG4_REG_6__SCAN_IN), .ZN(n1912) );
INV_X1 U1767 ( .A(DATA_IN_6_), .ZN(n1714) );
NAND3_X1 U1768 ( .A1(n2131), .A2(n2132), .A3(n2133), .ZN(n2129) );
XOR2_X1 U1769 ( .A(KEYINPUT57), .B(n2134), .Z(n2133) );
NOR2_X1 U1770 ( .A1(n2135), .A2(n2136), .ZN(n2134) );
XOR2_X1 U1771 ( .A(KEYINPUT13), .B(n2137), .Z(n2136) );
NOR2_X1 U1772 ( .A1(DATA_IN_4_), .A2(REG4_REG_4__SCAN_IN), .ZN(n2137) );
NOR2_X1 U1773 ( .A1(n2138), .A2(n2139), .ZN(n2135) );
NOR2_X1 U1774 ( .A1(n1711), .A2(n1841), .ZN(n2139) );
INV_X1 U1775 ( .A(REG4_REG_3__SCAN_IN), .ZN(n1841) );
INV_X1 U1776 ( .A(DATA_IN_3_), .ZN(n1711) );
NOR2_X1 U1777 ( .A1(n2140), .A2(n2141), .ZN(n2138) );
NOR2_X1 U1778 ( .A1(n2142), .A2(n2143), .ZN(n2141) );
NOR2_X1 U1779 ( .A1(n1703), .A2(n2071), .ZN(n2143) );
INV_X1 U1780 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2071) );
INV_X1 U1781 ( .A(DATA_IN_2_), .ZN(n1703) );
NOR3_X1 U1782 ( .A1(n2144), .A2(n2145), .A3(n2146), .ZN(n2142) );
NOR2_X1 U1783 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2146) );
NOR2_X1 U1784 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2145) );
NOR2_X1 U1785 ( .A1(n2147), .A2(n2148), .ZN(n2144) );
AND2_X1 U1786 ( .A1(DATA_IN_1_), .A2(REG4_REG_1__SCAN_IN), .ZN(n2148) );
NOR2_X1 U1787 ( .A1(n1705), .A2(n2149), .ZN(n2147) );
NOR2_X1 U1788 ( .A1(DATA_IN_3_), .A2(REG4_REG_3__SCAN_IN), .ZN(n2140) );
NAND2_X1 U1789 ( .A1(REG4_REG_5__SCAN_IN), .A2(n2150), .ZN(n2132) );
XNOR2_X1 U1790 ( .A(KEYINPUT54), .B(n1687), .ZN(n2150) );
NAND2_X1 U1791 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2131) );
NAND2_X1 U1792 ( .A1(n1687), .A2(n1970), .ZN(n2128) );
INV_X1 U1793 ( .A(REG4_REG_5__SCAN_IN), .ZN(n1970) );
INV_X1 U1794 ( .A(DATA_IN_5_), .ZN(n1687) );
OR2_X1 U1795 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2122) );
INV_X1 U1796 ( .A(n2084), .ZN(n2085) );
XNOR2_X1 U1797 ( .A(n2151), .B(n2063), .ZN(n2084) );
AND2_X1 U1798 ( .A1(n2152), .A2(n2153), .ZN(n2063) );
NAND2_X1 U1799 ( .A1(RESTART), .A2(n2116), .ZN(n2153) );
INV_X1 U1800 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n2116) );
NAND2_X1 U1801 ( .A1(n2154), .A2(n1911), .ZN(n2152) );
XNOR2_X1 U1802 ( .A(REG4_REG_1__SCAN_IN), .B(KEYINPUT22), .ZN(n2154) );
XNOR2_X1 U1803 ( .A(n2067), .B(n2066), .ZN(n2151) );
NAND2_X1 U1804 ( .A1(n2155), .A2(n2156), .ZN(n2066) );
NAND2_X1 U1805 ( .A1(RESTART), .A2(n1743), .ZN(n2156) );
INV_X1 U1806 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1743) );
NAND2_X1 U1807 ( .A1(n1708), .A2(n1911), .ZN(n2155) );
INV_X1 U1808 ( .A(DATA_IN_1_), .ZN(n1708) );
NAND3_X1 U1809 ( .A1(n2157), .A2(n2158), .A3(n2159), .ZN(n2067) );
INV_X1 U1810 ( .A(n2089), .ZN(n2159) );
NAND3_X1 U1811 ( .A1(n2160), .A2(n2161), .A3(n2162), .ZN(n2089) );
NAND2_X1 U1812 ( .A1(n2163), .A2(n1742), .ZN(n2162) );
INV_X1 U1813 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1742) );
NAND2_X1 U1814 ( .A1(DATA_IN_0_), .A2(n1911), .ZN(n2163) );
NAND3_X1 U1815 ( .A1(KEYINPUT46), .A2(n1705), .A3(n1911), .ZN(n2161) );
INV_X1 U1816 ( .A(DATA_IN_0_), .ZN(n1705) );
OR2_X1 U1817 ( .A1(n1911), .A2(KEYINPUT46), .ZN(n2160) );
OR2_X1 U1818 ( .A1(n1911), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2158) );
NAND2_X1 U1819 ( .A1(n2149), .A2(n1911), .ZN(n2157) );
INV_X1 U1820 ( .A(REG4_REG_0__SCAN_IN), .ZN(n2149) );
NAND2_X1 U1821 ( .A1(n1862), .A2(REG4_REG_0__SCAN_IN), .ZN(n2075) );
NOR3_X1 U1822 ( .A1(n1771), .A2(n2080), .A3(n2121), .ZN(n1862) );
INV_X1 U1823 ( .A(AVERAGE), .ZN(n2121) );
NAND3_X1 U1824 ( .A1(U280), .A2(n1911), .A3(STATO_REG_1__SCAN_IN), .ZN(n2080) );
INV_X1 U1825 ( .A(RESTART), .ZN(n1911) );
INV_X1 U1826 ( .A(ENABLE), .ZN(n1771) );
NAND2_X1 U1827 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1775), .ZN(n2074) );
NAND2_X1 U1828 ( .A1(n1624), .A2(n2164), .ZN(U280) );
NAND2_X1 U1829 ( .A1(STATO_REG_0__SCAN_IN), .A2(n1772), .ZN(n2164) );
INV_X1 U1830 ( .A(STATO_REG_1__SCAN_IN), .ZN(n1772) );
endmodule


