//Key = 1111000000000101010001100100001110010000101010011111000000111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404;

XNOR2_X1 U782 ( .A(G107), .B(n1074), .ZN(G9) );
NAND2_X1 U783 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U784 ( .A1(n1077), .A2(n1078), .ZN(G75) );
XOR2_X1 U785 ( .A(KEYINPUT16), .B(n1079), .Z(n1078) );
NOR3_X1 U786 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U787 ( .A1(n1083), .A2(n1084), .ZN(n1081) );
NOR2_X1 U788 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR3_X1 U789 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NOR2_X1 U790 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U791 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U792 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U794 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NOR2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(n1094) );
NOR2_X1 U796 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U797 ( .A1(n1104), .A2(n1105), .ZN(n1102) );
NOR3_X1 U798 ( .A1(n1097), .A2(n1106), .A3(n1101), .ZN(n1090) );
NOR4_X1 U799 ( .A1(n1107), .A2(n1101), .A3(n1097), .A4(n1093), .ZN(n1085) );
INV_X1 U800 ( .A(n1108), .ZN(n1093) );
INV_X1 U801 ( .A(n1109), .ZN(n1097) );
NOR2_X1 U802 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
NOR2_X1 U803 ( .A1(n1089), .A2(n1112), .ZN(n1110) );
NOR2_X1 U804 ( .A1(G952), .A2(n1082), .ZN(n1077) );
NAND2_X1 U805 ( .A1(n1113), .A2(n1114), .ZN(n1082) );
NAND4_X1 U806 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .ZN(n1114) );
NOR4_X1 U807 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
INV_X1 U808 ( .A(n1112), .ZN(n1122) );
NAND2_X1 U809 ( .A1(n1123), .A2(n1124), .ZN(n1119) );
NOR3_X1 U810 ( .A1(n1125), .A2(n1126), .A3(n1089), .ZN(n1117) );
XOR2_X1 U811 ( .A(n1127), .B(KEYINPUT32), .Z(n1126) );
XOR2_X1 U812 ( .A(n1128), .B(n1129), .Z(n1125) );
XOR2_X1 U813 ( .A(n1130), .B(KEYINPUT13), .Z(n1129) );
NAND2_X1 U814 ( .A1(KEYINPUT2), .A2(n1131), .ZN(n1128) );
XOR2_X1 U815 ( .A(n1132), .B(G475), .Z(n1116) );
NAND2_X1 U816 ( .A1(KEYINPUT42), .A2(n1133), .ZN(n1132) );
XOR2_X1 U817 ( .A(n1134), .B(G478), .Z(n1115) );
NAND2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(G72) );
NAND2_X1 U819 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U820 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
NAND2_X1 U821 ( .A1(n1141), .A2(n1140), .ZN(n1135) );
NAND2_X1 U822 ( .A1(G953), .A2(n1142), .ZN(n1140) );
INV_X1 U823 ( .A(G227), .ZN(n1142) );
INV_X1 U824 ( .A(n1138), .ZN(n1141) );
NAND2_X1 U825 ( .A1(KEYINPUT0), .A2(n1143), .ZN(n1138) );
XOR2_X1 U826 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND2_X1 U827 ( .A1(n1113), .A2(n1146), .ZN(n1145) );
NAND2_X1 U828 ( .A1(n1147), .A2(n1139), .ZN(n1144) );
INV_X1 U829 ( .A(n1148), .ZN(n1139) );
XOR2_X1 U830 ( .A(n1149), .B(n1150), .Z(n1147) );
XOR2_X1 U831 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U832 ( .A(n1153), .B(G137), .Z(n1152) );
NAND2_X1 U833 ( .A1(KEYINPUT47), .A2(n1154), .ZN(n1151) );
XOR2_X1 U834 ( .A(n1155), .B(n1156), .Z(n1149) );
XOR2_X1 U835 ( .A(n1157), .B(n1158), .Z(n1155) );
XOR2_X1 U836 ( .A(n1159), .B(n1160), .Z(G69) );
XOR2_X1 U837 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U838 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XOR2_X1 U839 ( .A(KEYINPUT9), .B(G953), .Z(n1164) );
NOR2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
XOR2_X1 U841 ( .A(n1167), .B(KEYINPUT14), .Z(n1165) );
NAND2_X1 U842 ( .A1(n1168), .A2(n1169), .ZN(n1161) );
NAND2_X1 U843 ( .A1(G953), .A2(n1170), .ZN(n1169) );
XOR2_X1 U844 ( .A(KEYINPUT31), .B(G898), .Z(n1170) );
XOR2_X1 U845 ( .A(n1171), .B(n1172), .Z(n1168) );
XOR2_X1 U846 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U847 ( .A(n1175), .B(n1176), .Z(n1171) );
NOR2_X1 U848 ( .A1(KEYINPUT53), .A2(n1177), .ZN(n1176) );
INV_X1 U849 ( .A(n1178), .ZN(n1177) );
XNOR2_X1 U850 ( .A(KEYINPUT19), .B(KEYINPUT12), .ZN(n1175) );
NAND2_X1 U851 ( .A1(G953), .A2(n1179), .ZN(n1159) );
NAND2_X1 U852 ( .A1(G898), .A2(G224), .ZN(n1179) );
NOR3_X1 U853 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(G66) );
NOR3_X1 U854 ( .A1(n1183), .A2(G953), .A3(G952), .ZN(n1182) );
INV_X1 U855 ( .A(KEYINPUT5), .ZN(n1183) );
NOR2_X1 U856 ( .A1(KEYINPUT5), .A2(n1184), .ZN(n1181) );
XNOR2_X1 U857 ( .A(n1185), .B(n1186), .ZN(n1180) );
NOR2_X1 U858 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NOR2_X1 U859 ( .A1(n1189), .A2(n1190), .ZN(G63) );
XOR2_X1 U860 ( .A(n1191), .B(n1192), .Z(n1190) );
NOR2_X1 U861 ( .A1(n1193), .A2(n1188), .ZN(n1191) );
NOR2_X1 U862 ( .A1(n1189), .A2(n1194), .ZN(G60) );
NOR3_X1 U863 ( .A1(n1195), .A2(n1133), .A3(n1196), .ZN(n1194) );
NOR2_X1 U864 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NOR2_X1 U865 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
XOR2_X1 U866 ( .A(KEYINPUT54), .B(n1201), .Z(n1195) );
NOR3_X1 U867 ( .A1(n1202), .A2(n1200), .A3(n1188), .ZN(n1201) );
XNOR2_X1 U868 ( .A(G104), .B(n1203), .ZN(G6) );
NOR2_X1 U869 ( .A1(n1189), .A2(n1204), .ZN(G57) );
XOR2_X1 U870 ( .A(n1205), .B(n1206), .Z(n1204) );
XNOR2_X1 U871 ( .A(G101), .B(n1207), .ZN(n1206) );
XNOR2_X1 U872 ( .A(n1208), .B(n1209), .ZN(n1205) );
NOR2_X1 U873 ( .A1(n1130), .A2(n1188), .ZN(n1209) );
INV_X1 U874 ( .A(G472), .ZN(n1130) );
NOR3_X1 U875 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(G54) );
NOR3_X1 U876 ( .A1(n1213), .A2(G953), .A3(G952), .ZN(n1212) );
INV_X1 U877 ( .A(KEYINPUT11), .ZN(n1213) );
NOR2_X1 U878 ( .A1(KEYINPUT11), .A2(n1184), .ZN(n1211) );
INV_X1 U879 ( .A(n1189), .ZN(n1184) );
XOR2_X1 U880 ( .A(n1214), .B(n1215), .Z(n1210) );
NOR2_X1 U881 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
AND3_X1 U882 ( .A1(KEYINPUT52), .A2(n1218), .A3(G140), .ZN(n1217) );
NOR2_X1 U883 ( .A1(KEYINPUT52), .A2(n1219), .ZN(n1216) );
XOR2_X1 U884 ( .A(n1220), .B(n1221), .Z(n1214) );
NOR2_X1 U885 ( .A1(n1222), .A2(n1188), .ZN(n1221) );
INV_X1 U886 ( .A(G469), .ZN(n1222) );
NOR2_X1 U887 ( .A1(n1189), .A2(n1223), .ZN(G51) );
XOR2_X1 U888 ( .A(n1224), .B(n1225), .Z(n1223) );
XOR2_X1 U889 ( .A(n1226), .B(n1227), .Z(n1225) );
NOR2_X1 U890 ( .A1(n1228), .A2(n1188), .ZN(n1227) );
NAND2_X1 U891 ( .A1(G902), .A2(n1080), .ZN(n1188) );
INV_X1 U892 ( .A(n1199), .ZN(n1080) );
NOR3_X1 U893 ( .A1(n1167), .A2(n1166), .A3(n1146), .ZN(n1199) );
NAND4_X1 U894 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1146) );
NOR4_X1 U895 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1232) );
INV_X1 U896 ( .A(n1237), .ZN(n1235) );
NOR3_X1 U897 ( .A1(n1111), .A2(KEYINPUT60), .A3(n1238), .ZN(n1234) );
NOR2_X1 U898 ( .A1(n1239), .A2(n1240), .ZN(n1233) );
NOR2_X1 U899 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
NOR2_X1 U900 ( .A1(n1238), .A2(n1243), .ZN(n1242) );
INV_X1 U901 ( .A(KEYINPUT60), .ZN(n1243) );
NOR3_X1 U902 ( .A1(n1244), .A2(n1106), .A3(n1245), .ZN(n1241) );
NOR2_X1 U903 ( .A1(n1246), .A2(n1075), .ZN(n1106) );
NAND4_X1 U904 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1166) );
NAND4_X1 U905 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1109), .ZN(n1247) );
XOR2_X1 U906 ( .A(n1240), .B(KEYINPUT40), .Z(n1252) );
XOR2_X1 U907 ( .A(n1254), .B(KEYINPUT8), .Z(n1251) );
NAND4_X1 U908 ( .A1(n1255), .A2(n1203), .A3(n1256), .A4(n1257), .ZN(n1167) );
NAND2_X1 U909 ( .A1(n1246), .A2(n1076), .ZN(n1203) );
NOR2_X1 U910 ( .A1(n1258), .A2(n1101), .ZN(n1076) );
INV_X1 U911 ( .A(n1259), .ZN(n1101) );
NAND4_X1 U912 ( .A1(n1075), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1255) );
OR2_X1 U913 ( .A1(n1262), .A2(KEYINPUT57), .ZN(n1261) );
NAND2_X1 U914 ( .A1(KEYINPUT57), .A2(n1263), .ZN(n1260) );
NAND3_X1 U915 ( .A1(n1240), .A2(n1254), .A3(n1103), .ZN(n1263) );
XOR2_X1 U916 ( .A(n1264), .B(n1265), .Z(n1224) );
XOR2_X1 U917 ( .A(KEYINPUT7), .B(KEYINPUT18), .Z(n1265) );
NAND2_X1 U918 ( .A1(KEYINPUT58), .A2(n1266), .ZN(n1264) );
NOR2_X1 U919 ( .A1(n1113), .A2(G952), .ZN(n1189) );
XNOR2_X1 U920 ( .A(G146), .B(n1267), .ZN(G48) );
NAND4_X1 U921 ( .A1(n1268), .A2(n1269), .A3(n1246), .A4(n1270), .ZN(n1267) );
XOR2_X1 U922 ( .A(KEYINPUT45), .B(n1111), .Z(n1270) );
XOR2_X1 U923 ( .A(G143), .B(n1271), .Z(G45) );
NOR3_X1 U924 ( .A1(n1238), .A2(KEYINPUT26), .A3(n1240), .ZN(n1271) );
NAND4_X1 U925 ( .A1(n1099), .A2(n1269), .A3(n1272), .A4(n1273), .ZN(n1238) );
INV_X1 U926 ( .A(n1245), .ZN(n1269) );
XOR2_X1 U927 ( .A(G140), .B(n1236), .Z(G42) );
AND3_X1 U928 ( .A1(n1246), .A2(n1098), .A3(n1274), .ZN(n1236) );
XOR2_X1 U929 ( .A(n1275), .B(n1237), .Z(G39) );
NAND3_X1 U930 ( .A1(n1268), .A2(n1274), .A3(n1108), .ZN(n1237) );
NAND2_X1 U931 ( .A1(n1276), .A2(n1277), .ZN(G36) );
OR2_X1 U932 ( .A1(n1231), .A2(G134), .ZN(n1277) );
XOR2_X1 U933 ( .A(n1278), .B(KEYINPUT34), .Z(n1276) );
NAND2_X1 U934 ( .A1(G134), .A2(n1231), .ZN(n1278) );
NAND2_X1 U935 ( .A1(n1253), .A2(n1274), .ZN(n1231) );
XOR2_X1 U936 ( .A(n1229), .B(n1279), .Z(G33) );
NAND2_X1 U937 ( .A1(KEYINPUT3), .A2(G131), .ZN(n1279) );
NAND3_X1 U938 ( .A1(n1274), .A2(n1246), .A3(n1099), .ZN(n1229) );
NOR3_X1 U939 ( .A1(n1087), .A2(n1089), .A3(n1245), .ZN(n1274) );
NAND2_X1 U940 ( .A1(n1103), .A2(n1280), .ZN(n1245) );
XNOR2_X1 U941 ( .A(n1112), .B(KEYINPUT39), .ZN(n1087) );
NAND2_X1 U942 ( .A1(n1281), .A2(n1282), .ZN(G30) );
NAND2_X1 U943 ( .A1(G128), .A2(n1283), .ZN(n1282) );
XOR2_X1 U944 ( .A(KEYINPUT44), .B(n1284), .Z(n1281) );
NOR2_X1 U945 ( .A1(G128), .A2(n1283), .ZN(n1284) );
NAND4_X1 U946 ( .A1(n1285), .A2(n1280), .A3(n1111), .A4(n1286), .ZN(n1283) );
AND2_X1 U947 ( .A1(n1075), .A2(n1268), .ZN(n1286) );
XOR2_X1 U948 ( .A(KEYINPUT43), .B(n1103), .Z(n1285) );
XNOR2_X1 U949 ( .A(G101), .B(n1256), .ZN(G3) );
NAND3_X1 U950 ( .A1(n1099), .A2(n1262), .A3(n1108), .ZN(n1256) );
XNOR2_X1 U951 ( .A(G125), .B(n1230), .ZN(G27) );
NAND4_X1 U952 ( .A1(n1246), .A2(n1109), .A3(n1287), .A4(n1098), .ZN(n1230) );
AND2_X1 U953 ( .A1(n1280), .A2(n1111), .ZN(n1287) );
NAND2_X1 U954 ( .A1(n1288), .A2(n1084), .ZN(n1280) );
NAND3_X1 U955 ( .A1(G902), .A2(n1289), .A3(n1148), .ZN(n1288) );
NOR2_X1 U956 ( .A1(G900), .A2(n1113), .ZN(n1148) );
XNOR2_X1 U957 ( .A(G122), .B(n1248), .ZN(G24) );
NAND4_X1 U958 ( .A1(n1290), .A2(n1259), .A3(n1272), .A4(n1273), .ZN(n1248) );
NOR2_X1 U959 ( .A1(n1291), .A2(n1292), .ZN(n1259) );
XNOR2_X1 U960 ( .A(G119), .B(n1249), .ZN(G21) );
NAND3_X1 U961 ( .A1(n1108), .A2(n1268), .A3(n1290), .ZN(n1249) );
INV_X1 U962 ( .A(n1244), .ZN(n1268) );
NAND2_X1 U963 ( .A1(n1292), .A2(n1291), .ZN(n1244) );
INV_X1 U964 ( .A(n1293), .ZN(n1292) );
NAND3_X1 U965 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(G18) );
NAND2_X1 U966 ( .A1(G116), .A2(n1297), .ZN(n1296) );
NAND2_X1 U967 ( .A1(KEYINPUT55), .A2(n1298), .ZN(n1295) );
NAND2_X1 U968 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
INV_X1 U969 ( .A(n1297), .ZN(n1300) );
XNOR2_X1 U970 ( .A(KEYINPUT28), .B(G116), .ZN(n1299) );
NAND2_X1 U971 ( .A1(n1301), .A2(n1302), .ZN(n1294) );
INV_X1 U972 ( .A(KEYINPUT55), .ZN(n1302) );
NAND2_X1 U973 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
OR3_X1 U974 ( .A1(n1297), .A2(G116), .A3(KEYINPUT28), .ZN(n1304) );
NAND2_X1 U975 ( .A1(n1290), .A2(n1253), .ZN(n1297) );
AND2_X1 U976 ( .A1(n1099), .A2(n1075), .ZN(n1253) );
NOR2_X1 U977 ( .A1(n1273), .A2(n1305), .ZN(n1075) );
NAND2_X1 U978 ( .A1(KEYINPUT28), .A2(G116), .ZN(n1303) );
XNOR2_X1 U979 ( .A(G113), .B(n1250), .ZN(G15) );
NAND3_X1 U980 ( .A1(n1099), .A2(n1246), .A3(n1290), .ZN(n1250) );
AND3_X1 U981 ( .A1(n1111), .A2(n1254), .A3(n1109), .ZN(n1290) );
NOR2_X1 U982 ( .A1(n1104), .A2(n1121), .ZN(n1109) );
INV_X1 U983 ( .A(n1105), .ZN(n1121) );
AND2_X1 U984 ( .A1(n1305), .A2(n1273), .ZN(n1246) );
NOR2_X1 U985 ( .A1(n1291), .A2(n1293), .ZN(n1099) );
XNOR2_X1 U986 ( .A(G110), .B(n1257), .ZN(G12) );
NAND3_X1 U987 ( .A1(n1098), .A2(n1262), .A3(n1108), .ZN(n1257) );
NOR2_X1 U988 ( .A1(n1272), .A2(n1273), .ZN(n1108) );
NAND3_X1 U989 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1273) );
NAND2_X1 U990 ( .A1(G475), .A2(n1309), .ZN(n1308) );
NAND2_X1 U991 ( .A1(KEYINPUT38), .A2(n1310), .ZN(n1307) );
NAND2_X1 U992 ( .A1(n1311), .A2(n1200), .ZN(n1310) );
INV_X1 U993 ( .A(G475), .ZN(n1200) );
XOR2_X1 U994 ( .A(KEYINPUT24), .B(n1133), .Z(n1311) );
INV_X1 U995 ( .A(n1309), .ZN(n1133) );
NAND2_X1 U996 ( .A1(n1312), .A2(n1313), .ZN(n1306) );
INV_X1 U997 ( .A(KEYINPUT38), .ZN(n1313) );
NAND2_X1 U998 ( .A1(n1314), .A2(n1315), .ZN(n1312) );
OR3_X1 U999 ( .A1(n1309), .A2(G475), .A3(KEYINPUT24), .ZN(n1315) );
NAND2_X1 U1000 ( .A1(KEYINPUT24), .A2(n1309), .ZN(n1314) );
NAND2_X1 U1001 ( .A1(n1202), .A2(n1316), .ZN(n1309) );
INV_X1 U1002 ( .A(n1198), .ZN(n1202) );
XOR2_X1 U1003 ( .A(n1317), .B(n1318), .Z(n1198) );
XOR2_X1 U1004 ( .A(n1319), .B(n1320), .Z(n1318) );
XOR2_X1 U1005 ( .A(G122), .B(G113), .Z(n1320) );
XOR2_X1 U1006 ( .A(G143), .B(G131), .Z(n1319) );
XOR2_X1 U1007 ( .A(n1321), .B(n1322), .Z(n1317) );
XOR2_X1 U1008 ( .A(G104), .B(n1323), .Z(n1322) );
NOR2_X1 U1009 ( .A1(KEYINPUT29), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1010 ( .A(n1154), .B(n1158), .Z(n1324) );
INV_X1 U1011 ( .A(G140), .ZN(n1154) );
XOR2_X1 U1012 ( .A(n1325), .B(n1326), .Z(n1321) );
NAND2_X1 U1013 ( .A1(G214), .A2(n1327), .ZN(n1325) );
INV_X1 U1014 ( .A(n1305), .ZN(n1272) );
XOR2_X1 U1015 ( .A(n1193), .B(n1328), .Z(n1305) );
NOR2_X1 U1016 ( .A1(KEYINPUT46), .A2(n1134), .ZN(n1328) );
OR2_X1 U1017 ( .A1(n1192), .A2(G902), .ZN(n1134) );
XNOR2_X1 U1018 ( .A(n1329), .B(n1330), .ZN(n1192) );
XOR2_X1 U1019 ( .A(G107), .B(n1331), .Z(n1330) );
XOR2_X1 U1020 ( .A(G122), .B(G116), .Z(n1331) );
XOR2_X1 U1021 ( .A(n1332), .B(n1333), .Z(n1329) );
AND2_X1 U1022 ( .A1(n1334), .A2(G217), .ZN(n1333) );
NAND2_X1 U1023 ( .A1(n1335), .A2(KEYINPUT35), .ZN(n1332) );
XOR2_X1 U1024 ( .A(n1336), .B(n1337), .Z(n1335) );
NOR2_X1 U1025 ( .A1(KEYINPUT37), .A2(n1153), .ZN(n1337) );
XOR2_X1 U1026 ( .A(G128), .B(n1338), .Z(n1336) );
INV_X1 U1027 ( .A(G478), .ZN(n1193) );
INV_X1 U1028 ( .A(n1258), .ZN(n1262) );
NAND3_X1 U1029 ( .A1(n1111), .A2(n1254), .A3(n1103), .ZN(n1258) );
AND2_X1 U1030 ( .A1(n1105), .A2(n1104), .ZN(n1103) );
NAND2_X1 U1031 ( .A1(n1127), .A2(n1124), .ZN(n1104) );
NAND2_X1 U1032 ( .A1(G469), .A2(n1339), .ZN(n1124) );
OR2_X1 U1033 ( .A1(n1339), .A2(G469), .ZN(n1127) );
NAND2_X1 U1034 ( .A1(n1340), .A2(n1316), .ZN(n1339) );
XNOR2_X1 U1035 ( .A(n1220), .B(n1219), .ZN(n1340) );
XOR2_X1 U1036 ( .A(G140), .B(n1341), .Z(n1219) );
XOR2_X1 U1037 ( .A(n1342), .B(n1343), .Z(n1220) );
XOR2_X1 U1038 ( .A(n1344), .B(n1345), .Z(n1343) );
XNOR2_X1 U1039 ( .A(KEYINPUT41), .B(KEYINPUT27), .ZN(n1345) );
NAND2_X1 U1040 ( .A1(G227), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1041 ( .A(KEYINPUT15), .B(G953), .Z(n1346) );
XOR2_X1 U1042 ( .A(n1347), .B(n1156), .Z(n1342) );
XOR2_X1 U1043 ( .A(G143), .B(KEYINPUT25), .Z(n1156) );
XOR2_X1 U1044 ( .A(n1348), .B(n1349), .Z(n1347) );
NAND2_X1 U1045 ( .A1(G221), .A2(n1350), .ZN(n1105) );
NAND2_X1 U1046 ( .A1(n1084), .A2(n1351), .ZN(n1254) );
NAND4_X1 U1047 ( .A1(G902), .A2(G953), .A3(n1289), .A4(n1352), .ZN(n1351) );
INV_X1 U1048 ( .A(G898), .ZN(n1352) );
NAND3_X1 U1049 ( .A1(n1289), .A2(n1113), .A3(G952), .ZN(n1084) );
NAND2_X1 U1050 ( .A1(G237), .A2(G234), .ZN(n1289) );
INV_X1 U1051 ( .A(n1240), .ZN(n1111) );
NAND2_X1 U1052 ( .A1(n1089), .A2(n1112), .ZN(n1240) );
NAND2_X1 U1053 ( .A1(G214), .A2(n1353), .ZN(n1112) );
XOR2_X1 U1054 ( .A(n1354), .B(n1228), .Z(n1089) );
NAND2_X1 U1055 ( .A1(G210), .A2(n1353), .ZN(n1228) );
NAND2_X1 U1056 ( .A1(n1355), .A2(n1316), .ZN(n1353) );
XOR2_X1 U1057 ( .A(KEYINPUT30), .B(G237), .Z(n1355) );
NAND2_X1 U1058 ( .A1(n1356), .A2(n1316), .ZN(n1354) );
XOR2_X1 U1059 ( .A(n1226), .B(n1266), .Z(n1356) );
XOR2_X1 U1060 ( .A(n1357), .B(n1358), .Z(n1266) );
NOR2_X1 U1061 ( .A1(KEYINPUT36), .A2(n1173), .ZN(n1358) );
XNOR2_X1 U1062 ( .A(n1359), .B(n1218), .ZN(n1173) );
XNOR2_X1 U1063 ( .A(G122), .B(KEYINPUT59), .ZN(n1359) );
NAND2_X1 U1064 ( .A1(n1360), .A2(n1361), .ZN(n1357) );
NAND2_X1 U1065 ( .A1(n1178), .A2(n1174), .ZN(n1361) );
XOR2_X1 U1066 ( .A(KEYINPUT49), .B(n1362), .Z(n1360) );
NOR2_X1 U1067 ( .A1(n1178), .A2(n1174), .ZN(n1362) );
XNOR2_X1 U1068 ( .A(G113), .B(n1363), .ZN(n1174) );
XNOR2_X1 U1069 ( .A(n1349), .B(n1364), .ZN(n1178) );
XOR2_X1 U1070 ( .A(KEYINPUT63), .B(KEYINPUT22), .Z(n1364) );
XOR2_X1 U1071 ( .A(G101), .B(n1365), .Z(n1349) );
XOR2_X1 U1072 ( .A(G107), .B(G104), .Z(n1365) );
XOR2_X1 U1073 ( .A(n1366), .B(n1367), .Z(n1226) );
XOR2_X1 U1074 ( .A(n1368), .B(n1158), .Z(n1367) );
XOR2_X1 U1075 ( .A(n1369), .B(n1370), .Z(n1366) );
AND2_X1 U1076 ( .A1(n1113), .A2(G224), .ZN(n1370) );
AND2_X1 U1077 ( .A1(n1293), .A2(n1291), .ZN(n1098) );
NAND2_X1 U1078 ( .A1(n1371), .A2(n1123), .ZN(n1291) );
NAND2_X1 U1079 ( .A1(n1372), .A2(n1373), .ZN(n1123) );
XOR2_X1 U1080 ( .A(KEYINPUT50), .B(n1120), .Z(n1371) );
NOR2_X1 U1081 ( .A1(n1373), .A2(n1372), .ZN(n1120) );
INV_X1 U1082 ( .A(n1187), .ZN(n1372) );
NAND2_X1 U1083 ( .A1(G217), .A2(n1350), .ZN(n1187) );
NAND2_X1 U1084 ( .A1(G234), .A2(n1316), .ZN(n1350) );
NAND2_X1 U1085 ( .A1(n1185), .A2(n1316), .ZN(n1373) );
XNOR2_X1 U1086 ( .A(n1374), .B(n1375), .ZN(n1185) );
XOR2_X1 U1087 ( .A(n1376), .B(n1377), .Z(n1375) );
NAND2_X1 U1088 ( .A1(KEYINPUT1), .A2(n1378), .ZN(n1377) );
XOR2_X1 U1089 ( .A(n1275), .B(n1379), .Z(n1378) );
NAND2_X1 U1090 ( .A1(G221), .A2(n1334), .ZN(n1379) );
AND2_X1 U1091 ( .A1(G234), .A2(n1113), .ZN(n1334) );
INV_X1 U1092 ( .A(G953), .ZN(n1113) );
NAND3_X1 U1093 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n1376) );
OR2_X1 U1094 ( .A1(n1383), .A2(n1341), .ZN(n1382) );
NAND2_X1 U1095 ( .A1(n1384), .A2(n1385), .ZN(n1381) );
INV_X1 U1096 ( .A(KEYINPUT48), .ZN(n1385) );
NAND2_X1 U1097 ( .A1(n1383), .A2(n1386), .ZN(n1384) );
XOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1218), .Z(n1386) );
INV_X1 U1099 ( .A(n1341), .ZN(n1218) );
NAND2_X1 U1100 ( .A1(KEYINPUT48), .A2(n1387), .ZN(n1380) );
NAND2_X1 U1101 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
NAND3_X1 U1102 ( .A1(KEYINPUT62), .A2(n1383), .A3(n1341), .ZN(n1389) );
XNOR2_X1 U1103 ( .A(G128), .B(n1390), .ZN(n1383) );
NOR2_X1 U1104 ( .A1(G119), .A2(KEYINPUT6), .ZN(n1390) );
OR2_X1 U1105 ( .A1(n1341), .A2(KEYINPUT62), .ZN(n1388) );
XNOR2_X1 U1106 ( .A(G110), .B(KEYINPUT21), .ZN(n1341) );
XOR2_X1 U1107 ( .A(n1391), .B(n1326), .Z(n1374) );
XOR2_X1 U1108 ( .A(G146), .B(KEYINPUT56), .Z(n1326) );
NAND2_X1 U1109 ( .A1(KEYINPUT17), .A2(n1392), .ZN(n1391) );
XOR2_X1 U1110 ( .A(G140), .B(n1158), .Z(n1392) );
XOR2_X1 U1111 ( .A(G125), .B(KEYINPUT23), .Z(n1158) );
XOR2_X1 U1112 ( .A(n1131), .B(G472), .Z(n1293) );
NAND2_X1 U1113 ( .A1(n1316), .A2(n1393), .ZN(n1131) );
NAND2_X1 U1114 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
OR2_X1 U1115 ( .A1(n1208), .A2(n1396), .ZN(n1395) );
XOR2_X1 U1116 ( .A(n1397), .B(KEYINPUT20), .Z(n1394) );
NAND2_X1 U1117 ( .A1(n1396), .A2(n1208), .ZN(n1397) );
XNOR2_X1 U1118 ( .A(n1398), .B(n1399), .ZN(n1208) );
XNOR2_X1 U1119 ( .A(G113), .B(n1369), .ZN(n1399) );
NAND2_X1 U1120 ( .A1(n1400), .A2(n1338), .ZN(n1369) );
INV_X1 U1121 ( .A(G143), .ZN(n1338) );
XNOR2_X1 U1122 ( .A(KEYINPUT61), .B(KEYINPUT10), .ZN(n1400) );
XOR2_X1 U1123 ( .A(n1348), .B(n1401), .Z(n1398) );
NOR2_X1 U1124 ( .A1(KEYINPUT4), .A2(n1363), .ZN(n1401) );
XNOR2_X1 U1125 ( .A(G119), .B(G116), .ZN(n1363) );
XOR2_X1 U1126 ( .A(n1157), .B(n1402), .Z(n1348) );
XOR2_X1 U1127 ( .A(n1153), .B(n1403), .Z(n1402) );
NAND2_X1 U1128 ( .A1(KEYINPUT51), .A2(n1275), .ZN(n1403) );
INV_X1 U1129 ( .A(G137), .ZN(n1275) );
INV_X1 U1130 ( .A(G134), .ZN(n1153) );
XNOR2_X1 U1131 ( .A(G131), .B(n1368), .ZN(n1157) );
XOR2_X1 U1132 ( .A(G146), .B(G128), .Z(n1368) );
XNOR2_X1 U1133 ( .A(n1207), .B(n1404), .ZN(n1396) );
NOR2_X1 U1134 ( .A1(G101), .A2(KEYINPUT33), .ZN(n1404) );
NAND2_X1 U1135 ( .A1(G210), .A2(n1327), .ZN(n1207) );
NOR2_X1 U1136 ( .A1(G953), .A2(G237), .ZN(n1327) );
INV_X1 U1137 ( .A(G902), .ZN(n1316) );
endmodule


