//Key = 1111101001101011111000110101100010000111111101111100100010111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352;

NAND2_X1 U733 ( .A1(n1025), .A2(n1026), .ZN(G9) );
NAND2_X1 U734 ( .A1(G107), .A2(n1027), .ZN(n1026) );
XOR2_X1 U735 ( .A(KEYINPUT4), .B(n1028), .Z(n1025) );
NOR2_X1 U736 ( .A1(G107), .A2(n1027), .ZN(n1028) );
NOR2_X1 U737 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
XOR2_X1 U739 ( .A(KEYINPUT28), .B(n1035), .Z(n1032) );
NOR3_X1 U740 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
INV_X1 U742 ( .A(n1041), .ZN(n1040) );
NOR2_X1 U743 ( .A1(n1042), .A2(n1043), .ZN(n1039) );
AND2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U745 ( .A1(n1046), .A2(n1047), .ZN(n1042) );
NOR4_X1 U746 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1037) );
XOR2_X1 U747 ( .A(KEYINPUT57), .B(n1052), .Z(n1036) );
NOR4_X1 U748 ( .A1(n1053), .A2(n1054), .A3(n1048), .A4(n1051), .ZN(n1052) );
INV_X1 U749 ( .A(n1055), .ZN(n1051) );
NAND4_X1 U750 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1031) );
NAND3_X1 U751 ( .A1(n1060), .A2(n1061), .A3(n1055), .ZN(n1057) );
NAND2_X1 U752 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND3_X1 U753 ( .A1(n1044), .A2(n1064), .A3(n1065), .ZN(n1063) );
NAND2_X1 U754 ( .A1(n1066), .A2(n1067), .ZN(n1062) );
XOR2_X1 U755 ( .A(KEYINPUT7), .B(n1068), .Z(n1067) );
NOR2_X1 U756 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U757 ( .A1(n1044), .A2(n1071), .ZN(n1056) );
NAND2_X1 U758 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND3_X1 U759 ( .A1(n1066), .A2(n1074), .A3(n1055), .ZN(n1073) );
NOR2_X1 U760 ( .A1(n1075), .A2(n1047), .ZN(n1055) );
NAND2_X1 U761 ( .A1(n1041), .A2(n1076), .ZN(n1072) );
NOR3_X1 U762 ( .A1(n1050), .A2(n1054), .A3(n1075), .ZN(n1041) );
INV_X1 U763 ( .A(n1066), .ZN(n1050) );
NOR3_X1 U764 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1029) );
INV_X1 U765 ( .A(n1058), .ZN(n1077) );
NAND4_X1 U766 ( .A1(n1078), .A2(n1060), .A3(n1079), .A4(n1080), .ZN(n1058) );
NOR4_X1 U767 ( .A1(n1064), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1080) );
XNOR2_X1 U768 ( .A(n1084), .B(n1085), .ZN(n1083) );
NAND2_X1 U769 ( .A1(KEYINPUT18), .A2(n1086), .ZN(n1084) );
XOR2_X1 U770 ( .A(n1087), .B(n1088), .Z(n1082) );
NAND2_X1 U771 ( .A1(KEYINPUT56), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U772 ( .A(G469), .B(n1090), .ZN(n1079) );
NOR2_X1 U773 ( .A1(KEYINPUT13), .A2(n1091), .ZN(n1090) );
XOR2_X1 U774 ( .A(n1092), .B(n1093), .Z(G72) );
NOR2_X1 U775 ( .A1(n1094), .A2(n1059), .ZN(n1093) );
NOR2_X1 U776 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U777 ( .A1(KEYINPUT29), .A2(n1097), .ZN(n1092) );
XOR2_X1 U778 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U779 ( .A1(n1100), .A2(G953), .ZN(n1099) );
NAND2_X1 U780 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U781 ( .A1(G953), .A2(n1096), .ZN(n1102) );
XOR2_X1 U782 ( .A(n1103), .B(n1104), .Z(n1101) );
XNOR2_X1 U783 ( .A(n1105), .B(n1106), .ZN(n1104) );
XOR2_X1 U784 ( .A(KEYINPUT6), .B(n1107), .Z(n1103) );
NOR2_X1 U785 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U786 ( .A(n1110), .B(KEYINPUT15), .Z(n1109) );
NAND2_X1 U787 ( .A1(G131), .A2(n1111), .ZN(n1110) );
NOR2_X1 U788 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
XNOR2_X1 U789 ( .A(KEYINPUT24), .B(n1113), .ZN(n1112) );
NAND2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U791 ( .A1(G134), .A2(n1116), .ZN(n1115) );
XOR2_X1 U792 ( .A(KEYINPUT48), .B(n1117), .Z(n1114) );
NOR2_X1 U793 ( .A1(G134), .A2(n1116), .ZN(n1117) );
XOR2_X1 U794 ( .A(n1118), .B(n1119), .Z(G69) );
NOR2_X1 U795 ( .A1(n1120), .A2(G953), .ZN(n1119) );
XOR2_X1 U796 ( .A(n1121), .B(n1122), .Z(n1118) );
NOR2_X1 U797 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U798 ( .A1(G224), .A2(n1059), .ZN(n1123) );
NAND2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(n1121) );
INV_X1 U800 ( .A(n1124), .ZN(n1126) );
XOR2_X1 U801 ( .A(n1127), .B(n1128), .Z(n1125) );
NOR2_X1 U802 ( .A1(KEYINPUT5), .A2(n1129), .ZN(n1127) );
NOR2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(G66) );
XNOR2_X1 U804 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR3_X1 U805 ( .A1(n1134), .A2(KEYINPUT35), .A3(n1135), .ZN(n1133) );
NOR2_X1 U806 ( .A1(n1130), .A2(n1136), .ZN(G63) );
XNOR2_X1 U807 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U808 ( .A1(n1139), .A2(n1134), .ZN(n1138) );
NOR3_X1 U809 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(G60) );
AND3_X1 U810 ( .A1(KEYINPUT34), .A2(G952), .A3(G953), .ZN(n1142) );
NOR2_X1 U811 ( .A1(KEYINPUT34), .A2(n1143), .ZN(n1141) );
INV_X1 U812 ( .A(n1130), .ZN(n1143) );
XOR2_X1 U813 ( .A(n1144), .B(n1145), .Z(n1140) );
NOR2_X1 U814 ( .A1(n1089), .A2(n1134), .ZN(n1145) );
NAND3_X1 U815 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(G6) );
NAND2_X1 U816 ( .A1(KEYINPUT36), .A2(n1149), .ZN(n1148) );
OR3_X1 U817 ( .A1(n1149), .A2(KEYINPUT36), .A3(G104), .ZN(n1147) );
NAND2_X1 U818 ( .A1(G104), .A2(n1150), .ZN(n1146) );
NAND2_X1 U819 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
INV_X1 U820 ( .A(KEYINPUT36), .ZN(n1152) );
XOR2_X1 U821 ( .A(n1149), .B(KEYINPUT12), .Z(n1151) );
NAND3_X1 U822 ( .A1(n1153), .A2(n1045), .A3(n1154), .ZN(n1149) );
NOR3_X1 U823 ( .A1(n1054), .A2(n1155), .A3(n1046), .ZN(n1154) );
XNOR2_X1 U824 ( .A(n1156), .B(KEYINPUT3), .ZN(n1153) );
NOR2_X1 U825 ( .A1(n1130), .A2(n1157), .ZN(G57) );
XOR2_X1 U826 ( .A(n1158), .B(n1159), .Z(n1157) );
XNOR2_X1 U827 ( .A(n1160), .B(n1161), .ZN(n1159) );
XOR2_X1 U828 ( .A(KEYINPUT30), .B(n1162), .Z(n1158) );
NOR2_X1 U829 ( .A1(n1163), .A2(n1134), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1130), .A2(n1164), .ZN(G54) );
NOR2_X1 U831 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
XOR2_X1 U832 ( .A(KEYINPUT50), .B(n1167), .Z(n1166) );
AND2_X1 U833 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U834 ( .A1(n1169), .A2(n1168), .ZN(n1165) );
XNOR2_X1 U835 ( .A(n1170), .B(n1171), .ZN(n1168) );
XOR2_X1 U836 ( .A(KEYINPUT23), .B(n1172), .Z(n1171) );
NOR2_X1 U837 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NOR2_X1 U838 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XNOR2_X1 U839 ( .A(KEYINPUT27), .B(n1177), .ZN(n1176) );
XNOR2_X1 U840 ( .A(n1178), .B(n1179), .ZN(n1170) );
NAND2_X1 U841 ( .A1(n1180), .A2(n1181), .ZN(n1178) );
NAND2_X1 U842 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U843 ( .A(KEYINPUT22), .B(n1184), .ZN(n1183) );
XNOR2_X1 U844 ( .A(n1185), .B(KEYINPUT10), .ZN(n1182) );
NAND2_X1 U845 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
XNOR2_X1 U846 ( .A(KEYINPUT10), .B(n1105), .ZN(n1187) );
INV_X1 U847 ( .A(n1185), .ZN(n1105) );
XNOR2_X1 U848 ( .A(n1188), .B(KEYINPUT37), .ZN(n1186) );
NOR2_X1 U849 ( .A1(n1134), .A2(n1189), .ZN(n1169) );
INV_X1 U850 ( .A(G469), .ZN(n1189) );
NOR3_X1 U851 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(G51) );
AND2_X1 U852 ( .A1(n1130), .A2(KEYINPUT52), .ZN(n1192) );
NOR2_X1 U853 ( .A1(n1059), .A2(G952), .ZN(n1130) );
NOR3_X1 U854 ( .A1(KEYINPUT52), .A2(G953), .A3(G952), .ZN(n1191) );
XOR2_X1 U855 ( .A(n1193), .B(n1194), .Z(n1190) );
XOR2_X1 U856 ( .A(n1195), .B(n1196), .Z(n1193) );
NOR2_X1 U857 ( .A1(n1086), .A2(n1134), .ZN(n1196) );
NAND2_X1 U858 ( .A1(G902), .A2(n1197), .ZN(n1134) );
NAND2_X1 U859 ( .A1(n1120), .A2(n1100), .ZN(n1197) );
INV_X1 U860 ( .A(n1033), .ZN(n1100) );
NAND4_X1 U861 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1033) );
AND4_X1 U862 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
NAND3_X1 U863 ( .A1(n1076), .A2(n1206), .A3(n1207), .ZN(n1200) );
XNOR2_X1 U864 ( .A(KEYINPUT61), .B(n1049), .ZN(n1206) );
NAND3_X1 U865 ( .A1(n1156), .A2(n1208), .A3(n1045), .ZN(n1198) );
NAND2_X1 U866 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
INV_X1 U867 ( .A(n1034), .ZN(n1120) );
NAND4_X1 U868 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1034) );
NOR4_X1 U869 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NOR3_X1 U870 ( .A1(n1219), .A2(n1046), .A3(n1054), .ZN(n1218) );
INV_X1 U871 ( .A(n1060), .ZN(n1054) );
NAND3_X1 U872 ( .A1(n1220), .A2(n1221), .A3(n1045), .ZN(n1219) );
OR2_X1 U873 ( .A1(n1222), .A2(KEYINPUT11), .ZN(n1221) );
NAND2_X1 U874 ( .A1(KEYINPUT11), .A2(n1223), .ZN(n1220) );
NAND2_X1 U875 ( .A1(n1155), .A2(n1156), .ZN(n1223) );
AND2_X1 U876 ( .A1(n1027), .A2(n1224), .ZN(n1213) );
NAND4_X1 U877 ( .A1(n1222), .A2(n1076), .A3(n1060), .A4(n1225), .ZN(n1027) );
NAND2_X1 U878 ( .A1(KEYINPUT32), .A2(n1226), .ZN(n1195) );
XNOR2_X1 U879 ( .A(G146), .B(n1227), .ZN(G48) );
NAND3_X1 U880 ( .A1(n1228), .A2(n1045), .A3(n1229), .ZN(n1227) );
XNOR2_X1 U881 ( .A(n1156), .B(KEYINPUT42), .ZN(n1229) );
XNOR2_X1 U882 ( .A(G143), .B(n1199), .ZN(G45) );
NAND4_X1 U883 ( .A1(n1225), .A2(n1156), .A3(n1230), .A4(n1231), .ZN(n1199) );
AND3_X1 U884 ( .A1(n1232), .A2(n1233), .A3(n1234), .ZN(n1231) );
XOR2_X1 U885 ( .A(G140), .B(n1235), .Z(G42) );
NOR2_X1 U886 ( .A1(KEYINPUT20), .A2(n1205), .ZN(n1235) );
NAND3_X1 U887 ( .A1(n1045), .A2(n1074), .A3(n1207), .ZN(n1205) );
XNOR2_X1 U888 ( .A(n1236), .B(n1116), .ZN(G39) );
INV_X1 U889 ( .A(G137), .ZN(n1116) );
NAND2_X1 U890 ( .A1(KEYINPUT9), .A2(n1204), .ZN(n1236) );
NAND3_X1 U891 ( .A1(n1228), .A2(n1237), .A3(n1066), .ZN(n1204) );
NAND2_X1 U892 ( .A1(n1238), .A2(n1239), .ZN(G36) );
NAND2_X1 U893 ( .A1(G134), .A2(n1240), .ZN(n1239) );
XOR2_X1 U894 ( .A(KEYINPUT62), .B(n1241), .Z(n1238) );
NOR2_X1 U895 ( .A1(G134), .A2(n1240), .ZN(n1241) );
NAND3_X1 U896 ( .A1(n1230), .A2(n1076), .A3(n1207), .ZN(n1240) );
XNOR2_X1 U897 ( .A(G131), .B(n1203), .ZN(G33) );
NAND3_X1 U898 ( .A1(n1045), .A2(n1230), .A3(n1207), .ZN(n1203) );
AND3_X1 U899 ( .A1(n1225), .A2(n1233), .A3(n1066), .ZN(n1207) );
NOR2_X1 U900 ( .A1(n1242), .A2(n1243), .ZN(n1066) );
XNOR2_X1 U901 ( .A(G128), .B(n1202), .ZN(G30) );
NAND3_X1 U902 ( .A1(n1076), .A2(n1156), .A3(n1228), .ZN(n1202) );
INV_X1 U903 ( .A(n1210), .ZN(n1228) );
NAND4_X1 U904 ( .A1(n1225), .A2(n1244), .A3(n1245), .A4(n1233), .ZN(n1210) );
INV_X1 U905 ( .A(n1046), .ZN(n1225) );
XOR2_X1 U906 ( .A(n1246), .B(n1217), .Z(G3) );
AND2_X1 U907 ( .A1(n1230), .A2(n1247), .ZN(n1217) );
XNOR2_X1 U908 ( .A(G101), .B(KEYINPUT25), .ZN(n1246) );
XNOR2_X1 U909 ( .A(G125), .B(n1248), .ZN(G27) );
NAND3_X1 U910 ( .A1(n1249), .A2(n1045), .A3(n1250), .ZN(n1248) );
XNOR2_X1 U911 ( .A(n1156), .B(KEYINPUT59), .ZN(n1250) );
INV_X1 U912 ( .A(n1209), .ZN(n1249) );
NAND3_X1 U913 ( .A1(n1074), .A2(n1233), .A3(n1044), .ZN(n1209) );
NAND2_X1 U914 ( .A1(n1075), .A2(n1251), .ZN(n1233) );
NAND4_X1 U915 ( .A1(G902), .A2(G953), .A3(n1252), .A4(n1096), .ZN(n1251) );
INV_X1 U916 ( .A(G900), .ZN(n1096) );
XNOR2_X1 U917 ( .A(G122), .B(n1211), .ZN(G24) );
NAND4_X1 U918 ( .A1(n1253), .A2(n1060), .A3(n1232), .A4(n1234), .ZN(n1211) );
NOR2_X1 U919 ( .A1(n1245), .A2(n1244), .ZN(n1060) );
XNOR2_X1 U920 ( .A(G119), .B(n1212), .ZN(G21) );
NAND4_X1 U921 ( .A1(n1253), .A2(n1237), .A3(n1244), .A4(n1245), .ZN(n1212) );
XOR2_X1 U922 ( .A(G116), .B(n1216), .Z(G18) );
AND3_X1 U923 ( .A1(n1253), .A2(n1076), .A3(n1230), .ZN(n1216) );
NOR2_X1 U924 ( .A1(n1234), .A2(n1078), .ZN(n1076) );
XOR2_X1 U925 ( .A(G113), .B(n1254), .Z(G15) );
NOR2_X1 U926 ( .A1(KEYINPUT26), .A2(n1224), .ZN(n1254) );
NAND3_X1 U927 ( .A1(n1230), .A2(n1253), .A3(n1045), .ZN(n1224) );
AND2_X1 U928 ( .A1(n1078), .A2(n1234), .ZN(n1045) );
INV_X1 U929 ( .A(n1232), .ZN(n1078) );
NOR2_X1 U930 ( .A1(n1048), .A2(n1255), .ZN(n1253) );
INV_X1 U931 ( .A(n1044), .ZN(n1048) );
NOR2_X1 U932 ( .A1(n1069), .A2(n1081), .ZN(n1044) );
INV_X1 U933 ( .A(n1070), .ZN(n1081) );
XNOR2_X1 U934 ( .A(n1256), .B(KEYINPUT46), .ZN(n1069) );
INV_X1 U935 ( .A(n1049), .ZN(n1230) );
NAND2_X1 U936 ( .A1(n1257), .A2(n1245), .ZN(n1049) );
XNOR2_X1 U937 ( .A(G110), .B(n1258), .ZN(G12) );
NAND2_X1 U938 ( .A1(KEYINPUT43), .A2(n1215), .ZN(n1258) );
AND2_X1 U939 ( .A1(n1247), .A2(n1074), .ZN(n1215) );
NOR2_X1 U940 ( .A1(n1245), .A2(n1257), .ZN(n1074) );
INV_X1 U941 ( .A(n1244), .ZN(n1257) );
XOR2_X1 U942 ( .A(n1259), .B(n1135), .Z(n1244) );
NAND2_X1 U943 ( .A1(G217), .A2(n1260), .ZN(n1135) );
NAND2_X1 U944 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
NAND2_X1 U945 ( .A1(n1132), .A2(n1262), .ZN(n1259) );
XNOR2_X1 U946 ( .A(n1263), .B(n1264), .ZN(n1132) );
XOR2_X1 U947 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U948 ( .A(n1267), .B(G125), .Z(n1266) );
NAND2_X1 U949 ( .A1(G221), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U950 ( .A(G137), .B(G146), .ZN(n1265) );
XOR2_X1 U951 ( .A(n1269), .B(n1270), .Z(n1263) );
XNOR2_X1 U952 ( .A(n1271), .B(n1177), .ZN(n1269) );
NAND2_X1 U953 ( .A1(KEYINPUT17), .A2(G128), .ZN(n1271) );
XOR2_X1 U954 ( .A(n1272), .B(n1163), .Z(n1245) );
INV_X1 U955 ( .A(G472), .ZN(n1163) );
NAND2_X1 U956 ( .A1(n1273), .A2(n1262), .ZN(n1272) );
XOR2_X1 U957 ( .A(n1274), .B(n1161), .Z(n1273) );
XOR2_X1 U958 ( .A(n1275), .B(n1276), .Z(n1161) );
XNOR2_X1 U959 ( .A(n1277), .B(n1278), .ZN(n1276) );
NOR2_X1 U960 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U961 ( .A(G210), .ZN(n1279) );
XOR2_X1 U962 ( .A(n1281), .B(n1282), .Z(n1275) );
NAND2_X1 U963 ( .A1(n1283), .A2(n1284), .ZN(n1274) );
NAND2_X1 U964 ( .A1(n1160), .A2(n1285), .ZN(n1284) );
INV_X1 U965 ( .A(KEYINPUT55), .ZN(n1285) );
XOR2_X1 U966 ( .A(n1286), .B(n1287), .Z(n1160) );
NAND3_X1 U967 ( .A1(n1286), .A2(n1287), .A3(KEYINPUT55), .ZN(n1283) );
NOR3_X1 U968 ( .A1(n1255), .A2(n1046), .A3(n1047), .ZN(n1247) );
INV_X1 U969 ( .A(n1237), .ZN(n1047) );
NOR2_X1 U970 ( .A1(n1232), .A2(n1234), .ZN(n1237) );
XOR2_X1 U971 ( .A(n1088), .B(n1288), .Z(n1234) );
XNOR2_X1 U972 ( .A(KEYINPUT53), .B(n1089), .ZN(n1288) );
INV_X1 U973 ( .A(G475), .ZN(n1089) );
NOR2_X1 U974 ( .A1(n1144), .A2(G902), .ZN(n1088) );
XOR2_X1 U975 ( .A(n1289), .B(n1290), .Z(n1144) );
XNOR2_X1 U976 ( .A(n1282), .B(n1291), .ZN(n1290) );
XOR2_X1 U977 ( .A(n1292), .B(n1293), .Z(n1289) );
NAND2_X1 U978 ( .A1(n1294), .A2(KEYINPUT38), .ZN(n1292) );
XOR2_X1 U979 ( .A(n1295), .B(n1296), .Z(n1294) );
XNOR2_X1 U980 ( .A(n1113), .B(n1297), .ZN(n1296) );
NOR2_X1 U981 ( .A1(n1298), .A2(n1280), .ZN(n1297) );
NAND2_X1 U982 ( .A1(n1299), .A2(n1059), .ZN(n1280) );
XNOR2_X1 U983 ( .A(KEYINPUT45), .B(n1300), .ZN(n1299) );
INV_X1 U984 ( .A(G214), .ZN(n1298) );
INV_X1 U985 ( .A(G131), .ZN(n1113) );
XNOR2_X1 U986 ( .A(n1106), .B(n1301), .ZN(n1295) );
XOR2_X1 U987 ( .A(G140), .B(G125), .Z(n1106) );
XOR2_X1 U988 ( .A(n1302), .B(n1139), .Z(n1232) );
INV_X1 U989 ( .A(G478), .ZN(n1139) );
NAND2_X1 U990 ( .A1(n1137), .A2(n1262), .ZN(n1302) );
XNOR2_X1 U991 ( .A(n1303), .B(n1304), .ZN(n1137) );
XNOR2_X1 U992 ( .A(n1305), .B(n1306), .ZN(n1304) );
XOR2_X1 U993 ( .A(n1307), .B(n1308), .Z(n1306) );
NOR2_X1 U994 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U995 ( .A(n1311), .B(KEYINPUT1), .Z(n1310) );
NAND2_X1 U996 ( .A1(G134), .A2(n1312), .ZN(n1311) );
NOR2_X1 U997 ( .A1(G134), .A2(n1312), .ZN(n1309) );
XNOR2_X1 U998 ( .A(n1313), .B(n1314), .ZN(n1312) );
INV_X1 U999 ( .A(G128), .ZN(n1314) );
NAND2_X1 U1000 ( .A1(KEYINPUT40), .A2(n1315), .ZN(n1313) );
NAND2_X1 U1001 ( .A1(G217), .A2(n1268), .ZN(n1307) );
AND2_X1 U1002 ( .A1(G234), .A2(n1059), .ZN(n1268) );
XOR2_X1 U1003 ( .A(n1316), .B(n1317), .Z(n1303) );
NOR2_X1 U1004 ( .A1(KEYINPUT44), .A2(G107), .ZN(n1317) );
XNOR2_X1 U1005 ( .A(G116), .B(KEYINPUT8), .ZN(n1316) );
NAND2_X1 U1006 ( .A1(n1256), .A2(n1070), .ZN(n1046) );
NAND2_X1 U1007 ( .A1(G221), .A2(n1318), .ZN(n1070) );
XOR2_X1 U1008 ( .A(KEYINPUT39), .B(n1319), .Z(n1318) );
AND2_X1 U1009 ( .A1(n1262), .A2(n1261), .ZN(n1319) );
XNOR2_X1 U1010 ( .A(n1091), .B(G469), .ZN(n1256) );
NAND2_X1 U1011 ( .A1(n1320), .A2(n1262), .ZN(n1091) );
XOR2_X1 U1012 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1013 ( .A(n1184), .B(n1185), .ZN(n1322) );
XOR2_X1 U1014 ( .A(G128), .B(n1301), .Z(n1185) );
INV_X1 U1015 ( .A(n1188), .ZN(n1184) );
XOR2_X1 U1016 ( .A(G101), .B(n1323), .Z(n1188) );
NOR2_X1 U1017 ( .A1(n1324), .A2(n1325), .ZN(n1321) );
NOR2_X1 U1018 ( .A1(n1287), .A2(n1326), .ZN(n1325) );
XNOR2_X1 U1019 ( .A(n1175), .B(n1177), .ZN(n1326) );
NOR2_X1 U1020 ( .A1(n1327), .A2(n1179), .ZN(n1324) );
INV_X1 U1021 ( .A(n1287), .ZN(n1179) );
XOR2_X1 U1022 ( .A(G131), .B(n1328), .Z(n1287) );
NOR2_X1 U1023 ( .A1(KEYINPUT21), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1024 ( .A(G137), .B(G134), .ZN(n1329) );
NOR2_X1 U1025 ( .A1(n1330), .A2(n1173), .ZN(n1327) );
AND2_X1 U1026 ( .A1(n1175), .A2(n1177), .ZN(n1173) );
NOR2_X1 U1027 ( .A1(n1175), .A2(n1177), .ZN(n1330) );
XNOR2_X1 U1028 ( .A(G110), .B(G140), .ZN(n1177) );
NOR2_X1 U1029 ( .A1(n1095), .A2(G953), .ZN(n1175) );
INV_X1 U1030 ( .A(G227), .ZN(n1095) );
INV_X1 U1031 ( .A(n1222), .ZN(n1255) );
NOR2_X1 U1032 ( .A1(n1053), .A2(n1155), .ZN(n1222) );
AND2_X1 U1033 ( .A1(n1331), .A2(n1075), .ZN(n1155) );
NAND3_X1 U1034 ( .A1(n1252), .A2(n1059), .A3(G952), .ZN(n1075) );
NAND3_X1 U1035 ( .A1(n1124), .A2(n1252), .A3(G902), .ZN(n1331) );
NAND2_X1 U1036 ( .A1(G237), .A2(n1261), .ZN(n1252) );
XNOR2_X1 U1037 ( .A(G234), .B(KEYINPUT49), .ZN(n1261) );
NOR2_X1 U1038 ( .A1(G898), .A2(n1059), .ZN(n1124) );
INV_X1 U1039 ( .A(n1156), .ZN(n1053) );
NOR2_X1 U1040 ( .A1(n1243), .A2(n1065), .ZN(n1156) );
INV_X1 U1041 ( .A(n1242), .ZN(n1065) );
XOR2_X1 U1042 ( .A(n1085), .B(n1086), .Z(n1242) );
NAND2_X1 U1043 ( .A1(G210), .A2(n1332), .ZN(n1086) );
NAND2_X1 U1044 ( .A1(n1333), .A2(n1262), .ZN(n1085) );
XOR2_X1 U1045 ( .A(n1226), .B(n1194), .Z(n1333) );
XNOR2_X1 U1046 ( .A(n1334), .B(n1335), .ZN(n1194) );
XOR2_X1 U1047 ( .A(G125), .B(n1336), .Z(n1335) );
AND2_X1 U1048 ( .A1(n1059), .A2(G224), .ZN(n1336) );
INV_X1 U1049 ( .A(G953), .ZN(n1059) );
INV_X1 U1050 ( .A(n1286), .ZN(n1334) );
XOR2_X1 U1051 ( .A(G128), .B(n1337), .Z(n1286) );
NOR2_X1 U1052 ( .A1(n1338), .A2(n1339), .ZN(n1337) );
NOR3_X1 U1053 ( .A1(n1340), .A2(G146), .A3(n1315), .ZN(n1339) );
INV_X1 U1054 ( .A(KEYINPUT31), .ZN(n1340) );
NOR2_X1 U1055 ( .A1(KEYINPUT31), .A2(n1301), .ZN(n1338) );
XNOR2_X1 U1056 ( .A(n1315), .B(G146), .ZN(n1301) );
INV_X1 U1057 ( .A(G143), .ZN(n1315) );
XNOR2_X1 U1058 ( .A(n1341), .B(n1129), .ZN(n1226) );
XOR2_X1 U1059 ( .A(n1281), .B(n1342), .Z(n1129) );
XOR2_X1 U1060 ( .A(n1343), .B(n1344), .Z(n1342) );
NAND2_X1 U1061 ( .A1(KEYINPUT58), .A2(n1282), .ZN(n1344) );
XOR2_X1 U1062 ( .A(G113), .B(KEYINPUT60), .Z(n1282) );
NAND2_X1 U1063 ( .A1(n1345), .A2(n1346), .ZN(n1343) );
OR2_X1 U1064 ( .A1(n1277), .A2(n1347), .ZN(n1346) );
XOR2_X1 U1065 ( .A(n1348), .B(KEYINPUT33), .Z(n1345) );
NAND2_X1 U1066 ( .A1(n1347), .A2(n1277), .ZN(n1348) );
INV_X1 U1067 ( .A(G101), .ZN(n1277) );
XNOR2_X1 U1068 ( .A(n1349), .B(n1323), .ZN(n1347) );
XNOR2_X1 U1069 ( .A(n1350), .B(n1293), .ZN(n1323) );
XOR2_X1 U1070 ( .A(G104), .B(KEYINPUT41), .Z(n1293) );
XNOR2_X1 U1071 ( .A(G107), .B(KEYINPUT2), .ZN(n1350) );
XNOR2_X1 U1072 ( .A(KEYINPUT19), .B(KEYINPUT14), .ZN(n1349) );
XNOR2_X1 U1073 ( .A(G116), .B(n1270), .ZN(n1281) );
XOR2_X1 U1074 ( .A(G119), .B(KEYINPUT51), .Z(n1270) );
XOR2_X1 U1075 ( .A(n1351), .B(KEYINPUT54), .Z(n1341) );
NAND2_X1 U1076 ( .A1(KEYINPUT47), .A2(n1128), .ZN(n1351) );
XNOR2_X1 U1077 ( .A(n1352), .B(G110), .ZN(n1128) );
NAND2_X1 U1078 ( .A1(KEYINPUT0), .A2(n1291), .ZN(n1352) );
INV_X1 U1079 ( .A(n1305), .ZN(n1291) );
XOR2_X1 U1080 ( .A(G122), .B(KEYINPUT63), .Z(n1305) );
XNOR2_X1 U1081 ( .A(n1064), .B(KEYINPUT16), .ZN(n1243) );
AND2_X1 U1082 ( .A1(G214), .A2(n1332), .ZN(n1064) );
NAND2_X1 U1083 ( .A1(n1300), .A2(n1262), .ZN(n1332) );
INV_X1 U1084 ( .A(G902), .ZN(n1262) );
INV_X1 U1085 ( .A(G237), .ZN(n1300) );
endmodule


