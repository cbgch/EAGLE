//Key = 0100111011001111001111001100011101101001101110000001000001110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366;

XOR2_X1 U743 ( .A(n1035), .B(n1036), .Z(G9) );
NOR2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(G75) );
XOR2_X1 U745 ( .A(n1039), .B(KEYINPUT43), .Z(n1038) );
NAND4_X1 U746 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NAND4_X1 U747 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
NAND2_X1 U748 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U749 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U750 ( .A1(n1052), .A2(n1053), .ZN(n1042) );
NAND3_X1 U751 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
XOR2_X1 U752 ( .A(n1057), .B(KEYINPUT54), .Z(n1056) );
NAND3_X1 U753 ( .A1(n1058), .A2(n1059), .A3(n1044), .ZN(n1057) );
NAND2_X1 U754 ( .A1(n1060), .A2(n1061), .ZN(n1055) );
INV_X1 U755 ( .A(KEYINPUT1), .ZN(n1061) );
NAND2_X1 U756 ( .A1(n1044), .A2(n1062), .ZN(n1060) );
NOR2_X1 U757 ( .A1(n1063), .A2(n1064), .ZN(n1044) );
NAND2_X1 U758 ( .A1(n1065), .A2(n1066), .ZN(n1054) );
NAND2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U760 ( .A1(n1046), .A2(n1069), .A3(n1045), .ZN(n1068) );
NAND2_X1 U761 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U762 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U763 ( .A1(n1074), .A2(n1075), .ZN(n1067) );
NAND2_X1 U764 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U765 ( .A1(n1046), .A2(n1078), .ZN(n1077) );
NAND2_X1 U766 ( .A1(KEYINPUT1), .A2(n1062), .ZN(n1076) );
INV_X1 U767 ( .A(n1063), .ZN(n1065) );
INV_X1 U768 ( .A(n1079), .ZN(n1041) );
NOR2_X1 U769 ( .A1(G952), .A2(n1079), .ZN(n1037) );
NAND2_X1 U770 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U771 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR4_X1 U772 ( .A1(n1050), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1083) );
XOR2_X1 U773 ( .A(n1051), .B(KEYINPUT14), .Z(n1085) );
AND2_X1 U774 ( .A1(n1087), .A2(n1088), .ZN(n1084) );
NOR4_X1 U775 ( .A1(n1064), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1082) );
XOR2_X1 U776 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U777 ( .A(KEYINPUT9), .B(n1094), .Z(n1093) );
NOR2_X1 U778 ( .A1(KEYINPUT16), .A2(n1095), .ZN(n1092) );
INV_X1 U779 ( .A(n1096), .ZN(n1095) );
XOR2_X1 U780 ( .A(KEYINPUT37), .B(n1097), .Z(n1090) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1087), .ZN(n1097) );
XOR2_X1 U782 ( .A(n1098), .B(n1099), .Z(G72) );
XOR2_X1 U783 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U784 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U785 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U786 ( .A(n1106), .B(n1107), .Z(n1105) );
XOR2_X1 U787 ( .A(n1108), .B(n1109), .Z(n1104) );
XOR2_X1 U788 ( .A(KEYINPUT41), .B(G140), .Z(n1109) );
NAND2_X1 U789 ( .A1(KEYINPUT21), .A2(G125), .ZN(n1108) );
NOR2_X1 U790 ( .A1(G900), .A2(n1080), .ZN(n1102) );
NAND2_X1 U791 ( .A1(n1080), .A2(n1110), .ZN(n1100) );
NAND2_X1 U792 ( .A1(G953), .A2(n1111), .ZN(n1098) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1111) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U795 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U796 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U797 ( .A(KEYINPUT53), .B(G953), .Z(n1117) );
INV_X1 U798 ( .A(n1118), .ZN(n1116) );
NOR2_X1 U799 ( .A1(KEYINPUT60), .A2(n1119), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1120), .A2(n1080), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND4_X1 U802 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1112) );
NAND2_X1 U803 ( .A1(KEYINPUT45), .A2(n1127), .ZN(n1126) );
NAND2_X1 U804 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XNOR2_X1 U805 ( .A(KEYINPUT36), .B(n1130), .ZN(n1128) );
NAND2_X1 U806 ( .A1(n1131), .A2(n1132), .ZN(n1125) );
INV_X1 U807 ( .A(KEYINPUT45), .ZN(n1132) );
NAND2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
OR2_X1 U809 ( .A1(n1130), .A2(KEYINPUT36), .ZN(n1134) );
NAND3_X1 U810 ( .A1(n1130), .A2(n1129), .A3(KEYINPUT36), .ZN(n1133) );
OR2_X1 U811 ( .A1(n1129), .A2(n1130), .ZN(n1124) );
NAND2_X1 U812 ( .A1(G953), .A2(n1122), .ZN(n1123) );
NOR2_X1 U813 ( .A1(n1135), .A2(n1136), .ZN(G66) );
XNOR2_X1 U814 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(n1135) );
XOR2_X1 U817 ( .A(KEYINPUT56), .B(G952), .Z(n1142) );
NOR2_X1 U818 ( .A1(n1143), .A2(n1144), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1145), .A2(n1094), .A3(n1146), .ZN(n1144) );
NOR4_X1 U820 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1140), .ZN(n1146) );
NOR2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1145) );
NOR2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(n1151) );
INV_X1 U823 ( .A(n1152), .ZN(n1148) );
INV_X1 U824 ( .A(n1153), .ZN(n1147) );
NOR2_X1 U825 ( .A1(n1040), .A2(n1149), .ZN(n1150) );
NOR2_X1 U826 ( .A1(n1143), .A2(n1154), .ZN(G60) );
NOR3_X1 U827 ( .A1(n1088), .A2(n1155), .A3(n1156), .ZN(n1154) );
NOR3_X1 U828 ( .A1(n1157), .A2(n1087), .A3(n1140), .ZN(n1156) );
INV_X1 U829 ( .A(n1158), .ZN(n1157) );
NOR2_X1 U830 ( .A1(n1159), .A2(n1158), .ZN(n1155) );
NOR2_X1 U831 ( .A1(n1040), .A2(n1087), .ZN(n1159) );
XOR2_X1 U832 ( .A(n1160), .B(G104), .Z(G6) );
NAND2_X1 U833 ( .A1(KEYINPUT20), .A2(n1161), .ZN(n1160) );
NAND3_X1 U834 ( .A1(n1162), .A2(n1046), .A3(n1163), .ZN(n1161) );
NOR2_X1 U835 ( .A1(n1143), .A2(n1164), .ZN(G57) );
XOR2_X1 U836 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U838 ( .A1(n1169), .A2(n1140), .ZN(n1168) );
INV_X1 U839 ( .A(G472), .ZN(n1169) );
NOR2_X1 U840 ( .A1(n1170), .A2(n1171), .ZN(n1167) );
NOR2_X1 U841 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NOR2_X1 U842 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
INV_X1 U843 ( .A(KEYINPUT5), .ZN(n1175) );
NOR2_X1 U844 ( .A1(KEYINPUT2), .A2(n1176), .ZN(n1174) );
INV_X1 U845 ( .A(n1177), .ZN(n1176) );
NOR2_X1 U846 ( .A1(n1178), .A2(n1177), .ZN(n1170) );
XNOR2_X1 U847 ( .A(n1179), .B(KEYINPUT22), .ZN(n1177) );
NOR2_X1 U848 ( .A1(n1180), .A2(KEYINPUT2), .ZN(n1178) );
AND2_X1 U849 ( .A1(n1173), .A2(KEYINPUT5), .ZN(n1180) );
NOR2_X1 U850 ( .A1(n1143), .A2(n1181), .ZN(G54) );
XOR2_X1 U851 ( .A(n1182), .B(n1183), .Z(n1181) );
XOR2_X1 U852 ( .A(n1184), .B(n1185), .Z(n1183) );
NOR2_X1 U853 ( .A1(n1186), .A2(n1140), .ZN(n1184) );
INV_X1 U854 ( .A(G469), .ZN(n1186) );
XOR2_X1 U855 ( .A(KEYINPUT39), .B(n1187), .Z(n1182) );
NOR2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U857 ( .A1(n1143), .A2(n1190), .ZN(G51) );
XOR2_X1 U858 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U859 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U860 ( .A1(n1195), .A2(n1140), .ZN(n1193) );
OR2_X1 U861 ( .A1(n1196), .A2(n1040), .ZN(n1140) );
NOR2_X1 U862 ( .A1(n1118), .A2(n1110), .ZN(n1040) );
NAND4_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1110) );
NOR3_X1 U864 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
NAND2_X1 U865 ( .A1(n1052), .A2(n1204), .ZN(n1199) );
NAND2_X1 U866 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
NAND2_X1 U867 ( .A1(n1207), .A2(n1078), .ZN(n1206) );
OR2_X1 U868 ( .A1(n1163), .A2(n1208), .ZN(n1078) );
XNOR2_X1 U869 ( .A(n1209), .B(KEYINPUT35), .ZN(n1205) );
NAND4_X1 U870 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1118) );
AND4_X1 U871 ( .A1(n1036), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1213) );
NAND3_X1 U872 ( .A1(n1162), .A2(n1046), .A3(n1208), .ZN(n1036) );
NOR2_X1 U873 ( .A1(n1217), .A2(n1218), .ZN(n1212) );
NAND4_X1 U874 ( .A1(KEYINPUT32), .A2(n1219), .A3(n1220), .A4(n1062), .ZN(n1211) );
NOR2_X1 U875 ( .A1(n1221), .A2(n1070), .ZN(n1220) );
NAND2_X1 U876 ( .A1(n1162), .A2(n1222), .ZN(n1210) );
NAND2_X1 U877 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NAND2_X1 U878 ( .A1(n1163), .A2(n1225), .ZN(n1224) );
XOR2_X1 U879 ( .A(KEYINPUT27), .B(n1046), .Z(n1225) );
OR2_X1 U880 ( .A1(n1226), .A2(KEYINPUT32), .ZN(n1223) );
INV_X1 U881 ( .A(G210), .ZN(n1195) );
NOR2_X1 U882 ( .A1(n1141), .A2(G952), .ZN(n1143) );
XOR2_X1 U883 ( .A(KEYINPUT61), .B(n1080), .Z(n1141) );
XNOR2_X1 U884 ( .A(n1227), .B(n1197), .ZN(G48) );
NAND3_X1 U885 ( .A1(n1163), .A2(n1228), .A3(n1229), .ZN(n1197) );
NAND2_X1 U886 ( .A1(KEYINPUT19), .A2(n1230), .ZN(n1227) );
XNOR2_X1 U887 ( .A(G143), .B(n1198), .ZN(G45) );
NAND2_X1 U888 ( .A1(n1207), .A2(n1231), .ZN(n1198) );
XNOR2_X1 U889 ( .A(G140), .B(n1232), .ZN(G42) );
NAND2_X1 U890 ( .A1(n1209), .A2(n1052), .ZN(n1232) );
AND2_X1 U891 ( .A1(n1233), .A2(n1234), .ZN(n1209) );
XNOR2_X1 U892 ( .A(n1201), .B(n1235), .ZN(G39) );
NAND2_X1 U893 ( .A1(KEYINPUT6), .A2(G137), .ZN(n1235) );
AND3_X1 U894 ( .A1(n1229), .A2(n1045), .A3(n1052), .ZN(n1201) );
XOR2_X1 U895 ( .A(n1236), .B(n1237), .Z(G36) );
XNOR2_X1 U896 ( .A(G134), .B(KEYINPUT49), .ZN(n1237) );
NAND4_X1 U897 ( .A1(KEYINPUT31), .A2(n1207), .A3(n1052), .A4(n1208), .ZN(n1236) );
INV_X1 U898 ( .A(n1238), .ZN(n1207) );
XOR2_X1 U899 ( .A(n1239), .B(n1240), .Z(G33) );
NAND2_X1 U900 ( .A1(n1052), .A2(n1241), .ZN(n1240) );
XOR2_X1 U901 ( .A(KEYINPUT50), .B(n1242), .Z(n1241) );
NOR2_X1 U902 ( .A1(n1243), .A2(n1238), .ZN(n1242) );
NAND3_X1 U903 ( .A1(n1234), .A2(n1244), .A3(n1245), .ZN(n1238) );
NOR2_X1 U904 ( .A1(n1246), .A2(n1050), .ZN(n1052) );
INV_X1 U905 ( .A(n1051), .ZN(n1246) );
XOR2_X1 U906 ( .A(G128), .B(n1203), .Z(G30) );
AND3_X1 U907 ( .A1(n1208), .A2(n1228), .A3(n1229), .ZN(n1203) );
AND4_X1 U908 ( .A1(n1247), .A2(n1234), .A3(n1248), .A4(n1244), .ZN(n1229) );
XOR2_X1 U909 ( .A(G101), .B(n1249), .Z(G3) );
AND2_X1 U910 ( .A1(n1162), .A2(n1062), .ZN(n1249) );
INV_X1 U911 ( .A(n1226), .ZN(n1062) );
NAND2_X1 U912 ( .A1(n1245), .A2(n1045), .ZN(n1226) );
XOR2_X1 U913 ( .A(G125), .B(n1202), .Z(G27) );
AND3_X1 U914 ( .A1(n1074), .A2(n1228), .A3(n1233), .ZN(n1202) );
AND4_X1 U915 ( .A1(n1247), .A2(n1163), .A3(n1058), .A4(n1244), .ZN(n1233) );
NAND2_X1 U916 ( .A1(n1063), .A2(n1250), .ZN(n1244) );
NAND3_X1 U917 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1250) );
XOR2_X1 U918 ( .A(n1080), .B(KEYINPUT42), .Z(n1253) );
INV_X1 U919 ( .A(G900), .ZN(n1252) );
INV_X1 U920 ( .A(n1064), .ZN(n1074) );
XOR2_X1 U921 ( .A(n1254), .B(n1255), .Z(G24) );
NAND2_X1 U922 ( .A1(KEYINPUT63), .A2(n1218), .ZN(n1255) );
AND3_X1 U923 ( .A1(n1256), .A2(n1046), .A3(n1231), .ZN(n1218) );
AND3_X1 U924 ( .A1(n1228), .A2(n1257), .A3(n1258), .ZN(n1231) );
NOR2_X1 U925 ( .A1(n1089), .A2(n1247), .ZN(n1046) );
XNOR2_X1 U926 ( .A(n1217), .B(n1259), .ZN(G21) );
NAND2_X1 U927 ( .A1(KEYINPUT40), .A2(G119), .ZN(n1259) );
AND4_X1 U928 ( .A1(n1256), .A2(n1059), .A3(n1248), .A4(n1228), .ZN(n1217) );
XOR2_X1 U929 ( .A(n1260), .B(n1216), .Z(G18) );
NAND4_X1 U930 ( .A1(n1256), .A2(n1245), .A3(n1208), .A4(n1228), .ZN(n1216) );
INV_X1 U931 ( .A(n1048), .ZN(n1228) );
XOR2_X1 U932 ( .A(n1221), .B(KEYINPUT26), .Z(n1048) );
NOR2_X1 U933 ( .A1(n1257), .A2(n1261), .ZN(n1208) );
XNOR2_X1 U934 ( .A(G113), .B(n1215), .ZN(G15) );
NAND4_X1 U935 ( .A1(n1163), .A2(n1256), .A3(n1245), .A4(n1262), .ZN(n1215) );
NOR2_X1 U936 ( .A1(n1263), .A2(n1247), .ZN(n1245) );
INV_X1 U937 ( .A(n1248), .ZN(n1263) );
XOR2_X1 U938 ( .A(n1089), .B(KEYINPUT38), .Z(n1248) );
INV_X1 U939 ( .A(n1058), .ZN(n1089) );
NOR2_X1 U940 ( .A1(n1064), .A2(n1219), .ZN(n1256) );
NAND2_X1 U941 ( .A1(n1073), .A2(n1264), .ZN(n1064) );
INV_X1 U942 ( .A(n1243), .ZN(n1163) );
NAND2_X1 U943 ( .A1(n1261), .A2(n1257), .ZN(n1243) );
INV_X1 U944 ( .A(n1258), .ZN(n1261) );
XNOR2_X1 U945 ( .A(G110), .B(n1214), .ZN(G12) );
NAND3_X1 U946 ( .A1(n1058), .A2(n1162), .A3(n1059), .ZN(n1214) );
AND2_X1 U947 ( .A1(n1045), .A2(n1247), .ZN(n1059) );
XNOR2_X1 U948 ( .A(n1086), .B(KEYINPUT8), .ZN(n1247) );
XOR2_X1 U949 ( .A(n1265), .B(n1139), .Z(n1086) );
NAND2_X1 U950 ( .A1(G217), .A2(n1266), .ZN(n1139) );
NAND2_X1 U951 ( .A1(n1196), .A2(n1137), .ZN(n1265) );
NAND3_X1 U952 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1137) );
NAND2_X1 U953 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
NAND2_X1 U954 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XOR2_X1 U955 ( .A(KEYINPUT3), .B(n1274), .Z(n1272) );
INV_X1 U956 ( .A(n1275), .ZN(n1270) );
NAND3_X1 U957 ( .A1(n1274), .A2(n1275), .A3(n1273), .ZN(n1268) );
NAND3_X1 U958 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1275) );
NAND2_X1 U959 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U960 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND3_X1 U961 ( .A1(n1283), .A2(n1282), .A3(n1284), .ZN(n1277) );
INV_X1 U962 ( .A(n1281), .ZN(n1283) );
XOR2_X1 U963 ( .A(n1279), .B(n1285), .Z(n1281) );
XOR2_X1 U964 ( .A(KEYINPUT23), .B(KEYINPUT0), .Z(n1285) );
XNOR2_X1 U965 ( .A(G125), .B(n1286), .ZN(n1279) );
XOR2_X1 U966 ( .A(G146), .B(G140), .Z(n1286) );
OR2_X1 U967 ( .A1(n1284), .A2(n1282), .ZN(n1276) );
XNOR2_X1 U968 ( .A(n1287), .B(n1288), .ZN(n1282) );
XOR2_X1 U969 ( .A(G128), .B(G119), .Z(n1288) );
NAND2_X1 U970 ( .A1(KEYINPUT25), .A2(G110), .ZN(n1287) );
INV_X1 U971 ( .A(KEYINPUT52), .ZN(n1284) );
OR2_X1 U972 ( .A1(n1273), .A2(n1274), .ZN(n1267) );
XNOR2_X1 U973 ( .A(n1289), .B(G137), .ZN(n1274) );
NAND3_X1 U974 ( .A1(G234), .A2(n1080), .A3(G221), .ZN(n1289) );
INV_X1 U975 ( .A(KEYINPUT46), .ZN(n1273) );
NOR2_X1 U976 ( .A1(n1257), .A2(n1258), .ZN(n1045) );
XOR2_X1 U977 ( .A(n1290), .B(n1094), .Z(n1258) );
AND2_X1 U978 ( .A1(n1291), .A2(n1196), .ZN(n1094) );
NAND2_X1 U979 ( .A1(n1153), .A2(n1152), .ZN(n1291) );
NAND4_X1 U980 ( .A1(n1292), .A2(G217), .A3(n1293), .A4(n1080), .ZN(n1152) );
XOR2_X1 U981 ( .A(n1294), .B(n1295), .Z(n1293) );
NAND2_X1 U982 ( .A1(n1296), .A2(n1297), .ZN(n1153) );
NAND3_X1 U983 ( .A1(n1292), .A2(n1080), .A3(G217), .ZN(n1297) );
XNOR2_X1 U984 ( .A(G234), .B(KEYINPUT34), .ZN(n1292) );
XOR2_X1 U985 ( .A(n1298), .B(n1295), .Z(n1296) );
XNOR2_X1 U986 ( .A(n1299), .B(G122), .ZN(n1295) );
NAND2_X1 U987 ( .A1(KEYINPUT4), .A2(n1260), .ZN(n1299) );
INV_X1 U988 ( .A(G116), .ZN(n1260) );
INV_X1 U989 ( .A(n1294), .ZN(n1298) );
NAND2_X1 U990 ( .A1(KEYINPUT24), .A2(n1096), .ZN(n1290) );
XOR2_X1 U991 ( .A(n1149), .B(KEYINPUT10), .Z(n1096) );
INV_X1 U992 ( .A(G478), .ZN(n1149) );
XOR2_X1 U993 ( .A(n1088), .B(n1300), .Z(n1257) );
NOR2_X1 U994 ( .A1(KEYINPUT48), .A2(n1087), .ZN(n1300) );
INV_X1 U995 ( .A(G475), .ZN(n1087) );
NOR2_X1 U996 ( .A1(n1158), .A2(G902), .ZN(n1088) );
XOR2_X1 U997 ( .A(n1301), .B(n1302), .Z(n1158) );
XOR2_X1 U998 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U999 ( .A(n1305), .B(G104), .Z(n1304) );
NAND2_X1 U1000 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XNOR2_X1 U1001 ( .A(G214), .B(KEYINPUT15), .ZN(n1306) );
NAND2_X1 U1002 ( .A1(n1308), .A2(n1309), .ZN(n1303) );
NAND2_X1 U1003 ( .A1(n1310), .A2(n1230), .ZN(n1309) );
XOR2_X1 U1004 ( .A(KEYINPUT30), .B(n1311), .Z(n1308) );
NOR2_X1 U1005 ( .A1(n1310), .A2(n1230), .ZN(n1311) );
XOR2_X1 U1006 ( .A(G140), .B(n1312), .Z(n1310) );
NOR2_X1 U1007 ( .A1(G125), .A2(KEYINPUT28), .ZN(n1312) );
XOR2_X1 U1008 ( .A(n1313), .B(n1314), .Z(n1301) );
XOR2_X1 U1009 ( .A(G143), .B(G131), .Z(n1314) );
XOR2_X1 U1010 ( .A(G113), .B(n1254), .Z(n1313) );
NOR3_X1 U1011 ( .A1(n1221), .A2(n1219), .A3(n1070), .ZN(n1162) );
INV_X1 U1012 ( .A(n1234), .ZN(n1070) );
NOR2_X1 U1013 ( .A1(n1073), .A2(n1072), .ZN(n1234) );
INV_X1 U1014 ( .A(n1264), .ZN(n1072) );
NAND2_X1 U1015 ( .A1(n1315), .A2(n1266), .ZN(n1264) );
NAND2_X1 U1016 ( .A1(G234), .A2(n1196), .ZN(n1266) );
XOR2_X1 U1017 ( .A(KEYINPUT11), .B(G221), .Z(n1315) );
XOR2_X1 U1018 ( .A(n1316), .B(G469), .Z(n1073) );
NAND2_X1 U1019 ( .A1(n1317), .A2(n1196), .ZN(n1316) );
XOR2_X1 U1020 ( .A(n1318), .B(n1319), .Z(n1317) );
NAND2_X1 U1021 ( .A1(KEYINPUT62), .A2(n1185), .ZN(n1319) );
XNOR2_X1 U1022 ( .A(n1320), .B(n1321), .ZN(n1185) );
XOR2_X1 U1023 ( .A(G101), .B(n1322), .Z(n1321) );
XOR2_X1 U1024 ( .A(KEYINPUT44), .B(G104), .Z(n1322) );
XOR2_X1 U1025 ( .A(n1106), .B(n1294), .Z(n1320) );
XOR2_X1 U1026 ( .A(n1107), .B(G107), .Z(n1294) );
XOR2_X1 U1027 ( .A(G128), .B(n1323), .Z(n1107) );
XOR2_X1 U1028 ( .A(G143), .B(G134), .Z(n1323) );
XNOR2_X1 U1029 ( .A(n1324), .B(n1325), .ZN(n1106) );
XOR2_X1 U1030 ( .A(KEYINPUT57), .B(n1326), .Z(n1325) );
INV_X1 U1031 ( .A(n1327), .ZN(n1326) );
NAND3_X1 U1032 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1318) );
INV_X1 U1033 ( .A(n1188), .ZN(n1330) );
NOR2_X1 U1034 ( .A1(n1331), .A2(n1332), .ZN(n1188) );
NAND2_X1 U1035 ( .A1(n1189), .A2(KEYINPUT33), .ZN(n1329) );
AND2_X1 U1036 ( .A1(n1332), .A2(n1331), .ZN(n1189) );
NAND2_X1 U1037 ( .A1(G227), .A2(n1080), .ZN(n1331) );
OR2_X1 U1038 ( .A1(n1332), .A2(KEYINPUT33), .ZN(n1328) );
XOR2_X1 U1039 ( .A(G110), .B(G140), .Z(n1332) );
AND2_X1 U1040 ( .A1(n1333), .A2(n1063), .ZN(n1219) );
NAND3_X1 U1041 ( .A1(n1334), .A2(n1080), .A3(G952), .ZN(n1063) );
INV_X1 U1042 ( .A(G953), .ZN(n1080) );
NAND3_X1 U1043 ( .A1(n1251), .A2(n1122), .A3(G953), .ZN(n1333) );
INV_X1 U1044 ( .A(G898), .ZN(n1122) );
AND2_X1 U1045 ( .A1(n1335), .A2(n1334), .ZN(n1251) );
NAND2_X1 U1046 ( .A1(G237), .A2(G234), .ZN(n1334) );
XOR2_X1 U1047 ( .A(KEYINPUT55), .B(G902), .Z(n1335) );
INV_X1 U1048 ( .A(n1262), .ZN(n1221) );
NOR2_X1 U1049 ( .A1(n1051), .A2(n1050), .ZN(n1262) );
AND2_X1 U1050 ( .A1(G214), .A2(n1336), .ZN(n1050) );
XOR2_X1 U1051 ( .A(n1337), .B(n1338), .Z(n1051) );
AND2_X1 U1052 ( .A1(n1336), .A2(G210), .ZN(n1338) );
NAND2_X1 U1053 ( .A1(n1339), .A2(n1196), .ZN(n1336) );
XOR2_X1 U1054 ( .A(KEYINPUT12), .B(G237), .Z(n1339) );
NAND2_X1 U1055 ( .A1(n1340), .A2(n1196), .ZN(n1337) );
XOR2_X1 U1056 ( .A(n1341), .B(n1342), .Z(n1340) );
INV_X1 U1057 ( .A(n1191), .ZN(n1342) );
XOR2_X1 U1058 ( .A(n1343), .B(n1344), .Z(n1191) );
XNOR2_X1 U1059 ( .A(n1129), .B(n1130), .ZN(n1344) );
XNOR2_X1 U1060 ( .A(n1345), .B(n1346), .ZN(n1130) );
XOR2_X1 U1061 ( .A(G101), .B(n1347), .Z(n1346) );
NOR2_X1 U1062 ( .A1(KEYINPUT47), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1063 ( .A(n1035), .B(G104), .Z(n1348) );
INV_X1 U1064 ( .A(G107), .ZN(n1035) );
NAND3_X1 U1065 ( .A1(n1349), .A2(n1350), .A3(n1351), .ZN(n1129) );
OR2_X1 U1066 ( .A1(n1254), .A2(n1352), .ZN(n1351) );
NAND3_X1 U1067 ( .A1(n1352), .A2(n1254), .A3(KEYINPUT58), .ZN(n1350) );
INV_X1 U1068 ( .A(G122), .ZN(n1254) );
NOR2_X1 U1069 ( .A1(G110), .A2(KEYINPUT17), .ZN(n1352) );
NAND2_X1 U1070 ( .A1(G110), .A2(n1353), .ZN(n1349) );
INV_X1 U1071 ( .A(KEYINPUT58), .ZN(n1353) );
XOR2_X1 U1072 ( .A(n1354), .B(n1355), .Z(n1343) );
XNOR2_X1 U1073 ( .A(G125), .B(KEYINPUT7), .ZN(n1354) );
XOR2_X1 U1074 ( .A(n1356), .B(KEYINPUT13), .Z(n1341) );
NAND2_X1 U1075 ( .A1(KEYINPUT18), .A2(n1194), .ZN(n1356) );
NOR2_X1 U1076 ( .A1(n1121), .A2(G953), .ZN(n1194) );
INV_X1 U1077 ( .A(G224), .ZN(n1121) );
XOR2_X1 U1078 ( .A(n1357), .B(G472), .Z(n1058) );
NAND2_X1 U1079 ( .A1(n1358), .A2(n1196), .ZN(n1357) );
INV_X1 U1080 ( .A(G902), .ZN(n1196) );
XOR2_X1 U1081 ( .A(n1359), .B(n1165), .Z(n1358) );
XNOR2_X1 U1082 ( .A(n1360), .B(G101), .ZN(n1165) );
NAND2_X1 U1083 ( .A1(G210), .A2(n1307), .ZN(n1360) );
NOR2_X1 U1084 ( .A1(G953), .A2(G237), .ZN(n1307) );
XNOR2_X1 U1085 ( .A(n1173), .B(n1179), .ZN(n1359) );
XNOR2_X1 U1086 ( .A(n1327), .B(n1361), .ZN(n1179) );
XOR2_X1 U1087 ( .A(G134), .B(n1355), .Z(n1361) );
AND2_X1 U1088 ( .A1(n1362), .A2(n1363), .ZN(n1355) );
NAND2_X1 U1089 ( .A1(n1364), .A2(G128), .ZN(n1363) );
XOR2_X1 U1090 ( .A(KEYINPUT29), .B(n1365), .Z(n1362) );
NOR2_X1 U1091 ( .A1(G128), .A2(n1364), .ZN(n1365) );
XNOR2_X1 U1092 ( .A(G143), .B(n1324), .ZN(n1364) );
XNOR2_X1 U1093 ( .A(n1230), .B(KEYINPUT51), .ZN(n1324) );
INV_X1 U1094 ( .A(G146), .ZN(n1230) );
XOR2_X1 U1095 ( .A(n1239), .B(G137), .Z(n1327) );
INV_X1 U1096 ( .A(G131), .ZN(n1239) );
XNOR2_X1 U1097 ( .A(n1345), .B(KEYINPUT59), .ZN(n1173) );
XNOR2_X1 U1098 ( .A(G113), .B(n1366), .ZN(n1345) );
XOR2_X1 U1099 ( .A(G119), .B(G116), .Z(n1366) );
endmodule


