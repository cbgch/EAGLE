//Key = 11101001001100110111110011100010001000011001000100101110101001111110010010000001101100
module c3540 ( G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, 
        G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, 
        G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, 
        G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, 
        G1698, G2897, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, G353, G355, G361, G358, G351, G372, 
        G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, 
        G407, G409, G405, G402 );
  input G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
         G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
         G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
         G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330,
         G343, G1698, G2897, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
         G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire   n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260;

  NOR3_X2 U1667 ( .A1(n2918), .A2(n2919), .A3(n2920), .ZN(n2567) );
  NOR3_X2 U1668 ( .A1(n2921), .A2(n2922), .A3(n2920), .ZN(n2518) );
  XNOR2_X2 U1669 ( .A(keyinput15), .B(G200), .ZN(n2922) );
  XNOR2_X2 U1670 ( .A(keyinput7), .B(G77), .ZN(n2538) );
  NOR3_X2 U1671 ( .A1(n2918), .A2(n2921), .A3(n2920), .ZN(n2573) );
  NAND3_X1 U1672 ( .A1(n2431), .A2(G407), .A3(G213), .ZN(G409) );
  OR3_X1 U1673 ( .A1(n2432), .A2(G343), .A3(n2433), .ZN(n2431) );
  NAND2_X1 U1674 ( .A1(n2434), .A2(n2435), .ZN(G407) );
  NOR4_X1 U1675 ( .A1(n2436), .A2(n2432), .A3(n2437), .A4(n2438), .ZN(n2435) );
  NOR4_X1 U1676 ( .A1(n2439), .A2(n2433), .A3(n2440), .A4(n2441), .ZN(n2434) );
  XOR2_X1 U1677 ( .A(n2442), .B(n2443), .Z(G405) );
  XOR2_X1 U1678 ( .A(n2444), .B(n2445), .Z(n2443) );
  NOR2_X1 U1679 ( .A1(n2446), .A2(n2447), .ZN(n2445) );
  NAND2_X1 U1680 ( .A1(n2448), .A2(n2449), .ZN(n2442) );
  NAND2_X1 U1681 ( .A1(G375), .A2(n2450), .ZN(n2449) );
  NAND2_X1 U1682 ( .A1(G2897), .A2(n2446), .ZN(n2448) );
  INV_X1 U1683 ( .A(n2450), .ZN(n2446) );
  NAND2_X1 U1684 ( .A1(G213), .A2(n2451), .ZN(n2450) );
  XOR2_X1 U1685 ( .A(n2447), .B(n2452), .Z(G402) );
  XNOR2_X1 U1686 ( .A(n2444), .B(G375), .ZN(n2452) );
  XOR2_X1 U1687 ( .A(n2453), .B(n2454), .Z(n2444) );
  XOR2_X1 U1688 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR2_X1 U1689 ( .A(n2457), .B(n2458), .Z(n2456) );
  XOR2_X1 U1690 ( .A(n2459), .B(n2460), .Z(n2453) );
  XNOR2_X1 U1691 ( .A(n2461), .B(n2462), .ZN(n2460) );
  NOR2_X1 U1692 ( .A1(n2463), .A2(n2457), .ZN(G396) );
  XNOR2_X1 U1693 ( .A(n2436), .B(keyinput73), .ZN(n2457) );
  INV_X1 U1694 ( .A(n2436), .ZN(n2463) );
  NAND3_X1 U1695 ( .A1(n2464), .A2(n2465), .A3(n2466), .ZN(n2436) );
  NAND2_X1 U1696 ( .A1(n2467), .A2(n2468), .ZN(n2466) );
  INV_X1 U1697 ( .A(keyinput72), .ZN(n2468) );
  NAND3_X1 U1698 ( .A1(n2469), .A2(n2470), .A3(n2471), .ZN(n2467) );
  NAND4_X1 U1699 ( .A1(n2472), .A2(n2473), .A3(n2474), .A4(n2475), .ZN(n2465) );
  NOR2_X1 U1700 ( .A1(n2476), .A2(n2477), .ZN(n2475) );
  NOR2_X1 U1701 ( .A1(n2478), .A2(n2479), .ZN(n2476) );
  NAND2_X1 U1702 ( .A1(n2480), .A2(n2481), .ZN(n2474) );
  NAND3_X1 U1703 ( .A1(n2482), .A2(n2483), .A3(n2484), .ZN(n2481) );
  NAND2_X1 U1704 ( .A1(n2485), .A2(G355), .ZN(n2484) );
  NAND3_X1 U1705 ( .A1(n2486), .A2(n2487), .A3(n2488), .ZN(n2483) );
  NAND2_X1 U1706 ( .A1(n2489), .A2(n2490), .ZN(n2482) );
  NAND2_X1 U1707 ( .A1(n2491), .A2(n2492), .ZN(n2489) );
  NAND2_X1 U1708 ( .A1(n2493), .A2(n2494), .ZN(n2492) );
  NAND2_X1 U1709 ( .A1(n2495), .A2(G45), .ZN(n2491) );
  NAND4_X1 U1710 ( .A1(n2496), .A2(n2497), .A3(n2498), .A4(n2499), .ZN(n2473) );
  NOR4_X1 U1711 ( .A1(n2500), .A2(n2501), .A3(n2502), .A4(n2503), .ZN(n2499) );
  AND2_X1 U1712 ( .A1(n2504), .A2(G326), .ZN(n2502) );
  NOR2_X1 U1713 ( .A1(n2505), .A2(n2506), .ZN(n2501) );
  NOR2_X1 U1714 ( .A1(n2507), .A2(n2508), .ZN(n2500) );
  NOR3_X1 U1715 ( .A1(n2509), .A2(n2510), .A3(n2511), .ZN(n2498) );
  NOR2_X1 U1716 ( .A1(n2512), .A2(n2513), .ZN(n2511) );
  NOR2_X1 U1717 ( .A1(n2514), .A2(n2515), .ZN(n2510) );
  NOR2_X1 U1718 ( .A1(n2516), .A2(n2517), .ZN(n2509) );
  NAND2_X1 U1719 ( .A1(G311), .A2(n2518), .ZN(n2497) );
  NAND2_X1 U1720 ( .A1(G329), .A2(n2519), .ZN(n2496) );
  NAND4_X1 U1721 ( .A1(n2520), .A2(n2521), .A3(n2522), .A4(n2523), .ZN(n2472) );
  NOR4_X1 U1722 ( .A1(n2524), .A2(n2525), .A3(n2526), .A4(n2527), .ZN(n2523) );
  NOR2_X1 U1723 ( .A1(n2528), .A2(n2529), .ZN(n2526) );
  NOR2_X1 U1724 ( .A1(n2530), .A2(n2512), .ZN(n2524) );
  NOR3_X1 U1725 ( .A1(n2531), .A2(n2532), .A3(n2533), .ZN(n2522) );
  NOR2_X1 U1726 ( .A1(n2534), .A2(n2535), .ZN(n2533) );
  NOR2_X1 U1727 ( .A1(n2536), .A2(n2516), .ZN(n2532) );
  NOR2_X1 U1728 ( .A1(n2537), .A2(n2514), .ZN(n2531) );
  NAND2_X1 U1729 ( .A1(n2538), .A2(n2518), .ZN(n2521) );
  NAND2_X1 U1730 ( .A1(n2539), .A2(n2540), .ZN(n2520) );
  NAND3_X1 U1731 ( .A1(n2469), .A2(n2470), .A3(n2541), .ZN(n2464) );
  NAND2_X1 U1732 ( .A1(n2542), .A2(n2543), .ZN(n2541) );
  NAND2_X1 U1733 ( .A1(keyinput72), .A2(n2471), .ZN(n2543) );
  NAND2_X1 U1734 ( .A1(n2544), .A2(n2545), .ZN(n2469) );
  NOR2_X1 U1735 ( .A1(n2546), .A2(n2455), .ZN(G393) );
  XOR2_X1 U1736 ( .A(n2546), .B(keyinput81), .Z(n2455) );
  INV_X1 U1737 ( .A(n2437), .ZN(n2546) );
  NAND3_X1 U1738 ( .A1(n2547), .A2(n2548), .A3(n2549), .ZN(n2437) );
  XOR2_X1 U1739 ( .A(n2550), .B(keyinput75), .Z(n2549) );
  NAND2_X1 U1740 ( .A1(n2551), .A2(n2471), .ZN(n2550) );
  NAND4_X1 U1741 ( .A1(n2552), .A2(n2553), .A3(n2554), .A4(n2555), .ZN(n2548) );
  NOR3_X1 U1742 ( .A1(n2556), .A2(n2557), .A3(n2558), .ZN(n2555) );
  NOR4_X1 U1743 ( .A1(n2559), .A2(n2560), .A3(n2561), .A4(n2562), .ZN(n2558) );
  NOR2_X1 U1744 ( .A1(n2514), .A2(n2517), .ZN(n2562) );
  NOR2_X1 U1745 ( .A1(n2507), .A2(n2513), .ZN(n2561) );
  NAND3_X1 U1746 ( .A1(n2563), .A2(n2564), .A3(n2565), .ZN(n2560) );
  NAND2_X1 U1747 ( .A1(G326), .A2(n2519), .ZN(n2565) );
  NAND2_X1 U1748 ( .A1(n2566), .A2(n2567), .ZN(n2564) );
  NAND2_X1 U1749 ( .A1(G322), .A2(n2504), .ZN(n2563) );
  NAND4_X1 U1750 ( .A1(n2568), .A2(n2569), .A3(n2570), .A4(n2571), .ZN(n2559) );
  NAND2_X1 U1751 ( .A1(G283), .A2(n2572), .ZN(n2571) );
  NAND2_X1 U1752 ( .A1(G311), .A2(n2573), .ZN(n2570) );
  NAND2_X1 U1753 ( .A1(G303), .A2(n2518), .ZN(n2569) );
  NOR4_X1 U1754 ( .A1(n2574), .A2(n2575), .A3(n2576), .A4(n2577), .ZN(n2557) );
  NOR2_X1 U1755 ( .A1(n2514), .A2(n2535), .ZN(n2577) );
  NAND3_X1 U1756 ( .A1(n2578), .A2(n2579), .A3(n2580), .ZN(n2575) );
  NAND2_X1 U1757 ( .A1(n2519), .A2(G150), .ZN(n2580) );
  NAND2_X1 U1758 ( .A1(G159), .A2(n2504), .ZN(n2578) );
  NAND4_X1 U1759 ( .A1(n2581), .A2(n2582), .A3(n2583), .A4(n2584), .ZN(n2574) );
  NAND2_X1 U1760 ( .A1(n2573), .A2(n2585), .ZN(n2583) );
  NAND2_X1 U1761 ( .A1(n2518), .A2(n2586), .ZN(n2582) );
  NOR3_X1 U1762 ( .A1(n2488), .A2(G45), .A3(n2587), .ZN(n2556) );
  NOR4_X1 U1763 ( .A1(n2588), .A2(n2537), .A3(n2589), .A4(n2590), .ZN(n2587) );
  NOR2_X1 U1764 ( .A1(n2536), .A2(n2591), .ZN(n2588) );
  NAND2_X1 U1765 ( .A1(n2592), .A2(n2593), .ZN(n2553) );
  XOR2_X1 U1766 ( .A(n2594), .B(n2595), .Z(n2593) );
  INV_X1 U1767 ( .A(n2478), .ZN(n2592) );
  NAND2_X1 U1768 ( .A1(n2480), .A2(n2596), .ZN(n2552) );
  NAND3_X1 U1769 ( .A1(n2597), .A2(n2598), .A3(n2599), .ZN(n2596) );
  NAND2_X1 U1770 ( .A1(n2485), .A2(n2590), .ZN(n2599) );
  INV_X1 U1771 ( .A(n2487), .ZN(n2485) );
  NAND3_X1 U1772 ( .A1(n2600), .A2(n2487), .A3(n2488), .ZN(n2598) );
  NAND3_X1 U1773 ( .A1(G45), .A2(n2601), .A3(n2490), .ZN(n2597) );
  INV_X1 U1774 ( .A(n2602), .ZN(n2480) );
  NAND2_X1 U1775 ( .A1(n2603), .A2(n2604), .ZN(n2547) );
  XOR2_X1 U1776 ( .A(n2605), .B(n2551), .Z(n2603) );
  NOR2_X1 U1777 ( .A1(n2606), .A2(n2459), .ZN(G390) );
  XOR2_X1 U1778 ( .A(n2438), .B(keyinput82), .Z(n2459) );
  INV_X1 U1779 ( .A(n2438), .ZN(n2606) );
  NAND3_X1 U1780 ( .A1(n2607), .A2(n2608), .A3(n2609), .ZN(n2438) );
  XOR2_X1 U1781 ( .A(n2610), .B(keyinput76), .Z(n2609) );
  NAND2_X1 U1782 ( .A1(n2611), .A2(n2471), .ZN(n2610) );
  NAND4_X1 U1783 ( .A1(n2612), .A2(n2487), .A3(n2613), .A4(n2614), .ZN(n2608) );
  NOR4_X1 U1784 ( .A1(n2615), .A2(n2616), .A3(n2617), .A4(n2477), .ZN(n2614) );
  NOR2_X1 U1785 ( .A1(n2618), .A2(n2478), .ZN(n2617) );
  NOR2_X1 U1786 ( .A1(n2488), .A2(n2619), .ZN(n2616) );
  NOR3_X1 U1787 ( .A1(n2490), .A2(n2620), .A3(n2602), .ZN(n2615) );
  NAND4_X1 U1788 ( .A1(n2621), .A2(n2622), .A3(n2623), .A4(n2624), .ZN(n2613) );
  NOR4_X1 U1789 ( .A1(n2625), .A2(n2525), .A3(n2626), .A4(n2503), .ZN(n2624) );
  NOR2_X1 U1790 ( .A1(n2529), .A2(n2515), .ZN(n2626) );
  INV_X1 U1791 ( .A(G322), .ZN(n2515) );
  NOR2_X1 U1792 ( .A1(n2505), .A2(n2600), .ZN(n2525) );
  NOR2_X1 U1793 ( .A1(n2512), .A2(n2486), .ZN(n2625) );
  NOR3_X1 U1794 ( .A1(n2627), .A2(n2628), .A3(n2629), .ZN(n2623) );
  NOR2_X1 U1795 ( .A1(n2534), .A2(n2517), .ZN(n2629) );
  NOR2_X1 U1796 ( .A1(n2516), .A2(n2508), .ZN(n2628) );
  INV_X1 U1797 ( .A(G303), .ZN(n2508) );
  NOR2_X1 U1798 ( .A1(n2514), .A2(n2630), .ZN(n2627) );
  NAND2_X1 U1799 ( .A1(G294), .A2(n2518), .ZN(n2622) );
  NAND2_X1 U1800 ( .A1(G283), .A2(n2539), .ZN(n2621) );
  NAND4_X1 U1801 ( .A1(n2631), .A2(n2632), .A3(n2633), .A4(n2634), .ZN(n2612) );
  NOR4_X1 U1802 ( .A1(n2635), .A2(n2636), .A3(n2637), .A4(n2527), .ZN(n2634) );
  NOR2_X1 U1803 ( .A1(n2638), .A2(n2529), .ZN(n2637) );
  NOR2_X1 U1804 ( .A1(n2639), .A2(n2505), .ZN(n2636) );
  NOR2_X1 U1805 ( .A1(n2512), .A2(n2591), .ZN(n2635) );
  NOR3_X1 U1806 ( .A1(n2640), .A2(n2641), .A3(n2642), .ZN(n2633) );
  NOR2_X1 U1807 ( .A1(n2534), .A2(n2643), .ZN(n2642) );
  NOR2_X1 U1808 ( .A1(n2516), .A2(n2535), .ZN(n2641) );
  NOR2_X1 U1809 ( .A1(n2514), .A2(n2528), .ZN(n2640) );
  NAND2_X1 U1810 ( .A1(n2518), .A2(n2585), .ZN(n2632) );
  NAND2_X1 U1811 ( .A1(n2539), .A2(n2586), .ZN(n2631) );
  NAND2_X1 U1812 ( .A1(n2644), .A2(n2604), .ZN(n2607) );
  XNOR2_X1 U1813 ( .A(n2611), .B(n2645), .ZN(n2644) );
  NAND2_X1 U1814 ( .A1(n2605), .A2(n2551), .ZN(n2645) );
  NOR2_X1 U1815 ( .A1(n2646), .A2(n2461), .ZN(G387) );
  XOR2_X1 U1816 ( .A(n2439), .B(keyinput80), .Z(n2461) );
  INV_X1 U1817 ( .A(n2439), .ZN(n2646) );
  NAND3_X1 U1818 ( .A1(n2647), .A2(n2648), .A3(n2649), .ZN(n2439) );
  XOR2_X1 U1819 ( .A(keyinput79), .B(n2650), .Z(n2649) );
  NOR2_X1 U1820 ( .A1(n2651), .A2(n2652), .ZN(n2650) );
  XOR2_X1 U1821 ( .A(n2653), .B(n2654), .Z(n2652) );
  NAND3_X1 U1822 ( .A1(n2604), .A2(n2655), .A3(n2656), .ZN(n2648) );
  XOR2_X1 U1823 ( .A(n2657), .B(n2654), .Z(n2656) );
  XNOR2_X1 U1824 ( .A(n2658), .B(n2659), .ZN(n2654) );
  NAND2_X1 U1825 ( .A1(n2660), .A2(n2661), .ZN(n2658) );
  OR2_X1 U1826 ( .A1(n2662), .A2(n2663), .ZN(n2661) );
  NAND2_X1 U1827 ( .A1(n2618), .A2(n2664), .ZN(n2660) );
  INV_X1 U1828 ( .A(n2653), .ZN(n2657) );
  NAND2_X1 U1829 ( .A1(n2605), .A2(n2665), .ZN(n2655) );
  NAND2_X1 U1830 ( .A1(n2611), .A2(n2551), .ZN(n2665) );
  XOR2_X1 U1831 ( .A(n2666), .B(n2470), .Z(n2551) );
  NAND2_X1 U1832 ( .A1(n2667), .A2(n2668), .ZN(n2666) );
  OR2_X1 U1833 ( .A1(n2669), .A2(n2670), .ZN(n2668) );
  AND3_X1 U1834 ( .A1(n2671), .A2(n2672), .A3(n2673), .ZN(n2611) );
  OR2_X1 U1835 ( .A1(n2618), .A2(G399), .ZN(n2673) );
  NAND2_X1 U1836 ( .A1(n2674), .A2(n2675), .ZN(G399) );
  NAND2_X1 U1837 ( .A1(n2676), .A2(n2669), .ZN(n2675) );
  OR3_X1 U1838 ( .A1(n2674), .A2(n2677), .A3(n2659), .ZN(n2672) );
  NOR2_X1 U1839 ( .A1(n2618), .A2(n2678), .ZN(n2677) );
  AND2_X1 U1840 ( .A1(n2676), .A2(n2669), .ZN(n2678) );
  NAND2_X1 U1841 ( .A1(n2659), .A2(n2674), .ZN(n2671) );
  XNOR2_X1 U1842 ( .A(n2664), .B(keyinput70), .ZN(n2674) );
  NAND2_X1 U1843 ( .A1(n2679), .A2(n2667), .ZN(n2664) );
  NAND2_X1 U1844 ( .A1(n2670), .A2(n2669), .ZN(n2667) );
  XNOR2_X1 U1845 ( .A(n2680), .B(keyinput59), .ZN(n2670) );
  NAND2_X1 U1846 ( .A1(n2681), .A2(n2682), .ZN(n2680) );
  NAND2_X1 U1847 ( .A1(n2683), .A2(n2682), .ZN(n2679) );
  XOR2_X1 U1848 ( .A(n2684), .B(keyinput32), .Z(n2683) );
  AND3_X1 U1849 ( .A1(n2618), .A2(n2669), .A3(n2676), .ZN(n2659) );
  INV_X1 U1850 ( .A(n2470), .ZN(n2676) );
  NAND2_X1 U1851 ( .A1(n2685), .A2(n2479), .ZN(n2470) );
  INV_X1 U1852 ( .A(n2545), .ZN(n2479) );
  XOR2_X1 U1853 ( .A(n2686), .B(n2687), .Z(n2545) );
  XOR2_X1 U1854 ( .A(keyinput64), .B(keyinput37), .Z(n2687) );
  XNOR2_X1 U1855 ( .A(n2688), .B(n2689), .ZN(n2686) );
  NAND2_X1 U1856 ( .A1(n2663), .A2(n2690), .ZN(n2688) );
  XNOR2_X1 U1857 ( .A(n2691), .B(keyinput69), .ZN(n2669) );
  NAND2_X1 U1858 ( .A1(n2692), .A2(n2693), .ZN(n2691) );
  NAND2_X1 U1859 ( .A1(n2694), .A2(n2695), .ZN(n2693) );
  XOR2_X1 U1860 ( .A(keyinput49), .B(n2594), .Z(n2695) );
  XNOR2_X1 U1861 ( .A(keyinput65), .B(n2595), .ZN(n2694) );
  XOR2_X1 U1862 ( .A(n2696), .B(keyinput67), .Z(n2692) );
  NAND2_X1 U1863 ( .A1(n2697), .A2(n2698), .ZN(n2696) );
  XOR2_X1 U1864 ( .A(keyinput65), .B(n2595), .Z(n2698) );
  XOR2_X1 U1865 ( .A(n2699), .B(keyinput63), .Z(n2595) );
  XNOR2_X1 U1866 ( .A(n2594), .B(keyinput49), .ZN(n2697) );
  XNOR2_X1 U1867 ( .A(n2700), .B(keyinput36), .ZN(n2594) );
  NAND2_X1 U1868 ( .A1(n2663), .A2(n2701), .ZN(n2700) );
  XNOR2_X1 U1869 ( .A(n2702), .B(n2703), .ZN(n2618) );
  NAND2_X1 U1870 ( .A1(n2663), .A2(n2704), .ZN(n2702) );
  NAND4_X1 U1871 ( .A1(n2705), .A2(n2487), .A3(n2706), .A4(n2707), .ZN(n2647) );
  NOR4_X1 U1872 ( .A1(n2708), .A2(n2709), .A3(n2710), .A4(n2477), .ZN(n2707) );
  NOR2_X1 U1873 ( .A1(n2653), .A2(n2478), .ZN(n2710) );
  XNOR2_X1 U1874 ( .A(n2711), .B(n2712), .ZN(n2653) );
  NAND2_X1 U1875 ( .A1(n2663), .A2(n2713), .ZN(n2711) );
  NOR2_X1 U1876 ( .A1(n2488), .A2(n2714), .ZN(n2709) );
  NOR3_X1 U1877 ( .A1(n2490), .A2(n2540), .A3(n2602), .ZN(n2708) );
  NAND2_X1 U1878 ( .A1(n2478), .A2(n2715), .ZN(n2602) );
  NAND2_X1 U1879 ( .A1(n2716), .A2(n2717), .ZN(n2478) );
  INV_X1 U1880 ( .A(n2488), .ZN(n2490) );
  NAND2_X1 U1881 ( .A1(n2718), .A2(n2719), .ZN(n2488) );
  NAND4_X1 U1882 ( .A1(n2720), .A2(n2721), .A3(n2722), .A4(n2723), .ZN(n2706) );
  NOR4_X1 U1883 ( .A1(n2724), .A2(n2725), .A3(n2726), .A4(n2503), .ZN(n2723) );
  NOR2_X1 U1884 ( .A1(n2529), .A2(n2517), .ZN(n2726) );
  INV_X1 U1885 ( .A(G317), .ZN(n2517) );
  NOR2_X1 U1886 ( .A1(n2512), .A2(n2600), .ZN(n2725) );
  NOR2_X1 U1887 ( .A1(n2507), .A2(n2486), .ZN(n2724) );
  NOR3_X1 U1888 ( .A1(n2727), .A2(n2728), .A3(n2729), .ZN(n2722) );
  INV_X1 U1889 ( .A(n2579), .ZN(n2729) );
  NAND2_X1 U1890 ( .A1(n2567), .A2(n2620), .ZN(n2579) );
  NOR2_X1 U1891 ( .A1(n2516), .A2(n2513), .ZN(n2728) );
  INV_X1 U1892 ( .A(G294), .ZN(n2513) );
  NOR2_X1 U1893 ( .A1(n2534), .A2(n2630), .ZN(n2727) );
  INV_X1 U1894 ( .A(G311), .ZN(n2630) );
  NAND2_X1 U1895 ( .A1(G303), .A2(n2730), .ZN(n2721) );
  NAND2_X1 U1896 ( .A1(G283), .A2(n2518), .ZN(n2720) );
  NAND2_X1 U1897 ( .A1(n2731), .A2(n2718), .ZN(n2487) );
  NAND4_X1 U1898 ( .A1(n2732), .A2(n2733), .A3(n2734), .A4(n2735), .ZN(n2705) );
  NOR4_X1 U1899 ( .A1(n2736), .A2(n2737), .A3(n2738), .A4(n2527), .ZN(n2735) );
  NOR2_X1 U1900 ( .A1(n2739), .A2(n2529), .ZN(n2738) );
  NOR2_X1 U1901 ( .A1(n2505), .A2(n2591), .ZN(n2737) );
  NOR2_X1 U1902 ( .A1(n2536), .A2(n2512), .ZN(n2736) );
  INV_X1 U1903 ( .A(n2572), .ZN(n2512) );
  NOR3_X1 U1904 ( .A1(n2740), .A2(n2741), .A3(n2742), .ZN(n2734) );
  NOR2_X1 U1905 ( .A1(n2638), .A2(n2534), .ZN(n2742) );
  NOR2_X1 U1906 ( .A1(n2516), .A2(n2528), .ZN(n2741) );
  NOR2_X1 U1907 ( .A1(n2514), .A2(n2643), .ZN(n2740) );
  NAND2_X1 U1908 ( .A1(n2589), .A2(n2518), .ZN(n2733) );
  NAND2_X1 U1909 ( .A1(n2539), .A2(n2585), .ZN(n2732) );
  INV_X1 U1910 ( .A(n2507), .ZN(n2539) );
  NOR2_X1 U1911 ( .A1(n2743), .A2(n2458), .ZN(G384) );
  XNOR2_X1 U1912 ( .A(n2440), .B(keyinput77), .ZN(n2458) );
  INV_X1 U1913 ( .A(n2440), .ZN(n2743) );
  NAND3_X1 U1914 ( .A1(n2744), .A2(n2745), .A3(n2746), .ZN(n2440) );
  XOR2_X1 U1915 ( .A(n2747), .B(keyinput74), .Z(n2746) );
  NAND2_X1 U1916 ( .A1(n2471), .A2(n2748), .ZN(n2747) );
  NAND3_X1 U1917 ( .A1(n2554), .A2(n2749), .A3(n2750), .ZN(n2745) );
  NOR3_X1 U1918 ( .A1(n2751), .A2(n2752), .A3(n2753), .ZN(n2750) );
  NOR4_X1 U1919 ( .A1(n2754), .A2(n2755), .A3(n2756), .A4(n2757), .ZN(n2753) );
  NOR2_X1 U1920 ( .A1(n2507), .A2(n2535), .ZN(n2757) );
  NOR2_X1 U1921 ( .A1(n2758), .A2(n2528), .ZN(n2756) );
  NAND3_X1 U1922 ( .A1(n2759), .A2(n2760), .A3(n2761), .ZN(n2755) );
  NAND2_X1 U1923 ( .A1(n2730), .A2(G143), .ZN(n2761) );
  NAND2_X1 U1924 ( .A1(G150), .A2(n2573), .ZN(n2760) );
  NAND2_X1 U1925 ( .A1(G137), .A2(n2504), .ZN(n2759) );
  NAND4_X1 U1926 ( .A1(n2581), .A2(n2762), .A3(n2763), .A4(n2764), .ZN(n2754) );
  NAND2_X1 U1927 ( .A1(n2572), .A2(n2585), .ZN(n2764) );
  NAND2_X1 U1928 ( .A1(n2519), .A2(G132), .ZN(n2762) );
  NOR4_X1 U1929 ( .A1(n2765), .A2(n2766), .A3(n2767), .A4(n2768), .ZN(n2752) );
  NOR2_X1 U1930 ( .A1(n2507), .A2(n2600), .ZN(n2768) );
  NOR2_X1 U1931 ( .A1(n2758), .A2(n2486), .ZN(n2767) );
  NAND3_X1 U1932 ( .A1(n2769), .A2(n2770), .A3(n2771), .ZN(n2766) );
  NAND2_X1 U1933 ( .A1(G294), .A2(n2730), .ZN(n2771) );
  NAND2_X1 U1934 ( .A1(G283), .A2(n2573), .ZN(n2770) );
  NAND2_X1 U1935 ( .A1(G303), .A2(n2504), .ZN(n2769) );
  NAND4_X1 U1936 ( .A1(n2568), .A2(n2772), .A3(n2773), .A4(n2774), .ZN(n2765) );
  NAND2_X1 U1937 ( .A1(n2572), .A2(n2620), .ZN(n2774) );
  NAND2_X1 U1938 ( .A1(n2567), .A2(n2540), .ZN(n2773) );
  NAND2_X1 U1939 ( .A1(G311), .A2(n2519), .ZN(n2772) );
  NOR2_X1 U1940 ( .A1(n2538), .A2(n2775), .ZN(n2751) );
  NAND2_X1 U1941 ( .A1(n2776), .A2(n2716), .ZN(n2749) );
  NAND2_X1 U1942 ( .A1(n2604), .A2(n2748), .ZN(n2744) );
  NAND3_X1 U1943 ( .A1(n2777), .A2(n2778), .A3(n2779), .ZN(n2748) );
  NAND2_X1 U1944 ( .A1(n2605), .A2(n2780), .ZN(n2779) );
  OR3_X1 U1945 ( .A1(n2781), .A2(n2780), .A3(n2782), .ZN(n2778) );
  NAND2_X1 U1946 ( .A1(n2782), .A2(n2783), .ZN(n2777) );
  NAND2_X1 U1947 ( .A1(n2784), .A2(n2785), .ZN(n2783) );
  NAND2_X1 U1948 ( .A1(n2776), .A2(n2781), .ZN(n2785) );
  NOR2_X1 U1949 ( .A1(n2786), .A2(n2462), .ZN(G381) );
  XNOR2_X1 U1950 ( .A(n2441), .B(keyinput84), .ZN(n2462) );
  INV_X1 U1951 ( .A(n2441), .ZN(n2786) );
  NAND3_X1 U1952 ( .A1(n2787), .A2(n2788), .A3(n2789), .ZN(n2441) );
  XOR2_X1 U1953 ( .A(n2790), .B(keyinput78), .Z(n2789) );
  NAND2_X1 U1954 ( .A1(n2471), .A2(n2791), .ZN(n2790) );
  NAND3_X1 U1955 ( .A1(n2554), .A2(n2792), .A3(n2793), .ZN(n2788) );
  NOR3_X1 U1956 ( .A1(n2794), .A2(n2795), .A3(n2796), .ZN(n2793) );
  NOR4_X1 U1957 ( .A1(n2797), .A2(n2798), .A3(n2799), .A4(n2800), .ZN(n2796) );
  NOR2_X1 U1958 ( .A1(n2530), .A2(n2507), .ZN(n2800) );
  NOR2_X1 U1959 ( .A1(n2758), .A2(n2600), .ZN(n2799) );
  NAND3_X1 U1960 ( .A1(n2801), .A2(n2802), .A3(n2803), .ZN(n2798) );
  NAND2_X1 U1961 ( .A1(G283), .A2(n2730), .ZN(n2803) );
  NAND2_X1 U1962 ( .A1(n2566), .A2(n2573), .ZN(n2802) );
  NAND2_X1 U1963 ( .A1(G294), .A2(n2504), .ZN(n2801) );
  NAND4_X1 U1964 ( .A1(n2568), .A2(n2804), .A3(n2805), .A4(n2584), .ZN(n2797) );
  NAND2_X1 U1965 ( .A1(n2572), .A2(n2540), .ZN(n2584) );
  NAND2_X1 U1966 ( .A1(n2538), .A2(n2567), .ZN(n2805) );
  NAND2_X1 U1967 ( .A1(G303), .A2(n2519), .ZN(n2804) );
  NOR4_X1 U1968 ( .A1(n2806), .A2(n2807), .A3(n2808), .A4(n2809), .ZN(n2795) );
  NOR2_X1 U1969 ( .A1(n2507), .A2(n2528), .ZN(n2809) );
  NOR2_X1 U1970 ( .A1(n2758), .A2(n2643), .ZN(n2808) );
  NAND3_X1 U1971 ( .A1(n2810), .A2(n2811), .A3(n2812), .ZN(n2807) );
  NAND2_X1 U1972 ( .A1(G137), .A2(n2730), .ZN(n2812) );
  NAND2_X1 U1973 ( .A1(G143), .A2(n2573), .ZN(n2811) );
  NAND2_X1 U1974 ( .A1(G132), .A2(n2504), .ZN(n2810) );
  NAND4_X1 U1975 ( .A1(n2581), .A2(n2813), .A3(n2814), .A4(n2815), .ZN(n2806) );
  NAND2_X1 U1976 ( .A1(n2572), .A2(n2589), .ZN(n2815) );
  NAND2_X1 U1977 ( .A1(n2567), .A2(n2585), .ZN(n2814) );
  NAND2_X1 U1978 ( .A1(G128), .A2(n2519), .ZN(n2813) );
  NOR2_X1 U1979 ( .A1(n2586), .A2(n2775), .ZN(n2794) );
  NAND2_X1 U1980 ( .A1(n2716), .A2(n2816), .ZN(n2792) );
  NAND2_X1 U1981 ( .A1(n2817), .A2(n2604), .ZN(n2787) );
  XOR2_X1 U1982 ( .A(n2791), .B(n2818), .Z(n2817) );
  INV_X1 U1983 ( .A(n2447), .ZN(G378) );
  XOR2_X1 U1984 ( .A(n2433), .B(keyinput83), .Z(n2447) );
  NAND3_X1 U1985 ( .A1(n2819), .A2(n2820), .A3(n2821), .ZN(n2433) );
  NAND2_X1 U1986 ( .A1(n2822), .A2(n2471), .ZN(n2821) );
  INV_X1 U1987 ( .A(n2651), .ZN(n2471) );
  NAND3_X1 U1988 ( .A1(n2554), .A2(n2823), .A3(n2824), .ZN(n2820) );
  NOR3_X1 U1989 ( .A1(n2825), .A2(n2826), .A3(n2827), .ZN(n2824) );
  NOR4_X1 U1990 ( .A1(n2828), .A2(n2829), .A3(n2830), .A4(n2831), .ZN(n2827) );
  NOR2_X1 U1991 ( .A1(n2639), .A2(n2507), .ZN(n2831) );
  NOR2_X1 U1992 ( .A1(n2530), .A2(n2758), .ZN(n2830) );
  NAND3_X1 U1993 ( .A1(n2832), .A2(n2833), .A3(n2834), .ZN(n2829) );
  NAND2_X1 U1994 ( .A1(n2566), .A2(n2730), .ZN(n2834) );
  NAND2_X1 U1995 ( .A1(n2835), .A2(n2573), .ZN(n2833) );
  NAND2_X1 U1996 ( .A1(G283), .A2(n2504), .ZN(n2832) );
  NAND4_X1 U1997 ( .A1(n2568), .A2(n2836), .A3(n2763), .A4(n2837), .ZN(n2828) );
  NAND2_X1 U1998 ( .A1(n2538), .A2(n2572), .ZN(n2837) );
  NAND2_X1 U1999 ( .A1(n2567), .A2(n2586), .ZN(n2763) );
  NAND2_X1 U2000 ( .A1(G294), .A2(n2519), .ZN(n2836) );
  INV_X1 U2001 ( .A(n2503), .ZN(n2568) );
  NOR4_X1 U2002 ( .A1(n2838), .A2(n2839), .A3(n2840), .A4(n2841), .ZN(n2826) );
  NOR2_X1 U2003 ( .A1(n2643), .A2(n2507), .ZN(n2841) );
  NOR2_X1 U2004 ( .A1(n2638), .A2(n2758), .ZN(n2840) );
  NAND3_X1 U2005 ( .A1(n2842), .A2(n2843), .A3(n2844), .ZN(n2839) );
  NAND2_X1 U2006 ( .A1(n2730), .A2(G132), .ZN(n2844) );
  NAND2_X1 U2007 ( .A1(G137), .A2(n2573), .ZN(n2843) );
  NAND2_X1 U2008 ( .A1(G128), .A2(n2504), .ZN(n2842) );
  NAND4_X1 U2009 ( .A1(n2581), .A2(n2845), .A3(n2846), .A4(n2847), .ZN(n2838) );
  NAND2_X1 U2010 ( .A1(n2572), .A2(G159), .ZN(n2847) );
  NAND2_X1 U2011 ( .A1(n2567), .A2(n2589), .ZN(n2846) );
  NAND2_X1 U2012 ( .A1(G125), .A2(n2519), .ZN(n2845) );
  INV_X1 U2013 ( .A(n2527), .ZN(n2581) );
  NOR2_X1 U2014 ( .A1(n2775), .A2(n2585), .ZN(n2825) );
  NAND2_X1 U2015 ( .A1(n2848), .A2(n2716), .ZN(n2823) );
  NAND2_X1 U2016 ( .A1(n2849), .A2(n2604), .ZN(n2819) );
  INV_X1 U2017 ( .A(n2542), .ZN(n2604) );
  XNOR2_X1 U2018 ( .A(n2822), .B(n2850), .ZN(n2849) );
  NAND2_X1 U2019 ( .A1(n2818), .A2(n2791), .ZN(n2850) );
  XOR2_X1 U2020 ( .A(n2432), .B(keyinput85), .Z(G375) );
  NAND2_X1 U2021 ( .A1(n2851), .A2(n2852), .ZN(n2432) );
  NAND3_X1 U2022 ( .A1(n2853), .A2(n2854), .A3(n2477), .ZN(n2852) );
  NAND3_X1 U2023 ( .A1(n2651), .A2(n2855), .A3(n2818), .ZN(n2854) );
  NOR2_X1 U2024 ( .A1(n2856), .A2(n2857), .ZN(n2818) );
  NOR2_X1 U2025 ( .A1(n2781), .A2(n2858), .ZN(n2857) );
  NAND2_X1 U2026 ( .A1(n2822), .A2(n2791), .ZN(n2855) );
  NAND3_X1 U2027 ( .A1(n2859), .A2(n2860), .A3(n2861), .ZN(n2791) );
  NAND2_X1 U2028 ( .A1(n2862), .A2(n2863), .ZN(n2861) );
  INV_X1 U2029 ( .A(n2864), .ZN(n2862) );
  OR3_X1 U2030 ( .A1(n2863), .A2(n2865), .A3(n2816), .ZN(n2860) );
  NAND2_X1 U2031 ( .A1(n2866), .A2(n2816), .ZN(n2859) );
  INV_X1 U2032 ( .A(n2867), .ZN(n2816) );
  XOR2_X1 U2033 ( .A(n2863), .B(n2865), .Z(n2866) );
  AND3_X1 U2034 ( .A1(n2868), .A2(n2869), .A3(n2870), .ZN(n2822) );
  NAND2_X1 U2035 ( .A1(n2848), .A2(n2871), .ZN(n2870) );
  XOR2_X1 U2036 ( .A(n2864), .B(n2872), .Z(n2871) );
  NAND3_X1 U2037 ( .A1(n2873), .A2(n2864), .A3(n2872), .ZN(n2869) );
  NAND2_X1 U2038 ( .A1(n2874), .A2(n2875), .ZN(n2868) );
  INV_X1 U2039 ( .A(n2872), .ZN(n2875) );
  XOR2_X1 U2040 ( .A(n2876), .B(n2877), .Z(n2853) );
  XNOR2_X1 U2041 ( .A(n2874), .B(n2878), .ZN(n2877) );
  NAND4_X1 U2042 ( .A1(n2879), .A2(n2880), .A3(n2881), .A4(n2554), .ZN(n2851) );
  INV_X1 U2043 ( .A(n2477), .ZN(n2554) );
  NAND2_X1 U2044 ( .A1(n2542), .A2(n2651), .ZN(n2477) );
  XOR2_X1 U2045 ( .A(n2882), .B(keyinput24), .Z(n2651) );
  NAND2_X1 U2046 ( .A1(n2883), .A2(n2884), .ZN(n2882) );
  NAND3_X1 U2047 ( .A1(n2885), .A2(n2717), .A3(G45), .ZN(n2884) );
  XNOR2_X1 U2048 ( .A(n2886), .B(keyinput26), .ZN(n2542) );
  NAND2_X1 U2049 ( .A1(n2878), .A2(n2716), .ZN(n2881) );
  XNOR2_X1 U2050 ( .A(n2887), .B(n2888), .ZN(n2878) );
  NOR2_X1 U2051 ( .A1(n2889), .A2(n2890), .ZN(n2888) );
  NAND2_X1 U2052 ( .A1(n2535), .A2(n2891), .ZN(n2880) );
  NAND2_X1 U2053 ( .A1(n2775), .A2(n2892), .ZN(n2891) );
  NAND2_X1 U2054 ( .A1(G41), .A2(n2893), .ZN(n2892) );
  OR2_X1 U2055 ( .A1(n2893), .A2(n2716), .ZN(n2775) );
  NOR2_X1 U2056 ( .A1(n2719), .A2(n2885), .ZN(n2716) );
  NAND2_X1 U2057 ( .A1(n2894), .A2(n2895), .ZN(n2879) );
  NAND2_X1 U2058 ( .A1(n2896), .A2(n2897), .ZN(n2894) );
  NAND4_X1 U2059 ( .A1(n2898), .A2(n2899), .A3(n2900), .A4(n2901), .ZN(n2897) );
  NOR4_X1 U2060 ( .A1(n2902), .A2(n2903), .A3(n2904), .A4(n2503), .ZN(n2901) );
  NAND2_X1 U2061 ( .A1(n2893), .A2(n2719), .ZN(n2503) );
  NOR2_X1 U2062 ( .A1(n2537), .A2(n2505), .ZN(n2904) );
  NOR2_X1 U2063 ( .A1(n2639), .A2(n2758), .ZN(n2903) );
  NOR2_X1 U2064 ( .A1(n2530), .A2(n2516), .ZN(n2902) );
  INV_X1 U2065 ( .A(n2573), .ZN(n2516) );
  NOR3_X1 U2066 ( .A1(n2576), .A2(n2905), .A3(n2906), .ZN(n2900) );
  NOR2_X1 U2067 ( .A1(n2529), .A2(n2506), .ZN(n2906) );
  INV_X1 U2068 ( .A(G283), .ZN(n2506) );
  INV_X1 U2069 ( .A(n2519), .ZN(n2529) );
  NOR2_X1 U2070 ( .A1(n2534), .A2(n2486), .ZN(n2905) );
  NOR2_X1 U2071 ( .A1(n2507), .A2(n2591), .ZN(n2576) );
  NAND2_X1 U2072 ( .A1(n2835), .A2(n2730), .ZN(n2899) );
  NAND2_X1 U2073 ( .A1(n2572), .A2(n2586), .ZN(n2898) );
  NAND4_X1 U2074 ( .A1(n2907), .A2(n2908), .A3(n2909), .A4(n2910), .ZN(n2896) );
  NOR4_X1 U2075 ( .A1(n2911), .A2(n2912), .A3(n2913), .A4(n2527), .ZN(n2910) );
  NAND2_X1 U2076 ( .A1(n2893), .A2(n2731), .ZN(n2527) );
  INV_X1 U2077 ( .A(n2715), .ZN(n2893) );
  NAND2_X1 U2078 ( .A1(n2914), .A2(n2915), .ZN(n2715) );
  NAND2_X1 U2079 ( .A1(n2916), .A2(n2917), .ZN(n2915) );
  NOR2_X1 U2080 ( .A1(n2528), .A2(n2505), .ZN(n2913) );
  INV_X1 U2081 ( .A(n2567), .ZN(n2505) );
  NOR2_X1 U2082 ( .A1(n2739), .A2(n2758), .ZN(n2912) );
  INV_X1 U2083 ( .A(n2518), .ZN(n2758) );
  INV_X1 U2084 ( .A(G137), .ZN(n2739) );
  AND2_X1 U2085 ( .A1(n2573), .A2(G132), .ZN(n2911) );
  NOR3_X1 U2086 ( .A1(n2923), .A2(n2924), .A3(n2925), .ZN(n2909) );
  AND2_X1 U2087 ( .A1(G124), .A2(n2519), .ZN(n2925) );
  NOR2_X1 U2088 ( .A1(n2926), .A2(n2920), .ZN(n2519) );
  AND2_X1 U2089 ( .A1(n2504), .A2(G125), .ZN(n2924) );
  INV_X1 U2090 ( .A(n2534), .ZN(n2504) );
  NAND3_X1 U2091 ( .A1(n2922), .A2(n2920), .A3(n2919), .ZN(n2534) );
  NOR2_X1 U2092 ( .A1(n2638), .A2(n2507), .ZN(n2923) );
  NAND4_X1 U2093 ( .A1(n2922), .A2(n2917), .A3(n2921), .A4(n2920), .ZN(n2507) );
  INV_X1 U2094 ( .A(G143), .ZN(n2638) );
  NAND2_X1 U2095 ( .A1(G128), .A2(n2730), .ZN(n2908) );
  INV_X1 U2096 ( .A(n2514), .ZN(n2730) );
  NAND3_X1 U2097 ( .A1(n2918), .A2(n2920), .A3(n2919), .ZN(n2514) );
  INV_X1 U2098 ( .A(n2921), .ZN(n2919) );
  INV_X1 U2099 ( .A(n2927), .ZN(n2920) );
  INV_X1 U2100 ( .A(n2922), .ZN(n2918) );
  NAND2_X1 U2101 ( .A1(n2572), .A2(G150), .ZN(n2907) );
  NOR2_X1 U2102 ( .A1(n2926), .A2(n2927), .ZN(n2572) );
  NOR2_X1 U2103 ( .A1(n2717), .A2(n2928), .ZN(n2927) );
  NAND2_X1 U2104 ( .A1(n2921), .A2(n2929), .ZN(n2926) );
  NAND2_X1 U2105 ( .A1(n2922), .A2(n2917), .ZN(n2929) );
  NAND2_X1 U2106 ( .A1(n2917), .A2(n2930), .ZN(n2921) );
  NOR2_X1 U2107 ( .A1(n2858), .A2(n2931), .ZN(G372) );
  NAND2_X1 U2108 ( .A1(n2932), .A2(n2933), .ZN(G369) );
  NAND2_X1 U2109 ( .A1(n2934), .A2(n2935), .ZN(n2933) );
  NAND3_X1 U2110 ( .A1(n2936), .A2(n2937), .A3(n2938), .ZN(G367) );
  NAND3_X1 U2111 ( .A1(n2939), .A2(n2940), .A3(n2941), .ZN(n2938) );
  NAND2_X1 U2112 ( .A1(n2942), .A2(n2536), .ZN(n2940) );
  NAND3_X1 U2113 ( .A1(n2538), .A2(n2589), .A3(n2585), .ZN(n2942) );
  NAND3_X1 U2114 ( .A1(n2589), .A2(n2943), .A3(n2586), .ZN(n2939) );
  NAND2_X1 U2115 ( .A1(n2537), .A2(n2538), .ZN(n2943) );
  NAND3_X1 U2116 ( .A1(n2944), .A2(n2945), .A3(n2946), .ZN(n2937) );
  INV_X1 U2117 ( .A(n2941), .ZN(n2945) );
  XOR2_X1 U2118 ( .A(n2947), .B(n2948), .Z(n2944) );
  XOR2_X1 U2119 ( .A(n2856), .B(n2876), .Z(n2948) );
  XOR2_X1 U2120 ( .A(n2949), .B(keyinput71), .Z(n2876) );
  NAND2_X1 U2121 ( .A1(n2950), .A2(n2951), .ZN(n2949) );
  NAND2_X1 U2122 ( .A1(n2873), .A2(n2872), .ZN(n2951) );
  NAND2_X1 U2123 ( .A1(n2952), .A2(n2953), .ZN(n2872) );
  NAND2_X1 U2124 ( .A1(n2867), .A2(n2863), .ZN(n2953) );
  NAND2_X1 U2125 ( .A1(n2954), .A2(n2955), .ZN(n2863) );
  NAND2_X1 U2126 ( .A1(n2780), .A2(n2782), .ZN(n2955) );
  NAND2_X1 U2127 ( .A1(n2956), .A2(n2682), .ZN(n2954) );
  NAND2_X1 U2128 ( .A1(n2957), .A2(n2682), .ZN(n2952) );
  NAND2_X1 U2129 ( .A1(n2890), .A2(n2958), .ZN(n2950) );
  NAND2_X1 U2130 ( .A1(n2932), .A2(n2959), .ZN(n2856) );
  NAND2_X1 U2131 ( .A1(n2934), .A2(n2782), .ZN(n2959) );
  AND3_X1 U2132 ( .A1(n2960), .A2(n2961), .A3(n2962), .ZN(n2932) );
  NAND2_X1 U2133 ( .A1(n2887), .A2(n2963), .ZN(n2961) );
  NAND2_X1 U2134 ( .A1(n2964), .A2(n2965), .ZN(n2963) );
  NAND2_X1 U2135 ( .A1(n2966), .A2(n2967), .ZN(n2965) );
  NAND2_X1 U2136 ( .A1(n2968), .A2(n2969), .ZN(n2967) );
  NAND2_X1 U2137 ( .A1(n2970), .A2(n2956), .ZN(n2969) );
  NAND2_X1 U2138 ( .A1(n2971), .A2(n2972), .ZN(n2947) );
  NAND2_X1 U2139 ( .A1(n2874), .A2(n2858), .ZN(n2972) );
  NOR2_X1 U2140 ( .A1(n2864), .A2(n2848), .ZN(n2874) );
  NAND2_X1 U2141 ( .A1(n2867), .A2(n2865), .ZN(n2864) );
  INV_X1 U2142 ( .A(n2784), .ZN(n2865) );
  NAND2_X1 U2143 ( .A1(n2973), .A2(n2780), .ZN(n2784) );
  NAND3_X1 U2144 ( .A1(n2973), .A2(n2974), .A3(n2934), .ZN(n2971) );
  INV_X1 U2145 ( .A(n2858), .ZN(n2934) );
  NAND4_X1 U2146 ( .A1(n2975), .A2(n2966), .A3(n2970), .A4(n2887), .ZN(n2858) );
  XNOR2_X1 U2147 ( .A(n2976), .B(keyinput51), .ZN(n2887) );
  NAND3_X1 U2148 ( .A1(n2960), .A2(n2977), .A3(n2962), .ZN(n2976) );
  XOR2_X1 U2149 ( .A(n2978), .B(keyinput38), .Z(n2962) );
  NAND3_X1 U2150 ( .A1(n2979), .A2(n2980), .A3(n2981), .ZN(n2978) );
  NAND3_X1 U2151 ( .A1(n2982), .A2(n2983), .A3(n2889), .ZN(n2977) );
  INV_X1 U2152 ( .A(n2980), .ZN(n2889) );
  NAND2_X1 U2153 ( .A1(n2922), .A2(n2979), .ZN(n2983) );
  NAND2_X1 U2154 ( .A1(n2928), .A2(n2984), .ZN(n2982) );
  XNOR2_X1 U2155 ( .A(n2985), .B(keyinput39), .ZN(n2960) );
  NAND3_X1 U2156 ( .A1(n2930), .A2(n2980), .A3(n2984), .ZN(n2985) );
  INV_X1 U2157 ( .A(n2979), .ZN(n2984) );
  NAND3_X1 U2158 ( .A1(n2986), .A2(n2987), .A3(n2988), .ZN(n2979) );
  NAND2_X1 U2159 ( .A1(n2989), .A2(G226), .ZN(n2988) );
  NAND2_X1 U2160 ( .A1(n2990), .A2(n2991), .ZN(n2986) );
  NAND3_X1 U2161 ( .A1(n2992), .A2(n2993), .A3(n2994), .ZN(n2991) );
  NAND2_X1 U2162 ( .A1(n2538), .A2(n2719), .ZN(n2994) );
  NAND2_X1 U2163 ( .A1(G223), .A2(n2995), .ZN(n2993) );
  NAND2_X1 U2164 ( .A1(G222), .A2(n2996), .ZN(n2992) );
  NAND4_X1 U2165 ( .A1(n2997), .A2(n2998), .A3(n2999), .A4(n3000), .ZN(n2980) );
  NOR2_X1 U2166 ( .A1(n3001), .A2(n3002), .ZN(n3000) );
  NOR2_X1 U2167 ( .A1(n2643), .A2(n3003), .ZN(n3002) );
  INV_X1 U2168 ( .A(G150), .ZN(n2643) );
  AND2_X1 U2169 ( .A1(n3004), .A2(n2585), .ZN(n3001) );
  NAND2_X1 U2170 ( .A1(n3005), .A2(n2586), .ZN(n2999) );
  NAND2_X1 U2171 ( .A1(n3006), .A2(n2535), .ZN(n2998) );
  NAND2_X1 U2172 ( .A1(n2589), .A2(n3007), .ZN(n2997) );
  NAND3_X1 U2173 ( .A1(n2873), .A2(n2780), .A3(n2867), .ZN(n2974) );
  XOR2_X1 U2174 ( .A(n3008), .B(n3009), .Z(n2867) );
  XNOR2_X1 U2175 ( .A(n3010), .B(n2970), .ZN(n3009) );
  XOR2_X1 U2176 ( .A(n3011), .B(keyinput52), .Z(n2970) );
  NAND2_X1 U2177 ( .A1(n2968), .A2(n3012), .ZN(n3011) );
  NAND3_X1 U2178 ( .A1(n3013), .A2(n3014), .A3(n3015), .ZN(n3012) );
  NAND2_X1 U2179 ( .A1(n2922), .A2(n3016), .ZN(n3014) );
  NAND2_X1 U2180 ( .A1(n2928), .A2(n3017), .ZN(n3013) );
  INV_X1 U2181 ( .A(n2957), .ZN(n2968) );
  NAND2_X1 U2182 ( .A1(n3018), .A2(n3019), .ZN(n2957) );
  XOR2_X1 U2183 ( .A(keyinput40), .B(n3020), .Z(n3019) );
  NOR3_X1 U2184 ( .A1(n2916), .A2(n3015), .A3(n3017), .ZN(n3020) );
  XOR2_X1 U2185 ( .A(n3021), .B(keyinput41), .Z(n3018) );
  NAND3_X1 U2186 ( .A1(n2930), .A2(n3022), .A3(n3017), .ZN(n3021) );
  INV_X1 U2187 ( .A(n3016), .ZN(n3017) );
  NAND3_X1 U2188 ( .A1(n3023), .A2(n2987), .A3(n3024), .ZN(n3016) );
  NAND2_X1 U2189 ( .A1(G238), .A2(n2989), .ZN(n3024) );
  NAND2_X1 U2190 ( .A1(n2990), .A2(n3025), .ZN(n3023) );
  NAND3_X1 U2191 ( .A1(n3026), .A2(n3027), .A3(n3028), .ZN(n3025) );
  NAND2_X1 U2192 ( .A1(n2620), .A2(n2719), .ZN(n3028) );
  NAND2_X1 U2193 ( .A1(G232), .A2(n2995), .ZN(n3027) );
  NAND2_X1 U2194 ( .A1(G226), .A2(n2996), .ZN(n3026) );
  NOR2_X1 U2195 ( .A1(n3015), .A2(n2682), .ZN(n3010) );
  INV_X1 U2196 ( .A(n3022), .ZN(n3015) );
  NAND4_X1 U2197 ( .A1(n3029), .A2(n3030), .A3(n3031), .A4(n3032), .ZN(n3022) );
  NAND2_X1 U2198 ( .A1(n3033), .A2(n2586), .ZN(n3032) );
  NAND2_X1 U2199 ( .A1(n2536), .A2(n3034), .ZN(n3031) );
  NAND2_X1 U2200 ( .A1(n3035), .A2(n2538), .ZN(n3030) );
  NAND2_X1 U2201 ( .A1(n3036), .A2(n2589), .ZN(n3029) );
  XNOR2_X1 U2202 ( .A(keyinput61), .B(keyinput34), .ZN(n3008) );
  INV_X1 U2203 ( .A(n2776), .ZN(n2780) );
  XOR2_X1 U2204 ( .A(n3037), .B(n3038), .Z(n2776) );
  XNOR2_X1 U2205 ( .A(n3039), .B(n2975), .ZN(n3038) );
  XOR2_X1 U2206 ( .A(n3040), .B(keyinput53), .Z(n2975) );
  NAND2_X1 U2207 ( .A1(n3041), .A2(n3042), .ZN(n3040) );
  NAND3_X1 U2208 ( .A1(n3043), .A2(n3044), .A3(n3045), .ZN(n3042) );
  NAND2_X1 U2209 ( .A1(n2922), .A2(n3046), .ZN(n3044) );
  NAND2_X1 U2210 ( .A1(n2928), .A2(n3047), .ZN(n3043) );
  INV_X1 U2211 ( .A(n2956), .ZN(n3041) );
  NAND2_X1 U2212 ( .A1(n3048), .A2(n3049), .ZN(n2956) );
  NAND3_X1 U2213 ( .A1(n3046), .A2(n3050), .A3(n2981), .ZN(n3049) );
  XOR2_X1 U2214 ( .A(n3051), .B(keyinput42), .Z(n3048) );
  NAND3_X1 U2215 ( .A1(n2930), .A2(n3050), .A3(n3047), .ZN(n3051) );
  INV_X1 U2216 ( .A(n3046), .ZN(n3047) );
  NAND3_X1 U2217 ( .A1(n3052), .A2(n2987), .A3(n3053), .ZN(n3046) );
  NAND2_X1 U2218 ( .A1(G244), .A2(n2989), .ZN(n3053) );
  NAND2_X1 U2219 ( .A1(n2990), .A2(n3054), .ZN(n3052) );
  NAND3_X1 U2220 ( .A1(n3055), .A2(n3056), .A3(n3057), .ZN(n3054) );
  NAND2_X1 U2221 ( .A1(n2835), .A2(n2719), .ZN(n3057) );
  NAND2_X1 U2222 ( .A1(G238), .A2(n2995), .ZN(n3056) );
  NAND2_X1 U2223 ( .A1(n2996), .A2(G232), .ZN(n3055) );
  NOR2_X1 U2224 ( .A1(n3045), .A2(n2682), .ZN(n3039) );
  INV_X1 U2225 ( .A(n3050), .ZN(n3045) );
  NAND4_X1 U2226 ( .A1(n3058), .A2(n3059), .A3(n3060), .A4(n3061), .ZN(n3050) );
  NAND2_X1 U2227 ( .A1(n3006), .A2(n2591), .ZN(n3061) );
  NAND2_X1 U2228 ( .A1(n2538), .A2(n3007), .ZN(n3060) );
  NAND2_X1 U2229 ( .A1(n3062), .A2(n3063), .ZN(n3007) );
  NAND2_X1 U2230 ( .A1(n3035), .A2(n2540), .ZN(n3059) );
  NAND2_X1 U2231 ( .A1(n3036), .A2(n2585), .ZN(n3058) );
  XNOR2_X1 U2232 ( .A(keyinput62), .B(keyinput35), .ZN(n3037) );
  INV_X1 U2233 ( .A(n2848), .ZN(n2873) );
  XNOR2_X1 U2234 ( .A(n2966), .B(n3064), .ZN(n2848) );
  NOR2_X1 U2235 ( .A1(n3065), .A2(n2890), .ZN(n3064) );
  AND2_X1 U2236 ( .A1(n2964), .A2(n3066), .ZN(n2966) );
  NAND3_X1 U2237 ( .A1(n3067), .A2(n3068), .A3(n3065), .ZN(n3066) );
  NAND2_X1 U2238 ( .A1(n2922), .A2(n3069), .ZN(n3068) );
  NAND2_X1 U2239 ( .A1(n2928), .A2(n3070), .ZN(n3067) );
  INV_X1 U2240 ( .A(n3069), .ZN(n3070) );
  INV_X1 U2241 ( .A(n2958), .ZN(n2964) );
  NAND2_X1 U2242 ( .A1(n3071), .A2(n3072), .ZN(n2958) );
  NAND3_X1 U2243 ( .A1(n3073), .A2(n3069), .A3(n2981), .ZN(n3072) );
  XOR2_X1 U2244 ( .A(keyinput50), .B(n3074), .Z(n3071) );
  NOR3_X1 U2245 ( .A1(n3069), .A2(n3065), .A3(n3075), .ZN(n3074) );
  INV_X1 U2246 ( .A(n3073), .ZN(n3065) );
  NAND4_X1 U2247 ( .A1(n3076), .A2(n3077), .A3(n3078), .A4(n3079), .ZN(n3073) );
  NOR2_X1 U2248 ( .A1(n3080), .A2(n3081), .ZN(n3079) );
  NOR2_X1 U2249 ( .A1(n2528), .A2(n3003), .ZN(n3081) );
  INV_X1 U2250 ( .A(G159), .ZN(n2528) );
  NOR2_X1 U2251 ( .A1(n2536), .A2(n3082), .ZN(n3080) );
  OR2_X1 U2252 ( .A1(n3062), .A2(n3083), .ZN(n3078) );
  NAND2_X1 U2253 ( .A1(n3006), .A2(n2537), .ZN(n3077) );
  NAND2_X1 U2254 ( .A1(n3033), .A2(n2585), .ZN(n3076) );
  INV_X1 U2255 ( .A(n3063), .ZN(n3033) );
  NAND3_X1 U2256 ( .A1(n3084), .A2(n3085), .A3(n3086), .ZN(n3063) );
  NAND2_X1 U2257 ( .A1(n2917), .A2(n3087), .ZN(n3085) );
  NAND3_X1 U2258 ( .A1(n3088), .A2(n2987), .A3(n3089), .ZN(n3069) );
  NAND2_X1 U2259 ( .A1(n2989), .A2(G232), .ZN(n3089) );
  NOR2_X1 U2260 ( .A1(n3090), .A2(n2990), .ZN(n2989) );
  NAND2_X1 U2261 ( .A1(G274), .A2(n3090), .ZN(n2987) );
  AND2_X1 U2262 ( .A1(n3087), .A2(n3091), .ZN(n3090) );
  NAND2_X1 U2263 ( .A1(n2895), .A2(n2494), .ZN(n3091) );
  INV_X1 U2264 ( .A(G45), .ZN(n2494) );
  NAND2_X1 U2265 ( .A1(n2990), .A2(n3092), .ZN(n3088) );
  NAND3_X1 U2266 ( .A1(n3093), .A2(n3094), .A3(n3095), .ZN(n3092) );
  NAND2_X1 U2267 ( .A1(n2540), .A2(n2719), .ZN(n3095) );
  NAND2_X1 U2268 ( .A1(G226), .A2(n2995), .ZN(n3094) );
  NAND2_X1 U2269 ( .A1(G223), .A2(n2996), .ZN(n3093) );
  OR3_X1 U2270 ( .A1(n3096), .A2(n2486), .A3(n2946), .ZN(n2936) );
  NAND3_X1 U2271 ( .A1(n3097), .A2(n3098), .A3(n3099), .ZN(G364) );
  OR2_X1 U2272 ( .A1(n2493), .A2(n2886), .ZN(n3099) );
  NAND3_X1 U2273 ( .A1(n3100), .A2(n2886), .A3(n2883), .ZN(n3098) );
  XNOR2_X1 U2274 ( .A(n3101), .B(keyinput25), .ZN(n2886) );
  NAND2_X1 U2275 ( .A1(n2718), .A2(n2895), .ZN(n3101) );
  INV_X1 U2276 ( .A(G41), .ZN(n2895) );
  INV_X1 U2277 ( .A(n2590), .ZN(n3100) );
  NAND4_X1 U2278 ( .A1(n2639), .A2(n2530), .A3(n2486), .A4(n2600), .ZN(n2590) );
  OR2_X1 U2279 ( .A1(n2883), .A2(n2605), .ZN(n3097) );
  NOR2_X1 U2280 ( .A1(n2782), .A2(n2973), .ZN(n2605) );
  INV_X1 U2281 ( .A(n2781), .ZN(n2973) );
  NAND3_X1 U2282 ( .A1(n3102), .A2(n3103), .A3(n2685), .ZN(n2781) );
  INV_X1 U2283 ( .A(n2544), .ZN(n2685) );
  XNOR2_X1 U2284 ( .A(keyinput16), .B(G330), .ZN(n2544) );
  NAND2_X1 U2285 ( .A1(n2931), .A2(n2682), .ZN(n3103) );
  NAND4_X1 U2286 ( .A1(n2689), .A2(n2712), .A3(n2703), .A4(n2699), .ZN(n2931) );
  XOR2_X1 U2287 ( .A(n3104), .B(keyinput56), .Z(n2689) );
  NAND2_X1 U2288 ( .A1(n3105), .A2(n3106), .ZN(n3104) );
  XOR2_X1 U2289 ( .A(n3107), .B(keyinput28), .Z(n3105) );
  NAND3_X1 U2290 ( .A1(n3108), .A2(n3109), .A3(n3110), .ZN(n3107) );
  NAND2_X1 U2291 ( .A1(n2922), .A2(n3111), .ZN(n3109) );
  NAND2_X1 U2292 ( .A1(n2928), .A2(n3112), .ZN(n3108) );
  NAND2_X1 U2293 ( .A1(n3113), .A2(n2663), .ZN(n3102) );
  NAND2_X1 U2294 ( .A1(n3114), .A2(n3115), .ZN(n3113) );
  NAND2_X1 U2295 ( .A1(n2930), .A2(n3116), .ZN(n3115) );
  NAND4_X1 U2296 ( .A1(n3117), .A2(n3118), .A3(n3112), .A4(n3119), .ZN(n3116) );
  NAND2_X1 U2297 ( .A1(n3075), .A2(n3120), .ZN(n3114) );
  NAND4_X1 U2298 ( .A1(n3111), .A2(n3121), .A3(n3122), .A4(n3123), .ZN(n3120) );
  XNOR2_X1 U2299 ( .A(n3124), .B(keyinput68), .ZN(n2782) );
  NAND2_X1 U2300 ( .A1(n2935), .A2(n2682), .ZN(n3124) );
  INV_X1 U2301 ( .A(n2663), .ZN(n2682) );
  NOR2_X1 U2302 ( .A1(n2451), .A2(n2890), .ZN(n2663) );
  NAND4_X1 U2303 ( .A1(n2885), .A2(G213), .A3(n2717), .A4(n3087), .ZN(n2890) );
  INV_X1 U2304 ( .A(G343), .ZN(n2451) );
  XNOR2_X1 U2305 ( .A(keyinput66), .B(n3125), .ZN(n2935) );
  NAND2_X1 U2306 ( .A1(n3126), .A2(n3127), .ZN(n3125) );
  NAND2_X1 U2307 ( .A1(n2712), .A2(n3128), .ZN(n3127) );
  NAND2_X1 U2308 ( .A1(n2662), .A2(n3129), .ZN(n3128) );
  NAND2_X1 U2309 ( .A1(n2703), .A2(n3130), .ZN(n3129) );
  NAND2_X1 U2310 ( .A1(n3131), .A2(n3132), .ZN(n3130) );
  NAND2_X1 U2311 ( .A1(n2681), .A2(n2699), .ZN(n3132) );
  XNOR2_X1 U2312 ( .A(n3133), .B(keyinput55), .ZN(n2699) );
  NAND2_X1 U2313 ( .A1(n3134), .A2(n3135), .ZN(n3133) );
  XOR2_X1 U2314 ( .A(n3136), .B(keyinput27), .Z(n3134) );
  NAND3_X1 U2315 ( .A1(n3137), .A2(n3138), .A3(n3139), .ZN(n3136) );
  INV_X1 U2316 ( .A(n2701), .ZN(n3139) );
  NAND2_X1 U2317 ( .A1(n2922), .A2(n3121), .ZN(n3138) );
  NAND2_X1 U2318 ( .A1(n2928), .A2(n3119), .ZN(n3137) );
  XNOR2_X1 U2319 ( .A(n3106), .B(keyinput33), .ZN(n2681) );
  AND2_X1 U2320 ( .A1(n3140), .A2(n3141), .ZN(n3106) );
  XOR2_X1 U2321 ( .A(keyinput47), .B(n3142), .Z(n3141) );
  NOR3_X1 U2322 ( .A1(n2916), .A2(n3110), .A3(n3112), .ZN(n3142) );
  INV_X1 U2323 ( .A(n2690), .ZN(n3110) );
  XOR2_X1 U2324 ( .A(n3143), .B(keyinput48), .Z(n3140) );
  NAND3_X1 U2325 ( .A1(n2930), .A2(n2690), .A3(n3112), .ZN(n3143) );
  INV_X1 U2326 ( .A(n3111), .ZN(n3112) );
  NAND3_X1 U2327 ( .A1(n3144), .A2(n3145), .A3(n3146), .ZN(n3111) );
  NAND2_X1 U2328 ( .A1(n2990), .A2(n3147), .ZN(n3146) );
  NAND3_X1 U2329 ( .A1(n3148), .A2(n3149), .A3(n3150), .ZN(n3147) );
  NAND2_X1 U2330 ( .A1(G303), .A2(n2719), .ZN(n3150) );
  NAND2_X1 U2331 ( .A1(G264), .A2(n2995), .ZN(n3149) );
  NAND2_X1 U2332 ( .A1(G257), .A2(n2996), .ZN(n3148) );
  NAND2_X1 U2333 ( .A1(G270), .A2(n3151), .ZN(n3144) );
  NAND4_X1 U2334 ( .A1(n3152), .A2(n3153), .A3(n3154), .A4(n3155), .ZN(n2690) );
  NAND2_X1 U2335 ( .A1(n3006), .A2(n2486), .ZN(n3155) );
  OR2_X1 U2336 ( .A1(n2486), .A2(n3156), .ZN(n3154) );
  NAND2_X1 U2337 ( .A1(n3035), .A2(G283), .ZN(n3153) );
  NAND2_X1 U2338 ( .A1(n3036), .A2(n2620), .ZN(n3152) );
  XOR2_X1 U2339 ( .A(keyinput32), .B(n3135), .Z(n3131) );
  INV_X1 U2340 ( .A(n2684), .ZN(n3135) );
  NAND2_X1 U2341 ( .A1(n3157), .A2(n3158), .ZN(n2684) );
  XOR2_X1 U2342 ( .A(n3159), .B(keyinput45), .Z(n3158) );
  NAND3_X1 U2343 ( .A1(n3121), .A2(n2701), .A3(n2981), .ZN(n3159) );
  INV_X1 U2344 ( .A(n2916), .ZN(n2981) );
  XOR2_X1 U2345 ( .A(n3160), .B(keyinput46), .Z(n3157) );
  NAND3_X1 U2346 ( .A1(n2930), .A2(n2701), .A3(n3119), .ZN(n3160) );
  INV_X1 U2347 ( .A(n3121), .ZN(n3119) );
  NAND3_X1 U2348 ( .A1(n3161), .A2(n3145), .A3(n3162), .ZN(n3121) );
  NAND2_X1 U2349 ( .A1(n2990), .A2(n3163), .ZN(n3162) );
  NAND3_X1 U2350 ( .A1(n3164), .A2(n3165), .A3(n3166), .ZN(n3163) );
  NAND2_X1 U2351 ( .A1(G294), .A2(n2719), .ZN(n3166) );
  NAND2_X1 U2352 ( .A1(G257), .A2(n2995), .ZN(n3165) );
  NAND2_X1 U2353 ( .A1(G250), .A2(n2996), .ZN(n3164) );
  NAND2_X1 U2354 ( .A1(G264), .A2(n3151), .ZN(n3161) );
  NAND4_X1 U2355 ( .A1(n3167), .A2(n3168), .A3(n3169), .A4(n3170), .ZN(n2701) );
  NAND2_X1 U2356 ( .A1(n2600), .A2(n3034), .ZN(n3170) );
  NAND2_X1 U2357 ( .A1(n3086), .A2(n3062), .ZN(n3034) );
  NAND2_X1 U2358 ( .A1(n3171), .A2(n2835), .ZN(n3169) );
  NAND2_X1 U2359 ( .A1(n3035), .A2(n2566), .ZN(n3168) );
  INV_X1 U2360 ( .A(n3082), .ZN(n3035) );
  NAND2_X1 U2361 ( .A1(n3036), .A2(n2540), .ZN(n3167) );
  XNOR2_X1 U2362 ( .A(n3172), .B(keyinput60), .ZN(n2703) );
  NAND2_X1 U2363 ( .A1(n3173), .A2(n3174), .ZN(n3172) );
  NAND3_X1 U2364 ( .A1(n3175), .A2(n3176), .A3(n3177), .ZN(n3174) );
  NAND2_X1 U2365 ( .A1(n2922), .A2(n3122), .ZN(n3176) );
  NAND2_X1 U2366 ( .A1(n2928), .A2(n3118), .ZN(n3175) );
  XNOR2_X1 U2367 ( .A(n3173), .B(keyinput58), .ZN(n2662) );
  AND2_X1 U2368 ( .A1(n3178), .A2(n3179), .ZN(n3173) );
  XOR2_X1 U2369 ( .A(keyinput30), .B(n3180), .Z(n3179) );
  NOR3_X1 U2370 ( .A1(n2916), .A2(n3177), .A3(n3118), .ZN(n3180) );
  INV_X1 U2371 ( .A(n2704), .ZN(n3177) );
  XOR2_X1 U2372 ( .A(n3181), .B(keyinput31), .Z(n3178) );
  NAND3_X1 U2373 ( .A1(n2930), .A2(n2704), .A3(n3118), .ZN(n3181) );
  INV_X1 U2374 ( .A(n3122), .ZN(n3118) );
  NAND3_X1 U2375 ( .A1(n3182), .A2(n3145), .A3(n3183), .ZN(n3122) );
  NAND2_X1 U2376 ( .A1(n2990), .A2(n3184), .ZN(n3183) );
  NAND3_X1 U2377 ( .A1(n3185), .A2(n3186), .A3(n3187), .ZN(n3184) );
  NAND2_X1 U2378 ( .A1(G283), .A2(n2719), .ZN(n3187) );
  NAND2_X1 U2379 ( .A1(G250), .A2(n2995), .ZN(n3186) );
  NAND2_X1 U2380 ( .A1(G244), .A2(n2996), .ZN(n3185) );
  NAND2_X1 U2381 ( .A1(n3188), .A2(G274), .ZN(n3145) );
  NAND2_X1 U2382 ( .A1(G257), .A2(n3151), .ZN(n3182) );
  NOR2_X1 U2383 ( .A1(n3188), .A2(n2990), .ZN(n3151) );
  NOR2_X1 U2384 ( .A1(n3189), .A2(G41), .ZN(n3188) );
  NAND4_X1 U2385 ( .A1(n3190), .A2(n3191), .A3(n3192), .A4(n3193), .ZN(n2704) );
  NOR2_X1 U2386 ( .A1(n3194), .A2(n3195), .ZN(n3193) );
  NOR2_X1 U2387 ( .A1(n2591), .A2(n3003), .ZN(n3195) );
  INV_X1 U2388 ( .A(n2538), .ZN(n2591) );
  NOR2_X1 U2389 ( .A1(n2600), .A2(n3082), .ZN(n3194) );
  NAND3_X1 U2390 ( .A1(n2719), .A2(n2717), .A3(n3196), .ZN(n3082) );
  NAND2_X1 U2391 ( .A1(n3005), .A2(n3096), .ZN(n3192) );
  NAND2_X1 U2392 ( .A1(n3006), .A2(n2530), .ZN(n3191) );
  INV_X1 U2393 ( .A(n3086), .ZN(n3006) );
  NAND2_X1 U2394 ( .A1(n3171), .A2(n2620), .ZN(n3190) );
  XOR2_X1 U2395 ( .A(n3197), .B(keyinput54), .Z(n2712) );
  NAND2_X1 U2396 ( .A1(n3198), .A2(n3199), .ZN(n3197) );
  NAND3_X1 U2397 ( .A1(n3200), .A2(n3201), .A3(n3202), .ZN(n3199) );
  NAND2_X1 U2398 ( .A1(n2922), .A2(n3123), .ZN(n3201) );
  NAND2_X1 U2399 ( .A1(n2928), .A2(n3117), .ZN(n3200) );
  XNOR2_X1 U2400 ( .A(keyinput14), .B(G190), .ZN(n2928) );
  XNOR2_X1 U2401 ( .A(n3198), .B(n3203), .ZN(n3126) );
  XNOR2_X1 U2402 ( .A(keyinput57), .B(keyinput29), .ZN(n3203) );
  AND2_X1 U2403 ( .A1(n3204), .A2(n3205), .ZN(n3198) );
  XOR2_X1 U2404 ( .A(keyinput43), .B(n3206), .Z(n3205) );
  NOR3_X1 U2405 ( .A1(n2916), .A2(n3202), .A3(n3117), .ZN(n3206) );
  INV_X1 U2406 ( .A(n2713), .ZN(n3202) );
  XNOR2_X1 U2407 ( .A(keyinput12), .B(G169), .ZN(n2916) );
  XOR2_X1 U2408 ( .A(n3207), .B(keyinput44), .Z(n3204) );
  NAND3_X1 U2409 ( .A1(n2930), .A2(n2713), .A3(n3117), .ZN(n3207) );
  INV_X1 U2410 ( .A(n3123), .ZN(n3117) );
  NAND3_X1 U2411 ( .A1(n3208), .A2(n3209), .A3(n3210), .ZN(n3123) );
  NAND2_X1 U2412 ( .A1(n3211), .A2(G274), .ZN(n3210) );
  INV_X1 U2413 ( .A(n3189), .ZN(n3211) );
  NAND3_X1 U2414 ( .A1(G250), .A2(n3189), .A3(n3212), .ZN(n3209) );
  NAND2_X1 U2415 ( .A1(G45), .A2(n3087), .ZN(n3189) );
  NAND2_X1 U2416 ( .A1(n2990), .A2(n3213), .ZN(n3208) );
  NAND3_X1 U2417 ( .A1(n3214), .A2(n3215), .A3(n3216), .ZN(n3213) );
  NAND2_X1 U2418 ( .A1(n2566), .A2(n2719), .ZN(n3216) );
  NAND2_X1 U2419 ( .A1(G244), .A2(n2995), .ZN(n3215) );
  NOR2_X1 U2420 ( .A1(n2719), .A2(n2996), .ZN(n2995) );
  NAND2_X1 U2421 ( .A1(G238), .A2(n2996), .ZN(n3214) );
  NOR2_X1 U2422 ( .A1(G1698), .A2(n2719), .ZN(n2996) );
  INV_X1 U2423 ( .A(n3212), .ZN(n2990) );
  NAND2_X1 U2424 ( .A1(n2914), .A2(n3217), .ZN(n3212) );
  NAND2_X1 U2425 ( .A1(G41), .A2(n2719), .ZN(n3217) );
  NAND4_X1 U2426 ( .A1(n3218), .A2(n3219), .A3(n3220), .A4(n3221), .ZN(n2713) );
  NAND2_X1 U2427 ( .A1(n2620), .A2(n3004), .ZN(n3221) );
  NAND2_X1 U2428 ( .A1(n3062), .A2(n3222), .ZN(n3004) );
  NAND2_X1 U2429 ( .A1(n3196), .A2(n2719), .ZN(n3222) );
  NAND2_X1 U2430 ( .A1(n3036), .A2(n2586), .ZN(n3220) );
  INV_X1 U2431 ( .A(n3003), .ZN(n3036) );
  NAND3_X1 U2432 ( .A1(n2731), .A2(n2717), .A3(n3196), .ZN(n3003) );
  NAND2_X1 U2433 ( .A1(n3005), .A2(n2835), .ZN(n3219) );
  NOR2_X1 U2434 ( .A1(n3223), .A2(n3224), .ZN(n3218) );
  NOR2_X1 U2435 ( .A1(n2540), .A2(n3086), .ZN(n3224) );
  NOR2_X1 U2436 ( .A1(n3156), .A2(n2639), .ZN(n3223) );
  NOR2_X1 U2437 ( .A1(n3171), .A2(n3005), .ZN(n3156) );
  INV_X1 U2438 ( .A(n3062), .ZN(n3005) );
  NAND2_X1 U2439 ( .A1(n3196), .A2(n2917), .ZN(n3062) );
  AND3_X1 U2440 ( .A1(n3084), .A2(n3225), .A3(n3086), .ZN(n3171) );
  XOR2_X1 U2441 ( .A(n3226), .B(keyinput23), .Z(n3086) );
  NAND2_X1 U2442 ( .A1(n3227), .A2(n3087), .ZN(n3226) );
  XOR2_X1 U2443 ( .A(n3228), .B(n3229), .Z(n3227) );
  XNOR2_X1 U2444 ( .A(keyinput18), .B(keyinput17), .ZN(n3229) );
  NAND2_X1 U2445 ( .A1(n2885), .A2(n2917), .ZN(n3228) );
  NAND2_X1 U2446 ( .A1(n2719), .A2(n3087), .ZN(n3225) );
  INV_X1 U2447 ( .A(n2731), .ZN(n2719) );
  INV_X1 U2448 ( .A(n3196), .ZN(n3084) );
  XOR2_X1 U2449 ( .A(n3230), .B(keyinput22), .Z(n3196) );
  NAND2_X1 U2450 ( .A1(n3231), .A2(n3232), .ZN(n3230) );
  XOR2_X1 U2451 ( .A(keyinput21), .B(n3233), .Z(n3232) );
  NOR3_X1 U2452 ( .A1(n2717), .A2(n2731), .A3(n3087), .ZN(n3233) );
  XNOR2_X1 U2453 ( .A(keyinput3), .B(G33), .ZN(n2731) );
  INV_X1 U2454 ( .A(n2917), .ZN(n2717) );
  XOR2_X1 U2455 ( .A(keyinput20), .B(n2914), .Z(n3231) );
  INV_X1 U2456 ( .A(n3075), .ZN(n2930) );
  XNOR2_X1 U2457 ( .A(keyinput13), .B(G179), .ZN(n3075) );
  XOR2_X1 U2458 ( .A(n3087), .B(keyinput19), .Z(n2883) );
  NOR3_X1 U2459 ( .A1(n3234), .A2(n3235), .A3(n3236), .ZN(G361) );
  NOR3_X1 U2460 ( .A1(n3237), .A2(n3238), .A3(n3239), .ZN(n3236) );
  INV_X1 U2461 ( .A(G250), .ZN(n3239) );
  NOR2_X1 U2462 ( .A1(G257), .A2(G264), .ZN(n3238) );
  NOR3_X1 U2463 ( .A1(n2718), .A2(n3240), .A3(n3241), .ZN(n3235) );
  NOR2_X1 U2464 ( .A1(n3242), .A2(n3243), .ZN(n3241) );
  NAND4_X1 U2465 ( .A1(n3244), .A2(n3245), .A3(n3246), .A4(n3247), .ZN(n3243) );
  NAND2_X1 U2466 ( .A1(G264), .A2(n2835), .ZN(n3247) );
  NAND2_X1 U2467 ( .A1(G257), .A2(n2620), .ZN(n3246) );
  INV_X1 U2468 ( .A(n2530), .ZN(n2620) );
  NAND2_X1 U2469 ( .A1(G270), .A2(n2566), .ZN(n3245) );
  NAND2_X1 U2470 ( .A1(G250), .A2(n2540), .ZN(n3244) );
  NAND4_X1 U2471 ( .A1(n3248), .A2(n3249), .A3(n3250), .A4(n3251), .ZN(n3242) );
  NAND2_X1 U2472 ( .A1(G244), .A2(n2538), .ZN(n3251) );
  NAND2_X1 U2473 ( .A1(G232), .A2(n2585), .ZN(n3250) );
  NAND2_X1 U2474 ( .A1(G238), .A2(n2586), .ZN(n3249) );
  NAND2_X1 U2475 ( .A1(G226), .A2(n2589), .ZN(n3248) );
  INV_X1 U2476 ( .A(n2946), .ZN(n3240) );
  INV_X1 U2477 ( .A(n3237), .ZN(n2718) );
  NAND2_X1 U2478 ( .A1(n2941), .A2(n2917), .ZN(n3237) );
  NOR2_X1 U2479 ( .A1(n3087), .A2(n2885), .ZN(n2941) );
  NOR2_X1 U2480 ( .A1(n2493), .A2(n2946), .ZN(n3234) );
  NAND2_X1 U2481 ( .A1(n2914), .A2(n2917), .ZN(n2946) );
  XNOR2_X1 U2482 ( .A(keyinput2), .B(G20), .ZN(n2917) );
  NOR2_X1 U2483 ( .A1(n3252), .A2(n3087), .ZN(n2914) );
  XOR2_X1 U2484 ( .A(keyinput0), .B(G1), .Z(n3087) );
  INV_X1 U2485 ( .A(n2885), .ZN(n3252) );
  XNOR2_X1 U2486 ( .A(keyinput1), .B(G13), .ZN(n2885) );
  NAND2_X1 U2487 ( .A1(n2589), .A2(n3253), .ZN(n2493) );
  NAND2_X1 U2488 ( .A1(n2537), .A2(n2536), .ZN(n3253) );
  XOR2_X1 U2489 ( .A(n2714), .B(n2601), .Z(G358) );
  XNOR2_X1 U2490 ( .A(n3254), .B(n3255), .ZN(n2601) );
  XOR2_X1 U2491 ( .A(G244), .B(G238), .Z(n3255) );
  XNOR2_X1 U2492 ( .A(G226), .B(G232), .ZN(n3254) );
  XOR2_X1 U2493 ( .A(n3256), .B(n3257), .Z(n2714) );
  XOR2_X1 U2494 ( .A(G257), .B(G250), .Z(n3257) );
  XNOR2_X1 U2495 ( .A(G270), .B(G264), .ZN(n3256) );
  NAND2_X1 U2496 ( .A1(n2540), .A2(n3258), .ZN(G355) );
  NAND2_X1 U2497 ( .A1(n2530), .A2(n2600), .ZN(n3258) );
  INV_X1 U2498 ( .A(n2639), .ZN(n2540) );
  NOR4_X1 U2499 ( .A1(n2589), .A2(n2538), .A3(n2586), .A4(n2585), .ZN(G353) );
  INV_X1 U2500 ( .A(n2537), .ZN(n2585) );
  INV_X1 U2501 ( .A(n2536), .ZN(n2586) );
  XOR2_X1 U2502 ( .A(n2619), .B(n2495), .Z(G351) );
  XNOR2_X1 U2503 ( .A(n3259), .B(n3083), .ZN(n2495) );
  XOR2_X1 U2504 ( .A(n2536), .B(n2537), .Z(n3083) );
  XNOR2_X1 U2505 ( .A(keyinput5), .B(G58), .ZN(n2537) );
  XNOR2_X1 U2506 ( .A(keyinput6), .B(G68), .ZN(n2536) );
  XOR2_X1 U2507 ( .A(n2538), .B(n2535), .Z(n3259) );
  INV_X1 U2508 ( .A(n2589), .ZN(n2535) );
  XNOR2_X1 U2509 ( .A(keyinput4), .B(G50), .ZN(n2589) );
  XOR2_X1 U2510 ( .A(n3260), .B(n3096), .Z(n2619) );
  XNOR2_X1 U2511 ( .A(n2530), .B(n2600), .ZN(n3096) );
  INV_X1 U2512 ( .A(n2835), .ZN(n2600) );
  XNOR2_X1 U2513 ( .A(keyinput10), .B(G107), .ZN(n2835) );
  XNOR2_X1 U2514 ( .A(keyinput9), .B(G97), .ZN(n2530) );
  XOR2_X1 U2515 ( .A(n2639), .B(n2486), .Z(n3260) );
  INV_X1 U2516 ( .A(n2566), .ZN(n2486) );
  XNOR2_X1 U2517 ( .A(keyinput11), .B(G116), .ZN(n2566) );
  XNOR2_X1 U2518 ( .A(keyinput8), .B(G87), .ZN(n2639) );
endmodule

