//Key = 1000011111010111001001100101010010001001000110011001000111001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370;

XOR2_X1 U750 ( .A(n1036), .B(n1037), .Z(G9) );
AND2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U752 ( .A1(KEYINPUT40), .A2(n1040), .ZN(n1036) );
NOR2_X1 U753 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1043), .A2(n1044), .A3(G953), .A4(n1045), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U756 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U757 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
NOR2_X1 U761 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U764 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
XOR2_X1 U765 ( .A(n1066), .B(KEYINPUT51), .Z(n1064) );
NOR2_X1 U766 ( .A1(n1067), .A2(n1054), .ZN(n1058) );
NOR2_X1 U767 ( .A1(n1039), .A2(n1068), .ZN(n1067) );
NOR3_X1 U768 ( .A1(n1061), .A2(n1069), .A3(n1054), .ZN(n1048) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
INV_X1 U771 ( .A(n1074), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1051), .B(KEYINPUT1), .Z(n1072) );
NOR2_X1 U773 ( .A1(n1075), .A2(n1057), .ZN(n1070) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
INV_X1 U776 ( .A(n1080), .ZN(n1061) );
NAND2_X1 U777 ( .A1(KEYINPUT27), .A2(n1081), .ZN(n1043) );
NOR3_X1 U778 ( .A1(n1045), .A2(G953), .A3(G952), .ZN(n1041) );
AND4_X1 U779 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1045) );
NOR4_X1 U780 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1085) );
NOR2_X1 U781 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U782 ( .A(KEYINPUT35), .B(G472), .Z(n1090) );
AND2_X1 U783 ( .A1(n1091), .A2(G472), .ZN(n1088) );
XOR2_X1 U784 ( .A(G475), .B(n1092), .Z(n1087) );
NAND3_X1 U785 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1086) );
XOR2_X1 U786 ( .A(n1096), .B(G469), .Z(n1095) );
XOR2_X1 U787 ( .A(KEYINPUT43), .B(n1097), .Z(n1094) );
NOR2_X1 U788 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
AND3_X1 U789 ( .A1(n1100), .A2(n1079), .A3(n1065), .ZN(n1084) );
NAND2_X1 U790 ( .A1(n1101), .A2(n1099), .ZN(n1083) );
XOR2_X1 U791 ( .A(KEYINPUT49), .B(n1098), .Z(n1101) );
OR2_X1 U792 ( .A1(n1102), .A2(n1103), .ZN(n1082) );
NAND2_X1 U793 ( .A1(n1104), .A2(n1105), .ZN(G72) );
NAND2_X1 U794 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
INV_X1 U798 ( .A(n1111), .ZN(n1113) );
NAND2_X1 U799 ( .A1(n1114), .A2(G953), .ZN(n1104) );
XOR2_X1 U800 ( .A(n1115), .B(n1112), .Z(n1114) );
XOR2_X1 U801 ( .A(n1110), .B(KEYINPUT60), .Z(n1112) );
NAND2_X1 U802 ( .A1(n1116), .A2(n1117), .ZN(n1110) );
NAND2_X1 U803 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XOR2_X1 U804 ( .A(n1119), .B(n1120), .Z(n1116) );
XOR2_X1 U805 ( .A(KEYINPUT50), .B(G140), .Z(n1120) );
XOR2_X1 U806 ( .A(n1121), .B(G125), .Z(n1119) );
NAND3_X1 U807 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
NAND2_X1 U808 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U809 ( .A1(KEYINPUT31), .A2(n1127), .ZN(n1123) );
NAND2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U811 ( .A(n1130), .B(KEYINPUT4), .Z(n1128) );
NAND2_X1 U812 ( .A1(n1131), .A2(n1132), .ZN(n1122) );
INV_X1 U813 ( .A(KEYINPUT31), .ZN(n1132) );
NAND2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
OR3_X1 U815 ( .A1(n1125), .A2(n1126), .A3(KEYINPUT4), .ZN(n1134) );
INV_X1 U816 ( .A(n1129), .ZN(n1125) );
XNOR2_X1 U817 ( .A(n1135), .B(n1136), .ZN(n1129) );
XOR2_X1 U818 ( .A(n1137), .B(KEYINPUT23), .Z(n1135) );
INV_X1 U819 ( .A(G131), .ZN(n1137) );
NAND2_X1 U820 ( .A1(KEYINPUT4), .A2(n1126), .ZN(n1133) );
NAND2_X1 U821 ( .A1(G900), .A2(G227), .ZN(n1115) );
XOR2_X1 U822 ( .A(n1138), .B(n1139), .Z(G69) );
XOR2_X1 U823 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U824 ( .A1(n1142), .A2(G953), .ZN(n1141) );
NOR2_X1 U825 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U826 ( .A(n1145), .B(KEYINPUT5), .Z(n1143) );
NOR2_X1 U827 ( .A1(n1146), .A2(n1147), .ZN(n1140) );
XOR2_X1 U828 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U829 ( .A(n1150), .B(n1151), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1152), .B(KEYINPUT0), .Z(n1148) );
NOR2_X1 U831 ( .A1(G898), .A2(n1107), .ZN(n1146) );
NOR2_X1 U832 ( .A1(n1153), .A2(n1107), .ZN(n1138) );
NOR2_X1 U833 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NOR2_X1 U834 ( .A1(n1156), .A2(n1157), .ZN(G66) );
XOR2_X1 U835 ( .A(n1158), .B(n1159), .Z(n1157) );
AND2_X1 U836 ( .A1(G217), .A2(n1160), .ZN(n1159) );
NAND2_X1 U837 ( .A1(n1161), .A2(KEYINPUT7), .ZN(n1158) );
NOR2_X1 U838 ( .A1(n1156), .A2(n1162), .ZN(G63) );
XOR2_X1 U839 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U840 ( .A1(n1165), .A2(KEYINPUT12), .ZN(n1164) );
AND2_X1 U841 ( .A1(G478), .A2(n1160), .ZN(n1165) );
NOR2_X1 U842 ( .A1(n1156), .A2(n1166), .ZN(G60) );
NOR3_X1 U843 ( .A1(n1092), .A2(n1167), .A3(n1168), .ZN(n1166) );
AND4_X1 U844 ( .A1(n1169), .A2(KEYINPUT9), .A3(G475), .A4(n1160), .ZN(n1168) );
NOR2_X1 U845 ( .A1(n1170), .A2(n1169), .ZN(n1167) );
AND3_X1 U846 ( .A1(KEYINPUT9), .A2(n1171), .A3(G475), .ZN(n1170) );
INV_X1 U847 ( .A(n1081), .ZN(n1171) );
XOR2_X1 U848 ( .A(n1172), .B(G104), .Z(G6) );
NAND2_X1 U849 ( .A1(KEYINPUT48), .A2(n1173), .ZN(n1172) );
NOR2_X1 U850 ( .A1(n1156), .A2(n1174), .ZN(G57) );
XOR2_X1 U851 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U852 ( .A(n1177), .B(KEYINPUT26), .Z(n1175) );
NAND2_X1 U853 ( .A1(n1160), .A2(G472), .ZN(n1177) );
NOR2_X1 U854 ( .A1(n1156), .A2(n1178), .ZN(G54) );
XOR2_X1 U855 ( .A(n1179), .B(n1180), .Z(n1178) );
XNOR2_X1 U856 ( .A(n1181), .B(n1182), .ZN(n1180) );
XOR2_X1 U857 ( .A(n1183), .B(n1184), .Z(n1179) );
NOR2_X1 U858 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U859 ( .A(KEYINPUT24), .B(n1187), .Z(n1186) );
NOR2_X1 U860 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
AND2_X1 U861 ( .A1(n1188), .A2(n1189), .ZN(n1185) );
XNOR2_X1 U862 ( .A(n1190), .B(n1191), .ZN(n1189) );
XOR2_X1 U863 ( .A(KEYINPUT2), .B(G140), .Z(n1191) );
NAND2_X1 U864 ( .A1(n1160), .A2(G469), .ZN(n1183) );
NOR2_X1 U865 ( .A1(n1156), .A2(n1192), .ZN(G51) );
XOR2_X1 U866 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U867 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U868 ( .A(n1197), .B(n1198), .Z(n1193) );
NAND2_X1 U869 ( .A1(n1160), .A2(n1098), .ZN(n1197) );
NOR2_X1 U870 ( .A1(n1199), .A2(n1081), .ZN(n1160) );
NOR3_X1 U871 ( .A1(n1144), .A2(n1200), .A3(n1111), .ZN(n1081) );
NAND4_X1 U872 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1111) );
NOR3_X1 U873 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1204) );
INV_X1 U874 ( .A(n1208), .ZN(n1206) );
NAND2_X1 U875 ( .A1(n1068), .A2(n1209), .ZN(n1203) );
NAND2_X1 U876 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NAND2_X1 U877 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U878 ( .A(KEYINPUT39), .B(n1054), .Z(n1212) );
NAND2_X1 U879 ( .A1(n1214), .A2(n1063), .ZN(n1210) );
NAND2_X1 U880 ( .A1(n1215), .A2(n1216), .ZN(n1201) );
NAND2_X1 U881 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
NAND2_X1 U882 ( .A1(n1213), .A2(n1039), .ZN(n1218) );
NAND4_X1 U883 ( .A1(n1173), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1144) );
NOR4_X1 U884 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
NOR4_X1 U885 ( .A1(n1226), .A2(n1057), .A3(n1227), .A4(n1228), .ZN(n1225) );
INV_X1 U886 ( .A(n1229), .ZN(n1057) );
NAND2_X1 U887 ( .A1(n1230), .A2(n1039), .ZN(n1226) );
XOR2_X1 U888 ( .A(n1231), .B(KEYINPUT56), .Z(n1230) );
INV_X1 U889 ( .A(n1232), .ZN(n1224) );
INV_X1 U890 ( .A(n1233), .ZN(n1222) );
NAND4_X1 U891 ( .A1(n1074), .A2(n1068), .A3(n1234), .A4(n1235), .ZN(n1219) );
NOR2_X1 U892 ( .A1(n1227), .A2(n1236), .ZN(n1234) );
XOR2_X1 U893 ( .A(n1228), .B(KEYINPUT61), .Z(n1236) );
NAND2_X1 U894 ( .A1(n1068), .A2(n1038), .ZN(n1173) );
AND2_X1 U895 ( .A1(n1237), .A2(n1229), .ZN(n1038) );
NOR2_X1 U896 ( .A1(n1107), .A2(G952), .ZN(n1156) );
XOR2_X1 U897 ( .A(G146), .B(n1238), .Z(G48) );
NOR4_X1 U898 ( .A1(KEYINPUT45), .A2(n1228), .A3(n1239), .A4(n1240), .ZN(n1238) );
XOR2_X1 U899 ( .A(n1241), .B(n1202), .Z(G45) );
NAND4_X1 U900 ( .A1(n1242), .A2(n1213), .A3(n1063), .A4(n1243), .ZN(n1202) );
INV_X1 U901 ( .A(n1244), .ZN(n1213) );
XOR2_X1 U902 ( .A(G140), .B(n1205), .Z(G42) );
AND3_X1 U903 ( .A1(n1077), .A2(n1215), .A3(n1245), .ZN(n1205) );
XOR2_X1 U904 ( .A(G137), .B(n1246), .Z(G39) );
NOR2_X1 U905 ( .A1(n1054), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U906 ( .A(KEYINPUT18), .B(n1217), .ZN(n1247) );
NAND2_X1 U907 ( .A1(n1080), .A2(n1214), .ZN(n1217) );
NAND2_X1 U908 ( .A1(n1248), .A2(n1249), .ZN(G36) );
NAND2_X1 U909 ( .A1(G134), .A2(n1250), .ZN(n1249) );
XOR2_X1 U910 ( .A(KEYINPUT14), .B(n1251), .Z(n1248) );
NOR2_X1 U911 ( .A1(G134), .A2(n1250), .ZN(n1251) );
NAND4_X1 U912 ( .A1(n1252), .A2(n1039), .A3(n1253), .A4(n1215), .ZN(n1250) );
XOR2_X1 U913 ( .A(KEYINPUT52), .B(n1074), .Z(n1253) );
XOR2_X1 U914 ( .A(G131), .B(n1254), .Z(G33) );
NOR3_X1 U915 ( .A1(n1244), .A2(n1054), .A3(n1239), .ZN(n1254) );
INV_X1 U916 ( .A(n1215), .ZN(n1054) );
NAND2_X1 U917 ( .A1(n1255), .A2(n1256), .ZN(n1215) );
OR2_X1 U918 ( .A1(n1228), .A2(KEYINPUT51), .ZN(n1256) );
NAND3_X1 U919 ( .A1(n1066), .A2(n1065), .A3(KEYINPUT51), .ZN(n1255) );
NAND2_X1 U920 ( .A1(n1074), .A2(n1252), .ZN(n1244) );
XOR2_X1 U921 ( .A(n1257), .B(n1258), .Z(G30) );
NAND2_X1 U922 ( .A1(KEYINPUT6), .A2(n1207), .ZN(n1258) );
AND3_X1 U923 ( .A1(n1039), .A2(n1063), .A3(n1214), .ZN(n1207) );
INV_X1 U924 ( .A(n1240), .ZN(n1214) );
NAND3_X1 U925 ( .A1(n1259), .A2(n1260), .A3(n1252), .ZN(n1240) );
AND2_X1 U926 ( .A1(n1077), .A2(n1261), .ZN(n1252) );
INV_X1 U927 ( .A(n1231), .ZN(n1077) );
NAND2_X1 U928 ( .A1(n1262), .A2(n1263), .ZN(G3) );
NAND2_X1 U929 ( .A1(n1223), .A2(n1264), .ZN(n1263) );
XOR2_X1 U930 ( .A(KEYINPUT25), .B(n1265), .Z(n1262) );
NOR2_X1 U931 ( .A1(n1223), .A2(n1264), .ZN(n1265) );
XOR2_X1 U932 ( .A(KEYINPUT36), .B(G101), .Z(n1264) );
AND3_X1 U933 ( .A1(n1074), .A2(n1237), .A3(n1080), .ZN(n1223) );
XOR2_X1 U934 ( .A(G125), .B(n1266), .Z(G27) );
NOR2_X1 U935 ( .A1(KEYINPUT53), .A2(n1208), .ZN(n1266) );
NAND3_X1 U936 ( .A1(n1235), .A2(n1063), .A3(n1245), .ZN(n1208) );
AND4_X1 U937 ( .A1(n1267), .A2(n1068), .A3(n1260), .A4(n1261), .ZN(n1245) );
NAND2_X1 U938 ( .A1(n1268), .A2(n1047), .ZN(n1261) );
NAND2_X1 U939 ( .A1(n1269), .A2(n1118), .ZN(n1268) );
INV_X1 U940 ( .A(G900), .ZN(n1118) );
INV_X1 U941 ( .A(n1228), .ZN(n1063) );
INV_X1 U942 ( .A(n1051), .ZN(n1235) );
XOR2_X1 U943 ( .A(G122), .B(n1200), .Z(G24) );
INV_X1 U944 ( .A(n1145), .ZN(n1200) );
NAND4_X1 U945 ( .A1(n1242), .A2(n1270), .A3(n1229), .A4(n1243), .ZN(n1145) );
NOR2_X1 U946 ( .A1(n1260), .A2(n1259), .ZN(n1229) );
NAND2_X1 U947 ( .A1(n1271), .A2(n1272), .ZN(G21) );
OR2_X1 U948 ( .A1(n1232), .A2(G119), .ZN(n1272) );
XOR2_X1 U949 ( .A(n1273), .B(KEYINPUT46), .Z(n1271) );
NAND2_X1 U950 ( .A1(G119), .A2(n1232), .ZN(n1273) );
NAND4_X1 U951 ( .A1(n1080), .A2(n1270), .A3(n1259), .A4(n1260), .ZN(n1232) );
XOR2_X1 U952 ( .A(n1274), .B(n1233), .Z(G18) );
NAND3_X1 U953 ( .A1(n1270), .A2(n1039), .A3(n1074), .ZN(n1233) );
NOR2_X1 U954 ( .A1(n1242), .A2(n1093), .ZN(n1039) );
XNOR2_X1 U955 ( .A(G113), .B(n1275), .ZN(G15) );
NAND4_X1 U956 ( .A1(KEYINPUT55), .A2(n1074), .A3(n1270), .A4(n1276), .ZN(n1275) );
XOR2_X1 U957 ( .A(KEYINPUT41), .B(n1068), .Z(n1276) );
INV_X1 U958 ( .A(n1239), .ZN(n1068) );
NAND2_X1 U959 ( .A1(n1242), .A2(n1093), .ZN(n1239) );
NOR3_X1 U960 ( .A1(n1228), .A2(n1227), .A3(n1051), .ZN(n1270) );
NAND2_X1 U961 ( .A1(n1277), .A2(n1079), .ZN(n1051) );
INV_X1 U962 ( .A(n1078), .ZN(n1277) );
NOR2_X1 U963 ( .A1(n1260), .A2(n1267), .ZN(n1074) );
XOR2_X1 U964 ( .A(n1190), .B(n1220), .Z(G12) );
NAND2_X1 U965 ( .A1(n1278), .A2(n1237), .ZN(n1220) );
NOR3_X1 U966 ( .A1(n1228), .A2(n1227), .A3(n1231), .ZN(n1237) );
NAND2_X1 U967 ( .A1(n1078), .A2(n1079), .ZN(n1231) );
NAND2_X1 U968 ( .A1(G221), .A2(n1279), .ZN(n1079) );
XNOR2_X1 U969 ( .A(n1280), .B(n1096), .ZN(n1078) );
NAND2_X1 U970 ( .A1(n1281), .A2(n1199), .ZN(n1096) );
XOR2_X1 U971 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U972 ( .A(n1188), .B(n1182), .ZN(n1283) );
NAND2_X1 U973 ( .A1(G227), .A2(n1107), .ZN(n1188) );
XOR2_X1 U974 ( .A(n1284), .B(n1285), .Z(n1282) );
NOR2_X1 U975 ( .A1(KEYINPUT17), .A2(n1181), .ZN(n1285) );
XNOR2_X1 U976 ( .A(n1286), .B(n1126), .ZN(n1181) );
INV_X1 U977 ( .A(n1130), .ZN(n1126) );
XNOR2_X1 U978 ( .A(n1287), .B(n1288), .ZN(n1130) );
NOR2_X1 U979 ( .A1(KEYINPUT16), .A2(n1289), .ZN(n1288) );
NAND2_X1 U980 ( .A1(n1290), .A2(n1291), .ZN(n1286) );
NAND2_X1 U981 ( .A1(n1292), .A2(n1293), .ZN(n1291) );
XOR2_X1 U982 ( .A(KEYINPUT62), .B(n1294), .Z(n1290) );
NOR2_X1 U983 ( .A1(n1292), .A2(n1293), .ZN(n1294) );
NOR2_X1 U984 ( .A1(n1295), .A2(n1296), .ZN(n1284) );
XOR2_X1 U985 ( .A(n1297), .B(KEYINPUT32), .Z(n1296) );
NAND2_X1 U986 ( .A1(G140), .A2(n1190), .ZN(n1297) );
NOR2_X1 U987 ( .A1(G140), .A2(n1190), .ZN(n1295) );
NAND2_X1 U988 ( .A1(KEYINPUT21), .A2(n1298), .ZN(n1280) );
INV_X1 U989 ( .A(G469), .ZN(n1298) );
AND2_X1 U990 ( .A1(n1299), .A2(n1047), .ZN(n1227) );
NAND3_X1 U991 ( .A1(n1300), .A2(n1107), .A3(G952), .ZN(n1047) );
NAND2_X1 U992 ( .A1(n1269), .A2(n1155), .ZN(n1299) );
INV_X1 U993 ( .A(G898), .ZN(n1155) );
AND3_X1 U994 ( .A1(G902), .A2(n1300), .A3(G953), .ZN(n1269) );
NAND2_X1 U995 ( .A1(G237), .A2(G234), .ZN(n1300) );
NAND2_X1 U996 ( .A1(n1301), .A2(n1065), .ZN(n1228) );
NAND2_X1 U997 ( .A1(G214), .A2(n1302), .ZN(n1065) );
INV_X1 U998 ( .A(n1066), .ZN(n1301) );
XOR2_X1 U999 ( .A(n1303), .B(n1098), .Z(n1066) );
AND2_X1 U1000 ( .A1(G210), .A2(n1302), .ZN(n1098) );
NAND2_X1 U1001 ( .A1(n1304), .A2(n1199), .ZN(n1302) );
INV_X1 U1002 ( .A(G237), .ZN(n1304) );
NAND2_X1 U1003 ( .A1(KEYINPUT57), .A2(n1305), .ZN(n1303) );
INV_X1 U1004 ( .A(n1099), .ZN(n1305) );
NAND2_X1 U1005 ( .A1(n1306), .A2(n1199), .ZN(n1099) );
XNOR2_X1 U1006 ( .A(n1195), .B(n1307), .ZN(n1306) );
XOR2_X1 U1007 ( .A(n1152), .B(n1308), .Z(n1307) );
NOR2_X1 U1008 ( .A1(KEYINPUT54), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1009 ( .A(n1196), .B(n1310), .ZN(n1309) );
XNOR2_X1 U1010 ( .A(n1311), .B(n1312), .ZN(n1196) );
NOR2_X1 U1011 ( .A1(G953), .A2(n1154), .ZN(n1312) );
INV_X1 U1012 ( .A(G224), .ZN(n1154) );
XOR2_X1 U1013 ( .A(n1150), .B(n1313), .Z(n1195) );
NOR2_X1 U1014 ( .A1(KEYINPUT59), .A2(n1151), .ZN(n1313) );
XOR2_X1 U1015 ( .A(G122), .B(n1190), .Z(n1151) );
XNOR2_X1 U1016 ( .A(n1314), .B(n1315), .ZN(n1150) );
NOR2_X1 U1017 ( .A1(KEYINPUT20), .A2(n1316), .ZN(n1315) );
XNOR2_X1 U1018 ( .A(n1292), .B(KEYINPUT38), .ZN(n1316) );
XOR2_X1 U1019 ( .A(n1317), .B(n1318), .Z(n1292) );
NAND2_X1 U1020 ( .A1(KEYINPUT8), .A2(n1274), .ZN(n1314) );
INV_X1 U1021 ( .A(G116), .ZN(n1274) );
INV_X1 U1022 ( .A(n1055), .ZN(n1278) );
NAND3_X1 U1023 ( .A1(n1267), .A2(n1260), .A3(n1080), .ZN(n1055) );
NOR2_X1 U1024 ( .A1(n1243), .A2(n1242), .ZN(n1080) );
XNOR2_X1 U1025 ( .A(n1092), .B(n1319), .ZN(n1242) );
NOR2_X1 U1026 ( .A1(G475), .A2(KEYINPUT3), .ZN(n1319) );
NOR2_X1 U1027 ( .A1(n1169), .A2(G902), .ZN(n1092) );
NAND3_X1 U1028 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1169) );
NAND2_X1 U1029 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
OR3_X1 U1030 ( .A1(n1324), .A2(n1323), .A3(KEYINPUT42), .ZN(n1321) );
XOR2_X1 U1031 ( .A(n1325), .B(n1318), .Z(n1323) );
XOR2_X1 U1032 ( .A(G104), .B(KEYINPUT13), .Z(n1318) );
XNOR2_X1 U1033 ( .A(G113), .B(G122), .ZN(n1325) );
NAND2_X1 U1034 ( .A1(KEYINPUT11), .A2(n1326), .ZN(n1324) );
NAND2_X1 U1035 ( .A1(KEYINPUT42), .A2(n1327), .ZN(n1320) );
INV_X1 U1036 ( .A(n1326), .ZN(n1327) );
XNOR2_X1 U1037 ( .A(n1328), .B(n1329), .ZN(n1326) );
XNOR2_X1 U1038 ( .A(n1330), .B(n1289), .ZN(n1329) );
XNOR2_X1 U1039 ( .A(n1241), .B(G146), .ZN(n1289) );
INV_X1 U1040 ( .A(G143), .ZN(n1241) );
NAND2_X1 U1041 ( .A1(G214), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1042 ( .A(n1332), .B(G131), .Z(n1328) );
NAND2_X1 U1043 ( .A1(n1333), .A2(n1334), .ZN(n1332) );
NAND2_X1 U1044 ( .A1(G140), .A2(n1311), .ZN(n1334) );
XOR2_X1 U1045 ( .A(KEYINPUT29), .B(n1335), .Z(n1333) );
NOR2_X1 U1046 ( .A1(G140), .A2(n1311), .ZN(n1335) );
INV_X1 U1047 ( .A(G125), .ZN(n1311) );
INV_X1 U1048 ( .A(n1093), .ZN(n1243) );
XOR2_X1 U1049 ( .A(n1336), .B(G478), .Z(n1093) );
NAND2_X1 U1050 ( .A1(n1163), .A2(n1199), .ZN(n1336) );
XOR2_X1 U1051 ( .A(n1337), .B(n1338), .Z(n1163) );
XOR2_X1 U1052 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1053 ( .A(G134), .B(G128), .Z(n1340) );
XOR2_X1 U1054 ( .A(KEYINPUT22), .B(G143), .Z(n1339) );
XOR2_X1 U1055 ( .A(n1341), .B(n1342), .Z(n1337) );
XNOR2_X1 U1056 ( .A(G122), .B(n1343), .ZN(n1342) );
NAND2_X1 U1057 ( .A1(KEYINPUT15), .A2(G116), .ZN(n1343) );
XOR2_X1 U1058 ( .A(n1344), .B(n1345), .Z(n1341) );
AND2_X1 U1059 ( .A1(n1346), .A2(G217), .ZN(n1345) );
NAND2_X1 U1060 ( .A1(KEYINPUT63), .A2(n1317), .ZN(n1344) );
XNOR2_X1 U1061 ( .A(n1040), .B(KEYINPUT33), .ZN(n1317) );
INV_X1 U1062 ( .A(G107), .ZN(n1040) );
NAND3_X1 U1063 ( .A1(n1347), .A2(n1348), .A3(n1100), .ZN(n1260) );
NAND2_X1 U1064 ( .A1(n1103), .A2(n1102), .ZN(n1100) );
OR3_X1 U1065 ( .A1(n1102), .A2(n1103), .A3(KEYINPUT58), .ZN(n1348) );
NAND2_X1 U1066 ( .A1(n1349), .A2(G217), .ZN(n1102) );
XOR2_X1 U1067 ( .A(n1279), .B(KEYINPUT19), .Z(n1349) );
NAND2_X1 U1068 ( .A1(G234), .A2(n1199), .ZN(n1279) );
NAND2_X1 U1069 ( .A1(KEYINPUT58), .A2(n1103), .ZN(n1347) );
AND2_X1 U1070 ( .A1(n1161), .A2(n1199), .ZN(n1103) );
XOR2_X1 U1071 ( .A(n1350), .B(n1351), .Z(n1161) );
XOR2_X1 U1072 ( .A(n1352), .B(n1353), .Z(n1351) );
NOR2_X1 U1073 ( .A1(KEYINPUT34), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1074 ( .A(n1355), .B(n1356), .Z(n1354) );
XOR2_X1 U1075 ( .A(G119), .B(G110), .Z(n1356) );
XOR2_X1 U1076 ( .A(KEYINPUT10), .B(G128), .Z(n1355) );
NAND2_X1 U1077 ( .A1(G221), .A2(n1346), .ZN(n1352) );
AND2_X1 U1078 ( .A1(G234), .A2(n1107), .ZN(n1346) );
INV_X1 U1079 ( .A(G953), .ZN(n1107) );
NAND2_X1 U1080 ( .A1(n1357), .A2(n1358), .ZN(n1350) );
NAND2_X1 U1081 ( .A1(n1359), .A2(G140), .ZN(n1358) );
NAND2_X1 U1082 ( .A1(n1360), .A2(n1361), .ZN(n1357) );
INV_X1 U1083 ( .A(G140), .ZN(n1361) );
XNOR2_X1 U1084 ( .A(KEYINPUT30), .B(n1359), .ZN(n1360) );
XNOR2_X1 U1085 ( .A(G125), .B(n1362), .ZN(n1359) );
XOR2_X1 U1086 ( .A(G146), .B(G137), .Z(n1362) );
INV_X1 U1087 ( .A(n1259), .ZN(n1267) );
XNOR2_X1 U1088 ( .A(n1091), .B(G472), .ZN(n1259) );
NAND2_X1 U1089 ( .A1(n1176), .A2(n1199), .ZN(n1091) );
INV_X1 U1090 ( .A(G902), .ZN(n1199) );
XNOR2_X1 U1091 ( .A(n1363), .B(n1364), .ZN(n1176) );
XOR2_X1 U1092 ( .A(n1182), .B(n1198), .Z(n1364) );
XNOR2_X1 U1093 ( .A(n1152), .B(n1310), .ZN(n1198) );
XNOR2_X1 U1094 ( .A(n1365), .B(n1366), .ZN(n1310) );
XOR2_X1 U1095 ( .A(G143), .B(n1367), .Z(n1366) );
NOR2_X1 U1096 ( .A1(KEYINPUT28), .A2(n1287), .ZN(n1367) );
XNOR2_X1 U1097 ( .A(n1257), .B(KEYINPUT47), .ZN(n1287) );
INV_X1 U1098 ( .A(G128), .ZN(n1257) );
NAND2_X1 U1099 ( .A1(KEYINPUT44), .A2(G146), .ZN(n1365) );
XOR2_X1 U1100 ( .A(n1293), .B(n1368), .Z(n1152) );
XOR2_X1 U1101 ( .A(G119), .B(G113), .Z(n1368) );
INV_X1 U1102 ( .A(G101), .ZN(n1293) );
XOR2_X1 U1103 ( .A(G131), .B(n1369), .Z(n1182) );
NOR2_X1 U1104 ( .A1(KEYINPUT37), .A2(n1136), .ZN(n1369) );
XNOR2_X1 U1105 ( .A(G137), .B(G134), .ZN(n1136) );
XOR2_X1 U1106 ( .A(n1370), .B(G116), .Z(n1363) );
NAND2_X1 U1107 ( .A1(G210), .A2(n1331), .ZN(n1370) );
NOR2_X1 U1108 ( .A1(G953), .A2(G237), .ZN(n1331) );
INV_X1 U1109 ( .A(G110), .ZN(n1190) );
endmodule


