//Key = 1101111111001110000001001010011011011111111100000001100101101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317;

XNOR2_X1 U721 ( .A(n996), .B(n997), .ZN(G9) );
NOR2_X1 U722 ( .A1(n998), .A2(n999), .ZN(n997) );
XNOR2_X1 U723 ( .A(n1000), .B(KEYINPUT48), .ZN(n998) );
NOR2_X1 U724 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR4_X1 U725 ( .A1(G953), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1002) );
NOR2_X1 U726 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U727 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR3_X1 U728 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1009) );
NOR2_X1 U729 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR3_X1 U730 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NOR2_X1 U731 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
XOR2_X1 U732 ( .A(KEYINPUT47), .B(n1020), .Z(n1019) );
NOR2_X1 U733 ( .A1(n1021), .A2(n1022), .ZN(n1018) );
NOR3_X1 U734 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1013) );
NOR3_X1 U735 ( .A1(n1016), .A2(n1026), .A3(n1027), .ZN(n1025) );
NOR2_X1 U736 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NOR2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1024) );
NOR3_X1 U738 ( .A1(n1023), .A2(n1032), .A3(n1015), .ZN(n1008) );
INV_X1 U739 ( .A(n1030), .ZN(n1015) );
NOR2_X1 U740 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NOR2_X1 U741 ( .A1(n1012), .A2(n1035), .ZN(n1034) );
INV_X1 U742 ( .A(n1036), .ZN(n1012) );
NOR3_X1 U743 ( .A1(n1010), .A2(n1021), .A3(n1016), .ZN(n1033) );
AND3_X1 U744 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1021) );
XNOR2_X1 U745 ( .A(KEYINPUT1), .B(n1040), .ZN(n1039) );
NOR3_X1 U746 ( .A1(n1003), .A2(G953), .A3(G952), .ZN(n1001) );
AND4_X1 U747 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1003) );
NOR4_X1 U748 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1044) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1046) );
XOR2_X1 U750 ( .A(n1051), .B(KEYINPUT43), .Z(n1049) );
NAND3_X1 U751 ( .A1(n1052), .A2(n1037), .A3(n1031), .ZN(n1045) );
NOR3_X1 U752 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1043) );
XNOR2_X1 U753 ( .A(KEYINPUT20), .B(n1056), .ZN(n1055) );
AND2_X1 U754 ( .A1(n1057), .A2(n1058), .ZN(n1054) );
XNOR2_X1 U755 ( .A(n1059), .B(n1060), .ZN(n1053) );
NAND2_X1 U756 ( .A1(n1061), .A2(n1062), .ZN(n1042) );
XOR2_X1 U757 ( .A(n1063), .B(KEYINPUT30), .Z(n1061) );
NOR2_X1 U758 ( .A1(n1064), .A2(n1065), .ZN(n1041) );
INV_X1 U759 ( .A(n1066), .ZN(n1064) );
XOR2_X1 U760 ( .A(n1067), .B(n1068), .Z(G72) );
NOR2_X1 U761 ( .A1(KEYINPUT25), .A2(n1069), .ZN(n1068) );
XOR2_X1 U762 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U763 ( .A1(n1072), .A2(G953), .ZN(n1071) );
NAND3_X1 U764 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1070) );
XOR2_X1 U765 ( .A(KEYINPUT41), .B(n1076), .Z(n1075) );
NOR2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U767 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
XNOR2_X1 U768 ( .A(n1079), .B(n1080), .ZN(n1078) );
XOR2_X1 U769 ( .A(n1081), .B(n1082), .Z(n1080) );
NAND2_X1 U770 ( .A1(KEYINPUT12), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U771 ( .A(G131), .B(KEYINPUT40), .ZN(n1079) );
XNOR2_X1 U772 ( .A(G140), .B(G125), .ZN(n1077) );
INV_X1 U773 ( .A(n1084), .ZN(n1073) );
NOR2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1067) );
XOR2_X1 U775 ( .A(n1087), .B(KEYINPUT14), .Z(n1085) );
NAND2_X1 U776 ( .A1(G900), .A2(G227), .ZN(n1087) );
XOR2_X1 U777 ( .A(n1088), .B(n1089), .Z(G69) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NAND2_X1 U780 ( .A1(n1094), .A2(n1086), .ZN(n1093) );
XOR2_X1 U781 ( .A(KEYINPUT51), .B(n1095), .Z(n1094) );
NOR2_X1 U782 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND3_X1 U783 ( .A1(KEYINPUT6), .A2(n1098), .A3(G953), .ZN(n1092) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1098) );
NOR2_X1 U785 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XNOR2_X1 U786 ( .A(n1101), .B(KEYINPUT7), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1099) );
XOR2_X1 U788 ( .A(n1104), .B(KEYINPUT59), .Z(n1103) );
NAND2_X1 U789 ( .A1(n1057), .A2(n1105), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U791 ( .A1(n1058), .A2(n1005), .ZN(n1107) );
NOR3_X1 U792 ( .A1(n1108), .A2(n1109), .A3(n1106), .ZN(n1102) );
NOR2_X1 U793 ( .A1(n1101), .A2(n1110), .ZN(G63) );
NOR2_X1 U794 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U795 ( .A(KEYINPUT45), .B(n1113), .Z(n1112) );
NOR2_X1 U796 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
AND2_X1 U797 ( .A1(n1115), .A2(n1114), .ZN(n1111) );
NAND2_X1 U798 ( .A1(n1116), .A2(G478), .ZN(n1115) );
NOR2_X1 U799 ( .A1(n1117), .A2(n1118), .ZN(G60) );
XNOR2_X1 U800 ( .A(n1119), .B(n1120), .ZN(n1118) );
NOR2_X1 U801 ( .A1(n1121), .A2(n1108), .ZN(n1119) );
XNOR2_X1 U802 ( .A(n1101), .B(KEYINPUT3), .ZN(n1117) );
XOR2_X1 U803 ( .A(G104), .B(n1122), .Z(G6) );
NOR2_X1 U804 ( .A1(n999), .A2(n1038), .ZN(n1122) );
NOR2_X1 U805 ( .A1(n1101), .A2(n1123), .ZN(G57) );
XOR2_X1 U806 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U808 ( .A1(n1050), .A2(n1108), .ZN(n1127) );
INV_X1 U809 ( .A(G472), .ZN(n1050) );
NOR2_X1 U810 ( .A1(KEYINPUT62), .A2(n1128), .ZN(n1126) );
XOR2_X1 U811 ( .A(KEYINPUT42), .B(n1129), .Z(n1128) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1124) );
NOR2_X1 U813 ( .A1(n1101), .A2(n1132), .ZN(G54) );
XOR2_X1 U814 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U815 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U816 ( .A1(KEYINPUT44), .A2(n1137), .ZN(n1136) );
INV_X1 U817 ( .A(n1138), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1059), .A2(n1108), .ZN(n1135) );
INV_X1 U819 ( .A(G469), .ZN(n1059) );
NOR2_X1 U820 ( .A1(n1101), .A2(n1139), .ZN(G51) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U822 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U823 ( .A1(KEYINPUT8), .A2(n1144), .ZN(n1142) );
NAND2_X1 U824 ( .A1(n1116), .A2(n1145), .ZN(n1144) );
INV_X1 U825 ( .A(n1108), .ZN(n1116) );
NAND2_X1 U826 ( .A1(G902), .A2(n1005), .ZN(n1108) );
NAND3_X1 U827 ( .A1(n1072), .A2(n1146), .A3(n1147), .ZN(n1005) );
XOR2_X1 U828 ( .A(n1096), .B(KEYINPUT33), .Z(n1147) );
NAND3_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1096) );
OR2_X1 U830 ( .A1(n1151), .A2(n1035), .ZN(n1150) );
NAND2_X1 U831 ( .A1(n1152), .A2(n1153), .ZN(n1148) );
NAND2_X1 U832 ( .A1(n1038), .A2(n1040), .ZN(n1153) );
INV_X1 U833 ( .A(n999), .ZN(n1152) );
NAND3_X1 U834 ( .A1(n1154), .A2(n1155), .A3(n1030), .ZN(n999) );
INV_X1 U835 ( .A(n1097), .ZN(n1146) );
NAND4_X1 U836 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1097) );
NAND3_X1 U837 ( .A1(n1026), .A2(n1000), .A3(n1160), .ZN(n1157) );
NOR2_X1 U838 ( .A1(n1161), .A2(n1162), .ZN(n1156) );
NOR2_X1 U839 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
INV_X1 U840 ( .A(KEYINPUT26), .ZN(n1163) );
NOR2_X1 U841 ( .A1(KEYINPUT26), .A2(n1165), .ZN(n1161) );
NAND4_X1 U842 ( .A1(n1166), .A2(n1167), .A3(n1155), .A4(n1035), .ZN(n1165) );
AND4_X1 U843 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1072) );
AND4_X1 U844 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
NAND2_X1 U845 ( .A1(n1176), .A2(n1177), .ZN(n1170) );
NAND2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U847 ( .A1(n1180), .A2(n1029), .A3(n1036), .ZN(n1179) );
NOR2_X1 U848 ( .A1(n1181), .A2(n1182), .ZN(n1140) );
AND2_X1 U849 ( .A1(KEYINPUT21), .A2(n1183), .ZN(n1182) );
NOR3_X1 U850 ( .A1(KEYINPUT21), .A2(n1184), .A3(n1185), .ZN(n1181) );
AND2_X1 U851 ( .A1(G953), .A2(n1186), .ZN(n1101) );
XOR2_X1 U852 ( .A(KEYINPUT52), .B(G952), .Z(n1186) );
XNOR2_X1 U853 ( .A(G146), .B(n1168), .ZN(G48) );
NAND2_X1 U854 ( .A1(n1187), .A2(n1188), .ZN(n1168) );
XNOR2_X1 U855 ( .A(G143), .B(n1169), .ZN(G45) );
NAND4_X1 U856 ( .A1(n1189), .A2(n1026), .A3(n1190), .A4(n1154), .ZN(n1169) );
NOR2_X1 U857 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U858 ( .A(n1193), .B(n1194), .ZN(G42) );
NOR2_X1 U859 ( .A1(KEYINPUT46), .A2(n1175), .ZN(n1194) );
NAND2_X1 U860 ( .A1(n1176), .A2(n1195), .ZN(n1175) );
XNOR2_X1 U861 ( .A(G137), .B(n1196), .ZN(G39) );
NAND4_X1 U862 ( .A1(n1197), .A2(n1176), .A3(n1180), .A4(n1029), .ZN(n1196) );
XNOR2_X1 U863 ( .A(KEYINPUT63), .B(n1036), .ZN(n1197) );
XOR2_X1 U864 ( .A(G134), .B(n1198), .Z(G36) );
NOR2_X1 U865 ( .A1(KEYINPUT16), .A2(n1174), .ZN(n1198) );
NAND3_X1 U866 ( .A1(n1176), .A2(n1000), .A3(n1026), .ZN(n1174) );
XOR2_X1 U867 ( .A(G131), .B(n1199), .Z(G33) );
NOR3_X1 U868 ( .A1(n1178), .A2(KEYINPUT23), .A3(n1200), .ZN(n1199) );
INV_X1 U869 ( .A(n1176), .ZN(n1200) );
NOR4_X1 U870 ( .A1(n1010), .A2(n1201), .A3(n1192), .A4(n1016), .ZN(n1176) );
INV_X1 U871 ( .A(n1031), .ZN(n1016) );
INV_X1 U872 ( .A(n1202), .ZN(n1192) );
XNOR2_X1 U873 ( .A(G128), .B(n1173), .ZN(G30) );
NAND2_X1 U874 ( .A1(n1187), .A2(n1000), .ZN(n1173) );
INV_X1 U875 ( .A(n1040), .ZN(n1000) );
AND3_X1 U876 ( .A1(n1202), .A2(n1029), .A3(n1203), .ZN(n1187) );
XNOR2_X1 U877 ( .A(n1204), .B(n1205), .ZN(G3) );
NOR2_X1 U878 ( .A1(n1206), .A2(n1035), .ZN(n1205) );
XOR2_X1 U879 ( .A(n1151), .B(KEYINPUT50), .Z(n1206) );
NAND4_X1 U880 ( .A1(n1026), .A2(n1020), .A3(n1036), .A4(n1155), .ZN(n1151) );
INV_X1 U881 ( .A(n1201), .ZN(n1020) );
XNOR2_X1 U882 ( .A(G125), .B(n1172), .ZN(G27) );
NAND3_X1 U883 ( .A1(n1207), .A2(n1202), .A3(n1195), .ZN(n1172) );
NOR3_X1 U884 ( .A1(n1029), .A2(n1028), .A3(n1038), .ZN(n1195) );
NAND2_X1 U885 ( .A1(n1007), .A2(n1208), .ZN(n1202) );
NAND3_X1 U886 ( .A1(n1084), .A2(n1209), .A3(n1210), .ZN(n1208) );
XNOR2_X1 U887 ( .A(G902), .B(KEYINPUT5), .ZN(n1210) );
NOR2_X1 U888 ( .A1(n1086), .A2(G900), .ZN(n1084) );
XNOR2_X1 U889 ( .A(G122), .B(n1158), .ZN(G24) );
NAND4_X1 U890 ( .A1(n1189), .A2(n1160), .A3(n1030), .A4(n1211), .ZN(n1158) );
NOR2_X1 U891 ( .A1(n1029), .A2(n1180), .ZN(n1030) );
XNOR2_X1 U892 ( .A(G119), .B(n1159), .ZN(G21) );
NAND4_X1 U893 ( .A1(n1160), .A2(n1036), .A3(n1180), .A4(n1029), .ZN(n1159) );
INV_X1 U894 ( .A(n1212), .ZN(n1029) );
NAND2_X1 U895 ( .A1(n1213), .A2(n1214), .ZN(G18) );
NAND2_X1 U896 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U897 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
NAND2_X1 U898 ( .A1(KEYINPUT11), .A2(n1219), .ZN(n1218) );
OR2_X1 U899 ( .A1(n1220), .A2(KEYINPUT11), .ZN(n1217) );
NAND2_X1 U900 ( .A1(G116), .A2(n1220), .ZN(n1213) );
NOR2_X1 U901 ( .A1(n1221), .A2(KEYINPUT31), .ZN(n1220) );
INV_X1 U902 ( .A(n1219), .ZN(n1221) );
NAND3_X1 U903 ( .A1(n1026), .A2(n1222), .A3(n1160), .ZN(n1219) );
XNOR2_X1 U904 ( .A(KEYINPUT34), .B(n1040), .ZN(n1222) );
NAND2_X1 U905 ( .A1(n1223), .A2(n1189), .ZN(n1040) );
XNOR2_X1 U906 ( .A(n1224), .B(KEYINPUT9), .ZN(n1189) );
XNOR2_X1 U907 ( .A(n1191), .B(KEYINPUT39), .ZN(n1223) );
XNOR2_X1 U908 ( .A(n1225), .B(n1164), .ZN(G15) );
NAND2_X1 U909 ( .A1(n1166), .A2(n1160), .ZN(n1164) );
AND2_X1 U910 ( .A1(n1207), .A2(n1155), .ZN(n1160) );
NOR2_X1 U911 ( .A1(n1023), .A2(n1035), .ZN(n1207) );
INV_X1 U912 ( .A(n1167), .ZN(n1023) );
NOR2_X1 U913 ( .A1(n1022), .A2(n1226), .ZN(n1167) );
INV_X1 U914 ( .A(n1037), .ZN(n1226) );
INV_X1 U915 ( .A(n1178), .ZN(n1166) );
NAND2_X1 U916 ( .A1(n1026), .A2(n1188), .ZN(n1178) );
NOR2_X1 U917 ( .A1(n1180), .A2(n1212), .ZN(n1026) );
NAND2_X1 U918 ( .A1(KEYINPUT37), .A2(n1227), .ZN(n1225) );
XNOR2_X1 U919 ( .A(G110), .B(n1149), .ZN(G12) );
NAND4_X1 U920 ( .A1(n1203), .A2(n1212), .A3(n1036), .A4(n1155), .ZN(n1149) );
NAND2_X1 U921 ( .A1(n1007), .A2(n1228), .ZN(n1155) );
NAND3_X1 U922 ( .A1(n1090), .A2(n1209), .A3(G902), .ZN(n1228) );
NOR2_X1 U923 ( .A1(n1086), .A2(G898), .ZN(n1090) );
NAND3_X1 U924 ( .A1(n1209), .A2(n1086), .A3(G952), .ZN(n1007) );
NAND2_X1 U925 ( .A1(G237), .A2(G234), .ZN(n1209) );
NAND2_X1 U926 ( .A1(n1229), .A2(n1230), .ZN(n1036) );
OR2_X1 U927 ( .A1(n1038), .A2(KEYINPUT39), .ZN(n1230) );
INV_X1 U928 ( .A(n1188), .ZN(n1038) );
NOR2_X1 U929 ( .A1(n1224), .A2(n1191), .ZN(n1188) );
NAND3_X1 U930 ( .A1(n1191), .A2(n1056), .A3(KEYINPUT39), .ZN(n1229) );
INV_X1 U931 ( .A(n1224), .ZN(n1056) );
XNOR2_X1 U932 ( .A(n1231), .B(G478), .ZN(n1224) );
NAND2_X1 U933 ( .A1(n1232), .A2(n1114), .ZN(n1231) );
XNOR2_X1 U934 ( .A(n1233), .B(n1234), .ZN(n1114) );
XOR2_X1 U935 ( .A(n1235), .B(n1236), .Z(n1234) );
XNOR2_X1 U936 ( .A(n1237), .B(G122), .ZN(n1236) );
XOR2_X1 U937 ( .A(G143), .B(G134), .Z(n1235) );
XOR2_X1 U938 ( .A(n1238), .B(n1239), .Z(n1233) );
XNOR2_X1 U939 ( .A(n1216), .B(G107), .ZN(n1239) );
NAND3_X1 U940 ( .A1(G234), .A2(n1086), .A3(G217), .ZN(n1238) );
XNOR2_X1 U941 ( .A(KEYINPUT13), .B(n1240), .ZN(n1232) );
INV_X1 U942 ( .A(n1211), .ZN(n1191) );
NAND3_X1 U943 ( .A1(n1241), .A2(n1242), .A3(n1066), .ZN(n1211) );
NAND3_X1 U944 ( .A1(n1121), .A2(n1240), .A3(n1120), .ZN(n1066) );
INV_X1 U945 ( .A(G475), .ZN(n1121) );
OR2_X1 U946 ( .A1(G475), .A2(KEYINPUT29), .ZN(n1242) );
NAND2_X1 U947 ( .A1(n1065), .A2(KEYINPUT29), .ZN(n1241) );
AND2_X1 U948 ( .A1(G475), .A2(n1243), .ZN(n1065) );
NAND2_X1 U949 ( .A1(n1120), .A2(n1240), .ZN(n1243) );
XOR2_X1 U950 ( .A(n1244), .B(n1245), .Z(n1120) );
XOR2_X1 U951 ( .A(G104), .B(n1246), .Z(n1245) );
NOR2_X1 U952 ( .A1(KEYINPUT17), .A2(n1247), .ZN(n1246) );
XOR2_X1 U953 ( .A(n1248), .B(n1249), .Z(n1247) );
XNOR2_X1 U954 ( .A(n1250), .B(n1251), .ZN(n1249) );
NOR2_X1 U955 ( .A1(n1252), .A2(KEYINPUT53), .ZN(n1250) );
AND3_X1 U956 ( .A1(G214), .A2(n1086), .A3(n1253), .ZN(n1252) );
XNOR2_X1 U957 ( .A(G131), .B(n1254), .ZN(n1248) );
NAND3_X1 U958 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1254) );
NAND2_X1 U959 ( .A1(KEYINPUT18), .A2(n1185), .ZN(n1257) );
OR3_X1 U960 ( .A1(n1185), .A2(KEYINPUT18), .A3(n1258), .ZN(n1256) );
NAND2_X1 U961 ( .A1(n1258), .A2(n1259), .ZN(n1255) );
NAND2_X1 U962 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U963 ( .A(KEYINPUT18), .ZN(n1261) );
XNOR2_X1 U964 ( .A(KEYINPUT61), .B(n1185), .ZN(n1260) );
XNOR2_X1 U965 ( .A(KEYINPUT28), .B(n1193), .ZN(n1258) );
XNOR2_X1 U966 ( .A(G113), .B(G122), .ZN(n1244) );
NOR2_X1 U967 ( .A1(n1262), .A2(n1047), .ZN(n1212) );
NOR2_X1 U968 ( .A1(n1051), .A2(G472), .ZN(n1047) );
AND2_X1 U969 ( .A1(G472), .A2(n1051), .ZN(n1262) );
NAND2_X1 U970 ( .A1(n1263), .A2(n1240), .ZN(n1051) );
XOR2_X1 U971 ( .A(n1264), .B(n1265), .Z(n1263) );
NOR2_X1 U972 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
AND2_X1 U973 ( .A1(KEYINPUT57), .A2(n1131), .ZN(n1267) );
XOR2_X1 U974 ( .A(n1268), .B(n1204), .Z(n1131) );
NOR3_X1 U975 ( .A1(KEYINPUT57), .A2(n1204), .A3(n1268), .ZN(n1266) );
NAND3_X1 U976 ( .A1(n1253), .A2(n1086), .A3(n1269), .ZN(n1268) );
XOR2_X1 U977 ( .A(KEYINPUT22), .B(G210), .Z(n1269) );
XOR2_X1 U978 ( .A(n1130), .B(n1129), .Z(n1264) );
XOR2_X1 U979 ( .A(n1184), .B(n1270), .Z(n1130) );
AND2_X1 U980 ( .A1(n1154), .A2(n1180), .ZN(n1203) );
INV_X1 U981 ( .A(n1028), .ZN(n1180) );
NOR2_X1 U982 ( .A1(n1271), .A2(n1048), .ZN(n1028) );
NOR2_X1 U983 ( .A1(n1057), .A2(n1058), .ZN(n1048) );
AND2_X1 U984 ( .A1(n1058), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U985 ( .A(KEYINPUT60), .B(n1057), .ZN(n1272) );
NAND2_X1 U986 ( .A1(n1106), .A2(n1240), .ZN(n1057) );
XNOR2_X1 U987 ( .A(n1273), .B(n1274), .ZN(n1106) );
XOR2_X1 U988 ( .A(n1275), .B(n1276), .Z(n1274) );
XNOR2_X1 U989 ( .A(n1185), .B(G119), .ZN(n1276) );
INV_X1 U990 ( .A(G125), .ZN(n1185) );
XOR2_X1 U991 ( .A(KEYINPUT28), .B(G137), .Z(n1275) );
XOR2_X1 U992 ( .A(n1277), .B(n1278), .Z(n1273) );
XOR2_X1 U993 ( .A(n1279), .B(n1280), .Z(n1278) );
NOR2_X1 U994 ( .A1(G128), .A2(KEYINPUT2), .ZN(n1279) );
XOR2_X1 U995 ( .A(n1281), .B(n1282), .Z(n1277) );
AND3_X1 U996 ( .A1(G221), .A2(n1086), .A3(G234), .ZN(n1282) );
NAND2_X1 U997 ( .A1(KEYINPUT0), .A2(n1283), .ZN(n1281) );
INV_X1 U998 ( .A(G146), .ZN(n1283) );
INV_X1 U999 ( .A(n1109), .ZN(n1058) );
NAND2_X1 U1000 ( .A1(G217), .A2(n1284), .ZN(n1109) );
NOR2_X1 U1001 ( .A1(n1201), .A2(n1035), .ZN(n1154) );
NAND2_X1 U1002 ( .A1(n1031), .A2(n1010), .ZN(n1035) );
NAND2_X1 U1003 ( .A1(n1052), .A2(n1285), .ZN(n1010) );
OR2_X1 U1004 ( .A1(n1063), .A2(n1145), .ZN(n1285) );
NAND2_X1 U1005 ( .A1(n1145), .A2(n1063), .ZN(n1052) );
NAND2_X1 U1006 ( .A1(n1286), .A2(n1240), .ZN(n1063) );
XOR2_X1 U1007 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U1008 ( .A(n1143), .B(n1183), .Z(n1288) );
XNOR2_X1 U1009 ( .A(n1184), .B(G125), .ZN(n1183) );
XNOR2_X1 U1010 ( .A(n1289), .B(n1251), .ZN(n1184) );
NAND2_X1 U1011 ( .A1(KEYINPUT35), .A2(n1237), .ZN(n1289) );
XNOR2_X1 U1012 ( .A(n1091), .B(n1290), .ZN(n1143) );
XOR2_X1 U1013 ( .A(KEYINPUT27), .B(n1291), .Z(n1290) );
NOR2_X1 U1014 ( .A1(G953), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1015 ( .A(KEYINPUT38), .B(G224), .Z(n1292) );
XNOR2_X1 U1016 ( .A(n1293), .B(n1294), .ZN(n1091) );
XOR2_X1 U1017 ( .A(G122), .B(G110), .Z(n1294) );
XOR2_X1 U1018 ( .A(n1295), .B(n1129), .Z(n1293) );
XNOR2_X1 U1019 ( .A(n1227), .B(n1296), .ZN(n1129) );
XNOR2_X1 U1020 ( .A(G119), .B(n1216), .ZN(n1296) );
INV_X1 U1021 ( .A(G116), .ZN(n1216) );
INV_X1 U1022 ( .A(G113), .ZN(n1227) );
NAND2_X1 U1023 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
NAND2_X1 U1024 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1025 ( .A(KEYINPUT24), .B(n1301), .Z(n1297) );
NOR2_X1 U1026 ( .A1(n1299), .A2(n1300), .ZN(n1301) );
XNOR2_X1 U1027 ( .A(G104), .B(n996), .ZN(n1300) );
XNOR2_X1 U1028 ( .A(KEYINPUT36), .B(G101), .ZN(n1299) );
XNOR2_X1 U1029 ( .A(KEYINPUT58), .B(KEYINPUT15), .ZN(n1287) );
INV_X1 U1030 ( .A(n1062), .ZN(n1145) );
NAND2_X1 U1031 ( .A1(G210), .A2(n1302), .ZN(n1062) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1302), .ZN(n1031) );
NAND2_X1 U1033 ( .A1(n1253), .A2(n1240), .ZN(n1302) );
INV_X1 U1034 ( .A(G237), .ZN(n1253) );
NAND2_X1 U1035 ( .A1(n1022), .A2(n1037), .ZN(n1201) );
NAND2_X1 U1036 ( .A1(G221), .A2(n1284), .ZN(n1037) );
NAND2_X1 U1037 ( .A1(G234), .A2(n1303), .ZN(n1284) );
XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(n1240), .ZN(n1303) );
NAND2_X1 U1039 ( .A1(n1304), .A2(n1305), .ZN(n1022) );
OR2_X1 U1040 ( .A1(n1306), .A2(n1060), .ZN(n1305) );
XOR2_X1 U1041 ( .A(n1307), .B(KEYINPUT56), .Z(n1304) );
NAND2_X1 U1042 ( .A1(n1060), .A2(n1306), .ZN(n1307) );
XOR2_X1 U1043 ( .A(G469), .B(KEYINPUT4), .Z(n1306) );
AND2_X1 U1044 ( .A1(n1308), .A2(n1240), .ZN(n1060) );
INV_X1 U1045 ( .A(G902), .ZN(n1240) );
XOR2_X1 U1046 ( .A(n1133), .B(n1309), .Z(n1308) );
NOR2_X1 U1047 ( .A1(KEYINPUT49), .A2(n1138), .ZN(n1309) );
XNOR2_X1 U1048 ( .A(n1310), .B(n1311), .ZN(n1138) );
XNOR2_X1 U1049 ( .A(n1204), .B(n1312), .ZN(n1311) );
XOR2_X1 U1050 ( .A(KEYINPUT54), .B(G104), .Z(n1312) );
INV_X1 U1051 ( .A(G101), .ZN(n1204) );
XOR2_X1 U1052 ( .A(n1082), .B(n1313), .Z(n1310) );
XOR2_X1 U1053 ( .A(n1314), .B(n1270), .Z(n1313) );
XOR2_X1 U1054 ( .A(n1083), .B(n1315), .Z(n1270) );
NOR2_X1 U1055 ( .A1(G131), .A2(KEYINPUT19), .ZN(n1315) );
XOR2_X1 U1056 ( .A(G134), .B(G137), .Z(n1083) );
NOR2_X1 U1057 ( .A1(KEYINPUT10), .A2(n996), .ZN(n1314) );
INV_X1 U1058 ( .A(G107), .ZN(n996) );
XNOR2_X1 U1059 ( .A(n1316), .B(n1237), .ZN(n1082) );
INV_X1 U1060 ( .A(G128), .ZN(n1237) );
NAND2_X1 U1061 ( .A1(KEYINPUT32), .A2(n1251), .ZN(n1316) );
XNOR2_X1 U1062 ( .A(G143), .B(G146), .ZN(n1251) );
XOR2_X1 U1063 ( .A(n1317), .B(n1280), .Z(n1133) );
XNOR2_X1 U1064 ( .A(G110), .B(n1193), .ZN(n1280) );
INV_X1 U1065 ( .A(G140), .ZN(n1193) );
NAND2_X1 U1066 ( .A1(G227), .A2(n1086), .ZN(n1317) );
INV_X1 U1067 ( .A(G953), .ZN(n1086) );
endmodule


