//Key = 0010110111011010010100100010100111010010000101111111100011100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369;

XOR2_X1 U749 ( .A(n1033), .B(n1034), .Z(G9) );
NAND2_X1 U750 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U751 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
INV_X1 U752 ( .A(KEYINPUT25), .ZN(n1038) );
NAND3_X1 U753 ( .A1(n1039), .A2(n1040), .A3(KEYINPUT25), .ZN(n1035) );
NAND2_X1 U754 ( .A1(KEYINPUT2), .A2(n1041), .ZN(n1033) );
NOR2_X1 U755 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR3_X1 U756 ( .A1(n1044), .A2(G953), .A3(n1045), .ZN(n1043) );
XOR2_X1 U757 ( .A(KEYINPUT56), .B(n1046), .Z(n1044) );
NOR4_X1 U758 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
XOR2_X1 U759 ( .A(n1051), .B(KEYINPUT47), .Z(n1049) );
NAND3_X1 U760 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
NOR2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1048) );
NOR2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR3_X1 U764 ( .A1(n1061), .A2(n1039), .A3(n1062), .ZN(n1059) );
NOR2_X1 U765 ( .A1(KEYINPUT33), .A2(n1063), .ZN(n1062) );
NOR2_X1 U766 ( .A1(n1064), .A2(n1065), .ZN(n1061) );
NOR2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1057) );
NOR2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
NOR2_X1 U771 ( .A1(n1074), .A2(n1063), .ZN(n1073) );
NOR2_X1 U772 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
XNOR2_X1 U773 ( .A(KEYINPUT46), .B(n1063), .ZN(n1076) );
NOR3_X1 U774 ( .A1(n1063), .A2(n1077), .A3(n1078), .ZN(n1068) );
NOR2_X1 U775 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR3_X1 U776 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1079) );
INV_X1 U777 ( .A(KEYINPUT33), .ZN(n1081) );
NOR3_X1 U778 ( .A1(n1084), .A2(n1085), .A3(n1060), .ZN(n1047) );
INV_X1 U779 ( .A(n1052), .ZN(n1060) );
NOR3_X1 U780 ( .A1(n1078), .A2(n1071), .A3(n1067), .ZN(n1052) );
XNOR2_X1 U781 ( .A(n1053), .B(KEYINPUT27), .ZN(n1085) );
INV_X1 U782 ( .A(n1086), .ZN(n1084) );
NOR3_X1 U783 ( .A1(n1045), .A2(G953), .A3(G952), .ZN(n1042) );
AND4_X1 U784 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1045) );
NOR3_X1 U785 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
XOR2_X1 U786 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U787 ( .A1(G469), .A2(KEYINPUT37), .ZN(n1095) );
NOR2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
NAND3_X1 U789 ( .A1(n1064), .A2(n1098), .A3(n1082), .ZN(n1091) );
NOR3_X1 U790 ( .A1(n1065), .A2(n1099), .A3(n1100), .ZN(n1089) );
NOR2_X1 U791 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XNOR2_X1 U792 ( .A(KEYINPUT51), .B(n1103), .ZN(n1102) );
AND2_X1 U793 ( .A1(n1103), .A2(n1101), .ZN(n1099) );
XNOR2_X1 U794 ( .A(G478), .B(n1104), .ZN(n1088) );
NAND2_X1 U795 ( .A1(KEYINPUT17), .A2(n1105), .ZN(n1104) );
XOR2_X1 U796 ( .A(n1106), .B(n1107), .Z(G72) );
XOR2_X1 U797 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U798 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND2_X1 U799 ( .A1(G900), .A2(G227), .ZN(n1110) );
NAND2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U801 ( .A1(G953), .A2(n1113), .ZN(n1112) );
XOR2_X1 U802 ( .A(n1114), .B(n1115), .Z(n1111) );
XNOR2_X1 U803 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NAND2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U806 ( .A(KEYINPUT40), .B(n1122), .Z(n1120) );
XOR2_X1 U807 ( .A(n1123), .B(n1124), .Z(n1114) );
XNOR2_X1 U808 ( .A(n1125), .B(G140), .ZN(n1124) );
NOR2_X1 U809 ( .A1(KEYINPUT21), .A2(n1126), .ZN(n1123) );
NOR2_X1 U810 ( .A1(n1127), .A2(G953), .ZN(n1106) );
XOR2_X1 U811 ( .A(n1128), .B(n1129), .Z(G69) );
XOR2_X1 U812 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U813 ( .A1(n1132), .A2(G953), .ZN(n1131) );
NOR2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
XOR2_X1 U815 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U816 ( .A1(G898), .A2(n1137), .ZN(n1133) );
XNOR2_X1 U817 ( .A(G953), .B(KEYINPUT18), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1138), .A2(n1139), .ZN(n1128) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NOR2_X1 U820 ( .A1(n1142), .A2(n1143), .ZN(G66) );
XOR2_X1 U821 ( .A(KEYINPUT63), .B(n1144), .Z(n1143) );
XOR2_X1 U822 ( .A(n1145), .B(n1146), .Z(n1142) );
NAND3_X1 U823 ( .A1(n1147), .A2(G217), .A3(KEYINPUT50), .ZN(n1145) );
NOR2_X1 U824 ( .A1(n1144), .A2(n1148), .ZN(G63) );
NOR3_X1 U825 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
NOR3_X1 U826 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
NOR2_X1 U827 ( .A1(n1155), .A2(n1156), .ZN(n1150) );
AND2_X1 U828 ( .A1(n1050), .A2(G478), .ZN(n1155) );
NOR2_X1 U829 ( .A1(n1144), .A2(n1157), .ZN(G60) );
XOR2_X1 U830 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U831 ( .A1(n1103), .A2(n1154), .ZN(n1158) );
XOR2_X1 U832 ( .A(G104), .B(n1160), .Z(G6) );
NOR2_X1 U833 ( .A1(n1144), .A2(n1161), .ZN(G57) );
XNOR2_X1 U834 ( .A(n1162), .B(n1163), .ZN(n1161) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
AND2_X1 U836 ( .A1(G472), .A2(n1147), .ZN(n1164) );
NOR2_X1 U837 ( .A1(n1144), .A2(n1166), .ZN(G54) );
XOR2_X1 U838 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U839 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U840 ( .A(n1171), .B(n1172), .Z(n1167) );
XNOR2_X1 U841 ( .A(n1173), .B(n1174), .ZN(n1172) );
AND2_X1 U842 ( .A1(G469), .A2(n1147), .ZN(n1171) );
INV_X1 U843 ( .A(n1154), .ZN(n1147) );
NOR2_X1 U844 ( .A1(n1144), .A2(n1175), .ZN(G51) );
XOR2_X1 U845 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U846 ( .A1(KEYINPUT54), .A2(n1178), .ZN(n1177) );
XNOR2_X1 U847 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U848 ( .A1(n1154), .A2(n1181), .ZN(n1176) );
XOR2_X1 U849 ( .A(KEYINPUT12), .B(G210), .Z(n1181) );
NAND2_X1 U850 ( .A1(G902), .A2(n1050), .ZN(n1154) );
NAND2_X1 U851 ( .A1(n1127), .A2(n1132), .ZN(n1050) );
AND4_X1 U852 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1132) );
NOR4_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
INV_X1 U854 ( .A(n1190), .ZN(n1188) );
NOR2_X1 U855 ( .A1(n1037), .A2(n1160), .ZN(n1184) );
AND4_X1 U856 ( .A1(n1191), .A2(n1192), .A3(n1080), .A4(n1193), .ZN(n1160) );
NOR2_X1 U857 ( .A1(n1194), .A2(n1075), .ZN(n1193) );
NOR2_X1 U858 ( .A1(n1040), .A2(n1194), .ZN(n1037) );
NAND4_X1 U859 ( .A1(n1080), .A2(n1191), .A3(n1195), .A4(n1192), .ZN(n1040) );
AND4_X1 U860 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1127) );
NOR4_X1 U861 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
INV_X1 U862 ( .A(n1204), .ZN(n1201) );
NOR2_X1 U863 ( .A1(n1205), .A2(n1206), .ZN(n1200) );
NOR3_X1 U864 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1198) );
NOR2_X1 U865 ( .A1(n1210), .A2(n1194), .ZN(n1209) );
NOR4_X1 U866 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
NOR2_X1 U867 ( .A1(KEYINPUT19), .A2(n1215), .ZN(n1214) );
NOR3_X1 U868 ( .A1(n1216), .A2(n1075), .A3(n1217), .ZN(n1213) );
NAND3_X1 U869 ( .A1(n1218), .A2(n1206), .A3(n1219), .ZN(n1216) );
INV_X1 U870 ( .A(KEYINPUT22), .ZN(n1206) );
NOR2_X1 U871 ( .A1(KEYINPUT19), .A2(n1220), .ZN(n1212) );
AND3_X1 U872 ( .A1(n1220), .A2(n1215), .A3(KEYINPUT19), .ZN(n1211) );
XOR2_X1 U873 ( .A(n1219), .B(KEYINPUT20), .Z(n1215) );
NOR4_X1 U874 ( .A1(n1039), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1208) );
AND2_X1 U875 ( .A1(n1221), .A2(n1224), .ZN(n1207) );
INV_X1 U876 ( .A(KEYINPUT44), .ZN(n1221) );
NOR2_X1 U877 ( .A1(n1139), .A2(G952), .ZN(n1144) );
XNOR2_X1 U878 ( .A(G146), .B(n1205), .ZN(G48) );
NAND4_X1 U879 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1080), .ZN(n1205) );
XOR2_X1 U880 ( .A(n1228), .B(n1224), .Z(G45) );
NOR2_X1 U881 ( .A1(n1223), .A2(n1229), .ZN(n1224) );
INV_X1 U882 ( .A(n1225), .ZN(n1229) );
NAND4_X1 U883 ( .A1(n1086), .A2(n1080), .A3(n1230), .A4(n1231), .ZN(n1223) );
XNOR2_X1 U884 ( .A(G143), .B(KEYINPUT5), .ZN(n1228) );
XOR2_X1 U885 ( .A(n1196), .B(n1232), .Z(G42) );
NAND2_X1 U886 ( .A1(KEYINPUT38), .A2(G140), .ZN(n1232) );
NAND3_X1 U887 ( .A1(n1054), .A2(n1227), .A3(n1233), .ZN(n1196) );
XNOR2_X1 U888 ( .A(n1197), .B(n1234), .ZN(G39) );
XOR2_X1 U889 ( .A(KEYINPUT15), .B(G137), .Z(n1234) );
NAND3_X1 U890 ( .A1(n1226), .A2(n1235), .A3(n1233), .ZN(n1197) );
XOR2_X1 U891 ( .A(G134), .B(n1203), .Z(G36) );
AND3_X1 U892 ( .A1(n1086), .A2(n1195), .A3(n1233), .ZN(n1203) );
XOR2_X1 U893 ( .A(G131), .B(n1202), .Z(G33) );
AND3_X1 U894 ( .A1(n1227), .A2(n1086), .A3(n1233), .ZN(n1202) );
NOR3_X1 U895 ( .A1(n1218), .A2(n1222), .A3(n1063), .ZN(n1233) );
INV_X1 U896 ( .A(n1053), .ZN(n1063) );
NOR2_X1 U897 ( .A1(n1065), .A2(n1236), .ZN(n1053) );
INV_X1 U898 ( .A(n1237), .ZN(n1236) );
XOR2_X1 U899 ( .A(n1238), .B(n1239), .Z(G30) );
NOR2_X1 U900 ( .A1(KEYINPUT41), .A2(G128), .ZN(n1239) );
NAND2_X1 U901 ( .A1(n1220), .A2(n1225), .ZN(n1238) );
NOR3_X1 U902 ( .A1(n1218), .A2(n1074), .A3(n1217), .ZN(n1220) );
XNOR2_X1 U903 ( .A(G101), .B(n1182), .ZN(G3) );
NAND2_X1 U904 ( .A1(n1240), .A2(n1086), .ZN(n1182) );
XNOR2_X1 U905 ( .A(G125), .B(n1204), .ZN(G27) );
NAND4_X1 U906 ( .A1(n1054), .A2(n1225), .A3(n1227), .A4(n1241), .ZN(n1204) );
NOR2_X1 U907 ( .A1(n1194), .A2(n1222), .ZN(n1225) );
INV_X1 U908 ( .A(n1219), .ZN(n1222) );
NAND2_X1 U909 ( .A1(n1067), .A2(n1242), .ZN(n1219) );
NAND4_X1 U910 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1113), .ZN(n1242) );
INV_X1 U911 ( .A(G900), .ZN(n1113) );
XNOR2_X1 U912 ( .A(G122), .B(n1183), .ZN(G24) );
NAND4_X1 U913 ( .A1(n1244), .A2(n1191), .A3(n1230), .A4(n1231), .ZN(n1183) );
INV_X1 U914 ( .A(n1056), .ZN(n1191) );
NAND2_X1 U915 ( .A1(n1245), .A2(n1087), .ZN(n1056) );
INV_X1 U916 ( .A(n1246), .ZN(n1245) );
NAND2_X1 U917 ( .A1(n1247), .A2(n1248), .ZN(G21) );
NAND2_X1 U918 ( .A1(n1189), .A2(n1249), .ZN(n1248) );
INV_X1 U919 ( .A(n1250), .ZN(n1189) );
XOR2_X1 U920 ( .A(n1251), .B(KEYINPUT59), .Z(n1247) );
NAND2_X1 U921 ( .A1(G119), .A2(n1250), .ZN(n1251) );
NAND3_X1 U922 ( .A1(n1226), .A2(n1235), .A3(n1244), .ZN(n1250) );
INV_X1 U923 ( .A(n1217), .ZN(n1226) );
NAND2_X1 U924 ( .A1(n1252), .A2(n1246), .ZN(n1217) );
XNOR2_X1 U925 ( .A(KEYINPUT39), .B(n1087), .ZN(n1252) );
XNOR2_X1 U926 ( .A(G116), .B(n1190), .ZN(G18) );
NAND3_X1 U927 ( .A1(n1086), .A2(n1195), .A3(n1244), .ZN(n1190) );
INV_X1 U928 ( .A(n1074), .ZN(n1195) );
NAND2_X1 U929 ( .A1(n1230), .A2(n1253), .ZN(n1074) );
XOR2_X1 U930 ( .A(n1254), .B(KEYINPUT49), .Z(n1230) );
NAND2_X1 U931 ( .A1(n1255), .A2(n1256), .ZN(G15) );
NAND2_X1 U932 ( .A1(n1187), .A2(n1257), .ZN(n1256) );
XOR2_X1 U933 ( .A(KEYINPUT43), .B(n1258), .Z(n1255) );
NOR2_X1 U934 ( .A1(n1187), .A2(n1257), .ZN(n1258) );
AND3_X1 U935 ( .A1(n1227), .A2(n1086), .A3(n1244), .ZN(n1187) );
AND3_X1 U936 ( .A1(n1039), .A2(n1192), .A3(n1241), .ZN(n1244) );
INV_X1 U937 ( .A(n1071), .ZN(n1241) );
NAND2_X1 U938 ( .A1(n1259), .A2(n1082), .ZN(n1071) );
INV_X1 U939 ( .A(n1083), .ZN(n1259) );
NOR2_X1 U940 ( .A1(n1246), .A2(n1087), .ZN(n1086) );
INV_X1 U941 ( .A(n1075), .ZN(n1227) );
NAND2_X1 U942 ( .A1(n1231), .A2(n1254), .ZN(n1075) );
INV_X1 U943 ( .A(n1253), .ZN(n1231) );
XNOR2_X1 U944 ( .A(G110), .B(n1260), .ZN(G12) );
NOR2_X1 U945 ( .A1(n1186), .A2(KEYINPUT42), .ZN(n1260) );
AND2_X1 U946 ( .A1(n1240), .A2(n1054), .ZN(n1186) );
AND2_X1 U947 ( .A1(n1087), .A2(n1246), .ZN(n1054) );
NAND3_X1 U948 ( .A1(n1261), .A2(n1262), .A3(n1098), .ZN(n1246) );
NAND2_X1 U949 ( .A1(n1096), .A2(n1097), .ZN(n1098) );
NAND2_X1 U950 ( .A1(n1097), .A2(n1263), .ZN(n1262) );
OR3_X1 U951 ( .A1(n1097), .A2(n1096), .A3(n1263), .ZN(n1261) );
INV_X1 U952 ( .A(KEYINPUT4), .ZN(n1263) );
AND2_X1 U953 ( .A1(n1146), .A2(n1264), .ZN(n1096) );
XNOR2_X1 U954 ( .A(n1265), .B(n1266), .ZN(n1146) );
XOR2_X1 U955 ( .A(G137), .B(n1267), .Z(n1266) );
NOR2_X1 U956 ( .A1(KEYINPUT6), .A2(n1268), .ZN(n1267) );
XOR2_X1 U957 ( .A(n1269), .B(n1270), .Z(n1268) );
NAND3_X1 U958 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(n1269) );
NAND2_X1 U959 ( .A1(n1274), .A2(G140), .ZN(n1273) );
XNOR2_X1 U960 ( .A(n1275), .B(G125), .ZN(n1274) );
NAND3_X1 U961 ( .A1(n1126), .A2(n1173), .A3(n1275), .ZN(n1272) );
NAND2_X1 U962 ( .A1(n1276), .A2(n1277), .ZN(n1271) );
INV_X1 U963 ( .A(n1275), .ZN(n1277) );
XNOR2_X1 U964 ( .A(n1278), .B(G110), .ZN(n1275) );
NAND2_X1 U965 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND2_X1 U966 ( .A1(G128), .A2(n1249), .ZN(n1280) );
XOR2_X1 U967 ( .A(KEYINPUT52), .B(n1281), .Z(n1279) );
NOR2_X1 U968 ( .A1(G128), .A2(n1249), .ZN(n1281) );
NAND3_X1 U969 ( .A1(n1282), .A2(G221), .A3(KEYINPUT28), .ZN(n1265) );
NAND2_X1 U970 ( .A1(n1283), .A2(n1284), .ZN(n1097) );
XNOR2_X1 U971 ( .A(G217), .B(KEYINPUT45), .ZN(n1283) );
XOR2_X1 U972 ( .A(n1285), .B(G472), .Z(n1087) );
NAND2_X1 U973 ( .A1(n1286), .A2(n1264), .ZN(n1285) );
XOR2_X1 U974 ( .A(n1287), .B(n1165), .Z(n1286) );
XNOR2_X1 U975 ( .A(n1288), .B(n1289), .ZN(n1165) );
XOR2_X1 U976 ( .A(n1290), .B(n1291), .Z(n1289) );
NAND2_X1 U977 ( .A1(KEYINPUT58), .A2(n1292), .ZN(n1290) );
XOR2_X1 U978 ( .A(n1293), .B(n1294), .Z(n1288) );
NOR2_X1 U979 ( .A1(KEYINPUT30), .A2(n1295), .ZN(n1287) );
XNOR2_X1 U980 ( .A(KEYINPUT9), .B(n1296), .ZN(n1295) );
INV_X1 U981 ( .A(n1162), .ZN(n1296) );
XNOR2_X1 U982 ( .A(n1297), .B(G101), .ZN(n1162) );
NAND2_X1 U983 ( .A1(G210), .A2(n1298), .ZN(n1297) );
AND4_X1 U984 ( .A1(n1235), .A2(n1039), .A3(n1080), .A4(n1192), .ZN(n1240) );
NAND2_X1 U985 ( .A1(n1067), .A2(n1299), .ZN(n1192) );
NAND4_X1 U986 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1141), .ZN(n1299) );
INV_X1 U987 ( .A(G898), .ZN(n1141) );
NAND3_X1 U988 ( .A1(n1243), .A2(n1139), .A3(n1300), .ZN(n1067) );
XOR2_X1 U989 ( .A(KEYINPUT10), .B(G952), .Z(n1300) );
NAND2_X1 U990 ( .A1(G237), .A2(n1301), .ZN(n1243) );
INV_X1 U991 ( .A(n1218), .ZN(n1080) );
NAND2_X1 U992 ( .A1(n1083), .A2(n1082), .ZN(n1218) );
NAND2_X1 U993 ( .A1(G221), .A2(n1284), .ZN(n1082) );
NAND2_X1 U994 ( .A1(n1301), .A2(n1264), .ZN(n1284) );
XOR2_X1 U995 ( .A(G234), .B(KEYINPUT34), .Z(n1301) );
XNOR2_X1 U996 ( .A(n1094), .B(G469), .ZN(n1083) );
NAND3_X1 U997 ( .A1(n1302), .A2(n1303), .A3(n1264), .ZN(n1094) );
OR3_X1 U998 ( .A1(n1304), .A2(n1305), .A3(KEYINPUT48), .ZN(n1303) );
NAND2_X1 U999 ( .A1(n1306), .A2(KEYINPUT48), .ZN(n1302) );
XNOR2_X1 U1000 ( .A(n1307), .B(n1305), .ZN(n1306) );
XNOR2_X1 U1001 ( .A(n1308), .B(n1169), .ZN(n1305) );
XNOR2_X1 U1002 ( .A(n1293), .B(n1117), .ZN(n1169) );
XNOR2_X1 U1003 ( .A(n1309), .B(n1310), .ZN(n1117) );
XOR2_X1 U1004 ( .A(KEYINPUT53), .B(G128), .Z(n1310) );
NAND2_X1 U1005 ( .A1(KEYINPUT26), .A2(n1311), .ZN(n1309) );
XNOR2_X1 U1006 ( .A(n1312), .B(n1125), .ZN(n1293) );
NAND2_X1 U1007 ( .A1(n1118), .A2(n1313), .ZN(n1312) );
NAND2_X1 U1008 ( .A1(n1314), .A2(n1121), .ZN(n1313) );
XOR2_X1 U1009 ( .A(KEYINPUT29), .B(n1122), .Z(n1314) );
OR2_X1 U1010 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
XOR2_X1 U1011 ( .A(G131), .B(G137), .Z(n1122) );
NAND2_X1 U1012 ( .A1(KEYINPUT14), .A2(n1304), .ZN(n1307) );
XOR2_X1 U1013 ( .A(n1315), .B(n1316), .Z(n1304) );
XOR2_X1 U1014 ( .A(G110), .B(n1174), .Z(n1316) );
AND2_X1 U1015 ( .A1(G227), .A2(n1139), .ZN(n1174) );
NAND2_X1 U1016 ( .A1(KEYINPUT11), .A2(n1173), .ZN(n1315) );
INV_X1 U1017 ( .A(n1194), .ZN(n1039) );
NAND2_X1 U1018 ( .A1(n1237), .A2(n1065), .ZN(n1194) );
NAND2_X1 U1019 ( .A1(n1317), .A2(n1318), .ZN(n1065) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1319), .ZN(n1318) );
NAND2_X1 U1021 ( .A1(n1264), .A2(n1320), .ZN(n1319) );
NAND2_X1 U1022 ( .A1(G237), .A2(n1321), .ZN(n1320) );
NAND3_X1 U1023 ( .A1(n1322), .A2(n1264), .A3(n1323), .ZN(n1317) );
INV_X1 U1024 ( .A(n1321), .ZN(n1323) );
NAND2_X1 U1025 ( .A1(n1324), .A2(n1325), .ZN(n1321) );
NAND2_X1 U1026 ( .A1(n1179), .A2(n1326), .ZN(n1325) );
NAND2_X1 U1027 ( .A1(n1327), .A2(n1180), .ZN(n1324) );
INV_X1 U1028 ( .A(n1326), .ZN(n1180) );
XOR2_X1 U1029 ( .A(n1291), .B(n1125), .Z(n1326) );
INV_X1 U1030 ( .A(G146), .ZN(n1125) );
XNOR2_X1 U1031 ( .A(n1328), .B(n1311), .ZN(n1291) );
NAND2_X1 U1032 ( .A1(KEYINPUT32), .A2(G128), .ZN(n1328) );
XNOR2_X1 U1033 ( .A(n1179), .B(KEYINPUT24), .ZN(n1327) );
XNOR2_X1 U1034 ( .A(n1329), .B(n1330), .ZN(n1179) );
XOR2_X1 U1035 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1036 ( .A(KEYINPUT3), .B(n1126), .ZN(n1332) );
NOR2_X1 U1037 ( .A1(G953), .A2(n1140), .ZN(n1331) );
INV_X1 U1038 ( .A(G224), .ZN(n1140) );
XOR2_X1 U1039 ( .A(n1135), .B(n1333), .Z(n1329) );
NOR2_X1 U1040 ( .A1(KEYINPUT60), .A2(n1136), .ZN(n1333) );
XNOR2_X1 U1041 ( .A(n1294), .B(n1292), .ZN(n1136) );
XNOR2_X1 U1042 ( .A(G113), .B(KEYINPUT8), .ZN(n1292) );
XNOR2_X1 U1043 ( .A(G116), .B(n1249), .ZN(n1294) );
INV_X1 U1044 ( .A(G119), .ZN(n1249) );
XNOR2_X1 U1045 ( .A(n1170), .B(n1334), .ZN(n1135) );
XOR2_X1 U1046 ( .A(KEYINPUT1), .B(G122), .Z(n1334) );
XNOR2_X1 U1047 ( .A(n1308), .B(G110), .ZN(n1170) );
XNOR2_X1 U1048 ( .A(G101), .B(n1335), .ZN(n1308) );
XNOR2_X1 U1049 ( .A(n1041), .B(G104), .ZN(n1335) );
INV_X1 U1050 ( .A(G107), .ZN(n1041) );
INV_X1 U1051 ( .A(G902), .ZN(n1264) );
NAND2_X1 U1052 ( .A1(G237), .A2(G210), .ZN(n1322) );
XOR2_X1 U1053 ( .A(n1064), .B(KEYINPUT23), .Z(n1237) );
NAND2_X1 U1054 ( .A1(G214), .A2(n1336), .ZN(n1064) );
OR2_X1 U1055 ( .A1(G237), .A2(G902), .ZN(n1336) );
INV_X1 U1056 ( .A(n1078), .ZN(n1235) );
NAND2_X1 U1057 ( .A1(n1253), .A2(n1254), .ZN(n1078) );
NAND3_X1 U1058 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1254) );
NAND2_X1 U1059 ( .A1(n1340), .A2(n1153), .ZN(n1339) );
OR3_X1 U1060 ( .A1(n1153), .A2(n1340), .A3(KEYINPUT16), .ZN(n1338) );
NAND2_X1 U1061 ( .A1(KEYINPUT7), .A2(n1149), .ZN(n1340) );
INV_X1 U1062 ( .A(G478), .ZN(n1153) );
NAND2_X1 U1063 ( .A1(KEYINPUT16), .A2(n1105), .ZN(n1337) );
INV_X1 U1064 ( .A(n1149), .ZN(n1105) );
NOR2_X1 U1065 ( .A1(n1156), .A2(G902), .ZN(n1149) );
INV_X1 U1066 ( .A(n1152), .ZN(n1156) );
XNOR2_X1 U1067 ( .A(n1341), .B(n1342), .ZN(n1152) );
XOR2_X1 U1068 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1069 ( .A(G128), .B(G122), .Z(n1344) );
XNOR2_X1 U1070 ( .A(KEYINPUT62), .B(n1311), .ZN(n1343) );
XOR2_X1 U1071 ( .A(n1345), .B(n1346), .Z(n1341) );
XNOR2_X1 U1072 ( .A(n1347), .B(G107), .ZN(n1346) );
INV_X1 U1073 ( .A(G116), .ZN(n1347) );
XOR2_X1 U1074 ( .A(n1348), .B(n1121), .Z(n1345) );
XOR2_X1 U1075 ( .A(G134), .B(KEYINPUT0), .Z(n1121) );
NAND2_X1 U1076 ( .A1(n1282), .A2(G217), .ZN(n1348) );
AND2_X1 U1077 ( .A1(G234), .A2(n1139), .ZN(n1282) );
INV_X1 U1078 ( .A(G953), .ZN(n1139) );
XOR2_X1 U1079 ( .A(n1101), .B(n1103), .Z(n1253) );
INV_X1 U1080 ( .A(G475), .ZN(n1103) );
NOR2_X1 U1081 ( .A1(n1159), .A2(G902), .ZN(n1101) );
XNOR2_X1 U1082 ( .A(n1349), .B(n1350), .ZN(n1159) );
XNOR2_X1 U1083 ( .A(G122), .B(n1257), .ZN(n1350) );
INV_X1 U1084 ( .A(G113), .ZN(n1257) );
XOR2_X1 U1085 ( .A(n1351), .B(G104), .Z(n1349) );
NAND2_X1 U1086 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND4_X1 U1087 ( .A1(n1354), .A2(n1355), .A3(n1356), .A4(n1357), .ZN(n1353) );
NAND2_X1 U1088 ( .A1(n1358), .A2(n1359), .ZN(n1357) );
NAND2_X1 U1089 ( .A1(n1360), .A2(n1361), .ZN(n1356) );
NAND3_X1 U1090 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1352) );
NAND2_X1 U1091 ( .A1(n1354), .A2(n1355), .ZN(n1364) );
INV_X1 U1092 ( .A(KEYINPUT61), .ZN(n1355) );
XNOR2_X1 U1093 ( .A(KEYINPUT35), .B(n1311), .ZN(n1354) );
INV_X1 U1094 ( .A(G143), .ZN(n1311) );
NAND2_X1 U1095 ( .A1(n1360), .A2(n1358), .ZN(n1363) );
XOR2_X1 U1096 ( .A(n1365), .B(KEYINPUT13), .Z(n1358) );
NAND2_X1 U1097 ( .A1(n1361), .A2(n1359), .ZN(n1362) );
INV_X1 U1098 ( .A(n1360), .ZN(n1359) );
XNOR2_X1 U1099 ( .A(n1366), .B(G131), .ZN(n1360) );
NAND2_X1 U1100 ( .A1(G214), .A2(n1298), .ZN(n1366) );
NOR2_X1 U1101 ( .A1(G953), .A2(G237), .ZN(n1298) );
XOR2_X1 U1102 ( .A(n1365), .B(KEYINPUT57), .Z(n1361) );
XOR2_X1 U1103 ( .A(n1270), .B(n1367), .Z(n1365) );
NOR3_X1 U1104 ( .A1(n1368), .A2(KEYINPUT36), .A3(n1276), .ZN(n1367) );
NOR2_X1 U1105 ( .A1(n1126), .A2(G140), .ZN(n1276) );
INV_X1 U1106 ( .A(G125), .ZN(n1126) );
XOR2_X1 U1107 ( .A(KEYINPUT55), .B(n1369), .Z(n1368) );
NOR2_X1 U1108 ( .A1(G125), .A2(n1173), .ZN(n1369) );
INV_X1 U1109 ( .A(G140), .ZN(n1173) );
XNOR2_X1 U1110 ( .A(G146), .B(KEYINPUT31), .ZN(n1270) );
endmodule


