//Key = 0001110110111101011101100000000001010011101111100101100011111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330;

XNOR2_X1 U727 ( .A(G107), .B(n1005), .ZN(G9) );
NOR2_X1 U728 ( .A1(n1006), .A2(n1007), .ZN(G75) );
AND4_X1 U729 ( .A1(n1008), .A2(n1009), .A3(KEYINPUT13), .A4(n1010), .ZN(n1007) );
NOR4_X1 U730 ( .A1(G953), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1010) );
NOR2_X1 U731 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR2_X1 U732 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NOR3_X1 U733 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1017) );
NOR2_X1 U734 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U735 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U736 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NOR2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
AND2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U740 ( .A1(n1033), .A2(n1034), .ZN(n1025) );
NOR2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR3_X1 U743 ( .A1(n1034), .A2(n1039), .A3(n1028), .ZN(n1021) );
NOR2_X1 U744 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR4_X1 U745 ( .A1(n1042), .A2(n1028), .A3(n1034), .A4(n1024), .ZN(n1016) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U747 ( .A1(n1018), .A2(n1045), .ZN(n1043) );
INV_X1 U748 ( .A(n1046), .ZN(n1011) );
NOR3_X1 U749 ( .A1(n1012), .A2(G953), .A3(G952), .ZN(n1006) );
AND4_X1 U750 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1012) );
NOR3_X1 U751 ( .A1(n1032), .A2(n1051), .A3(n1019), .ZN(n1050) );
XOR2_X1 U752 ( .A(n1052), .B(KEYINPUT56), .Z(n1049) );
NAND4_X1 U753 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1037), .ZN(n1052) );
NAND2_X1 U754 ( .A1(n1056), .A2(n1057), .ZN(n1048) );
XOR2_X1 U755 ( .A(n1058), .B(n1059), .Z(n1047) );
XNOR2_X1 U756 ( .A(KEYINPUT57), .B(n1060), .ZN(n1059) );
NAND2_X1 U757 ( .A1(KEYINPUT22), .A2(n1061), .ZN(n1058) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(G72) );
NAND2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XOR2_X1 U760 ( .A(KEYINPUT52), .B(n1066), .Z(n1062) );
NOR2_X1 U761 ( .A1(n1067), .A2(n1065), .ZN(n1066) );
NAND2_X1 U762 ( .A1(G953), .A2(n1068), .ZN(n1065) );
NAND2_X1 U763 ( .A1(G900), .A2(G227), .ZN(n1068) );
XNOR2_X1 U764 ( .A(n1064), .B(KEYINPUT42), .ZN(n1067) );
XNOR2_X1 U765 ( .A(n1069), .B(n1070), .ZN(n1064) );
NOR2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
XOR2_X1 U767 ( .A(n1073), .B(n1074), .Z(n1072) );
XNOR2_X1 U768 ( .A(n1075), .B(n1076), .ZN(n1074) );
XOR2_X1 U769 ( .A(n1077), .B(n1078), .Z(n1073) );
XNOR2_X1 U770 ( .A(n1079), .B(G125), .ZN(n1078) );
NOR2_X1 U771 ( .A1(G900), .A2(n1080), .ZN(n1071) );
XNOR2_X1 U772 ( .A(G953), .B(KEYINPUT26), .ZN(n1080) );
NAND2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1069) );
NAND2_X1 U774 ( .A1(n1009), .A2(n1083), .ZN(n1081) );
XNOR2_X1 U775 ( .A(KEYINPUT40), .B(n1046), .ZN(n1083) );
XOR2_X1 U776 ( .A(n1084), .B(n1085), .Z(G69) );
NAND2_X1 U777 ( .A1(G953), .A2(n1086), .ZN(n1085) );
NAND2_X1 U778 ( .A1(G898), .A2(G224), .ZN(n1086) );
NAND2_X1 U779 ( .A1(KEYINPUT60), .A2(n1087), .ZN(n1084) );
XOR2_X1 U780 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U781 ( .A1(n1082), .A2(n1090), .ZN(n1089) );
NAND2_X1 U782 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
NAND2_X1 U783 ( .A1(n1093), .A2(G953), .ZN(n1092) );
XNOR2_X1 U784 ( .A(n1094), .B(n1095), .ZN(n1091) );
XNOR2_X1 U785 ( .A(n1096), .B(n1097), .ZN(n1095) );
NOR2_X1 U786 ( .A1(KEYINPUT53), .A2(n1098), .ZN(n1097) );
NOR2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(G66) );
XNOR2_X1 U788 ( .A(n1101), .B(n1102), .ZN(n1100) );
XNOR2_X1 U789 ( .A(KEYINPUT14), .B(n1103), .ZN(n1102) );
NOR3_X1 U790 ( .A1(n1104), .A2(KEYINPUT9), .A3(n1105), .ZN(n1103) );
NOR2_X1 U791 ( .A1(n1099), .A2(n1106), .ZN(G63) );
XNOR2_X1 U792 ( .A(n1107), .B(n1108), .ZN(n1106) );
NOR2_X1 U793 ( .A1(n1109), .A2(n1104), .ZN(n1108) );
NOR2_X1 U794 ( .A1(n1099), .A2(n1110), .ZN(G60) );
XNOR2_X1 U795 ( .A(n1111), .B(n1112), .ZN(n1110) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1104), .ZN(n1112) );
XOR2_X1 U797 ( .A(G104), .B(n1114), .Z(G6) );
NOR2_X1 U798 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1099), .A2(n1117), .ZN(G57) );
XOR2_X1 U800 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U801 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U802 ( .A1(n1122), .A2(n1104), .ZN(n1120) );
XOR2_X1 U803 ( .A(n1123), .B(KEYINPUT28), .Z(n1118) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U805 ( .A(KEYINPUT8), .B(n1126), .ZN(n1124) );
NOR2_X1 U806 ( .A1(n1099), .A2(n1127), .ZN(G54) );
NOR2_X1 U807 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1129) );
NOR2_X1 U809 ( .A1(n1060), .A2(n1104), .ZN(n1131) );
NOR2_X1 U810 ( .A1(KEYINPUT48), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U811 ( .A(n1133), .B(n1076), .ZN(n1132) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(n1128) );
INV_X1 U813 ( .A(KEYINPUT48), .ZN(n1135) );
XNOR2_X1 U814 ( .A(n1133), .B(n1136), .ZN(n1134) );
NOR2_X1 U815 ( .A1(n1099), .A2(n1137), .ZN(G51) );
XOR2_X1 U816 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U817 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U818 ( .A1(G125), .A2(KEYINPUT50), .ZN(n1140) );
XOR2_X1 U819 ( .A(n1142), .B(n1143), .Z(n1138) );
XNOR2_X1 U820 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1146), .A2(n1104), .ZN(n1142) );
NAND2_X1 U822 ( .A1(G902), .A2(n1147), .ZN(n1104) );
NAND3_X1 U823 ( .A1(n1009), .A2(n1046), .A3(n1008), .ZN(n1147) );
INV_X1 U824 ( .A(n1090), .ZN(n1008) );
NAND4_X1 U825 ( .A1(n1148), .A2(n1005), .A3(n1149), .A4(n1150), .ZN(n1090) );
NOR4_X1 U826 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
NAND2_X1 U827 ( .A1(n1040), .A2(n1155), .ZN(n1149) );
NAND2_X1 U828 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND3_X1 U829 ( .A1(n1036), .A2(n1158), .A3(n1159), .ZN(n1157) );
NAND2_X1 U830 ( .A1(n1160), .A2(n1161), .ZN(n1156) );
XNOR2_X1 U831 ( .A(KEYINPUT37), .B(n1028), .ZN(n1161) );
INV_X1 U832 ( .A(n1162), .ZN(n1028) );
NAND2_X1 U833 ( .A1(n1163), .A2(n1041), .ZN(n1005) );
INV_X1 U834 ( .A(n1115), .ZN(n1163) );
NAND2_X1 U835 ( .A1(n1160), .A2(n1162), .ZN(n1115) );
AND4_X1 U836 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1009) );
AND4_X1 U837 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1172), .A2(n1173), .ZN(n1166) );
INV_X1 U839 ( .A(n1174), .ZN(n1172) );
NAND3_X1 U840 ( .A1(n1175), .A2(n1176), .A3(n1177), .ZN(n1165) );
INV_X1 U841 ( .A(KEYINPUT38), .ZN(n1177) );
NAND2_X1 U842 ( .A1(n1178), .A2(KEYINPUT38), .ZN(n1164) );
NOR2_X1 U843 ( .A1(n1179), .A2(G952), .ZN(n1099) );
XNOR2_X1 U844 ( .A(n1082), .B(KEYINPUT45), .ZN(n1179) );
XOR2_X1 U845 ( .A(G146), .B(n1173), .Z(G48) );
AND2_X1 U846 ( .A1(n1180), .A2(n1040), .ZN(n1173) );
XOR2_X1 U847 ( .A(G143), .B(n1178), .Z(G45) );
AND2_X1 U848 ( .A1(n1175), .A2(n1044), .ZN(n1178) );
AND4_X1 U849 ( .A1(n1030), .A2(n1036), .A3(n1181), .A4(n1182), .ZN(n1175) );
XNOR2_X1 U850 ( .A(G140), .B(n1174), .ZN(G42) );
NAND4_X1 U851 ( .A1(n1183), .A2(n1040), .A3(n1184), .A4(n1185), .ZN(n1174) );
XNOR2_X1 U852 ( .A(G137), .B(n1171), .ZN(G39) );
NAND4_X1 U853 ( .A1(n1183), .A2(n1186), .A3(n1185), .A4(n1038), .ZN(n1171) );
INV_X1 U854 ( .A(n1034), .ZN(n1185) );
NAND2_X1 U855 ( .A1(n1187), .A2(n1188), .ZN(G36) );
NAND2_X1 U856 ( .A1(G134), .A2(n1170), .ZN(n1188) );
XOR2_X1 U857 ( .A(n1189), .B(KEYINPUT54), .Z(n1187) );
OR2_X1 U858 ( .A1(n1170), .A2(G134), .ZN(n1189) );
NAND2_X1 U859 ( .A1(n1190), .A2(n1041), .ZN(n1170) );
XNOR2_X1 U860 ( .A(G131), .B(n1046), .ZN(G33) );
NAND2_X1 U861 ( .A1(n1040), .A2(n1190), .ZN(n1046) );
NOR4_X1 U862 ( .A1(n1191), .A2(n1034), .A3(n1176), .A4(n1192), .ZN(n1190) );
NAND2_X1 U863 ( .A1(n1193), .A2(n1194), .ZN(n1034) );
XOR2_X1 U864 ( .A(KEYINPUT25), .B(n1031), .Z(n1193) );
INV_X1 U865 ( .A(n1036), .ZN(n1191) );
XNOR2_X1 U866 ( .A(n1169), .B(n1195), .ZN(G30) );
XOR2_X1 U867 ( .A(KEYINPUT6), .B(G128), .Z(n1195) );
NAND2_X1 U868 ( .A1(n1180), .A2(n1041), .ZN(n1169) );
AND3_X1 U869 ( .A1(n1030), .A2(n1038), .A3(n1183), .ZN(n1180) );
NOR3_X1 U870 ( .A1(n1192), .A2(n1037), .A3(n1176), .ZN(n1183) );
XNOR2_X1 U871 ( .A(G101), .B(n1196), .ZN(G3) );
NAND2_X1 U872 ( .A1(KEYINPUT59), .A2(n1154), .ZN(n1196) );
AND3_X1 U873 ( .A1(n1036), .A2(n1160), .A3(n1186), .ZN(n1154) );
XNOR2_X1 U874 ( .A(G125), .B(n1168), .ZN(G27) );
NAND4_X1 U875 ( .A1(n1184), .A2(n1040), .A3(n1030), .A4(n1197), .ZN(n1168) );
NOR4_X1 U876 ( .A1(n1019), .A2(n1037), .A3(n1192), .A4(n1018), .ZN(n1197) );
INV_X1 U877 ( .A(n1182), .ZN(n1192) );
NAND2_X1 U878 ( .A1(n1015), .A2(n1198), .ZN(n1182) );
NAND2_X1 U879 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
INV_X1 U880 ( .A(G900), .ZN(n1200) );
XOR2_X1 U881 ( .A(G122), .B(n1153), .Z(G24) );
AND4_X1 U882 ( .A1(n1030), .A2(n1159), .A3(n1181), .A4(n1162), .ZN(n1153) );
NOR2_X1 U883 ( .A1(n1201), .A2(n1038), .ZN(n1162) );
XNOR2_X1 U884 ( .A(n1152), .B(n1202), .ZN(G21) );
XNOR2_X1 U885 ( .A(KEYINPUT21), .B(n1203), .ZN(n1202) );
AND4_X1 U886 ( .A1(n1030), .A2(n1159), .A3(n1204), .A4(n1186), .ZN(n1152) );
NOR2_X1 U887 ( .A1(n1037), .A2(n1184), .ZN(n1204) );
INV_X1 U888 ( .A(n1201), .ZN(n1037) );
NAND2_X1 U889 ( .A1(n1205), .A2(n1206), .ZN(G18) );
NAND2_X1 U890 ( .A1(G116), .A2(n1207), .ZN(n1206) );
NAND2_X1 U891 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U892 ( .A1(KEYINPUT55), .A2(n1210), .ZN(n1209) );
NAND3_X1 U893 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1205) );
INV_X1 U894 ( .A(KEYINPUT55), .ZN(n1213) );
NAND2_X1 U895 ( .A1(n1148), .A2(n1210), .ZN(n1212) );
INV_X1 U896 ( .A(KEYINPUT23), .ZN(n1210) );
NAND2_X1 U897 ( .A1(n1208), .A2(n1214), .ZN(n1211) );
OR2_X1 U898 ( .A1(G116), .A2(KEYINPUT23), .ZN(n1214) );
INV_X1 U899 ( .A(n1148), .ZN(n1208) );
NAND4_X1 U900 ( .A1(n1030), .A2(n1159), .A3(n1036), .A4(n1041), .ZN(n1148) );
NAND2_X1 U901 ( .A1(n1215), .A2(n1216), .ZN(n1041) );
OR3_X1 U902 ( .A1(n1054), .A2(n1217), .A3(KEYINPUT20), .ZN(n1216) );
NAND2_X1 U903 ( .A1(KEYINPUT20), .A2(n1181), .ZN(n1215) );
NOR2_X1 U904 ( .A1(n1218), .A2(n1054), .ZN(n1181) );
XNOR2_X1 U905 ( .A(n1158), .B(KEYINPUT19), .ZN(n1030) );
XOR2_X1 U906 ( .A(n1219), .B(n1220), .Z(G15) );
XNOR2_X1 U907 ( .A(KEYINPUT12), .B(n1221), .ZN(n1220) );
NAND4_X1 U908 ( .A1(n1222), .A2(n1159), .A3(n1040), .A4(n1158), .ZN(n1219) );
INV_X1 U909 ( .A(n1116), .ZN(n1040) );
NAND2_X1 U910 ( .A1(n1054), .A2(n1223), .ZN(n1116) );
XOR2_X1 U911 ( .A(KEYINPUT62), .B(n1218), .Z(n1223) );
NOR3_X1 U912 ( .A1(n1224), .A2(n1019), .A3(n1018), .ZN(n1159) );
INV_X1 U913 ( .A(n1045), .ZN(n1019) );
INV_X1 U914 ( .A(n1225), .ZN(n1224) );
XNOR2_X1 U915 ( .A(n1036), .B(KEYINPUT58), .ZN(n1222) );
NOR2_X1 U916 ( .A1(n1201), .A2(n1184), .ZN(n1036) );
XNOR2_X1 U917 ( .A(G110), .B(n1226), .ZN(G12) );
NOR2_X1 U918 ( .A1(n1151), .A2(KEYINPUT1), .ZN(n1226) );
AND4_X1 U919 ( .A1(n1186), .A2(n1160), .A3(n1184), .A4(n1201), .ZN(n1151) );
NAND3_X1 U920 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1201) );
NAND2_X1 U921 ( .A1(n1230), .A2(n1101), .ZN(n1229) );
OR3_X1 U922 ( .A1(n1101), .A2(n1230), .A3(G902), .ZN(n1228) );
NOR2_X1 U923 ( .A1(n1105), .A2(G234), .ZN(n1230) );
INV_X1 U924 ( .A(G217), .ZN(n1105) );
XNOR2_X1 U925 ( .A(n1231), .B(n1232), .ZN(n1101) );
XNOR2_X1 U926 ( .A(n1233), .B(n1234), .ZN(n1232) );
XOR2_X1 U927 ( .A(KEYINPUT5), .B(G146), .Z(n1234) );
INV_X1 U928 ( .A(G125), .ZN(n1233) );
XOR2_X1 U929 ( .A(n1235), .B(n1236), .Z(n1231) );
XOR2_X1 U930 ( .A(n1237), .B(n1238), .Z(n1235) );
AND3_X1 U931 ( .A1(G221), .A2(n1082), .A3(G234), .ZN(n1238) );
NAND2_X1 U932 ( .A1(n1239), .A2(KEYINPUT3), .ZN(n1237) );
XNOR2_X1 U933 ( .A(G119), .B(n1240), .ZN(n1239) );
NOR2_X1 U934 ( .A1(G128), .A2(KEYINPUT29), .ZN(n1240) );
NAND2_X1 U935 ( .A1(G217), .A2(G902), .ZN(n1227) );
INV_X1 U936 ( .A(n1038), .ZN(n1184) );
XNOR2_X1 U937 ( .A(n1055), .B(KEYINPUT47), .ZN(n1038) );
XNOR2_X1 U938 ( .A(n1241), .B(n1122), .ZN(n1055) );
INV_X1 U939 ( .A(G472), .ZN(n1122) );
NAND2_X1 U940 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XNOR2_X1 U941 ( .A(n1244), .B(n1121), .ZN(n1242) );
XOR2_X1 U942 ( .A(n1245), .B(n1246), .Z(n1121) );
INV_X1 U943 ( .A(G101), .ZN(n1246) );
NAND2_X1 U944 ( .A1(n1247), .A2(G210), .ZN(n1245) );
NAND2_X1 U945 ( .A1(n1126), .A2(n1125), .ZN(n1244) );
NAND2_X1 U946 ( .A1(n1248), .A2(n1249), .ZN(n1125) );
NAND2_X1 U947 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
INV_X1 U948 ( .A(n1252), .ZN(n1248) );
NAND3_X1 U949 ( .A1(n1252), .A2(n1251), .A3(n1250), .ZN(n1126) );
XNOR2_X1 U950 ( .A(KEYINPUT17), .B(n1253), .ZN(n1250) );
NAND2_X1 U951 ( .A1(G113), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U952 ( .A(n1203), .B(G116), .ZN(n1254) );
NAND2_X1 U953 ( .A1(n1255), .A2(n1221), .ZN(n1251) );
XNOR2_X1 U954 ( .A(G116), .B(G119), .ZN(n1255) );
XNOR2_X1 U955 ( .A(n1256), .B(n1257), .ZN(n1252) );
XNOR2_X1 U956 ( .A(n1144), .B(n1258), .ZN(n1256) );
INV_X1 U957 ( .A(G137), .ZN(n1258) );
AND3_X1 U958 ( .A1(n1044), .A2(n1225), .A3(n1158), .ZN(n1160) );
NOR2_X1 U959 ( .A1(n1032), .A2(n1031), .ZN(n1158) );
NOR2_X1 U960 ( .A1(n1259), .A2(n1051), .ZN(n1031) );
NOR2_X1 U961 ( .A1(n1057), .A2(n1056), .ZN(n1051) );
AND2_X1 U962 ( .A1(n1260), .A2(n1057), .ZN(n1259) );
NAND2_X1 U963 ( .A1(n1261), .A2(n1243), .ZN(n1057) );
XOR2_X1 U964 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U965 ( .A(n1144), .B(n1264), .Z(n1263) );
XNOR2_X1 U966 ( .A(G125), .B(KEYINPUT61), .ZN(n1264) );
NAND3_X1 U967 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1144) );
NAND2_X1 U968 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U969 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XNOR2_X1 U970 ( .A(KEYINPUT0), .B(n1272), .ZN(n1270) );
NAND3_X1 U971 ( .A1(n1273), .A2(n1274), .A3(n1271), .ZN(n1266) );
INV_X1 U972 ( .A(KEYINPUT16), .ZN(n1271) );
NAND2_X1 U973 ( .A1(KEYINPUT16), .A2(n1272), .ZN(n1265) );
INV_X1 U974 ( .A(n1273), .ZN(n1272) );
XOR2_X1 U975 ( .A(n1275), .B(n1141), .Z(n1262) );
XNOR2_X1 U976 ( .A(n1276), .B(n1098), .ZN(n1141) );
XOR2_X1 U977 ( .A(G110), .B(n1277), .Z(n1098) );
XOR2_X1 U978 ( .A(KEYINPUT51), .B(G122), .Z(n1277) );
XNOR2_X1 U979 ( .A(n1278), .B(n1279), .ZN(n1276) );
INV_X1 U980 ( .A(n1094), .ZN(n1279) );
XOR2_X1 U981 ( .A(n1280), .B(n1221), .Z(n1094) );
NAND2_X1 U982 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND2_X1 U983 ( .A1(G116), .A2(n1203), .ZN(n1282) );
XOR2_X1 U984 ( .A(KEYINPUT10), .B(n1283), .Z(n1281) );
NOR2_X1 U985 ( .A1(G116), .A2(n1203), .ZN(n1283) );
INV_X1 U986 ( .A(G119), .ZN(n1203) );
NAND2_X1 U987 ( .A1(KEYINPUT49), .A2(n1096), .ZN(n1278) );
NAND2_X1 U988 ( .A1(KEYINPUT15), .A2(n1145), .ZN(n1275) );
AND2_X1 U989 ( .A1(G224), .A2(n1082), .ZN(n1145) );
XNOR2_X1 U990 ( .A(n1056), .B(KEYINPUT18), .ZN(n1260) );
INV_X1 U991 ( .A(n1146), .ZN(n1056) );
NAND2_X1 U992 ( .A1(G210), .A2(n1284), .ZN(n1146) );
INV_X1 U993 ( .A(n1194), .ZN(n1032) );
NAND2_X1 U994 ( .A1(G214), .A2(n1284), .ZN(n1194) );
NAND2_X1 U995 ( .A1(n1285), .A2(n1243), .ZN(n1284) );
INV_X1 U996 ( .A(G237), .ZN(n1285) );
NAND2_X1 U997 ( .A1(n1015), .A2(n1286), .ZN(n1225) );
NAND2_X1 U998 ( .A1(n1287), .A2(n1199), .ZN(n1286) );
AND3_X1 U999 ( .A1(G953), .A2(n1288), .A3(n1289), .ZN(n1199) );
XNOR2_X1 U1000 ( .A(G902), .B(KEYINPUT44), .ZN(n1289) );
XOR2_X1 U1001 ( .A(n1093), .B(KEYINPUT31), .Z(n1287) );
XNOR2_X1 U1002 ( .A(G898), .B(KEYINPUT34), .ZN(n1093) );
NAND3_X1 U1003 ( .A1(n1288), .A2(n1082), .A3(G952), .ZN(n1015) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1288) );
INV_X1 U1005 ( .A(n1176), .ZN(n1044) );
NAND2_X1 U1006 ( .A1(n1290), .A2(n1045), .ZN(n1176) );
NAND2_X1 U1007 ( .A1(G221), .A2(n1291), .ZN(n1045) );
NAND2_X1 U1008 ( .A1(G234), .A2(n1243), .ZN(n1291) );
XNOR2_X1 U1009 ( .A(n1018), .B(KEYINPUT46), .ZN(n1290) );
XOR2_X1 U1010 ( .A(n1061), .B(n1060), .Z(n1018) );
INV_X1 U1011 ( .A(G469), .ZN(n1060) );
NAND2_X1 U1012 ( .A1(n1292), .A2(n1243), .ZN(n1061) );
XNOR2_X1 U1013 ( .A(n1293), .B(n1294), .ZN(n1292) );
XNOR2_X1 U1014 ( .A(n1295), .B(KEYINPUT32), .ZN(n1294) );
NAND2_X1 U1015 ( .A1(KEYINPUT43), .A2(n1076), .ZN(n1295) );
INV_X1 U1016 ( .A(n1136), .ZN(n1076) );
XOR2_X1 U1017 ( .A(n1273), .B(n1296), .Z(n1136) );
NOR2_X1 U1018 ( .A1(KEYINPUT41), .A2(n1297), .ZN(n1296) );
XNOR2_X1 U1019 ( .A(KEYINPUT4), .B(n1274), .ZN(n1297) );
INV_X1 U1020 ( .A(n1268), .ZN(n1274) );
XOR2_X1 U1021 ( .A(G128), .B(KEYINPUT39), .Z(n1268) );
INV_X1 U1022 ( .A(n1133), .ZN(n1293) );
XNOR2_X1 U1023 ( .A(n1298), .B(n1299), .ZN(n1133) );
XNOR2_X1 U1024 ( .A(n1236), .B(n1300), .ZN(n1299) );
INV_X1 U1025 ( .A(n1096), .ZN(n1300) );
XOR2_X1 U1026 ( .A(G101), .B(n1301), .Z(n1096) );
XOR2_X1 U1027 ( .A(G107), .B(G104), .Z(n1301) );
XOR2_X1 U1028 ( .A(G110), .B(n1075), .Z(n1236) );
XNOR2_X1 U1029 ( .A(G137), .B(n1302), .ZN(n1075) );
XNOR2_X1 U1030 ( .A(n1257), .B(n1303), .ZN(n1298) );
AND2_X1 U1031 ( .A1(n1082), .A2(G227), .ZN(n1303) );
XNOR2_X1 U1032 ( .A(n1304), .B(n1077), .ZN(n1257) );
XOR2_X1 U1033 ( .A(G131), .B(KEYINPUT33), .Z(n1077) );
NAND2_X1 U1034 ( .A1(KEYINPUT11), .A2(n1079), .ZN(n1304) );
INV_X1 U1035 ( .A(n1024), .ZN(n1186) );
NAND2_X1 U1036 ( .A1(n1054), .A2(n1218), .ZN(n1024) );
INV_X1 U1037 ( .A(n1217), .ZN(n1218) );
XOR2_X1 U1038 ( .A(n1053), .B(n1305), .Z(n1217) );
XOR2_X1 U1039 ( .A(KEYINPUT35), .B(KEYINPUT2), .Z(n1305) );
XNOR2_X1 U1040 ( .A(n1306), .B(n1113), .ZN(n1053) );
INV_X1 U1041 ( .A(G475), .ZN(n1113) );
NAND2_X1 U1042 ( .A1(n1111), .A2(n1243), .ZN(n1306) );
XNOR2_X1 U1043 ( .A(n1307), .B(n1308), .ZN(n1111) );
XNOR2_X1 U1044 ( .A(n1273), .B(n1309), .ZN(n1308) );
XOR2_X1 U1045 ( .A(n1310), .B(n1311), .Z(n1309) );
NOR2_X1 U1046 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
XOR2_X1 U1047 ( .A(n1314), .B(KEYINPUT7), .Z(n1313) );
NAND2_X1 U1048 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U1049 ( .A(KEYINPUT24), .B(n1317), .Z(n1316) );
NOR2_X1 U1050 ( .A1(n1317), .A2(n1315), .ZN(n1312) );
XOR2_X1 U1051 ( .A(KEYINPUT63), .B(G104), .Z(n1315) );
XNOR2_X1 U1052 ( .A(n1221), .B(G122), .ZN(n1317) );
INV_X1 U1053 ( .A(G113), .ZN(n1221) );
NAND2_X1 U1054 ( .A1(n1247), .A2(G214), .ZN(n1310) );
NOR2_X1 U1055 ( .A1(G953), .A2(G237), .ZN(n1247) );
XOR2_X1 U1056 ( .A(G143), .B(G146), .Z(n1273) );
XNOR2_X1 U1057 ( .A(G125), .B(n1318), .ZN(n1307) );
XNOR2_X1 U1058 ( .A(n1302), .B(G131), .ZN(n1318) );
INV_X1 U1059 ( .A(G140), .ZN(n1302) );
XNOR2_X1 U1060 ( .A(n1319), .B(n1109), .ZN(n1054) );
INV_X1 U1061 ( .A(G478), .ZN(n1109) );
NAND2_X1 U1062 ( .A1(n1243), .A2(n1107), .ZN(n1319) );
NAND2_X1 U1063 ( .A1(n1320), .A2(n1321), .ZN(n1107) );
OR2_X1 U1064 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1065 ( .A(n1324), .B(KEYINPUT27), .Z(n1320) );
NAND2_X1 U1066 ( .A1(n1323), .A2(n1322), .ZN(n1324) );
NAND3_X1 U1067 ( .A1(G234), .A2(n1082), .A3(G217), .ZN(n1322) );
INV_X1 U1068 ( .A(G953), .ZN(n1082) );
XNOR2_X1 U1069 ( .A(n1325), .B(n1326), .ZN(n1323) );
XNOR2_X1 U1070 ( .A(n1079), .B(n1327), .ZN(n1326) );
XOR2_X1 U1071 ( .A(KEYINPUT36), .B(G143), .Z(n1327) );
INV_X1 U1072 ( .A(G134), .ZN(n1079) );
XOR2_X1 U1073 ( .A(n1328), .B(n1329), .Z(n1325) );
NOR2_X1 U1074 ( .A1(KEYINPUT30), .A2(n1330), .ZN(n1329) );
XNOR2_X1 U1075 ( .A(G122), .B(G116), .ZN(n1330) );
XNOR2_X1 U1076 ( .A(G107), .B(G128), .ZN(n1328) );
INV_X1 U1077 ( .A(G902), .ZN(n1243) );
endmodule


