//Key = 0001101110011011010110000011101110100000111111011011100110011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373;

XNOR2_X1 U764 ( .A(G107), .B(n1060), .ZN(G9) );
NOR2_X1 U765 ( .A1(n1061), .A2(KEYINPUT1), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1062), .A2(n1063), .ZN(G75) );
NOR4_X1 U767 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1063) );
NOR2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U770 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U771 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NOR2_X1 U772 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U773 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR2_X1 U774 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U775 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR2_X1 U776 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR2_X1 U777 ( .A1(n1086), .A2(n1087), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U779 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR3_X1 U780 ( .A1(n1087), .A2(n1092), .A3(n1081), .ZN(n1074) );
NOR3_X1 U781 ( .A1(n1087), .A2(n1093), .A3(n1081), .ZN(n1070) );
NOR3_X1 U782 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
AND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR3_X1 U784 ( .A1(n1099), .A2(n1073), .A3(n1100), .ZN(n1095) );
NOR2_X1 U785 ( .A1(n1077), .A2(n1101), .ZN(n1094) );
XNOR2_X1 U786 ( .A(KEYINPUT51), .B(n1102), .ZN(n1065) );
NAND3_X1 U787 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1064) );
NAND3_X1 U788 ( .A1(n1106), .A2(n1099), .A3(n1107), .ZN(n1105) );
INV_X1 U789 ( .A(KEYINPUT41), .ZN(n1099) );
OR4_X1 U790 ( .A1(n1100), .A2(n1069), .A3(n1081), .A4(n1073), .ZN(n1106) );
INV_X1 U791 ( .A(n1108), .ZN(n1073) );
XOR2_X1 U792 ( .A(n1109), .B(KEYINPUT40), .Z(n1100) );
AND3_X1 U793 ( .A1(n1103), .A2(n1104), .A3(n1110), .ZN(n1062) );
NAND4_X1 U794 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1103) );
NOR4_X1 U795 ( .A1(n1115), .A2(n1116), .A3(n1081), .A4(n1117), .ZN(n1114) );
XNOR2_X1 U796 ( .A(n1118), .B(n1119), .ZN(n1117) );
NOR2_X1 U797 ( .A1(KEYINPUT39), .A2(n1120), .ZN(n1119) );
INV_X1 U798 ( .A(n1121), .ZN(n1081) );
XOR2_X1 U799 ( .A(n1122), .B(n1123), .Z(n1116) );
XNOR2_X1 U800 ( .A(KEYINPUT58), .B(n1124), .ZN(n1123) );
NAND2_X1 U801 ( .A1(n1125), .A2(n1126), .ZN(n1122) );
XOR2_X1 U802 ( .A(KEYINPUT5), .B(KEYINPUT45), .Z(n1125) );
XOR2_X1 U803 ( .A(n1127), .B(KEYINPUT29), .Z(n1113) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1112) );
XNOR2_X1 U805 ( .A(n1130), .B(n1131), .ZN(n1111) );
NAND2_X1 U806 ( .A1(KEYINPUT48), .A2(n1132), .ZN(n1130) );
INV_X1 U807 ( .A(n1133), .ZN(n1132) );
XOR2_X1 U808 ( .A(n1134), .B(n1135), .Z(G72) );
NOR2_X1 U809 ( .A1(n1136), .A2(n1104), .ZN(n1135) );
AND2_X1 U810 ( .A1(G227), .A2(G900), .ZN(n1136) );
NAND2_X1 U811 ( .A1(n1137), .A2(n1138), .ZN(n1134) );
NAND2_X1 U812 ( .A1(n1139), .A2(n1104), .ZN(n1138) );
XOR2_X1 U813 ( .A(n1102), .B(n1140), .Z(n1139) );
NAND3_X1 U814 ( .A1(G900), .A2(n1140), .A3(G953), .ZN(n1137) );
XNOR2_X1 U815 ( .A(n1141), .B(n1142), .ZN(n1140) );
XOR2_X1 U816 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U817 ( .A(n1145), .B(n1146), .ZN(n1144) );
NAND2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
XNOR2_X1 U819 ( .A(KEYINPUT56), .B(KEYINPUT4), .ZN(n1147) );
XNOR2_X1 U820 ( .A(G137), .B(KEYINPUT38), .ZN(n1143) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(n1141) );
XNOR2_X1 U822 ( .A(n1151), .B(n1152), .ZN(n1149) );
NOR2_X1 U823 ( .A1(G140), .A2(KEYINPUT13), .ZN(n1152) );
NAND2_X1 U824 ( .A1(n1153), .A2(n1154), .ZN(G69) );
NAND2_X1 U825 ( .A1(n1155), .A2(n1104), .ZN(n1154) );
XNOR2_X1 U826 ( .A(n1156), .B(n1067), .ZN(n1155) );
NAND2_X1 U827 ( .A1(n1157), .A2(G953), .ZN(n1153) );
NAND2_X1 U828 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U829 ( .A1(n1156), .A2(n1160), .ZN(n1159) );
NAND2_X1 U830 ( .A1(G224), .A2(n1161), .ZN(n1158) );
NAND2_X1 U831 ( .A1(G898), .A2(n1156), .ZN(n1161) );
NAND2_X1 U832 ( .A1(n1162), .A2(n1163), .ZN(n1156) );
NAND2_X1 U833 ( .A1(G953), .A2(n1164), .ZN(n1163) );
XOR2_X1 U834 ( .A(n1165), .B(n1166), .Z(n1162) );
NOR2_X1 U835 ( .A1(KEYINPUT9), .A2(n1167), .ZN(n1165) );
XNOR2_X1 U836 ( .A(n1168), .B(n1169), .ZN(n1167) );
NOR2_X1 U837 ( .A1(KEYINPUT23), .A2(n1170), .ZN(n1169) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(G66) );
NOR3_X1 U839 ( .A1(n1128), .A2(n1173), .A3(n1174), .ZN(n1172) );
NOR3_X1 U840 ( .A1(n1175), .A2(n1129), .A3(n1176), .ZN(n1174) );
NOR2_X1 U841 ( .A1(n1177), .A2(n1178), .ZN(n1173) );
NOR2_X1 U842 ( .A1(n1179), .A2(n1129), .ZN(n1177) );
NOR2_X1 U843 ( .A1(n1102), .A2(n1067), .ZN(n1179) );
NOR2_X1 U844 ( .A1(n1171), .A2(n1180), .ZN(G63) );
XOR2_X1 U845 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1176), .ZN(n1182) );
INV_X1 U847 ( .A(G478), .ZN(n1183) );
NOR2_X1 U848 ( .A1(n1171), .A2(n1184), .ZN(G60) );
XNOR2_X1 U849 ( .A(n1185), .B(n1186), .ZN(n1184) );
NOR2_X1 U850 ( .A1(n1124), .A2(n1176), .ZN(n1186) );
XOR2_X1 U851 ( .A(G104), .B(n1187), .Z(G6) );
NOR2_X1 U852 ( .A1(n1171), .A2(n1188), .ZN(G57) );
XOR2_X1 U853 ( .A(n1189), .B(n1190), .Z(n1188) );
XOR2_X1 U854 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U855 ( .A(n1193), .B(n1194), .Z(n1189) );
NOR2_X1 U856 ( .A1(n1120), .A2(n1176), .ZN(n1194) );
NAND2_X1 U857 ( .A1(n1195), .A2(KEYINPUT28), .ZN(n1193) );
XNOR2_X1 U858 ( .A(n1196), .B(n1197), .ZN(n1195) );
NAND2_X1 U859 ( .A1(KEYINPUT43), .A2(n1198), .ZN(n1196) );
NOR2_X1 U860 ( .A1(n1199), .A2(n1200), .ZN(G54) );
XOR2_X1 U861 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U862 ( .A(n1203), .B(n1204), .Z(n1202) );
NOR2_X1 U863 ( .A1(n1205), .A2(n1176), .ZN(n1204) );
NOR2_X1 U864 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
XOR2_X1 U865 ( .A(n1208), .B(KEYINPUT11), .Z(n1207) );
NAND2_X1 U866 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U867 ( .A(KEYINPUT49), .B(n1211), .Z(n1209) );
XOR2_X1 U868 ( .A(n1212), .B(KEYINPUT2), .Z(n1199) );
NAND2_X1 U869 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
OR3_X1 U870 ( .A1(n1110), .A2(n1104), .A3(KEYINPUT60), .ZN(n1214) );
INV_X1 U871 ( .A(G952), .ZN(n1110) );
NAND2_X1 U872 ( .A1(n1171), .A2(KEYINPUT60), .ZN(n1213) );
NOR2_X1 U873 ( .A1(n1171), .A2(n1215), .ZN(G51) );
XOR2_X1 U874 ( .A(n1216), .B(n1217), .Z(n1215) );
NOR2_X1 U875 ( .A1(n1133), .A2(n1176), .ZN(n1217) );
NAND2_X1 U876 ( .A1(G902), .A2(n1218), .ZN(n1176) );
OR2_X1 U877 ( .A1(n1067), .A2(n1102), .ZN(n1218) );
NAND4_X1 U878 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1102) );
NOR4_X1 U879 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1222) );
INV_X1 U880 ( .A(n1227), .ZN(n1226) );
INV_X1 U881 ( .A(n1228), .ZN(n1225) );
OR2_X1 U882 ( .A1(n1229), .A2(n1230), .ZN(n1221) );
NAND3_X1 U883 ( .A1(n1231), .A2(n1232), .A3(n1107), .ZN(n1219) );
NAND2_X1 U884 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND3_X1 U885 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1233) );
XOR2_X1 U886 ( .A(KEYINPUT21), .B(n1089), .Z(n1235) );
NAND4_X1 U887 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1067) );
NOR4_X1 U888 ( .A1(n1061), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1241) );
AND3_X1 U889 ( .A1(n1237), .A2(n1108), .A3(n1245), .ZN(n1061) );
NOR2_X1 U890 ( .A1(n1187), .A2(n1246), .ZN(n1240) );
NOR2_X1 U891 ( .A1(n1230), .A2(n1247), .ZN(n1246) );
AND3_X1 U892 ( .A1(n1245), .A2(n1108), .A3(n1109), .ZN(n1187) );
NAND2_X1 U893 ( .A1(n1248), .A2(KEYINPUT15), .ZN(n1216) );
XOR2_X1 U894 ( .A(n1249), .B(n1250), .Z(n1248) );
XNOR2_X1 U895 ( .A(n1146), .B(n1251), .ZN(n1250) );
NOR2_X1 U896 ( .A1(KEYINPUT33), .A2(n1151), .ZN(n1251) );
XOR2_X1 U897 ( .A(n1252), .B(n1253), .Z(n1249) );
NOR2_X1 U898 ( .A1(KEYINPUT24), .A2(n1254), .ZN(n1253) );
NOR2_X1 U899 ( .A1(n1104), .A2(G952), .ZN(n1171) );
XNOR2_X1 U900 ( .A(G146), .B(n1255), .ZN(G48) );
NAND2_X1 U901 ( .A1(KEYINPUT7), .A2(n1224), .ZN(n1255) );
NOR4_X1 U902 ( .A1(n1256), .A2(n1234), .A3(n1230), .A4(n1097), .ZN(n1224) );
XNOR2_X1 U903 ( .A(G143), .B(n1257), .ZN(G45) );
NAND3_X1 U904 ( .A1(KEYINPUT44), .A2(n1083), .A3(n1258), .ZN(n1257) );
XOR2_X1 U905 ( .A(n1229), .B(KEYINPUT14), .Z(n1258) );
NAND4_X1 U906 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1231), .ZN(n1229) );
XNOR2_X1 U907 ( .A(G140), .B(n1262), .ZN(G42) );
NAND2_X1 U908 ( .A1(KEYINPUT8), .A2(n1223), .ZN(n1262) );
NOR4_X1 U909 ( .A1(n1234), .A2(n1087), .A3(n1263), .A4(n1256), .ZN(n1223) );
XNOR2_X1 U910 ( .A(G137), .B(n1220), .ZN(G39) );
NAND4_X1 U911 ( .A1(n1260), .A2(n1107), .A3(n1098), .A4(n1263), .ZN(n1220) );
XOR2_X1 U912 ( .A(n1264), .B(n1265), .Z(G36) );
NAND2_X1 U913 ( .A1(KEYINPUT32), .A2(G134), .ZN(n1265) );
NAND4_X1 U914 ( .A1(n1266), .A2(n1260), .A3(n1107), .A4(n1237), .ZN(n1264) );
XNOR2_X1 U915 ( .A(n1231), .B(KEYINPUT47), .ZN(n1266) );
XNOR2_X1 U916 ( .A(n1267), .B(n1148), .ZN(G33) );
NAND2_X1 U917 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND4_X1 U918 ( .A1(n1270), .A2(n1231), .A3(KEYINPUT62), .A4(n1087), .ZN(n1269) );
INV_X1 U919 ( .A(n1234), .ZN(n1270) );
OR4_X1 U920 ( .A1(n1101), .A2(KEYINPUT62), .A3(n1234), .A4(n1087), .ZN(n1268) );
INV_X1 U921 ( .A(n1107), .ZN(n1087) );
NOR2_X1 U922 ( .A1(n1084), .A2(n1115), .ZN(n1107) );
INV_X1 U923 ( .A(n1085), .ZN(n1115) );
NAND2_X1 U924 ( .A1(n1260), .A2(n1109), .ZN(n1234) );
INV_X1 U925 ( .A(n1231), .ZN(n1101) );
XOR2_X1 U926 ( .A(G128), .B(n1271), .Z(G30) );
NOR2_X1 U927 ( .A1(KEYINPUT18), .A2(n1227), .ZN(n1271) );
NAND3_X1 U928 ( .A1(n1272), .A2(n1260), .A3(n1273), .ZN(n1227) );
NOR3_X1 U929 ( .A1(n1092), .A2(n1097), .A3(n1230), .ZN(n1273) );
AND2_X1 U930 ( .A1(n1089), .A2(n1236), .ZN(n1260) );
XNOR2_X1 U931 ( .A(G101), .B(n1238), .ZN(G3) );
NAND3_X1 U932 ( .A1(n1274), .A2(n1245), .A3(n1231), .ZN(n1238) );
XNOR2_X1 U933 ( .A(G125), .B(n1228), .ZN(G27) );
NAND4_X1 U934 ( .A1(n1272), .A2(n1121), .A3(n1109), .A4(n1275), .ZN(n1228) );
AND3_X1 U935 ( .A1(n1097), .A2(n1236), .A3(n1083), .ZN(n1275) );
NAND2_X1 U936 ( .A1(n1276), .A2(n1069), .ZN(n1236) );
NAND4_X1 U937 ( .A1(G953), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1276) );
INV_X1 U938 ( .A(G900), .ZN(n1279) );
XNOR2_X1 U939 ( .A(KEYINPUT10), .B(n1280), .ZN(n1277) );
XNOR2_X1 U940 ( .A(G122), .B(n1239), .ZN(G24) );
NAND4_X1 U941 ( .A1(n1259), .A2(n1281), .A3(n1261), .A4(n1108), .ZN(n1239) );
NOR2_X1 U942 ( .A1(n1263), .A2(n1272), .ZN(n1108) );
XOR2_X1 U943 ( .A(G119), .B(n1244), .Z(G21) );
AND3_X1 U944 ( .A1(n1098), .A2(n1263), .A3(n1281), .ZN(n1244) );
XNOR2_X1 U945 ( .A(G116), .B(n1282), .ZN(G18) );
NAND2_X1 U946 ( .A1(KEYINPUT17), .A2(n1243), .ZN(n1282) );
AND3_X1 U947 ( .A1(n1281), .A2(n1237), .A3(n1231), .ZN(n1243) );
INV_X1 U948 ( .A(n1092), .ZN(n1237) );
NAND2_X1 U949 ( .A1(n1261), .A2(n1283), .ZN(n1092) );
AND3_X1 U950 ( .A1(n1083), .A2(n1284), .A3(n1121), .ZN(n1281) );
XNOR2_X1 U951 ( .A(G113), .B(n1285), .ZN(G15) );
NAND3_X1 U952 ( .A1(KEYINPUT27), .A2(n1083), .A3(n1286), .ZN(n1285) );
XOR2_X1 U953 ( .A(n1247), .B(KEYINPUT31), .Z(n1286) );
NAND4_X1 U954 ( .A1(n1109), .A2(n1231), .A3(n1121), .A4(n1284), .ZN(n1247) );
NOR2_X1 U955 ( .A1(n1090), .A2(n1287), .ZN(n1121) );
INV_X1 U956 ( .A(n1091), .ZN(n1287) );
NOR2_X1 U957 ( .A1(n1097), .A2(n1272), .ZN(n1231) );
INV_X1 U958 ( .A(n1256), .ZN(n1272) );
NOR2_X1 U959 ( .A1(n1283), .A2(n1261), .ZN(n1109) );
NAND2_X1 U960 ( .A1(n1288), .A2(n1289), .ZN(G12) );
NAND2_X1 U961 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U962 ( .A1(n1292), .A2(n1293), .ZN(n1290) );
NAND2_X1 U963 ( .A1(KEYINPUT57), .A2(n1294), .ZN(n1293) );
NAND3_X1 U964 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1288) );
INV_X1 U965 ( .A(KEYINPUT57), .ZN(n1297) );
NAND2_X1 U966 ( .A1(n1242), .A2(n1294), .ZN(n1296) );
INV_X1 U967 ( .A(n1292), .ZN(n1242) );
NAND2_X1 U968 ( .A1(n1298), .A2(n1292), .ZN(n1295) );
NAND3_X1 U969 ( .A1(n1097), .A2(n1245), .A3(n1098), .ZN(n1292) );
NOR2_X1 U970 ( .A1(n1077), .A2(n1256), .ZN(n1098) );
XNOR2_X1 U971 ( .A(n1299), .B(n1128), .ZN(n1256) );
NOR2_X1 U972 ( .A1(n1178), .A2(G902), .ZN(n1128) );
INV_X1 U973 ( .A(n1175), .ZN(n1178) );
XNOR2_X1 U974 ( .A(n1300), .B(n1301), .ZN(n1175) );
XOR2_X1 U975 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U976 ( .A(n1304), .B(n1291), .ZN(n1303) );
NAND2_X1 U977 ( .A1(KEYINPUT19), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U978 ( .A(n1306), .B(n1307), .ZN(n1305) );
XNOR2_X1 U979 ( .A(n1308), .B(n1309), .ZN(n1307) );
NOR2_X1 U980 ( .A1(KEYINPUT36), .A2(n1146), .ZN(n1309) );
NOR2_X1 U981 ( .A1(G146), .A2(KEYINPUT22), .ZN(n1308) );
NAND3_X1 U982 ( .A1(n1310), .A2(G221), .A3(KEYINPUT50), .ZN(n1302) );
XOR2_X1 U983 ( .A(n1311), .B(n1312), .Z(n1300) );
XOR2_X1 U984 ( .A(KEYINPUT34), .B(G137), .Z(n1312) );
XNOR2_X1 U985 ( .A(G119), .B(G128), .ZN(n1311) );
NAND2_X1 U986 ( .A1(KEYINPUT61), .A2(n1129), .ZN(n1299) );
NAND2_X1 U987 ( .A1(G217), .A2(n1313), .ZN(n1129) );
INV_X1 U988 ( .A(n1274), .ZN(n1077) );
NOR2_X1 U989 ( .A1(n1261), .A2(n1259), .ZN(n1274) );
INV_X1 U990 ( .A(n1283), .ZN(n1259) );
XOR2_X1 U991 ( .A(n1314), .B(n1124), .Z(n1283) );
INV_X1 U992 ( .A(G475), .ZN(n1124) );
NAND2_X1 U993 ( .A1(KEYINPUT42), .A2(n1126), .ZN(n1314) );
NAND2_X1 U994 ( .A1(n1185), .A2(n1280), .ZN(n1126) );
XNOR2_X1 U995 ( .A(n1315), .B(n1316), .ZN(n1185) );
XOR2_X1 U996 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U997 ( .A(G122), .B(G113), .Z(n1318) );
XNOR2_X1 U998 ( .A(n1148), .B(G125), .ZN(n1317) );
INV_X1 U999 ( .A(G131), .ZN(n1148) );
XOR2_X1 U1000 ( .A(n1319), .B(n1320), .Z(n1315) );
XNOR2_X1 U1001 ( .A(n1321), .B(n1322), .ZN(n1320) );
INV_X1 U1002 ( .A(n1306), .ZN(n1321) );
XOR2_X1 U1003 ( .A(G140), .B(KEYINPUT46), .Z(n1306) );
XNOR2_X1 U1004 ( .A(G104), .B(n1323), .ZN(n1319) );
AND3_X1 U1005 ( .A1(G214), .A2(n1104), .A3(n1324), .ZN(n1323) );
XOR2_X1 U1006 ( .A(n1127), .B(KEYINPUT12), .Z(n1261) );
XNOR2_X1 U1007 ( .A(G478), .B(n1325), .ZN(n1127) );
NOR2_X1 U1008 ( .A1(G902), .A2(n1181), .ZN(n1325) );
XOR2_X1 U1009 ( .A(n1326), .B(n1327), .Z(n1181) );
NOR2_X1 U1010 ( .A1(KEYINPUT16), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1011 ( .A(n1329), .B(n1330), .Z(n1328) );
XNOR2_X1 U1012 ( .A(n1331), .B(n1332), .ZN(n1330) );
XNOR2_X1 U1013 ( .A(n1333), .B(n1334), .ZN(n1332) );
NOR2_X1 U1014 ( .A1(G128), .A2(KEYINPUT25), .ZN(n1334) );
NAND2_X1 U1015 ( .A1(KEYINPUT26), .A2(n1150), .ZN(n1333) );
XOR2_X1 U1016 ( .A(n1335), .B(n1336), .Z(n1329) );
XOR2_X1 U1017 ( .A(KEYINPUT63), .B(G143), .Z(n1336) );
XNOR2_X1 U1018 ( .A(G107), .B(G122), .ZN(n1335) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1310), .ZN(n1326) );
AND2_X1 U1020 ( .A1(G234), .A2(n1104), .ZN(n1310) );
AND3_X1 U1021 ( .A1(n1089), .A2(n1284), .A3(n1083), .ZN(n1245) );
INV_X1 U1022 ( .A(n1230), .ZN(n1083) );
NAND2_X1 U1023 ( .A1(n1084), .A2(n1085), .ZN(n1230) );
NAND2_X1 U1024 ( .A1(G214), .A2(n1337), .ZN(n1085) );
XOR2_X1 U1025 ( .A(n1131), .B(n1133), .Z(n1084) );
NAND2_X1 U1026 ( .A1(G210), .A2(n1337), .ZN(n1133) );
NAND2_X1 U1027 ( .A1(n1324), .A2(n1280), .ZN(n1337) );
NAND2_X1 U1028 ( .A1(n1338), .A2(n1280), .ZN(n1131) );
XOR2_X1 U1029 ( .A(n1339), .B(n1340), .Z(n1338) );
XNOR2_X1 U1030 ( .A(n1146), .B(n1254), .ZN(n1340) );
NOR2_X1 U1031 ( .A1(n1160), .A2(G953), .ZN(n1254) );
INV_X1 U1032 ( .A(G224), .ZN(n1160) );
INV_X1 U1033 ( .A(G125), .ZN(n1146) );
XNOR2_X1 U1034 ( .A(n1252), .B(n1341), .ZN(n1339) );
XOR2_X1 U1035 ( .A(n1342), .B(n1166), .Z(n1252) );
XNOR2_X1 U1036 ( .A(n1291), .B(G122), .ZN(n1166) );
INV_X1 U1037 ( .A(G110), .ZN(n1291) );
XNOR2_X1 U1038 ( .A(n1343), .B(n1344), .ZN(n1342) );
INV_X1 U1039 ( .A(n1168), .ZN(n1344) );
NAND2_X1 U1040 ( .A1(KEYINPUT30), .A2(n1345), .ZN(n1343) );
INV_X1 U1041 ( .A(n1170), .ZN(n1345) );
XNOR2_X1 U1042 ( .A(n1346), .B(n1347), .ZN(n1170) );
NAND2_X1 U1043 ( .A1(KEYINPUT20), .A2(n1197), .ZN(n1346) );
NAND2_X1 U1044 ( .A1(n1069), .A2(n1348), .ZN(n1284) );
NAND4_X1 U1045 ( .A1(G953), .A2(G902), .A3(n1278), .A4(n1164), .ZN(n1348) );
INV_X1 U1046 ( .A(G898), .ZN(n1164) );
NAND3_X1 U1047 ( .A1(n1278), .A2(n1104), .A3(G952), .ZN(n1069) );
NAND2_X1 U1048 ( .A1(G237), .A2(G234), .ZN(n1278) );
AND2_X1 U1049 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U1050 ( .A1(G221), .A2(n1313), .ZN(n1091) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1280), .ZN(n1313) );
XOR2_X1 U1052 ( .A(n1349), .B(n1205), .Z(n1090) );
INV_X1 U1053 ( .A(G469), .ZN(n1205) );
NAND2_X1 U1054 ( .A1(n1350), .A2(n1280), .ZN(n1349) );
XOR2_X1 U1055 ( .A(n1351), .B(n1201), .Z(n1350) );
XOR2_X1 U1056 ( .A(n1347), .B(n1352), .Z(n1201) );
XNOR2_X1 U1057 ( .A(n1197), .B(n1192), .ZN(n1352) );
INV_X1 U1058 ( .A(G101), .ZN(n1197) );
XNOR2_X1 U1059 ( .A(G104), .B(n1353), .ZN(n1347) );
INV_X1 U1060 ( .A(G107), .ZN(n1353) );
NAND2_X1 U1061 ( .A1(n1354), .A2(n1355), .ZN(n1351) );
INV_X1 U1062 ( .A(n1206), .ZN(n1355) );
NOR2_X1 U1063 ( .A1(n1210), .A2(n1211), .ZN(n1206) );
NAND2_X1 U1064 ( .A1(n1211), .A2(n1210), .ZN(n1354) );
NAND2_X1 U1065 ( .A1(G227), .A2(n1104), .ZN(n1210) );
XNOR2_X1 U1066 ( .A(G110), .B(n1356), .ZN(n1211) );
INV_X1 U1067 ( .A(G140), .ZN(n1356) );
INV_X1 U1068 ( .A(n1263), .ZN(n1097) );
XOR2_X1 U1069 ( .A(n1118), .B(n1120), .Z(n1263) );
INV_X1 U1070 ( .A(G472), .ZN(n1120) );
NAND2_X1 U1071 ( .A1(n1357), .A2(n1280), .ZN(n1118) );
INV_X1 U1072 ( .A(G902), .ZN(n1280) );
XOR2_X1 U1073 ( .A(n1358), .B(n1359), .Z(n1357) );
XOR2_X1 U1074 ( .A(n1360), .B(n1191), .Z(n1359) );
XNOR2_X1 U1075 ( .A(n1168), .B(KEYINPUT59), .ZN(n1191) );
XNOR2_X1 U1076 ( .A(n1361), .B(n1331), .ZN(n1168) );
XOR2_X1 U1077 ( .A(G116), .B(KEYINPUT55), .Z(n1331) );
XNOR2_X1 U1078 ( .A(G113), .B(G119), .ZN(n1361) );
NAND2_X1 U1079 ( .A1(KEYINPUT52), .A2(n1362), .ZN(n1360) );
XNOR2_X1 U1080 ( .A(n1198), .B(n1363), .ZN(n1362) );
XNOR2_X1 U1081 ( .A(G101), .B(KEYINPUT0), .ZN(n1363) );
AND3_X1 U1082 ( .A1(n1324), .A2(n1104), .A3(G210), .ZN(n1198) );
INV_X1 U1083 ( .A(G953), .ZN(n1104) );
INV_X1 U1084 ( .A(G237), .ZN(n1324) );
NAND2_X1 U1085 ( .A1(n1364), .A2(n1365), .ZN(n1358) );
NAND3_X1 U1086 ( .A1(n1366), .A2(n1151), .A3(n1367), .ZN(n1365) );
INV_X1 U1087 ( .A(KEYINPUT6), .ZN(n1367) );
NAND2_X1 U1088 ( .A1(n1192), .A2(KEYINPUT6), .ZN(n1364) );
XNOR2_X1 U1089 ( .A(n1341), .B(n1366), .ZN(n1192) );
XNOR2_X1 U1090 ( .A(n1368), .B(KEYINPUT53), .ZN(n1366) );
NAND2_X1 U1091 ( .A1(n1369), .A2(n1370), .ZN(n1368) );
NAND2_X1 U1092 ( .A1(G131), .A2(n1371), .ZN(n1370) );
XOR2_X1 U1093 ( .A(n1372), .B(KEYINPUT35), .Z(n1369) );
OR2_X1 U1094 ( .A1(n1371), .A2(G131), .ZN(n1372) );
XOR2_X1 U1095 ( .A(n1150), .B(n1373), .Z(n1371) );
NOR2_X1 U1096 ( .A1(G137), .A2(KEYINPUT54), .ZN(n1373) );
XOR2_X1 U1097 ( .A(G134), .B(KEYINPUT3), .Z(n1150) );
INV_X1 U1098 ( .A(n1151), .ZN(n1341) );
XOR2_X1 U1099 ( .A(G128), .B(n1322), .Z(n1151) );
XOR2_X1 U1100 ( .A(G143), .B(G146), .Z(n1322) );
NAND2_X1 U1101 ( .A1(G110), .A2(n1294), .ZN(n1298) );
INV_X1 U1102 ( .A(KEYINPUT37), .ZN(n1294) );
endmodule


