//Key = 1010011011001111111011111000000000101111111010011000101110110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322;

XOR2_X1 U720 ( .A(G107), .B(n1001), .Z(G9) );
NOR2_X1 U721 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NAND4_X1 U722 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(G75) );
INV_X1 U723 ( .A(n1008), .ZN(n1007) );
NAND2_X1 U724 ( .A1(n1009), .A2(n1010), .ZN(n1006) );
NOR4_X1 U725 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
INV_X1 U726 ( .A(n1015), .ZN(n1014) );
NOR2_X1 U727 ( .A1(G469), .A2(n1016), .ZN(n1013) );
NOR4_X1 U728 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1009) );
XOR2_X1 U729 ( .A(n1021), .B(n1022), .Z(n1020) );
XOR2_X1 U730 ( .A(n1023), .B(n1024), .Z(n1019) );
XOR2_X1 U731 ( .A(KEYINPUT10), .B(n1025), .Z(n1018) );
AND2_X1 U732 ( .A1(n1016), .A2(G469), .ZN(n1025) );
NAND2_X1 U733 ( .A1(G952), .A2(n1026), .ZN(n1005) );
NAND3_X1 U734 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
NAND2_X1 U735 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
NAND2_X1 U736 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND3_X1 U737 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NAND2_X1 U738 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NAND2_X1 U739 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U740 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U741 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U742 ( .A1(n1015), .A2(n1045), .ZN(n1037) );
NAND2_X1 U743 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U744 ( .A1(n1012), .A2(n1048), .ZN(n1047) );
INV_X1 U745 ( .A(n1049), .ZN(n1012) );
NAND3_X1 U746 ( .A1(n1015), .A2(n1050), .A3(n1039), .ZN(n1032) );
NAND2_X1 U747 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND3_X1 U748 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
NAND2_X1 U749 ( .A1(n1011), .A2(n1056), .ZN(n1054) );
INV_X1 U750 ( .A(n1057), .ZN(n1011) );
NAND3_X1 U751 ( .A1(n1002), .A2(n1058), .A3(n1057), .ZN(n1053) );
INV_X1 U752 ( .A(n1059), .ZN(n1002) );
NAND2_X1 U753 ( .A1(n1034), .A2(n1060), .ZN(n1051) );
INV_X1 U754 ( .A(n1061), .ZN(n1030) );
OR2_X1 U755 ( .A1(G953), .A2(KEYINPUT55), .ZN(n1027) );
NAND2_X1 U756 ( .A1(KEYINPUT55), .A2(G953), .ZN(n1004) );
NAND2_X1 U757 ( .A1(n1062), .A2(n1063), .ZN(G72) );
NAND2_X1 U758 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U759 ( .A1(G953), .A2(n1066), .ZN(n1064) );
NAND2_X1 U760 ( .A1(G900), .A2(G227), .ZN(n1066) );
NAND2_X1 U761 ( .A1(n1067), .A2(n1068), .ZN(n1062) );
NAND2_X1 U762 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
OR2_X1 U763 ( .A1(n1071), .A2(G227), .ZN(n1070) );
INV_X1 U764 ( .A(n1072), .ZN(n1069) );
INV_X1 U765 ( .A(n1065), .ZN(n1067) );
NAND2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1065) );
NAND2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
OR2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U769 ( .A(KEYINPUT58), .B(n1079), .Z(n1073) );
NOR4_X1 U770 ( .A1(n1075), .A2(n1072), .A3(n1078), .A4(n1077), .ZN(n1079) );
XNOR2_X1 U771 ( .A(n1080), .B(KEYINPUT32), .ZN(n1077) );
NAND2_X1 U772 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U773 ( .A1(n1082), .A2(n1081), .ZN(n1078) );
XOR2_X1 U774 ( .A(n1083), .B(n1084), .Z(n1081) );
XNOR2_X1 U775 ( .A(n1085), .B(n1086), .ZN(n1082) );
XOR2_X1 U776 ( .A(n1087), .B(n1088), .Z(n1085) );
NAND2_X1 U777 ( .A1(KEYINPUT24), .A2(n1089), .ZN(n1087) );
NOR2_X1 U778 ( .A1(n1071), .A2(G900), .ZN(n1072) );
NOR2_X1 U779 ( .A1(n1090), .A2(G953), .ZN(n1075) );
XOR2_X1 U780 ( .A(n1091), .B(n1092), .Z(G69) );
XOR2_X1 U781 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U783 ( .A1(G953), .A2(n1097), .ZN(n1096) );
XOR2_X1 U784 ( .A(KEYINPUT7), .B(n1098), .Z(n1095) );
NAND2_X1 U785 ( .A1(n1099), .A2(n1071), .ZN(n1093) );
XOR2_X1 U786 ( .A(n1100), .B(KEYINPUT60), .Z(n1099) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U788 ( .A1(n1103), .A2(n1071), .ZN(n1091) );
NOR2_X1 U789 ( .A1(n1104), .A2(n1097), .ZN(n1103) );
NOR2_X1 U790 ( .A1(n1008), .A2(n1105), .ZN(G66) );
XOR2_X1 U791 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR2_X1 U793 ( .A1(n1008), .A2(n1110), .ZN(G63) );
XOR2_X1 U794 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1109), .ZN(n1111) );
INV_X1 U796 ( .A(G478), .ZN(n1113) );
NOR2_X1 U797 ( .A1(n1008), .A2(n1114), .ZN(G60) );
NOR3_X1 U798 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
NOR3_X1 U799 ( .A1(n1118), .A2(n1023), .A3(n1109), .ZN(n1117) );
NOR2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1116) );
INV_X1 U801 ( .A(n1118), .ZN(n1120) );
NOR2_X1 U802 ( .A1(n1029), .A2(n1023), .ZN(n1119) );
INV_X1 U803 ( .A(n1121), .ZN(n1029) );
XNOR2_X1 U804 ( .A(G104), .B(n1122), .ZN(G6) );
NOR2_X1 U805 ( .A1(n1008), .A2(n1123), .ZN(G57) );
XOR2_X1 U806 ( .A(n1124), .B(n1125), .Z(n1123) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U808 ( .A(n1128), .B(n1129), .Z(n1127) );
NAND2_X1 U809 ( .A1(KEYINPUT40), .A2(n1130), .ZN(n1128) );
XOR2_X1 U810 ( .A(n1131), .B(n1132), .Z(n1124) );
XOR2_X1 U811 ( .A(KEYINPUT44), .B(n1133), .Z(n1132) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1109), .ZN(n1133) );
INV_X1 U813 ( .A(G472), .ZN(n1134) );
NAND2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(n1131) );
NAND2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U816 ( .A(KEYINPUT12), .B(n1139), .Z(n1135) );
NOR2_X1 U817 ( .A1(n1138), .A2(n1137), .ZN(n1139) );
NOR2_X1 U818 ( .A1(n1008), .A2(n1140), .ZN(G54) );
XOR2_X1 U819 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U820 ( .A(n1143), .B(n1130), .ZN(n1142) );
XOR2_X1 U821 ( .A(G131), .B(n1089), .Z(n1130) );
NAND2_X1 U822 ( .A1(KEYINPUT48), .A2(n1144), .ZN(n1143) );
XOR2_X1 U823 ( .A(KEYINPUT56), .B(n1145), .Z(n1144) );
XOR2_X1 U824 ( .A(n1146), .B(n1147), .Z(n1141) );
NOR2_X1 U825 ( .A1(n1148), .A2(n1109), .ZN(n1147) );
INV_X1 U826 ( .A(G469), .ZN(n1148) );
NAND2_X1 U827 ( .A1(KEYINPUT37), .A2(n1149), .ZN(n1146) );
XOR2_X1 U828 ( .A(n1150), .B(n1151), .Z(n1149) );
NOR2_X1 U829 ( .A1(n1008), .A2(n1152), .ZN(G51) );
XOR2_X1 U830 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U831 ( .A(n1098), .B(n1155), .Z(n1154) );
XOR2_X1 U832 ( .A(n1156), .B(n1157), .Z(n1153) );
NOR2_X1 U833 ( .A1(n1158), .A2(KEYINPUT45), .ZN(n1157) );
NOR2_X1 U834 ( .A1(n1021), .A2(n1109), .ZN(n1158) );
NAND2_X1 U835 ( .A1(G902), .A2(n1121), .ZN(n1109) );
NAND3_X1 U836 ( .A1(n1090), .A2(n1159), .A3(n1101), .ZN(n1121) );
AND4_X1 U837 ( .A1(n1122), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1101) );
AND4_X1 U838 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
NAND4_X1 U839 ( .A1(n1167), .A2(n1015), .A3(n1168), .A4(n1169), .ZN(n1161) );
AND2_X1 U840 ( .A1(n1170), .A2(n1059), .ZN(n1168) );
XNOR2_X1 U841 ( .A(n1060), .B(KEYINPUT41), .ZN(n1167) );
OR2_X1 U842 ( .A1(n1058), .A2(n1003), .ZN(n1122) );
NAND2_X1 U843 ( .A1(n1171), .A2(n1015), .ZN(n1003) );
XNOR2_X1 U844 ( .A(KEYINPUT52), .B(n1102), .ZN(n1159) );
NAND4_X1 U845 ( .A1(n1172), .A2(n1173), .A3(n1036), .A4(n1170), .ZN(n1102) );
XOR2_X1 U846 ( .A(n1046), .B(KEYINPUT8), .Z(n1172) );
AND4_X1 U847 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1090) );
NOR4_X1 U848 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
INV_X1 U849 ( .A(n1182), .ZN(n1180) );
INV_X1 U850 ( .A(n1183), .ZN(n1179) );
NOR2_X1 U851 ( .A1(n1184), .A2(n1185), .ZN(n1176) );
NOR2_X1 U852 ( .A1(n1046), .A2(n1186), .ZN(n1185) );
INV_X1 U853 ( .A(n1187), .ZN(n1184) );
XNOR2_X1 U854 ( .A(n1188), .B(KEYINPUT34), .ZN(n1156) );
NOR2_X1 U855 ( .A1(n1071), .A2(G952), .ZN(n1008) );
XOR2_X1 U856 ( .A(G146), .B(n1189), .Z(G48) );
NOR2_X1 U857 ( .A1(KEYINPUT3), .A2(n1187), .ZN(n1189) );
NAND3_X1 U858 ( .A1(n1190), .A2(n1169), .A3(n1191), .ZN(n1187) );
XOR2_X1 U859 ( .A(n1192), .B(n1174), .Z(G45) );
NAND4_X1 U860 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1174) );
AND2_X1 U861 ( .A1(n1017), .A2(n1169), .ZN(n1195) );
XNOR2_X1 U862 ( .A(G140), .B(n1175), .ZN(G42) );
NAND2_X1 U863 ( .A1(n1197), .A2(n1198), .ZN(n1175) );
XOR2_X1 U864 ( .A(G137), .B(n1181), .Z(G39) );
AND3_X1 U865 ( .A1(n1191), .A2(n1034), .A3(n1039), .ZN(n1181) );
NAND2_X1 U866 ( .A1(n1199), .A2(n1200), .ZN(G36) );
NAND2_X1 U867 ( .A1(G134), .A2(n1182), .ZN(n1200) );
XOR2_X1 U868 ( .A(KEYINPUT0), .B(n1201), .Z(n1199) );
NOR2_X1 U869 ( .A1(G134), .A2(n1182), .ZN(n1201) );
NAND3_X1 U870 ( .A1(n1196), .A2(n1059), .A3(n1198), .ZN(n1182) );
XOR2_X1 U871 ( .A(n1202), .B(G131), .Z(G33) );
NAND2_X1 U872 ( .A1(KEYINPUT61), .A2(n1183), .ZN(n1202) );
NAND2_X1 U873 ( .A1(n1173), .A2(n1198), .ZN(n1183) );
AND2_X1 U874 ( .A1(n1039), .A2(n1194), .ZN(n1198) );
AND2_X1 U875 ( .A1(n1048), .A2(n1049), .ZN(n1039) );
XNOR2_X1 U876 ( .A(n1203), .B(KEYINPUT20), .ZN(n1048) );
XOR2_X1 U877 ( .A(n1204), .B(n1178), .Z(G30) );
AND3_X1 U878 ( .A1(n1169), .A2(n1059), .A3(n1191), .ZN(n1178) );
AND3_X1 U879 ( .A1(n1205), .A2(n1044), .A3(n1194), .ZN(n1191) );
AND2_X1 U880 ( .A1(n1060), .A2(n1206), .ZN(n1194) );
NAND2_X1 U881 ( .A1(KEYINPUT14), .A2(n1207), .ZN(n1204) );
XOR2_X1 U882 ( .A(n1138), .B(n1160), .Z(G3) );
NAND3_X1 U883 ( .A1(n1034), .A2(n1171), .A3(n1196), .ZN(n1160) );
XOR2_X1 U884 ( .A(n1083), .B(n1208), .Z(G27) );
NAND2_X1 U885 ( .A1(n1169), .A2(n1209), .ZN(n1208) );
XNOR2_X1 U886 ( .A(KEYINPUT46), .B(n1186), .ZN(n1209) );
NAND3_X1 U887 ( .A1(n1036), .A2(n1206), .A3(n1197), .ZN(n1186) );
AND3_X1 U888 ( .A1(n1043), .A2(n1044), .A3(n1190), .ZN(n1197) );
NAND2_X1 U889 ( .A1(n1210), .A2(n1061), .ZN(n1206) );
NAND4_X1 U890 ( .A1(n1211), .A2(G953), .A3(G902), .A4(n1212), .ZN(n1210) );
XNOR2_X1 U891 ( .A(G900), .B(KEYINPUT62), .ZN(n1211) );
XNOR2_X1 U892 ( .A(G122), .B(n1166), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1193), .A2(n1213), .A3(n1015), .A4(n1017), .ZN(n1166) );
NOR2_X1 U894 ( .A1(n1044), .A2(n1205), .ZN(n1015) );
XNOR2_X1 U895 ( .A(G119), .B(n1164), .ZN(G21) );
NAND4_X1 U896 ( .A1(n1213), .A2(n1034), .A3(n1205), .A4(n1044), .ZN(n1164) );
INV_X1 U897 ( .A(n1043), .ZN(n1205) );
XNOR2_X1 U898 ( .A(n1163), .B(n1214), .ZN(G18) );
NOR2_X1 U899 ( .A1(KEYINPUT31), .A2(n1215), .ZN(n1214) );
INV_X1 U900 ( .A(G116), .ZN(n1215) );
NAND3_X1 U901 ( .A1(n1213), .A2(n1059), .A3(n1196), .ZN(n1163) );
NAND2_X1 U902 ( .A1(n1216), .A2(n1217), .ZN(n1059) );
OR2_X1 U903 ( .A1(n1056), .A2(KEYINPUT6), .ZN(n1217) );
INV_X1 U904 ( .A(n1034), .ZN(n1056) );
NAND3_X1 U905 ( .A1(n1218), .A2(n1017), .A3(KEYINPUT6), .ZN(n1216) );
XOR2_X1 U906 ( .A(G113), .B(n1219), .Z(G15) );
AND2_X1 U907 ( .A1(n1213), .A2(n1173), .ZN(n1219) );
NOR2_X1 U908 ( .A1(n1058), .A2(n1041), .ZN(n1173) );
INV_X1 U909 ( .A(n1196), .ZN(n1041) );
NOR2_X1 U910 ( .A1(n1044), .A2(n1043), .ZN(n1196) );
INV_X1 U911 ( .A(n1190), .ZN(n1058) );
NOR2_X1 U912 ( .A1(n1218), .A2(n1017), .ZN(n1190) );
INV_X1 U913 ( .A(n1193), .ZN(n1218) );
AND3_X1 U914 ( .A1(n1169), .A2(n1170), .A3(n1036), .ZN(n1213) );
AND2_X1 U915 ( .A1(n1055), .A2(n1057), .ZN(n1036) );
NAND2_X1 U916 ( .A1(n1220), .A2(n1221), .ZN(G12) );
NAND2_X1 U917 ( .A1(G110), .A2(n1165), .ZN(n1221) );
XOR2_X1 U918 ( .A(n1222), .B(KEYINPUT49), .Z(n1220) );
OR2_X1 U919 ( .A1(n1165), .A2(G110), .ZN(n1222) );
NAND4_X1 U920 ( .A1(n1034), .A2(n1171), .A3(n1043), .A4(n1044), .ZN(n1165) );
NAND3_X1 U921 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1044) );
NAND2_X1 U922 ( .A1(n1226), .A2(n1107), .ZN(n1225) );
OR3_X1 U923 ( .A1(n1107), .A2(n1226), .A3(G902), .ZN(n1224) );
NOR2_X1 U924 ( .A1(n1108), .A2(G234), .ZN(n1226) );
INV_X1 U925 ( .A(G217), .ZN(n1108) );
XNOR2_X1 U926 ( .A(n1227), .B(n1228), .ZN(n1107) );
XOR2_X1 U927 ( .A(G125), .B(n1229), .Z(n1228) );
XOR2_X1 U928 ( .A(G146), .B(G128), .Z(n1229) );
XOR2_X1 U929 ( .A(n1230), .B(n1231), .Z(n1227) );
XNOR2_X1 U930 ( .A(n1232), .B(n1233), .ZN(n1230) );
NOR2_X1 U931 ( .A1(G119), .A2(KEYINPUT28), .ZN(n1233) );
NOR3_X1 U932 ( .A1(n1234), .A2(KEYINPUT63), .A3(n1235), .ZN(n1232) );
NOR4_X1 U933 ( .A1(G953), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1235) );
XNOR2_X1 U934 ( .A(G137), .B(KEYINPUT53), .ZN(n1236) );
NOR2_X1 U935 ( .A1(n1239), .A2(G137), .ZN(n1234) );
NOR3_X1 U936 ( .A1(n1238), .A2(G953), .A3(n1237), .ZN(n1239) );
INV_X1 U937 ( .A(G234), .ZN(n1237) );
INV_X1 U938 ( .A(G221), .ZN(n1238) );
NAND2_X1 U939 ( .A1(G217), .A2(G902), .ZN(n1223) );
XOR2_X1 U940 ( .A(n1240), .B(G472), .Z(n1043) );
NAND2_X1 U941 ( .A1(n1241), .A2(n1242), .ZN(n1240) );
XOR2_X1 U942 ( .A(n1243), .B(n1244), .Z(n1241) );
XOR2_X1 U943 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U944 ( .A(n1247), .B(n1129), .Z(n1246) );
NAND2_X1 U945 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND2_X1 U946 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NAND2_X1 U947 ( .A1(KEYINPUT17), .A2(n1252), .ZN(n1251) );
NAND2_X1 U948 ( .A1(KEYINPUT21), .A2(n1138), .ZN(n1252) );
INV_X1 U949 ( .A(n1137), .ZN(n1250) );
NAND2_X1 U950 ( .A1(G101), .A2(n1253), .ZN(n1248) );
NAND2_X1 U951 ( .A1(KEYINPUT21), .A2(n1254), .ZN(n1253) );
NAND2_X1 U952 ( .A1(KEYINPUT17), .A2(n1137), .ZN(n1254) );
NAND3_X1 U953 ( .A1(n1255), .A2(n1071), .A3(G210), .ZN(n1137) );
XNOR2_X1 U954 ( .A(n1256), .B(n1257), .ZN(n1243) );
XNOR2_X1 U955 ( .A(KEYINPUT57), .B(KEYINPUT16), .ZN(n1256) );
AND3_X1 U956 ( .A1(n1169), .A2(n1170), .A3(n1060), .ZN(n1171) );
NOR2_X1 U957 ( .A1(n1055), .A2(n1258), .ZN(n1060) );
XOR2_X1 U958 ( .A(KEYINPUT18), .B(n1057), .Z(n1258) );
NAND2_X1 U959 ( .A1(G221), .A2(n1259), .ZN(n1057) );
NAND2_X1 U960 ( .A1(G234), .A2(n1242), .ZN(n1259) );
XNOR2_X1 U961 ( .A(n1016), .B(n1260), .ZN(n1055) );
XOR2_X1 U962 ( .A(KEYINPUT42), .B(G469), .Z(n1260) );
NAND2_X1 U963 ( .A1(n1261), .A2(n1242), .ZN(n1016) );
XOR2_X1 U964 ( .A(n1262), .B(n1145), .Z(n1261) );
XNOR2_X1 U965 ( .A(n1263), .B(n1231), .ZN(n1145) );
XNOR2_X1 U966 ( .A(G110), .B(n1084), .ZN(n1231) );
NAND2_X1 U967 ( .A1(G227), .A2(n1071), .ZN(n1263) );
NOR2_X1 U968 ( .A1(KEYINPUT27), .A2(n1264), .ZN(n1262) );
XNOR2_X1 U969 ( .A(n1265), .B(n1151), .ZN(n1264) );
XOR2_X1 U970 ( .A(n1266), .B(n1086), .Z(n1151) );
XOR2_X1 U971 ( .A(n1267), .B(n1207), .Z(n1086) );
XNOR2_X1 U972 ( .A(KEYINPUT26), .B(KEYINPUT22), .ZN(n1267) );
XOR2_X1 U973 ( .A(n1268), .B(n1269), .Z(n1266) );
NAND2_X1 U974 ( .A1(KEYINPUT13), .A2(n1270), .ZN(n1268) );
XNOR2_X1 U975 ( .A(n1245), .B(KEYINPUT9), .ZN(n1265) );
XOR2_X1 U976 ( .A(n1088), .B(n1089), .Z(n1245) );
XOR2_X1 U977 ( .A(G134), .B(G137), .Z(n1089) );
NAND2_X1 U978 ( .A1(n1271), .A2(n1061), .ZN(n1170) );
NAND3_X1 U979 ( .A1(n1212), .A2(n1071), .A3(G952), .ZN(n1061) );
XOR2_X1 U980 ( .A(KEYINPUT2), .B(n1272), .Z(n1271) );
AND4_X1 U981 ( .A1(n1097), .A2(n1212), .A3(G902), .A4(G953), .ZN(n1272) );
NAND2_X1 U982 ( .A1(G237), .A2(G234), .ZN(n1212) );
INV_X1 U983 ( .A(G898), .ZN(n1097) );
INV_X1 U984 ( .A(n1046), .ZN(n1169) );
NAND2_X1 U985 ( .A1(n1273), .A2(n1049), .ZN(n1046) );
NAND2_X1 U986 ( .A1(G214), .A2(n1274), .ZN(n1049) );
XOR2_X1 U987 ( .A(n1203), .B(KEYINPUT23), .Z(n1273) );
XOR2_X1 U988 ( .A(n1021), .B(n1275), .Z(n1203) );
NOR2_X1 U989 ( .A1(KEYINPUT29), .A2(n1022), .ZN(n1275) );
NAND2_X1 U990 ( .A1(n1276), .A2(n1242), .ZN(n1022) );
XNOR2_X1 U991 ( .A(n1277), .B(n1098), .ZN(n1276) );
XNOR2_X1 U992 ( .A(n1278), .B(n1279), .ZN(n1098) );
XOR2_X1 U993 ( .A(n1280), .B(n1129), .Z(n1279) );
XOR2_X1 U994 ( .A(n1281), .B(n1282), .Z(n1129) );
XOR2_X1 U995 ( .A(G119), .B(G116), .Z(n1282) );
INV_X1 U996 ( .A(G113), .ZN(n1281) );
NAND2_X1 U997 ( .A1(n1283), .A2(n1284), .ZN(n1280) );
NAND2_X1 U998 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XNOR2_X1 U999 ( .A(KEYINPUT11), .B(n1270), .ZN(n1286) );
XNOR2_X1 U1000 ( .A(n1269), .B(KEYINPUT33), .ZN(n1285) );
XOR2_X1 U1001 ( .A(KEYINPUT39), .B(n1287), .Z(n1283) );
AND2_X1 U1002 ( .A1(n1269), .A2(n1270), .ZN(n1287) );
XNOR2_X1 U1003 ( .A(G104), .B(G107), .ZN(n1270) );
XNOR2_X1 U1004 ( .A(n1138), .B(KEYINPUT59), .ZN(n1269) );
INV_X1 U1005 ( .A(G101), .ZN(n1138) );
XNOR2_X1 U1006 ( .A(G110), .B(n1288), .ZN(n1278) );
NOR2_X1 U1007 ( .A1(G122), .A2(KEYINPUT25), .ZN(n1288) );
NAND2_X1 U1008 ( .A1(n1289), .A2(n1290), .ZN(n1277) );
OR2_X1 U1009 ( .A1(n1155), .A2(n1188), .ZN(n1290) );
XOR2_X1 U1010 ( .A(n1291), .B(KEYINPUT43), .Z(n1289) );
NAND2_X1 U1011 ( .A1(n1188), .A2(n1155), .ZN(n1291) );
XOR2_X1 U1012 ( .A(n1126), .B(G125), .Z(n1155) );
XOR2_X1 U1013 ( .A(n1257), .B(n1150), .Z(n1126) );
NAND2_X1 U1014 ( .A1(KEYINPUT38), .A2(n1207), .ZN(n1257) );
NOR2_X1 U1015 ( .A1(n1104), .A2(G953), .ZN(n1188) );
INV_X1 U1016 ( .A(G224), .ZN(n1104) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1274), .ZN(n1021) );
NAND2_X1 U1018 ( .A1(n1292), .A2(n1242), .ZN(n1274) );
INV_X1 U1019 ( .A(G237), .ZN(n1292) );
NOR2_X1 U1020 ( .A1(n1017), .A2(n1193), .ZN(n1034) );
XOR2_X1 U1021 ( .A(n1293), .B(n1115), .Z(n1193) );
INV_X1 U1022 ( .A(n1024), .ZN(n1115) );
NAND2_X1 U1023 ( .A1(n1118), .A2(n1242), .ZN(n1024) );
XOR2_X1 U1024 ( .A(n1294), .B(n1295), .Z(n1118) );
XNOR2_X1 U1025 ( .A(n1088), .B(n1296), .ZN(n1295) );
XOR2_X1 U1026 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U1027 ( .A1(G122), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1028 ( .A(KEYINPUT51), .B(KEYINPUT50), .Z(n1299) );
NAND2_X1 U1029 ( .A1(n1300), .A2(n1301), .ZN(n1297) );
NAND2_X1 U1030 ( .A1(n1084), .A2(n1302), .ZN(n1301) );
NAND2_X1 U1031 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U1032 ( .A1(n1083), .A2(n1305), .ZN(n1304) );
INV_X1 U1033 ( .A(G125), .ZN(n1083) );
INV_X1 U1034 ( .A(KEYINPUT30), .ZN(n1303) );
NAND2_X1 U1035 ( .A1(G125), .A2(n1306), .ZN(n1300) );
NAND2_X1 U1036 ( .A1(n1305), .A2(n1307), .ZN(n1306) );
OR2_X1 U1037 ( .A1(n1084), .A2(KEYINPUT30), .ZN(n1307) );
XNOR2_X1 U1038 ( .A(G140), .B(KEYINPUT4), .ZN(n1084) );
INV_X1 U1039 ( .A(KEYINPUT35), .ZN(n1305) );
XOR2_X1 U1040 ( .A(G131), .B(n1308), .Z(n1088) );
INV_X1 U1041 ( .A(n1150), .ZN(n1308) );
XOR2_X1 U1042 ( .A(n1192), .B(G146), .Z(n1150) );
INV_X1 U1043 ( .A(G143), .ZN(n1192) );
XOR2_X1 U1044 ( .A(n1309), .B(n1310), .Z(n1294) );
XOR2_X1 U1045 ( .A(G113), .B(G104), .Z(n1310) );
NAND3_X1 U1046 ( .A1(n1255), .A2(n1071), .A3(G214), .ZN(n1309) );
XOR2_X1 U1047 ( .A(G237), .B(KEYINPUT54), .Z(n1255) );
NAND2_X1 U1048 ( .A1(KEYINPUT15), .A2(n1023), .ZN(n1293) );
INV_X1 U1049 ( .A(G475), .ZN(n1023) );
XNOR2_X1 U1050 ( .A(n1311), .B(G478), .ZN(n1017) );
NAND2_X1 U1051 ( .A1(n1312), .A2(n1242), .ZN(n1311) );
INV_X1 U1052 ( .A(G902), .ZN(n1242) );
XOR2_X1 U1053 ( .A(KEYINPUT47), .B(n1112), .Z(n1312) );
XNOR2_X1 U1054 ( .A(n1313), .B(n1314), .ZN(n1112) );
XOR2_X1 U1055 ( .A(n1315), .B(n1316), .Z(n1314) );
XOR2_X1 U1056 ( .A(G143), .B(G134), .Z(n1316) );
XOR2_X1 U1057 ( .A(KEYINPUT5), .B(KEYINPUT19), .Z(n1315) );
XOR2_X1 U1058 ( .A(n1317), .B(n1318), .Z(n1313) );
XOR2_X1 U1059 ( .A(n1319), .B(n1320), .Z(n1318) );
NAND3_X1 U1060 ( .A1(n1321), .A2(n1071), .A3(G217), .ZN(n1320) );
INV_X1 U1061 ( .A(G953), .ZN(n1071) );
XOR2_X1 U1062 ( .A(KEYINPUT1), .B(G234), .Z(n1321) );
NAND2_X1 U1063 ( .A1(KEYINPUT36), .A2(n1322), .ZN(n1319) );
XOR2_X1 U1064 ( .A(G122), .B(G116), .Z(n1322) );
XOR2_X1 U1065 ( .A(G107), .B(n1207), .Z(n1317) );
INV_X1 U1066 ( .A(G128), .ZN(n1207) );
endmodule


