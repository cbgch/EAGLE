//Key = 1110100101110010001111110111101100000111111100000001000011111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327;

XNOR2_X1 U723 ( .A(G107), .B(n1014), .ZN(G9) );
NOR2_X1 U724 ( .A1(n1015), .A2(n1016), .ZN(G75) );
NOR3_X1 U725 ( .A1(n1017), .A2(n1018), .A3(n1019), .ZN(n1016) );
NOR3_X1 U726 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1018) );
NOR3_X1 U727 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1021) );
NOR2_X1 U728 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U729 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
AND2_X1 U730 ( .A1(n1030), .A2(KEYINPUT21), .ZN(n1028) );
NOR4_X1 U731 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1024) );
NOR2_X1 U732 ( .A1(n1035), .A2(n1036), .ZN(n1031) );
NOR2_X1 U733 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NOR2_X1 U734 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U735 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR2_X1 U736 ( .A1(n1043), .A2(n1044), .ZN(n1035) );
NOR2_X1 U737 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NOR2_X1 U738 ( .A1(n1047), .A2(KEYINPUT21), .ZN(n1023) );
NOR2_X1 U739 ( .A1(n1048), .A2(n1027), .ZN(n1047) );
INV_X1 U740 ( .A(n1049), .ZN(n1027) );
NAND3_X1 U741 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1017) );
NAND4_X1 U742 ( .A1(n1053), .A2(n1049), .A3(n1054), .A4(n1055), .ZN(n1052) );
NAND3_X1 U743 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
INV_X1 U744 ( .A(n1059), .ZN(n1058) );
NAND2_X1 U745 ( .A1(KEYINPUT45), .A2(n1060), .ZN(n1057) );
OR3_X1 U746 ( .A1(n1020), .A2(KEYINPUT45), .A3(n1060), .ZN(n1056) );
NOR3_X1 U747 ( .A1(n1044), .A2(n1038), .A3(n1033), .ZN(n1049) );
AND3_X1 U748 ( .A1(n1050), .A2(n1051), .A3(n1061), .ZN(n1015) );
NAND4_X1 U749 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1050) );
NOR4_X1 U750 ( .A1(n1066), .A2(n1067), .A3(n1020), .A4(n1068), .ZN(n1065) );
XNOR2_X1 U751 ( .A(G478), .B(n1069), .ZN(n1068) );
NAND2_X1 U752 ( .A1(KEYINPUT60), .A2(n1070), .ZN(n1069) );
NOR2_X1 U753 ( .A1(n1071), .A2(n1022), .ZN(n1064) );
XNOR2_X1 U754 ( .A(n1072), .B(n1073), .ZN(n1063) );
NAND2_X1 U755 ( .A1(KEYINPUT9), .A2(n1074), .ZN(n1073) );
XOR2_X1 U756 ( .A(G469), .B(n1075), .Z(n1062) );
NOR2_X1 U757 ( .A1(n1076), .A2(KEYINPUT32), .ZN(n1075) );
XOR2_X1 U758 ( .A(n1077), .B(n1078), .Z(G72) );
NOR2_X1 U759 ( .A1(n1079), .A2(n1051), .ZN(n1078) );
AND2_X1 U760 ( .A1(G227), .A2(G900), .ZN(n1079) );
NAND3_X1 U761 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1077) );
NAND2_X1 U762 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
OR3_X1 U763 ( .A1(n1084), .A2(n1083), .A3(n1085), .ZN(n1081) );
OR2_X1 U764 ( .A1(G953), .A2(n1086), .ZN(n1083) );
INV_X1 U765 ( .A(KEYINPUT23), .ZN(n1084) );
NAND3_X1 U766 ( .A1(n1086), .A2(n1087), .A3(n1085), .ZN(n1080) );
XNOR2_X1 U767 ( .A(n1088), .B(n1089), .ZN(n1085) );
XOR2_X1 U768 ( .A(n1090), .B(n1091), .Z(n1089) );
XNOR2_X1 U769 ( .A(G125), .B(G131), .ZN(n1091) );
NAND2_X1 U770 ( .A1(KEYINPUT38), .A2(G140), .ZN(n1090) );
XOR2_X1 U771 ( .A(n1092), .B(n1093), .Z(n1088) );
NAND2_X1 U772 ( .A1(G953), .A2(n1094), .ZN(n1087) );
XOR2_X1 U773 ( .A(n1095), .B(n1096), .Z(G69) );
XOR2_X1 U774 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U775 ( .A1(n1099), .A2(G953), .ZN(n1098) );
NOR2_X1 U776 ( .A1(n1100), .A2(n1101), .ZN(n1097) );
XNOR2_X1 U777 ( .A(G953), .B(KEYINPUT44), .ZN(n1101) );
AND2_X1 U778 ( .A1(G224), .A2(G898), .ZN(n1100) );
NOR2_X1 U779 ( .A1(n1102), .A2(n1103), .ZN(n1095) );
NOR2_X1 U780 ( .A1(KEYINPUT46), .A2(n1104), .ZN(n1103) );
INV_X1 U781 ( .A(n1105), .ZN(n1104) );
NOR2_X1 U782 ( .A1(KEYINPUT2), .A2(n1105), .ZN(n1102) );
NAND2_X1 U783 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U784 ( .A1(G953), .A2(n1108), .ZN(n1107) );
XOR2_X1 U785 ( .A(n1109), .B(n1110), .Z(n1106) );
XOR2_X1 U786 ( .A(KEYINPUT33), .B(n1111), .Z(n1110) );
NOR2_X1 U787 ( .A1(n1112), .A2(n1113), .ZN(G66) );
NOR3_X1 U788 ( .A1(n1072), .A2(n1114), .A3(n1115), .ZN(n1113) );
NOR2_X1 U789 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
AND3_X1 U790 ( .A1(n1117), .A2(G902), .A3(n1116), .ZN(n1114) );
NOR3_X1 U791 ( .A1(KEYINPUT16), .A2(n1118), .A3(n1119), .ZN(n1116) );
INV_X1 U792 ( .A(n1019), .ZN(n1118) );
NOR2_X1 U793 ( .A1(n1112), .A2(n1120), .ZN(G63) );
NOR3_X1 U794 ( .A1(n1070), .A2(n1121), .A3(n1122), .ZN(n1120) );
AND2_X1 U795 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR3_X1 U796 ( .A1(n1124), .A2(n1125), .A3(n1123), .ZN(n1121) );
NAND3_X1 U797 ( .A1(G478), .A2(n1019), .A3(KEYINPUT0), .ZN(n1123) );
NOR2_X1 U798 ( .A1(n1112), .A2(n1126), .ZN(G60) );
XOR2_X1 U799 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND4_X1 U800 ( .A1(KEYINPUT56), .A2(G475), .A3(n1129), .A4(n1019), .ZN(n1128) );
XNOR2_X1 U801 ( .A(KEYINPUT63), .B(n1125), .ZN(n1129) );
NAND2_X1 U802 ( .A1(n1130), .A2(n1131), .ZN(G6) );
NAND3_X1 U803 ( .A1(KEYINPUT4), .A2(n1132), .A3(n1133), .ZN(n1131) );
NAND2_X1 U804 ( .A1(n1134), .A2(G104), .ZN(n1130) );
NAND2_X1 U805 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U806 ( .A1(n1137), .A2(n1132), .ZN(n1136) );
NAND2_X1 U807 ( .A1(n1138), .A2(n1139), .ZN(n1135) );
NAND2_X1 U808 ( .A1(KEYINPUT4), .A2(n1132), .ZN(n1139) );
INV_X1 U809 ( .A(n1137), .ZN(n1138) );
XOR2_X1 U810 ( .A(KEYINPUT57), .B(KEYINPUT43), .Z(n1137) );
NOR2_X1 U811 ( .A1(n1112), .A2(n1140), .ZN(G57) );
XOR2_X1 U812 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U814 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U815 ( .A1(n1147), .A2(KEYINPUT13), .ZN(n1145) );
XOR2_X1 U816 ( .A(n1148), .B(n1149), .Z(n1141) );
XOR2_X1 U817 ( .A(KEYINPUT47), .B(KEYINPUT22), .Z(n1149) );
NAND3_X1 U818 ( .A1(G902), .A2(n1150), .A3(G472), .ZN(n1148) );
XNOR2_X1 U819 ( .A(KEYINPUT30), .B(n1019), .ZN(n1150) );
NOR3_X1 U820 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(G54) );
NOR3_X1 U821 ( .A1(n1154), .A2(n1051), .A3(n1061), .ZN(n1153) );
INV_X1 U822 ( .A(G952), .ZN(n1061) );
AND2_X1 U823 ( .A1(n1154), .A2(n1112), .ZN(n1152) );
INV_X1 U824 ( .A(KEYINPUT53), .ZN(n1154) );
XOR2_X1 U825 ( .A(n1155), .B(n1156), .Z(n1151) );
XNOR2_X1 U826 ( .A(n1157), .B(n1158), .ZN(n1156) );
NAND2_X1 U827 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U828 ( .A1(G140), .A2(n1161), .ZN(n1160) );
INV_X1 U829 ( .A(n1162), .ZN(n1159) );
XOR2_X1 U830 ( .A(n1163), .B(n1164), .Z(n1155) );
XNOR2_X1 U831 ( .A(n1147), .B(n1165), .ZN(n1164) );
INV_X1 U832 ( .A(n1166), .ZN(n1147) );
NAND4_X1 U833 ( .A1(KEYINPUT14), .A2(G902), .A3(G469), .A4(n1019), .ZN(n1163) );
NOR2_X1 U834 ( .A1(n1112), .A2(n1167), .ZN(G51) );
NOR2_X1 U835 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U836 ( .A(n1170), .B(KEYINPUT11), .Z(n1169) );
NAND2_X1 U837 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
XNOR2_X1 U839 ( .A(n1173), .B(KEYINPUT59), .ZN(n1172) );
AND3_X1 U840 ( .A1(n1174), .A2(n1019), .A3(G902), .ZN(n1171) );
NAND2_X1 U841 ( .A1(n1099), .A2(n1086), .ZN(n1019) );
AND4_X1 U842 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1086) );
NOR4_X1 U843 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1178) );
NOR3_X1 U844 ( .A1(n1183), .A2(n1184), .A3(n1185), .ZN(n1177) );
NOR2_X1 U845 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
INV_X1 U846 ( .A(KEYINPUT10), .ZN(n1186) );
NOR4_X1 U847 ( .A1(KEYINPUT10), .A2(n1188), .A3(n1029), .A4(n1189), .ZN(n1184) );
AND4_X1 U848 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1099) );
AND4_X1 U849 ( .A1(n1014), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1193) );
NAND3_X1 U850 ( .A1(n1045), .A2(n1197), .A3(n1040), .ZN(n1014) );
NOR2_X1 U851 ( .A1(n1132), .A2(n1198), .ZN(n1192) );
NOR2_X1 U852 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
AND3_X1 U853 ( .A1(n1040), .A2(n1197), .A3(n1046), .ZN(n1132) );
NOR2_X1 U854 ( .A1(n1051), .A2(G952), .ZN(n1112) );
XNOR2_X1 U855 ( .A(n1183), .B(n1201), .ZN(G48) );
NAND2_X1 U856 ( .A1(KEYINPUT1), .A2(G146), .ZN(n1201) );
AND4_X1 U857 ( .A1(n1202), .A2(n1046), .A3(n1032), .A4(n1034), .ZN(n1183) );
NAND2_X1 U858 ( .A1(n1203), .A2(n1204), .ZN(G45) );
OR2_X1 U859 ( .A1(n1205), .A2(G143), .ZN(n1204) );
NAND2_X1 U860 ( .A1(G143), .A2(n1206), .ZN(n1203) );
NAND2_X1 U861 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
OR2_X1 U862 ( .A1(n1176), .A2(KEYINPUT61), .ZN(n1208) );
NAND2_X1 U863 ( .A1(KEYINPUT61), .A2(n1205), .ZN(n1207) );
NAND2_X1 U864 ( .A1(n1209), .A2(n1210), .ZN(n1205) );
INV_X1 U865 ( .A(n1176), .ZN(n1210) );
NAND4_X1 U866 ( .A1(n1202), .A2(n1029), .A3(n1211), .A4(n1067), .ZN(n1176) );
XNOR2_X1 U867 ( .A(KEYINPUT25), .B(KEYINPUT19), .ZN(n1209) );
XOR2_X1 U868 ( .A(G140), .B(n1182), .Z(G42) );
NOR3_X1 U869 ( .A1(n1189), .A2(n1048), .A3(n1188), .ZN(n1182) );
INV_X1 U870 ( .A(n1030), .ZN(n1048) );
XNOR2_X1 U871 ( .A(G137), .B(n1175), .ZN(G39) );
NAND2_X1 U872 ( .A1(n1212), .A2(n1213), .ZN(n1175) );
XNOR2_X1 U873 ( .A(n1214), .B(n1181), .ZN(G36) );
AND3_X1 U874 ( .A1(n1029), .A2(n1045), .A3(n1212), .ZN(n1181) );
XOR2_X1 U875 ( .A(n1187), .B(n1215), .Z(G33) );
NAND2_X1 U876 ( .A1(KEYINPUT18), .A2(G131), .ZN(n1215) );
NAND3_X1 U877 ( .A1(n1029), .A2(n1046), .A3(n1212), .ZN(n1187) );
INV_X1 U878 ( .A(n1188), .ZN(n1212) );
NAND4_X1 U879 ( .A1(n1216), .A2(n1040), .A3(n1217), .A4(n1060), .ZN(n1188) );
XNOR2_X1 U880 ( .A(n1180), .B(n1218), .ZN(G30) );
NAND2_X1 U881 ( .A1(G128), .A2(n1219), .ZN(n1218) );
XOR2_X1 U882 ( .A(KEYINPUT48), .B(KEYINPUT42), .Z(n1219) );
AND4_X1 U883 ( .A1(n1202), .A2(n1045), .A3(n1032), .A4(n1034), .ZN(n1180) );
AND3_X1 U884 ( .A1(n1059), .A2(n1217), .A3(n1040), .ZN(n1202) );
INV_X1 U885 ( .A(n1220), .ZN(n1040) );
XOR2_X1 U886 ( .A(n1190), .B(n1221), .Z(G3) );
NOR2_X1 U887 ( .A1(G101), .A2(KEYINPUT6), .ZN(n1221) );
NAND2_X1 U888 ( .A1(n1029), .A2(n1222), .ZN(n1190) );
XOR2_X1 U889 ( .A(n1179), .B(n1223), .Z(G27) );
NOR2_X1 U890 ( .A1(KEYINPUT15), .A2(n1224), .ZN(n1223) );
AND4_X1 U891 ( .A1(n1059), .A2(n1217), .A3(n1030), .A4(n1225), .ZN(n1179) );
NOR2_X1 U892 ( .A1(n1189), .A2(n1044), .ZN(n1225) );
INV_X1 U893 ( .A(n1226), .ZN(n1044) );
NAND2_X1 U894 ( .A1(n1033), .A2(n1227), .ZN(n1217) );
NAND4_X1 U895 ( .A1(G953), .A2(G902), .A3(n1228), .A4(n1094), .ZN(n1227) );
INV_X1 U896 ( .A(G900), .ZN(n1094) );
NAND3_X1 U897 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(G24) );
NAND2_X1 U898 ( .A1(KEYINPUT49), .A2(G122), .ZN(n1231) );
OR3_X1 U899 ( .A1(G122), .A2(KEYINPUT49), .A3(n1191), .ZN(n1230) );
NAND2_X1 U900 ( .A1(n1232), .A2(n1191), .ZN(n1229) );
NAND4_X1 U901 ( .A1(n1226), .A2(n1197), .A3(n1211), .A4(n1067), .ZN(n1191) );
NOR3_X1 U902 ( .A1(n1034), .A2(n1032), .A3(n1199), .ZN(n1197) );
NAND2_X1 U903 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
INV_X1 U904 ( .A(KEYINPUT49), .ZN(n1234) );
XOR2_X1 U905 ( .A(KEYINPUT26), .B(G122), .Z(n1233) );
XNOR2_X1 U906 ( .A(G119), .B(n1196), .ZN(G21) );
NAND3_X1 U907 ( .A1(n1226), .A2(n1235), .A3(n1213), .ZN(n1196) );
NOR3_X1 U908 ( .A1(n1054), .A2(n1053), .A3(n1038), .ZN(n1213) );
XNOR2_X1 U909 ( .A(n1236), .B(n1237), .ZN(G18) );
NOR3_X1 U910 ( .A1(n1200), .A2(KEYINPUT3), .A3(n1199), .ZN(n1237) );
NAND3_X1 U911 ( .A1(n1226), .A2(n1045), .A3(n1029), .ZN(n1200) );
AND2_X1 U912 ( .A1(n1238), .A2(n1211), .ZN(n1045) );
XNOR2_X1 U913 ( .A(n1239), .B(KEYINPUT8), .ZN(n1211) );
XNOR2_X1 U914 ( .A(G113), .B(n1195), .ZN(G15) );
NAND4_X1 U915 ( .A1(n1029), .A2(n1226), .A3(n1046), .A4(n1235), .ZN(n1195) );
INV_X1 U916 ( .A(n1199), .ZN(n1235) );
INV_X1 U917 ( .A(n1189), .ZN(n1046) );
NAND2_X1 U918 ( .A1(n1067), .A2(n1239), .ZN(n1189) );
NOR2_X1 U919 ( .A1(n1042), .A2(n1071), .ZN(n1226) );
NOR2_X1 U920 ( .A1(n1034), .A2(n1054), .ZN(n1029) );
INV_X1 U921 ( .A(n1032), .ZN(n1054) );
XNOR2_X1 U922 ( .A(G110), .B(n1194), .ZN(G12) );
NAND2_X1 U923 ( .A1(n1030), .A2(n1222), .ZN(n1194) );
NOR3_X1 U924 ( .A1(n1220), .A2(n1199), .A3(n1038), .ZN(n1222) );
NAND2_X1 U925 ( .A1(n1238), .A2(n1239), .ZN(n1038) );
NAND3_X1 U926 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1239) );
NAND2_X1 U927 ( .A1(n1070), .A2(n1243), .ZN(n1242) );
INV_X1 U928 ( .A(KEYINPUT27), .ZN(n1243) );
NAND3_X1 U929 ( .A1(KEYINPUT27), .A2(n1244), .A3(n1245), .ZN(n1241) );
OR2_X1 U930 ( .A1(n1245), .A2(n1244), .ZN(n1240) );
NOR2_X1 U931 ( .A1(n1070), .A2(KEYINPUT17), .ZN(n1244) );
AND2_X1 U932 ( .A1(n1124), .A2(n1125), .ZN(n1070) );
XNOR2_X1 U933 ( .A(n1246), .B(n1247), .ZN(n1124) );
XNOR2_X1 U934 ( .A(n1248), .B(n1249), .ZN(n1247) );
XOR2_X1 U935 ( .A(n1250), .B(n1251), .Z(n1246) );
XNOR2_X1 U936 ( .A(n1214), .B(G107), .ZN(n1251) );
INV_X1 U937 ( .A(G134), .ZN(n1214) );
OR2_X1 U938 ( .A1(n1119), .A2(n1252), .ZN(n1250) );
INV_X1 U939 ( .A(G217), .ZN(n1119) );
INV_X1 U940 ( .A(G478), .ZN(n1245) );
INV_X1 U941 ( .A(n1067), .ZN(n1238) );
XOR2_X1 U942 ( .A(G475), .B(n1253), .Z(n1067) );
AND2_X1 U943 ( .A1(n1127), .A2(n1125), .ZN(n1253) );
NAND2_X1 U944 ( .A1(n1254), .A2(n1255), .ZN(n1127) );
NAND2_X1 U945 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U946 ( .A(KEYINPUT7), .B(n1258), .Z(n1254) );
NOR2_X1 U947 ( .A1(n1257), .A2(n1256), .ZN(n1258) );
XNOR2_X1 U948 ( .A(n1133), .B(n1259), .ZN(n1256) );
NOR2_X1 U949 ( .A1(KEYINPUT12), .A2(n1260), .ZN(n1259) );
NOR2_X1 U950 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U951 ( .A(KEYINPUT52), .B(n1263), .Z(n1262) );
AND2_X1 U952 ( .A1(n1264), .A2(G122), .ZN(n1263) );
NOR2_X1 U953 ( .A1(G122), .A2(n1264), .ZN(n1261) );
XNOR2_X1 U954 ( .A(n1265), .B(n1266), .ZN(n1257) );
XOR2_X1 U955 ( .A(G143), .B(G131), .Z(n1266) );
XOR2_X1 U956 ( .A(n1267), .B(n1268), .Z(n1265) );
AND3_X1 U957 ( .A1(G214), .A2(n1051), .A3(n1269), .ZN(n1268) );
NAND2_X1 U958 ( .A1(KEYINPUT39), .A2(n1270), .ZN(n1267) );
NAND2_X1 U959 ( .A1(n1059), .A2(n1271), .ZN(n1199) );
NAND2_X1 U960 ( .A1(n1033), .A2(n1272), .ZN(n1271) );
NAND4_X1 U961 ( .A1(G953), .A2(G902), .A3(n1228), .A4(n1108), .ZN(n1272) );
INV_X1 U962 ( .A(G898), .ZN(n1108) );
NAND3_X1 U963 ( .A1(n1228), .A2(n1051), .A3(G952), .ZN(n1033) );
NAND2_X1 U964 ( .A1(G237), .A2(G234), .ZN(n1228) );
NOR2_X1 U965 ( .A1(n1216), .A2(n1022), .ZN(n1059) );
INV_X1 U966 ( .A(n1060), .ZN(n1022) );
NAND2_X1 U967 ( .A1(G214), .A2(n1273), .ZN(n1060) );
INV_X1 U968 ( .A(n1020), .ZN(n1216) );
XNOR2_X1 U969 ( .A(n1274), .B(n1174), .ZN(n1020) );
AND2_X1 U970 ( .A1(G210), .A2(n1273), .ZN(n1174) );
NAND2_X1 U971 ( .A1(n1269), .A2(n1125), .ZN(n1273) );
NAND2_X1 U972 ( .A1(n1275), .A2(n1125), .ZN(n1274) );
XNOR2_X1 U973 ( .A(n1276), .B(n1173), .ZN(n1275) );
XOR2_X1 U974 ( .A(n1277), .B(n1278), .Z(n1173) );
XNOR2_X1 U975 ( .A(n1279), .B(n1109), .ZN(n1278) );
XOR2_X1 U976 ( .A(n1280), .B(n1249), .Z(n1109) );
XNOR2_X1 U977 ( .A(n1236), .B(G122), .ZN(n1249) );
XNOR2_X1 U978 ( .A(n1281), .B(n1161), .ZN(n1280) );
NAND2_X1 U979 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U980 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U981 ( .A(n1286), .B(KEYINPUT24), .Z(n1282) );
OR2_X1 U982 ( .A1(n1284), .A2(n1285), .ZN(n1286) );
INV_X1 U983 ( .A(G101), .ZN(n1285) );
NAND2_X1 U984 ( .A1(n1287), .A2(n1288), .ZN(n1284) );
OR2_X1 U985 ( .A1(n1289), .A2(KEYINPUT54), .ZN(n1288) );
NAND3_X1 U986 ( .A1(G104), .A2(n1290), .A3(KEYINPUT54), .ZN(n1287) );
INV_X1 U987 ( .A(G107), .ZN(n1290) );
XOR2_X1 U988 ( .A(n1291), .B(n1292), .Z(n1277) );
XNOR2_X1 U989 ( .A(KEYINPUT58), .B(n1224), .ZN(n1292) );
INV_X1 U990 ( .A(G125), .ZN(n1224) );
NAND2_X1 U991 ( .A1(G224), .A2(n1051), .ZN(n1291) );
XNOR2_X1 U992 ( .A(KEYINPUT35), .B(KEYINPUT28), .ZN(n1276) );
NAND2_X1 U993 ( .A1(n1293), .A2(n1042), .ZN(n1220) );
XOR2_X1 U994 ( .A(n1076), .B(G469), .Z(n1042) );
AND2_X1 U995 ( .A1(n1294), .A2(n1125), .ZN(n1076) );
XNOR2_X1 U996 ( .A(n1295), .B(n1165), .ZN(n1294) );
NAND2_X1 U997 ( .A1(G227), .A2(n1051), .ZN(n1165) );
XOR2_X1 U998 ( .A(n1296), .B(n1297), .Z(n1295) );
NOR2_X1 U999 ( .A1(n1162), .A2(n1298), .ZN(n1297) );
NOR2_X1 U1000 ( .A1(G110), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1001 ( .A(KEYINPUT51), .B(G140), .Z(n1299) );
NOR2_X1 U1002 ( .A1(n1161), .A2(G140), .ZN(n1162) );
NAND2_X1 U1003 ( .A1(n1300), .A2(n1301), .ZN(n1296) );
NAND2_X1 U1004 ( .A1(n1158), .A2(n1166), .ZN(n1301) );
XOR2_X1 U1005 ( .A(KEYINPUT62), .B(n1302), .Z(n1300) );
NOR2_X1 U1006 ( .A1(n1158), .A2(n1166), .ZN(n1302) );
XNOR2_X1 U1007 ( .A(n1303), .B(n1289), .ZN(n1158) );
XNOR2_X1 U1008 ( .A(G107), .B(n1133), .ZN(n1289) );
INV_X1 U1009 ( .A(G104), .ZN(n1133) );
XNOR2_X1 U1010 ( .A(G101), .B(n1093), .ZN(n1303) );
XNOR2_X1 U1011 ( .A(n1071), .B(KEYINPUT55), .ZN(n1293) );
INV_X1 U1012 ( .A(n1041), .ZN(n1071) );
NAND2_X1 U1013 ( .A1(G221), .A2(n1304), .ZN(n1041) );
NOR2_X1 U1014 ( .A1(n1032), .A2(n1053), .ZN(n1030) );
INV_X1 U1015 ( .A(n1034), .ZN(n1053) );
XNOR2_X1 U1016 ( .A(n1072), .B(n1074), .ZN(n1034) );
NAND2_X1 U1017 ( .A1(G217), .A2(n1304), .ZN(n1074) );
NAND2_X1 U1018 ( .A1(G234), .A2(n1125), .ZN(n1304) );
NOR2_X1 U1019 ( .A1(n1117), .A2(G902), .ZN(n1072) );
XOR2_X1 U1020 ( .A(n1305), .B(n1306), .Z(n1117) );
XOR2_X1 U1021 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U1022 ( .A(n1161), .B(n1309), .ZN(n1308) );
NOR2_X1 U1023 ( .A1(KEYINPUT50), .A2(n1310), .ZN(n1309) );
XOR2_X1 U1024 ( .A(n1311), .B(n1270), .Z(n1310) );
XNOR2_X1 U1025 ( .A(n1312), .B(n1313), .ZN(n1270) );
XNOR2_X1 U1026 ( .A(G125), .B(G140), .ZN(n1312) );
XNOR2_X1 U1027 ( .A(KEYINPUT5), .B(KEYINPUT41), .ZN(n1311) );
INV_X1 U1028 ( .A(G110), .ZN(n1161) );
NOR2_X1 U1029 ( .A1(n1314), .A2(n1252), .ZN(n1307) );
NAND2_X1 U1030 ( .A1(G234), .A2(n1051), .ZN(n1252) );
INV_X1 U1031 ( .A(G221), .ZN(n1314) );
XNOR2_X1 U1032 ( .A(G119), .B(n1315), .ZN(n1305) );
XOR2_X1 U1033 ( .A(G137), .B(G128), .Z(n1315) );
XOR2_X1 U1034 ( .A(n1066), .B(KEYINPUT36), .Z(n1032) );
XNOR2_X1 U1035 ( .A(n1316), .B(G472), .ZN(n1066) );
NAND2_X1 U1036 ( .A1(n1317), .A2(n1125), .ZN(n1316) );
INV_X1 U1037 ( .A(G902), .ZN(n1125) );
XNOR2_X1 U1038 ( .A(n1146), .B(n1318), .ZN(n1317) );
XNOR2_X1 U1039 ( .A(n1319), .B(KEYINPUT37), .ZN(n1318) );
NAND2_X1 U1040 ( .A1(KEYINPUT20), .A2(n1320), .ZN(n1319) );
XNOR2_X1 U1041 ( .A(n1166), .B(n1143), .ZN(n1320) );
XOR2_X1 U1042 ( .A(n1321), .B(n1322), .Z(n1143) );
INV_X1 U1043 ( .A(n1279), .ZN(n1322) );
XOR2_X1 U1044 ( .A(n1111), .B(n1093), .Z(n1279) );
XNOR2_X1 U1045 ( .A(n1248), .B(n1313), .ZN(n1093) );
XOR2_X1 U1046 ( .A(G146), .B(KEYINPUT40), .Z(n1313) );
XNOR2_X1 U1047 ( .A(G128), .B(G143), .ZN(n1248) );
XNOR2_X1 U1048 ( .A(G119), .B(n1264), .ZN(n1111) );
INV_X1 U1049 ( .A(G113), .ZN(n1264) );
NAND2_X1 U1050 ( .A1(KEYINPUT31), .A2(n1236), .ZN(n1321) );
INV_X1 U1051 ( .A(G116), .ZN(n1236) );
NAND2_X1 U1052 ( .A1(n1323), .A2(n1324), .ZN(n1166) );
OR2_X1 U1053 ( .A1(n1325), .A2(G131), .ZN(n1324) );
XOR2_X1 U1054 ( .A(n1326), .B(KEYINPUT34), .Z(n1323) );
NAND2_X1 U1055 ( .A1(G131), .A2(n1325), .ZN(n1326) );
XNOR2_X1 U1056 ( .A(n1092), .B(KEYINPUT29), .ZN(n1325) );
XNOR2_X1 U1057 ( .A(G134), .B(G137), .ZN(n1092) );
XOR2_X1 U1058 ( .A(G101), .B(n1327), .Z(n1146) );
AND3_X1 U1059 ( .A1(G210), .A2(n1051), .A3(n1269), .ZN(n1327) );
INV_X1 U1060 ( .A(G237), .ZN(n1269) );
INV_X1 U1061 ( .A(G953), .ZN(n1051) );
endmodule


