//Key = 1100111001100101101101101001001110100001011011101010001000101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292;

XNOR2_X1 U720 ( .A(G107), .B(n979), .ZN(G9) );
NAND2_X1 U721 ( .A1(n980), .A2(n981), .ZN(n979) );
XNOR2_X1 U722 ( .A(n982), .B(KEYINPUT22), .ZN(n980) );
NOR2_X1 U723 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR4_X1 U724 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n984) );
XOR2_X1 U725 ( .A(n989), .B(KEYINPUT63), .Z(n987) );
NAND2_X1 U726 ( .A1(n990), .A2(n991), .ZN(n989) );
NAND2_X1 U727 ( .A1(n992), .A2(n981), .ZN(n991) );
NAND2_X1 U728 ( .A1(n993), .A2(n994), .ZN(n990) );
NAND2_X1 U729 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U730 ( .A1(n997), .A2(n998), .ZN(n996) );
NAND2_X1 U731 ( .A1(n999), .A2(n1000), .ZN(n998) );
NAND2_X1 U732 ( .A1(n1001), .A2(n1002), .ZN(n1000) );
NAND2_X1 U733 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND3_X1 U734 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
INV_X1 U735 ( .A(KEYINPUT59), .ZN(n1006) );
NAND2_X1 U736 ( .A1(n1008), .A2(n1009), .ZN(n1003) );
NAND3_X1 U737 ( .A1(n1010), .A2(n1008), .A3(n1005), .ZN(n999) );
NAND2_X1 U738 ( .A1(KEYINPUT59), .A2(n1011), .ZN(n995) );
NAND2_X1 U739 ( .A1(n1012), .A2(n1007), .ZN(n1011) );
XOR2_X1 U740 ( .A(KEYINPUT7), .B(n1013), .Z(n986) );
NOR4_X1 U741 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
NAND3_X1 U742 ( .A1(n993), .A2(n1008), .A3(n1001), .ZN(n1014) );
NAND4_X1 U743 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n985) );
NAND4_X1 U744 ( .A1(n997), .A2(n1005), .A3(n993), .A4(n1022), .ZN(n1019) );
NAND2_X1 U745 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U746 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
XNOR2_X1 U747 ( .A(n1008), .B(KEYINPUT42), .ZN(n1025) );
NAND2_X1 U748 ( .A1(n1027), .A2(n1001), .ZN(n1023) );
NAND3_X1 U749 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1018) );
XOR2_X1 U750 ( .A(KEYINPUT2), .B(n992), .Z(n1029) );
AND2_X1 U751 ( .A1(n1012), .A2(n1008), .ZN(n992) );
AND3_X1 U752 ( .A1(n1005), .A2(n1001), .A3(n997), .ZN(n1012) );
INV_X1 U753 ( .A(n1016), .ZN(n997) );
NOR3_X1 U754 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n983) );
INV_X1 U755 ( .A(n1020), .ZN(n1031) );
NAND4_X1 U756 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1020) );
NOR3_X1 U757 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
AND2_X1 U758 ( .A1(n1039), .A2(G478), .ZN(n1038) );
XNOR2_X1 U759 ( .A(n1040), .B(G475), .ZN(n1034) );
XNOR2_X1 U760 ( .A(n1041), .B(n1042), .ZN(n1033) );
XOR2_X1 U761 ( .A(n1043), .B(KEYINPUT30), .Z(n1032) );
NAND3_X1 U762 ( .A1(n1044), .A2(n1015), .A3(n993), .ZN(n1043) );
XOR2_X1 U763 ( .A(G469), .B(n1045), .Z(n1044) );
NOR2_X1 U764 ( .A1(n1046), .A2(KEYINPUT26), .ZN(n1045) );
XOR2_X1 U765 ( .A(n1047), .B(n1048), .Z(G72) );
NOR2_X1 U766 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U767 ( .A1(n1021), .A2(n1051), .ZN(n1049) );
XOR2_X1 U768 ( .A(KEYINPUT28), .B(G227), .Z(n1051) );
XOR2_X1 U769 ( .A(n1052), .B(n1053), .Z(n1047) );
NOR2_X1 U770 ( .A1(G953), .A2(n1054), .ZN(n1053) );
NAND2_X1 U771 ( .A1(n1055), .A2(n1056), .ZN(n1052) );
INV_X1 U772 ( .A(n1050), .ZN(n1056) );
XOR2_X1 U773 ( .A(n1057), .B(n1058), .Z(n1055) );
XOR2_X1 U774 ( .A(n1059), .B(n1060), .Z(n1058) );
XNOR2_X1 U775 ( .A(n1061), .B(n1062), .ZN(n1057) );
NAND2_X1 U776 ( .A1(KEYINPUT24), .A2(n1063), .ZN(n1061) );
XOR2_X1 U777 ( .A(G125), .B(n1064), .Z(n1063) );
NOR2_X1 U778 ( .A1(KEYINPUT25), .A2(n1065), .ZN(n1064) );
XOR2_X1 U779 ( .A(n1066), .B(n1067), .Z(G69) );
NOR2_X1 U780 ( .A1(n1068), .A2(n1021), .ZN(n1067) );
NOR2_X1 U781 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U782 ( .A1(n1071), .A2(n1072), .ZN(n1066) );
NAND2_X1 U783 ( .A1(n1073), .A2(n1021), .ZN(n1072) );
XNOR2_X1 U784 ( .A(n1074), .B(n1075), .ZN(n1073) );
NAND3_X1 U785 ( .A1(G898), .A2(n1075), .A3(G953), .ZN(n1071) );
NAND2_X1 U786 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NAND2_X1 U787 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XNOR2_X1 U788 ( .A(n1080), .B(n1081), .ZN(n1079) );
XNOR2_X1 U789 ( .A(KEYINPUT23), .B(KEYINPUT9), .ZN(n1078) );
NAND2_X1 U790 ( .A1(n1082), .A2(n1083), .ZN(n1076) );
XOR2_X1 U791 ( .A(n1084), .B(n1085), .Z(n1083) );
XNOR2_X1 U792 ( .A(n1086), .B(n1087), .ZN(n1085) );
XOR2_X1 U793 ( .A(KEYINPUT9), .B(KEYINPUT23), .Z(n1082) );
NOR2_X1 U794 ( .A1(n1088), .A2(n1089), .ZN(G66) );
XOR2_X1 U795 ( .A(n1090), .B(n1091), .Z(n1089) );
NOR4_X1 U796 ( .A1(n1092), .A2(n1093), .A3(KEYINPUT37), .A4(n1094), .ZN(n1090) );
NOR2_X1 U797 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
INV_X1 U798 ( .A(KEYINPUT47), .ZN(n1096) );
NOR2_X1 U799 ( .A1(n1097), .A2(n988), .ZN(n1095) );
XNOR2_X1 U800 ( .A(KEYINPUT35), .B(G902), .ZN(n1097) );
NOR2_X1 U801 ( .A1(KEYINPUT47), .A2(n1098), .ZN(n1092) );
NOR2_X1 U802 ( .A1(n1088), .A2(n1099), .ZN(G63) );
XNOR2_X1 U803 ( .A(n1100), .B(n1101), .ZN(n1099) );
AND2_X1 U804 ( .A1(G478), .A2(n1098), .ZN(n1101) );
NOR2_X1 U805 ( .A1(n1088), .A2(n1102), .ZN(G60) );
XNOR2_X1 U806 ( .A(n1103), .B(n1104), .ZN(n1102) );
AND2_X1 U807 ( .A1(G475), .A2(n1098), .ZN(n1104) );
XNOR2_X1 U808 ( .A(G104), .B(n1105), .ZN(G6) );
NOR2_X1 U809 ( .A1(n1088), .A2(n1106), .ZN(G57) );
XOR2_X1 U810 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U811 ( .A(n1109), .B(n1110), .Z(n1107) );
XOR2_X1 U812 ( .A(n1111), .B(n1112), .Z(n1110) );
AND2_X1 U813 ( .A1(G472), .A2(n1098), .ZN(n1112) );
NOR2_X1 U814 ( .A1(KEYINPUT55), .A2(n1113), .ZN(n1111) );
NOR2_X1 U815 ( .A1(n1114), .A2(n1115), .ZN(G54) );
XOR2_X1 U816 ( .A(KEYINPUT12), .B(n1088), .Z(n1115) );
XOR2_X1 U817 ( .A(n1116), .B(n1117), .Z(n1114) );
XNOR2_X1 U818 ( .A(n1118), .B(n1119), .ZN(n1117) );
NAND2_X1 U819 ( .A1(KEYINPUT46), .A2(n1120), .ZN(n1119) );
NAND2_X1 U820 ( .A1(n1098), .A2(G469), .ZN(n1120) );
INV_X1 U821 ( .A(n1121), .ZN(n1098) );
NAND2_X1 U822 ( .A1(n1122), .A2(KEYINPUT10), .ZN(n1118) );
XOR2_X1 U823 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U824 ( .A1(n1125), .A2(KEYINPUT32), .ZN(n1123) );
XOR2_X1 U825 ( .A(n1126), .B(KEYINPUT50), .Z(n1125) );
NOR2_X1 U826 ( .A1(n1088), .A2(n1127), .ZN(G51) );
XOR2_X1 U827 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U828 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U829 ( .A1(n1132), .A2(KEYINPUT21), .ZN(n1131) );
XNOR2_X1 U830 ( .A(n1133), .B(n1134), .ZN(n1132) );
NOR2_X1 U831 ( .A1(n1135), .A2(n1121), .ZN(n1128) );
NAND2_X1 U832 ( .A1(n1136), .A2(n988), .ZN(n1121) );
NAND2_X1 U833 ( .A1(n1074), .A2(n1054), .ZN(n988) );
AND4_X1 U834 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1054) );
NOR4_X1 U835 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
NOR2_X1 U836 ( .A1(n1145), .A2(n1146), .ZN(n1139) );
NOR2_X1 U837 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XNOR2_X1 U838 ( .A(n1027), .B(KEYINPUT62), .ZN(n1147) );
NOR3_X1 U839 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1145) );
XNOR2_X1 U840 ( .A(n1027), .B(KEYINPUT56), .ZN(n1150) );
AND4_X1 U841 ( .A1(n1152), .A2(n1105), .A3(n1153), .A4(n1154), .ZN(n1074) );
NOR3_X1 U842 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1154) );
NOR2_X1 U843 ( .A1(n1158), .A2(n1159), .ZN(n1155) );
NOR2_X1 U844 ( .A1(n982), .A2(n1160), .ZN(n1158) );
NOR2_X1 U845 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U846 ( .A1(n1163), .A2(n1164), .ZN(n1161) );
AND4_X1 U847 ( .A1(n1008), .A2(n1009), .A3(n1026), .A4(n1165), .ZN(n982) );
NAND4_X1 U848 ( .A1(n1166), .A2(n1010), .A3(n1008), .A4(n1165), .ZN(n1105) );
XNOR2_X1 U849 ( .A(KEYINPUT35), .B(n1167), .ZN(n1136) );
NOR2_X1 U850 ( .A1(n1021), .A2(G952), .ZN(n1088) );
XNOR2_X1 U851 ( .A(G146), .B(n1137), .ZN(G48) );
NAND4_X1 U852 ( .A1(n1168), .A2(n1169), .A3(n1009), .A4(n1036), .ZN(n1137) );
INV_X1 U853 ( .A(n1149), .ZN(n1169) );
XNOR2_X1 U854 ( .A(G143), .B(n1170), .ZN(G45) );
NOR2_X1 U855 ( .A1(n1144), .A2(KEYINPUT52), .ZN(n1170) );
AND3_X1 U856 ( .A1(n1007), .A2(n1166), .A3(n1171), .ZN(n1144) );
NOR3_X1 U857 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
XNOR2_X1 U858 ( .A(G140), .B(n1175), .ZN(G42) );
OR2_X1 U859 ( .A1(n1148), .A2(n1176), .ZN(n1175) );
NAND2_X1 U860 ( .A1(n1177), .A2(n1010), .ZN(n1148) );
XOR2_X1 U861 ( .A(G137), .B(n1143), .Z(G39) );
AND2_X1 U862 ( .A1(n1163), .A2(n1177), .ZN(n1143) );
XOR2_X1 U863 ( .A(G134), .B(n1142), .Z(G36) );
AND3_X1 U864 ( .A1(n1007), .A2(n1026), .A3(n1177), .ZN(n1142) );
XOR2_X1 U865 ( .A(n1178), .B(G131), .Z(G33) );
NAND2_X1 U866 ( .A1(KEYINPUT18), .A2(n1138), .ZN(n1178) );
NAND2_X1 U867 ( .A1(n1164), .A2(n1177), .ZN(n1138) );
AND3_X1 U868 ( .A1(n1009), .A2(n1179), .A3(n993), .ZN(n1177) );
NOR2_X1 U869 ( .A1(n1180), .A2(n1030), .ZN(n993) );
XOR2_X1 U870 ( .A(n1141), .B(n1181), .Z(G30) );
NOR2_X1 U871 ( .A1(KEYINPUT38), .A2(n1182), .ZN(n1181) );
AND3_X1 U872 ( .A1(n1168), .A2(n1166), .A3(n1183), .ZN(n1141) );
NOR3_X1 U873 ( .A1(n1184), .A2(n1174), .A3(n1185), .ZN(n1183) );
INV_X1 U874 ( .A(n1179), .ZN(n1174) );
XOR2_X1 U875 ( .A(G101), .B(n1157), .Z(G3) );
AND2_X1 U876 ( .A1(n1007), .A2(n1186), .ZN(n1157) );
XOR2_X1 U877 ( .A(G125), .B(n1187), .Z(G27) );
NOR3_X1 U878 ( .A1(n1149), .A2(n1176), .A3(n1151), .ZN(n1187) );
NAND3_X1 U879 ( .A1(n981), .A2(n1179), .A3(n1010), .ZN(n1149) );
NAND2_X1 U880 ( .A1(n1016), .A2(n1188), .ZN(n1179) );
NAND3_X1 U881 ( .A1(G902), .A2(n1189), .A3(n1050), .ZN(n1188) );
NOR2_X1 U882 ( .A1(G900), .A2(n1021), .ZN(n1050) );
NAND2_X1 U883 ( .A1(n1190), .A2(n1191), .ZN(G24) );
NAND2_X1 U884 ( .A1(n1156), .A2(n1192), .ZN(n1191) );
XOR2_X1 U885 ( .A(n1193), .B(KEYINPUT20), .Z(n1190) );
OR2_X1 U886 ( .A1(n1192), .A2(n1156), .ZN(n1193) );
NOR4_X1 U887 ( .A1(n1172), .A2(n1162), .A3(n1194), .A4(n1159), .ZN(n1156) );
NAND2_X1 U888 ( .A1(n1195), .A2(n1008), .ZN(n1194) );
NOR2_X1 U889 ( .A1(n1036), .A2(n1168), .ZN(n1008) );
XNOR2_X1 U890 ( .A(G119), .B(n1196), .ZN(G21) );
NAND3_X1 U891 ( .A1(n1163), .A2(n1197), .A3(n1198), .ZN(n1196) );
XNOR2_X1 U892 ( .A(n981), .B(KEYINPUT61), .ZN(n1198) );
AND3_X1 U893 ( .A1(n1168), .A2(n1036), .A3(n1001), .ZN(n1163) );
XNOR2_X1 U894 ( .A(G116), .B(n1153), .ZN(G18) );
NAND4_X1 U895 ( .A1(n1007), .A2(n1197), .A3(n981), .A4(n1026), .ZN(n1153) );
INV_X1 U896 ( .A(n1184), .ZN(n1026) );
NAND2_X1 U897 ( .A1(n1199), .A2(n1195), .ZN(n1184) );
XNOR2_X1 U898 ( .A(G113), .B(n1200), .ZN(G15) );
NAND4_X1 U899 ( .A1(KEYINPUT41), .A2(n1164), .A3(n1197), .A4(n1201), .ZN(n1200) );
XNOR2_X1 U900 ( .A(KEYINPUT40), .B(n1159), .ZN(n1201) );
INV_X1 U901 ( .A(n981), .ZN(n1159) );
INV_X1 U902 ( .A(n1162), .ZN(n1197) );
NAND2_X1 U903 ( .A1(n1005), .A2(n1165), .ZN(n1162) );
INV_X1 U904 ( .A(n1151), .ZN(n1005) );
NAND2_X1 U905 ( .A1(n1202), .A2(n1015), .ZN(n1151) );
INV_X1 U906 ( .A(n1017), .ZN(n1202) );
XOR2_X1 U907 ( .A(n1203), .B(KEYINPUT57), .Z(n1017) );
AND2_X1 U908 ( .A1(n1007), .A2(n1010), .ZN(n1164) );
NOR2_X1 U909 ( .A1(n1195), .A2(n1172), .ZN(n1010) );
XNOR2_X1 U910 ( .A(n1204), .B(KEYINPUT16), .ZN(n1172) );
NOR2_X1 U911 ( .A1(n1168), .A2(n1185), .ZN(n1007) );
XNOR2_X1 U912 ( .A(G110), .B(n1152), .ZN(G12) );
NAND2_X1 U913 ( .A1(n1027), .A2(n1186), .ZN(n1152) );
AND3_X1 U914 ( .A1(n1166), .A2(n1165), .A3(n1001), .ZN(n1186) );
AND2_X1 U915 ( .A1(n1205), .A2(n1199), .ZN(n1001) );
XNOR2_X1 U916 ( .A(n1204), .B(KEYINPUT15), .ZN(n1199) );
XNOR2_X1 U917 ( .A(n1206), .B(n1207), .ZN(n1204) );
INV_X1 U918 ( .A(n1040), .ZN(n1207) );
NOR2_X1 U919 ( .A1(n1208), .A2(G902), .ZN(n1040) );
INV_X1 U920 ( .A(n1103), .ZN(n1208) );
XNOR2_X1 U921 ( .A(n1209), .B(n1210), .ZN(n1103) );
XNOR2_X1 U922 ( .A(n1211), .B(n1212), .ZN(n1210) );
XOR2_X1 U923 ( .A(n1213), .B(G131), .Z(n1212) );
NAND3_X1 U924 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1213) );
NAND2_X1 U925 ( .A1(n1217), .A2(G143), .ZN(n1216) );
NAND2_X1 U926 ( .A1(KEYINPUT8), .A2(n1218), .ZN(n1215) );
NAND2_X1 U927 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
INV_X1 U928 ( .A(G143), .ZN(n1220) );
XNOR2_X1 U929 ( .A(n1217), .B(KEYINPUT29), .ZN(n1219) );
NAND2_X1 U930 ( .A1(n1221), .A2(n1222), .ZN(n1214) );
INV_X1 U931 ( .A(KEYINPUT8), .ZN(n1222) );
NAND2_X1 U932 ( .A1(n1223), .A2(n1224), .ZN(n1221) );
OR3_X1 U933 ( .A1(n1217), .A2(G143), .A3(KEYINPUT29), .ZN(n1224) );
NAND2_X1 U934 ( .A1(KEYINPUT29), .A2(n1217), .ZN(n1223) );
AND3_X1 U935 ( .A1(n1225), .A2(n1021), .A3(G214), .ZN(n1217) );
XNOR2_X1 U936 ( .A(n1226), .B(n1086), .ZN(n1209) );
XNOR2_X1 U937 ( .A(G113), .B(n1192), .ZN(n1086) );
NAND2_X1 U938 ( .A1(KEYINPUT13), .A2(G475), .ZN(n1206) );
XNOR2_X1 U939 ( .A(n1173), .B(KEYINPUT45), .ZN(n1205) );
INV_X1 U940 ( .A(n1195), .ZN(n1173) );
NAND2_X1 U941 ( .A1(n1227), .A2(n1228), .ZN(n1195) );
NAND2_X1 U942 ( .A1(G478), .A2(n1039), .ZN(n1228) );
XOR2_X1 U943 ( .A(KEYINPUT6), .B(n1037), .Z(n1227) );
NOR2_X1 U944 ( .A1(n1039), .A2(G478), .ZN(n1037) );
NAND2_X1 U945 ( .A1(n1100), .A2(n1167), .ZN(n1039) );
XNOR2_X1 U946 ( .A(n1229), .B(n1230), .ZN(n1100) );
XOR2_X1 U947 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U948 ( .A(G107), .B(n1233), .Z(n1232) );
NOR2_X1 U949 ( .A1(KEYINPUT51), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U950 ( .A(n1235), .B(n1182), .ZN(n1234) );
NAND2_X1 U951 ( .A1(KEYINPUT58), .A2(G143), .ZN(n1235) );
AND3_X1 U952 ( .A1(G217), .A2(n1021), .A3(G234), .ZN(n1231) );
XNOR2_X1 U953 ( .A(G116), .B(n1236), .ZN(n1229) );
XNOR2_X1 U954 ( .A(G134), .B(n1192), .ZN(n1236) );
INV_X1 U955 ( .A(G122), .ZN(n1192) );
NAND2_X1 U956 ( .A1(n1016), .A2(n1237), .ZN(n1165) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1189), .A4(n1070), .ZN(n1237) );
INV_X1 U958 ( .A(G898), .ZN(n1070) );
NAND3_X1 U959 ( .A1(n1189), .A2(n1021), .A3(G952), .ZN(n1016) );
NAND2_X1 U960 ( .A1(G237), .A2(G234), .ZN(n1189) );
AND2_X1 U961 ( .A1(n981), .A2(n1009), .ZN(n1166) );
AND2_X1 U962 ( .A1(n1203), .A2(n1015), .ZN(n1009) );
NAND2_X1 U963 ( .A1(G221), .A2(n1238), .ZN(n1015) );
XOR2_X1 U964 ( .A(n1046), .B(G469), .Z(n1203) );
AND2_X1 U965 ( .A1(n1239), .A2(n1167), .ZN(n1046) );
XOR2_X1 U966 ( .A(n1240), .B(n1116), .Z(n1239) );
XOR2_X1 U967 ( .A(n1241), .B(n1242), .Z(n1116) );
XNOR2_X1 U968 ( .A(n1243), .B(n1244), .ZN(n1242) );
INV_X1 U969 ( .A(n1211), .ZN(n1243) );
XOR2_X1 U970 ( .A(G146), .B(n1245), .Z(n1211) );
XOR2_X1 U971 ( .A(n1246), .B(n1059), .Z(n1241) );
XNOR2_X1 U972 ( .A(n1247), .B(G143), .ZN(n1059) );
NAND2_X1 U973 ( .A1(KEYINPUT0), .A2(n1182), .ZN(n1247) );
NAND3_X1 U974 ( .A1(n1248), .A2(n1249), .A3(KEYINPUT4), .ZN(n1240) );
NAND2_X1 U975 ( .A1(n1124), .A2(n1126), .ZN(n1249) );
XOR2_X1 U976 ( .A(KEYINPUT39), .B(n1250), .Z(n1248) );
NOR2_X1 U977 ( .A1(n1124), .A2(n1126), .ZN(n1250) );
XNOR2_X1 U978 ( .A(n1087), .B(n1251), .ZN(n1126) );
XNOR2_X1 U979 ( .A(KEYINPUT33), .B(n1065), .ZN(n1251) );
AND2_X1 U980 ( .A1(G227), .A2(n1021), .ZN(n1124) );
NOR2_X1 U981 ( .A1(n1028), .A2(n1030), .ZN(n981) );
AND2_X1 U982 ( .A1(G214), .A2(n1252), .ZN(n1030) );
XOR2_X1 U983 ( .A(KEYINPUT44), .B(n1253), .Z(n1252) );
NOR2_X1 U984 ( .A1(G237), .A2(G902), .ZN(n1253) );
INV_X1 U985 ( .A(n1180), .ZN(n1028) );
XOR2_X1 U986 ( .A(n1254), .B(n1135), .Z(n1180) );
NAND2_X1 U987 ( .A1(G210), .A2(n1255), .ZN(n1135) );
NAND2_X1 U988 ( .A1(n1225), .A2(n1167), .ZN(n1255) );
NAND2_X1 U989 ( .A1(n1256), .A2(n1167), .ZN(n1254) );
XNOR2_X1 U990 ( .A(n1257), .B(n1258), .ZN(n1256) );
XOR2_X1 U991 ( .A(n1130), .B(n1259), .Z(n1258) );
NAND2_X1 U992 ( .A1(KEYINPUT60), .A2(n1134), .ZN(n1259) );
NOR2_X1 U993 ( .A1(n1069), .A2(G953), .ZN(n1134) );
INV_X1 U994 ( .A(G224), .ZN(n1069) );
NAND2_X1 U995 ( .A1(n1260), .A2(n1261), .ZN(n1130) );
OR2_X1 U996 ( .A1(n1081), .A2(n1080), .ZN(n1261) );
XOR2_X1 U997 ( .A(n1262), .B(KEYINPUT11), .Z(n1260) );
NAND2_X1 U998 ( .A1(n1080), .A2(n1081), .ZN(n1262) );
XOR2_X1 U999 ( .A(G122), .B(n1087), .Z(n1081) );
XOR2_X1 U1000 ( .A(n1084), .B(n1263), .Z(n1080) );
XOR2_X1 U1001 ( .A(n1264), .B(n1244), .Z(n1084) );
XOR2_X1 U1002 ( .A(G101), .B(G107), .Z(n1244) );
XOR2_X1 U1003 ( .A(n1265), .B(n1245), .Z(n1264) );
XOR2_X1 U1004 ( .A(G104), .B(KEYINPUT5), .Z(n1245) );
NAND2_X1 U1005 ( .A1(KEYINPUT1), .A2(n1266), .ZN(n1265) );
INV_X1 U1006 ( .A(n1133), .ZN(n1257) );
XOR2_X1 U1007 ( .A(G125), .B(n1113), .Z(n1133) );
INV_X1 U1008 ( .A(n1176), .ZN(n1027) );
NAND2_X1 U1009 ( .A1(n1168), .A2(n1185), .ZN(n1176) );
INV_X1 U1010 ( .A(n1036), .ZN(n1185) );
XNOR2_X1 U1011 ( .A(n1267), .B(G472), .ZN(n1036) );
NAND2_X1 U1012 ( .A1(n1268), .A2(n1167), .ZN(n1267) );
XOR2_X1 U1013 ( .A(n1269), .B(n1108), .Z(n1268) );
XOR2_X1 U1014 ( .A(n1270), .B(n1246), .Z(n1108) );
NAND2_X1 U1015 ( .A1(n1271), .A2(n1272), .ZN(n1246) );
NAND3_X1 U1016 ( .A1(G131), .A2(n1273), .A3(n1274), .ZN(n1272) );
INV_X1 U1017 ( .A(KEYINPUT27), .ZN(n1274) );
NAND2_X1 U1018 ( .A1(n1060), .A2(KEYINPUT27), .ZN(n1271) );
XOR2_X1 U1019 ( .A(G131), .B(n1273), .Z(n1060) );
XOR2_X1 U1020 ( .A(G134), .B(G137), .Z(n1273) );
XOR2_X1 U1021 ( .A(n1275), .B(G101), .Z(n1270) );
NAND3_X1 U1022 ( .A1(n1225), .A2(n1021), .A3(G210), .ZN(n1275) );
INV_X1 U1023 ( .A(G237), .ZN(n1225) );
XNOR2_X1 U1024 ( .A(n1113), .B(n1276), .ZN(n1269) );
XNOR2_X1 U1025 ( .A(n1277), .B(KEYINPUT54), .ZN(n1276) );
NAND2_X1 U1026 ( .A1(KEYINPUT19), .A2(n1109), .ZN(n1277) );
XNOR2_X1 U1027 ( .A(n1263), .B(n1278), .ZN(n1109) );
NOR2_X1 U1028 ( .A1(KEYINPUT17), .A2(n1266), .ZN(n1278) );
XNOR2_X1 U1029 ( .A(G116), .B(G119), .ZN(n1266) );
INV_X1 U1030 ( .A(G113), .ZN(n1263) );
XNOR2_X1 U1031 ( .A(n1279), .B(n1280), .ZN(n1113) );
NOR2_X1 U1032 ( .A1(G146), .A2(KEYINPUT43), .ZN(n1280) );
XNOR2_X1 U1033 ( .A(G143), .B(n1281), .ZN(n1279) );
NOR2_X1 U1034 ( .A1(KEYINPUT53), .A2(n1182), .ZN(n1281) );
INV_X1 U1035 ( .A(G128), .ZN(n1182) );
XNOR2_X1 U1036 ( .A(n1042), .B(n1282), .ZN(n1168) );
NOR2_X1 U1037 ( .A1(n1041), .A2(KEYINPUT36), .ZN(n1282) );
INV_X1 U1038 ( .A(n1094), .ZN(n1041) );
NAND2_X1 U1039 ( .A1(G217), .A2(n1238), .ZN(n1094) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1167), .ZN(n1238) );
AND2_X1 U1041 ( .A1(n1283), .A2(n1167), .ZN(n1042) );
INV_X1 U1042 ( .A(G902), .ZN(n1167) );
XNOR2_X1 U1043 ( .A(n1091), .B(KEYINPUT49), .ZN(n1283) );
XNOR2_X1 U1044 ( .A(n1284), .B(n1285), .ZN(n1091) );
XNOR2_X1 U1045 ( .A(n1286), .B(n1087), .ZN(n1285) );
XOR2_X1 U1046 ( .A(G110), .B(KEYINPUT34), .Z(n1087) );
NAND2_X1 U1047 ( .A1(KEYINPUT48), .A2(n1287), .ZN(n1286) );
XOR2_X1 U1048 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U1049 ( .A(G137), .B(KEYINPUT3), .ZN(n1289) );
NAND3_X1 U1050 ( .A1(G221), .A2(n1021), .A3(G234), .ZN(n1288) );
INV_X1 U1051 ( .A(G953), .ZN(n1021) );
XOR2_X1 U1052 ( .A(n1290), .B(n1291), .Z(n1284) );
NOR2_X1 U1053 ( .A1(KEYINPUT14), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U1054 ( .A(n1062), .B(n1226), .ZN(n1292) );
XNOR2_X1 U1055 ( .A(G125), .B(n1065), .ZN(n1226) );
XNOR2_X1 U1056 ( .A(G140), .B(KEYINPUT31), .ZN(n1065) );
INV_X1 U1057 ( .A(G146), .ZN(n1062) );
XNOR2_X1 U1058 ( .A(G119), .B(G128), .ZN(n1290) );
endmodule


