//Key = 1001010100011010101001110000010100111010110010010101110000110101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378;

XNOR2_X1 U750 ( .A(G107), .B(n1040), .ZN(G9) );
NOR2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(G75) );
NOR4_X1 U752 ( .A1(n1043), .A2(n1044), .A3(KEYINPUT25), .A4(G953), .ZN(n1042) );
NAND2_X1 U753 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND3_X1 U756 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NAND2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U760 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
INV_X1 U761 ( .A(KEYINPUT19), .ZN(n1061) );
NAND2_X1 U762 ( .A1(KEYINPUT35), .A2(n1062), .ZN(n1058) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1054) );
NAND3_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1064) );
INV_X1 U765 ( .A(n1068), .ZN(n1067) );
NAND3_X1 U766 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1066) );
NAND2_X1 U767 ( .A1(KEYINPUT56), .A2(n1072), .ZN(n1065) );
NAND2_X1 U768 ( .A1(n1056), .A2(n1073), .ZN(n1049) );
NAND3_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NAND2_X1 U770 ( .A1(n1063), .A2(n1077), .ZN(n1076) );
NAND2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U772 ( .A1(n1053), .A2(n1080), .ZN(n1079) );
OR2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1051), .A2(n1083), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NAND2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
INV_X1 U777 ( .A(n1088), .ZN(n1084) );
NAND4_X1 U778 ( .A1(n1053), .A2(n1060), .A3(KEYINPUT19), .A4(n1089), .ZN(n1075) );
INV_X1 U779 ( .A(n1051), .ZN(n1089) );
NAND4_X1 U780 ( .A1(n1090), .A2(n1091), .A3(n1062), .A4(n1051), .ZN(n1074) );
INV_X1 U781 ( .A(KEYINPUT35), .ZN(n1091) );
INV_X1 U782 ( .A(n1092), .ZN(n1045) );
NOR3_X1 U783 ( .A1(n1044), .A2(G953), .A3(G952), .ZN(n1041) );
AND4_X1 U784 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1044) );
NOR4_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1090), .A4(n1072), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1099), .B(n1100), .Z(n1097) );
NOR2_X1 U787 ( .A1(G475), .A2(KEYINPUT60), .ZN(n1100) );
NOR3_X1 U788 ( .A1(n1101), .A2(n1102), .A3(n1069), .ZN(n1095) );
NAND2_X1 U789 ( .A1(G472), .A2(n1103), .ZN(n1094) );
XOR2_X1 U790 ( .A(KEYINPUT51), .B(n1104), .Z(n1093) );
XOR2_X1 U791 ( .A(n1105), .B(n1106), .Z(G72) );
XOR2_X1 U792 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
INV_X1 U794 ( .A(n1111), .ZN(n1110) );
XOR2_X1 U795 ( .A(KEYINPUT42), .B(n1112), .Z(n1109) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U797 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U798 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U799 ( .A1(KEYINPUT58), .A2(n1119), .ZN(n1118) );
NOR2_X1 U800 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
NOR3_X1 U801 ( .A1(n1122), .A2(n1120), .A3(n1121), .ZN(n1113) );
XNOR2_X1 U802 ( .A(KEYINPUT27), .B(n1123), .ZN(n1121) );
INV_X1 U803 ( .A(KEYINPUT29), .ZN(n1120) );
XOR2_X1 U804 ( .A(n1117), .B(n1124), .Z(n1122) );
NAND2_X1 U805 ( .A1(KEYINPUT58), .A2(n1125), .ZN(n1124) );
INV_X1 U806 ( .A(n1119), .ZN(n1125) );
XOR2_X1 U807 ( .A(G125), .B(KEYINPUT1), .Z(n1119) );
NAND2_X1 U808 ( .A1(n1126), .A2(n1127), .ZN(n1117) );
NAND2_X1 U809 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U810 ( .A(KEYINPUT59), .B(n1130), .Z(n1126) );
NOR2_X1 U811 ( .A1(n1129), .A2(n1128), .ZN(n1130) );
XNOR2_X1 U812 ( .A(n1131), .B(n1132), .ZN(n1128) );
NAND2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1107) );
NAND2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XNOR2_X1 U815 ( .A(KEYINPUT5), .B(n1137), .ZN(n1136) );
XNOR2_X1 U816 ( .A(KEYINPUT12), .B(n1138), .ZN(n1133) );
NOR2_X1 U817 ( .A1(n1139), .A2(n1138), .ZN(n1105) );
AND2_X1 U818 ( .A1(G227), .A2(G900), .ZN(n1139) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(G69) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U821 ( .A1(G953), .A2(n1144), .ZN(n1143) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1144) );
NAND2_X1 U823 ( .A1(n1145), .A2(n1146), .ZN(n1142) );
NAND2_X1 U824 ( .A1(G953), .A2(n1147), .ZN(n1146) );
XOR2_X1 U825 ( .A(n1148), .B(n1149), .Z(n1145) );
XNOR2_X1 U826 ( .A(n1150), .B(G110), .ZN(n1149) );
NOR2_X1 U827 ( .A1(n1151), .A2(G953), .ZN(n1140) );
NOR3_X1 U828 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(G66) );
AND2_X1 U829 ( .A1(KEYINPUT44), .A2(n1155), .ZN(n1154) );
NOR2_X1 U830 ( .A1(KEYINPUT44), .A2(n1156), .ZN(n1153) );
XNOR2_X1 U831 ( .A(n1157), .B(n1158), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U833 ( .A1(n1155), .A2(n1161), .ZN(G63) );
XNOR2_X1 U834 ( .A(n1162), .B(n1163), .ZN(n1161) );
NOR2_X1 U835 ( .A1(n1164), .A2(n1160), .ZN(n1163) );
INV_X1 U836 ( .A(G478), .ZN(n1164) );
NOR3_X1 U837 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(G60) );
NOR2_X1 U838 ( .A1(n1156), .A2(n1168), .ZN(n1167) );
AND2_X1 U839 ( .A1(n1168), .A2(n1155), .ZN(n1166) );
INV_X1 U840 ( .A(KEYINPUT39), .ZN(n1168) );
XOR2_X1 U841 ( .A(n1169), .B(n1170), .Z(n1165) );
NOR2_X1 U842 ( .A1(n1171), .A2(KEYINPUT32), .ZN(n1169) );
NOR2_X1 U843 ( .A1(n1172), .A2(n1160), .ZN(n1171) );
XNOR2_X1 U844 ( .A(G104), .B(n1173), .ZN(G6) );
NOR2_X1 U845 ( .A1(n1155), .A2(n1174), .ZN(G57) );
XOR2_X1 U846 ( .A(n1175), .B(n1176), .Z(n1174) );
XOR2_X1 U847 ( .A(n1177), .B(n1178), .Z(n1176) );
NAND2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NAND2_X1 U849 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U850 ( .A(KEYINPUT14), .B(n1183), .Z(n1179) );
NOR2_X1 U851 ( .A1(n1181), .A2(n1182), .ZN(n1183) );
XNOR2_X1 U852 ( .A(KEYINPUT10), .B(n1184), .ZN(n1182) );
NAND2_X1 U853 ( .A1(KEYINPUT41), .A2(n1185), .ZN(n1177) );
XOR2_X1 U854 ( .A(n1186), .B(n1187), .Z(n1185) );
XOR2_X1 U855 ( .A(KEYINPUT8), .B(KEYINPUT2), .Z(n1187) );
NOR2_X1 U856 ( .A1(n1188), .A2(n1160), .ZN(n1175) );
INV_X1 U857 ( .A(G472), .ZN(n1188) );
NOR3_X1 U858 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(G54) );
AND2_X1 U859 ( .A1(n1155), .A2(KEYINPUT53), .ZN(n1191) );
NOR2_X1 U860 ( .A1(KEYINPUT53), .A2(n1156), .ZN(n1190) );
NAND2_X1 U861 ( .A1(G952), .A2(G953), .ZN(n1156) );
XOR2_X1 U862 ( .A(n1192), .B(n1193), .Z(n1189) );
NOR2_X1 U863 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U864 ( .A1(KEYINPUT48), .A2(n1196), .ZN(n1195) );
AND2_X1 U865 ( .A1(KEYINPUT57), .A2(n1196), .ZN(n1194) );
XNOR2_X1 U866 ( .A(n1197), .B(n1198), .ZN(n1196) );
XNOR2_X1 U867 ( .A(G110), .B(G140), .ZN(n1197) );
NOR2_X1 U868 ( .A1(n1199), .A2(n1160), .ZN(n1192) );
NOR2_X1 U869 ( .A1(n1155), .A2(n1200), .ZN(G51) );
XOR2_X1 U870 ( .A(n1201), .B(n1202), .Z(n1200) );
XNOR2_X1 U871 ( .A(n1203), .B(n1204), .ZN(n1202) );
NOR2_X1 U872 ( .A1(n1205), .A2(n1160), .ZN(n1204) );
NAND2_X1 U873 ( .A1(G902), .A2(n1092), .ZN(n1160) );
NAND3_X1 U874 ( .A1(n1135), .A2(n1137), .A3(n1151), .ZN(n1092) );
AND2_X1 U875 ( .A1(n1206), .A2(n1207), .ZN(n1151) );
AND4_X1 U876 ( .A1(n1173), .A2(n1040), .A3(n1208), .A4(n1209), .ZN(n1207) );
NAND4_X1 U877 ( .A1(n1210), .A2(n1068), .A3(n1060), .A4(n1051), .ZN(n1040) );
NAND4_X1 U878 ( .A1(n1062), .A2(n1210), .A3(n1068), .A4(n1051), .ZN(n1173) );
AND4_X1 U879 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1206) );
NAND2_X1 U880 ( .A1(n1056), .A2(n1215), .ZN(n1214) );
INV_X1 U881 ( .A(n1216), .ZN(n1215) );
AND4_X1 U882 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1135) );
NOR4_X1 U883 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1220) );
INV_X1 U884 ( .A(n1225), .ZN(n1224) );
NAND2_X1 U885 ( .A1(n1226), .A2(n1227), .ZN(n1219) );
XNOR2_X1 U886 ( .A(KEYINPUT4), .B(n1228), .ZN(n1227) );
INV_X1 U887 ( .A(n1229), .ZN(n1226) );
NAND4_X1 U888 ( .A1(n1230), .A2(n1068), .A3(n1231), .A4(n1232), .ZN(n1217) );
XNOR2_X1 U889 ( .A(KEYINPUT45), .B(n1090), .ZN(n1231) );
INV_X1 U890 ( .A(n1233), .ZN(n1230) );
XNOR2_X1 U891 ( .A(n1234), .B(n1235), .ZN(n1201) );
NOR2_X1 U892 ( .A1(n1138), .A2(G952), .ZN(n1155) );
XNOR2_X1 U893 ( .A(n1236), .B(n1237), .ZN(G48) );
NOR2_X1 U894 ( .A1(n1228), .A2(n1229), .ZN(n1237) );
NAND2_X1 U895 ( .A1(n1238), .A2(n1062), .ZN(n1229) );
INV_X1 U896 ( .A(n1239), .ZN(n1228) );
XNOR2_X1 U897 ( .A(n1240), .B(n1218), .ZN(G45) );
NAND4_X1 U898 ( .A1(n1238), .A2(n1081), .A3(n1241), .A4(n1242), .ZN(n1218) );
NAND2_X1 U899 ( .A1(KEYINPUT40), .A2(n1243), .ZN(n1240) );
NAND2_X1 U900 ( .A1(n1244), .A2(n1245), .ZN(G42) );
OR2_X1 U901 ( .A1(n1137), .A2(G140), .ZN(n1245) );
XOR2_X1 U902 ( .A(n1246), .B(KEYINPUT9), .Z(n1244) );
NAND2_X1 U903 ( .A1(G140), .A2(n1137), .ZN(n1246) );
NAND3_X1 U904 ( .A1(n1082), .A2(n1062), .A3(n1247), .ZN(n1137) );
XOR2_X1 U905 ( .A(G137), .B(n1248), .Z(G39) );
NOR2_X1 U906 ( .A1(n1249), .A2(n1233), .ZN(n1248) );
NAND2_X1 U907 ( .A1(n1239), .A2(n1063), .ZN(n1233) );
XNOR2_X1 U908 ( .A(n1250), .B(n1223), .ZN(G36) );
AND3_X1 U909 ( .A1(n1081), .A2(n1060), .A3(n1247), .ZN(n1223) );
XNOR2_X1 U910 ( .A(n1131), .B(n1222), .ZN(G33) );
AND3_X1 U911 ( .A1(n1081), .A2(n1062), .A3(n1247), .ZN(n1222) );
INV_X1 U912 ( .A(n1249), .ZN(n1247) );
NAND3_X1 U913 ( .A1(n1068), .A2(n1232), .A3(n1053), .ZN(n1249) );
INV_X1 U914 ( .A(n1090), .ZN(n1053) );
NAND2_X1 U915 ( .A1(n1087), .A2(n1251), .ZN(n1090) );
XNOR2_X1 U916 ( .A(n1252), .B(n1253), .ZN(G30) );
NAND2_X1 U917 ( .A1(KEYINPUT18), .A2(n1225), .ZN(n1252) );
NAND3_X1 U918 ( .A1(n1239), .A2(n1060), .A3(n1238), .ZN(n1225) );
AND3_X1 U919 ( .A1(n1088), .A2(n1232), .A3(n1068), .ZN(n1238) );
XNOR2_X1 U920 ( .A(G101), .B(n1213), .ZN(G3) );
NAND3_X1 U921 ( .A1(n1254), .A2(n1068), .A3(n1081), .ZN(n1213) );
XOR2_X1 U922 ( .A(G125), .B(n1221), .Z(G27) );
AND4_X1 U923 ( .A1(n1056), .A2(n1232), .A3(n1088), .A4(n1255), .ZN(n1221) );
AND2_X1 U924 ( .A1(n1062), .A2(n1082), .ZN(n1255) );
NAND2_X1 U925 ( .A1(n1256), .A2(n1257), .ZN(n1232) );
NAND3_X1 U926 ( .A1(G902), .A2(n1048), .A3(n1111), .ZN(n1257) );
NOR2_X1 U927 ( .A1(n1138), .A2(G900), .ZN(n1111) );
XNOR2_X1 U928 ( .A(G122), .B(n1212), .ZN(G24) );
NAND4_X1 U929 ( .A1(n1210), .A2(n1051), .A3(n1258), .A4(n1056), .ZN(n1212) );
NOR2_X1 U930 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
NOR2_X1 U931 ( .A1(n1261), .A2(n1098), .ZN(n1051) );
XNOR2_X1 U932 ( .A(G119), .B(n1211), .ZN(G21) );
NAND3_X1 U933 ( .A1(n1254), .A2(n1056), .A3(n1239), .ZN(n1211) );
NOR2_X1 U934 ( .A1(n1262), .A2(n1263), .ZN(n1239) );
NAND2_X1 U935 ( .A1(n1264), .A2(n1265), .ZN(G18) );
NAND2_X1 U936 ( .A1(G116), .A2(n1209), .ZN(n1265) );
XOR2_X1 U937 ( .A(KEYINPUT36), .B(n1266), .Z(n1264) );
NOR2_X1 U938 ( .A1(G116), .A2(n1209), .ZN(n1266) );
NAND4_X1 U939 ( .A1(n1081), .A2(n1210), .A3(n1060), .A4(n1056), .ZN(n1209) );
NOR2_X1 U940 ( .A1(n1241), .A2(n1259), .ZN(n1060) );
XOR2_X1 U941 ( .A(G113), .B(n1267), .Z(G15) );
NOR2_X1 U942 ( .A1(n1268), .A2(n1216), .ZN(n1267) );
NAND3_X1 U943 ( .A1(n1062), .A2(n1210), .A3(n1081), .ZN(n1216) );
NOR2_X1 U944 ( .A1(n1098), .A2(n1263), .ZN(n1081) );
NOR2_X1 U945 ( .A1(n1242), .A2(n1260), .ZN(n1062) );
INV_X1 U946 ( .A(n1241), .ZN(n1260) );
XNOR2_X1 U947 ( .A(KEYINPUT20), .B(n1056), .ZN(n1268) );
NAND2_X1 U948 ( .A1(n1269), .A2(n1270), .ZN(n1056) );
NAND3_X1 U949 ( .A1(n1070), .A2(n1271), .A3(n1071), .ZN(n1270) );
INV_X1 U950 ( .A(KEYINPUT56), .ZN(n1071) );
NAND2_X1 U951 ( .A1(KEYINPUT56), .A2(n1068), .ZN(n1269) );
XOR2_X1 U952 ( .A(n1208), .B(n1272), .Z(G12) );
XNOR2_X1 U953 ( .A(G110), .B(KEYINPUT24), .ZN(n1272) );
NAND3_X1 U954 ( .A1(n1082), .A2(n1068), .A3(n1254), .ZN(n1208) );
AND2_X1 U955 ( .A1(n1063), .A2(n1210), .ZN(n1254) );
AND2_X1 U956 ( .A1(n1088), .A2(n1273), .ZN(n1210) );
NAND2_X1 U957 ( .A1(n1256), .A2(n1274), .ZN(n1273) );
NAND4_X1 U958 ( .A1(G953), .A2(G902), .A3(n1048), .A4(n1147), .ZN(n1274) );
INV_X1 U959 ( .A(G898), .ZN(n1147) );
NAND3_X1 U960 ( .A1(G952), .A2(n1138), .A3(n1275), .ZN(n1256) );
XOR2_X1 U961 ( .A(n1048), .B(KEYINPUT28), .Z(n1275) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1048) );
NOR2_X1 U963 ( .A1(n1087), .A2(n1086), .ZN(n1088) );
INV_X1 U964 ( .A(n1251), .ZN(n1086) );
NAND2_X1 U965 ( .A1(G214), .A2(n1276), .ZN(n1251) );
XNOR2_X1 U966 ( .A(n1277), .B(n1205), .ZN(n1087) );
NAND2_X1 U967 ( .A1(G210), .A2(n1276), .ZN(n1205) );
NAND2_X1 U968 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
INV_X1 U969 ( .A(G237), .ZN(n1278) );
NAND2_X1 U970 ( .A1(n1280), .A2(n1279), .ZN(n1277) );
XOR2_X1 U971 ( .A(n1281), .B(n1282), .Z(n1280) );
XOR2_X1 U972 ( .A(n1283), .B(n1234), .Z(n1282) );
XOR2_X1 U973 ( .A(n1284), .B(n1285), .Z(n1234) );
XNOR2_X1 U974 ( .A(n1243), .B(n1286), .ZN(n1285) );
NOR2_X1 U975 ( .A1(n1150), .A2(KEYINPUT62), .ZN(n1286) );
AND2_X1 U976 ( .A1(n1287), .A2(n1288), .ZN(n1150) );
NAND2_X1 U977 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
XNOR2_X1 U978 ( .A(G113), .B(KEYINPUT6), .ZN(n1290) );
XNOR2_X1 U979 ( .A(G116), .B(G119), .ZN(n1289) );
NAND2_X1 U980 ( .A1(G113), .A2(n1291), .ZN(n1287) );
XNOR2_X1 U981 ( .A(n1292), .B(G116), .ZN(n1291) );
XNOR2_X1 U982 ( .A(n1148), .B(n1293), .ZN(n1284) );
INV_X1 U983 ( .A(n1294), .ZN(n1293) );
XNOR2_X1 U984 ( .A(n1295), .B(n1181), .ZN(n1148) );
INV_X1 U985 ( .A(n1296), .ZN(n1181) );
XNOR2_X1 U986 ( .A(n1297), .B(n1298), .ZN(n1295) );
NAND2_X1 U987 ( .A1(KEYINPUT34), .A2(n1299), .ZN(n1297) );
XNOR2_X1 U988 ( .A(G104), .B(n1300), .ZN(n1299) );
NAND2_X1 U989 ( .A1(KEYINPUT31), .A2(G107), .ZN(n1300) );
NAND2_X1 U990 ( .A1(KEYINPUT0), .A2(n1203), .ZN(n1283) );
NAND2_X1 U991 ( .A1(G224), .A2(n1138), .ZN(n1203) );
XOR2_X1 U992 ( .A(KEYINPUT7), .B(n1301), .Z(n1281) );
NOR2_X1 U993 ( .A1(KEYINPUT50), .A2(n1235), .ZN(n1301) );
XNOR2_X1 U994 ( .A(G125), .B(KEYINPUT30), .ZN(n1235) );
NOR2_X1 U995 ( .A1(n1242), .A2(n1241), .ZN(n1063) );
XOR2_X1 U996 ( .A(n1099), .B(n1172), .Z(n1241) );
INV_X1 U997 ( .A(G475), .ZN(n1172) );
NAND2_X1 U998 ( .A1(n1170), .A2(n1279), .ZN(n1099) );
XNOR2_X1 U999 ( .A(n1302), .B(n1303), .ZN(n1170) );
XOR2_X1 U1000 ( .A(n1304), .B(n1305), .Z(n1303) );
XOR2_X1 U1001 ( .A(n1306), .B(n1307), .Z(n1305) );
AND2_X1 U1002 ( .A1(G214), .A2(n1308), .ZN(n1307) );
NOR2_X1 U1003 ( .A1(KEYINPUT54), .A2(n1309), .ZN(n1306) );
XNOR2_X1 U1004 ( .A(G113), .B(G122), .ZN(n1309) );
XOR2_X1 U1005 ( .A(n1310), .B(n1311), .Z(n1302) );
XNOR2_X1 U1006 ( .A(n1312), .B(n1313), .ZN(n1311) );
NOR2_X1 U1007 ( .A1(KEYINPUT13), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U1008 ( .A(KEYINPUT38), .B(n1236), .ZN(n1314) );
INV_X1 U1009 ( .A(G104), .ZN(n1312) );
XNOR2_X1 U1010 ( .A(G131), .B(G143), .ZN(n1310) );
INV_X1 U1011 ( .A(n1259), .ZN(n1242) );
NOR2_X1 U1012 ( .A1(n1104), .A2(n1101), .ZN(n1259) );
AND2_X1 U1013 ( .A1(G478), .A2(n1315), .ZN(n1101) );
NAND2_X1 U1014 ( .A1(n1162), .A2(n1279), .ZN(n1315) );
NOR3_X1 U1015 ( .A1(G478), .A2(G902), .A3(n1316), .ZN(n1104) );
INV_X1 U1016 ( .A(n1162), .ZN(n1316) );
XNOR2_X1 U1017 ( .A(n1317), .B(n1318), .ZN(n1162) );
XOR2_X1 U1018 ( .A(n1319), .B(n1320), .Z(n1318) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1020 ( .A1(n1322), .A2(n1323), .ZN(n1319) );
NAND3_X1 U1021 ( .A1(KEYINPUT49), .A2(G143), .A3(n1324), .ZN(n1323) );
XNOR2_X1 U1022 ( .A(G134), .B(n1325), .ZN(n1324) );
NAND2_X1 U1023 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
NAND2_X1 U1024 ( .A1(KEYINPUT23), .A2(n1253), .ZN(n1327) );
NAND2_X1 U1025 ( .A1(KEYINPUT55), .A2(G128), .ZN(n1326) );
NAND2_X1 U1026 ( .A1(n1328), .A2(n1329), .ZN(n1322) );
NAND2_X1 U1027 ( .A1(KEYINPUT49), .A2(G143), .ZN(n1329) );
XNOR2_X1 U1028 ( .A(n1330), .B(n1250), .ZN(n1328) );
NAND2_X1 U1029 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
OR2_X1 U1030 ( .A1(n1253), .A2(KEYINPUT23), .ZN(n1332) );
OR2_X1 U1031 ( .A1(G128), .A2(KEYINPUT55), .ZN(n1331) );
XNOR2_X1 U1032 ( .A(G107), .B(n1333), .ZN(n1317) );
XNOR2_X1 U1033 ( .A(n1298), .B(G116), .ZN(n1333) );
INV_X1 U1034 ( .A(G122), .ZN(n1298) );
NOR2_X1 U1035 ( .A1(n1070), .A2(n1069), .ZN(n1068) );
INV_X1 U1036 ( .A(n1271), .ZN(n1069) );
NAND2_X1 U1037 ( .A1(G221), .A2(n1334), .ZN(n1271) );
INV_X1 U1038 ( .A(n1072), .ZN(n1070) );
XOR2_X1 U1039 ( .A(n1335), .B(n1199), .Z(n1072) );
INV_X1 U1040 ( .A(G469), .ZN(n1199) );
NAND2_X1 U1041 ( .A1(n1336), .A2(n1279), .ZN(n1335) );
XOR2_X1 U1042 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1043 ( .A(KEYINPUT61), .B(n1339), .ZN(n1338) );
INV_X1 U1044 ( .A(G110), .ZN(n1339) );
XOR2_X1 U1045 ( .A(n1340), .B(n1198), .Z(n1337) );
XNOR2_X1 U1046 ( .A(n1341), .B(n1342), .ZN(n1198) );
XNOR2_X1 U1047 ( .A(n1343), .B(n1129), .ZN(n1342) );
XNOR2_X1 U1048 ( .A(n1344), .B(n1345), .ZN(n1129) );
NOR2_X1 U1049 ( .A1(KEYINPUT37), .A2(n1253), .ZN(n1345) );
INV_X1 U1050 ( .A(G128), .ZN(n1253) );
XNOR2_X1 U1051 ( .A(G146), .B(G143), .ZN(n1344) );
INV_X1 U1052 ( .A(n1346), .ZN(n1343) );
XNOR2_X1 U1053 ( .A(n1296), .B(n1347), .ZN(n1341) );
XOR2_X1 U1054 ( .A(n1348), .B(n1349), .Z(n1347) );
NAND2_X1 U1055 ( .A1(G227), .A2(n1138), .ZN(n1349) );
NAND2_X1 U1056 ( .A1(KEYINPUT52), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1057 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
NAND2_X1 U1058 ( .A1(n1353), .A2(G104), .ZN(n1352) );
XOR2_X1 U1059 ( .A(KEYINPUT22), .B(n1354), .Z(n1351) );
NOR2_X1 U1060 ( .A1(G104), .A2(n1353), .ZN(n1354) );
XNOR2_X1 U1061 ( .A(KEYINPUT15), .B(G107), .ZN(n1353) );
NAND2_X1 U1062 ( .A1(KEYINPUT63), .A2(n1123), .ZN(n1340) );
NOR2_X1 U1063 ( .A1(n1261), .A2(n1262), .ZN(n1082) );
INV_X1 U1064 ( .A(n1098), .ZN(n1262) );
XOR2_X1 U1065 ( .A(n1355), .B(n1159), .Z(n1098) );
NAND2_X1 U1066 ( .A1(G217), .A2(n1334), .ZN(n1159) );
NAND2_X1 U1067 ( .A1(G234), .A2(n1356), .ZN(n1334) );
XNOR2_X1 U1068 ( .A(KEYINPUT11), .B(n1279), .ZN(n1356) );
NAND2_X1 U1069 ( .A1(n1357), .A2(n1157), .ZN(n1355) );
XNOR2_X1 U1070 ( .A(n1358), .B(n1359), .ZN(n1157) );
XOR2_X1 U1071 ( .A(n1360), .B(n1361), .Z(n1359) );
XOR2_X1 U1072 ( .A(G137), .B(n1362), .Z(n1361) );
NOR2_X1 U1073 ( .A1(KEYINPUT17), .A2(n1292), .ZN(n1362) );
AND2_X1 U1074 ( .A1(G221), .A2(n1321), .ZN(n1360) );
AND2_X1 U1075 ( .A1(G234), .A2(n1138), .ZN(n1321) );
INV_X1 U1076 ( .A(G953), .ZN(n1138) );
XNOR2_X1 U1077 ( .A(n1294), .B(n1304), .ZN(n1358) );
XNOR2_X1 U1078 ( .A(G125), .B(n1123), .ZN(n1304) );
INV_X1 U1079 ( .A(G140), .ZN(n1123) );
XOR2_X1 U1080 ( .A(G110), .B(n1363), .Z(n1294) );
XNOR2_X1 U1081 ( .A(KEYINPUT21), .B(n1279), .ZN(n1357) );
INV_X1 U1082 ( .A(n1263), .ZN(n1261) );
NOR2_X1 U1083 ( .A1(n1364), .A2(n1102), .ZN(n1263) );
NOR2_X1 U1084 ( .A1(n1103), .A2(G472), .ZN(n1102) );
AND2_X1 U1085 ( .A1(n1365), .A2(G472), .ZN(n1364) );
XOR2_X1 U1086 ( .A(n1103), .B(KEYINPUT26), .Z(n1365) );
NAND2_X1 U1087 ( .A1(n1366), .A2(n1279), .ZN(n1103) );
INV_X1 U1088 ( .A(G902), .ZN(n1279) );
XOR2_X1 U1089 ( .A(n1367), .B(n1368), .Z(n1366) );
XNOR2_X1 U1090 ( .A(n1186), .B(n1296), .ZN(n1368) );
XOR2_X1 U1091 ( .A(G101), .B(KEYINPUT47), .Z(n1296) );
XNOR2_X1 U1092 ( .A(n1369), .B(n1370), .ZN(n1186) );
XNOR2_X1 U1093 ( .A(n1346), .B(n1371), .ZN(n1370) );
XOR2_X1 U1094 ( .A(n1372), .B(n1363), .Z(n1371) );
XNOR2_X1 U1095 ( .A(n1236), .B(G128), .ZN(n1363) );
INV_X1 U1096 ( .A(G146), .ZN(n1236) );
NAND2_X1 U1097 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
NAND2_X1 U1098 ( .A1(G116), .A2(n1292), .ZN(n1374) );
XOR2_X1 U1099 ( .A(n1375), .B(KEYINPUT33), .Z(n1373) );
OR2_X1 U1100 ( .A1(n1292), .A2(G116), .ZN(n1375) );
INV_X1 U1101 ( .A(G119), .ZN(n1292) );
XOR2_X1 U1102 ( .A(n1132), .B(n1376), .Z(n1346) );
XNOR2_X1 U1103 ( .A(n1377), .B(KEYINPUT3), .ZN(n1376) );
NAND2_X1 U1104 ( .A1(KEYINPUT16), .A2(n1131), .ZN(n1377) );
INV_X1 U1105 ( .A(G131), .ZN(n1131) );
XNOR2_X1 U1106 ( .A(G137), .B(n1250), .ZN(n1132) );
INV_X1 U1107 ( .A(G134), .ZN(n1250) );
XNOR2_X1 U1108 ( .A(G113), .B(n1378), .ZN(n1369) );
XNOR2_X1 U1109 ( .A(KEYINPUT46), .B(n1243), .ZN(n1378) );
INV_X1 U1110 ( .A(G143), .ZN(n1243) );
XOR2_X1 U1111 ( .A(n1184), .B(KEYINPUT43), .Z(n1367) );
NAND2_X1 U1112 ( .A1(n1308), .A2(G210), .ZN(n1184) );
NOR2_X1 U1113 ( .A1(G953), .A2(G237), .ZN(n1308) );
endmodule


