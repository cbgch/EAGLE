//Key = 1110010000101110011001100000101010011001101111110101001111011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
n1449, n1450, n1451, n1452, n1453, n1454;

XOR2_X1 U796 ( .A(n1109), .B(n1110), .Z(G9) );
NOR2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(G75) );
NOR3_X1 U798 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NAND3_X1 U799 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1113) );
NAND2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND4_X1 U802 ( .A1(n1123), .A2(n1124), .A3(n1125), .A4(n1126), .ZN(n1122) );
OR2_X1 U803 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND3_X1 U804 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1121) );
NAND2_X1 U805 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NAND2_X1 U806 ( .A1(n1124), .A2(n1134), .ZN(n1133) );
NAND2_X1 U807 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND3_X1 U808 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
INV_X1 U809 ( .A(KEYINPUT55), .ZN(n1138) );
NAND2_X1 U810 ( .A1(n1125), .A2(n1140), .ZN(n1135) );
NAND2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NAND2_X1 U812 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U813 ( .A(n1145), .B(KEYINPUT53), .Z(n1141) );
NAND2_X1 U814 ( .A1(n1123), .A2(n1137), .ZN(n1132) );
NAND3_X1 U815 ( .A1(n1146), .A2(n1147), .A3(n1123), .ZN(n1137) );
NAND2_X1 U816 ( .A1(n1124), .A2(n1148), .ZN(n1147) );
NAND2_X1 U817 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NAND2_X1 U818 ( .A1(KEYINPUT55), .A2(n1139), .ZN(n1150) );
NAND2_X1 U819 ( .A1(n1125), .A2(n1151), .ZN(n1146) );
NAND2_X1 U820 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U822 ( .A(n1156), .B(KEYINPUT16), .Z(n1154) );
NOR3_X1 U823 ( .A1(n1157), .A2(G953), .A3(G952), .ZN(n1111) );
INV_X1 U824 ( .A(n1116), .ZN(n1157) );
NAND4_X1 U825 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1116) );
NOR4_X1 U826 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1161) );
XOR2_X1 U827 ( .A(KEYINPUT2), .B(n1166), .Z(n1165) );
NOR2_X1 U828 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NOR2_X1 U829 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U830 ( .A1(G902), .A2(n1171), .ZN(n1169) );
NOR3_X1 U831 ( .A1(n1155), .A2(n1143), .A3(n1172), .ZN(n1160) );
NAND2_X1 U832 ( .A1(n1173), .A2(n1174), .ZN(n1159) );
XNOR2_X1 U833 ( .A(n1175), .B(n1176), .ZN(n1158) );
NAND2_X1 U834 ( .A1(n1177), .A2(KEYINPUT51), .ZN(n1176) );
XNOR2_X1 U835 ( .A(G478), .B(KEYINPUT24), .ZN(n1177) );
XOR2_X1 U836 ( .A(n1178), .B(n1179), .Z(G72) );
NOR2_X1 U837 ( .A1(n1180), .A2(n1117), .ZN(n1179) );
NOR2_X1 U838 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND2_X1 U839 ( .A1(n1183), .A2(n1184), .ZN(n1178) );
NAND2_X1 U840 ( .A1(n1185), .A2(n1117), .ZN(n1184) );
XOR2_X1 U841 ( .A(n1114), .B(n1186), .Z(n1185) );
NAND3_X1 U842 ( .A1(G900), .A2(n1186), .A3(G953), .ZN(n1183) );
XNOR2_X1 U843 ( .A(n1187), .B(n1188), .ZN(n1186) );
XNOR2_X1 U844 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND2_X1 U845 ( .A1(KEYINPUT32), .A2(G140), .ZN(n1189) );
XOR2_X1 U846 ( .A(n1191), .B(n1192), .Z(n1187) );
XOR2_X1 U847 ( .A(KEYINPUT36), .B(G125), .Z(n1192) );
NAND2_X1 U848 ( .A1(n1193), .A2(n1194), .ZN(n1191) );
NAND2_X1 U849 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U850 ( .A(KEYINPUT60), .B(n1197), .Z(n1193) );
NOR2_X1 U851 ( .A1(n1196), .A2(n1195), .ZN(n1197) );
NAND2_X1 U852 ( .A1(n1198), .A2(n1199), .ZN(n1195) );
NAND2_X1 U853 ( .A1(KEYINPUT45), .A2(n1200), .ZN(n1199) );
OR3_X1 U854 ( .A1(n1201), .A2(G137), .A3(KEYINPUT45), .ZN(n1198) );
INV_X1 U855 ( .A(G134), .ZN(n1201) );
INV_X1 U856 ( .A(G131), .ZN(n1196) );
NAND2_X1 U857 ( .A1(n1202), .A2(n1203), .ZN(G69) );
NAND2_X1 U858 ( .A1(n1204), .A2(n1117), .ZN(n1203) );
XNOR2_X1 U859 ( .A(n1205), .B(n1115), .ZN(n1204) );
NAND2_X1 U860 ( .A1(n1206), .A2(G953), .ZN(n1202) );
NAND2_X1 U861 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U862 ( .A1(n1205), .A2(n1209), .ZN(n1208) );
NAND2_X1 U863 ( .A1(G224), .A2(n1210), .ZN(n1207) );
NAND2_X1 U864 ( .A1(G898), .A2(n1205), .ZN(n1210) );
NAND2_X1 U865 ( .A1(n1211), .A2(n1212), .ZN(n1205) );
NAND2_X1 U866 ( .A1(G953), .A2(n1213), .ZN(n1212) );
XNOR2_X1 U867 ( .A(n1214), .B(n1215), .ZN(n1211) );
NAND3_X1 U868 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1214) );
OR2_X1 U869 ( .A1(n1219), .A2(KEYINPUT44), .ZN(n1217) );
NAND3_X1 U870 ( .A1(n1219), .A2(n1220), .A3(KEYINPUT44), .ZN(n1216) );
NOR2_X1 U871 ( .A1(n1221), .A2(n1222), .ZN(G66) );
NOR2_X1 U872 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
XOR2_X1 U873 ( .A(n1225), .B(KEYINPUT57), .Z(n1224) );
NAND2_X1 U874 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
XOR2_X1 U875 ( .A(n1171), .B(n1228), .Z(n1227) );
XOR2_X1 U876 ( .A(KEYINPUT21), .B(KEYINPUT14), .Z(n1228) );
NOR2_X1 U877 ( .A1(n1226), .A2(n1171), .ZN(n1223) );
NOR2_X1 U878 ( .A1(n1229), .A2(n1170), .ZN(n1226) );
NOR2_X1 U879 ( .A1(n1221), .A2(n1230), .ZN(G63) );
XOR2_X1 U880 ( .A(n1231), .B(n1232), .Z(n1230) );
NAND2_X1 U881 ( .A1(KEYINPUT43), .A2(n1233), .ZN(n1231) );
NAND2_X1 U882 ( .A1(n1234), .A2(G478), .ZN(n1233) );
NOR2_X1 U883 ( .A1(n1221), .A2(n1235), .ZN(G60) );
XOR2_X1 U884 ( .A(n1236), .B(n1237), .Z(n1235) );
NOR2_X1 U885 ( .A1(n1238), .A2(KEYINPUT20), .ZN(n1236) );
AND2_X1 U886 ( .A1(G475), .A2(n1234), .ZN(n1238) );
XOR2_X1 U887 ( .A(G104), .B(n1239), .Z(G6) );
NOR2_X1 U888 ( .A1(n1221), .A2(n1240), .ZN(G57) );
XOR2_X1 U889 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U890 ( .A(n1243), .B(n1244), .Z(n1241) );
NOR2_X1 U891 ( .A1(KEYINPUT41), .A2(n1245), .ZN(n1244) );
XOR2_X1 U892 ( .A(n1246), .B(KEYINPUT49), .Z(n1245) );
NAND2_X1 U893 ( .A1(n1234), .A2(G472), .ZN(n1243) );
NOR3_X1 U894 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(G54) );
AND2_X1 U895 ( .A1(KEYINPUT46), .A2(n1221), .ZN(n1249) );
NOR3_X1 U896 ( .A1(KEYINPUT46), .A2(G953), .A3(G952), .ZN(n1248) );
XOR2_X1 U897 ( .A(n1250), .B(n1251), .Z(n1247) );
XOR2_X1 U898 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U899 ( .A(n1254), .B(n1255), .Z(n1250) );
XOR2_X1 U900 ( .A(n1256), .B(G110), .Z(n1255) );
NAND2_X1 U901 ( .A1(KEYINPUT18), .A2(n1257), .ZN(n1256) );
NAND2_X1 U902 ( .A1(n1234), .A2(G469), .ZN(n1254) );
NOR2_X1 U903 ( .A1(n1221), .A2(n1258), .ZN(G51) );
XOR2_X1 U904 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U905 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U906 ( .A(n1263), .B(n1264), .Z(n1259) );
XOR2_X1 U907 ( .A(n1265), .B(n1266), .Z(n1264) );
NOR2_X1 U908 ( .A1(KEYINPUT27), .A2(n1267), .ZN(n1266) );
NAND2_X1 U909 ( .A1(n1234), .A2(n1173), .ZN(n1265) );
INV_X1 U910 ( .A(n1229), .ZN(n1234) );
NAND2_X1 U911 ( .A1(G902), .A2(n1268), .ZN(n1229) );
OR2_X1 U912 ( .A1(n1115), .A2(n1114), .ZN(n1268) );
NAND4_X1 U913 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1114) );
AND4_X1 U914 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1272) );
NAND2_X1 U915 ( .A1(n1277), .A2(n1278), .ZN(n1271) );
NAND2_X1 U916 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
NAND4_X1 U917 ( .A1(n1128), .A2(n1124), .A3(n1281), .A4(n1282), .ZN(n1280) );
XOR2_X1 U918 ( .A(KEYINPUT30), .B(n1283), .Z(n1279) );
NAND4_X1 U919 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1115) );
AND4_X1 U920 ( .A1(n1288), .A2(n1110), .A3(n1289), .A4(n1290), .ZN(n1287) );
NAND2_X1 U921 ( .A1(n1139), .A2(n1291), .ZN(n1110) );
NOR3_X1 U922 ( .A1(n1239), .A2(n1292), .A3(n1293), .ZN(n1286) );
NOR3_X1 U923 ( .A1(n1294), .A2(n1295), .A3(n1145), .ZN(n1293) );
INV_X1 U924 ( .A(KEYINPUT38), .ZN(n1294) );
NOR2_X1 U925 ( .A1(KEYINPUT38), .A2(n1296), .ZN(n1292) );
AND2_X1 U926 ( .A1(n1281), .A2(n1291), .ZN(n1239) );
AND3_X1 U927 ( .A1(n1129), .A2(n1131), .A3(n1297), .ZN(n1291) );
NAND2_X1 U928 ( .A1(KEYINPUT0), .A2(n1298), .ZN(n1263) );
NOR2_X1 U929 ( .A1(n1117), .A2(G952), .ZN(n1221) );
XOR2_X1 U930 ( .A(n1299), .B(n1269), .Z(G48) );
NAND3_X1 U931 ( .A1(n1281), .A2(n1277), .A3(n1300), .ZN(n1269) );
NAND2_X1 U932 ( .A1(n1301), .A2(n1302), .ZN(G45) );
NAND2_X1 U933 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U934 ( .A1(G143), .A2(n1305), .ZN(n1301) );
NAND2_X1 U935 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
OR2_X1 U936 ( .A1(n1270), .A2(KEYINPUT5), .ZN(n1307) );
NAND2_X1 U937 ( .A1(KEYINPUT5), .A2(n1308), .ZN(n1306) );
INV_X1 U938 ( .A(n1303), .ZN(n1308) );
NOR2_X1 U939 ( .A1(KEYINPUT58), .A2(n1270), .ZN(n1303) );
NAND4_X1 U940 ( .A1(n1309), .A2(n1277), .A3(n1310), .A4(n1163), .ZN(n1270) );
XNOR2_X1 U941 ( .A(G140), .B(n1276), .ZN(G42) );
NAND4_X1 U942 ( .A1(n1311), .A2(n1282), .A3(n1281), .A4(n1312), .ZN(n1276) );
NOR2_X1 U943 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XNOR2_X1 U944 ( .A(G137), .B(n1275), .ZN(G39) );
NAND3_X1 U945 ( .A1(n1123), .A2(n1125), .A3(n1300), .ZN(n1275) );
NAND2_X1 U946 ( .A1(n1315), .A2(n1316), .ZN(G36) );
NAND2_X1 U947 ( .A1(G134), .A2(n1274), .ZN(n1316) );
XOR2_X1 U948 ( .A(KEYINPUT28), .B(n1317), .Z(n1315) );
NOR2_X1 U949 ( .A1(G134), .A2(n1274), .ZN(n1317) );
NAND3_X1 U950 ( .A1(n1309), .A2(n1139), .A3(n1123), .ZN(n1274) );
XOR2_X1 U951 ( .A(n1273), .B(n1318), .Z(G33) );
NAND2_X1 U952 ( .A1(KEYINPUT13), .A2(G131), .ZN(n1318) );
NAND3_X1 U953 ( .A1(n1309), .A2(n1281), .A3(n1123), .ZN(n1273) );
INV_X1 U954 ( .A(n1314), .ZN(n1123) );
NAND2_X1 U955 ( .A1(n1144), .A2(n1319), .ZN(n1314) );
AND3_X1 U956 ( .A1(n1311), .A2(n1282), .A3(n1127), .ZN(n1309) );
INV_X1 U957 ( .A(n1152), .ZN(n1311) );
XOR2_X1 U958 ( .A(n1320), .B(n1321), .Z(G30) );
NAND2_X1 U959 ( .A1(n1283), .A2(n1277), .ZN(n1321) );
AND2_X1 U960 ( .A1(n1300), .A2(n1139), .ZN(n1283) );
NOR4_X1 U961 ( .A1(n1322), .A2(n1152), .A3(n1129), .A4(n1323), .ZN(n1300) );
XNOR2_X1 U962 ( .A(G101), .B(n1284), .ZN(G3) );
NAND3_X1 U963 ( .A1(n1297), .A2(n1125), .A3(n1127), .ZN(n1284) );
XOR2_X1 U964 ( .A(n1324), .B(n1325), .Z(G27) );
NAND4_X1 U965 ( .A1(n1281), .A2(n1277), .A3(n1124), .A4(n1326), .ZN(n1325) );
NOR2_X1 U966 ( .A1(n1313), .A2(n1327), .ZN(n1326) );
XOR2_X1 U967 ( .A(KEYINPUT31), .B(n1323), .Z(n1327) );
INV_X1 U968 ( .A(n1282), .ZN(n1323) );
NAND2_X1 U969 ( .A1(n1328), .A2(n1329), .ZN(n1282) );
NAND4_X1 U970 ( .A1(G953), .A2(G902), .A3(n1330), .A4(n1182), .ZN(n1329) );
INV_X1 U971 ( .A(G900), .ZN(n1182) );
XOR2_X1 U972 ( .A(KEYINPUT62), .B(n1119), .Z(n1328) );
INV_X1 U973 ( .A(n1331), .ZN(n1119) );
INV_X1 U974 ( .A(n1128), .ZN(n1313) );
XNOR2_X1 U975 ( .A(n1296), .B(n1332), .ZN(G24) );
NOR2_X1 U976 ( .A1(KEYINPUT23), .A2(n1333), .ZN(n1332) );
NAND2_X1 U977 ( .A1(n1295), .A2(n1277), .ZN(n1296) );
AND4_X1 U978 ( .A1(n1129), .A2(n1131), .A3(n1124), .A4(n1334), .ZN(n1295) );
NOR3_X1 U979 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
INV_X1 U980 ( .A(n1338), .ZN(n1131) );
XNOR2_X1 U981 ( .A(G119), .B(n1288), .ZN(G21) );
NAND4_X1 U982 ( .A1(n1164), .A2(n1339), .A3(n1125), .A4(n1340), .ZN(n1288) );
NOR3_X1 U983 ( .A1(n1341), .A2(n1145), .A3(n1322), .ZN(n1340) );
XNOR2_X1 U984 ( .A(n1285), .B(n1342), .ZN(G18) );
NOR2_X1 U985 ( .A1(KEYINPUT9), .A2(n1343), .ZN(n1342) );
NAND2_X1 U986 ( .A1(n1344), .A2(n1139), .ZN(n1285) );
AND2_X1 U987 ( .A1(n1345), .A2(n1310), .ZN(n1139) );
INV_X1 U988 ( .A(n1335), .ZN(n1310) );
XOR2_X1 U989 ( .A(n1346), .B(n1163), .Z(n1345) );
XOR2_X1 U990 ( .A(n1347), .B(n1290), .Z(G15) );
NAND2_X1 U991 ( .A1(n1344), .A2(n1281), .ZN(n1290) );
AND4_X1 U992 ( .A1(n1127), .A2(n1124), .A3(n1277), .A4(n1339), .ZN(n1344) );
INV_X1 U993 ( .A(n1341), .ZN(n1124) );
NAND2_X1 U994 ( .A1(n1348), .A2(n1156), .ZN(n1341) );
NOR2_X1 U995 ( .A1(n1338), .A2(n1129), .ZN(n1127) );
XOR2_X1 U996 ( .A(n1349), .B(n1289), .Z(G12) );
NAND3_X1 U997 ( .A1(n1297), .A2(n1125), .A3(n1128), .ZN(n1289) );
NOR2_X1 U998 ( .A1(n1322), .A2(n1164), .ZN(n1128) );
INV_X1 U999 ( .A(n1129), .ZN(n1164) );
XOR2_X1 U1000 ( .A(n1350), .B(G472), .Z(n1129) );
NAND3_X1 U1001 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1350) );
NAND2_X1 U1002 ( .A1(n1354), .A2(n1355), .ZN(n1352) );
INV_X1 U1003 ( .A(KEYINPUT34), .ZN(n1355) );
XOR2_X1 U1004 ( .A(n1242), .B(n1356), .Z(n1354) );
NAND3_X1 U1005 ( .A1(n1356), .A2(n1242), .A3(KEYINPUT34), .ZN(n1351) );
XNOR2_X1 U1006 ( .A(n1357), .B(n1358), .ZN(n1242) );
XOR2_X1 U1007 ( .A(n1347), .B(n1359), .Z(n1358) );
XNOR2_X1 U1008 ( .A(n1261), .B(n1360), .ZN(n1357) );
INV_X1 U1009 ( .A(n1246), .ZN(n1356) );
XOR2_X1 U1010 ( .A(n1361), .B(G101), .Z(n1246) );
NAND2_X1 U1011 ( .A1(G210), .A2(n1362), .ZN(n1361) );
XNOR2_X1 U1012 ( .A(n1338), .B(KEYINPUT7), .ZN(n1322) );
NAND2_X1 U1013 ( .A1(n1363), .A2(n1364), .ZN(n1338) );
NAND2_X1 U1014 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
OR2_X1 U1015 ( .A1(n1171), .A2(G902), .ZN(n1366) );
XNOR2_X1 U1016 ( .A(n1167), .B(KEYINPUT4), .ZN(n1363) );
NOR3_X1 U1017 ( .A1(n1365), .A2(G902), .A3(n1171), .ZN(n1167) );
XNOR2_X1 U1018 ( .A(n1367), .B(n1368), .ZN(n1171) );
XOR2_X1 U1019 ( .A(n1369), .B(n1370), .Z(n1368) );
XOR2_X1 U1020 ( .A(n1371), .B(n1372), .Z(n1370) );
NAND2_X1 U1021 ( .A1(KEYINPUT59), .A2(n1373), .ZN(n1371) );
XNOR2_X1 U1022 ( .A(G137), .B(n1374), .ZN(n1373) );
NAND2_X1 U1023 ( .A1(G221), .A2(n1375), .ZN(n1374) );
XOR2_X1 U1024 ( .A(n1376), .B(n1377), .Z(n1367) );
XOR2_X1 U1025 ( .A(KEYINPUT15), .B(G119), .Z(n1377) );
NAND2_X1 U1026 ( .A1(KEYINPUT35), .A2(n1378), .ZN(n1376) );
XOR2_X1 U1027 ( .A(KEYINPUT17), .B(G110), .Z(n1378) );
INV_X1 U1028 ( .A(n1170), .ZN(n1365) );
NAND2_X1 U1029 ( .A1(G217), .A2(n1379), .ZN(n1170) );
NAND2_X1 U1030 ( .A1(n1380), .A2(n1381), .ZN(n1125) );
NAND3_X1 U1031 ( .A1(n1382), .A2(n1337), .A3(n1346), .ZN(n1381) );
INV_X1 U1032 ( .A(KEYINPUT6), .ZN(n1346) );
NAND2_X1 U1033 ( .A1(KEYINPUT6), .A2(n1281), .ZN(n1380) );
INV_X1 U1034 ( .A(n1149), .ZN(n1281) );
NAND2_X1 U1035 ( .A1(n1382), .A2(n1163), .ZN(n1149) );
INV_X1 U1036 ( .A(n1337), .ZN(n1163) );
XOR2_X1 U1037 ( .A(n1383), .B(G475), .Z(n1337) );
NAND2_X1 U1038 ( .A1(n1237), .A2(n1353), .ZN(n1383) );
XNOR2_X1 U1039 ( .A(n1384), .B(n1385), .ZN(n1237) );
XOR2_X1 U1040 ( .A(n1386), .B(n1387), .Z(n1385) );
XOR2_X1 U1041 ( .A(G131), .B(G104), .Z(n1387) );
XOR2_X1 U1042 ( .A(G146), .B(G143), .Z(n1386) );
XOR2_X1 U1043 ( .A(n1388), .B(n1389), .Z(n1384) );
AND2_X1 U1044 ( .A1(n1362), .A2(G214), .ZN(n1389) );
NOR2_X1 U1045 ( .A1(G953), .A2(G237), .ZN(n1362) );
XOR2_X1 U1046 ( .A(n1390), .B(n1391), .Z(n1388) );
NOR2_X1 U1047 ( .A1(KEYINPUT63), .A2(n1369), .ZN(n1391) );
XOR2_X1 U1048 ( .A(n1324), .B(G140), .Z(n1369) );
NAND2_X1 U1049 ( .A1(n1392), .A2(n1393), .ZN(n1390) );
NAND2_X1 U1050 ( .A1(n1394), .A2(n1347), .ZN(n1393) );
NAND2_X1 U1051 ( .A1(KEYINPUT42), .A2(n1395), .ZN(n1394) );
NAND2_X1 U1052 ( .A1(n1333), .A2(n1396), .ZN(n1395) );
NAND2_X1 U1053 ( .A1(G122), .A2(n1397), .ZN(n1392) );
NAND2_X1 U1054 ( .A1(n1396), .A2(n1398), .ZN(n1397) );
NAND2_X1 U1055 ( .A1(G113), .A2(KEYINPUT42), .ZN(n1398) );
INV_X1 U1056 ( .A(KEYINPUT8), .ZN(n1396) );
XOR2_X1 U1057 ( .A(n1335), .B(KEYINPUT3), .Z(n1382) );
NAND3_X1 U1058 ( .A1(n1399), .A2(n1400), .A3(n1401), .ZN(n1335) );
NAND2_X1 U1059 ( .A1(KEYINPUT48), .A2(n1175), .ZN(n1401) );
OR4_X1 U1060 ( .A1(n1175), .A2(KEYINPUT48), .A3(n1402), .A4(G478), .ZN(n1400) );
NAND2_X1 U1061 ( .A1(G478), .A2(n1403), .ZN(n1399) );
OR2_X1 U1062 ( .A1(n1402), .A2(n1175), .ZN(n1403) );
NOR2_X1 U1063 ( .A1(n1232), .A2(G902), .ZN(n1175) );
XNOR2_X1 U1064 ( .A(n1404), .B(n1405), .ZN(n1232) );
XOR2_X1 U1065 ( .A(n1406), .B(n1407), .Z(n1405) );
NAND2_X1 U1066 ( .A1(KEYINPUT22), .A2(n1343), .ZN(n1407) );
NAND2_X1 U1067 ( .A1(G217), .A2(n1375), .ZN(n1406) );
AND2_X1 U1068 ( .A1(G234), .A2(n1117), .ZN(n1375) );
XOR2_X1 U1069 ( .A(n1408), .B(n1409), .Z(n1404) );
XOR2_X1 U1070 ( .A(G122), .B(G107), .Z(n1409) );
NAND2_X1 U1071 ( .A1(n1410), .A2(n1411), .ZN(n1408) );
NAND2_X1 U1072 ( .A1(G134), .A2(n1412), .ZN(n1411) );
XOR2_X1 U1073 ( .A(KEYINPUT10), .B(n1413), .Z(n1410) );
NOR2_X1 U1074 ( .A1(G134), .A2(n1412), .ZN(n1413) );
INV_X1 U1075 ( .A(KEYINPUT39), .ZN(n1402) );
NOR3_X1 U1076 ( .A1(n1152), .A2(n1336), .A3(n1145), .ZN(n1297) );
INV_X1 U1077 ( .A(n1277), .ZN(n1145) );
NOR2_X1 U1078 ( .A1(n1143), .A2(n1144), .ZN(n1277) );
NOR2_X1 U1079 ( .A1(n1172), .A2(n1414), .ZN(n1144) );
AND2_X1 U1080 ( .A1(n1415), .A2(n1174), .ZN(n1414) );
XOR2_X1 U1081 ( .A(KEYINPUT33), .B(n1173), .Z(n1415) );
NOR2_X1 U1082 ( .A1(n1174), .A2(n1173), .ZN(n1172) );
AND2_X1 U1083 ( .A1(G210), .A2(n1416), .ZN(n1173) );
NAND2_X1 U1084 ( .A1(n1417), .A2(n1418), .ZN(n1174) );
XOR2_X1 U1085 ( .A(KEYINPUT47), .B(G902), .Z(n1418) );
XOR2_X1 U1086 ( .A(n1419), .B(n1420), .Z(n1417) );
XNOR2_X1 U1087 ( .A(n1298), .B(n1421), .ZN(n1420) );
NAND2_X1 U1088 ( .A1(KEYINPUT12), .A2(n1262), .ZN(n1421) );
XOR2_X1 U1089 ( .A(n1324), .B(KEYINPUT29), .Z(n1262) );
INV_X1 U1090 ( .A(G125), .ZN(n1324) );
NOR2_X1 U1091 ( .A1(n1209), .A2(G953), .ZN(n1298) );
INV_X1 U1092 ( .A(G224), .ZN(n1209) );
XOR2_X1 U1093 ( .A(n1261), .B(n1267), .Z(n1419) );
XNOR2_X1 U1094 ( .A(n1422), .B(n1215), .ZN(n1267) );
XNOR2_X1 U1095 ( .A(n1333), .B(n1423), .ZN(n1215) );
NOR2_X1 U1096 ( .A1(G110), .A2(KEYINPUT25), .ZN(n1423) );
INV_X1 U1097 ( .A(G122), .ZN(n1333) );
NAND2_X1 U1098 ( .A1(n1218), .A2(n1424), .ZN(n1422) );
NAND2_X1 U1099 ( .A1(n1219), .A2(n1220), .ZN(n1424) );
OR2_X1 U1100 ( .A1(n1220), .A2(n1219), .ZN(n1218) );
AND2_X1 U1101 ( .A1(n1425), .A2(n1426), .ZN(n1219) );
XNOR2_X1 U1102 ( .A(n1347), .B(n1427), .ZN(n1220) );
NOR2_X1 U1103 ( .A1(KEYINPUT26), .A2(n1359), .ZN(n1427) );
XOR2_X1 U1104 ( .A(n1343), .B(G119), .Z(n1359) );
INV_X1 U1105 ( .A(G116), .ZN(n1343) );
INV_X1 U1106 ( .A(G113), .ZN(n1347) );
XOR2_X1 U1107 ( .A(n1428), .B(n1372), .Z(n1261) );
XOR2_X1 U1108 ( .A(G128), .B(G146), .Z(n1372) );
NAND2_X1 U1109 ( .A1(KEYINPUT40), .A2(n1304), .ZN(n1428) );
INV_X1 U1110 ( .A(n1319), .ZN(n1143) );
NAND2_X1 U1111 ( .A1(G214), .A2(n1416), .ZN(n1319) );
NAND2_X1 U1112 ( .A1(n1429), .A2(n1353), .ZN(n1416) );
INV_X1 U1113 ( .A(G237), .ZN(n1429) );
INV_X1 U1114 ( .A(n1339), .ZN(n1336) );
NAND2_X1 U1115 ( .A1(n1331), .A2(n1430), .ZN(n1339) );
NAND4_X1 U1116 ( .A1(G953), .A2(G902), .A3(n1330), .A4(n1213), .ZN(n1430) );
INV_X1 U1117 ( .A(G898), .ZN(n1213) );
NAND3_X1 U1118 ( .A1(n1330), .A2(n1117), .A3(G952), .ZN(n1331) );
INV_X1 U1119 ( .A(G953), .ZN(n1117) );
NAND2_X1 U1120 ( .A1(G237), .A2(G234), .ZN(n1330) );
NAND2_X1 U1121 ( .A1(n1348), .A2(n1431), .ZN(n1152) );
XOR2_X1 U1122 ( .A(KEYINPUT52), .B(n1432), .Z(n1431) );
INV_X1 U1123 ( .A(n1156), .ZN(n1432) );
XNOR2_X1 U1124 ( .A(n1162), .B(KEYINPUT11), .ZN(n1156) );
XNOR2_X1 U1125 ( .A(n1433), .B(G469), .ZN(n1162) );
NAND2_X1 U1126 ( .A1(n1434), .A2(n1353), .ZN(n1433) );
NAND2_X1 U1127 ( .A1(n1435), .A2(n1436), .ZN(n1434) );
NAND2_X1 U1128 ( .A1(n1437), .A2(n1438), .ZN(n1436) );
XOR2_X1 U1129 ( .A(n1439), .B(n1440), .Z(n1437) );
XOR2_X1 U1130 ( .A(n1441), .B(KEYINPUT61), .Z(n1435) );
NAND2_X1 U1131 ( .A1(n1442), .A2(n1443), .ZN(n1441) );
INV_X1 U1132 ( .A(n1438), .ZN(n1443) );
XOR2_X1 U1133 ( .A(n1257), .B(n1253), .Z(n1438) );
XNOR2_X1 U1134 ( .A(n1360), .B(n1190), .ZN(n1253) );
XOR2_X1 U1135 ( .A(n1412), .B(n1444), .Z(n1190) );
XNOR2_X1 U1136 ( .A(n1445), .B(KEYINPUT1), .ZN(n1444) );
NAND2_X1 U1137 ( .A1(KEYINPUT54), .A2(n1299), .ZN(n1445) );
INV_X1 U1138 ( .A(G146), .ZN(n1299) );
XOR2_X1 U1139 ( .A(n1320), .B(n1304), .Z(n1412) );
INV_X1 U1140 ( .A(G143), .ZN(n1304) );
INV_X1 U1141 ( .A(G128), .ZN(n1320) );
XOR2_X1 U1142 ( .A(G131), .B(n1200), .Z(n1360) );
XNOR2_X1 U1143 ( .A(G137), .B(G134), .ZN(n1200) );
NAND3_X1 U1144 ( .A1(n1446), .A2(n1447), .A3(n1426), .ZN(n1257) );
NAND3_X1 U1145 ( .A1(G104), .A2(n1109), .A3(G101), .ZN(n1426) );
OR2_X1 U1146 ( .A1(n1425), .A2(KEYINPUT37), .ZN(n1447) );
AND2_X1 U1147 ( .A1(n1448), .A2(n1449), .ZN(n1425) );
OR3_X1 U1148 ( .A1(G101), .A2(G104), .A3(G107), .ZN(n1449) );
NAND2_X1 U1149 ( .A1(n1450), .A2(G107), .ZN(n1448) );
XOR2_X1 U1150 ( .A(G104), .B(G101), .Z(n1450) );
NAND2_X1 U1151 ( .A1(n1451), .A2(KEYINPUT37), .ZN(n1446) );
XOR2_X1 U1152 ( .A(G101), .B(n1452), .Z(n1451) );
NOR2_X1 U1153 ( .A1(G104), .A2(n1109), .ZN(n1452) );
INV_X1 U1154 ( .A(G107), .ZN(n1109) );
XOR2_X1 U1155 ( .A(n1440), .B(n1252), .Z(n1442) );
INV_X1 U1156 ( .A(n1439), .ZN(n1252) );
XNOR2_X1 U1157 ( .A(G140), .B(n1453), .ZN(n1439) );
NOR2_X1 U1158 ( .A1(G953), .A2(n1181), .ZN(n1453) );
INV_X1 U1159 ( .A(G227), .ZN(n1181) );
NOR2_X1 U1160 ( .A1(KEYINPUT50), .A2(n1454), .ZN(n1440) );
XOR2_X1 U1161 ( .A(n1349), .B(KEYINPUT56), .Z(n1454) );
XNOR2_X1 U1162 ( .A(n1155), .B(KEYINPUT19), .ZN(n1348) );
AND2_X1 U1163 ( .A1(G221), .A2(n1379), .ZN(n1155) );
NAND2_X1 U1164 ( .A1(G234), .A2(n1353), .ZN(n1379) );
INV_X1 U1165 ( .A(G902), .ZN(n1353) );
INV_X1 U1166 ( .A(G110), .ZN(n1349) );
endmodule


