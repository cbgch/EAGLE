//Key = 1101110100111000001110110000100101010110101111101010110000001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
n1463, n1464, n1465, n1466, n1467, n1468;

XOR2_X1 U814 ( .A(G107), .B(n1133), .Z(G9) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U816 ( .A1(n1136), .A2(n1137), .ZN(G75) );
NOR4_X1 U817 ( .A1(G953), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NOR2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
NOR3_X1 U820 ( .A1(n1145), .A2(n1146), .A3(n1147), .ZN(n1144) );
NOR3_X1 U821 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NOR3_X1 U822 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR3_X1 U823 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
NOR2_X1 U824 ( .A1(n1157), .A2(n1158), .ZN(n1152) );
AND3_X1 U825 ( .A1(KEYINPUT52), .A2(n1159), .A3(n1157), .ZN(n1149) );
NOR2_X1 U826 ( .A1(n1160), .A2(n1161), .ZN(n1146) );
NOR3_X1 U827 ( .A1(n1162), .A2(KEYINPUT52), .A3(n1163), .ZN(n1161) );
NOR4_X1 U828 ( .A1(n1154), .A2(n1164), .A3(n1151), .A4(n1162), .ZN(n1143) );
INV_X1 U829 ( .A(n1157), .ZN(n1162) );
NOR3_X1 U830 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1164) );
NOR2_X1 U831 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NOR2_X1 U832 ( .A1(n1170), .A2(n1171), .ZN(n1168) );
NOR2_X1 U833 ( .A1(n1172), .A2(n1135), .ZN(n1171) );
NOR2_X1 U834 ( .A1(n1173), .A2(n1148), .ZN(n1170) );
INV_X1 U835 ( .A(n1160), .ZN(n1148) );
NOR2_X1 U836 ( .A1(n1172), .A2(n1174), .ZN(n1173) );
NOR4_X1 U837 ( .A1(n1175), .A2(n1145), .A3(n1176), .A4(n1174), .ZN(n1166) );
INV_X1 U838 ( .A(KEYINPUT1), .ZN(n1174) );
AND2_X1 U839 ( .A1(n1177), .A2(n1160), .ZN(n1165) );
NOR3_X1 U840 ( .A1(n1138), .A2(G953), .A3(G952), .ZN(n1136) );
AND4_X1 U841 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1138) );
NOR4_X1 U842 ( .A1(n1182), .A2(n1154), .A3(n1183), .A4(n1184), .ZN(n1181) );
XOR2_X1 U843 ( .A(n1185), .B(n1186), .Z(n1184) );
XOR2_X1 U844 ( .A(KEYINPUT60), .B(G472), .Z(n1186) );
NOR2_X1 U845 ( .A1(n1187), .A2(KEYINPUT24), .ZN(n1185) );
NOR3_X1 U846 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1180) );
NOR2_X1 U847 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U848 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U849 ( .A(KEYINPUT22), .B(KEYINPUT21), .Z(n1194) );
NOR2_X1 U850 ( .A1(n1195), .A2(n1193), .ZN(n1189) );
XNOR2_X1 U851 ( .A(n1196), .B(KEYINPUT49), .ZN(n1193) );
INV_X1 U852 ( .A(n1191), .ZN(n1195) );
XNOR2_X1 U853 ( .A(KEYINPUT45), .B(n1151), .ZN(n1188) );
XNOR2_X1 U854 ( .A(n1197), .B(n1198), .ZN(n1179) );
NAND2_X1 U855 ( .A1(KEYINPUT7), .A2(n1199), .ZN(n1197) );
XOR2_X1 U856 ( .A(n1200), .B(KEYINPUT5), .Z(n1178) );
NAND2_X1 U857 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
XOR2_X1 U858 ( .A(n1203), .B(n1204), .Z(G72) );
NOR2_X1 U859 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
AND2_X1 U860 ( .A1(G227), .A2(G900), .ZN(n1205) );
NAND2_X1 U861 ( .A1(n1207), .A2(n1208), .ZN(n1203) );
NAND3_X1 U862 ( .A1(n1209), .A2(n1210), .A3(n1211), .ZN(n1208) );
INV_X1 U863 ( .A(n1212), .ZN(n1210) );
OR2_X1 U864 ( .A1(n1211), .A2(n1209), .ZN(n1207) );
XNOR2_X1 U865 ( .A(n1213), .B(n1214), .ZN(n1209) );
XOR2_X1 U866 ( .A(n1215), .B(n1216), .Z(n1214) );
XOR2_X1 U867 ( .A(n1217), .B(KEYINPUT3), .Z(n1216) );
NAND2_X1 U868 ( .A1(n1218), .A2(n1219), .ZN(n1215) );
XNOR2_X1 U869 ( .A(n1220), .B(KEYINPUT30), .ZN(n1218) );
XOR2_X1 U870 ( .A(n1221), .B(n1222), .Z(n1213) );
NAND2_X1 U871 ( .A1(n1206), .A2(n1223), .ZN(n1211) );
NAND2_X1 U872 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND2_X1 U873 ( .A1(n1226), .A2(n1227), .ZN(G69) );
NAND2_X1 U874 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
XNOR2_X1 U875 ( .A(KEYINPUT8), .B(n1230), .ZN(n1229) );
XOR2_X1 U876 ( .A(n1231), .B(n1232), .Z(n1228) );
NAND2_X1 U877 ( .A1(n1233), .A2(n1234), .ZN(n1226) );
XNOR2_X1 U878 ( .A(n1232), .B(n1231), .ZN(n1234) );
NAND2_X1 U879 ( .A1(n1206), .A2(n1235), .ZN(n1231) );
NOR2_X1 U880 ( .A1(n1236), .A2(n1237), .ZN(n1232) );
XOR2_X1 U881 ( .A(n1238), .B(n1239), .Z(n1236) );
XOR2_X1 U882 ( .A(n1240), .B(n1241), .Z(n1238) );
NOR2_X1 U883 ( .A1(KEYINPUT29), .A2(n1242), .ZN(n1241) );
XOR2_X1 U884 ( .A(n1230), .B(KEYINPUT26), .Z(n1233) );
NAND2_X1 U885 ( .A1(G953), .A2(n1243), .ZN(n1230) );
NAND2_X1 U886 ( .A1(G898), .A2(G224), .ZN(n1243) );
NOR2_X1 U887 ( .A1(n1244), .A2(n1245), .ZN(G66) );
NOR2_X1 U888 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
XOR2_X1 U889 ( .A(n1248), .B(n1249), .Z(n1247) );
AND2_X1 U890 ( .A1(n1250), .A2(KEYINPUT42), .ZN(n1249) );
OR2_X1 U891 ( .A1(n1251), .A2(n1196), .ZN(n1248) );
NOR2_X1 U892 ( .A1(KEYINPUT42), .A2(n1250), .ZN(n1246) );
NOR2_X1 U893 ( .A1(n1252), .A2(n1253), .ZN(G63) );
XOR2_X1 U894 ( .A(KEYINPUT14), .B(n1244), .Z(n1253) );
XOR2_X1 U895 ( .A(n1254), .B(n1255), .Z(n1252) );
NAND2_X1 U896 ( .A1(n1256), .A2(G478), .ZN(n1254) );
NOR2_X1 U897 ( .A1(n1244), .A2(n1257), .ZN(G60) );
XOR2_X1 U898 ( .A(n1258), .B(n1259), .Z(n1257) );
NAND2_X1 U899 ( .A1(n1256), .A2(G475), .ZN(n1259) );
XOR2_X1 U900 ( .A(n1260), .B(n1261), .Z(G6) );
NOR2_X1 U901 ( .A1(n1244), .A2(n1262), .ZN(G57) );
XOR2_X1 U902 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U903 ( .A(n1265), .B(n1266), .Z(n1264) );
XOR2_X1 U904 ( .A(n1267), .B(n1268), .Z(n1263) );
NOR2_X1 U905 ( .A1(KEYINPUT56), .A2(n1269), .ZN(n1268) );
XOR2_X1 U906 ( .A(n1270), .B(n1271), .Z(n1269) );
NOR2_X1 U907 ( .A1(KEYINPUT16), .A2(n1272), .ZN(n1271) );
NAND2_X1 U908 ( .A1(n1256), .A2(G472), .ZN(n1267) );
NOR2_X1 U909 ( .A1(n1244), .A2(n1273), .ZN(G54) );
NOR2_X1 U910 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U911 ( .A(KEYINPUT55), .B(n1276), .Z(n1275) );
NOR2_X1 U912 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
AND2_X1 U913 ( .A1(n1278), .A2(n1277), .ZN(n1274) );
XOR2_X1 U914 ( .A(n1279), .B(n1280), .Z(n1277) );
XOR2_X1 U915 ( .A(G140), .B(G110), .Z(n1280) );
XOR2_X1 U916 ( .A(n1281), .B(n1282), .Z(n1279) );
NAND2_X1 U917 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
NAND2_X1 U918 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U919 ( .A1(KEYINPUT53), .A2(n1287), .ZN(n1286) );
NAND2_X1 U920 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
INV_X1 U921 ( .A(n1290), .ZN(n1285) );
NAND2_X1 U922 ( .A1(n1272), .A2(n1291), .ZN(n1283) );
NAND2_X1 U923 ( .A1(n1289), .A2(n1292), .ZN(n1291) );
NAND2_X1 U924 ( .A1(n1290), .A2(KEYINPUT53), .ZN(n1292) );
XOR2_X1 U925 ( .A(n1293), .B(n1294), .Z(n1290) );
XNOR2_X1 U926 ( .A(n1295), .B(KEYINPUT35), .ZN(n1294) );
NAND2_X1 U927 ( .A1(KEYINPUT0), .A2(n1221), .ZN(n1295) );
INV_X1 U928 ( .A(KEYINPUT9), .ZN(n1289) );
NAND2_X1 U929 ( .A1(n1256), .A2(G469), .ZN(n1278) );
INV_X1 U930 ( .A(n1251), .ZN(n1256) );
NOR2_X1 U931 ( .A1(n1244), .A2(n1296), .ZN(G51) );
XOR2_X1 U932 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U933 ( .A1(n1198), .A2(n1251), .ZN(n1298) );
NAND2_X1 U934 ( .A1(G902), .A2(n1140), .ZN(n1251) );
NAND3_X1 U935 ( .A1(n1299), .A2(n1224), .A3(n1300), .ZN(n1140) );
XOR2_X1 U936 ( .A(n1225), .B(KEYINPUT59), .Z(n1300) );
AND4_X1 U937 ( .A1(n1301), .A2(n1302), .A3(n1303), .A4(n1304), .ZN(n1224) );
NOR4_X1 U938 ( .A1(n1305), .A2(n1306), .A3(n1307), .A4(n1308), .ZN(n1304) );
INV_X1 U939 ( .A(n1309), .ZN(n1306) );
NAND2_X1 U940 ( .A1(n1160), .A2(n1310), .ZN(n1303) );
XOR2_X1 U941 ( .A(KEYINPUT39), .B(n1311), .Z(n1310) );
INV_X1 U942 ( .A(n1235), .ZN(n1299) );
NAND4_X1 U943 ( .A1(n1261), .A2(n1312), .A3(n1313), .A4(n1314), .ZN(n1235) );
AND4_X1 U944 ( .A1(n1315), .A2(n1316), .A3(n1317), .A4(n1318), .ZN(n1314) );
NAND2_X1 U945 ( .A1(n1319), .A2(n1320), .ZN(n1313) );
NAND2_X1 U946 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XNOR2_X1 U947 ( .A(KEYINPUT18), .B(n1134), .ZN(n1321) );
NAND3_X1 U948 ( .A1(n1323), .A2(n1324), .A3(n1156), .ZN(n1134) );
NAND4_X1 U949 ( .A1(n1155), .A2(n1319), .A3(n1323), .A4(n1324), .ZN(n1261) );
NAND2_X1 U950 ( .A1(n1325), .A2(KEYINPUT50), .ZN(n1297) );
XOR2_X1 U951 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U952 ( .A(n1328), .B(n1329), .ZN(n1326) );
NOR2_X1 U953 ( .A1(n1330), .A2(G952), .ZN(n1244) );
XOR2_X1 U954 ( .A(G953), .B(KEYINPUT10), .Z(n1330) );
XOR2_X1 U955 ( .A(n1331), .B(n1301), .Z(G48) );
NAND3_X1 U956 ( .A1(n1155), .A2(n1319), .A3(n1332), .ZN(n1301) );
XNOR2_X1 U957 ( .A(G143), .B(n1302), .ZN(G45) );
NAND4_X1 U958 ( .A1(n1333), .A2(n1183), .A3(n1334), .A4(n1335), .ZN(n1302) );
XOR2_X1 U959 ( .A(G140), .B(n1308), .Z(G42) );
AND2_X1 U960 ( .A1(n1336), .A2(n1337), .ZN(n1308) );
XNOR2_X1 U961 ( .A(G137), .B(n1338), .ZN(G39) );
NAND2_X1 U962 ( .A1(n1311), .A2(n1160), .ZN(n1338) );
AND2_X1 U963 ( .A1(n1332), .A2(n1157), .ZN(n1311) );
NAND3_X1 U964 ( .A1(n1339), .A2(n1340), .A3(n1341), .ZN(G36) );
NAND2_X1 U965 ( .A1(G134), .A2(n1342), .ZN(n1341) );
NAND2_X1 U966 ( .A1(n1343), .A2(n1344), .ZN(n1340) );
INV_X1 U967 ( .A(KEYINPUT19), .ZN(n1344) );
NAND2_X1 U968 ( .A1(n1345), .A2(n1307), .ZN(n1343) );
INV_X1 U969 ( .A(n1342), .ZN(n1307) );
XOR2_X1 U970 ( .A(KEYINPUT57), .B(n1217), .Z(n1345) );
NAND2_X1 U971 ( .A1(KEYINPUT19), .A2(n1346), .ZN(n1339) );
NAND2_X1 U972 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
OR3_X1 U973 ( .A1(n1342), .A2(G134), .A3(KEYINPUT57), .ZN(n1348) );
NAND3_X1 U974 ( .A1(n1177), .A2(n1156), .A3(n1337), .ZN(n1342) );
NAND2_X1 U975 ( .A1(KEYINPUT57), .A2(G134), .ZN(n1347) );
XOR2_X1 U976 ( .A(n1349), .B(n1309), .Z(G33) );
NAND3_X1 U977 ( .A1(n1155), .A2(n1177), .A3(n1337), .ZN(n1309) );
AND3_X1 U978 ( .A1(n1159), .A2(n1334), .A3(n1160), .ZN(n1337) );
NOR2_X1 U979 ( .A1(n1175), .A2(n1182), .ZN(n1160) );
INV_X1 U980 ( .A(n1176), .ZN(n1182) );
XNOR2_X1 U981 ( .A(n1350), .B(KEYINPUT40), .ZN(n1175) );
XOR2_X1 U982 ( .A(G128), .B(n1305), .Z(G30) );
AND3_X1 U983 ( .A1(n1319), .A2(n1156), .A3(n1332), .ZN(n1305) );
AND4_X1 U984 ( .A1(n1159), .A2(n1169), .A3(n1334), .A4(n1172), .ZN(n1332) );
XNOR2_X1 U985 ( .A(G101), .B(n1312), .ZN(G3) );
NAND3_X1 U986 ( .A1(n1157), .A2(n1351), .A3(n1333), .ZN(n1312) );
AND3_X1 U987 ( .A1(n1319), .A2(n1159), .A3(n1177), .ZN(n1333) );
INV_X1 U988 ( .A(n1135), .ZN(n1319) );
XOR2_X1 U989 ( .A(n1352), .B(n1353), .Z(G27) );
NAND2_X1 U990 ( .A1(KEYINPUT63), .A2(n1354), .ZN(n1353) );
INV_X1 U991 ( .A(n1225), .ZN(n1354) );
NAND3_X1 U992 ( .A1(n1355), .A2(n1334), .A3(n1336), .ZN(n1225) );
AND3_X1 U993 ( .A1(n1356), .A2(n1172), .A3(n1155), .ZN(n1336) );
NAND2_X1 U994 ( .A1(n1142), .A2(n1357), .ZN(n1334) );
NAND3_X1 U995 ( .A1(G902), .A2(n1358), .A3(n1212), .ZN(n1357) );
NOR2_X1 U996 ( .A1(n1206), .A2(G900), .ZN(n1212) );
XNOR2_X1 U997 ( .A(G122), .B(n1317), .ZN(G24) );
NAND4_X1 U998 ( .A1(n1359), .A2(n1360), .A3(n1183), .A4(n1335), .ZN(n1317) );
INV_X1 U999 ( .A(n1145), .ZN(n1359) );
NAND2_X1 U1000 ( .A1(n1323), .A2(n1356), .ZN(n1145) );
INV_X1 U1001 ( .A(n1172), .ZN(n1323) );
XOR2_X1 U1002 ( .A(n1361), .B(n1316), .Z(G21) );
NAND4_X1 U1003 ( .A1(n1157), .A2(n1360), .A3(n1169), .A4(n1172), .ZN(n1316) );
INV_X1 U1004 ( .A(n1356), .ZN(n1169) );
NAND2_X1 U1005 ( .A1(n1362), .A2(n1363), .ZN(G18) );
OR2_X1 U1006 ( .A1(n1364), .A2(G116), .ZN(n1363) );
NAND2_X1 U1007 ( .A1(G116), .A2(n1365), .ZN(n1362) );
NAND2_X1 U1008 ( .A1(n1366), .A2(n1367), .ZN(n1365) );
OR2_X1 U1009 ( .A1(n1318), .A2(KEYINPUT20), .ZN(n1367) );
NAND2_X1 U1010 ( .A1(KEYINPUT20), .A2(n1364), .ZN(n1366) );
OR2_X1 U1011 ( .A1(KEYINPUT58), .A2(n1318), .ZN(n1364) );
NAND3_X1 U1012 ( .A1(n1360), .A2(n1156), .A3(n1177), .ZN(n1318) );
NOR2_X1 U1013 ( .A1(n1183), .A2(n1368), .ZN(n1156) );
XOR2_X1 U1014 ( .A(n1315), .B(n1369), .Z(G15) );
NAND2_X1 U1015 ( .A1(KEYINPUT12), .A2(G113), .ZN(n1369) );
NAND3_X1 U1016 ( .A1(n1177), .A2(n1360), .A3(n1155), .ZN(n1315) );
AND2_X1 U1017 ( .A1(n1368), .A2(n1183), .ZN(n1155) );
INV_X1 U1018 ( .A(n1335), .ZN(n1368) );
AND2_X1 U1019 ( .A1(n1355), .A2(n1351), .ZN(n1360) );
NOR3_X1 U1020 ( .A1(n1151), .A2(n1154), .A3(n1135), .ZN(n1355) );
INV_X1 U1021 ( .A(n1158), .ZN(n1154) );
NOR2_X1 U1022 ( .A1(n1172), .A2(n1356), .ZN(n1177) );
XOR2_X1 U1023 ( .A(G110), .B(n1370), .Z(G12) );
NOR2_X1 U1024 ( .A1(n1371), .A2(n1135), .ZN(n1370) );
NAND2_X1 U1025 ( .A1(n1350), .A2(n1176), .ZN(n1135) );
NAND2_X1 U1026 ( .A1(n1372), .A2(n1373), .ZN(n1176) );
XNOR2_X1 U1027 ( .A(G214), .B(KEYINPUT44), .ZN(n1372) );
XNOR2_X1 U1028 ( .A(n1199), .B(n1198), .ZN(n1350) );
NAND2_X1 U1029 ( .A1(G210), .A2(n1373), .ZN(n1198) );
NAND2_X1 U1030 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
INV_X1 U1031 ( .A(G237), .ZN(n1374) );
AND2_X1 U1032 ( .A1(n1376), .A2(n1375), .ZN(n1199) );
XOR2_X1 U1033 ( .A(n1377), .B(n1327), .Z(n1376) );
AND2_X1 U1034 ( .A1(n1378), .A2(n1379), .ZN(n1327) );
NAND2_X1 U1035 ( .A1(n1380), .A2(n1239), .ZN(n1379) );
XOR2_X1 U1036 ( .A(n1381), .B(KEYINPUT25), .Z(n1380) );
NAND2_X1 U1037 ( .A1(n1382), .A2(n1383), .ZN(n1378) );
XOR2_X1 U1038 ( .A(n1381), .B(KEYINPUT43), .Z(n1383) );
XOR2_X1 U1039 ( .A(n1240), .B(n1242), .Z(n1381) );
XNOR2_X1 U1040 ( .A(n1384), .B(n1385), .ZN(n1242) );
NOR2_X1 U1041 ( .A1(G107), .A2(KEYINPUT41), .ZN(n1385) );
INV_X1 U1042 ( .A(n1239), .ZN(n1382) );
XNOR2_X1 U1043 ( .A(G110), .B(n1386), .ZN(n1239) );
XOR2_X1 U1044 ( .A(KEYINPUT13), .B(G122), .Z(n1386) );
NOR2_X1 U1045 ( .A1(KEYINPUT61), .A2(n1387), .ZN(n1377) );
XOR2_X1 U1046 ( .A(n1329), .B(n1388), .Z(n1387) );
NAND2_X1 U1047 ( .A1(n1389), .A2(n1390), .ZN(n1388) );
OR3_X1 U1048 ( .A1(n1352), .A2(n1391), .A3(KEYINPUT31), .ZN(n1390) );
NAND2_X1 U1049 ( .A1(n1328), .A2(KEYINPUT31), .ZN(n1389) );
XOR2_X1 U1050 ( .A(n1352), .B(n1391), .Z(n1328) );
INV_X1 U1051 ( .A(G125), .ZN(n1352) );
NAND2_X1 U1052 ( .A1(G224), .A2(n1392), .ZN(n1329) );
XOR2_X1 U1053 ( .A(KEYINPUT4), .B(G953), .Z(n1392) );
XOR2_X1 U1054 ( .A(n1322), .B(KEYINPUT27), .Z(n1371) );
NAND3_X1 U1055 ( .A1(n1324), .A2(n1172), .A3(n1157), .ZN(n1322) );
NOR2_X1 U1056 ( .A1(n1335), .A2(n1183), .ZN(n1157) );
XOR2_X1 U1057 ( .A(G475), .B(n1393), .Z(n1183) );
AND2_X1 U1058 ( .A1(n1258), .A2(n1375), .ZN(n1393) );
NAND2_X1 U1059 ( .A1(n1394), .A2(n1395), .ZN(n1258) );
NAND2_X1 U1060 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
XOR2_X1 U1061 ( .A(KEYINPUT38), .B(n1398), .Z(n1394) );
NOR2_X1 U1062 ( .A1(n1397), .A2(n1396), .ZN(n1398) );
XOR2_X1 U1063 ( .A(n1399), .B(n1400), .Z(n1396) );
XNOR2_X1 U1064 ( .A(n1401), .B(n1402), .ZN(n1400) );
AND2_X1 U1065 ( .A1(G214), .A2(n1403), .ZN(n1402) );
XOR2_X1 U1066 ( .A(n1404), .B(n1405), .Z(n1399) );
NOR2_X1 U1067 ( .A1(n1220), .A2(n1406), .ZN(n1405) );
XOR2_X1 U1068 ( .A(n1219), .B(KEYINPUT37), .Z(n1406) );
NAND2_X1 U1069 ( .A1(KEYINPUT62), .A2(n1349), .ZN(n1404) );
INV_X1 U1070 ( .A(G131), .ZN(n1349) );
XOR2_X1 U1071 ( .A(G104), .B(n1407), .Z(n1397) );
XOR2_X1 U1072 ( .A(G122), .B(G113), .Z(n1407) );
NAND2_X1 U1073 ( .A1(n1408), .A2(n1202), .ZN(n1335) );
NAND2_X1 U1074 ( .A1(G478), .A2(n1409), .ZN(n1202) );
XOR2_X1 U1075 ( .A(n1201), .B(KEYINPUT36), .Z(n1408) );
OR2_X1 U1076 ( .A1(n1409), .A2(G478), .ZN(n1201) );
NAND2_X1 U1077 ( .A1(n1255), .A2(n1375), .ZN(n1409) );
XOR2_X1 U1078 ( .A(n1410), .B(n1411), .Z(n1255) );
XOR2_X1 U1079 ( .A(n1412), .B(n1413), .Z(n1411) );
XOR2_X1 U1080 ( .A(G107), .B(n1414), .Z(n1413) );
NOR2_X1 U1081 ( .A1(n1415), .A2(n1416), .ZN(n1414) );
INV_X1 U1082 ( .A(G217), .ZN(n1416) );
XOR2_X1 U1083 ( .A(n1417), .B(n1418), .Z(n1410) );
XOR2_X1 U1084 ( .A(G134), .B(G128), .Z(n1418) );
XNOR2_X1 U1085 ( .A(G116), .B(G122), .ZN(n1417) );
NAND2_X1 U1086 ( .A1(n1419), .A2(n1420), .ZN(n1172) );
NAND2_X1 U1087 ( .A1(n1191), .A2(n1196), .ZN(n1420) );
XOR2_X1 U1088 ( .A(KEYINPUT48), .B(n1421), .Z(n1419) );
NOR2_X1 U1089 ( .A1(n1191), .A2(n1196), .ZN(n1421) );
NAND2_X1 U1090 ( .A1(G217), .A2(n1422), .ZN(n1196) );
NOR2_X1 U1091 ( .A1(n1250), .A2(n1423), .ZN(n1191) );
XOR2_X1 U1092 ( .A(KEYINPUT46), .B(n1375), .Z(n1423) );
XNOR2_X1 U1093 ( .A(n1424), .B(n1425), .ZN(n1250) );
XOR2_X1 U1094 ( .A(n1426), .B(n1427), .Z(n1425) );
XOR2_X1 U1095 ( .A(KEYINPUT6), .B(G137), .Z(n1427) );
NOR2_X1 U1096 ( .A1(n1428), .A2(n1220), .ZN(n1426) );
NOR2_X1 U1097 ( .A1(n1429), .A2(G125), .ZN(n1220) );
INV_X1 U1098 ( .A(n1219), .ZN(n1428) );
NAND2_X1 U1099 ( .A1(G125), .A2(n1429), .ZN(n1219) );
XOR2_X1 U1100 ( .A(n1430), .B(n1431), .Z(n1424) );
NOR2_X1 U1101 ( .A1(n1415), .A2(n1432), .ZN(n1431) );
INV_X1 U1102 ( .A(G221), .ZN(n1432) );
NAND2_X1 U1103 ( .A1(n1433), .A2(n1206), .ZN(n1415) );
XNOR2_X1 U1104 ( .A(G234), .B(KEYINPUT11), .ZN(n1433) );
XOR2_X1 U1105 ( .A(n1434), .B(n1435), .Z(n1430) );
NOR2_X1 U1106 ( .A1(KEYINPUT2), .A2(n1331), .ZN(n1435) );
NAND2_X1 U1107 ( .A1(n1436), .A2(n1437), .ZN(n1434) );
OR2_X1 U1108 ( .A1(n1438), .A2(G110), .ZN(n1437) );
XOR2_X1 U1109 ( .A(n1439), .B(KEYINPUT17), .Z(n1436) );
NAND2_X1 U1110 ( .A1(G110), .A2(n1438), .ZN(n1439) );
XNOR2_X1 U1111 ( .A(n1361), .B(G128), .ZN(n1438) );
INV_X1 U1112 ( .A(G119), .ZN(n1361) );
AND3_X1 U1113 ( .A1(n1356), .A2(n1351), .A3(n1159), .ZN(n1324) );
INV_X1 U1114 ( .A(n1163), .ZN(n1159) );
NAND2_X1 U1115 ( .A1(n1151), .A2(n1158), .ZN(n1163) );
NAND2_X1 U1116 ( .A1(G221), .A2(n1422), .ZN(n1158) );
NAND2_X1 U1117 ( .A1(G234), .A2(n1375), .ZN(n1422) );
XOR2_X1 U1118 ( .A(n1440), .B(n1441), .Z(n1151) );
XOR2_X1 U1119 ( .A(KEYINPUT23), .B(G469), .Z(n1441) );
NAND2_X1 U1120 ( .A1(n1442), .A2(n1375), .ZN(n1440) );
XOR2_X1 U1121 ( .A(n1443), .B(n1444), .Z(n1442) );
XOR2_X1 U1122 ( .A(n1429), .B(n1445), .Z(n1444) );
NAND2_X1 U1123 ( .A1(n1446), .A2(n1447), .ZN(n1445) );
OR2_X1 U1124 ( .A1(n1448), .A2(n1288), .ZN(n1447) );
XOR2_X1 U1125 ( .A(n1449), .B(KEYINPUT15), .Z(n1446) );
NAND2_X1 U1126 ( .A1(n1288), .A2(n1448), .ZN(n1449) );
XNOR2_X1 U1127 ( .A(n1450), .B(n1451), .ZN(n1448) );
INV_X1 U1128 ( .A(n1293), .ZN(n1451) );
XOR2_X1 U1129 ( .A(G107), .B(n1384), .Z(n1293) );
XOR2_X1 U1130 ( .A(G101), .B(n1260), .Z(n1384) );
INV_X1 U1131 ( .A(G104), .ZN(n1260) );
XNOR2_X1 U1132 ( .A(KEYINPUT54), .B(n1452), .ZN(n1450) );
NOR2_X1 U1133 ( .A1(KEYINPUT34), .A2(n1453), .ZN(n1452) );
INV_X1 U1134 ( .A(n1221), .ZN(n1453) );
XNOR2_X1 U1135 ( .A(n1401), .B(G128), .ZN(n1221) );
INV_X1 U1136 ( .A(G140), .ZN(n1429) );
XNOR2_X1 U1137 ( .A(n1282), .B(n1454), .ZN(n1443) );
NOR2_X1 U1138 ( .A1(G110), .A2(KEYINPUT51), .ZN(n1454) );
AND2_X1 U1139 ( .A1(G227), .A2(n1206), .ZN(n1282) );
NAND2_X1 U1140 ( .A1(n1142), .A2(n1455), .ZN(n1351) );
NAND3_X1 U1141 ( .A1(G902), .A2(n1358), .A3(n1237), .ZN(n1455) );
NOR2_X1 U1142 ( .A1(n1206), .A2(G898), .ZN(n1237) );
NAND3_X1 U1143 ( .A1(n1358), .A2(n1206), .A3(G952), .ZN(n1142) );
INV_X1 U1144 ( .A(G953), .ZN(n1206) );
NAND2_X1 U1145 ( .A1(G237), .A2(G234), .ZN(n1358) );
XNOR2_X1 U1146 ( .A(n1187), .B(G472), .ZN(n1356) );
AND3_X1 U1147 ( .A1(n1456), .A2(n1457), .A3(n1375), .ZN(n1187) );
INV_X1 U1148 ( .A(G902), .ZN(n1375) );
NAND2_X1 U1149 ( .A1(n1458), .A2(n1459), .ZN(n1457) );
INV_X1 U1150 ( .A(KEYINPUT47), .ZN(n1459) );
XOR2_X1 U1151 ( .A(n1265), .B(n1460), .Z(n1458) );
NAND3_X1 U1152 ( .A1(n1460), .A2(n1265), .A3(KEYINPUT47), .ZN(n1456) );
XNOR2_X1 U1153 ( .A(n1461), .B(G101), .ZN(n1265) );
NAND2_X1 U1154 ( .A1(n1403), .A2(G210), .ZN(n1461) );
NOR2_X1 U1155 ( .A1(G953), .A2(G237), .ZN(n1403) );
XOR2_X1 U1156 ( .A(n1266), .B(n1462), .Z(n1460) );
XOR2_X1 U1157 ( .A(n1391), .B(n1272), .Z(n1462) );
INV_X1 U1158 ( .A(n1288), .ZN(n1272) );
XOR2_X1 U1159 ( .A(n1463), .B(n1222), .Z(n1288) );
XOR2_X1 U1160 ( .A(G131), .B(G137), .Z(n1222) );
NAND2_X1 U1161 ( .A1(KEYINPUT33), .A2(n1217), .ZN(n1463) );
INV_X1 U1162 ( .A(G134), .ZN(n1217) );
INV_X1 U1163 ( .A(n1270), .ZN(n1391) );
XOR2_X1 U1164 ( .A(n1464), .B(G128), .Z(n1270) );
NAND2_X1 U1165 ( .A1(n1465), .A2(n1466), .ZN(n1464) );
NAND2_X1 U1166 ( .A1(n1401), .A2(n1467), .ZN(n1466) );
XNOR2_X1 U1167 ( .A(n1331), .B(n1412), .ZN(n1401) );
INV_X1 U1168 ( .A(G146), .ZN(n1331) );
OR3_X1 U1169 ( .A1(n1412), .A2(G146), .A3(n1467), .ZN(n1465) );
INV_X1 U1170 ( .A(KEYINPUT32), .ZN(n1467) );
XOR2_X1 U1171 ( .A(G143), .B(KEYINPUT28), .Z(n1412) );
INV_X1 U1172 ( .A(n1240), .ZN(n1266) );
XNOR2_X1 U1173 ( .A(G113), .B(n1468), .ZN(n1240) );
XOR2_X1 U1174 ( .A(G119), .B(G116), .Z(n1468) );
endmodule


