//Key = 0100000111000110000010100100011101011010000110100001110100000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;

XNOR2_X1 U755 ( .A(G107), .B(n1034), .ZN(G9) );
NOR2_X1 U756 ( .A1(n1035), .A2(n1036), .ZN(G75) );
NOR4_X1 U757 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
NOR2_X1 U758 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NOR3_X1 U759 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1041) );
NOR2_X1 U760 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NOR2_X1 U761 ( .A1(n1048), .A2(n1049), .ZN(n1046) );
NOR2_X1 U762 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U763 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U764 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR3_X1 U765 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1052) );
NOR3_X1 U766 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1048) );
NOR3_X1 U767 ( .A1(n1060), .A2(n1062), .A3(n1051), .ZN(n1044) );
INV_X1 U768 ( .A(n1063), .ZN(n1060) );
NOR2_X1 U769 ( .A1(n1064), .A2(n1065), .ZN(n1043) );
NAND3_X1 U770 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1037) );
NAND2_X1 U771 ( .A1(n1069), .A2(n1065), .ZN(n1068) );
INV_X1 U772 ( .A(KEYINPUT8), .ZN(n1065) );
OR2_X1 U773 ( .A1(n1042), .A2(n1064), .ZN(n1069) );
AND2_X1 U774 ( .A1(n1070), .A2(n1071), .ZN(n1064) );
NAND3_X1 U775 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1071) );
NAND2_X1 U776 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND3_X1 U777 ( .A1(n1056), .A2(n1058), .A3(n1077), .ZN(n1076) );
NAND2_X1 U778 ( .A1(n1078), .A2(n1079), .ZN(n1075) );
NAND2_X1 U779 ( .A1(n1063), .A2(n1080), .ZN(n1070) );
NAND2_X1 U780 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U782 ( .A(n1074), .B(KEYINPUT44), .ZN(n1083) );
NAND2_X1 U783 ( .A1(n1085), .A2(n1072), .ZN(n1081) );
NOR2_X1 U784 ( .A1(n1055), .A2(n1057), .ZN(n1063) );
INV_X1 U785 ( .A(n1077), .ZN(n1057) );
INV_X1 U786 ( .A(n1079), .ZN(n1055) );
NOR3_X1 U787 ( .A1(n1086), .A2(G953), .A3(G952), .ZN(n1035) );
INV_X1 U788 ( .A(n1066), .ZN(n1086) );
NAND4_X1 U789 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1066) );
NOR3_X1 U790 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
XOR2_X1 U791 ( .A(n1094), .B(KEYINPUT45), .Z(n1093) );
NAND4_X1 U792 ( .A1(n1072), .A2(n1095), .A3(n1056), .A4(n1096), .ZN(n1094) );
NAND2_X1 U793 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
XNOR2_X1 U794 ( .A(n1099), .B(KEYINPUT52), .ZN(n1097) );
NOR3_X1 U795 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1092) );
NOR2_X1 U796 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U797 ( .A1(KEYINPUT24), .A2(n1105), .ZN(n1103) );
NOR4_X1 U798 ( .A1(G478), .A2(n1106), .A3(KEYINPUT24), .A4(n1105), .ZN(n1101) );
AND2_X1 U799 ( .A1(n1106), .A2(n1105), .ZN(n1100) );
XOR2_X1 U800 ( .A(KEYINPUT60), .B(KEYINPUT6), .Z(n1106) );
XNOR2_X1 U801 ( .A(n1107), .B(n1108), .ZN(n1089) );
NOR2_X1 U802 ( .A1(KEYINPUT47), .A2(n1109), .ZN(n1108) );
NAND2_X1 U803 ( .A1(n1110), .A2(n1111), .ZN(n1088) );
NAND2_X1 U804 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NAND3_X1 U805 ( .A1(n1112), .A2(n1113), .A3(G472), .ZN(n1087) );
INV_X1 U806 ( .A(KEYINPUT21), .ZN(n1113) );
XOR2_X1 U807 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U808 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U809 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR2_X1 U810 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NOR2_X1 U811 ( .A1(n1120), .A2(n1122), .ZN(n1116) );
INV_X1 U812 ( .A(n1118), .ZN(n1122) );
NOR2_X1 U813 ( .A1(n1123), .A2(n1121), .ZN(n1118) );
XOR2_X1 U814 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U815 ( .A1(KEYINPUT32), .A2(n1126), .ZN(n1125) );
XOR2_X1 U816 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U817 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U818 ( .A1(KEYINPUT41), .A2(n1131), .ZN(n1129) );
NOR2_X1 U819 ( .A1(G227), .A2(n1067), .ZN(n1120) );
NAND2_X1 U820 ( .A1(n1067), .A2(n1038), .ZN(n1114) );
XOR2_X1 U821 ( .A(n1132), .B(n1133), .Z(G69) );
NOR2_X1 U822 ( .A1(n1134), .A2(n1067), .ZN(n1133) );
NOR2_X1 U823 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U824 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NAND2_X1 U825 ( .A1(n1139), .A2(n1067), .ZN(n1138) );
XOR2_X1 U826 ( .A(n1040), .B(n1140), .Z(n1139) );
NAND3_X1 U827 ( .A1(G898), .A2(n1140), .A3(G953), .ZN(n1137) );
XNOR2_X1 U828 ( .A(n1141), .B(n1142), .ZN(n1140) );
XNOR2_X1 U829 ( .A(n1143), .B(G110), .ZN(n1141) );
NOR2_X1 U830 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XOR2_X1 U831 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR3_X1 U832 ( .A1(n1148), .A2(KEYINPUT2), .A3(n1109), .ZN(n1147) );
NOR2_X1 U833 ( .A1(n1144), .A2(n1149), .ZN(G63) );
NOR3_X1 U834 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1149) );
AND2_X1 U835 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U836 ( .A1(n1155), .A2(n1153), .ZN(n1151) );
NOR2_X1 U837 ( .A1(n1156), .A2(n1105), .ZN(n1155) );
NOR2_X1 U838 ( .A1(n1157), .A2(n1154), .ZN(n1156) );
NOR2_X1 U839 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U840 ( .A1(n1040), .A2(n1038), .ZN(n1158) );
NOR3_X1 U841 ( .A1(n1159), .A2(n1160), .A3(n1148), .ZN(n1150) );
NOR2_X1 U842 ( .A1(n1154), .A2(n1153), .ZN(n1160) );
INV_X1 U843 ( .A(KEYINPUT43), .ZN(n1153) );
XNOR2_X1 U844 ( .A(n1104), .B(KEYINPUT9), .ZN(n1159) );
NOR2_X1 U845 ( .A1(n1144), .A2(n1161), .ZN(G60) );
XOR2_X1 U846 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U847 ( .A1(n1164), .A2(G475), .ZN(n1162) );
XNOR2_X1 U848 ( .A(G104), .B(n1165), .ZN(G6) );
NOR2_X1 U849 ( .A1(n1144), .A2(n1166), .ZN(G57) );
XOR2_X1 U850 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U851 ( .A(n1169), .B(n1170), .Z(n1167) );
NOR2_X1 U852 ( .A1(n1111), .A2(n1148), .ZN(n1170) );
NAND2_X1 U853 ( .A1(KEYINPUT13), .A2(n1171), .ZN(n1169) );
XOR2_X1 U854 ( .A(G101), .B(n1172), .Z(n1171) );
NOR2_X1 U855 ( .A1(n1144), .A2(n1173), .ZN(G54) );
XOR2_X1 U856 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U857 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR2_X1 U858 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U859 ( .A(KEYINPUT15), .B(n1180), .Z(n1179) );
NOR2_X1 U860 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
AND2_X1 U861 ( .A1(n1182), .A2(n1181), .ZN(n1178) );
XNOR2_X1 U862 ( .A(n1127), .B(KEYINPUT14), .ZN(n1182) );
NOR3_X1 U863 ( .A1(n1148), .A2(KEYINPUT58), .A3(n1183), .ZN(n1176) );
INV_X1 U864 ( .A(G469), .ZN(n1183) );
XOR2_X1 U865 ( .A(n1184), .B(n1185), .Z(n1174) );
NAND2_X1 U866 ( .A1(KEYINPUT63), .A2(n1186), .ZN(n1184) );
XOR2_X1 U867 ( .A(n1187), .B(n1188), .Z(n1186) );
NAND2_X1 U868 ( .A1(KEYINPUT55), .A2(n1189), .ZN(n1188) );
NOR2_X1 U869 ( .A1(n1144), .A2(n1190), .ZN(G51) );
XOR2_X1 U870 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U871 ( .A(n1193), .B(n1194), .Z(n1191) );
NAND2_X1 U872 ( .A1(n1164), .A2(n1195), .ZN(n1193) );
INV_X1 U873 ( .A(n1148), .ZN(n1164) );
NAND2_X1 U874 ( .A1(G902), .A2(n1196), .ZN(n1148) );
OR2_X1 U875 ( .A1(n1038), .A2(n1040), .ZN(n1196) );
NAND4_X1 U876 ( .A1(n1165), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1040) );
AND4_X1 U877 ( .A1(n1034), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1199) );
NAND3_X1 U878 ( .A1(n1203), .A2(n1077), .A3(n1204), .ZN(n1034) );
NOR2_X1 U879 ( .A1(n1205), .A2(n1206), .ZN(n1198) );
NOR2_X1 U880 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U881 ( .A(n1209), .B(KEYINPUT18), .Z(n1207) );
AND3_X1 U882 ( .A1(n1210), .A2(n1077), .A3(n1211), .ZN(n1205) );
NAND3_X1 U883 ( .A1(n1204), .A2(n1077), .A3(n1085), .ZN(n1165) );
NAND2_X1 U884 ( .A1(n1212), .A2(n1213), .ZN(n1038) );
NOR4_X1 U885 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1213) );
NOR4_X1 U886 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1212) );
NOR2_X1 U887 ( .A1(KEYINPUT50), .A2(n1222), .ZN(n1221) );
NOR2_X1 U888 ( .A1(n1223), .A2(n1224), .ZN(n1220) );
NOR2_X1 U889 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
NOR2_X1 U890 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XNOR2_X1 U891 ( .A(n1203), .B(KEYINPUT59), .ZN(n1227) );
AND4_X1 U892 ( .A1(n1208), .A2(n1229), .A3(n1211), .A4(KEYINPUT50), .ZN(n1225) );
NOR3_X1 U893 ( .A1(n1047), .A2(n1230), .A3(n1228), .ZN(n1219) );
AND2_X1 U894 ( .A1(n1231), .A2(G953), .ZN(n1144) );
XNOR2_X1 U895 ( .A(G952), .B(KEYINPUT56), .ZN(n1231) );
XOR2_X1 U896 ( .A(G146), .B(n1218), .Z(G48) );
NOR4_X1 U897 ( .A1(n1230), .A2(n1232), .A3(n1233), .A4(n1208), .ZN(n1218) );
XNOR2_X1 U898 ( .A(G143), .B(n1222), .ZN(G45) );
NAND4_X1 U899 ( .A1(n1211), .A2(n1078), .A3(n1229), .A4(n1084), .ZN(n1222) );
XOR2_X1 U900 ( .A(G140), .B(n1217), .Z(G42) );
NOR3_X1 U901 ( .A1(n1233), .A2(n1054), .A3(n1228), .ZN(n1217) );
NAND3_X1 U902 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(G39) );
NAND3_X1 U903 ( .A1(n1237), .A2(n1238), .A3(KEYINPUT38), .ZN(n1236) );
NAND3_X1 U904 ( .A1(G137), .A2(n1239), .A3(n1240), .ZN(n1235) );
INV_X1 U905 ( .A(KEYINPUT10), .ZN(n1240) );
NAND2_X1 U906 ( .A1(KEYINPUT38), .A2(n1237), .ZN(n1239) );
NAND2_X1 U907 ( .A1(KEYINPUT10), .A2(n1241), .ZN(n1234) );
OR2_X1 U908 ( .A1(n1238), .A2(n1237), .ZN(n1241) );
NOR3_X1 U909 ( .A1(n1228), .A2(n1242), .A3(n1047), .ZN(n1237) );
XOR2_X1 U910 ( .A(KEYINPUT5), .B(n1230), .Z(n1242) );
XNOR2_X1 U911 ( .A(G134), .B(n1243), .ZN(G36) );
NAND2_X1 U912 ( .A1(n1244), .A2(n1203), .ZN(n1243) );
NAND2_X1 U913 ( .A1(n1245), .A2(n1246), .ZN(G33) );
NAND2_X1 U914 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND2_X1 U915 ( .A1(n1131), .A2(n1249), .ZN(n1247) );
NAND2_X1 U916 ( .A1(KEYINPUT57), .A2(n1250), .ZN(n1249) );
NAND3_X1 U917 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1245) );
INV_X1 U918 ( .A(KEYINPUT57), .ZN(n1253) );
NAND2_X1 U919 ( .A1(G131), .A2(n1250), .ZN(n1252) );
NAND2_X1 U920 ( .A1(n1254), .A2(n1131), .ZN(n1251) );
NAND2_X1 U921 ( .A1(n1216), .A2(n1250), .ZN(n1254) );
INV_X1 U922 ( .A(KEYINPUT23), .ZN(n1250) );
INV_X1 U923 ( .A(n1248), .ZN(n1216) );
NAND2_X1 U924 ( .A1(n1244), .A2(n1085), .ZN(n1248) );
NOR2_X1 U925 ( .A1(n1224), .A2(n1228), .ZN(n1244) );
NAND2_X1 U926 ( .A1(n1229), .A2(n1072), .ZN(n1228) );
INV_X1 U927 ( .A(n1051), .ZN(n1072) );
NAND2_X1 U928 ( .A1(n1255), .A2(n1059), .ZN(n1051) );
INV_X1 U929 ( .A(n1061), .ZN(n1255) );
INV_X1 U930 ( .A(n1232), .ZN(n1229) );
INV_X1 U931 ( .A(n1078), .ZN(n1224) );
XOR2_X1 U932 ( .A(G128), .B(n1215), .Z(G30) );
NOR4_X1 U933 ( .A1(n1230), .A2(n1232), .A3(n1062), .A4(n1208), .ZN(n1215) );
INV_X1 U934 ( .A(n1203), .ZN(n1062) );
NAND3_X1 U935 ( .A1(n1056), .A2(n1058), .A3(n1256), .ZN(n1232) );
XNOR2_X1 U936 ( .A(G101), .B(n1197), .ZN(G3) );
NAND3_X1 U937 ( .A1(n1078), .A2(n1204), .A3(n1074), .ZN(n1197) );
XNOR2_X1 U938 ( .A(G125), .B(n1257), .ZN(G27) );
NAND2_X1 U939 ( .A1(KEYINPUT1), .A2(n1214), .ZN(n1257) );
AND4_X1 U940 ( .A1(n1085), .A2(n1079), .A3(n1258), .A4(n1259), .ZN(n1214) );
AND2_X1 U941 ( .A1(n1256), .A2(n1084), .ZN(n1258) );
NAND2_X1 U942 ( .A1(n1042), .A2(n1260), .ZN(n1256) );
NAND2_X1 U943 ( .A1(n1121), .A2(n1261), .ZN(n1260) );
NOR2_X1 U944 ( .A1(G900), .A2(n1067), .ZN(n1121) );
XNOR2_X1 U945 ( .A(G122), .B(n1262), .ZN(G24) );
NAND4_X1 U946 ( .A1(KEYINPUT51), .A2(n1210), .A3(n1211), .A4(n1077), .ZN(n1262) );
NOR2_X1 U947 ( .A1(n1263), .A2(n1264), .ZN(n1077) );
NOR2_X1 U948 ( .A1(n1265), .A2(n1266), .ZN(n1211) );
XNOR2_X1 U949 ( .A(G119), .B(n1202), .ZN(G21) );
OR3_X1 U950 ( .A1(n1047), .A2(n1230), .A3(n1267), .ZN(n1202) );
NAND2_X1 U951 ( .A1(n1264), .A2(n1263), .ZN(n1230) );
XOR2_X1 U952 ( .A(n1268), .B(n1269), .Z(G18) );
NAND2_X1 U953 ( .A1(n1270), .A2(KEYINPUT25), .ZN(n1269) );
XNOR2_X1 U954 ( .A(G116), .B(KEYINPUT7), .ZN(n1270) );
NAND2_X1 U955 ( .A1(n1084), .A2(n1271), .ZN(n1268) );
XNOR2_X1 U956 ( .A(KEYINPUT27), .B(n1209), .ZN(n1271) );
NAND3_X1 U957 ( .A1(n1078), .A2(n1203), .A3(n1272), .ZN(n1209) );
NOR2_X1 U958 ( .A1(n1091), .A2(n1266), .ZN(n1203) );
XNOR2_X1 U959 ( .A(G113), .B(n1201), .ZN(G15) );
NAND3_X1 U960 ( .A1(n1078), .A2(n1085), .A3(n1210), .ZN(n1201) );
INV_X1 U961 ( .A(n1267), .ZN(n1210) );
NAND2_X1 U962 ( .A1(n1272), .A2(n1084), .ZN(n1267) );
AND2_X1 U963 ( .A1(n1079), .A2(n1273), .ZN(n1272) );
NOR2_X1 U964 ( .A1(n1058), .A2(n1274), .ZN(n1079) );
INV_X1 U965 ( .A(n1056), .ZN(n1274) );
INV_X1 U966 ( .A(n1233), .ZN(n1085) );
NAND2_X1 U967 ( .A1(n1266), .A2(n1091), .ZN(n1233) );
NOR2_X1 U968 ( .A1(n1263), .A2(n1275), .ZN(n1078) );
XNOR2_X1 U969 ( .A(n1200), .B(n1276), .ZN(G12) );
NOR2_X1 U970 ( .A1(KEYINPUT28), .A2(n1277), .ZN(n1276) );
NAND3_X1 U971 ( .A1(n1259), .A2(n1204), .A3(n1074), .ZN(n1200) );
INV_X1 U972 ( .A(n1047), .ZN(n1074) );
NAND2_X1 U973 ( .A1(n1266), .A2(n1265), .ZN(n1047) );
INV_X1 U974 ( .A(n1091), .ZN(n1265) );
XNOR2_X1 U975 ( .A(n1278), .B(G475), .ZN(n1091) );
NAND2_X1 U976 ( .A1(n1163), .A2(n1279), .ZN(n1278) );
XNOR2_X1 U977 ( .A(n1280), .B(n1281), .ZN(n1163) );
XOR2_X1 U978 ( .A(n1282), .B(n1283), .Z(n1281) );
XNOR2_X1 U979 ( .A(G143), .B(G131), .ZN(n1283) );
NAND2_X1 U980 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
OR2_X1 U981 ( .A1(n1124), .A2(n1286), .ZN(n1285) );
XOR2_X1 U982 ( .A(n1287), .B(KEYINPUT39), .Z(n1284) );
NAND2_X1 U983 ( .A1(n1124), .A2(n1286), .ZN(n1287) );
XOR2_X1 U984 ( .A(G125), .B(G140), .Z(n1124) );
XOR2_X1 U985 ( .A(n1288), .B(n1143), .Z(n1280) );
XOR2_X1 U986 ( .A(n1289), .B(G122), .Z(n1143) );
NAND2_X1 U987 ( .A1(KEYINPUT30), .A2(n1290), .ZN(n1288) );
NAND3_X1 U988 ( .A1(n1291), .A2(n1067), .A3(G214), .ZN(n1290) );
XOR2_X1 U989 ( .A(n1105), .B(n1104), .Z(n1266) );
INV_X1 U990 ( .A(G478), .ZN(n1104) );
NOR2_X1 U991 ( .A1(n1154), .A2(G902), .ZN(n1105) );
XOR2_X1 U992 ( .A(n1292), .B(n1293), .Z(n1154) );
XOR2_X1 U993 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U994 ( .A(G107), .B(G116), .ZN(n1295) );
NAND3_X1 U995 ( .A1(G234), .A2(n1067), .A3(G217), .ZN(n1294) );
XOR2_X1 U996 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U997 ( .A(G128), .B(G122), .Z(n1297) );
XNOR2_X1 U998 ( .A(G134), .B(G143), .ZN(n1296) );
AND4_X1 U999 ( .A1(n1084), .A2(n1273), .A3(n1056), .A4(n1058), .ZN(n1204) );
NAND2_X1 U1000 ( .A1(n1096), .A2(n1298), .ZN(n1058) );
NAND2_X1 U1001 ( .A1(n1099), .A2(n1098), .ZN(n1298) );
OR2_X1 U1002 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
XOR2_X1 U1003 ( .A(G469), .B(KEYINPUT19), .Z(n1099) );
NAND2_X1 U1004 ( .A1(n1299), .A2(n1279), .ZN(n1098) );
XOR2_X1 U1005 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U1006 ( .A(n1302), .B(n1303), .Z(n1301) );
XNOR2_X1 U1007 ( .A(KEYINPUT61), .B(n1187), .ZN(n1303) );
NAND2_X1 U1008 ( .A1(G227), .A2(n1067), .ZN(n1187) );
NOR2_X1 U1009 ( .A1(KEYINPUT49), .A2(n1189), .ZN(n1302) );
XNOR2_X1 U1010 ( .A(G110), .B(G140), .ZN(n1189) );
XNOR2_X1 U1011 ( .A(n1304), .B(n1181), .ZN(n1300) );
XNOR2_X1 U1012 ( .A(G104), .B(n1305), .ZN(n1181) );
XOR2_X1 U1013 ( .A(n1127), .B(n1185), .Z(n1304) );
XOR2_X1 U1014 ( .A(n1306), .B(n1307), .Z(n1127) );
XNOR2_X1 U1015 ( .A(KEYINPUT22), .B(n1308), .ZN(n1307) );
INV_X1 U1016 ( .A(G143), .ZN(n1308) );
XOR2_X1 U1017 ( .A(n1309), .B(G128), .Z(n1306) );
NAND2_X1 U1018 ( .A1(KEYINPUT33), .A2(n1310), .ZN(n1309) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1311), .ZN(n1056) );
NAND2_X1 U1020 ( .A1(n1042), .A2(n1312), .ZN(n1273) );
NAND3_X1 U1021 ( .A1(n1261), .A2(n1136), .A3(G953), .ZN(n1312) );
INV_X1 U1022 ( .A(G898), .ZN(n1136) );
AND2_X1 U1023 ( .A1(n1313), .A2(n1314), .ZN(n1261) );
XNOR2_X1 U1024 ( .A(KEYINPUT48), .B(n1279), .ZN(n1313) );
NAND3_X1 U1025 ( .A1(n1314), .A2(n1067), .A3(G952), .ZN(n1042) );
NAND2_X1 U1026 ( .A1(G237), .A2(G234), .ZN(n1314) );
INV_X1 U1027 ( .A(n1208), .ZN(n1084) );
NAND2_X1 U1028 ( .A1(n1061), .A2(n1059), .ZN(n1208) );
NAND2_X1 U1029 ( .A1(n1315), .A2(n1316), .ZN(n1059) );
XOR2_X1 U1030 ( .A(KEYINPUT62), .B(G214), .Z(n1315) );
XNOR2_X1 U1031 ( .A(n1317), .B(n1195), .ZN(n1061) );
AND2_X1 U1032 ( .A1(G210), .A2(n1316), .ZN(n1195) );
NAND2_X1 U1033 ( .A1(n1279), .A2(n1291), .ZN(n1316) );
NAND2_X1 U1034 ( .A1(n1318), .A2(n1279), .ZN(n1317) );
XNOR2_X1 U1035 ( .A(n1194), .B(n1319), .ZN(n1318) );
NOR2_X1 U1036 ( .A1(KEYINPUT37), .A2(n1192), .ZN(n1319) );
XNOR2_X1 U1037 ( .A(n1320), .B(n1321), .ZN(n1192) );
XNOR2_X1 U1038 ( .A(G125), .B(n1322), .ZN(n1320) );
NOR2_X1 U1039 ( .A1(G953), .A2(n1135), .ZN(n1322) );
INV_X1 U1040 ( .A(G224), .ZN(n1135) );
XOR2_X1 U1041 ( .A(n1142), .B(n1323), .Z(n1194) );
XOR2_X1 U1042 ( .A(n1324), .B(n1289), .Z(n1323) );
XNOR2_X1 U1043 ( .A(G104), .B(n1325), .ZN(n1289) );
INV_X1 U1044 ( .A(n1326), .ZN(n1325) );
NOR2_X1 U1045 ( .A1(KEYINPUT0), .A2(n1327), .ZN(n1324) );
XNOR2_X1 U1046 ( .A(G122), .B(n1277), .ZN(n1327) );
INV_X1 U1047 ( .A(G110), .ZN(n1277) );
XOR2_X1 U1048 ( .A(n1305), .B(n1328), .Z(n1142) );
XOR2_X1 U1049 ( .A(KEYINPUT3), .B(n1329), .Z(n1328) );
XOR2_X1 U1050 ( .A(G107), .B(G101), .Z(n1305) );
INV_X1 U1051 ( .A(n1054), .ZN(n1259) );
NAND2_X1 U1052 ( .A1(n1275), .A2(n1263), .ZN(n1054) );
NAND2_X1 U1053 ( .A1(n1330), .A2(n1331), .ZN(n1263) );
NAND2_X1 U1054 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XNOR2_X1 U1055 ( .A(n1334), .B(KEYINPUT26), .ZN(n1332) );
XOR2_X1 U1056 ( .A(n1335), .B(KEYINPUT54), .Z(n1330) );
NAND2_X1 U1057 ( .A1(n1107), .A2(n1336), .ZN(n1335) );
XNOR2_X1 U1058 ( .A(KEYINPUT17), .B(n1337), .ZN(n1336) );
INV_X1 U1059 ( .A(n1334), .ZN(n1337) );
XNOR2_X1 U1060 ( .A(n1109), .B(KEYINPUT35), .ZN(n1334) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1311), .ZN(n1109) );
NAND2_X1 U1062 ( .A1(G234), .A2(n1279), .ZN(n1311) );
INV_X1 U1063 ( .A(n1333), .ZN(n1107) );
NAND2_X1 U1064 ( .A1(n1338), .A2(n1279), .ZN(n1333) );
XOR2_X1 U1065 ( .A(n1146), .B(KEYINPUT46), .Z(n1338) );
XOR2_X1 U1066 ( .A(n1339), .B(n1340), .Z(n1146) );
XNOR2_X1 U1067 ( .A(n1238), .B(n1341), .ZN(n1340) );
NOR2_X1 U1068 ( .A1(KEYINPUT4), .A2(n1342), .ZN(n1341) );
XOR2_X1 U1069 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1070 ( .A(G110), .B(n1345), .ZN(n1344) );
NOR2_X1 U1071 ( .A1(KEYINPUT40), .A2(n1346), .ZN(n1345) );
XOR2_X1 U1072 ( .A(G128), .B(G119), .Z(n1346) );
NAND2_X1 U1073 ( .A1(n1347), .A2(n1348), .ZN(n1343) );
NAND2_X1 U1074 ( .A1(n1349), .A2(n1286), .ZN(n1348) );
XOR2_X1 U1075 ( .A(KEYINPUT36), .B(n1350), .Z(n1347) );
NOR2_X1 U1076 ( .A1(n1349), .A2(n1286), .ZN(n1350) );
XNOR2_X1 U1077 ( .A(G125), .B(n1351), .ZN(n1349) );
NOR2_X1 U1078 ( .A1(G140), .A2(KEYINPUT11), .ZN(n1351) );
NAND3_X1 U1079 ( .A1(G234), .A2(n1067), .A3(G221), .ZN(n1339) );
INV_X1 U1080 ( .A(n1264), .ZN(n1275) );
XOR2_X1 U1081 ( .A(n1112), .B(n1111), .Z(n1264) );
INV_X1 U1082 ( .A(G472), .ZN(n1111) );
NAND2_X1 U1083 ( .A1(n1352), .A2(n1279), .ZN(n1112) );
INV_X1 U1084 ( .A(G902), .ZN(n1279) );
XOR2_X1 U1085 ( .A(n1353), .B(n1354), .Z(n1352) );
XNOR2_X1 U1086 ( .A(n1355), .B(n1168), .ZN(n1354) );
XNOR2_X1 U1087 ( .A(n1356), .B(n1357), .ZN(n1168) );
XNOR2_X1 U1088 ( .A(n1321), .B(n1358), .ZN(n1357) );
XNOR2_X1 U1089 ( .A(n1326), .B(KEYINPUT42), .ZN(n1358) );
XOR2_X1 U1090 ( .A(G113), .B(KEYINPUT53), .Z(n1326) );
XOR2_X1 U1091 ( .A(n1359), .B(n1310), .Z(n1321) );
INV_X1 U1092 ( .A(n1286), .ZN(n1310) );
XOR2_X1 U1093 ( .A(G146), .B(KEYINPUT16), .Z(n1286) );
XOR2_X1 U1094 ( .A(n1360), .B(G128), .Z(n1359) );
NAND2_X1 U1095 ( .A1(KEYINPUT29), .A2(G143), .ZN(n1360) );
XNOR2_X1 U1096 ( .A(n1185), .B(n1329), .ZN(n1356) );
XNOR2_X1 U1097 ( .A(n1361), .B(G119), .ZN(n1329) );
INV_X1 U1098 ( .A(G116), .ZN(n1361) );
XOR2_X1 U1099 ( .A(n1130), .B(n1362), .Z(n1185) );
XNOR2_X1 U1100 ( .A(n1363), .B(KEYINPUT34), .ZN(n1362) );
NAND2_X1 U1101 ( .A1(KEYINPUT31), .A2(n1131), .ZN(n1363) );
INV_X1 U1102 ( .A(G131), .ZN(n1131) );
XNOR2_X1 U1103 ( .A(G134), .B(n1238), .ZN(n1130) );
INV_X1 U1104 ( .A(G137), .ZN(n1238) );
NAND2_X1 U1105 ( .A1(KEYINPUT20), .A2(n1172), .ZN(n1355) );
AND3_X1 U1106 ( .A1(n1291), .A2(n1067), .A3(G210), .ZN(n1172) );
INV_X1 U1107 ( .A(G953), .ZN(n1067) );
INV_X1 U1108 ( .A(G237), .ZN(n1291) );
XOR2_X1 U1109 ( .A(KEYINPUT12), .B(G101), .Z(n1353) );
endmodule


