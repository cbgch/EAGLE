//Key = 1111111000101011110001000100111110111011111010111010010100011100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412;

XNOR2_X1 U771 ( .A(n1072), .B(n1073), .ZN(G9) );
XNOR2_X1 U772 ( .A(KEYINPUT36), .B(n1074), .ZN(n1073) );
NOR2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR3_X1 U774 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
NAND3_X1 U775 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1077) );
NAND2_X1 U776 ( .A1(n1083), .A2(n1084), .ZN(n1080) );
NAND2_X1 U777 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND4_X1 U778 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1089) );
NAND2_X1 U780 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U782 ( .A1(n1097), .A2(n1098), .ZN(n1091) );
XNOR2_X1 U783 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND3_X1 U784 ( .A1(n1097), .A2(n1101), .A3(n1093), .ZN(n1085) );
NAND2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND3_X1 U786 ( .A1(n1104), .A2(n1105), .A3(n1088), .ZN(n1103) );
NAND2_X1 U787 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND3_X1 U788 ( .A1(n1108), .A2(n1109), .A3(n1090), .ZN(n1104) );
NAND2_X1 U789 ( .A1(n1087), .A2(n1110), .ZN(n1102) );
INV_X1 U790 ( .A(n1111), .ZN(n1083) );
AND3_X1 U791 ( .A1(n1112), .A2(n1081), .A3(n1082), .ZN(n1075) );
NAND4_X1 U792 ( .A1(n1113), .A2(n1097), .A3(n1093), .A4(n1114), .ZN(n1081) );
NOR4_X1 U793 ( .A1(n1115), .A2(n1106), .A3(n1116), .A4(n1117), .ZN(n1114) );
NOR2_X1 U794 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
INV_X1 U795 ( .A(n1120), .ZN(n1115) );
XNOR2_X1 U796 ( .A(KEYINPUT54), .B(G952), .ZN(n1112) );
XOR2_X1 U797 ( .A(n1121), .B(n1122), .Z(G72) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U800 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U801 ( .A(G953), .B(KEYINPUT50), .ZN(n1127) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1125) );
NOR2_X1 U803 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
NOR2_X1 U804 ( .A1(G140), .A2(n1133), .ZN(n1132) );
NOR2_X1 U805 ( .A1(KEYINPUT23), .A2(n1134), .ZN(n1133) );
NOR3_X1 U806 ( .A1(n1135), .A2(KEYINPUT23), .A3(n1136), .ZN(n1131) );
XNOR2_X1 U807 ( .A(KEYINPUT63), .B(n1137), .ZN(n1129) );
NOR2_X1 U808 ( .A1(KEYINPUT7), .A2(n1138), .ZN(n1137) );
XOR2_X1 U809 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U810 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U811 ( .A(G137), .B(n1143), .ZN(n1139) );
NAND2_X1 U812 ( .A1(KEYINPUT46), .A2(n1144), .ZN(n1143) );
NAND2_X1 U813 ( .A1(n1145), .A2(n1146), .ZN(n1123) );
NAND2_X1 U814 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XNOR2_X1 U815 ( .A(KEYINPUT4), .B(n1149), .ZN(n1145) );
NOR2_X1 U816 ( .A1(n1150), .A2(n1149), .ZN(n1121) );
AND2_X1 U817 ( .A1(G227), .A2(G900), .ZN(n1150) );
XOR2_X1 U818 ( .A(n1151), .B(n1152), .Z(G69) );
XOR2_X1 U819 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U820 ( .A1(n1155), .A2(G953), .ZN(n1154) );
NOR2_X1 U821 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
XOR2_X1 U822 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U823 ( .A1(KEYINPUT56), .A2(n1160), .ZN(n1158) );
NOR2_X1 U824 ( .A1(G898), .A2(n1149), .ZN(n1156) );
NOR2_X1 U825 ( .A1(n1161), .A2(n1149), .ZN(n1151) );
AND2_X1 U826 ( .A1(G224), .A2(G898), .ZN(n1161) );
NOR2_X1 U827 ( .A1(n1162), .A2(n1163), .ZN(G66) );
XOR2_X1 U828 ( .A(n1164), .B(n1165), .Z(n1163) );
NOR2_X1 U829 ( .A1(n1119), .A2(n1166), .ZN(n1164) );
NOR2_X1 U830 ( .A1(n1167), .A2(n1168), .ZN(G63) );
XOR2_X1 U831 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U832 ( .A(n1171), .B(KEYINPUT6), .Z(n1169) );
NAND2_X1 U833 ( .A1(n1172), .A2(G478), .ZN(n1171) );
NOR2_X1 U834 ( .A1(n1149), .A2(n1173), .ZN(n1167) );
XNOR2_X1 U835 ( .A(KEYINPUT33), .B(n1078), .ZN(n1173) );
INV_X1 U836 ( .A(G952), .ZN(n1078) );
NOR2_X1 U837 ( .A1(n1162), .A2(n1174), .ZN(G60) );
XOR2_X1 U838 ( .A(n1175), .B(n1176), .Z(n1174) );
AND2_X1 U839 ( .A1(G475), .A2(n1172), .ZN(n1175) );
XNOR2_X1 U840 ( .A(n1177), .B(n1178), .ZN(G6) );
NOR2_X1 U841 ( .A1(n1179), .A2(n1095), .ZN(n1178) );
NOR2_X1 U842 ( .A1(n1162), .A2(n1180), .ZN(G57) );
XOR2_X1 U843 ( .A(n1181), .B(n1182), .Z(n1180) );
NAND2_X1 U844 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
NAND2_X1 U845 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U846 ( .A1(n1172), .A2(G472), .ZN(n1186) );
XOR2_X1 U847 ( .A(n1187), .B(KEYINPUT24), .Z(n1183) );
NAND3_X1 U848 ( .A1(n1172), .A2(G472), .A3(n1188), .ZN(n1187) );
INV_X1 U849 ( .A(n1185), .ZN(n1188) );
XNOR2_X1 U850 ( .A(n1189), .B(n1190), .ZN(n1185) );
XNOR2_X1 U851 ( .A(n1191), .B(KEYINPUT44), .ZN(n1189) );
NOR2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(G54) );
XNOR2_X1 U853 ( .A(n1162), .B(KEYINPUT1), .ZN(n1193) );
XOR2_X1 U854 ( .A(n1194), .B(n1195), .Z(n1192) );
XOR2_X1 U855 ( .A(n1196), .B(n1197), .Z(n1195) );
NAND2_X1 U856 ( .A1(KEYINPUT60), .A2(n1198), .ZN(n1197) );
NAND2_X1 U857 ( .A1(KEYINPUT10), .A2(n1199), .ZN(n1196) );
XNOR2_X1 U858 ( .A(n1200), .B(G110), .ZN(n1199) );
INV_X1 U859 ( .A(G140), .ZN(n1200) );
XNOR2_X1 U860 ( .A(n1201), .B(n1202), .ZN(n1194) );
NOR2_X1 U861 ( .A1(KEYINPUT52), .A2(n1203), .ZN(n1202) );
AND2_X1 U862 ( .A1(G469), .A2(n1172), .ZN(n1203) );
INV_X1 U863 ( .A(n1166), .ZN(n1172) );
NOR2_X1 U864 ( .A1(n1162), .A2(n1204), .ZN(G51) );
XOR2_X1 U865 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U866 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR4_X1 U867 ( .A1(n1209), .A2(n1210), .A3(KEYINPUT27), .A4(n1166), .ZN(n1208) );
NAND2_X1 U868 ( .A1(n1211), .A2(n1079), .ZN(n1166) );
NAND3_X1 U869 ( .A1(n1147), .A2(n1212), .A3(n1155), .ZN(n1079) );
AND4_X1 U870 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1155) );
NOR4_X1 U871 ( .A1(n1217), .A2(n1218), .A3(n1072), .A4(n1219), .ZN(n1216) );
NOR2_X1 U872 ( .A1(n1096), .A2(n1179), .ZN(n1072) );
NAND3_X1 U873 ( .A1(n1220), .A2(n1221), .A3(n1087), .ZN(n1179) );
NOR3_X1 U874 ( .A1(n1222), .A2(n1223), .A3(n1224), .ZN(n1218) );
XNOR2_X1 U875 ( .A(n1225), .B(KEYINPUT62), .ZN(n1223) );
NOR4_X1 U876 ( .A1(n1226), .A2(n1107), .A3(n1095), .A4(n1227), .ZN(n1217) );
XNOR2_X1 U877 ( .A(KEYINPUT19), .B(n1221), .ZN(n1227) );
INV_X1 U878 ( .A(n1087), .ZN(n1107) );
NOR2_X1 U879 ( .A1(n1228), .A2(n1229), .ZN(n1215) );
XNOR2_X1 U880 ( .A(KEYINPUT0), .B(n1148), .ZN(n1212) );
AND4_X1 U881 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1147) );
NOR4_X1 U882 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1233) );
INV_X1 U883 ( .A(n1238), .ZN(n1236) );
NAND3_X1 U884 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1232) );
XNOR2_X1 U885 ( .A(G902), .B(KEYINPUT16), .ZN(n1211) );
NOR2_X1 U886 ( .A1(n1242), .A2(n1243), .ZN(n1210) );
INV_X1 U887 ( .A(KEYINPUT43), .ZN(n1243) );
AND3_X1 U888 ( .A1(G210), .A2(n1244), .A3(n1245), .ZN(n1242) );
NOR2_X1 U889 ( .A1(KEYINPUT43), .A2(n1246), .ZN(n1209) );
NOR2_X1 U890 ( .A1(n1149), .A2(G952), .ZN(n1162) );
NAND2_X1 U891 ( .A1(n1247), .A2(n1248), .ZN(G48) );
NAND2_X1 U892 ( .A1(G146), .A2(n1230), .ZN(n1248) );
XOR2_X1 U893 ( .A(KEYINPUT48), .B(n1249), .Z(n1247) );
NOR2_X1 U894 ( .A1(G146), .A2(n1230), .ZN(n1249) );
NAND4_X1 U895 ( .A1(n1225), .A2(n1250), .A3(n1220), .A4(n1251), .ZN(n1230) );
XNOR2_X1 U896 ( .A(G143), .B(n1231), .ZN(G45) );
NAND4_X1 U897 ( .A1(n1252), .A2(n1251), .A3(n1253), .A4(n1254), .ZN(n1231) );
NOR2_X1 U898 ( .A1(n1226), .A2(n1109), .ZN(n1254) );
XNOR2_X1 U899 ( .A(G140), .B(n1238), .ZN(G42) );
NAND3_X1 U900 ( .A1(n1255), .A2(n1250), .A3(n1241), .ZN(n1238) );
XOR2_X1 U901 ( .A(n1235), .B(n1256), .Z(G39) );
NOR2_X1 U902 ( .A1(KEYINPUT58), .A2(n1257), .ZN(n1256) );
AND3_X1 U903 ( .A1(n1225), .A2(n1097), .A3(n1241), .ZN(n1235) );
INV_X1 U904 ( .A(n1258), .ZN(n1225) );
XNOR2_X1 U905 ( .A(n1144), .B(n1259), .ZN(G36) );
NOR4_X1 U906 ( .A1(n1260), .A2(n1096), .A3(n1109), .A4(n1261), .ZN(n1259) );
XNOR2_X1 U907 ( .A(n1262), .B(KEYINPUT47), .ZN(n1260) );
XNOR2_X1 U908 ( .A(G131), .B(n1148), .ZN(G33) );
NAND3_X1 U909 ( .A1(n1250), .A2(n1239), .A3(n1241), .ZN(n1148) );
NOR2_X1 U910 ( .A1(n1261), .A2(n1262), .ZN(n1241) );
NAND4_X1 U911 ( .A1(n1088), .A2(n1100), .A3(n1090), .A4(n1099), .ZN(n1261) );
INV_X1 U912 ( .A(n1095), .ZN(n1250) );
NAND2_X1 U913 ( .A1(n1263), .A2(n1264), .ZN(G30) );
OR2_X1 U914 ( .A1(n1265), .A2(G128), .ZN(n1264) );
NAND2_X1 U915 ( .A1(G128), .A2(n1266), .ZN(n1263) );
NAND2_X1 U916 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U917 ( .A1(n1234), .A2(n1269), .ZN(n1268) );
INV_X1 U918 ( .A(KEYINPUT12), .ZN(n1269) );
NAND2_X1 U919 ( .A1(KEYINPUT12), .A2(n1265), .ZN(n1267) );
NAND2_X1 U920 ( .A1(KEYINPUT40), .A2(n1234), .ZN(n1265) );
NOR4_X1 U921 ( .A1(n1258), .A2(n1096), .A3(n1226), .A4(n1262), .ZN(n1234) );
INV_X1 U922 ( .A(n1251), .ZN(n1262) );
XNOR2_X1 U923 ( .A(G101), .B(n1213), .ZN(G3) );
NAND4_X1 U924 ( .A1(n1239), .A2(n1097), .A3(n1220), .A4(n1221), .ZN(n1213) );
INV_X1 U925 ( .A(n1109), .ZN(n1239) );
NAND3_X1 U926 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(G27) );
NAND2_X1 U927 ( .A1(KEYINPUT45), .A2(n1273), .ZN(n1272) );
OR3_X1 U928 ( .A1(n1273), .A2(KEYINPUT45), .A3(G125), .ZN(n1271) );
NAND2_X1 U929 ( .A1(G125), .A2(n1274), .ZN(n1270) );
NAND2_X1 U930 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
INV_X1 U931 ( .A(KEYINPUT45), .ZN(n1276) );
XNOR2_X1 U932 ( .A(n1237), .B(KEYINPUT28), .ZN(n1275) );
INV_X1 U933 ( .A(n1273), .ZN(n1237) );
NAND4_X1 U934 ( .A1(n1110), .A2(n1251), .A3(n1093), .A4(n1277), .ZN(n1273) );
NOR2_X1 U935 ( .A1(n1095), .A2(n1108), .ZN(n1277) );
INV_X1 U936 ( .A(n1255), .ZN(n1108) );
NAND2_X1 U937 ( .A1(n1111), .A2(n1278), .ZN(n1251) );
NAND4_X1 U938 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1128), .ZN(n1278) );
INV_X1 U939 ( .A(G900), .ZN(n1128) );
XNOR2_X1 U940 ( .A(G122), .B(n1214), .ZN(G24) );
NAND4_X1 U941 ( .A1(n1280), .A2(n1087), .A3(n1253), .A4(n1252), .ZN(n1214) );
NOR2_X1 U942 ( .A1(n1281), .A2(n1117), .ZN(n1087) );
INV_X1 U943 ( .A(n1222), .ZN(n1280) );
XNOR2_X1 U944 ( .A(G119), .B(n1282), .ZN(G21) );
NOR2_X1 U945 ( .A1(n1283), .A2(KEYINPUT11), .ZN(n1282) );
NOR3_X1 U946 ( .A1(n1258), .A2(n1224), .A3(n1222), .ZN(n1283) );
INV_X1 U947 ( .A(n1097), .ZN(n1224) );
NAND2_X1 U948 ( .A1(n1117), .A2(n1281), .ZN(n1258) );
NAND2_X1 U949 ( .A1(n1284), .A2(n1285), .ZN(G18) );
NAND2_X1 U950 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
INV_X1 U951 ( .A(n1229), .ZN(n1287) );
NAND2_X1 U952 ( .A1(n1288), .A2(n1289), .ZN(n1286) );
NAND2_X1 U953 ( .A1(KEYINPUT30), .A2(n1290), .ZN(n1289) );
INV_X1 U954 ( .A(KEYINPUT35), .ZN(n1290) );
NAND3_X1 U955 ( .A1(n1291), .A2(n1292), .A3(KEYINPUT35), .ZN(n1284) );
OR2_X1 U956 ( .A1(G116), .A2(KEYINPUT30), .ZN(n1292) );
NAND2_X1 U957 ( .A1(KEYINPUT30), .A2(n1293), .ZN(n1291) );
NAND2_X1 U958 ( .A1(n1229), .A2(n1288), .ZN(n1293) );
INV_X1 U959 ( .A(G116), .ZN(n1288) );
NOR3_X1 U960 ( .A1(n1222), .A2(n1096), .A3(n1109), .ZN(n1229) );
INV_X1 U961 ( .A(n1240), .ZN(n1096) );
NOR2_X1 U962 ( .A1(n1252), .A2(n1294), .ZN(n1240) );
XNOR2_X1 U963 ( .A(n1295), .B(n1228), .ZN(G15) );
NOR3_X1 U964 ( .A1(n1109), .A2(n1222), .A3(n1095), .ZN(n1228) );
NAND2_X1 U965 ( .A1(n1294), .A2(n1252), .ZN(n1095) );
INV_X1 U966 ( .A(n1253), .ZN(n1294) );
NAND3_X1 U967 ( .A1(n1110), .A2(n1221), .A3(n1093), .ZN(n1222) );
AND2_X1 U968 ( .A1(n1296), .A2(n1099), .ZN(n1093) );
INV_X1 U969 ( .A(n1100), .ZN(n1296) );
NAND2_X1 U970 ( .A1(n1297), .A2(n1117), .ZN(n1109) );
XOR2_X1 U971 ( .A(G110), .B(n1219), .Z(G12) );
AND4_X1 U972 ( .A1(n1255), .A2(n1097), .A3(n1220), .A4(n1221), .ZN(n1219) );
NAND2_X1 U973 ( .A1(n1111), .A2(n1298), .ZN(n1221) );
NAND4_X1 U974 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1299), .ZN(n1298) );
INV_X1 U975 ( .A(G898), .ZN(n1299) );
NAND3_X1 U976 ( .A1(n1082), .A2(n1279), .A3(G952), .ZN(n1111) );
NAND2_X1 U977 ( .A1(G237), .A2(G234), .ZN(n1279) );
XOR2_X1 U978 ( .A(G953), .B(KEYINPUT3), .Z(n1082) );
INV_X1 U979 ( .A(n1226), .ZN(n1220) );
NAND3_X1 U980 ( .A1(n1100), .A2(n1099), .A3(n1110), .ZN(n1226) );
NOR2_X1 U981 ( .A1(n1088), .A2(n1106), .ZN(n1110) );
INV_X1 U982 ( .A(n1090), .ZN(n1106) );
NAND2_X1 U983 ( .A1(G214), .A2(n1300), .ZN(n1090) );
XNOR2_X1 U984 ( .A(n1113), .B(KEYINPUT41), .ZN(n1088) );
XOR2_X1 U985 ( .A(n1301), .B(n1246), .Z(n1113) );
AND2_X1 U986 ( .A1(G210), .A2(n1300), .ZN(n1246) );
NAND2_X1 U987 ( .A1(n1245), .A2(n1244), .ZN(n1300) );
INV_X1 U988 ( .A(G237), .ZN(n1245) );
NAND2_X1 U989 ( .A1(n1302), .A2(n1244), .ZN(n1301) );
XOR2_X1 U990 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U991 ( .A(n1205), .B(KEYINPUT61), .Z(n1304) );
XOR2_X1 U992 ( .A(n1305), .B(n1306), .Z(n1205) );
XOR2_X1 U993 ( .A(n1159), .B(n1160), .Z(n1306) );
XOR2_X1 U994 ( .A(G110), .B(n1307), .Z(n1160) );
NOR2_X1 U995 ( .A1(KEYINPUT22), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U996 ( .A(n1309), .B(n1310), .ZN(n1159) );
XOR2_X1 U997 ( .A(n1311), .B(n1312), .Z(n1310) );
NAND2_X1 U998 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
NAND2_X1 U999 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1000 ( .A1(G104), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1001 ( .A(G101), .B(G107), .ZN(n1315) );
NAND2_X1 U1002 ( .A1(n1318), .A2(n1317), .ZN(n1313) );
INV_X1 U1003 ( .A(KEYINPUT26), .ZN(n1317) );
NAND2_X1 U1004 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
XNOR2_X1 U1005 ( .A(G113), .B(KEYINPUT21), .ZN(n1309) );
XOR2_X1 U1006 ( .A(n1321), .B(KEYINPUT18), .Z(n1305) );
NAND2_X1 U1007 ( .A1(G224), .A2(n1149), .ZN(n1321) );
NAND2_X1 U1008 ( .A1(n1322), .A2(n1323), .ZN(n1303) );
NAND2_X1 U1009 ( .A1(KEYINPUT55), .A2(n1207), .ZN(n1323) );
XNOR2_X1 U1010 ( .A(n1324), .B(n1325), .ZN(n1207) );
NAND3_X1 U1011 ( .A1(n1325), .A2(n1135), .A3(n1326), .ZN(n1322) );
INV_X1 U1012 ( .A(KEYINPUT55), .ZN(n1326) );
XNOR2_X1 U1013 ( .A(n1327), .B(G128), .ZN(n1325) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1328), .ZN(n1099) );
XNOR2_X1 U1015 ( .A(n1329), .B(G469), .ZN(n1100) );
NAND3_X1 U1016 ( .A1(n1330), .A2(n1331), .A3(n1244), .ZN(n1329) );
NAND2_X1 U1017 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
XNOR2_X1 U1018 ( .A(n1334), .B(n1198), .ZN(n1332) );
NAND2_X1 U1019 ( .A1(KEYINPUT42), .A2(n1335), .ZN(n1334) );
NAND2_X1 U1020 ( .A1(n1336), .A2(n1201), .ZN(n1330) );
INV_X1 U1021 ( .A(n1333), .ZN(n1201) );
NAND2_X1 U1022 ( .A1(G227), .A2(n1149), .ZN(n1333) );
XNOR2_X1 U1023 ( .A(n1337), .B(n1198), .ZN(n1336) );
XNOR2_X1 U1024 ( .A(n1338), .B(n1339), .ZN(n1198) );
XOR2_X1 U1025 ( .A(n1340), .B(n1141), .Z(n1338) );
XNOR2_X1 U1026 ( .A(n1341), .B(n1342), .ZN(n1141) );
XNOR2_X1 U1027 ( .A(n1343), .B(KEYINPUT59), .ZN(n1342) );
NAND2_X1 U1028 ( .A1(KEYINPUT29), .A2(n1344), .ZN(n1343) );
NAND4_X1 U1029 ( .A1(n1320), .A2(n1319), .A3(n1345), .A4(n1346), .ZN(n1340) );
NAND3_X1 U1030 ( .A1(n1347), .A2(n1177), .A3(n1074), .ZN(n1346) );
NAND3_X1 U1031 ( .A1(G101), .A2(n1177), .A3(G107), .ZN(n1345) );
INV_X1 U1032 ( .A(G104), .ZN(n1177) );
NAND3_X1 U1033 ( .A1(G104), .A2(n1347), .A3(G107), .ZN(n1319) );
INV_X1 U1034 ( .A(G101), .ZN(n1347) );
NAND3_X1 U1035 ( .A1(G104), .A2(n1074), .A3(G101), .ZN(n1320) );
NAND2_X1 U1036 ( .A1(n1348), .A2(KEYINPUT42), .ZN(n1337) );
XOR2_X1 U1037 ( .A(n1335), .B(KEYINPUT53), .Z(n1348) );
XNOR2_X1 U1038 ( .A(G110), .B(n1349), .ZN(n1335) );
NOR2_X1 U1039 ( .A1(KEYINPUT9), .A2(n1350), .ZN(n1349) );
XNOR2_X1 U1040 ( .A(G140), .B(KEYINPUT38), .ZN(n1350) );
NOR2_X1 U1041 ( .A1(n1253), .A2(n1252), .ZN(n1097) );
XOR2_X1 U1042 ( .A(G475), .B(n1351), .Z(n1252) );
NOR2_X1 U1043 ( .A1(n1176), .A2(n1352), .ZN(n1351) );
XNOR2_X1 U1044 ( .A(KEYINPUT49), .B(n1244), .ZN(n1352) );
XNOR2_X1 U1045 ( .A(n1353), .B(n1354), .ZN(n1176) );
XOR2_X1 U1046 ( .A(n1355), .B(n1356), .Z(n1354) );
NOR2_X1 U1047 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
XOR2_X1 U1048 ( .A(KEYINPUT13), .B(n1359), .Z(n1358) );
AND2_X1 U1049 ( .A1(n1344), .A2(n1360), .ZN(n1359) );
NOR2_X1 U1050 ( .A1(n1360), .A2(n1344), .ZN(n1357) );
NAND2_X1 U1051 ( .A1(n1134), .A2(n1361), .ZN(n1360) );
NAND2_X1 U1052 ( .A1(G140), .A2(n1135), .ZN(n1361) );
INV_X1 U1053 ( .A(n1136), .ZN(n1134) );
NOR2_X1 U1054 ( .A1(KEYINPUT20), .A2(n1362), .ZN(n1355) );
XOR2_X1 U1055 ( .A(n1363), .B(n1364), .Z(n1362) );
XNOR2_X1 U1056 ( .A(G122), .B(G104), .ZN(n1364) );
NAND2_X1 U1057 ( .A1(KEYINPUT15), .A2(n1295), .ZN(n1363) );
INV_X1 U1058 ( .A(G113), .ZN(n1295) );
NAND2_X1 U1059 ( .A1(KEYINPUT17), .A2(n1365), .ZN(n1353) );
XNOR2_X1 U1060 ( .A(n1366), .B(n1367), .ZN(n1365) );
XOR2_X1 U1061 ( .A(n1368), .B(G131), .Z(n1367) );
NAND2_X1 U1062 ( .A1(G214), .A2(n1369), .ZN(n1368) );
XNOR2_X1 U1063 ( .A(n1370), .B(G478), .ZN(n1253) );
OR2_X1 U1064 ( .A1(n1170), .A2(G902), .ZN(n1370) );
XNOR2_X1 U1065 ( .A(n1371), .B(n1372), .ZN(n1170) );
XOR2_X1 U1066 ( .A(n1373), .B(n1374), .Z(n1372) );
XNOR2_X1 U1067 ( .A(n1308), .B(G116), .ZN(n1374) );
INV_X1 U1068 ( .A(G122), .ZN(n1308) );
XNOR2_X1 U1069 ( .A(n1144), .B(G128), .ZN(n1373) );
INV_X1 U1070 ( .A(G134), .ZN(n1144) );
XNOR2_X1 U1071 ( .A(n1375), .B(n1341), .ZN(n1371) );
XNOR2_X1 U1072 ( .A(n1376), .B(n1074), .ZN(n1375) );
INV_X1 U1073 ( .A(G107), .ZN(n1074) );
NAND2_X1 U1074 ( .A1(G217), .A2(n1377), .ZN(n1376) );
NOR2_X1 U1075 ( .A1(n1117), .A2(n1297), .ZN(n1255) );
INV_X1 U1076 ( .A(n1281), .ZN(n1297) );
NAND3_X1 U1077 ( .A1(n1378), .A2(n1379), .A3(n1120), .ZN(n1281) );
NAND2_X1 U1078 ( .A1(n1118), .A2(n1119), .ZN(n1120) );
NAND2_X1 U1079 ( .A1(n1119), .A2(n1380), .ZN(n1379) );
OR3_X1 U1080 ( .A1(n1119), .A2(n1118), .A3(n1380), .ZN(n1378) );
INV_X1 U1081 ( .A(KEYINPUT32), .ZN(n1380) );
NOR2_X1 U1082 ( .A1(n1165), .A2(G902), .ZN(n1118) );
XNOR2_X1 U1083 ( .A(n1381), .B(n1382), .ZN(n1165) );
AND2_X1 U1084 ( .A1(n1377), .A2(G221), .ZN(n1382) );
AND2_X1 U1085 ( .A1(G234), .A2(n1149), .ZN(n1377) );
INV_X1 U1086 ( .A(G953), .ZN(n1149) );
XNOR2_X1 U1087 ( .A(n1383), .B(n1257), .ZN(n1381) );
INV_X1 U1088 ( .A(G137), .ZN(n1257) );
NAND2_X1 U1089 ( .A1(n1384), .A2(n1385), .ZN(n1383) );
NAND2_X1 U1090 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
XOR2_X1 U1091 ( .A(KEYINPUT2), .B(n1388), .Z(n1384) );
NOR2_X1 U1092 ( .A1(n1386), .A2(n1387), .ZN(n1388) );
XOR2_X1 U1093 ( .A(G110), .B(n1389), .Z(n1387) );
XNOR2_X1 U1094 ( .A(n1390), .B(G119), .ZN(n1389) );
XNOR2_X1 U1095 ( .A(n1391), .B(n1344), .ZN(n1386) );
NAND2_X1 U1096 ( .A1(n1392), .A2(n1393), .ZN(n1391) );
NAND2_X1 U1097 ( .A1(G140), .A2(n1394), .ZN(n1393) );
NAND2_X1 U1098 ( .A1(n1324), .A2(n1395), .ZN(n1394) );
NAND2_X1 U1099 ( .A1(n1136), .A2(n1395), .ZN(n1392) );
INV_X1 U1100 ( .A(KEYINPUT8), .ZN(n1395) );
NOR2_X1 U1101 ( .A1(n1135), .A2(G140), .ZN(n1136) );
INV_X1 U1102 ( .A(n1324), .ZN(n1135) );
XOR2_X1 U1103 ( .A(G125), .B(KEYINPUT31), .Z(n1324) );
NAND2_X1 U1104 ( .A1(G217), .A2(n1328), .ZN(n1119) );
NAND2_X1 U1105 ( .A1(G234), .A2(n1244), .ZN(n1328) );
XNOR2_X1 U1106 ( .A(n1396), .B(G472), .ZN(n1117) );
NAND2_X1 U1107 ( .A1(n1397), .A2(n1244), .ZN(n1396) );
INV_X1 U1108 ( .A(G902), .ZN(n1244) );
XOR2_X1 U1109 ( .A(n1398), .B(n1182), .Z(n1397) );
XNOR2_X1 U1110 ( .A(n1399), .B(G101), .ZN(n1182) );
NAND2_X1 U1111 ( .A1(G210), .A2(n1369), .ZN(n1399) );
NOR2_X1 U1112 ( .A1(G953), .A2(G237), .ZN(n1369) );
NAND3_X1 U1113 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n1398) );
OR2_X1 U1114 ( .A1(n1403), .A2(KEYINPUT14), .ZN(n1402) );
INV_X1 U1115 ( .A(n1191), .ZN(n1403) );
NAND3_X1 U1116 ( .A1(KEYINPUT14), .A2(n1404), .A3(n1190), .ZN(n1401) );
OR2_X1 U1117 ( .A1(n1190), .A2(n1404), .ZN(n1400) );
NOR2_X1 U1118 ( .A1(KEYINPUT37), .A2(n1191), .ZN(n1404) );
XNOR2_X1 U1119 ( .A(n1405), .B(n1406), .ZN(n1191) );
NOR2_X1 U1120 ( .A1(KEYINPUT51), .A2(n1312), .ZN(n1406) );
XNOR2_X1 U1121 ( .A(G119), .B(G116), .ZN(n1312) );
XNOR2_X1 U1122 ( .A(G113), .B(KEYINPUT25), .ZN(n1405) );
XNOR2_X1 U1123 ( .A(n1327), .B(n1339), .ZN(n1190) );
XNOR2_X1 U1124 ( .A(n1407), .B(n1142), .ZN(n1339) );
XNOR2_X1 U1125 ( .A(G131), .B(n1390), .ZN(n1142) );
INV_X1 U1126 ( .A(G128), .ZN(n1390) );
NAND2_X1 U1127 ( .A1(KEYINPUT5), .A2(n1408), .ZN(n1407) );
XNOR2_X1 U1128 ( .A(G134), .B(n1409), .ZN(n1408) );
NAND2_X1 U1129 ( .A1(KEYINPUT39), .A2(G137), .ZN(n1409) );
NAND2_X1 U1130 ( .A1(n1410), .A2(n1411), .ZN(n1327) );
NAND2_X1 U1131 ( .A1(G146), .A2(n1366), .ZN(n1411) );
XOR2_X1 U1132 ( .A(n1412), .B(KEYINPUT57), .Z(n1410) );
NAND2_X1 U1133 ( .A1(n1341), .A2(n1344), .ZN(n1412) );
INV_X1 U1134 ( .A(G146), .ZN(n1344) );
INV_X1 U1135 ( .A(n1366), .ZN(n1341) );
XOR2_X1 U1136 ( .A(G143), .B(KEYINPUT34), .Z(n1366) );
endmodule


