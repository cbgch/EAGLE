//Key = 1100011110110000111110000101101000000100110001000110010000100001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;

XOR2_X1 U745 ( .A(G107), .B(n1024), .Z(G9) );
NOR2_X1 U746 ( .A1(KEYINPUT47), .A2(n1025), .ZN(n1024) );
NOR2_X1 U747 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR4_X1 U748 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
XOR2_X1 U749 ( .A(KEYINPUT2), .B(n1032), .Z(n1029) );
AND4_X1 U750 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
NAND4_X1 U751 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1028) );
NAND4_X1 U752 ( .A1(n1041), .A2(n1042), .A3(n1034), .A4(n1043), .ZN(n1038) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1035), .A2(n1046), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
INV_X1 U757 ( .A(n1051), .ZN(n1047) );
NAND2_X1 U758 ( .A1(n1052), .A2(n1053), .ZN(n1044) );
NAND2_X1 U759 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
INV_X1 U761 ( .A(n1058), .ZN(n1041) );
NAND2_X1 U762 ( .A1(n1035), .A2(n1059), .ZN(n1037) );
NAND2_X1 U763 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U764 ( .A1(n1036), .A2(n1062), .ZN(n1061) );
NAND2_X1 U765 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U766 ( .A1(n1034), .A2(n1065), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1042), .A2(n1066), .ZN(n1063) );
XOR2_X1 U768 ( .A(n1067), .B(KEYINPUT15), .Z(n1060) );
NAND4_X1 U769 ( .A1(n1036), .A2(n1042), .A3(n1068), .A4(n1069), .ZN(n1067) );
NAND2_X1 U770 ( .A1(KEYINPUT48), .A2(n1070), .ZN(n1069) );
NAND2_X1 U771 ( .A1(n1071), .A2(n1072), .ZN(n1068) );
INV_X1 U772 ( .A(KEYINPUT48), .ZN(n1072) );
NAND2_X1 U773 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U774 ( .A1(n1058), .A2(n1075), .ZN(n1036) );
NOR3_X1 U775 ( .A1(n1076), .A2(G953), .A3(G952), .ZN(n1026) );
INV_X1 U776 ( .A(n1039), .ZN(n1076) );
NAND4_X1 U777 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1039) );
NOR4_X1 U778 ( .A1(n1081), .A2(n1082), .A3(n1075), .A4(n1083), .ZN(n1080) );
XOR2_X1 U779 ( .A(KEYINPUT59), .B(n1084), .Z(n1083) );
NOR2_X1 U780 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR3_X1 U781 ( .A1(n1056), .A2(n1087), .A3(n1073), .ZN(n1079) );
NAND2_X1 U782 ( .A1(n1088), .A2(n1089), .ZN(n1078) );
NAND2_X1 U783 ( .A1(n1085), .A2(n1086), .ZN(n1077) );
NAND2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(G72) );
NAND2_X1 U785 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U786 ( .A1(G953), .A2(n1094), .ZN(n1093) );
NAND3_X1 U787 ( .A1(G953), .A2(n1095), .A3(n1096), .ZN(n1090) );
INV_X1 U788 ( .A(n1092), .ZN(n1096) );
NOR2_X1 U789 ( .A1(KEYINPUT36), .A2(n1097), .ZN(n1092) );
XOR2_X1 U790 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR3_X1 U791 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
XNOR2_X1 U793 ( .A(n1105), .B(n1106), .ZN(n1104) );
XOR2_X1 U794 ( .A(KEYINPUT54), .B(n1107), .Z(n1100) );
NOR2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U796 ( .A(n1105), .B(n1110), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(n1105) );
OR2_X1 U798 ( .A1(n1113), .A2(KEYINPUT38), .ZN(n1112) );
NAND3_X1 U799 ( .A1(G131), .A2(n1114), .A3(KEYINPUT38), .ZN(n1111) );
NAND2_X1 U800 ( .A1(n1040), .A2(n1031), .ZN(n1098) );
NAND2_X1 U801 ( .A1(G900), .A2(G227), .ZN(n1095) );
XOR2_X1 U802 ( .A(n1115), .B(n1116), .Z(G69) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1040), .ZN(n1116) );
NOR2_X1 U804 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U805 ( .A1(n1120), .A2(n1121), .ZN(n1115) );
OR3_X1 U806 ( .A1(n1122), .A2(G953), .A3(n1123), .ZN(n1121) );
NAND2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
NAND2_X1 U808 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U809 ( .A1(n1122), .A2(n1040), .ZN(n1126) );
INV_X1 U810 ( .A(n1030), .ZN(n1122) );
NAND2_X1 U811 ( .A1(n1127), .A2(G953), .ZN(n1125) );
XNOR2_X1 U812 ( .A(KEYINPUT24), .B(n1119), .ZN(n1127) );
NOR2_X1 U813 ( .A1(KEYINPUT35), .A2(n1128), .ZN(n1123) );
NOR2_X1 U814 ( .A1(n1129), .A2(n1130), .ZN(G66) );
XNOR2_X1 U815 ( .A(n1131), .B(n1132), .ZN(n1130) );
NOR2_X1 U816 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U817 ( .A1(n1129), .A2(n1135), .ZN(G63) );
NOR3_X1 U818 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
NOR2_X1 U819 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U820 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
XOR2_X1 U821 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U822 ( .A(KEYINPUT31), .B(KEYINPUT19), .Z(n1144) );
INV_X1 U823 ( .A(KEYINPUT49), .ZN(n1141) );
AND3_X1 U824 ( .A1(n1140), .A2(n1143), .A3(KEYINPUT49), .ZN(n1137) );
NAND2_X1 U825 ( .A1(n1145), .A2(G478), .ZN(n1140) );
NOR2_X1 U826 ( .A1(KEYINPUT49), .A2(n1143), .ZN(n1136) );
NOR2_X1 U827 ( .A1(n1129), .A2(n1146), .ZN(G60) );
NOR3_X1 U828 ( .A1(n1147), .A2(n1148), .A3(n1149), .ZN(n1146) );
NOR2_X1 U829 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NOR2_X1 U830 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
XNOR2_X1 U831 ( .A(KEYINPUT51), .B(n1154), .ZN(n1153) );
INV_X1 U832 ( .A(KEYINPUT30), .ZN(n1152) );
AND3_X1 U833 ( .A1(n1151), .A2(n1154), .A3(KEYINPUT30), .ZN(n1148) );
NOR2_X1 U834 ( .A1(KEYINPUT30), .A2(n1154), .ZN(n1147) );
NAND2_X1 U835 ( .A1(n1145), .A2(G475), .ZN(n1154) );
XOR2_X1 U836 ( .A(G104), .B(n1155), .Z(G6) );
NOR2_X1 U837 ( .A1(n1129), .A2(n1156), .ZN(G57) );
XOR2_X1 U838 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U839 ( .A(n1113), .B(n1159), .ZN(n1158) );
XOR2_X1 U840 ( .A(n1160), .B(n1161), .Z(n1157) );
AND2_X1 U841 ( .A1(G472), .A2(n1145), .ZN(n1161) );
INV_X1 U842 ( .A(n1134), .ZN(n1145) );
XNOR2_X1 U843 ( .A(n1162), .B(n1163), .ZN(n1160) );
NOR2_X1 U844 ( .A1(KEYINPUT32), .A2(n1164), .ZN(n1163) );
NOR2_X1 U845 ( .A1(KEYINPUT4), .A2(n1165), .ZN(n1162) );
XOR2_X1 U846 ( .A(n1166), .B(KEYINPUT37), .Z(n1165) );
NOR2_X1 U847 ( .A1(n1129), .A2(n1167), .ZN(G54) );
XOR2_X1 U848 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U849 ( .A(n1170), .B(n1171), .Z(n1169) );
NOR2_X1 U850 ( .A1(n1086), .A2(n1134), .ZN(n1171) );
NOR2_X1 U851 ( .A1(n1172), .A2(n1173), .ZN(n1170) );
NOR2_X1 U852 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U853 ( .A1(n1129), .A2(n1176), .ZN(G51) );
XOR2_X1 U854 ( .A(n1177), .B(n1178), .Z(n1176) );
NOR2_X1 U855 ( .A1(n1179), .A2(n1134), .ZN(n1178) );
NAND2_X1 U856 ( .A1(G902), .A2(n1180), .ZN(n1134) );
OR2_X1 U857 ( .A1(n1031), .A2(n1030), .ZN(n1180) );
NAND2_X1 U858 ( .A1(n1181), .A2(n1182), .ZN(n1030) );
AND4_X1 U859 ( .A1(n1183), .A2(n1184), .A3(n1025), .A4(n1185), .ZN(n1182) );
NAND3_X1 U860 ( .A1(n1052), .A2(n1186), .A3(n1065), .ZN(n1025) );
NOR4_X1 U861 ( .A1(n1187), .A2(n1155), .A3(n1188), .A4(n1189), .ZN(n1181) );
NOR2_X1 U862 ( .A1(n1054), .A2(n1190), .ZN(n1189) );
NOR3_X1 U863 ( .A1(n1191), .A2(n1075), .A3(n1192), .ZN(n1188) );
INV_X1 U864 ( .A(n1052), .ZN(n1075) );
AND3_X1 U865 ( .A1(n1052), .A2(n1186), .A3(n1033), .ZN(n1155) );
NAND2_X1 U866 ( .A1(n1193), .A2(n1194), .ZN(n1031) );
NOR4_X1 U867 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NOR4_X1 U868 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1193) );
NOR2_X1 U869 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
INV_X1 U870 ( .A(KEYINPUT45), .ZN(n1204) );
NOR2_X1 U871 ( .A1(n1205), .A2(n1206), .ZN(n1201) );
NOR2_X1 U872 ( .A1(n1207), .A2(n1208), .ZN(n1205) );
AND2_X1 U873 ( .A1(n1065), .A2(n1209), .ZN(n1208) );
NOR3_X1 U874 ( .A1(n1210), .A2(KEYINPUT45), .A3(n1066), .ZN(n1207) );
NOR2_X1 U875 ( .A1(n1211), .A2(n1212), .ZN(n1177) );
XOR2_X1 U876 ( .A(n1213), .B(KEYINPUT16), .Z(n1212) );
NAND2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NOR2_X1 U878 ( .A1(n1215), .A2(n1214), .ZN(n1211) );
XOR2_X1 U879 ( .A(KEYINPUT60), .B(n1216), .Z(n1214) );
NOR2_X1 U880 ( .A1(n1040), .A2(G952), .ZN(n1129) );
XNOR2_X1 U881 ( .A(n1217), .B(n1199), .ZN(G48) );
AND3_X1 U882 ( .A1(n1033), .A2(n1218), .A3(n1219), .ZN(n1199) );
XOR2_X1 U883 ( .A(n1198), .B(n1220), .Z(G45) );
XOR2_X1 U884 ( .A(KEYINPUT33), .B(G143), .Z(n1220) );
NOR3_X1 U885 ( .A1(n1221), .A2(n1054), .A3(n1192), .ZN(n1198) );
XNOR2_X1 U886 ( .A(G140), .B(n1203), .ZN(G42) );
NAND3_X1 U887 ( .A1(n1222), .A2(n1066), .A3(n1035), .ZN(n1203) );
INV_X1 U888 ( .A(n1210), .ZN(n1222) );
XOR2_X1 U889 ( .A(n1197), .B(n1223), .Z(G39) );
NOR2_X1 U890 ( .A1(KEYINPUT46), .A2(n1224), .ZN(n1223) );
AND3_X1 U891 ( .A1(n1035), .A2(n1219), .A3(n1042), .ZN(n1197) );
XNOR2_X1 U892 ( .A(G134), .B(n1225), .ZN(G36) );
NAND3_X1 U893 ( .A1(n1065), .A2(n1226), .A3(n1209), .ZN(n1225) );
INV_X1 U894 ( .A(n1221), .ZN(n1209) );
XNOR2_X1 U895 ( .A(KEYINPUT29), .B(n1206), .ZN(n1226) );
XOR2_X1 U896 ( .A(G131), .B(n1200), .Z(G33) );
NOR3_X1 U897 ( .A1(n1206), .A2(n1227), .A3(n1221), .ZN(n1200) );
NAND3_X1 U898 ( .A1(n1066), .A2(n1228), .A3(n1051), .ZN(n1221) );
INV_X1 U899 ( .A(n1035), .ZN(n1206) );
NOR2_X1 U900 ( .A1(n1229), .A2(n1056), .ZN(n1035) );
XNOR2_X1 U901 ( .A(n1230), .B(n1196), .ZN(G30) );
AND3_X1 U902 ( .A1(n1065), .A2(n1218), .A3(n1219), .ZN(n1196) );
AND4_X1 U903 ( .A1(n1066), .A2(n1231), .A3(n1050), .A4(n1228), .ZN(n1219) );
XOR2_X1 U904 ( .A(G101), .B(n1232), .Z(G3) );
NOR2_X1 U905 ( .A1(n1233), .A2(n1054), .ZN(n1232) );
XOR2_X1 U906 ( .A(n1190), .B(KEYINPUT43), .Z(n1233) );
NAND4_X1 U907 ( .A1(n1051), .A2(n1042), .A3(n1066), .A4(n1234), .ZN(n1190) );
XNOR2_X1 U908 ( .A(n1235), .B(n1195), .ZN(G27) );
NOR3_X1 U909 ( .A1(n1210), .A2(n1054), .A3(n1070), .ZN(n1195) );
INV_X1 U910 ( .A(n1218), .ZN(n1054) );
NAND4_X1 U911 ( .A1(n1049), .A2(n1033), .A3(n1050), .A4(n1228), .ZN(n1210) );
NAND2_X1 U912 ( .A1(n1058), .A2(n1236), .ZN(n1228) );
NAND3_X1 U913 ( .A1(n1237), .A2(n1238), .A3(n1102), .ZN(n1236) );
NOR2_X1 U914 ( .A1(n1040), .A2(G900), .ZN(n1102) );
XOR2_X1 U915 ( .A(KEYINPUT23), .B(n1239), .Z(n1237) );
XNOR2_X1 U916 ( .A(G122), .B(n1240), .ZN(G24) );
NAND3_X1 U917 ( .A1(n1052), .A2(n1241), .A3(n1242), .ZN(n1240) );
XNOR2_X1 U918 ( .A(KEYINPUT44), .B(n1192), .ZN(n1241) );
NAND2_X1 U919 ( .A1(n1243), .A2(n1082), .ZN(n1192) );
NOR2_X1 U920 ( .A1(n1050), .A2(n1231), .ZN(n1052) );
XOR2_X1 U921 ( .A(n1187), .B(n1244), .Z(G21) );
NOR2_X1 U922 ( .A1(KEYINPUT3), .A2(n1245), .ZN(n1244) );
AND4_X1 U923 ( .A1(n1242), .A2(n1042), .A3(n1231), .A4(n1050), .ZN(n1187) );
XOR2_X1 U924 ( .A(n1184), .B(n1246), .Z(G18) );
NAND2_X1 U925 ( .A1(KEYINPUT10), .A2(G116), .ZN(n1246) );
NAND3_X1 U926 ( .A1(n1051), .A2(n1065), .A3(n1242), .ZN(n1184) );
NOR2_X1 U927 ( .A1(n1082), .A2(n1247), .ZN(n1065) );
XOR2_X1 U928 ( .A(n1183), .B(n1248), .Z(G15) );
NOR2_X1 U929 ( .A1(G113), .A2(KEYINPUT56), .ZN(n1248) );
NAND3_X1 U930 ( .A1(n1051), .A2(n1033), .A3(n1242), .ZN(n1183) );
INV_X1 U931 ( .A(n1191), .ZN(n1242) );
NAND3_X1 U932 ( .A1(n1218), .A2(n1234), .A3(n1034), .ZN(n1191) );
INV_X1 U933 ( .A(n1070), .ZN(n1034) );
NAND2_X1 U934 ( .A1(n1074), .A2(n1249), .ZN(n1070) );
INV_X1 U935 ( .A(n1227), .ZN(n1033) );
NAND2_X1 U936 ( .A1(n1247), .A2(n1082), .ZN(n1227) );
NOR2_X1 U937 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
XNOR2_X1 U938 ( .A(G110), .B(n1185), .ZN(G12) );
NAND4_X1 U939 ( .A1(n1042), .A2(n1186), .A3(n1049), .A4(n1050), .ZN(n1185) );
XOR2_X1 U940 ( .A(n1250), .B(n1133), .Z(n1050) );
NAND2_X1 U941 ( .A1(G217), .A2(n1251), .ZN(n1133) );
NAND2_X1 U942 ( .A1(n1131), .A2(n1252), .ZN(n1250) );
XNOR2_X1 U943 ( .A(n1253), .B(n1254), .ZN(n1131) );
XOR2_X1 U944 ( .A(G110), .B(n1255), .Z(n1254) );
XNOR2_X1 U945 ( .A(n1230), .B(G119), .ZN(n1255) );
XOR2_X1 U946 ( .A(n1256), .B(n1257), .Z(n1253) );
NOR2_X1 U947 ( .A1(G137), .A2(KEYINPUT13), .ZN(n1257) );
XOR2_X1 U948 ( .A(n1258), .B(n1259), .Z(n1256) );
NOR2_X1 U949 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
INV_X1 U950 ( .A(G221), .ZN(n1261) );
NAND3_X1 U951 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1258) );
NAND2_X1 U952 ( .A1(KEYINPUT34), .A2(n1103), .ZN(n1264) );
NAND3_X1 U953 ( .A1(n1265), .A2(n1266), .A3(n1217), .ZN(n1263) );
INV_X1 U954 ( .A(KEYINPUT34), .ZN(n1266) );
OR2_X1 U955 ( .A1(n1217), .A2(n1265), .ZN(n1262) );
NOR2_X1 U956 ( .A1(KEYINPUT62), .A2(n1103), .ZN(n1265) );
INV_X1 U957 ( .A(n1108), .ZN(n1103) );
XOR2_X1 U958 ( .A(G125), .B(G140), .Z(n1108) );
INV_X1 U959 ( .A(n1231), .ZN(n1049) );
XNOR2_X1 U960 ( .A(n1267), .B(G472), .ZN(n1231) );
NAND2_X1 U961 ( .A1(n1268), .A2(n1252), .ZN(n1267) );
XOR2_X1 U962 ( .A(n1269), .B(n1159), .Z(n1268) );
XNOR2_X1 U963 ( .A(n1270), .B(G101), .ZN(n1159) );
NAND2_X1 U964 ( .A1(G210), .A2(n1271), .ZN(n1270) );
XOR2_X1 U965 ( .A(n1166), .B(n1272), .Z(n1269) );
NOR2_X1 U966 ( .A1(KEYINPUT42), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U967 ( .A(n1164), .B(n1113), .ZN(n1273) );
INV_X1 U968 ( .A(n1274), .ZN(n1113) );
XOR2_X1 U969 ( .A(n1275), .B(n1276), .Z(n1166) );
XOR2_X1 U970 ( .A(n1277), .B(KEYINPUT14), .Z(n1275) );
NAND3_X1 U971 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
OR2_X1 U972 ( .A1(G119), .A2(KEYINPUT58), .ZN(n1280) );
NAND3_X1 U973 ( .A1(KEYINPUT58), .A2(G119), .A3(n1281), .ZN(n1279) );
NAND2_X1 U974 ( .A1(n1282), .A2(n1283), .ZN(n1278) );
NAND2_X1 U975 ( .A1(KEYINPUT58), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U976 ( .A(KEYINPUT9), .B(n1245), .ZN(n1284) );
INV_X1 U977 ( .A(G119), .ZN(n1245) );
AND3_X1 U978 ( .A1(n1218), .A2(n1234), .A3(n1066), .ZN(n1186) );
NOR2_X1 U979 ( .A1(n1074), .A2(n1073), .ZN(n1066) );
INV_X1 U980 ( .A(n1249), .ZN(n1073) );
NAND2_X1 U981 ( .A1(G221), .A2(n1251), .ZN(n1249) );
NAND2_X1 U982 ( .A1(G234), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U983 ( .A(n1085), .B(n1285), .ZN(n1074) );
XNOR2_X1 U984 ( .A(KEYINPUT12), .B(n1086), .ZN(n1285) );
INV_X1 U985 ( .A(G469), .ZN(n1086) );
AND2_X1 U986 ( .A1(n1286), .A2(n1252), .ZN(n1085) );
XNOR2_X1 U987 ( .A(n1168), .B(n1287), .ZN(n1286) );
NOR2_X1 U988 ( .A1(n1172), .A2(n1288), .ZN(n1287) );
NOR2_X1 U989 ( .A1(n1175), .A2(n1289), .ZN(n1288) );
XNOR2_X1 U990 ( .A(n1174), .B(KEYINPUT41), .ZN(n1289) );
AND2_X1 U991 ( .A1(n1174), .A2(n1175), .ZN(n1172) );
XNOR2_X1 U992 ( .A(G110), .B(G140), .ZN(n1175) );
NOR2_X1 U993 ( .A1(n1094), .A2(G953), .ZN(n1174) );
INV_X1 U994 ( .A(G227), .ZN(n1094) );
XNOR2_X1 U995 ( .A(n1290), .B(n1291), .ZN(n1168) );
XOR2_X1 U996 ( .A(n1292), .B(n1293), .Z(n1291) );
XOR2_X1 U997 ( .A(KEYINPUT8), .B(KEYINPUT0), .Z(n1293) );
XNOR2_X1 U998 ( .A(n1294), .B(n1110), .ZN(n1290) );
INV_X1 U999 ( .A(n1106), .ZN(n1110) );
XOR2_X1 U1000 ( .A(n1295), .B(n1296), .Z(n1106) );
XNOR2_X1 U1001 ( .A(G146), .B(KEYINPUT63), .ZN(n1295) );
XNOR2_X1 U1002 ( .A(n1274), .B(n1297), .ZN(n1294) );
XOR2_X1 U1003 ( .A(G131), .B(n1114), .Z(n1274) );
XNOR2_X1 U1004 ( .A(n1224), .B(G134), .ZN(n1114) );
INV_X1 U1005 ( .A(G137), .ZN(n1224) );
NAND2_X1 U1006 ( .A1(n1058), .A2(n1298), .ZN(n1234) );
NAND4_X1 U1007 ( .A1(G953), .A2(n1239), .A3(n1238), .A4(n1119), .ZN(n1298) );
INV_X1 U1008 ( .A(G898), .ZN(n1119) );
XNOR2_X1 U1009 ( .A(n1252), .B(KEYINPUT52), .ZN(n1239) );
NAND3_X1 U1010 ( .A1(n1238), .A2(n1040), .A3(G952), .ZN(n1058) );
NAND2_X1 U1011 ( .A1(G237), .A2(G234), .ZN(n1238) );
NOR2_X1 U1012 ( .A1(n1056), .A2(n1057), .ZN(n1218) );
INV_X1 U1013 ( .A(n1229), .ZN(n1057) );
NAND3_X1 U1014 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1229) );
INV_X1 U1015 ( .A(n1087), .ZN(n1301) );
NOR2_X1 U1016 ( .A1(n1089), .A2(n1088), .ZN(n1087) );
NAND2_X1 U1017 ( .A1(KEYINPUT55), .A2(n1179), .ZN(n1300) );
NAND3_X1 U1018 ( .A1(n1089), .A2(n1302), .A3(n1088), .ZN(n1299) );
INV_X1 U1019 ( .A(n1179), .ZN(n1088) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1303), .ZN(n1179) );
INV_X1 U1021 ( .A(KEYINPUT55), .ZN(n1302) );
NAND2_X1 U1022 ( .A1(n1304), .A2(n1252), .ZN(n1089) );
XNOR2_X1 U1023 ( .A(n1216), .B(n1305), .ZN(n1304) );
XNOR2_X1 U1024 ( .A(n1215), .B(KEYINPUT25), .ZN(n1305) );
XNOR2_X1 U1025 ( .A(n1128), .B(KEYINPUT53), .ZN(n1215) );
XOR2_X1 U1026 ( .A(n1306), .B(n1307), .Z(n1128) );
XOR2_X1 U1027 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1028 ( .A(G119), .B(n1310), .ZN(n1309) );
NOR2_X1 U1029 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XOR2_X1 U1030 ( .A(n1313), .B(KEYINPUT6), .Z(n1312) );
NAND2_X1 U1031 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XOR2_X1 U1032 ( .A(KEYINPUT39), .B(G110), .Z(n1314) );
NOR2_X1 U1033 ( .A1(G110), .A2(n1315), .ZN(n1311) );
NAND2_X1 U1034 ( .A1(KEYINPUT18), .A2(n1292), .ZN(n1308) );
XOR2_X1 U1035 ( .A(G101), .B(KEYINPUT11), .Z(n1292) );
XNOR2_X1 U1036 ( .A(n1297), .B(n1316), .ZN(n1306) );
XNOR2_X1 U1037 ( .A(n1276), .B(n1282), .ZN(n1316) );
XNOR2_X1 U1038 ( .A(n1317), .B(KEYINPUT22), .ZN(n1276) );
XOR2_X1 U1039 ( .A(G104), .B(G107), .Z(n1297) );
XNOR2_X1 U1040 ( .A(n1318), .B(n1164), .ZN(n1216) );
XNOR2_X1 U1041 ( .A(n1319), .B(n1320), .ZN(n1164) );
XNOR2_X1 U1042 ( .A(G143), .B(n1321), .ZN(n1320) );
NAND2_X1 U1043 ( .A1(KEYINPUT50), .A2(G146), .ZN(n1321) );
NAND2_X1 U1044 ( .A1(KEYINPUT5), .A2(n1230), .ZN(n1319) );
XNOR2_X1 U1045 ( .A(G125), .B(n1322), .ZN(n1318) );
NOR2_X1 U1046 ( .A1(G953), .A2(n1118), .ZN(n1322) );
INV_X1 U1047 ( .A(G224), .ZN(n1118) );
AND2_X1 U1048 ( .A1(G214), .A2(n1303), .ZN(n1056) );
NAND2_X1 U1049 ( .A1(n1323), .A2(n1252), .ZN(n1303) );
INV_X1 U1050 ( .A(G237), .ZN(n1323) );
NOR2_X1 U1051 ( .A1(n1082), .A2(n1243), .ZN(n1042) );
INV_X1 U1052 ( .A(n1247), .ZN(n1243) );
XOR2_X1 U1053 ( .A(n1081), .B(KEYINPUT40), .Z(n1247) );
XNOR2_X1 U1054 ( .A(n1324), .B(G478), .ZN(n1081) );
NAND2_X1 U1055 ( .A1(n1143), .A2(n1252), .ZN(n1324) );
XNOR2_X1 U1056 ( .A(n1325), .B(n1326), .ZN(n1143) );
XOR2_X1 U1057 ( .A(G107), .B(n1327), .Z(n1326) );
XNOR2_X1 U1058 ( .A(KEYINPUT7), .B(n1315), .ZN(n1327) );
XNOR2_X1 U1059 ( .A(n1328), .B(n1282), .ZN(n1325) );
INV_X1 U1060 ( .A(n1281), .ZN(n1282) );
XOR2_X1 U1061 ( .A(G116), .B(KEYINPUT27), .Z(n1281) );
XOR2_X1 U1062 ( .A(n1329), .B(n1330), .Z(n1328) );
NOR2_X1 U1063 ( .A1(n1260), .A2(n1331), .ZN(n1330) );
INV_X1 U1064 ( .A(G217), .ZN(n1331) );
NAND2_X1 U1065 ( .A1(G234), .A2(n1040), .ZN(n1260) );
INV_X1 U1066 ( .A(G953), .ZN(n1040) );
NAND2_X1 U1067 ( .A1(n1332), .A2(n1333), .ZN(n1329) );
NAND2_X1 U1068 ( .A1(n1296), .A2(n1334), .ZN(n1333) );
XOR2_X1 U1069 ( .A(KEYINPUT17), .B(n1335), .Z(n1332) );
NOR2_X1 U1070 ( .A1(n1296), .A2(n1334), .ZN(n1335) );
INV_X1 U1071 ( .A(G134), .ZN(n1334) );
XOR2_X1 U1072 ( .A(n1230), .B(G143), .Z(n1296) );
INV_X1 U1073 ( .A(G128), .ZN(n1230) );
XNOR2_X1 U1074 ( .A(n1336), .B(G475), .ZN(n1082) );
NAND2_X1 U1075 ( .A1(n1151), .A2(n1252), .ZN(n1336) );
INV_X1 U1076 ( .A(G902), .ZN(n1252) );
XNOR2_X1 U1077 ( .A(n1337), .B(n1338), .ZN(n1151) );
XOR2_X1 U1078 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1079 ( .A(n1341), .B(n1342), .Z(n1340) );
NAND2_X1 U1080 ( .A1(KEYINPUT1), .A2(n1235), .ZN(n1342) );
INV_X1 U1081 ( .A(G125), .ZN(n1235) );
NAND2_X1 U1082 ( .A1(n1343), .A2(KEYINPUT28), .ZN(n1341) );
XOR2_X1 U1083 ( .A(n1344), .B(G143), .Z(n1343) );
NAND2_X1 U1084 ( .A1(G214), .A2(n1271), .ZN(n1344) );
NOR2_X1 U1085 ( .A1(G953), .A2(G237), .ZN(n1271) );
NOR2_X1 U1086 ( .A1(G104), .A2(KEYINPUT61), .ZN(n1339) );
XOR2_X1 U1087 ( .A(n1345), .B(n1346), .Z(n1337) );
XNOR2_X1 U1088 ( .A(n1217), .B(G140), .ZN(n1346) );
INV_X1 U1089 ( .A(G146), .ZN(n1217) );
XOR2_X1 U1090 ( .A(n1347), .B(G131), .Z(n1345) );
NAND3_X1 U1091 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1347) );
NAND2_X1 U1092 ( .A1(n1317), .A2(n1351), .ZN(n1350) );
NAND3_X1 U1093 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1351) );
NAND2_X1 U1094 ( .A1(KEYINPUT26), .A2(n1355), .ZN(n1354) );
OR2_X1 U1095 ( .A1(G122), .A2(KEYINPUT20), .ZN(n1353) );
NAND2_X1 U1096 ( .A1(KEYINPUT20), .A2(n1356), .ZN(n1352) );
NAND2_X1 U1097 ( .A1(n1315), .A2(n1357), .ZN(n1356) );
NAND2_X1 U1098 ( .A1(KEYINPUT57), .A2(n1358), .ZN(n1357) );
INV_X1 U1099 ( .A(n1359), .ZN(n1317) );
NAND4_X1 U1100 ( .A1(n1315), .A2(n1355), .A3(n1359), .A4(n1358), .ZN(n1349) );
INV_X1 U1101 ( .A(KEYINPUT26), .ZN(n1358) );
INV_X1 U1102 ( .A(KEYINPUT57), .ZN(n1355) );
NAND2_X1 U1103 ( .A1(KEYINPUT26), .A2(n1360), .ZN(n1348) );
NAND2_X1 U1104 ( .A1(n1315), .A2(n1361), .ZN(n1360) );
NAND2_X1 U1105 ( .A1(KEYINPUT57), .A2(n1359), .ZN(n1361) );
XOR2_X1 U1106 ( .A(G113), .B(KEYINPUT21), .Z(n1359) );
INV_X1 U1107 ( .A(G122), .ZN(n1315) );
endmodule


