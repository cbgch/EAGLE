//Key = 1000110100001001100111010000100010011001110010101111101000110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U734 ( .A(G107), .B(n1024), .ZN(G9) );
NAND2_X1 U735 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
XOR2_X1 U736 ( .A(n1027), .B(KEYINPUT15), .Z(n1025) );
NOR2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U738 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
NAND3_X1 U739 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1030) );
NAND2_X1 U740 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND4_X1 U742 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1040) );
NOR2_X1 U743 ( .A1(n1045), .A2(n1046), .ZN(n1041) );
NOR3_X1 U744 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NOR2_X1 U745 ( .A1(n1050), .A2(n1051), .ZN(n1045) );
NOR2_X1 U746 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NAND3_X1 U747 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1039) );
NAND2_X1 U748 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND3_X1 U749 ( .A1(n1059), .A2(n1051), .A3(n1042), .ZN(n1058) );
NAND2_X1 U750 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U751 ( .A1(n1043), .A2(n1062), .ZN(n1061) );
NAND2_X1 U752 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1065), .ZN(n1060) );
NAND3_X1 U754 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
OR3_X1 U755 ( .A1(n1069), .A2(n1070), .A3(KEYINPUT61), .ZN(n1067) );
NAND2_X1 U756 ( .A1(KEYINPUT61), .A2(n1043), .ZN(n1066) );
NAND2_X1 U757 ( .A1(n1071), .A2(n1044), .ZN(n1057) );
INV_X1 U758 ( .A(n1072), .ZN(n1037) );
NOR3_X1 U759 ( .A1(n1073), .A2(G953), .A3(n1074), .ZN(n1028) );
INV_X1 U760 ( .A(n1034), .ZN(n1074) );
NAND4_X1 U761 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1034) );
NOR4_X1 U762 ( .A1(n1052), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1078) );
XOR2_X1 U763 ( .A(KEYINPUT5), .B(n1082), .Z(n1081) );
NOR2_X1 U764 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U765 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U766 ( .A(n1087), .B(KEYINPUT21), .Z(n1085) );
XOR2_X1 U767 ( .A(n1088), .B(n1089), .Z(n1080) );
NOR2_X1 U768 ( .A1(KEYINPUT9), .A2(n1090), .ZN(n1089) );
NOR3_X1 U769 ( .A1(n1091), .A2(n1092), .A3(n1047), .ZN(n1077) );
NAND2_X1 U770 ( .A1(n1093), .A2(n1094), .ZN(n1076) );
XNOR2_X1 U771 ( .A(KEYINPUT13), .B(n1032), .ZN(n1073) );
XOR2_X1 U772 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U773 ( .A(n1097), .B(n1098), .Z(n1096) );
NOR2_X1 U774 ( .A1(n1099), .A2(n1035), .ZN(n1098) );
NOR2_X1 U775 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
XNOR2_X1 U776 ( .A(G900), .B(KEYINPUT56), .ZN(n1100) );
NAND2_X1 U777 ( .A1(n1102), .A2(n1103), .ZN(n1097) );
NAND2_X1 U778 ( .A1(G953), .A2(n1104), .ZN(n1103) );
XOR2_X1 U779 ( .A(n1105), .B(n1106), .Z(n1102) );
XOR2_X1 U780 ( .A(n1107), .B(n1108), .Z(n1106) );
NAND2_X1 U781 ( .A1(KEYINPUT44), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U782 ( .A(G140), .B(n1110), .ZN(n1109) );
NAND2_X1 U783 ( .A1(KEYINPUT52), .A2(G125), .ZN(n1110) );
XOR2_X1 U784 ( .A(n1111), .B(G137), .Z(n1105) );
NAND2_X1 U785 ( .A1(n1035), .A2(n1033), .ZN(n1095) );
NAND2_X1 U786 ( .A1(n1112), .A2(n1113), .ZN(G69) );
OR2_X1 U787 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U788 ( .A(n1116), .B(KEYINPUT38), .Z(n1112) );
NAND2_X1 U789 ( .A1(n1115), .A2(n1114), .ZN(n1116) );
NAND2_X1 U790 ( .A1(n1117), .A2(G953), .ZN(n1114) );
XOR2_X1 U791 ( .A(n1118), .B(KEYINPUT55), .Z(n1117) );
NAND2_X1 U792 ( .A1(G898), .A2(G224), .ZN(n1118) );
XNOR2_X1 U793 ( .A(n1119), .B(n1120), .ZN(n1115) );
NOR2_X1 U794 ( .A1(G953), .A2(n1121), .ZN(n1120) );
XOR2_X1 U795 ( .A(n1031), .B(KEYINPUT23), .Z(n1121) );
NAND2_X1 U796 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
INV_X1 U797 ( .A(n1124), .ZN(n1123) );
XOR2_X1 U798 ( .A(n1125), .B(n1126), .Z(n1122) );
NOR2_X1 U799 ( .A1(KEYINPUT30), .A2(n1127), .ZN(n1125) );
NOR3_X1 U800 ( .A1(n1128), .A2(n1129), .A3(n1130), .ZN(G66) );
AND2_X1 U801 ( .A1(KEYINPUT49), .A2(n1131), .ZN(n1130) );
NOR3_X1 U802 ( .A1(KEYINPUT49), .A2(n1035), .A3(n1032), .ZN(n1129) );
INV_X1 U803 ( .A(G952), .ZN(n1032) );
XOR2_X1 U804 ( .A(n1132), .B(n1133), .Z(n1128) );
NAND2_X1 U805 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NOR2_X1 U806 ( .A1(n1131), .A2(n1136), .ZN(G63) );
XOR2_X1 U807 ( .A(n1137), .B(n1138), .Z(n1136) );
AND2_X1 U808 ( .A1(G478), .A2(n1134), .ZN(n1137) );
NOR2_X1 U809 ( .A1(n1131), .A2(n1139), .ZN(G60) );
XOR2_X1 U810 ( .A(KEYINPUT47), .B(n1140), .Z(n1139) );
NOR2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U812 ( .A(KEYINPUT17), .B(n1143), .Z(n1142) );
NOR2_X1 U813 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U814 ( .A(KEYINPUT29), .B(n1146), .Z(n1145) );
AND2_X1 U815 ( .A1(n1144), .A2(n1146), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1147), .A2(n1090), .ZN(n1144) );
XOR2_X1 U817 ( .A(n1148), .B(n1149), .Z(G6) );
NAND2_X1 U818 ( .A1(KEYINPUT19), .A2(G104), .ZN(n1149) );
NOR2_X1 U819 ( .A1(n1131), .A2(n1150), .ZN(G57) );
XOR2_X1 U820 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U821 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U822 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U823 ( .A1(n1086), .A2(n1147), .ZN(n1155) );
NOR3_X1 U824 ( .A1(n1147), .A2(n1157), .A3(n1086), .ZN(n1153) );
INV_X1 U825 ( .A(G472), .ZN(n1086) );
XOR2_X1 U826 ( .A(n1156), .B(KEYINPUT48), .Z(n1157) );
NAND2_X1 U827 ( .A1(KEYINPUT32), .A2(n1158), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1131), .A2(n1159), .ZN(G54) );
XOR2_X1 U829 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U830 ( .A1(n1134), .A2(G469), .ZN(n1160) );
INV_X1 U831 ( .A(n1147), .ZN(n1134) );
NOR2_X1 U832 ( .A1(n1131), .A2(n1162), .ZN(G51) );
XOR2_X1 U833 ( .A(n1163), .B(n1164), .Z(n1162) );
NOR2_X1 U834 ( .A1(n1094), .A2(n1147), .ZN(n1164) );
NAND2_X1 U835 ( .A1(G902), .A2(n1165), .ZN(n1147) );
OR2_X1 U836 ( .A1(n1031), .A2(n1033), .ZN(n1165) );
NAND2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1033) );
NOR4_X1 U838 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NOR4_X1 U839 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1166) );
NOR3_X1 U840 ( .A1(n1176), .A2(n1177), .A3(n1063), .ZN(n1175) );
NOR4_X1 U841 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1174) );
XNOR2_X1 U842 ( .A(n1182), .B(KEYINPUT53), .ZN(n1180) );
NAND4_X1 U843 ( .A1(n1183), .A2(n1148), .A3(n1184), .A4(n1185), .ZN(n1031) );
AND3_X1 U844 ( .A1(n1186), .A2(n1187), .A3(n1188), .ZN(n1185) );
NAND2_X1 U845 ( .A1(n1189), .A2(n1190), .ZN(n1184) );
NAND2_X1 U846 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NAND2_X1 U847 ( .A1(n1071), .A2(n1193), .ZN(n1192) );
NAND3_X1 U848 ( .A1(n1194), .A2(n1195), .A3(n1048), .ZN(n1191) );
NAND2_X1 U849 ( .A1(KEYINPUT54), .A2(n1181), .ZN(n1195) );
NAND2_X1 U850 ( .A1(n1196), .A2(n1197), .ZN(n1194) );
INV_X1 U851 ( .A(KEYINPUT54), .ZN(n1197) );
NAND2_X1 U852 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
NAND3_X1 U853 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1148) );
NAND2_X1 U854 ( .A1(n1026), .A2(n1203), .ZN(n1183) );
NAND2_X1 U855 ( .A1(n1204), .A2(n1027), .ZN(n1203) );
NAND3_X1 U856 ( .A1(n1198), .A2(n1201), .A3(n1182), .ZN(n1027) );
NOR2_X1 U857 ( .A1(n1205), .A2(n1206), .ZN(n1163) );
XOR2_X1 U858 ( .A(KEYINPUT31), .B(n1207), .Z(n1206) );
NOR2_X1 U859 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XOR2_X1 U860 ( .A(n1210), .B(KEYINPUT1), .Z(n1208) );
AND2_X1 U861 ( .A1(n1209), .A2(n1210), .ZN(n1205) );
XOR2_X1 U862 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U863 ( .A(G125), .B(n1213), .Z(n1212) );
NAND2_X1 U864 ( .A1(n1214), .A2(n1215), .ZN(n1211) );
XOR2_X1 U865 ( .A(KEYINPUT46), .B(KEYINPUT10), .Z(n1214) );
NOR2_X1 U866 ( .A1(n1035), .A2(G952), .ZN(n1131) );
XNOR2_X1 U867 ( .A(n1173), .B(n1216), .ZN(G48) );
NOR2_X1 U868 ( .A1(G146), .A2(KEYINPUT11), .ZN(n1216) );
NOR4_X1 U869 ( .A1(n1063), .A2(n1181), .A3(n1179), .A4(n1178), .ZN(n1173) );
INV_X1 U870 ( .A(n1193), .ZN(n1179) );
NAND2_X1 U871 ( .A1(n1217), .A2(n1218), .ZN(G45) );
NAND2_X1 U872 ( .A1(n1171), .A2(n1219), .ZN(n1218) );
XOR2_X1 U873 ( .A(KEYINPUT39), .B(n1220), .Z(n1217) );
NOR2_X1 U874 ( .A1(n1171), .A2(n1219), .ZN(n1220) );
AND3_X1 U875 ( .A1(n1221), .A2(n1048), .A3(n1222), .ZN(n1171) );
NOR3_X1 U876 ( .A1(n1181), .A2(n1178), .A3(n1223), .ZN(n1222) );
INV_X1 U877 ( .A(n1224), .ZN(n1178) );
INV_X1 U878 ( .A(n1200), .ZN(n1181) );
XOR2_X1 U879 ( .A(n1170), .B(n1225), .Z(G42) );
XNOR2_X1 U880 ( .A(KEYINPUT60), .B(n1226), .ZN(n1225) );
AND3_X1 U881 ( .A1(n1202), .A2(n1049), .A3(n1227), .ZN(n1170) );
XOR2_X1 U882 ( .A(G137), .B(n1169), .Z(G39) );
AND3_X1 U883 ( .A1(n1044), .A2(n1193), .A3(n1227), .ZN(n1169) );
INV_X1 U884 ( .A(n1176), .ZN(n1227) );
XOR2_X1 U885 ( .A(G134), .B(n1168), .Z(G36) );
NOR3_X1 U886 ( .A1(n1177), .A2(n1064), .A3(n1176), .ZN(n1168) );
INV_X1 U887 ( .A(n1182), .ZN(n1064) );
XOR2_X1 U888 ( .A(G131), .B(n1228), .Z(G33) );
NOR4_X1 U889 ( .A1(KEYINPUT22), .A2(n1177), .A3(n1063), .A4(n1176), .ZN(n1228) );
NAND4_X1 U890 ( .A1(n1042), .A2(n1198), .A3(n1224), .A4(n1051), .ZN(n1176) );
INV_X1 U891 ( .A(n1068), .ZN(n1198) );
XNOR2_X1 U892 ( .A(G128), .B(n1229), .ZN(G30) );
NAND4_X1 U893 ( .A1(n1200), .A2(n1182), .A3(n1230), .A4(n1193), .ZN(n1229) );
XNOR2_X1 U894 ( .A(KEYINPUT28), .B(n1224), .ZN(n1230) );
XNOR2_X1 U895 ( .A(G101), .B(n1231), .ZN(G3) );
NAND2_X1 U896 ( .A1(n1048), .A2(n1232), .ZN(n1231) );
XOR2_X1 U897 ( .A(G125), .B(n1172), .Z(G27) );
AND4_X1 U898 ( .A1(n1202), .A2(n1071), .A3(n1049), .A4(n1224), .ZN(n1172) );
NAND2_X1 U899 ( .A1(n1072), .A2(n1233), .ZN(n1224) );
NAND4_X1 U900 ( .A1(G902), .A2(G953), .A3(n1234), .A4(n1104), .ZN(n1233) );
INV_X1 U901 ( .A(G900), .ZN(n1104) );
XNOR2_X1 U902 ( .A(G122), .B(n1186), .ZN(G24) );
NAND4_X1 U903 ( .A1(n1221), .A2(n1071), .A3(n1201), .A4(n1235), .ZN(n1186) );
AND3_X1 U904 ( .A1(n1054), .A2(n1236), .A3(n1056), .ZN(n1201) );
INV_X1 U905 ( .A(n1052), .ZN(n1054) );
AND2_X1 U906 ( .A1(n1043), .A2(n1026), .ZN(n1071) );
XNOR2_X1 U907 ( .A(G119), .B(n1237), .ZN(G21) );
NAND4_X1 U908 ( .A1(n1043), .A2(n1189), .A3(n1238), .A4(n1193), .ZN(n1237) );
NAND2_X1 U909 ( .A1(n1239), .A2(n1240), .ZN(n1193) );
OR2_X1 U910 ( .A1(n1177), .A2(KEYINPUT35), .ZN(n1240) );
INV_X1 U911 ( .A(n1048), .ZN(n1177) );
NAND3_X1 U912 ( .A1(n1052), .A2(n1053), .A3(KEYINPUT35), .ZN(n1239) );
INV_X1 U913 ( .A(n1056), .ZN(n1053) );
XNOR2_X1 U914 ( .A(KEYINPUT26), .B(n1199), .ZN(n1238) );
XNOR2_X1 U915 ( .A(G116), .B(n1188), .ZN(G18) );
NAND3_X1 U916 ( .A1(n1026), .A2(n1182), .A3(n1241), .ZN(n1188) );
NOR2_X1 U917 ( .A1(n1221), .A2(n1223), .ZN(n1182) );
XOR2_X1 U918 ( .A(n1242), .B(n1243), .Z(G15) );
NOR2_X1 U919 ( .A1(KEYINPUT37), .A2(n1244), .ZN(n1243) );
NOR2_X1 U920 ( .A1(n1245), .A2(n1199), .ZN(n1242) );
XOR2_X1 U921 ( .A(n1204), .B(KEYINPUT57), .Z(n1245) );
NAND2_X1 U922 ( .A1(n1202), .A2(n1241), .ZN(n1204) );
AND3_X1 U923 ( .A1(n1048), .A2(n1236), .A3(n1043), .ZN(n1241) );
NOR2_X1 U924 ( .A1(n1070), .A2(n1091), .ZN(n1043) );
NOR2_X1 U925 ( .A1(n1052), .A2(n1056), .ZN(n1048) );
INV_X1 U926 ( .A(n1063), .ZN(n1202) );
NAND2_X1 U927 ( .A1(n1246), .A2(n1223), .ZN(n1063) );
INV_X1 U928 ( .A(n1235), .ZN(n1223) );
XNOR2_X1 U929 ( .A(n1247), .B(KEYINPUT43), .ZN(n1246) );
XNOR2_X1 U930 ( .A(G110), .B(n1187), .ZN(G12) );
NAND2_X1 U931 ( .A1(n1049), .A2(n1232), .ZN(n1187) );
AND2_X1 U932 ( .A1(n1200), .A2(n1189), .ZN(n1232) );
AND2_X1 U933 ( .A1(n1044), .A2(n1236), .ZN(n1189) );
NAND2_X1 U934 ( .A1(n1072), .A2(n1248), .ZN(n1236) );
NAND3_X1 U935 ( .A1(n1124), .A2(n1234), .A3(G902), .ZN(n1248) );
NOR2_X1 U936 ( .A1(n1035), .A2(G898), .ZN(n1124) );
NAND3_X1 U937 ( .A1(n1234), .A2(n1035), .A3(G952), .ZN(n1072) );
NAND2_X1 U938 ( .A1(G237), .A2(G234), .ZN(n1234) );
NOR2_X1 U939 ( .A1(n1235), .A2(n1221), .ZN(n1044) );
INV_X1 U940 ( .A(n1247), .ZN(n1221) );
XOR2_X1 U941 ( .A(n1088), .B(n1249), .Z(n1247) );
XNOR2_X1 U942 ( .A(KEYINPUT41), .B(n1090), .ZN(n1249) );
INV_X1 U943 ( .A(G475), .ZN(n1090) );
NOR2_X1 U944 ( .A1(n1146), .A2(G902), .ZN(n1088) );
AND2_X1 U945 ( .A1(n1250), .A2(n1251), .ZN(n1146) );
NAND2_X1 U946 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U947 ( .A(n1254), .ZN(n1253) );
XNOR2_X1 U948 ( .A(n1255), .B(n1256), .ZN(n1252) );
XOR2_X1 U949 ( .A(n1257), .B(KEYINPUT2), .Z(n1250) );
NAND2_X1 U950 ( .A1(n1258), .A2(n1254), .ZN(n1257) );
XNOR2_X1 U951 ( .A(n1259), .B(n1260), .ZN(n1254) );
XNOR2_X1 U952 ( .A(n1244), .B(G104), .ZN(n1260) );
XOR2_X1 U953 ( .A(n1261), .B(G122), .Z(n1259) );
XNOR2_X1 U954 ( .A(KEYINPUT42), .B(KEYINPUT33), .ZN(n1261) );
XNOR2_X1 U955 ( .A(n1256), .B(n1262), .ZN(n1258) );
INV_X1 U956 ( .A(n1255), .ZN(n1262) );
XOR2_X1 U957 ( .A(G131), .B(n1263), .Z(n1255) );
XNOR2_X1 U958 ( .A(n1219), .B(G140), .ZN(n1263) );
XNOR2_X1 U959 ( .A(n1264), .B(n1265), .ZN(n1256) );
XOR2_X1 U960 ( .A(G125), .B(n1266), .Z(n1265) );
NOR2_X1 U961 ( .A1(KEYINPUT63), .A2(n1267), .ZN(n1266) );
NAND2_X1 U962 ( .A1(n1268), .A2(G214), .ZN(n1264) );
XNOR2_X1 U963 ( .A(n1075), .B(KEYINPUT27), .ZN(n1235) );
XNOR2_X1 U964 ( .A(G478), .B(n1269), .ZN(n1075) );
NOR2_X1 U965 ( .A1(G902), .A2(n1138), .ZN(n1269) );
XNOR2_X1 U966 ( .A(n1270), .B(n1271), .ZN(n1138) );
XNOR2_X1 U967 ( .A(n1272), .B(n1273), .ZN(n1271) );
XNOR2_X1 U968 ( .A(n1219), .B(G134), .ZN(n1273) );
XOR2_X1 U969 ( .A(n1274), .B(n1275), .Z(n1270) );
NOR2_X1 U970 ( .A1(KEYINPUT8), .A2(n1276), .ZN(n1275) );
XOR2_X1 U971 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U972 ( .A(G116), .B(G107), .Z(n1278) );
XOR2_X1 U973 ( .A(KEYINPUT3), .B(G122), .Z(n1277) );
NAND2_X1 U974 ( .A1(G217), .A2(n1279), .ZN(n1274) );
NOR2_X1 U975 ( .A1(n1199), .A2(n1068), .ZN(n1200) );
NAND2_X1 U976 ( .A1(n1280), .A2(n1070), .ZN(n1068) );
XOR2_X1 U977 ( .A(n1079), .B(KEYINPUT34), .Z(n1070) );
XNOR2_X1 U978 ( .A(n1281), .B(G469), .ZN(n1079) );
NAND2_X1 U979 ( .A1(n1161), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U980 ( .A(n1283), .B(n1284), .ZN(n1161) );
XNOR2_X1 U981 ( .A(n1285), .B(n1286), .ZN(n1284) );
XNOR2_X1 U982 ( .A(n1287), .B(n1288), .ZN(n1286) );
XOR2_X1 U983 ( .A(n1289), .B(n1290), .Z(n1283) );
XNOR2_X1 U984 ( .A(KEYINPUT36), .B(n1291), .ZN(n1290) );
XOR2_X1 U985 ( .A(n1111), .B(n1292), .Z(n1289) );
NOR2_X1 U986 ( .A1(G953), .A2(n1101), .ZN(n1292) );
INV_X1 U987 ( .A(G227), .ZN(n1101) );
NAND2_X1 U988 ( .A1(n1293), .A2(n1294), .ZN(n1111) );
NAND2_X1 U989 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XOR2_X1 U990 ( .A(n1297), .B(KEYINPUT20), .Z(n1295) );
XNOR2_X1 U991 ( .A(n1091), .B(KEYINPUT6), .ZN(n1280) );
INV_X1 U992 ( .A(n1069), .ZN(n1091) );
NAND2_X1 U993 ( .A1(G221), .A2(n1298), .ZN(n1069) );
INV_X1 U994 ( .A(n1026), .ZN(n1199) );
NOR2_X1 U995 ( .A1(n1047), .A2(n1042), .ZN(n1026) );
NOR2_X1 U996 ( .A1(n1299), .A2(n1092), .ZN(n1042) );
NOR2_X1 U997 ( .A1(n1094), .A2(n1093), .ZN(n1092) );
XNOR2_X1 U998 ( .A(KEYINPUT4), .B(n1300), .ZN(n1299) );
NOR2_X1 U999 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
XOR2_X1 U1000 ( .A(KEYINPUT12), .B(n1093), .Z(n1302) );
AND3_X1 U1001 ( .A1(n1303), .A2(n1282), .A3(n1304), .ZN(n1093) );
XOR2_X1 U1002 ( .A(n1305), .B(KEYINPUT62), .Z(n1304) );
NAND2_X1 U1003 ( .A1(n1209), .A2(n1306), .ZN(n1305) );
OR2_X1 U1004 ( .A1(n1306), .A2(n1209), .ZN(n1303) );
XNOR2_X1 U1005 ( .A(n1127), .B(n1126), .ZN(n1209) );
XNOR2_X1 U1006 ( .A(n1307), .B(G122), .ZN(n1126) );
INV_X1 U1007 ( .A(G110), .ZN(n1307) );
XOR2_X1 U1008 ( .A(n1308), .B(n1285), .Z(n1127) );
XNOR2_X1 U1009 ( .A(G107), .B(n1309), .ZN(n1285) );
XOR2_X1 U1010 ( .A(n1310), .B(n1311), .Z(n1308) );
NAND2_X1 U1011 ( .A1(KEYINPUT7), .A2(n1291), .ZN(n1310) );
INV_X1 U1012 ( .A(G104), .ZN(n1291) );
XNOR2_X1 U1013 ( .A(n1312), .B(n1313), .ZN(n1306) );
XOR2_X1 U1014 ( .A(KEYINPUT51), .B(n1213), .Z(n1313) );
AND2_X1 U1015 ( .A1(G224), .A2(n1035), .ZN(n1213) );
NAND2_X1 U1016 ( .A1(n1314), .A2(KEYINPUT50), .ZN(n1312) );
XOR2_X1 U1017 ( .A(n1215), .B(n1315), .Z(n1314) );
XOR2_X1 U1018 ( .A(KEYINPUT0), .B(G125), .Z(n1315) );
INV_X1 U1019 ( .A(n1094), .ZN(n1301) );
NAND2_X1 U1020 ( .A1(G210), .A2(n1316), .ZN(n1094) );
INV_X1 U1021 ( .A(n1051), .ZN(n1047) );
NAND2_X1 U1022 ( .A1(G214), .A2(n1316), .ZN(n1051) );
NAND2_X1 U1023 ( .A1(n1317), .A2(n1282), .ZN(n1316) );
INV_X1 U1024 ( .A(G237), .ZN(n1317) );
AND2_X1 U1025 ( .A1(n1318), .A2(n1056), .ZN(n1049) );
NOR2_X1 U1026 ( .A1(n1319), .A2(n1083), .ZN(n1056) );
NOR2_X1 U1027 ( .A1(n1087), .A2(G472), .ZN(n1083) );
AND2_X1 U1028 ( .A1(G472), .A2(n1087), .ZN(n1319) );
NAND2_X1 U1029 ( .A1(n1320), .A2(n1282), .ZN(n1087) );
XOR2_X1 U1030 ( .A(n1156), .B(n1158), .Z(n1320) );
AND2_X1 U1031 ( .A1(n1321), .A2(n1322), .ZN(n1158) );
NAND2_X1 U1032 ( .A1(n1323), .A2(n1309), .ZN(n1322) );
INV_X1 U1033 ( .A(G101), .ZN(n1309) );
NAND2_X1 U1034 ( .A1(n1268), .A2(G210), .ZN(n1323) );
NAND3_X1 U1035 ( .A1(n1268), .A2(G210), .A3(G101), .ZN(n1321) );
NOR2_X1 U1036 ( .A1(G953), .A2(G237), .ZN(n1268) );
XOR2_X1 U1037 ( .A(n1324), .B(n1325), .Z(n1156) );
XOR2_X1 U1038 ( .A(n1311), .B(n1288), .Z(n1325) );
XNOR2_X1 U1039 ( .A(n1108), .B(n1326), .ZN(n1288) );
NOR2_X1 U1040 ( .A1(G137), .A2(KEYINPUT25), .ZN(n1326) );
XNOR2_X1 U1041 ( .A(G131), .B(G134), .ZN(n1108) );
XNOR2_X1 U1042 ( .A(n1244), .B(n1327), .ZN(n1311) );
XOR2_X1 U1043 ( .A(G119), .B(G116), .Z(n1327) );
INV_X1 U1044 ( .A(G113), .ZN(n1244) );
XOR2_X1 U1045 ( .A(n1215), .B(KEYINPUT18), .Z(n1324) );
NAND2_X1 U1046 ( .A1(n1293), .A2(n1328), .ZN(n1215) );
NAND2_X1 U1047 ( .A1(n1329), .A2(n1296), .ZN(n1328) );
XNOR2_X1 U1048 ( .A(KEYINPUT24), .B(n1297), .ZN(n1329) );
NAND2_X1 U1049 ( .A1(G146), .A2(n1297), .ZN(n1293) );
XNOR2_X1 U1050 ( .A(G128), .B(n1330), .ZN(n1297) );
XNOR2_X1 U1051 ( .A(KEYINPUT59), .B(n1219), .ZN(n1330) );
INV_X1 U1052 ( .A(G143), .ZN(n1219) );
XNOR2_X1 U1053 ( .A(KEYINPUT35), .B(n1052), .ZN(n1318) );
XNOR2_X1 U1054 ( .A(n1331), .B(n1135), .ZN(n1052) );
AND2_X1 U1055 ( .A1(G217), .A2(n1298), .ZN(n1135) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1282), .ZN(n1298) );
NAND2_X1 U1057 ( .A1(n1133), .A2(n1282), .ZN(n1331) );
INV_X1 U1058 ( .A(G902), .ZN(n1282) );
XNOR2_X1 U1059 ( .A(n1332), .B(n1333), .ZN(n1133) );
XOR2_X1 U1060 ( .A(KEYINPUT40), .B(KEYINPUT16), .Z(n1333) );
XOR2_X1 U1061 ( .A(n1334), .B(n1335), .Z(n1332) );
XOR2_X1 U1062 ( .A(n1336), .B(n1337), .Z(n1335) );
XNOR2_X1 U1063 ( .A(n1272), .B(G125), .ZN(n1337) );
INV_X1 U1064 ( .A(G128), .ZN(n1272) );
XOR2_X1 U1065 ( .A(KEYINPUT14), .B(G137), .Z(n1336) );
XOR2_X1 U1066 ( .A(n1338), .B(n1339), .Z(n1334) );
XOR2_X1 U1067 ( .A(n1267), .B(n1287), .Z(n1339) );
XNOR2_X1 U1068 ( .A(G110), .B(n1226), .ZN(n1287) );
INV_X1 U1069 ( .A(G140), .ZN(n1226) );
XNOR2_X1 U1070 ( .A(n1296), .B(KEYINPUT45), .ZN(n1267) );
INV_X1 U1071 ( .A(G146), .ZN(n1296) );
XOR2_X1 U1072 ( .A(n1340), .B(G119), .Z(n1338) );
NAND2_X1 U1073 ( .A1(n1341), .A2(n1279), .ZN(n1340) );
AND2_X1 U1074 ( .A1(G234), .A2(n1035), .ZN(n1279) );
INV_X1 U1075 ( .A(G953), .ZN(n1035) );
XNOR2_X1 U1076 ( .A(G221), .B(KEYINPUT58), .ZN(n1341) );
endmodule


