//Key = 1010011010100000011101000010001010011100111011011110101110010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;

XOR2_X1 U715 ( .A(n981), .B(n982), .Z(G9) );
NOR2_X1 U716 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR4_X1 U717 ( .A1(G953), .A2(n985), .A3(n986), .A4(n987), .ZN(n984) );
NOR2_X1 U718 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR2_X1 U719 ( .A1(n990), .A2(n991), .ZN(n988) );
NOR2_X1 U720 ( .A1(n992), .A2(n993), .ZN(n991) );
NOR2_X1 U721 ( .A1(n994), .A2(n995), .ZN(n992) );
NOR2_X1 U722 ( .A1(n996), .A2(n997), .ZN(n995) );
NOR3_X1 U723 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n996) );
NOR3_X1 U724 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n1000) );
NOR2_X1 U725 ( .A1(n1004), .A2(n1005), .ZN(n998) );
NOR2_X1 U726 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U727 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR3_X1 U728 ( .A1(n1002), .A2(n1010), .A3(n1005), .ZN(n994) );
XOR2_X1 U729 ( .A(n1011), .B(n1012), .Z(n1010) );
NOR4_X1 U730 ( .A1(n1013), .A2(n997), .A3(n1005), .A4(n1002), .ZN(n990) );
INV_X1 U731 ( .A(n1014), .ZN(n1002) );
NOR2_X1 U732 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR3_X1 U733 ( .A1(n985), .A2(G953), .A3(G952), .ZN(n983) );
AND4_X1 U734 ( .A1(n1017), .A2(n1009), .A3(n1011), .A4(n1018), .ZN(n985) );
NOR4_X1 U735 ( .A1(n1019), .A2(n1020), .A3(n1005), .A4(n1012), .ZN(n1018) );
NOR2_X1 U736 ( .A1(KEYINPUT63), .A2(n1016), .ZN(n1020) );
AND2_X1 U737 ( .A1(n993), .A2(KEYINPUT63), .ZN(n1019) );
XNOR2_X1 U738 ( .A(n1021), .B(n1022), .ZN(n1017) );
NOR2_X1 U739 ( .A1(KEYINPUT24), .A2(n1023), .ZN(n1021) );
XOR2_X1 U740 ( .A(n1024), .B(KEYINPUT14), .Z(n1023) );
XOR2_X1 U741 ( .A(n1025), .B(n1026), .Z(G72) );
NAND2_X1 U742 ( .A1(G953), .A2(n1027), .ZN(n1026) );
NAND2_X1 U743 ( .A1(G900), .A2(G227), .ZN(n1027) );
NAND4_X1 U744 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1025) );
NAND3_X1 U745 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
INV_X1 U746 ( .A(KEYINPUT15), .ZN(n1033) );
OR2_X1 U747 ( .A1(n1034), .A2(n1032), .ZN(n1030) );
NOR2_X1 U748 ( .A1(n1035), .A2(n1036), .ZN(n1032) );
INV_X1 U749 ( .A(KEYINPUT48), .ZN(n1035) );
XNOR2_X1 U750 ( .A(n1037), .B(n1038), .ZN(n1034) );
XNOR2_X1 U751 ( .A(n1039), .B(KEYINPUT53), .ZN(n1038) );
NAND2_X1 U752 ( .A1(n1040), .A2(KEYINPUT62), .ZN(n1039) );
XOR2_X1 U753 ( .A(n1041), .B(n1042), .Z(n1040) );
NAND2_X1 U754 ( .A1(G953), .A2(n1043), .ZN(n1029) );
NAND2_X1 U755 ( .A1(KEYINPUT15), .A2(n1036), .ZN(n1028) );
NAND2_X1 U756 ( .A1(n1044), .A2(n1045), .ZN(n1036) );
XOR2_X1 U757 ( .A(n1046), .B(n1047), .Z(G69) );
NOR2_X1 U758 ( .A1(n1048), .A2(n1044), .ZN(n1047) );
NOR2_X1 U759 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U760 ( .A1(KEYINPUT60), .A2(n1051), .ZN(n1046) );
XOR2_X1 U761 ( .A(n1052), .B(n1053), .Z(n1051) );
NOR2_X1 U762 ( .A1(n1054), .A2(G953), .ZN(n1053) );
NOR3_X1 U763 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
INV_X1 U764 ( .A(n982), .ZN(n1056) );
NAND2_X1 U765 ( .A1(n1058), .A2(n1059), .ZN(n1052) );
NAND2_X1 U766 ( .A1(G953), .A2(n1050), .ZN(n1059) );
XOR2_X1 U767 ( .A(n1060), .B(n1061), .Z(n1058) );
XOR2_X1 U768 ( .A(n1062), .B(n1063), .Z(n1061) );
XOR2_X1 U769 ( .A(n1064), .B(KEYINPUT11), .Z(n1060) );
NOR3_X1 U770 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(G66) );
NOR3_X1 U771 ( .A1(n1068), .A2(G953), .A3(G952), .ZN(n1067) );
AND2_X1 U772 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
INV_X1 U773 ( .A(KEYINPUT22), .ZN(n1068) );
XOR2_X1 U774 ( .A(n1070), .B(n1071), .Z(n1065) );
NAND3_X1 U775 ( .A1(G902), .A2(n1072), .A3(n1073), .ZN(n1070) );
XNOR2_X1 U776 ( .A(KEYINPUT36), .B(n987), .ZN(n1072) );
NOR2_X1 U777 ( .A1(n1069), .A2(n1074), .ZN(G63) );
XNOR2_X1 U778 ( .A(n1075), .B(n1076), .ZN(n1074) );
NOR2_X1 U779 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
INV_X1 U780 ( .A(G478), .ZN(n1077) );
NOR2_X1 U781 ( .A1(n1069), .A2(n1079), .ZN(G60) );
XOR2_X1 U782 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U783 ( .A1(n1082), .A2(n1078), .ZN(n1080) );
INV_X1 U784 ( .A(G475), .ZN(n1082) );
XOR2_X1 U785 ( .A(n1083), .B(n1084), .Z(G6) );
NOR2_X1 U786 ( .A1(n1069), .A2(n1085), .ZN(G57) );
XOR2_X1 U787 ( .A(n1086), .B(n1087), .Z(n1085) );
XOR2_X1 U788 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U789 ( .A1(n1090), .A2(n1078), .ZN(n1088) );
INV_X1 U790 ( .A(G472), .ZN(n1090) );
XOR2_X1 U791 ( .A(n1091), .B(n1092), .Z(n1086) );
NOR2_X1 U792 ( .A1(KEYINPUT28), .A2(n1093), .ZN(n1092) );
XNOR2_X1 U793 ( .A(KEYINPUT43), .B(KEYINPUT16), .ZN(n1091) );
NOR2_X1 U794 ( .A1(n1069), .A2(n1094), .ZN(G54) );
XOR2_X1 U795 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR2_X1 U796 ( .A1(n1097), .A2(n1078), .ZN(n1096) );
NOR2_X1 U797 ( .A1(n1098), .A2(n1099), .ZN(n1095) );
XOR2_X1 U798 ( .A(n1100), .B(KEYINPUT32), .Z(n1099) );
NAND2_X1 U799 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XNOR2_X1 U800 ( .A(n1103), .B(KEYINPUT5), .ZN(n1102) );
NOR2_X1 U801 ( .A1(n1103), .A2(n1101), .ZN(n1098) );
XOR2_X1 U802 ( .A(n1104), .B(KEYINPUT27), .Z(n1101) );
AND3_X1 U803 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1103) );
NAND2_X1 U804 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U805 ( .A1(KEYINPUT2), .A2(n1110), .ZN(n1109) );
XOR2_X1 U806 ( .A(n1111), .B(n1112), .Z(n1108) );
NAND4_X1 U807 ( .A1(n1113), .A2(KEYINPUT2), .A3(KEYINPUT10), .A4(n1110), .ZN(n1106) );
XNOR2_X1 U808 ( .A(n1111), .B(n1112), .ZN(n1113) );
OR2_X1 U809 ( .A1(n1110), .A2(KEYINPUT10), .ZN(n1105) );
NOR2_X1 U810 ( .A1(n1069), .A2(n1114), .ZN(G51) );
XOR2_X1 U811 ( .A(n1115), .B(n1116), .Z(n1114) );
XNOR2_X1 U812 ( .A(n1117), .B(n1118), .ZN(n1116) );
NOR2_X1 U813 ( .A1(KEYINPUT4), .A2(n1119), .ZN(n1118) );
NAND2_X1 U814 ( .A1(KEYINPUT59), .A2(n1120), .ZN(n1117) );
XOR2_X1 U815 ( .A(n1121), .B(n1122), .Z(n1115) );
NOR2_X1 U816 ( .A1(n1123), .A2(n1078), .ZN(n1122) );
NAND2_X1 U817 ( .A1(G902), .A2(n987), .ZN(n1078) );
OR4_X1 U818 ( .A1(n1045), .A2(n1055), .A3(n1124), .A4(n1125), .ZN(n987) );
XNOR2_X1 U819 ( .A(KEYINPUT41), .B(n1057), .ZN(n1125) );
AND3_X1 U820 ( .A1(n1014), .A2(n1126), .A3(n1127), .ZN(n1057) );
XOR2_X1 U821 ( .A(KEYINPUT57), .B(n1128), .Z(n1126) );
XOR2_X1 U822 ( .A(KEYINPUT54), .B(n982), .Z(n1124) );
NAND3_X1 U823 ( .A1(n1015), .A2(n1129), .A3(n1130), .ZN(n982) );
NAND4_X1 U824 ( .A1(n1131), .A2(n1132), .A3(n1084), .A4(n1133), .ZN(n1055) );
NOR3_X1 U825 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
INV_X1 U826 ( .A(n1137), .ZN(n1134) );
NAND3_X1 U827 ( .A1(n1130), .A2(n1129), .A3(n1016), .ZN(n1084) );
INV_X1 U828 ( .A(n997), .ZN(n1129) );
NAND4_X1 U829 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1045) );
NOR4_X1 U830 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
NOR2_X1 U831 ( .A1(n1146), .A2(n1147), .ZN(n1140) );
NOR2_X1 U832 ( .A1(n1005), .A2(n1148), .ZN(n1147) );
XNOR2_X1 U833 ( .A(KEYINPUT52), .B(n1149), .ZN(n1148) );
NOR2_X1 U834 ( .A1(n1044), .A2(G952), .ZN(n1069) );
XOR2_X1 U835 ( .A(n1142), .B(n1150), .Z(G48) );
NOR2_X1 U836 ( .A1(KEYINPUT58), .A2(n1151), .ZN(n1150) );
AND3_X1 U837 ( .A1(n1152), .A2(n1128), .A3(n1016), .ZN(n1142) );
XOR2_X1 U838 ( .A(G143), .B(n1146), .Z(G45) );
AND4_X1 U839 ( .A1(n1153), .A2(n1154), .A3(n1128), .A4(n1155), .ZN(n1146) );
XNOR2_X1 U840 ( .A(G140), .B(n1138), .ZN(G42) );
NAND3_X1 U841 ( .A1(n1156), .A2(n1007), .A3(n1157), .ZN(n1138) );
XOR2_X1 U842 ( .A(n1139), .B(n1158), .Z(G39) );
NAND2_X1 U843 ( .A1(KEYINPUT47), .A2(G137), .ZN(n1158) );
NAND3_X1 U844 ( .A1(n1152), .A2(n1156), .A3(n1159), .ZN(n1139) );
XOR2_X1 U845 ( .A(G134), .B(n1160), .Z(G36) );
NOR3_X1 U846 ( .A1(n1149), .A2(KEYINPUT39), .A3(n1005), .ZN(n1160) );
NAND2_X1 U847 ( .A1(n1154), .A2(n1015), .ZN(n1149) );
XOR2_X1 U848 ( .A(G131), .B(n1145), .Z(G33) );
AND3_X1 U849 ( .A1(n1016), .A2(n1156), .A3(n1154), .ZN(n1145) );
AND4_X1 U850 ( .A1(n1011), .A2(n1007), .A3(n1012), .A4(n1161), .ZN(n1154) );
INV_X1 U851 ( .A(n1005), .ZN(n1156) );
NAND2_X1 U852 ( .A1(n1162), .A2(n1001), .ZN(n1005) );
XOR2_X1 U853 ( .A(G128), .B(n1144), .Z(G30) );
AND3_X1 U854 ( .A1(n1015), .A2(n1128), .A3(n1152), .ZN(n1144) );
AND4_X1 U855 ( .A1(n1007), .A2(n1163), .A3(n1012), .A4(n1161), .ZN(n1152) );
NAND3_X1 U856 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(G3) );
NAND2_X1 U857 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
OR3_X1 U858 ( .A1(n1168), .A2(n1167), .A3(n1131), .ZN(n1165) );
INV_X1 U859 ( .A(KEYINPUT49), .ZN(n1168) );
NAND2_X1 U860 ( .A1(n1169), .A2(n1131), .ZN(n1164) );
NAND4_X1 U861 ( .A1(n1159), .A2(n1130), .A3(n1011), .A4(n1012), .ZN(n1131) );
INV_X1 U862 ( .A(n1170), .ZN(n1012) );
NAND2_X1 U863 ( .A1(n1171), .A2(KEYINPUT49), .ZN(n1169) );
XOR2_X1 U864 ( .A(n1167), .B(KEYINPUT30), .Z(n1171) );
XOR2_X1 U865 ( .A(n1172), .B(KEYINPUT8), .Z(n1167) );
XOR2_X1 U866 ( .A(G125), .B(n1143), .Z(G27) );
AND2_X1 U867 ( .A1(n999), .A2(n1157), .ZN(n1143) );
AND4_X1 U868 ( .A1(n1170), .A2(n1016), .A3(n1163), .A4(n1161), .ZN(n1157) );
NAND2_X1 U869 ( .A1(n989), .A2(n1173), .ZN(n1161) );
NAND4_X1 U870 ( .A1(G953), .A2(G902), .A3(n1174), .A4(n1043), .ZN(n1173) );
INV_X1 U871 ( .A(G900), .ZN(n1043) );
XOR2_X1 U872 ( .A(n1175), .B(G122), .Z(G24) );
NAND2_X1 U873 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND3_X1 U874 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1177) );
INV_X1 U875 ( .A(KEYINPUT0), .ZN(n1180) );
NAND2_X1 U876 ( .A1(n1136), .A2(KEYINPUT0), .ZN(n1176) );
AND2_X1 U877 ( .A1(n1179), .A2(n1181), .ZN(n1136) );
NOR4_X1 U878 ( .A1(n1182), .A2(n1183), .A3(n997), .A4(n1184), .ZN(n1179) );
NAND2_X1 U879 ( .A1(n1170), .A2(n1185), .ZN(n997) );
XOR2_X1 U880 ( .A(KEYINPUT61), .B(n1163), .Z(n1185) );
XOR2_X1 U881 ( .A(G119), .B(n1186), .Z(G21) );
AND2_X1 U882 ( .A1(n999), .A2(n1127), .ZN(n1186) );
NOR4_X1 U883 ( .A1(n993), .A2(n1011), .A3(n1170), .A4(n1178), .ZN(n1127) );
INV_X1 U884 ( .A(n1183), .ZN(n999) );
XOR2_X1 U885 ( .A(n1132), .B(n1187), .Z(G18) );
NOR2_X1 U886 ( .A1(G116), .A2(KEYINPUT29), .ZN(n1187) );
NAND2_X1 U887 ( .A1(n1188), .A2(n1015), .ZN(n1132) );
NOR2_X1 U888 ( .A1(n1153), .A2(n1184), .ZN(n1015) );
XOR2_X1 U889 ( .A(G113), .B(n1189), .Z(G15) );
NOR2_X1 U890 ( .A1(KEYINPUT3), .A2(n1137), .ZN(n1189) );
NAND2_X1 U891 ( .A1(n1188), .A2(n1016), .ZN(n1137) );
NOR2_X1 U892 ( .A1(n1155), .A2(n1182), .ZN(n1016) );
INV_X1 U893 ( .A(n1184), .ZN(n1155) );
NOR4_X1 U894 ( .A1(n1163), .A2(n1183), .A3(n1170), .A4(n1178), .ZN(n1188) );
INV_X1 U895 ( .A(n1181), .ZN(n1178) );
NAND2_X1 U896 ( .A1(n1014), .A2(n1128), .ZN(n1183) );
NOR2_X1 U897 ( .A1(n1190), .A2(n1008), .ZN(n1014) );
XOR2_X1 U898 ( .A(KEYINPUT56), .B(n1009), .Z(n1190) );
NAND2_X1 U899 ( .A1(n1191), .A2(n1192), .ZN(G12) );
OR2_X1 U900 ( .A1(n1193), .A2(G110), .ZN(n1192) );
NAND2_X1 U901 ( .A1(G110), .A2(n1194), .ZN(n1191) );
NAND2_X1 U902 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND2_X1 U903 ( .A1(KEYINPUT9), .A2(n1135), .ZN(n1196) );
NAND2_X1 U904 ( .A1(n1193), .A2(n1197), .ZN(n1195) );
INV_X1 U905 ( .A(KEYINPUT9), .ZN(n1197) );
NAND2_X1 U906 ( .A1(KEYINPUT42), .A2(n1135), .ZN(n1193) );
AND4_X1 U907 ( .A1(n1159), .A2(n1130), .A3(n1170), .A4(n1163), .ZN(n1135) );
INV_X1 U908 ( .A(n1011), .ZN(n1163) );
XOR2_X1 U909 ( .A(n1198), .B(n1073), .Z(n1011) );
AND2_X1 U910 ( .A1(G217), .A2(n1199), .ZN(n1073) );
NAND2_X1 U911 ( .A1(n1071), .A2(n1200), .ZN(n1198) );
XOR2_X1 U912 ( .A(n1201), .B(n1202), .Z(n1071) );
XNOR2_X1 U913 ( .A(n1203), .B(n1204), .ZN(n1202) );
NAND2_X1 U914 ( .A1(n1205), .A2(KEYINPUT55), .ZN(n1203) );
XOR2_X1 U915 ( .A(n1206), .B(G137), .Z(n1205) );
NAND2_X1 U916 ( .A1(n1207), .A2(G221), .ZN(n1206) );
XOR2_X1 U917 ( .A(n1208), .B(n1209), .Z(n1201) );
NOR2_X1 U918 ( .A1(KEYINPUT38), .A2(n1210), .ZN(n1209) );
NOR2_X1 U919 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U920 ( .A(KEYINPUT34), .B(n1213), .Z(n1212) );
NOR2_X1 U921 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U922 ( .A(KEYINPUT7), .B(n1037), .Z(n1215) );
NOR2_X1 U923 ( .A1(n1216), .A2(n1217), .ZN(n1211) );
INV_X1 U924 ( .A(n1214), .ZN(n1217) );
XOR2_X1 U925 ( .A(n1218), .B(KEYINPUT7), .Z(n1216) );
INV_X1 U926 ( .A(n1037), .ZN(n1218) );
XNOR2_X1 U927 ( .A(G128), .B(G119), .ZN(n1208) );
XOR2_X1 U928 ( .A(n1219), .B(G472), .Z(n1170) );
NAND2_X1 U929 ( .A1(n1220), .A2(n1200), .ZN(n1219) );
XNOR2_X1 U930 ( .A(n1093), .B(n1089), .ZN(n1220) );
XNOR2_X1 U931 ( .A(n1221), .B(n1222), .ZN(n1089) );
XOR2_X1 U932 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U933 ( .A(KEYINPUT31), .B(G119), .Z(n1224) );
NOR2_X1 U934 ( .A1(KEYINPUT51), .A2(n1225), .ZN(n1223) );
XOR2_X1 U935 ( .A(n1226), .B(n1227), .Z(n1221) );
NAND2_X1 U936 ( .A1(n1228), .A2(G210), .ZN(n1093) );
AND3_X1 U937 ( .A1(n1007), .A2(n1181), .A3(n1128), .ZN(n1130) );
AND2_X1 U938 ( .A1(n1003), .A2(n1001), .ZN(n1128) );
NAND2_X1 U939 ( .A1(G214), .A2(n1229), .ZN(n1001) );
INV_X1 U940 ( .A(n1162), .ZN(n1003) );
XNOR2_X1 U941 ( .A(n1230), .B(n1123), .ZN(n1162) );
NAND2_X1 U942 ( .A1(G210), .A2(n1229), .ZN(n1123) );
NAND2_X1 U943 ( .A1(n1231), .A2(n1200), .ZN(n1229) );
INV_X1 U944 ( .A(G237), .ZN(n1231) );
NAND2_X1 U945 ( .A1(n1232), .A2(n1200), .ZN(n1230) );
XOR2_X1 U946 ( .A(n1233), .B(n1120), .Z(n1232) );
XOR2_X1 U947 ( .A(n1064), .B(n1234), .Z(n1120) );
NOR2_X1 U948 ( .A1(KEYINPUT46), .A2(n1235), .ZN(n1234) );
XOR2_X1 U949 ( .A(n1236), .B(n1063), .Z(n1235) );
XNOR2_X1 U950 ( .A(n1237), .B(n1227), .ZN(n1063) );
XOR2_X1 U951 ( .A(G113), .B(KEYINPUT17), .Z(n1227) );
XOR2_X1 U952 ( .A(n1225), .B(G119), .Z(n1237) );
INV_X1 U953 ( .A(G116), .ZN(n1225) );
NAND2_X1 U954 ( .A1(KEYINPUT35), .A2(n1062), .ZN(n1236) );
XOR2_X1 U955 ( .A(n1238), .B(G101), .Z(n1062) );
NAND3_X1 U956 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1238) );
OR2_X1 U957 ( .A1(n981), .A2(KEYINPUT18), .ZN(n1241) );
NAND3_X1 U958 ( .A1(KEYINPUT18), .A2(n981), .A3(G104), .ZN(n1240) );
INV_X1 U959 ( .A(G107), .ZN(n981) );
NAND2_X1 U960 ( .A1(n1242), .A2(n1083), .ZN(n1239) );
INV_X1 U961 ( .A(G104), .ZN(n1083) );
NAND2_X1 U962 ( .A1(KEYINPUT18), .A2(n1243), .ZN(n1242) );
XOR2_X1 U963 ( .A(KEYINPUT21), .B(G107), .Z(n1243) );
NAND2_X1 U964 ( .A1(n1244), .A2(n1245), .ZN(n1064) );
NAND2_X1 U965 ( .A1(G122), .A2(n1204), .ZN(n1245) );
XOR2_X1 U966 ( .A(n1246), .B(KEYINPUT20), .Z(n1244) );
OR2_X1 U967 ( .A1(n1204), .A2(G122), .ZN(n1246) );
NAND2_X1 U968 ( .A1(KEYINPUT19), .A2(n1247), .ZN(n1233) );
XOR2_X1 U969 ( .A(n1119), .B(n1248), .Z(n1247) );
XNOR2_X1 U970 ( .A(n1121), .B(KEYINPUT13), .ZN(n1248) );
NOR2_X1 U971 ( .A1(n1049), .A2(G953), .ZN(n1121) );
INV_X1 U972 ( .A(G224), .ZN(n1049) );
XOR2_X1 U973 ( .A(n1249), .B(n1042), .Z(n1119) );
XOR2_X1 U974 ( .A(n1250), .B(KEYINPUT44), .Z(n1249) );
NAND2_X1 U975 ( .A1(n989), .A2(n1251), .ZN(n1181) );
NAND4_X1 U976 ( .A1(G953), .A2(G902), .A3(n1174), .A4(n1050), .ZN(n1251) );
INV_X1 U977 ( .A(G898), .ZN(n1050) );
NAND3_X1 U978 ( .A1(n1174), .A2(n1044), .A3(G952), .ZN(n989) );
NAND2_X1 U979 ( .A1(G237), .A2(G234), .ZN(n1174) );
AND2_X1 U980 ( .A1(n1008), .A2(n1252), .ZN(n1007) );
XNOR2_X1 U981 ( .A(KEYINPUT56), .B(n1009), .ZN(n1252) );
NAND2_X1 U982 ( .A1(G221), .A2(n1199), .ZN(n1009) );
NAND2_X1 U983 ( .A1(G234), .A2(n1200), .ZN(n1199) );
XOR2_X1 U984 ( .A(n1022), .B(n1253), .Z(n1008) );
INV_X1 U985 ( .A(n1024), .ZN(n1253) );
XOR2_X1 U986 ( .A(n1097), .B(KEYINPUT50), .Z(n1024) );
INV_X1 U987 ( .A(G469), .ZN(n1097) );
NAND2_X1 U988 ( .A1(n1254), .A2(n1200), .ZN(n1022) );
XOR2_X1 U989 ( .A(n1104), .B(n1255), .Z(n1254) );
XOR2_X1 U990 ( .A(n1226), .B(n1112), .Z(n1255) );
XNOR2_X1 U991 ( .A(n1256), .B(n1257), .ZN(n1112) );
XOR2_X1 U992 ( .A(G107), .B(G104), .Z(n1257) );
XNOR2_X1 U993 ( .A(KEYINPUT25), .B(KEYINPUT1), .ZN(n1256) );
XOR2_X1 U994 ( .A(n1110), .B(n1111), .Z(n1226) );
XNOR2_X1 U995 ( .A(n1172), .B(n1042), .ZN(n1111) );
XOR2_X1 U996 ( .A(n1258), .B(n1214), .Z(n1042) );
INV_X1 U997 ( .A(G101), .ZN(n1172) );
XOR2_X1 U998 ( .A(n1041), .B(KEYINPUT26), .Z(n1110) );
XOR2_X1 U999 ( .A(n1259), .B(n1260), .Z(n1041) );
XOR2_X1 U1000 ( .A(G137), .B(G134), .Z(n1260) );
INV_X1 U1001 ( .A(G131), .ZN(n1259) );
XNOR2_X1 U1002 ( .A(n1204), .B(n1261), .ZN(n1104) );
XOR2_X1 U1003 ( .A(G140), .B(n1262), .Z(n1261) );
AND2_X1 U1004 ( .A1(n1044), .A2(G227), .ZN(n1262) );
XOR2_X1 U1005 ( .A(G110), .B(KEYINPUT37), .Z(n1204) );
INV_X1 U1006 ( .A(n993), .ZN(n1159) );
NAND2_X1 U1007 ( .A1(n1184), .A2(n1182), .ZN(n993) );
INV_X1 U1008 ( .A(n1153), .ZN(n1182) );
XOR2_X1 U1009 ( .A(n1263), .B(n1264), .Z(n1153) );
XOR2_X1 U1010 ( .A(KEYINPUT6), .B(G475), .Z(n1264) );
OR2_X1 U1011 ( .A1(n1081), .A2(G902), .ZN(n1263) );
XNOR2_X1 U1012 ( .A(n1265), .B(n1266), .ZN(n1081) );
XOR2_X1 U1013 ( .A(n1267), .B(n1268), .Z(n1266) );
XOR2_X1 U1014 ( .A(G113), .B(G104), .Z(n1268) );
XOR2_X1 U1015 ( .A(G131), .B(G122), .Z(n1267) );
XOR2_X1 U1016 ( .A(n1269), .B(n1270), .Z(n1265) );
XOR2_X1 U1017 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U1018 ( .A1(G143), .A2(KEYINPUT33), .ZN(n1272) );
AND2_X1 U1019 ( .A1(G214), .A2(n1228), .ZN(n1271) );
NOR2_X1 U1020 ( .A1(G953), .A2(G237), .ZN(n1228) );
XOR2_X1 U1021 ( .A(n1273), .B(n1037), .Z(n1269) );
XOR2_X1 U1022 ( .A(G140), .B(n1274), .Z(n1037) );
INV_X1 U1023 ( .A(n1250), .ZN(n1274) );
XNOR2_X1 U1024 ( .A(G125), .B(KEYINPUT40), .ZN(n1250) );
NAND2_X1 U1025 ( .A1(KEYINPUT45), .A2(n1214), .ZN(n1273) );
XOR2_X1 U1026 ( .A(n1151), .B(KEYINPUT23), .Z(n1214) );
INV_X1 U1027 ( .A(G146), .ZN(n1151) );
XOR2_X1 U1028 ( .A(n1275), .B(G478), .Z(n1184) );
NAND2_X1 U1029 ( .A1(n1075), .A2(n1200), .ZN(n1275) );
INV_X1 U1030 ( .A(G902), .ZN(n1200) );
XNOR2_X1 U1031 ( .A(n1276), .B(n1277), .ZN(n1075) );
XOR2_X1 U1032 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U1033 ( .A(G122), .B(G116), .Z(n1279) );
XOR2_X1 U1034 ( .A(KEYINPUT12), .B(G134), .Z(n1278) );
XNOR2_X1 U1035 ( .A(n1280), .B(n1258), .ZN(n1276) );
XNOR2_X1 U1036 ( .A(G128), .B(G143), .ZN(n1258) );
XOR2_X1 U1037 ( .A(n1281), .B(G107), .Z(n1280) );
NAND2_X1 U1038 ( .A1(G217), .A2(n1207), .ZN(n1281) );
AND2_X1 U1039 ( .A1(G234), .A2(n1044), .ZN(n1207) );
INV_X1 U1040 ( .A(G953), .ZN(n1044) );
endmodule


