//Key = 1010101110110001100100001101100001010101111110101110111101111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;

XOR2_X1 U729 ( .A(G107), .B(n1010), .Z(G9) );
NOR2_X1 U730 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .ZN(n1012) );
NOR4_X1 U732 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1015) );
INV_X1 U733 ( .A(n1021), .ZN(n1019) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1017) );
NOR2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
INV_X1 U736 ( .A(n1026), .ZN(n1025) );
NOR2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1024) );
NOR2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1022) );
NOR2_X1 U740 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NAND4_X1 U742 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1013) );
NAND4_X1 U743 ( .A1(n1041), .A2(n1026), .A3(n1042), .A4(n1043), .ZN(n1037) );
NAND2_X1 U744 ( .A1(n1044), .A2(n1020), .ZN(n1043) );
NAND2_X1 U745 ( .A1(KEYINPUT17), .A2(n1045), .ZN(n1044) );
NAND4_X1 U746 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1042) );
INV_X1 U747 ( .A(n1020), .ZN(n1049) );
NAND2_X1 U748 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND2_X1 U749 ( .A1(n1021), .A2(n1052), .ZN(n1047) );
NAND2_X1 U750 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1055), .ZN(n1046) );
INV_X1 U752 ( .A(KEYINPUT17), .ZN(n1055) );
NOR3_X1 U753 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1011) );
INV_X1 U754 ( .A(n1039), .ZN(n1056) );
NAND4_X1 U755 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1039) );
NOR4_X1 U756 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1035), .ZN(n1060) );
XNOR2_X1 U757 ( .A(n1029), .B(KEYINPUT61), .ZN(n1062) );
XNOR2_X1 U758 ( .A(n1064), .B(KEYINPUT11), .ZN(n1061) );
NOR3_X1 U759 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1059) );
XNOR2_X1 U760 ( .A(KEYINPUT39), .B(n1068), .ZN(n1057) );
XOR2_X1 U761 ( .A(n1069), .B(n1070), .Z(G72) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1040), .ZN(n1070) );
NOR2_X1 U763 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U764 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
NAND2_X1 U765 ( .A1(n1076), .A2(n1040), .ZN(n1075) );
XNOR2_X1 U766 ( .A(n1077), .B(n1078), .ZN(n1076) );
NAND3_X1 U767 ( .A1(G900), .A2(n1078), .A3(G953), .ZN(n1074) );
XNOR2_X1 U768 ( .A(n1079), .B(n1080), .ZN(n1078) );
NOR2_X1 U769 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NOR2_X1 U770 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U771 ( .A(G125), .B(KEYINPUT36), .ZN(n1083) );
XOR2_X1 U772 ( .A(n1085), .B(n1086), .Z(G69) );
NOR2_X1 U773 ( .A1(KEYINPUT1), .A2(n1087), .ZN(n1086) );
XOR2_X1 U774 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1040), .ZN(n1089) );
NAND2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U777 ( .A(n1038), .B(KEYINPUT23), .Z(n1091) );
NAND3_X1 U778 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1088) );
OR2_X1 U779 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
NAND2_X1 U780 ( .A1(n1096), .A2(n1098), .ZN(n1093) );
XNOR2_X1 U781 ( .A(n1097), .B(KEYINPUT16), .ZN(n1098) );
XOR2_X1 U782 ( .A(n1099), .B(n1100), .Z(n1096) );
NAND2_X1 U783 ( .A1(G953), .A2(n1101), .ZN(n1085) );
NAND2_X1 U784 ( .A1(G898), .A2(n1102), .ZN(n1101) );
XOR2_X1 U785 ( .A(KEYINPUT3), .B(G224), .Z(n1102) );
NOR2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(G66) );
XNOR2_X1 U787 ( .A(n1105), .B(n1106), .ZN(n1104) );
NOR2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR2_X1 U789 ( .A1(n1103), .A2(n1109), .ZN(G63) );
XOR2_X1 U790 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U791 ( .A1(n1112), .A2(n1108), .ZN(n1111) );
NAND2_X1 U792 ( .A1(n1113), .A2(KEYINPUT0), .ZN(n1110) );
XOR2_X1 U793 ( .A(n1114), .B(KEYINPUT5), .Z(n1113) );
NOR2_X1 U794 ( .A1(n1103), .A2(n1115), .ZN(G60) );
XOR2_X1 U795 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U796 ( .A1(n1118), .A2(n1108), .ZN(n1116) );
XOR2_X1 U797 ( .A(G104), .B(n1119), .Z(G6) );
NOR2_X1 U798 ( .A1(n1103), .A2(n1120), .ZN(G57) );
XOR2_X1 U799 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U800 ( .A(n1123), .B(n1124), .ZN(n1121) );
NOR2_X1 U801 ( .A1(n1125), .A2(n1108), .ZN(n1124) );
NOR2_X1 U802 ( .A1(n1103), .A2(n1126), .ZN(G54) );
XOR2_X1 U803 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U804 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U805 ( .A1(n1131), .A2(n1108), .ZN(n1129) );
XOR2_X1 U806 ( .A(n1132), .B(n1133), .Z(n1127) );
XNOR2_X1 U807 ( .A(KEYINPUT20), .B(n1084), .ZN(n1133) );
NOR2_X1 U808 ( .A1(n1103), .A2(n1134), .ZN(G51) );
XOR2_X1 U809 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U810 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR3_X1 U811 ( .A1(n1108), .A2(KEYINPUT29), .A3(n1139), .ZN(n1138) );
NAND2_X1 U812 ( .A1(n1140), .A2(n1141), .ZN(n1108) );
NAND3_X1 U813 ( .A1(n1077), .A2(n1038), .A3(n1092), .ZN(n1141) );
INV_X1 U814 ( .A(n1014), .ZN(n1092) );
NAND4_X1 U815 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1014) );
NOR4_X1 U816 ( .A1(n1146), .A2(n1147), .A3(n1119), .A4(n1010), .ZN(n1145) );
AND3_X1 U817 ( .A1(n1148), .A2(n1149), .A3(n1021), .ZN(n1010) );
AND3_X1 U818 ( .A1(n1021), .A2(n1148), .A3(n1150), .ZN(n1119) );
NAND2_X1 U819 ( .A1(n1028), .A2(n1151), .ZN(n1144) );
XNOR2_X1 U820 ( .A(KEYINPUT31), .B(n1152), .ZN(n1151) );
INV_X1 U821 ( .A(n1016), .ZN(n1077) );
NAND4_X1 U822 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1016) );
NOR4_X1 U823 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
NAND2_X1 U824 ( .A1(KEYINPUT10), .A2(n1161), .ZN(n1155) );
INV_X1 U825 ( .A(n1162), .ZN(n1161) );
NAND2_X1 U826 ( .A1(n1041), .A2(n1163), .ZN(n1154) );
NAND2_X1 U827 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U828 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND2_X1 U829 ( .A1(n1028), .A2(n1168), .ZN(n1153) );
NAND2_X1 U830 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND3_X1 U831 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1170) );
NOR3_X1 U832 ( .A1(n1068), .A2(KEYINPUT10), .A3(n1167), .ZN(n1173) );
NAND4_X1 U833 ( .A1(n1050), .A2(n1150), .A3(n1026), .A4(n1174), .ZN(n1169) );
XNOR2_X1 U834 ( .A(KEYINPUT62), .B(n1175), .ZN(n1140) );
NAND2_X1 U835 ( .A1(KEYINPUT55), .A2(n1176), .ZN(n1137) );
XNOR2_X1 U836 ( .A(G125), .B(n1177), .ZN(n1176) );
XOR2_X1 U837 ( .A(n1178), .B(n1179), .Z(n1135) );
NOR2_X1 U838 ( .A1(n1040), .A2(G952), .ZN(n1103) );
XNOR2_X1 U839 ( .A(n1160), .B(n1180), .ZN(G48) );
XOR2_X1 U840 ( .A(KEYINPUT60), .B(G146), .Z(n1180) );
AND3_X1 U841 ( .A1(n1181), .A2(n1028), .A3(n1166), .ZN(n1160) );
XNOR2_X1 U842 ( .A(G143), .B(n1162), .ZN(G45) );
NAND3_X1 U843 ( .A1(n1171), .A2(n1172), .A3(n1182), .ZN(n1162) );
NOR3_X1 U844 ( .A1(n1183), .A2(n1068), .A3(n1184), .ZN(n1182) );
XOR2_X1 U845 ( .A(n1185), .B(n1159), .Z(G42) );
AND3_X1 U846 ( .A1(n1041), .A2(n1050), .A3(n1166), .ZN(n1159) );
INV_X1 U847 ( .A(n1186), .ZN(n1166) );
NAND2_X1 U848 ( .A1(KEYINPUT54), .A2(n1084), .ZN(n1185) );
NAND2_X1 U849 ( .A1(n1187), .A2(n1188), .ZN(G39) );
NAND2_X1 U850 ( .A1(n1158), .A2(n1189), .ZN(n1188) );
XOR2_X1 U851 ( .A(KEYINPUT41), .B(n1190), .Z(n1187) );
NOR2_X1 U852 ( .A1(n1158), .A2(n1189), .ZN(n1190) );
INV_X1 U853 ( .A(G137), .ZN(n1189) );
AND4_X1 U854 ( .A1(n1172), .A2(n1041), .A3(n1181), .A4(n1051), .ZN(n1158) );
XOR2_X1 U855 ( .A(G134), .B(n1191), .Z(G36) );
NOR3_X1 U856 ( .A1(n1192), .A2(KEYINPUT18), .A3(n1032), .ZN(n1191) );
INV_X1 U857 ( .A(n1041), .ZN(n1032) );
XNOR2_X1 U858 ( .A(KEYINPUT50), .B(n1164), .ZN(n1192) );
NAND3_X1 U859 ( .A1(n1167), .A2(n1149), .A3(n1172), .ZN(n1164) );
XOR2_X1 U860 ( .A(n1193), .B(n1194), .Z(G33) );
NOR2_X1 U861 ( .A1(KEYINPUT13), .A2(n1195), .ZN(n1194) );
NOR3_X1 U862 ( .A1(n1186), .A2(n1196), .A3(n1183), .ZN(n1193) );
XNOR2_X1 U863 ( .A(n1041), .B(KEYINPUT47), .ZN(n1196) );
NOR2_X1 U864 ( .A1(n1029), .A2(n1066), .ZN(n1041) );
NAND2_X1 U865 ( .A1(n1172), .A2(n1150), .ZN(n1186) );
AND2_X1 U866 ( .A1(n1034), .A2(n1174), .ZN(n1172) );
XOR2_X1 U867 ( .A(G128), .B(n1157), .Z(G30) );
AND3_X1 U868 ( .A1(n1197), .A2(n1181), .A3(n1198), .ZN(n1157) );
NOR3_X1 U869 ( .A1(n1184), .A2(n1199), .A3(n1053), .ZN(n1198) );
INV_X1 U870 ( .A(n1149), .ZN(n1053) );
XOR2_X1 U871 ( .A(G101), .B(n1147), .Z(G3) );
AND2_X1 U872 ( .A1(n1045), .A2(n1148), .ZN(n1147) );
NOR2_X1 U873 ( .A1(n1183), .A2(n1018), .ZN(n1045) );
INV_X1 U874 ( .A(n1167), .ZN(n1183) );
XNOR2_X1 U875 ( .A(G125), .B(n1200), .ZN(G27) );
NAND3_X1 U876 ( .A1(n1201), .A2(n1050), .A3(n1202), .ZN(n1200) );
NOR3_X1 U877 ( .A1(n1054), .A2(n1199), .A3(n1184), .ZN(n1202) );
INV_X1 U878 ( .A(n1174), .ZN(n1199) );
NAND2_X1 U879 ( .A1(n1020), .A2(n1203), .ZN(n1174) );
NAND4_X1 U880 ( .A1(G902), .A2(G953), .A3(n1204), .A4(n1073), .ZN(n1203) );
INV_X1 U881 ( .A(G900), .ZN(n1073) );
INV_X1 U882 ( .A(n1150), .ZN(n1054) );
XNOR2_X1 U883 ( .A(KEYINPUT4), .B(n1026), .ZN(n1201) );
NAND2_X1 U884 ( .A1(n1205), .A2(n1206), .ZN(G24) );
NAND2_X1 U885 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U886 ( .A1(G122), .A2(n1209), .ZN(n1205) );
NAND2_X1 U887 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
OR2_X1 U888 ( .A1(n1143), .A2(KEYINPUT28), .ZN(n1211) );
NAND2_X1 U889 ( .A1(KEYINPUT28), .A2(n1212), .ZN(n1210) );
INV_X1 U890 ( .A(n1207), .ZN(n1212) );
NOR2_X1 U891 ( .A1(KEYINPUT38), .A2(n1143), .ZN(n1207) );
NAND4_X1 U892 ( .A1(n1026), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1143) );
AND2_X1 U893 ( .A1(n1021), .A2(n1171), .ZN(n1215) );
XNOR2_X1 U894 ( .A(n1063), .B(KEYINPUT48), .ZN(n1171) );
NOR2_X1 U895 ( .A1(n1216), .A2(n1064), .ZN(n1021) );
NAND2_X1 U896 ( .A1(n1217), .A2(n1218), .ZN(G21) );
NAND2_X1 U897 ( .A1(n1146), .A2(n1219), .ZN(n1218) );
XOR2_X1 U898 ( .A(KEYINPUT15), .B(n1220), .Z(n1217) );
NOR2_X1 U899 ( .A1(n1146), .A2(n1219), .ZN(n1220) );
AND4_X1 U900 ( .A1(n1181), .A2(n1051), .A3(n1214), .A4(n1026), .ZN(n1146) );
AND2_X1 U901 ( .A1(n1064), .A2(n1216), .ZN(n1181) );
XNOR2_X1 U902 ( .A(G116), .B(n1038), .ZN(G18) );
NAND4_X1 U903 ( .A1(n1167), .A2(n1214), .A3(n1026), .A4(n1149), .ZN(n1038) );
NAND2_X1 U904 ( .A1(n1221), .A2(n1222), .ZN(n1149) );
OR2_X1 U905 ( .A1(n1018), .A2(KEYINPUT48), .ZN(n1222) );
INV_X1 U906 ( .A(n1051), .ZN(n1018) );
NAND3_X1 U907 ( .A1(n1063), .A2(n1068), .A3(KEYINPUT48), .ZN(n1221) );
XNOR2_X1 U908 ( .A(n1223), .B(n1224), .ZN(G15) );
NOR2_X1 U909 ( .A1(n1184), .A2(n1152), .ZN(n1224) );
NAND4_X1 U910 ( .A1(n1150), .A2(n1167), .A3(n1026), .A4(n1225), .ZN(n1152) );
NAND2_X1 U911 ( .A1(n1226), .A2(n1227), .ZN(n1026) );
NAND2_X1 U912 ( .A1(n1034), .A2(n1228), .ZN(n1227) );
INV_X1 U913 ( .A(KEYINPUT35), .ZN(n1228) );
NAND3_X1 U914 ( .A1(n1229), .A2(n1036), .A3(KEYINPUT35), .ZN(n1226) );
NOR2_X1 U915 ( .A1(n1216), .A2(n1230), .ZN(n1167) );
NOR2_X1 U916 ( .A1(n1063), .A2(n1068), .ZN(n1150) );
INV_X1 U917 ( .A(n1213), .ZN(n1068) );
INV_X1 U918 ( .A(n1028), .ZN(n1184) );
XNOR2_X1 U919 ( .A(G110), .B(n1142), .ZN(G12) );
NAND3_X1 U920 ( .A1(n1148), .A2(n1051), .A3(n1050), .ZN(n1142) );
AND2_X1 U921 ( .A1(n1230), .A2(n1216), .ZN(n1050) );
NAND2_X1 U922 ( .A1(n1231), .A2(n1058), .ZN(n1216) );
NAND2_X1 U923 ( .A1(n1232), .A2(n1233), .ZN(n1058) );
XNOR2_X1 U924 ( .A(n1067), .B(KEYINPUT26), .ZN(n1231) );
NOR2_X1 U925 ( .A1(n1233), .A2(n1232), .ZN(n1067) );
INV_X1 U926 ( .A(n1107), .ZN(n1232) );
NAND2_X1 U927 ( .A1(G217), .A2(n1234), .ZN(n1107) );
NAND2_X1 U928 ( .A1(n1105), .A2(n1175), .ZN(n1233) );
XNOR2_X1 U929 ( .A(n1235), .B(n1236), .ZN(n1105) );
XOR2_X1 U930 ( .A(n1237), .B(n1238), .Z(n1236) );
XNOR2_X1 U931 ( .A(G119), .B(G137), .ZN(n1238) );
NAND3_X1 U932 ( .A1(G234), .A2(n1040), .A3(G221), .ZN(n1237) );
XOR2_X1 U933 ( .A(n1239), .B(n1240), .Z(n1235) );
XOR2_X1 U934 ( .A(n1241), .B(n1242), .Z(n1239) );
NAND2_X1 U935 ( .A1(n1243), .A2(n1244), .ZN(n1241) );
NAND2_X1 U936 ( .A1(G140), .A2(G125), .ZN(n1244) );
INV_X1 U937 ( .A(n1064), .ZN(n1230) );
XOR2_X1 U938 ( .A(n1245), .B(n1125), .Z(n1064) );
INV_X1 U939 ( .A(G472), .ZN(n1125) );
NAND2_X1 U940 ( .A1(n1246), .A2(n1175), .ZN(n1245) );
XNOR2_X1 U941 ( .A(n1247), .B(n1122), .ZN(n1246) );
XNOR2_X1 U942 ( .A(n1248), .B(n1249), .ZN(n1122) );
XNOR2_X1 U943 ( .A(n1250), .B(n1251), .ZN(n1249) );
NAND2_X1 U944 ( .A1(G210), .A2(n1252), .ZN(n1250) );
XOR2_X1 U945 ( .A(n1177), .B(n1253), .Z(n1248) );
NAND2_X1 U946 ( .A1(KEYINPUT7), .A2(n1123), .ZN(n1247) );
AND2_X1 U947 ( .A1(n1254), .A2(n1255), .ZN(n1123) );
NAND2_X1 U948 ( .A1(n1256), .A2(G113), .ZN(n1255) );
XNOR2_X1 U949 ( .A(G116), .B(n1257), .ZN(n1256) );
XOR2_X1 U950 ( .A(n1258), .B(KEYINPUT21), .Z(n1254) );
NAND2_X1 U951 ( .A1(n1259), .A2(n1223), .ZN(n1258) );
XNOR2_X1 U952 ( .A(n1260), .B(n1257), .ZN(n1259) );
NOR2_X1 U953 ( .A1(G119), .A2(KEYINPUT45), .ZN(n1257) );
INV_X1 U954 ( .A(G116), .ZN(n1260) );
NOR2_X1 U955 ( .A1(n1063), .A2(n1213), .ZN(n1051) );
XOR2_X1 U956 ( .A(n1261), .B(n1118), .Z(n1213) );
INV_X1 U957 ( .A(G475), .ZN(n1118) );
OR2_X1 U958 ( .A1(n1117), .A2(G902), .ZN(n1261) );
XOR2_X1 U959 ( .A(n1262), .B(n1208), .Z(n1117) );
XOR2_X1 U960 ( .A(n1263), .B(n1264), .Z(n1262) );
XOR2_X1 U961 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U962 ( .A(n1223), .B(G104), .ZN(n1266) );
INV_X1 U963 ( .A(G113), .ZN(n1223) );
XNOR2_X1 U964 ( .A(KEYINPUT51), .B(n1267), .ZN(n1265) );
XOR2_X1 U965 ( .A(n1268), .B(n1269), .Z(n1263) );
XOR2_X1 U966 ( .A(n1270), .B(n1271), .Z(n1269) );
NAND2_X1 U967 ( .A1(G214), .A2(n1252), .ZN(n1271) );
NOR2_X1 U968 ( .A1(G953), .A2(G237), .ZN(n1252) );
NAND2_X1 U969 ( .A1(KEYINPUT19), .A2(n1272), .ZN(n1270) );
XOR2_X1 U970 ( .A(KEYINPUT42), .B(G146), .Z(n1272) );
XOR2_X1 U971 ( .A(n1273), .B(n1274), .Z(n1268) );
NAND2_X1 U972 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND3_X1 U973 ( .A1(n1243), .A2(n1084), .A3(KEYINPUT43), .ZN(n1276) );
INV_X1 U974 ( .A(G140), .ZN(n1084) );
INV_X1 U975 ( .A(n1081), .ZN(n1243) );
NAND2_X1 U976 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
INV_X1 U977 ( .A(G125), .ZN(n1278) );
NAND2_X1 U978 ( .A1(n1081), .A2(KEYINPUT43), .ZN(n1277) );
NOR2_X1 U979 ( .A1(G125), .A2(G140), .ZN(n1081) );
XOR2_X1 U980 ( .A(n1279), .B(n1112), .Z(n1063) );
INV_X1 U981 ( .A(G478), .ZN(n1112) );
NAND2_X1 U982 ( .A1(n1175), .A2(n1114), .ZN(n1279) );
NAND3_X1 U983 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1114) );
NAND4_X1 U984 ( .A1(G217), .A2(G234), .A3(n1283), .A4(n1040), .ZN(n1282) );
NAND2_X1 U985 ( .A1(KEYINPUT44), .A2(n1284), .ZN(n1283) );
NAND2_X1 U986 ( .A1(KEYINPUT57), .A2(n1285), .ZN(n1284) );
INV_X1 U987 ( .A(n1286), .ZN(n1285) );
OR2_X1 U988 ( .A1(n1286), .A2(KEYINPUT44), .ZN(n1281) );
NAND3_X1 U989 ( .A1(n1286), .A2(n1287), .A3(KEYINPUT44), .ZN(n1280) );
NAND4_X1 U990 ( .A1(KEYINPUT57), .A2(G217), .A3(G234), .A4(n1040), .ZN(n1287) );
XNOR2_X1 U991 ( .A(n1288), .B(n1289), .ZN(n1286) );
XNOR2_X1 U992 ( .A(G107), .B(n1290), .ZN(n1289) );
NAND2_X1 U993 ( .A1(KEYINPUT8), .A2(n1291), .ZN(n1290) );
XNOR2_X1 U994 ( .A(n1267), .B(G128), .ZN(n1291) );
INV_X1 U995 ( .A(G143), .ZN(n1267) );
XNOR2_X1 U996 ( .A(G116), .B(n1292), .ZN(n1288) );
XNOR2_X1 U997 ( .A(G134), .B(n1208), .ZN(n1292) );
INV_X1 U998 ( .A(G122), .ZN(n1208) );
AND2_X1 U999 ( .A1(n1214), .A2(n1197), .ZN(n1148) );
XNOR2_X1 U1000 ( .A(n1034), .B(KEYINPUT40), .ZN(n1197) );
NOR2_X1 U1001 ( .A1(n1229), .A2(n1065), .ZN(n1034) );
INV_X1 U1002 ( .A(n1036), .ZN(n1065) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1234), .ZN(n1036) );
NAND2_X1 U1004 ( .A1(G234), .A2(n1175), .ZN(n1234) );
INV_X1 U1005 ( .A(n1035), .ZN(n1229) );
XOR2_X1 U1006 ( .A(n1293), .B(n1131), .Z(n1035) );
INV_X1 U1007 ( .A(G469), .ZN(n1131) );
NAND2_X1 U1008 ( .A1(n1294), .A2(n1175), .ZN(n1293) );
XOR2_X1 U1009 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1010 ( .A(n1297), .B(n1130), .Z(n1296) );
XNOR2_X1 U1011 ( .A(n1298), .B(n1299), .ZN(n1130) );
XNOR2_X1 U1012 ( .A(n1300), .B(n1079), .ZN(n1299) );
XOR2_X1 U1013 ( .A(n1301), .B(n1253), .Z(n1079) );
XNOR2_X1 U1014 ( .A(n1302), .B(n1274), .ZN(n1253) );
XNOR2_X1 U1015 ( .A(n1195), .B(KEYINPUT49), .ZN(n1274) );
INV_X1 U1016 ( .A(G131), .ZN(n1195) );
XNOR2_X1 U1017 ( .A(G134), .B(G137), .ZN(n1302) );
XOR2_X1 U1018 ( .A(n1303), .B(KEYINPUT34), .Z(n1301) );
NAND2_X1 U1019 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U1020 ( .A1(G128), .A2(n1306), .ZN(n1305) );
XOR2_X1 U1021 ( .A(KEYINPUT37), .B(n1307), .Z(n1304) );
NOR2_X1 U1022 ( .A1(G128), .A2(n1306), .ZN(n1307) );
XNOR2_X1 U1023 ( .A(G143), .B(n1308), .ZN(n1306) );
NAND2_X1 U1024 ( .A1(KEYINPUT52), .A2(G146), .ZN(n1308) );
XOR2_X1 U1025 ( .A(n1309), .B(n1242), .Z(n1298) );
XNOR2_X1 U1026 ( .A(KEYINPUT59), .B(n1310), .ZN(n1309) );
NOR2_X1 U1027 ( .A1(KEYINPUT12), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1028 ( .A1(n1312), .A2(KEYINPUT46), .ZN(n1297) );
XNOR2_X1 U1029 ( .A(n1132), .B(KEYINPUT63), .ZN(n1312) );
NOR2_X1 U1030 ( .A1(n1072), .A2(G953), .ZN(n1132) );
INV_X1 U1031 ( .A(G227), .ZN(n1072) );
XOR2_X1 U1032 ( .A(n1313), .B(n1314), .Z(n1295) );
NOR2_X1 U1033 ( .A1(G140), .A2(KEYINPUT32), .ZN(n1314) );
XNOR2_X1 U1034 ( .A(KEYINPUT6), .B(KEYINPUT27), .ZN(n1313) );
AND2_X1 U1035 ( .A1(n1028), .A2(n1225), .ZN(n1214) );
NAND2_X1 U1036 ( .A1(n1020), .A2(n1315), .ZN(n1225) );
NAND3_X1 U1037 ( .A1(n1316), .A2(n1204), .A3(G902), .ZN(n1315) );
INV_X1 U1038 ( .A(n1095), .ZN(n1316) );
NAND2_X1 U1039 ( .A1(n1317), .A2(G953), .ZN(n1095) );
XNOR2_X1 U1040 ( .A(G898), .B(KEYINPUT56), .ZN(n1317) );
NAND3_X1 U1041 ( .A1(n1204), .A2(n1040), .A3(G952), .ZN(n1020) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1204) );
NOR2_X1 U1043 ( .A1(n1318), .A2(n1066), .ZN(n1028) );
INV_X1 U1044 ( .A(n1030), .ZN(n1066) );
NAND2_X1 U1045 ( .A1(n1319), .A2(G214), .ZN(n1030) );
XOR2_X1 U1046 ( .A(n1320), .B(KEYINPUT30), .Z(n1319) );
INV_X1 U1047 ( .A(n1029), .ZN(n1318) );
XOR2_X1 U1048 ( .A(n1321), .B(n1139), .Z(n1029) );
NAND2_X1 U1049 ( .A1(G210), .A2(n1320), .ZN(n1139) );
OR2_X1 U1050 ( .A1(G902), .A2(G237), .ZN(n1320) );
NAND3_X1 U1051 ( .A1(n1322), .A2(n1175), .A3(n1323), .ZN(n1321) );
XOR2_X1 U1052 ( .A(n1324), .B(KEYINPUT14), .Z(n1323) );
NAND2_X1 U1053 ( .A1(n1325), .A2(n1178), .ZN(n1324) );
INV_X1 U1054 ( .A(G902), .ZN(n1175) );
OR2_X1 U1055 ( .A1(n1178), .A2(n1325), .ZN(n1322) );
XNOR2_X1 U1056 ( .A(n1326), .B(n1179), .ZN(n1325) );
NAND2_X1 U1057 ( .A1(G224), .A2(n1040), .ZN(n1179) );
INV_X1 U1058 ( .A(G953), .ZN(n1040) );
NAND2_X1 U1059 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
NAND2_X1 U1060 ( .A1(n1177), .A2(G125), .ZN(n1328) );
XOR2_X1 U1061 ( .A(KEYINPUT24), .B(n1329), .Z(n1327) );
NOR2_X1 U1062 ( .A1(G125), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1063 ( .A(n1177), .B(n1331), .Z(n1330) );
XOR2_X1 U1064 ( .A(KEYINPUT25), .B(KEYINPUT2), .Z(n1331) );
XNOR2_X1 U1065 ( .A(G143), .B(n1240), .ZN(n1177) );
XOR2_X1 U1066 ( .A(G128), .B(G146), .Z(n1240) );
NAND2_X1 U1067 ( .A1(n1332), .A2(n1333), .ZN(n1178) );
NAND2_X1 U1068 ( .A1(n1334), .A2(n1097), .ZN(n1333) );
XOR2_X1 U1069 ( .A(KEYINPUT58), .B(n1335), .Z(n1332) );
NOR2_X1 U1070 ( .A1(n1334), .A2(n1097), .ZN(n1335) );
XOR2_X1 U1071 ( .A(G122), .B(n1242), .Z(n1097) );
XOR2_X1 U1072 ( .A(G110), .B(KEYINPUT22), .Z(n1242) );
XNOR2_X1 U1073 ( .A(n1100), .B(n1336), .ZN(n1334) );
NOR2_X1 U1074 ( .A1(KEYINPUT9), .A2(n1099), .ZN(n1336) );
XOR2_X1 U1075 ( .A(G113), .B(n1337), .Z(n1099) );
XNOR2_X1 U1076 ( .A(n1219), .B(G116), .ZN(n1337) );
INV_X1 U1077 ( .A(G119), .ZN(n1219) );
XOR2_X1 U1078 ( .A(n1338), .B(n1311), .Z(n1100) );
INV_X1 U1079 ( .A(n1251), .ZN(n1311) );
XOR2_X1 U1080 ( .A(G101), .B(KEYINPUT33), .Z(n1251) );
NAND2_X1 U1081 ( .A1(KEYINPUT53), .A2(n1300), .ZN(n1338) );
XOR2_X1 U1082 ( .A(G104), .B(G107), .Z(n1300) );
endmodule


