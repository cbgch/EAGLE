//Key = 0111000111100001101101110001101111110001110011100001010000110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282;

XOR2_X1 U706 ( .A(G107), .B(n967), .Z(G9) );
NOR2_X1 U707 ( .A1(n968), .A2(n969), .ZN(n967) );
NOR2_X1 U708 ( .A1(n970), .A2(n971), .ZN(G75) );
NOR4_X1 U709 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(n971) );
NOR3_X1 U710 ( .A1(n976), .A2(n977), .A3(n978), .ZN(n975) );
NOR2_X1 U711 ( .A1(n979), .A2(n980), .ZN(n978) );
XOR2_X1 U712 ( .A(KEYINPUT54), .B(n981), .Z(n979) );
NOR2_X1 U713 ( .A1(n982), .A2(n983), .ZN(n977) );
NOR2_X1 U714 ( .A1(n984), .A2(n985), .ZN(n983) );
NOR2_X1 U715 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U716 ( .A1(n988), .A2(n989), .ZN(n987) );
NOR2_X1 U717 ( .A1(n990), .A2(n991), .ZN(n988) );
NOR2_X1 U718 ( .A1(n992), .A2(n993), .ZN(n991) );
NOR2_X1 U719 ( .A1(n994), .A2(n995), .ZN(n992) );
NOR2_X1 U720 ( .A1(n996), .A2(n997), .ZN(n995) );
NOR2_X1 U721 ( .A1(n998), .A2(n999), .ZN(n990) );
NOR2_X1 U722 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR2_X1 U723 ( .A1(n1002), .A2(n999), .ZN(n986) );
NOR2_X1 U724 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NOR2_X1 U725 ( .A1(n993), .A2(n1005), .ZN(n1004) );
NOR2_X1 U726 ( .A1(n1006), .A2(n1007), .ZN(n1003) );
XNOR2_X1 U727 ( .A(KEYINPUT23), .B(n993), .ZN(n1007) );
AND2_X1 U728 ( .A1(n1008), .A2(n981), .ZN(n973) );
NOR4_X1 U729 ( .A1(n985), .A2(n989), .A3(n999), .A4(n993), .ZN(n981) );
INV_X1 U730 ( .A(n1009), .ZN(n993) );
INV_X1 U731 ( .A(n1010), .ZN(n989) );
NAND2_X1 U732 ( .A1(n1011), .A2(n1012), .ZN(n972) );
NOR3_X1 U733 ( .A1(n1013), .A2(G952), .A3(n974), .ZN(n970) );
AND4_X1 U734 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n974) );
NOR4_X1 U735 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
XNOR2_X1 U736 ( .A(G469), .B(n1022), .ZN(n1021) );
NAND2_X1 U737 ( .A1(KEYINPUT32), .A2(n1023), .ZN(n1022) );
XNOR2_X1 U738 ( .A(KEYINPUT13), .B(n1024), .ZN(n1020) );
XNOR2_X1 U739 ( .A(n1025), .B(KEYINPUT62), .ZN(n1018) );
NOR3_X1 U740 ( .A1(n1026), .A2(n982), .A3(n1027), .ZN(n1016) );
NOR2_X1 U741 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
XNOR2_X1 U742 ( .A(n1030), .B(KEYINPUT60), .ZN(n1029) );
XNOR2_X1 U743 ( .A(KEYINPUT30), .B(n1031), .ZN(n1015) );
XOR2_X1 U744 ( .A(KEYINPUT19), .B(n1032), .Z(n1014) );
NOR2_X1 U745 ( .A1(n1030), .A2(n1033), .ZN(n1032) );
INV_X1 U746 ( .A(n1012), .ZN(n1013) );
NAND2_X1 U747 ( .A1(n1034), .A2(n1035), .ZN(G72) );
NAND3_X1 U748 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
XOR2_X1 U749 ( .A(n1039), .B(n1040), .Z(n1038) );
INV_X1 U750 ( .A(KEYINPUT56), .ZN(n1037) );
XNOR2_X1 U751 ( .A(KEYINPUT40), .B(n1041), .ZN(n1036) );
NAND2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1034) );
NAND2_X1 U753 ( .A1(n1044), .A2(n1041), .ZN(n1043) );
NAND2_X1 U754 ( .A1(G953), .A2(n1045), .ZN(n1041) );
NAND2_X1 U755 ( .A1(G900), .A2(G227), .ZN(n1045) );
NAND2_X1 U756 ( .A1(KEYINPUT56), .A2(KEYINPUT40), .ZN(n1044) );
XNOR2_X1 U757 ( .A(n1040), .B(n1039), .ZN(n1042) );
NAND2_X1 U758 ( .A1(n1046), .A2(n1047), .ZN(n1039) );
NAND2_X1 U759 ( .A1(G953), .A2(n1048), .ZN(n1047) );
XNOR2_X1 U760 ( .A(KEYINPUT44), .B(n1049), .ZN(n1048) );
XOR2_X1 U761 ( .A(n1050), .B(n1051), .Z(n1046) );
XNOR2_X1 U762 ( .A(n1052), .B(n1053), .ZN(n1051) );
XNOR2_X1 U763 ( .A(n1054), .B(KEYINPUT57), .ZN(n1050) );
NAND2_X1 U764 ( .A1(n1055), .A2(KEYINPUT45), .ZN(n1054) );
XOR2_X1 U765 ( .A(n1056), .B(n1057), .Z(n1055) );
NAND2_X1 U766 ( .A1(KEYINPUT33), .A2(n1058), .ZN(n1056) );
NAND2_X1 U767 ( .A1(n1059), .A2(n1060), .ZN(n1040) );
XOR2_X1 U768 ( .A(n1061), .B(n1062), .Z(G69) );
NAND2_X1 U769 ( .A1(G953), .A2(n1063), .ZN(n1062) );
NAND2_X1 U770 ( .A1(G898), .A2(G224), .ZN(n1063) );
NAND2_X1 U771 ( .A1(KEYINPUT3), .A2(n1064), .ZN(n1061) );
XOR2_X1 U772 ( .A(n1065), .B(n1066), .Z(n1064) );
NAND2_X1 U773 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XNOR2_X1 U774 ( .A(G953), .B(KEYINPUT20), .ZN(n1067) );
NAND2_X1 U775 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
XOR2_X1 U776 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U777 ( .A1(KEYINPUT27), .A2(n1073), .ZN(n1072) );
NAND2_X1 U778 ( .A1(n1074), .A2(n1075), .ZN(n1071) );
OR2_X1 U779 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U780 ( .A(n1078), .B(KEYINPUT14), .Z(n1074) );
NAND2_X1 U781 ( .A1(n1076), .A2(n1077), .ZN(n1078) );
XOR2_X1 U782 ( .A(G119), .B(n1079), .Z(n1076) );
XOR2_X1 U783 ( .A(n1080), .B(KEYINPUT24), .Z(n1069) );
NAND2_X1 U784 ( .A1(G953), .A2(n1081), .ZN(n1080) );
NOR2_X1 U785 ( .A1(n1082), .A2(n1083), .ZN(G66) );
XOR2_X1 U786 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND3_X1 U787 ( .A1(n1086), .A2(n1030), .A3(KEYINPUT63), .ZN(n1084) );
NOR2_X1 U788 ( .A1(n1082), .A2(n1087), .ZN(G63) );
XOR2_X1 U789 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U790 ( .A1(n1086), .A2(G478), .ZN(n1088) );
NOR2_X1 U791 ( .A1(n1082), .A2(n1090), .ZN(G60) );
XNOR2_X1 U792 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR3_X1 U793 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NOR2_X1 U794 ( .A1(KEYINPUT9), .A2(n1096), .ZN(n1095) );
NOR2_X1 U795 ( .A1(G902), .A2(n1011), .ZN(n1096) );
AND2_X1 U796 ( .A1(n1097), .A2(KEYINPUT9), .ZN(n1094) );
XOR2_X1 U797 ( .A(G104), .B(n1098), .Z(G6) );
NOR2_X1 U798 ( .A1(n969), .A2(n1099), .ZN(n1098) );
NOR2_X1 U799 ( .A1(n1082), .A2(n1100), .ZN(G57) );
XOR2_X1 U800 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U801 ( .A(n1103), .B(n1104), .Z(n1102) );
XNOR2_X1 U802 ( .A(n1105), .B(n1106), .ZN(n1103) );
NOR3_X1 U803 ( .A1(n1097), .A2(KEYINPUT25), .A3(n1107), .ZN(n1106) );
NOR2_X1 U804 ( .A1(KEYINPUT42), .A2(n1108), .ZN(n1105) );
XOR2_X1 U805 ( .A(n1109), .B(n1110), .Z(n1101) );
NOR2_X1 U806 ( .A1(KEYINPUT12), .A2(n1111), .ZN(n1110) );
XOR2_X1 U807 ( .A(n1112), .B(n1113), .Z(n1111) );
XNOR2_X1 U808 ( .A(KEYINPUT1), .B(n1114), .ZN(n1113) );
XNOR2_X1 U809 ( .A(G101), .B(G119), .ZN(n1109) );
NOR2_X1 U810 ( .A1(n1082), .A2(n1115), .ZN(G54) );
XOR2_X1 U811 ( .A(n1116), .B(n1117), .Z(n1115) );
XNOR2_X1 U812 ( .A(n1118), .B(n1119), .ZN(n1117) );
XOR2_X1 U813 ( .A(n1120), .B(n1121), .Z(n1116) );
XOR2_X1 U814 ( .A(KEYINPUT47), .B(n1122), .Z(n1121) );
NAND2_X1 U815 ( .A1(n1086), .A2(G469), .ZN(n1120) );
NOR2_X1 U816 ( .A1(n1082), .A2(n1123), .ZN(G51) );
XOR2_X1 U817 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U818 ( .A1(n1126), .A2(n1097), .ZN(n1125) );
INV_X1 U819 ( .A(n1086), .ZN(n1097) );
NOR2_X1 U820 ( .A1(n1127), .A2(n1011), .ZN(n1086) );
NOR2_X1 U821 ( .A1(n1060), .A2(n1068), .ZN(n1011) );
NAND4_X1 U822 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1068) );
AND4_X1 U823 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1131) );
NAND2_X1 U824 ( .A1(n1008), .A2(n1136), .ZN(n1130) );
NAND2_X1 U825 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XNOR2_X1 U826 ( .A(KEYINPUT58), .B(n1099), .ZN(n1138) );
NAND2_X1 U827 ( .A1(n1139), .A2(n1140), .ZN(n1099) );
XNOR2_X1 U828 ( .A(KEYINPUT34), .B(n968), .ZN(n1137) );
NAND2_X1 U829 ( .A1(n1141), .A2(n1140), .ZN(n968) );
AND3_X1 U830 ( .A1(n994), .A2(n1142), .A3(n1009), .ZN(n1140) );
NAND3_X1 U831 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1128) );
INV_X1 U832 ( .A(n1146), .ZN(n1145) );
NAND2_X1 U833 ( .A1(KEYINPUT7), .A2(n1147), .ZN(n1144) );
NAND2_X1 U834 ( .A1(n1148), .A2(n1149), .ZN(n1143) );
INV_X1 U835 ( .A(KEYINPUT7), .ZN(n1149) );
NAND3_X1 U836 ( .A1(n1142), .A2(n969), .A3(n1150), .ZN(n1148) );
INV_X1 U837 ( .A(n1008), .ZN(n969) );
NAND4_X1 U838 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1060) );
NOR4_X1 U839 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1154) );
INV_X1 U840 ( .A(n1159), .ZN(n1158) );
NOR3_X1 U841 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1153) );
NOR4_X1 U842 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1162) );
INV_X1 U843 ( .A(KEYINPUT37), .ZN(n1163) );
NOR2_X1 U844 ( .A1(KEYINPUT37), .A2(n1167), .ZN(n1161) );
NOR2_X1 U845 ( .A1(n1168), .A2(n1146), .ZN(n1160) );
NAND4_X1 U846 ( .A1(n1169), .A2(n1141), .A3(n1170), .A4(n1171), .ZN(n1151) );
OR2_X1 U847 ( .A1(n1172), .A2(KEYINPUT48), .ZN(n1171) );
NAND2_X1 U848 ( .A1(KEYINPUT48), .A2(n1173), .ZN(n1170) );
NAND3_X1 U849 ( .A1(n1174), .A2(n1175), .A3(n1008), .ZN(n1173) );
NAND2_X1 U850 ( .A1(KEYINPUT59), .A2(n1176), .ZN(n1124) );
XNOR2_X1 U851 ( .A(G125), .B(n1177), .ZN(n1176) );
NOR2_X1 U852 ( .A1(n1059), .A2(G952), .ZN(n1082) );
XOR2_X1 U853 ( .A(G146), .B(n1157), .Z(G48) );
AND3_X1 U854 ( .A1(n1172), .A2(n1139), .A3(n1169), .ZN(n1157) );
NAND2_X1 U855 ( .A1(n1178), .A2(n1179), .ZN(G45) );
NAND2_X1 U856 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U857 ( .A(KEYINPUT41), .B(n1182), .Z(n1178) );
NOR2_X1 U858 ( .A1(n1180), .A2(n1181), .ZN(n1182) );
INV_X1 U859 ( .A(n1167), .ZN(n1180) );
NAND3_X1 U860 ( .A1(n1172), .A2(n1001), .A3(n1165), .ZN(n1167) );
XOR2_X1 U861 ( .A(G140), .B(n1156), .Z(G42) );
NOR3_X1 U862 ( .A1(n1005), .A2(n1168), .A3(n1183), .ZN(n1156) );
XNOR2_X1 U863 ( .A(n1058), .B(n1184), .ZN(G39) );
NOR3_X1 U864 ( .A1(n1146), .A2(KEYINPUT29), .A3(n1168), .ZN(n1184) );
XNOR2_X1 U865 ( .A(G134), .B(n1152), .ZN(G36) );
OR3_X1 U866 ( .A1(n1168), .A2(n1006), .A3(n1166), .ZN(n1152) );
INV_X1 U867 ( .A(n1141), .ZN(n1006) );
XOR2_X1 U868 ( .A(n1155), .B(n1185), .Z(G33) );
XOR2_X1 U869 ( .A(KEYINPUT61), .B(G131), .Z(n1185) );
NOR3_X1 U870 ( .A1(n1166), .A2(n1168), .A3(n1005), .ZN(n1155) );
INV_X1 U871 ( .A(n1139), .ZN(n1005) );
NAND4_X1 U872 ( .A1(n1024), .A2(n994), .A3(n1174), .A4(n980), .ZN(n1168) );
INV_X1 U873 ( .A(n982), .ZN(n980) );
XNOR2_X1 U874 ( .A(G128), .B(n1186), .ZN(G30) );
NAND3_X1 U875 ( .A1(n1172), .A2(n1141), .A3(n1169), .ZN(n1186) );
INV_X1 U876 ( .A(n1164), .ZN(n1172) );
NAND3_X1 U877 ( .A1(n994), .A2(n1174), .A3(n1008), .ZN(n1164) );
XNOR2_X1 U878 ( .A(G101), .B(n1135), .ZN(G3) );
NAND3_X1 U879 ( .A1(n1001), .A2(n994), .A3(n1187), .ZN(n1135) );
XNOR2_X1 U880 ( .A(G125), .B(n1159), .ZN(G27) );
NAND4_X1 U881 ( .A1(n1008), .A2(n1174), .A3(n1139), .A4(n1188), .ZN(n1159) );
NOR2_X1 U882 ( .A1(n1183), .A2(n999), .ZN(n1188) );
INV_X1 U883 ( .A(n1150), .ZN(n999) );
INV_X1 U884 ( .A(n1000), .ZN(n1183) );
NAND2_X1 U885 ( .A1(n985), .A2(n1189), .ZN(n1174) );
NAND4_X1 U886 ( .A1(G953), .A2(G902), .A3(n1190), .A4(n1049), .ZN(n1189) );
INV_X1 U887 ( .A(G900), .ZN(n1049) );
XNOR2_X1 U888 ( .A(G122), .B(n1129), .ZN(G24) );
NAND3_X1 U889 ( .A1(n1165), .A2(n1009), .A3(n1191), .ZN(n1129) );
NOR2_X1 U890 ( .A1(n1019), .A2(n1192), .ZN(n1009) );
INV_X1 U891 ( .A(n1193), .ZN(n1192) );
NOR2_X1 U892 ( .A1(n1194), .A2(n1031), .ZN(n1165) );
XNOR2_X1 U893 ( .A(n1195), .B(n1196), .ZN(G21) );
NOR2_X1 U894 ( .A1(n1146), .A2(n1147), .ZN(n1196) );
NAND2_X1 U895 ( .A1(n1010), .A2(n1169), .ZN(n1146) );
NOR2_X1 U896 ( .A1(n1193), .A2(n1197), .ZN(n1169) );
INV_X1 U897 ( .A(n1019), .ZN(n1197) );
XNOR2_X1 U898 ( .A(G116), .B(n1134), .ZN(G18) );
NAND3_X1 U899 ( .A1(n1001), .A2(n1141), .A3(n1191), .ZN(n1134) );
NOR2_X1 U900 ( .A1(n1198), .A2(n1194), .ZN(n1141) );
INV_X1 U901 ( .A(n1025), .ZN(n1194) );
XOR2_X1 U902 ( .A(n1199), .B(G113), .Z(G15) );
NAND2_X1 U903 ( .A1(KEYINPUT51), .A2(n1133), .ZN(n1199) );
NAND3_X1 U904 ( .A1(n1139), .A2(n1001), .A3(n1191), .ZN(n1133) );
INV_X1 U905 ( .A(n1147), .ZN(n1191) );
NAND3_X1 U906 ( .A1(n1008), .A2(n1142), .A3(n1150), .ZN(n1147) );
NOR2_X1 U907 ( .A1(n996), .A2(n1027), .ZN(n1150) );
INV_X1 U908 ( .A(n997), .ZN(n1027) );
INV_X1 U909 ( .A(n1166), .ZN(n1001) );
NAND2_X1 U910 ( .A1(n1200), .A2(n1019), .ZN(n1166) );
XNOR2_X1 U911 ( .A(n1193), .B(KEYINPUT18), .ZN(n1200) );
NOR2_X1 U912 ( .A1(n1025), .A2(n1031), .ZN(n1139) );
INV_X1 U913 ( .A(n1198), .ZN(n1031) );
XNOR2_X1 U914 ( .A(G110), .B(n1132), .ZN(G12) );
NAND3_X1 U915 ( .A1(n1000), .A2(n994), .A3(n1187), .ZN(n1132) );
AND3_X1 U916 ( .A1(n1008), .A2(n1142), .A3(n1010), .ZN(n1187) );
NOR2_X1 U917 ( .A1(n1025), .A2(n1198), .ZN(n1010) );
XOR2_X1 U918 ( .A(n1201), .B(n1093), .Z(n1198) );
INV_X1 U919 ( .A(G475), .ZN(n1093) );
NAND2_X1 U920 ( .A1(n1202), .A2(n1091), .ZN(n1201) );
XNOR2_X1 U921 ( .A(n1203), .B(n1204), .ZN(n1091) );
XNOR2_X1 U922 ( .A(n1181), .B(n1205), .ZN(n1204) );
XOR2_X1 U923 ( .A(KEYINPUT52), .B(G146), .Z(n1205) );
XNOR2_X1 U924 ( .A(n1206), .B(n1207), .ZN(n1203) );
INV_X1 U925 ( .A(n1053), .ZN(n1207) );
XOR2_X1 U926 ( .A(G131), .B(n1208), .Z(n1053) );
XOR2_X1 U927 ( .A(n1209), .B(n1210), .Z(n1206) );
NOR3_X1 U928 ( .A1(n1211), .A2(G953), .A3(G237), .ZN(n1210) );
NAND2_X1 U929 ( .A1(n1212), .A2(n1213), .ZN(n1209) );
NAND2_X1 U930 ( .A1(n1214), .A2(G104), .ZN(n1213) );
XOR2_X1 U931 ( .A(n1215), .B(KEYINPUT36), .Z(n1212) );
OR2_X1 U932 ( .A1(n1214), .A2(G104), .ZN(n1215) );
XOR2_X1 U933 ( .A(G113), .B(n1216), .Z(n1214) );
XNOR2_X1 U934 ( .A(n1217), .B(KEYINPUT39), .ZN(n1202) );
XNOR2_X1 U935 ( .A(n1218), .B(G478), .ZN(n1025) );
NAND2_X1 U936 ( .A1(n1089), .A2(n1217), .ZN(n1218) );
XNOR2_X1 U937 ( .A(n1219), .B(n1220), .ZN(n1089) );
XOR2_X1 U938 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U939 ( .A(n1223), .B(n1224), .ZN(n1222) );
NAND2_X1 U940 ( .A1(KEYINPUT2), .A2(n1225), .ZN(n1224) );
NAND3_X1 U941 ( .A1(G217), .A2(n1226), .A3(KEYINPUT16), .ZN(n1223) );
XNOR2_X1 U942 ( .A(G107), .B(KEYINPUT55), .ZN(n1221) );
XOR2_X1 U943 ( .A(n1216), .B(n1227), .Z(n1219) );
XOR2_X1 U944 ( .A(n1057), .B(n1228), .Z(n1227) );
NAND2_X1 U945 ( .A1(n985), .A2(n1229), .ZN(n1142) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1190), .A4(n1081), .ZN(n1229) );
INV_X1 U947 ( .A(G898), .ZN(n1081) );
NAND3_X1 U948 ( .A1(n1012), .A2(n1190), .A3(G952), .ZN(n985) );
NAND2_X1 U949 ( .A1(G237), .A2(G234), .ZN(n1190) );
XOR2_X1 U950 ( .A(G953), .B(KEYINPUT22), .Z(n1012) );
NOR2_X1 U951 ( .A1(n1024), .A2(n982), .ZN(n1008) );
NOR2_X1 U952 ( .A1(n1211), .A2(n1230), .ZN(n982) );
INV_X1 U953 ( .A(G214), .ZN(n1211) );
INV_X1 U954 ( .A(n976), .ZN(n1024) );
XNOR2_X1 U955 ( .A(n1231), .B(n1232), .ZN(n976) );
NOR2_X1 U956 ( .A1(n1230), .A2(n1233), .ZN(n1232) );
XNOR2_X1 U957 ( .A(KEYINPUT46), .B(n1126), .ZN(n1233) );
NOR2_X1 U958 ( .A1(G902), .A2(G237), .ZN(n1230) );
NAND2_X1 U959 ( .A1(n1234), .A2(n1217), .ZN(n1231) );
XNOR2_X1 U960 ( .A(n1235), .B(n1177), .ZN(n1234) );
XOR2_X1 U961 ( .A(n1236), .B(n1237), .Z(n1177) );
XOR2_X1 U962 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U963 ( .A(KEYINPUT10), .B(n1240), .Z(n1239) );
AND2_X1 U964 ( .A1(n1059), .A2(G224), .ZN(n1240) );
NOR2_X1 U965 ( .A1(KEYINPUT5), .A2(n1241), .ZN(n1238) );
XOR2_X1 U966 ( .A(n1242), .B(n1073), .Z(n1236) );
XNOR2_X1 U967 ( .A(G110), .B(n1216), .ZN(n1073) );
XNOR2_X1 U968 ( .A(G122), .B(KEYINPUT28), .ZN(n1216) );
XOR2_X1 U969 ( .A(n1243), .B(n1079), .Z(n1242) );
XNOR2_X1 U970 ( .A(n1225), .B(n1244), .ZN(n1079) );
NOR2_X1 U971 ( .A1(KEYINPUT4), .A2(n1245), .ZN(n1244) );
XOR2_X1 U972 ( .A(KEYINPUT53), .B(G113), .Z(n1245) );
INV_X1 U973 ( .A(G116), .ZN(n1225) );
NAND2_X1 U974 ( .A1(KEYINPUT31), .A2(n1246), .ZN(n1235) );
INV_X1 U975 ( .A(n1175), .ZN(n994) );
NAND2_X1 U976 ( .A1(n996), .A2(n997), .ZN(n1175) );
NAND2_X1 U977 ( .A1(G221), .A2(n1247), .ZN(n997) );
XOR2_X1 U978 ( .A(n1023), .B(G469), .Z(n996) );
AND2_X1 U979 ( .A1(n1248), .A2(n1217), .ZN(n1023) );
XNOR2_X1 U980 ( .A(n1249), .B(n1114), .ZN(n1248) );
XNOR2_X1 U981 ( .A(n1250), .B(n1251), .ZN(n1249) );
NOR2_X1 U982 ( .A1(KEYINPUT38), .A2(n1119), .ZN(n1251) );
XNOR2_X1 U983 ( .A(n1252), .B(n1241), .ZN(n1119) );
INV_X1 U984 ( .A(n1077), .ZN(n1241) );
XOR2_X1 U985 ( .A(G101), .B(n1253), .Z(n1077) );
XOR2_X1 U986 ( .A(G107), .B(G104), .Z(n1253) );
XOR2_X1 U987 ( .A(n1052), .B(KEYINPUT43), .Z(n1252) );
XOR2_X1 U988 ( .A(n1112), .B(KEYINPUT15), .Z(n1052) );
NOR2_X1 U989 ( .A1(n1122), .A2(KEYINPUT0), .ZN(n1250) );
AND2_X1 U990 ( .A1(n1254), .A2(n1255), .ZN(n1122) );
NAND3_X1 U991 ( .A1(G227), .A2(n1059), .A3(n1256), .ZN(n1255) );
XNOR2_X1 U992 ( .A(G110), .B(G140), .ZN(n1256) );
NAND2_X1 U993 ( .A1(n1257), .A2(n1258), .ZN(n1254) );
NAND2_X1 U994 ( .A1(G227), .A2(n1059), .ZN(n1258) );
XNOR2_X1 U995 ( .A(G140), .B(n1259), .ZN(n1257) );
NOR2_X1 U996 ( .A1(n1193), .A2(n1019), .ZN(n1000) );
XOR2_X1 U997 ( .A(n1260), .B(n1107), .Z(n1019) );
INV_X1 U998 ( .A(G472), .ZN(n1107) );
NAND2_X1 U999 ( .A1(n1261), .A2(n1217), .ZN(n1260) );
XOR2_X1 U1000 ( .A(n1262), .B(n1263), .Z(n1261) );
NOR2_X1 U1001 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
XOR2_X1 U1002 ( .A(n1266), .B(KEYINPUT35), .Z(n1265) );
NAND2_X1 U1003 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NOR2_X1 U1004 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
INV_X1 U1005 ( .A(n1108), .ZN(n1268) );
NOR3_X1 U1006 ( .A1(G237), .A2(G953), .A3(n1126), .ZN(n1108) );
INV_X1 U1007 ( .A(G210), .ZN(n1126) );
INV_X1 U1008 ( .A(G101), .ZN(n1267) );
NAND2_X1 U1009 ( .A1(KEYINPUT21), .A2(n1269), .ZN(n1262) );
XNOR2_X1 U1010 ( .A(n1104), .B(n1270), .ZN(n1269) );
XNOR2_X1 U1011 ( .A(n1243), .B(n1114), .ZN(n1270) );
INV_X1 U1012 ( .A(n1118), .ZN(n1114) );
XNOR2_X1 U1013 ( .A(n1271), .B(n1057), .ZN(n1118) );
XOR2_X1 U1014 ( .A(G134), .B(KEYINPUT50), .Z(n1057) );
XNOR2_X1 U1015 ( .A(G131), .B(G137), .ZN(n1271) );
XNOR2_X1 U1016 ( .A(n1112), .B(n1195), .ZN(n1243) );
XNOR2_X1 U1017 ( .A(G146), .B(n1228), .ZN(n1112) );
XNOR2_X1 U1018 ( .A(G128), .B(n1181), .ZN(n1228) );
INV_X1 U1019 ( .A(G143), .ZN(n1181) );
XOR2_X1 U1020 ( .A(G113), .B(n1272), .Z(n1104) );
NOR2_X1 U1021 ( .A1(G116), .A2(KEYINPUT11), .ZN(n1272) );
XOR2_X1 U1022 ( .A(n1028), .B(n1273), .Z(n1193) );
NOR2_X1 U1023 ( .A1(n1030), .A2(KEYINPUT6), .ZN(n1273) );
AND2_X1 U1024 ( .A1(G217), .A2(n1247), .ZN(n1030) );
NAND2_X1 U1025 ( .A1(G234), .A2(n1127), .ZN(n1247) );
INV_X1 U1026 ( .A(G902), .ZN(n1127) );
INV_X1 U1027 ( .A(n1033), .ZN(n1028) );
NAND2_X1 U1028 ( .A1(n1274), .A2(n1217), .ZN(n1033) );
XOR2_X1 U1029 ( .A(G902), .B(KEYINPUT8), .Z(n1217) );
XOR2_X1 U1030 ( .A(KEYINPUT26), .B(n1085), .Z(n1274) );
XNOR2_X1 U1031 ( .A(n1275), .B(n1276), .ZN(n1085) );
XNOR2_X1 U1032 ( .A(n1058), .B(n1277), .ZN(n1276) );
NOR2_X1 U1033 ( .A1(KEYINPUT17), .A2(n1278), .ZN(n1277) );
XOR2_X1 U1034 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U1035 ( .A(n1281), .B(n1208), .Z(n1280) );
XNOR2_X1 U1036 ( .A(n1246), .B(G140), .ZN(n1208) );
INV_X1 U1037 ( .A(G125), .ZN(n1246) );
NOR2_X1 U1038 ( .A1(G146), .A2(KEYINPUT49), .ZN(n1281) );
XNOR2_X1 U1039 ( .A(n1259), .B(n1282), .ZN(n1279) );
XNOR2_X1 U1040 ( .A(G128), .B(n1195), .ZN(n1282) );
INV_X1 U1041 ( .A(G119), .ZN(n1195) );
INV_X1 U1042 ( .A(G110), .ZN(n1259) );
INV_X1 U1043 ( .A(G137), .ZN(n1058) );
NAND2_X1 U1044 ( .A1(G221), .A2(n1226), .ZN(n1275) );
AND2_X1 U1045 ( .A1(G234), .A2(n1059), .ZN(n1226) );
INV_X1 U1046 ( .A(G953), .ZN(n1059) );
endmodule


