//Key = 1101001111000100101000100110000010101011010001100001111011101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421, n1422, n1423, n1424, n1425;

XNOR2_X1 U777 ( .A(G107), .B(n1079), .ZN(G9) );
NAND3_X1 U778 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NOR2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(G75) );
NOR3_X1 U780 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NOR4_X1 U781 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1086) );
NOR2_X1 U782 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NOR3_X1 U784 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1092) );
NOR3_X1 U785 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
NOR2_X1 U786 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NOR2_X1 U787 ( .A1(n1104), .A2(n1081), .ZN(n1097) );
NAND3_X1 U788 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1085) );
NAND4_X1 U789 ( .A1(n1108), .A2(n1109), .A3(n1104), .A4(n1110), .ZN(n1107) );
NOR2_X1 U790 ( .A1(n1099), .A2(n1096), .ZN(n1110) );
NAND2_X1 U791 ( .A1(n1111), .A2(n1091), .ZN(n1109) );
NAND3_X1 U792 ( .A1(n1112), .A2(n1082), .A3(KEYINPUT62), .ZN(n1111) );
NAND3_X1 U793 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1108) );
INV_X1 U794 ( .A(n1091), .ZN(n1115) );
NAND2_X1 U795 ( .A1(n1112), .A2(n1116), .ZN(n1114) );
NAND2_X1 U796 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
OR2_X1 U797 ( .A1(n1119), .A2(KEYINPUT62), .ZN(n1118) );
NAND2_X1 U798 ( .A1(n1120), .A2(n1121), .ZN(n1113) );
NAND3_X1 U799 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
NAND2_X1 U800 ( .A1(KEYINPUT21), .A2(n1125), .ZN(n1123) );
OR3_X1 U801 ( .A1(n1126), .A2(KEYINPUT21), .A3(n1125), .ZN(n1122) );
NOR3_X1 U802 ( .A1(n1127), .A2(G953), .A3(G952), .ZN(n1083) );
INV_X1 U803 ( .A(n1105), .ZN(n1127) );
NAND4_X1 U804 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1105) );
NOR4_X1 U805 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1131) );
XNOR2_X1 U806 ( .A(n1136), .B(n1137), .ZN(n1134) );
XNOR2_X1 U807 ( .A(KEYINPUT32), .B(n1138), .ZN(n1137) );
INV_X1 U808 ( .A(n1126), .ZN(n1132) );
NOR2_X1 U809 ( .A1(n1139), .A2(n1140), .ZN(n1130) );
XNOR2_X1 U810 ( .A(G472), .B(n1141), .ZN(n1140) );
XNOR2_X1 U811 ( .A(G469), .B(n1142), .ZN(n1139) );
XOR2_X1 U812 ( .A(n1143), .B(n1144), .Z(n1129) );
XOR2_X1 U813 ( .A(KEYINPUT5), .B(KEYINPUT17), .Z(n1144) );
XNOR2_X1 U814 ( .A(n1145), .B(n1146), .ZN(n1128) );
NAND2_X1 U815 ( .A1(n1147), .A2(n1148), .ZN(G72) );
NAND2_X1 U816 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
OR2_X1 U817 ( .A1(n1106), .A2(G227), .ZN(n1150) );
NAND3_X1 U818 ( .A1(G953), .A2(n1151), .A3(n1152), .ZN(n1147) );
INV_X1 U819 ( .A(n1149), .ZN(n1152) );
XNOR2_X1 U820 ( .A(n1153), .B(n1154), .ZN(n1149) );
NOR2_X1 U821 ( .A1(n1155), .A2(G953), .ZN(n1154) );
NOR2_X1 U822 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U823 ( .A1(n1158), .A2(n1159), .ZN(n1153) );
NAND2_X1 U824 ( .A1(G953), .A2(n1160), .ZN(n1159) );
XOR2_X1 U825 ( .A(KEYINPUT50), .B(n1161), .Z(n1158) );
NOR2_X1 U826 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U827 ( .A(n1164), .B(KEYINPUT52), .Z(n1163) );
NAND2_X1 U828 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NOR2_X1 U829 ( .A1(n1167), .A2(n1165), .ZN(n1162) );
XOR2_X1 U830 ( .A(n1168), .B(n1169), .Z(n1165) );
NAND2_X1 U831 ( .A1(n1170), .A2(n1171), .ZN(n1168) );
NAND2_X1 U832 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
XOR2_X1 U833 ( .A(KEYINPUT41), .B(n1174), .Z(n1172) );
NAND2_X1 U834 ( .A1(n1174), .A2(G137), .ZN(n1170) );
XOR2_X1 U835 ( .A(KEYINPUT20), .B(n1166), .Z(n1167) );
XNOR2_X1 U836 ( .A(n1175), .B(G140), .ZN(n1166) );
NAND2_X1 U837 ( .A1(KEYINPUT25), .A2(G125), .ZN(n1175) );
NAND2_X1 U838 ( .A1(G900), .A2(G227), .ZN(n1151) );
XOR2_X1 U839 ( .A(n1176), .B(n1177), .Z(G69) );
NAND2_X1 U840 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
OR3_X1 U841 ( .A1(n1106), .A2(G224), .A3(n1180), .ZN(n1179) );
NAND2_X1 U842 ( .A1(n1181), .A2(n1180), .ZN(n1178) );
OR2_X1 U843 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
XNOR2_X1 U844 ( .A(n1184), .B(n1185), .ZN(n1182) );
XNOR2_X1 U845 ( .A(n1186), .B(n1187), .ZN(n1185) );
NOR2_X1 U846 ( .A1(KEYINPUT49), .A2(n1188), .ZN(n1187) );
NOR2_X1 U847 ( .A1(KEYINPUT11), .A2(n1189), .ZN(n1186) );
NAND2_X1 U848 ( .A1(G953), .A2(n1190), .ZN(n1181) );
NAND2_X1 U849 ( .A1(G898), .A2(G224), .ZN(n1190) );
NAND2_X1 U850 ( .A1(n1106), .A2(n1191), .ZN(n1176) );
NAND2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XNOR2_X1 U852 ( .A(n1194), .B(KEYINPUT31), .ZN(n1192) );
NOR2_X1 U853 ( .A1(n1195), .A2(n1196), .ZN(G66) );
NOR3_X1 U854 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
NOR3_X1 U855 ( .A1(n1200), .A2(n1201), .A3(n1202), .ZN(n1199) );
INV_X1 U856 ( .A(n1203), .ZN(n1200) );
NOR2_X1 U857 ( .A1(n1204), .A2(n1203), .ZN(n1198) );
NOR2_X1 U858 ( .A1(n1205), .A2(n1201), .ZN(n1204) );
NOR2_X1 U859 ( .A1(n1195), .A2(n1206), .ZN(G63) );
XOR2_X1 U860 ( .A(n1207), .B(n1208), .Z(n1206) );
NAND3_X1 U861 ( .A1(n1209), .A2(n1210), .A3(G478), .ZN(n1207) );
NAND2_X1 U862 ( .A1(KEYINPUT61), .A2(n1202), .ZN(n1210) );
NAND2_X1 U863 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
INV_X1 U864 ( .A(KEYINPUT61), .ZN(n1212) );
NAND2_X1 U865 ( .A1(n1205), .A2(G902), .ZN(n1211) );
NOR2_X1 U866 ( .A1(n1195), .A2(n1213), .ZN(G60) );
NOR3_X1 U867 ( .A1(n1136), .A2(n1214), .A3(n1215), .ZN(n1213) );
NOR3_X1 U868 ( .A1(n1216), .A2(n1138), .A3(n1202), .ZN(n1215) );
INV_X1 U869 ( .A(n1217), .ZN(n1216) );
NOR2_X1 U870 ( .A1(n1218), .A2(n1217), .ZN(n1214) );
NOR2_X1 U871 ( .A1(n1205), .A2(n1138), .ZN(n1218) );
INV_X1 U872 ( .A(n1087), .ZN(n1205) );
XNOR2_X1 U873 ( .A(G104), .B(n1219), .ZN(G6) );
NOR2_X1 U874 ( .A1(n1195), .A2(n1220), .ZN(G57) );
XOR2_X1 U875 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U876 ( .A(n1223), .B(n1224), .ZN(n1222) );
XOR2_X1 U877 ( .A(n1225), .B(n1226), .Z(n1221) );
XOR2_X1 U878 ( .A(n1227), .B(n1228), .Z(n1226) );
NOR2_X1 U879 ( .A1(KEYINPUT28), .A2(n1229), .ZN(n1228) );
NOR2_X1 U880 ( .A1(n1230), .A2(n1202), .ZN(n1225) );
INV_X1 U881 ( .A(G472), .ZN(n1230) );
NOR2_X1 U882 ( .A1(n1195), .A2(n1231), .ZN(G54) );
XOR2_X1 U883 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U884 ( .A(n1234), .B(n1235), .Z(n1233) );
XNOR2_X1 U885 ( .A(n1236), .B(G110), .ZN(n1235) );
NOR2_X1 U886 ( .A1(n1237), .A2(n1202), .ZN(n1234) );
INV_X1 U887 ( .A(G469), .ZN(n1237) );
XOR2_X1 U888 ( .A(n1238), .B(n1239), .Z(n1232) );
NOR2_X1 U889 ( .A1(n1240), .A2(KEYINPUT4), .ZN(n1239) );
NAND2_X1 U890 ( .A1(KEYINPUT16), .A2(n1241), .ZN(n1238) );
NOR2_X1 U891 ( .A1(n1195), .A2(n1242), .ZN(G51) );
XOR2_X1 U892 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U893 ( .A(n1245), .B(n1246), .Z(n1244) );
XOR2_X1 U894 ( .A(G125), .B(n1247), .Z(n1246) );
NOR2_X1 U895 ( .A1(KEYINPUT37), .A2(n1248), .ZN(n1247) );
NOR2_X1 U896 ( .A1(n1146), .A2(n1202), .ZN(n1245) );
NAND2_X1 U897 ( .A1(G902), .A2(n1087), .ZN(n1202) );
NAND4_X1 U898 ( .A1(n1249), .A2(n1193), .A3(n1250), .A4(n1251), .ZN(n1087) );
INV_X1 U899 ( .A(n1157), .ZN(n1250) );
NAND4_X1 U900 ( .A1(n1252), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1157) );
NAND3_X1 U901 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1253) );
XNOR2_X1 U902 ( .A(KEYINPUT48), .B(n1259), .ZN(n1257) );
NAND2_X1 U903 ( .A1(n1260), .A2(n1104), .ZN(n1252) );
XNOR2_X1 U904 ( .A(n1261), .B(KEYINPUT9), .ZN(n1260) );
AND4_X1 U905 ( .A1(n1262), .A2(n1263), .A3(n1219), .A4(n1264), .ZN(n1193) );
AND4_X1 U906 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1264) );
NAND3_X1 U907 ( .A1(n1080), .A2(n1081), .A3(n1269), .ZN(n1219) );
NAND4_X1 U908 ( .A1(n1082), .A2(n1270), .A3(n1271), .A4(n1081), .ZN(n1262) );
XNOR2_X1 U909 ( .A(KEYINPUT39), .B(n1272), .ZN(n1271) );
XOR2_X1 U910 ( .A(n1156), .B(KEYINPUT1), .Z(n1249) );
NAND4_X1 U911 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1156) );
NAND2_X1 U912 ( .A1(n1082), .A2(n1277), .ZN(n1274) );
NAND2_X1 U913 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NAND3_X1 U914 ( .A1(n1280), .A2(n1259), .A3(KEYINPUT35), .ZN(n1279) );
NAND2_X1 U915 ( .A1(n1258), .A2(n1104), .ZN(n1278) );
OR2_X1 U916 ( .A1(n1281), .A2(KEYINPUT35), .ZN(n1273) );
XNOR2_X1 U917 ( .A(n1282), .B(n1223), .ZN(n1243) );
NOR2_X1 U918 ( .A1(n1106), .A2(G952), .ZN(n1195) );
XNOR2_X1 U919 ( .A(G146), .B(n1254), .ZN(G48) );
NAND3_X1 U920 ( .A1(n1269), .A2(n1100), .A3(n1280), .ZN(n1254) );
XOR2_X1 U921 ( .A(G143), .B(n1283), .Z(G45) );
NOR3_X1 U922 ( .A1(n1284), .A2(n1285), .A3(n1259), .ZN(n1283) );
XNOR2_X1 U923 ( .A(n1256), .B(KEYINPUT14), .ZN(n1285) );
XNOR2_X1 U924 ( .A(G140), .B(n1286), .ZN(G42) );
NAND2_X1 U925 ( .A1(n1261), .A2(n1104), .ZN(n1286) );
AND2_X1 U926 ( .A1(n1287), .A2(n1288), .ZN(n1261) );
XNOR2_X1 U927 ( .A(n1289), .B(n1255), .ZN(G39) );
NAND3_X1 U928 ( .A1(n1104), .A2(n1120), .A3(n1280), .ZN(n1255) );
XNOR2_X1 U929 ( .A(G137), .B(KEYINPUT34), .ZN(n1289) );
XOR2_X1 U930 ( .A(G134), .B(n1290), .Z(G36) );
NOR4_X1 U931 ( .A1(KEYINPUT59), .A2(n1119), .A3(n1095), .A4(n1284), .ZN(n1290) );
INV_X1 U932 ( .A(n1104), .ZN(n1095) );
XOR2_X1 U933 ( .A(n1275), .B(n1291), .Z(G33) );
XNOR2_X1 U934 ( .A(G131), .B(KEYINPUT42), .ZN(n1291) );
NAND3_X1 U935 ( .A1(n1104), .A2(n1269), .A3(n1258), .ZN(n1275) );
INV_X1 U936 ( .A(n1284), .ZN(n1258) );
NAND3_X1 U937 ( .A1(n1288), .A2(n1292), .A3(n1293), .ZN(n1284) );
NOR2_X1 U938 ( .A1(n1102), .A2(n1133), .ZN(n1104) );
INV_X1 U939 ( .A(n1103), .ZN(n1133) );
NAND3_X1 U940 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(G30) );
NAND2_X1 U941 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
NAND2_X1 U942 ( .A1(KEYINPUT19), .A2(n1299), .ZN(n1295) );
NAND2_X1 U943 ( .A1(n1300), .A2(G128), .ZN(n1299) );
XNOR2_X1 U944 ( .A(KEYINPUT23), .B(n1297), .ZN(n1300) );
NAND2_X1 U945 ( .A1(n1301), .A2(n1302), .ZN(n1294) );
INV_X1 U946 ( .A(KEYINPUT19), .ZN(n1302) );
NAND2_X1 U947 ( .A1(n1303), .A2(n1304), .ZN(n1301) );
OR3_X1 U948 ( .A1(n1298), .A2(n1297), .A3(KEYINPUT23), .ZN(n1304) );
NAND2_X1 U949 ( .A1(KEYINPUT23), .A2(n1297), .ZN(n1303) );
INV_X1 U950 ( .A(n1281), .ZN(n1297) );
NAND3_X1 U951 ( .A1(n1082), .A2(n1100), .A3(n1280), .ZN(n1281) );
AND4_X1 U952 ( .A1(n1099), .A2(n1288), .A3(n1305), .A4(n1292), .ZN(n1280) );
XNOR2_X1 U953 ( .A(n1263), .B(n1306), .ZN(G3) );
NOR2_X1 U954 ( .A1(KEYINPUT63), .A2(n1307), .ZN(n1306) );
NAND4_X1 U955 ( .A1(n1120), .A2(n1293), .A3(n1308), .A4(n1288), .ZN(n1263) );
INV_X1 U956 ( .A(n1124), .ZN(n1288) );
AND2_X1 U957 ( .A1(n1272), .A2(n1100), .ZN(n1308) );
XNOR2_X1 U958 ( .A(G125), .B(n1276), .ZN(G27) );
NAND3_X1 U959 ( .A1(n1112), .A2(n1100), .A3(n1287), .ZN(n1276) );
AND4_X1 U960 ( .A1(n1099), .A2(n1269), .A3(n1309), .A4(n1292), .ZN(n1287) );
NAND2_X1 U961 ( .A1(n1091), .A2(n1310), .ZN(n1292) );
NAND4_X1 U962 ( .A1(G902), .A2(G953), .A3(n1311), .A4(n1160), .ZN(n1310) );
INV_X1 U963 ( .A(G900), .ZN(n1160) );
XNOR2_X1 U964 ( .A(G122), .B(n1268), .ZN(G24) );
NAND4_X1 U965 ( .A1(n1256), .A2(n1312), .A3(n1309), .A4(n1081), .ZN(n1268) );
INV_X1 U966 ( .A(n1096), .ZN(n1309) );
AND2_X1 U967 ( .A1(n1313), .A2(n1314), .ZN(n1256) );
XNOR2_X1 U968 ( .A(G119), .B(n1267), .ZN(G21) );
NAND4_X1 U969 ( .A1(n1099), .A2(n1120), .A3(n1305), .A4(n1312), .ZN(n1267) );
XOR2_X1 U970 ( .A(n1266), .B(n1315), .Z(G18) );
NAND2_X1 U971 ( .A1(KEYINPUT36), .A2(G116), .ZN(n1315) );
NAND3_X1 U972 ( .A1(n1293), .A2(n1082), .A3(n1312), .ZN(n1266) );
INV_X1 U973 ( .A(n1119), .ZN(n1082) );
NAND2_X1 U974 ( .A1(n1316), .A2(n1317), .ZN(n1119) );
XOR2_X1 U975 ( .A(KEYINPUT15), .B(n1314), .Z(n1316) );
XNOR2_X1 U976 ( .A(n1143), .B(KEYINPUT24), .ZN(n1314) );
XNOR2_X1 U977 ( .A(G113), .B(n1265), .ZN(G15) );
NAND3_X1 U978 ( .A1(n1293), .A2(n1269), .A3(n1312), .ZN(n1265) );
AND3_X1 U979 ( .A1(n1100), .A2(n1272), .A3(n1112), .ZN(n1312) );
INV_X1 U980 ( .A(n1089), .ZN(n1112) );
NAND2_X1 U981 ( .A1(n1318), .A2(n1126), .ZN(n1089) );
XNOR2_X1 U982 ( .A(KEYINPUT21), .B(n1125), .ZN(n1318) );
INV_X1 U983 ( .A(n1259), .ZN(n1100) );
INV_X1 U984 ( .A(n1117), .ZN(n1269) );
NAND2_X1 U985 ( .A1(n1313), .A2(n1143), .ZN(n1117) );
INV_X1 U986 ( .A(n1317), .ZN(n1313) );
INV_X1 U987 ( .A(n1094), .ZN(n1293) );
NAND2_X1 U988 ( .A1(n1305), .A2(n1081), .ZN(n1094) );
XNOR2_X1 U989 ( .A(G110), .B(n1319), .ZN(G12) );
NAND2_X1 U990 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U991 ( .A1(KEYINPUT55), .A2(n1194), .ZN(n1321) );
OR2_X1 U992 ( .A1(KEYINPUT43), .A2(n1194), .ZN(n1320) );
INV_X1 U993 ( .A(n1251), .ZN(n1194) );
NAND3_X1 U994 ( .A1(n1099), .A2(n1080), .A3(n1120), .ZN(n1251) );
INV_X1 U995 ( .A(n1090), .ZN(n1120) );
NAND2_X1 U996 ( .A1(n1143), .A2(n1317), .ZN(n1090) );
XOR2_X1 U997 ( .A(n1322), .B(n1323), .Z(n1317) );
INV_X1 U998 ( .A(n1136), .ZN(n1323) );
NOR2_X1 U999 ( .A1(n1217), .A2(G902), .ZN(n1136) );
XNOR2_X1 U1000 ( .A(n1324), .B(n1325), .ZN(n1217) );
XOR2_X1 U1001 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1002 ( .A(n1328), .B(n1329), .Z(n1327) );
NOR2_X1 U1003 ( .A1(KEYINPUT47), .A2(n1330), .ZN(n1329) );
NAND2_X1 U1004 ( .A1(G214), .A2(n1331), .ZN(n1328) );
XOR2_X1 U1005 ( .A(n1332), .B(n1333), .Z(n1324) );
XNOR2_X1 U1006 ( .A(G131), .B(n1334), .ZN(n1333) );
XNOR2_X1 U1007 ( .A(G104), .B(G113), .ZN(n1332) );
NAND2_X1 U1008 ( .A1(KEYINPUT3), .A2(n1138), .ZN(n1322) );
INV_X1 U1009 ( .A(G475), .ZN(n1138) );
XOR2_X1 U1010 ( .A(n1335), .B(G478), .Z(n1143) );
NAND2_X1 U1011 ( .A1(n1208), .A2(n1336), .ZN(n1335) );
XNOR2_X1 U1012 ( .A(n1337), .B(n1338), .ZN(n1208) );
XOR2_X1 U1013 ( .A(n1339), .B(n1340), .Z(n1338) );
XOR2_X1 U1014 ( .A(G107), .B(n1341), .Z(n1340) );
AND3_X1 U1015 ( .A1(G234), .A2(n1106), .A3(G217), .ZN(n1341) );
XNOR2_X1 U1016 ( .A(G116), .B(n1342), .ZN(n1337) );
XNOR2_X1 U1017 ( .A(G134), .B(n1334), .ZN(n1342) );
INV_X1 U1018 ( .A(G122), .ZN(n1334) );
AND2_X1 U1019 ( .A1(n1270), .A2(n1272), .ZN(n1080) );
NAND2_X1 U1020 ( .A1(n1091), .A2(n1343), .ZN(n1272) );
NAND3_X1 U1021 ( .A1(n1183), .A2(n1311), .A3(G902), .ZN(n1343) );
NOR2_X1 U1022 ( .A1(n1106), .A2(G898), .ZN(n1183) );
NAND3_X1 U1023 ( .A1(n1311), .A2(n1106), .A3(G952), .ZN(n1091) );
NAND2_X1 U1024 ( .A1(G237), .A2(n1344), .ZN(n1311) );
NOR3_X1 U1025 ( .A1(n1096), .A2(n1259), .A3(n1124), .ZN(n1270) );
NAND2_X1 U1026 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U1027 ( .A1(G221), .A2(n1345), .ZN(n1126) );
XNOR2_X1 U1028 ( .A(G469), .B(n1346), .ZN(n1125) );
NOR2_X1 U1029 ( .A1(n1347), .A2(KEYINPUT44), .ZN(n1346) );
INV_X1 U1030 ( .A(n1142), .ZN(n1347) );
NAND2_X1 U1031 ( .A1(n1348), .A2(n1336), .ZN(n1142) );
XOR2_X1 U1032 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1033 ( .A(n1241), .B(KEYINPUT7), .Z(n1350) );
XOR2_X1 U1034 ( .A(n1351), .B(n1169), .Z(n1241) );
XNOR2_X1 U1035 ( .A(n1352), .B(n1339), .ZN(n1169) );
XOR2_X1 U1036 ( .A(G143), .B(G128), .Z(n1339) );
XOR2_X1 U1037 ( .A(n1224), .B(n1188), .Z(n1351) );
NAND2_X1 U1038 ( .A1(n1353), .A2(n1354), .ZN(n1349) );
NAND2_X1 U1039 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1040 ( .A1(n1357), .A2(n1358), .ZN(n1355) );
NAND2_X1 U1041 ( .A1(n1240), .A2(G110), .ZN(n1358) );
NAND2_X1 U1042 ( .A1(n1359), .A2(n1360), .ZN(n1357) );
NAND2_X1 U1043 ( .A1(n1361), .A2(n1362), .ZN(n1353) );
NAND2_X1 U1044 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
NAND2_X1 U1045 ( .A1(n1240), .A2(n1360), .ZN(n1364) );
NAND2_X1 U1046 ( .A1(G110), .A2(n1359), .ZN(n1363) );
XNOR2_X1 U1047 ( .A(n1240), .B(n1365), .ZN(n1359) );
XOR2_X1 U1048 ( .A(KEYINPUT6), .B(KEYINPUT38), .Z(n1365) );
AND2_X1 U1049 ( .A1(n1366), .A2(n1106), .ZN(n1240) );
XNOR2_X1 U1050 ( .A(G227), .B(KEYINPUT26), .ZN(n1366) );
INV_X1 U1051 ( .A(n1356), .ZN(n1361) );
NAND2_X1 U1052 ( .A1(KEYINPUT53), .A2(n1236), .ZN(n1356) );
NAND2_X1 U1053 ( .A1(n1102), .A2(n1103), .ZN(n1259) );
NAND2_X1 U1054 ( .A1(G214), .A2(n1367), .ZN(n1103) );
XOR2_X1 U1055 ( .A(n1145), .B(n1368), .Z(n1102) );
NOR2_X1 U1056 ( .A1(KEYINPUT10), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1057 ( .A(n1146), .B(KEYINPUT56), .Z(n1369) );
NAND2_X1 U1058 ( .A1(G210), .A2(n1367), .ZN(n1146) );
NAND2_X1 U1059 ( .A1(n1370), .A2(n1336), .ZN(n1367) );
INV_X1 U1060 ( .A(G237), .ZN(n1370) );
NAND2_X1 U1061 ( .A1(n1371), .A2(n1336), .ZN(n1145) );
XOR2_X1 U1062 ( .A(n1282), .B(n1372), .Z(n1371) );
XOR2_X1 U1063 ( .A(n1373), .B(n1248), .Z(n1372) );
NAND2_X1 U1064 ( .A1(G224), .A2(n1106), .ZN(n1248) );
NAND2_X1 U1065 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
NAND2_X1 U1066 ( .A1(n1223), .A2(G125), .ZN(n1375) );
XOR2_X1 U1067 ( .A(KEYINPUT46), .B(n1376), .Z(n1374) );
NOR2_X1 U1068 ( .A1(G125), .A2(n1223), .ZN(n1376) );
XNOR2_X1 U1069 ( .A(n1189), .B(n1377), .ZN(n1282) );
NOR2_X1 U1070 ( .A1(n1378), .A2(n1379), .ZN(n1377) );
XOR2_X1 U1071 ( .A(n1380), .B(KEYINPUT60), .Z(n1379) );
NAND2_X1 U1072 ( .A1(n1381), .A2(n1184), .ZN(n1380) );
XOR2_X1 U1073 ( .A(n1188), .B(KEYINPUT40), .Z(n1381) );
NOR2_X1 U1074 ( .A1(n1188), .A2(n1184), .ZN(n1378) );
XNOR2_X1 U1075 ( .A(G113), .B(n1382), .ZN(n1184) );
XOR2_X1 U1076 ( .A(G119), .B(G116), .Z(n1382) );
XNOR2_X1 U1077 ( .A(G101), .B(n1383), .ZN(n1188) );
XOR2_X1 U1078 ( .A(G107), .B(G104), .Z(n1383) );
XNOR2_X1 U1079 ( .A(G122), .B(n1360), .ZN(n1189) );
XNOR2_X1 U1080 ( .A(n1305), .B(KEYINPUT57), .ZN(n1096) );
XOR2_X1 U1081 ( .A(n1384), .B(n1385), .Z(n1305) );
NOR2_X1 U1082 ( .A1(KEYINPUT30), .A2(n1141), .ZN(n1385) );
NAND3_X1 U1083 ( .A1(n1386), .A2(n1336), .A3(n1387), .ZN(n1141) );
NAND3_X1 U1084 ( .A1(n1388), .A2(n1389), .A3(n1227), .ZN(n1387) );
XNOR2_X1 U1085 ( .A(n1390), .B(n1391), .ZN(n1388) );
NAND2_X1 U1086 ( .A1(KEYINPUT18), .A2(n1392), .ZN(n1390) );
NAND2_X1 U1087 ( .A1(n1393), .A2(n1394), .ZN(n1386) );
NAND2_X1 U1088 ( .A1(n1227), .A2(n1389), .ZN(n1394) );
INV_X1 U1089 ( .A(KEYINPUT27), .ZN(n1389) );
AND2_X1 U1090 ( .A1(n1395), .A2(n1396), .ZN(n1227) );
OR2_X1 U1091 ( .A1(n1397), .A2(n1398), .ZN(n1396) );
XOR2_X1 U1092 ( .A(n1399), .B(KEYINPUT12), .Z(n1395) );
NAND2_X1 U1093 ( .A1(n1397), .A2(n1398), .ZN(n1399) );
INV_X1 U1094 ( .A(G113), .ZN(n1398) );
XOR2_X1 U1095 ( .A(G116), .B(n1400), .Z(n1397) );
NOR2_X1 U1096 ( .A1(G119), .A2(KEYINPUT2), .ZN(n1400) );
XNOR2_X1 U1097 ( .A(n1401), .B(n1402), .ZN(n1393) );
INV_X1 U1098 ( .A(n1391), .ZN(n1402) );
XOR2_X1 U1099 ( .A(n1229), .B(KEYINPUT0), .Z(n1391) );
XOR2_X1 U1100 ( .A(n1403), .B(n1307), .Z(n1229) );
INV_X1 U1101 ( .A(G101), .ZN(n1307) );
NAND2_X1 U1102 ( .A1(G210), .A2(n1331), .ZN(n1403) );
NOR2_X1 U1103 ( .A1(G953), .A2(G237), .ZN(n1331) );
NOR2_X1 U1104 ( .A1(n1392), .A2(n1404), .ZN(n1401) );
INV_X1 U1105 ( .A(KEYINPUT18), .ZN(n1404) );
NAND3_X1 U1106 ( .A1(n1405), .A2(n1406), .A3(n1407), .ZN(n1392) );
NAND2_X1 U1107 ( .A1(KEYINPUT29), .A2(n1408), .ZN(n1407) );
OR3_X1 U1108 ( .A1(n1408), .A2(KEYINPUT29), .A3(n1224), .ZN(n1406) );
NAND2_X1 U1109 ( .A1(n1224), .A2(n1409), .ZN(n1405) );
NAND2_X1 U1110 ( .A1(n1410), .A2(n1411), .ZN(n1409) );
INV_X1 U1111 ( .A(KEYINPUT29), .ZN(n1411) );
XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1223), .ZN(n1410) );
INV_X1 U1113 ( .A(n1408), .ZN(n1223) );
XOR2_X1 U1114 ( .A(n1412), .B(n1298), .Z(n1408) );
NAND3_X1 U1115 ( .A1(n1413), .A2(n1414), .A3(KEYINPUT45), .ZN(n1412) );
NAND2_X1 U1116 ( .A1(n1326), .A2(n1415), .ZN(n1414) );
INV_X1 U1117 ( .A(KEYINPUT33), .ZN(n1415) );
XNOR2_X1 U1118 ( .A(G143), .B(G146), .ZN(n1326) );
NAND3_X1 U1119 ( .A1(G143), .A2(n1352), .A3(KEYINPUT33), .ZN(n1413) );
INV_X1 U1120 ( .A(G146), .ZN(n1352) );
XOR2_X1 U1121 ( .A(G137), .B(n1174), .Z(n1224) );
XOR2_X1 U1122 ( .A(G131), .B(G134), .Z(n1174) );
XNOR2_X1 U1123 ( .A(G472), .B(KEYINPUT51), .ZN(n1384) );
INV_X1 U1124 ( .A(n1081), .ZN(n1099) );
XOR2_X1 U1125 ( .A(n1135), .B(KEYINPUT22), .Z(n1081) );
XNOR2_X1 U1126 ( .A(n1197), .B(n1201), .ZN(n1135) );
NAND2_X1 U1127 ( .A1(G217), .A2(n1345), .ZN(n1201) );
NAND2_X1 U1128 ( .A1(n1344), .A2(n1336), .ZN(n1345) );
INV_X1 U1129 ( .A(G902), .ZN(n1336) );
XNOR2_X1 U1130 ( .A(G234), .B(KEYINPUT54), .ZN(n1344) );
NOR2_X1 U1131 ( .A1(n1203), .A2(G902), .ZN(n1197) );
XNOR2_X1 U1132 ( .A(n1416), .B(n1417), .ZN(n1203) );
NOR2_X1 U1133 ( .A1(n1418), .A2(n1419), .ZN(n1417) );
XOR2_X1 U1134 ( .A(n1420), .B(KEYINPUT8), .Z(n1419) );
NAND2_X1 U1135 ( .A1(n1421), .A2(n1422), .ZN(n1420) );
NOR2_X1 U1136 ( .A1(n1421), .A2(n1422), .ZN(n1418) );
XNOR2_X1 U1137 ( .A(n1360), .B(n1423), .ZN(n1422) );
XNOR2_X1 U1138 ( .A(n1298), .B(G119), .ZN(n1423) );
INV_X1 U1139 ( .A(G128), .ZN(n1298) );
INV_X1 U1140 ( .A(G110), .ZN(n1360) );
XNOR2_X1 U1141 ( .A(G146), .B(n1330), .ZN(n1421) );
XNOR2_X1 U1142 ( .A(n1236), .B(G125), .ZN(n1330) );
INV_X1 U1143 ( .A(G140), .ZN(n1236) );
XNOR2_X1 U1144 ( .A(n1424), .B(n1173), .ZN(n1416) );
INV_X1 U1145 ( .A(G137), .ZN(n1173) );
NAND3_X1 U1146 ( .A1(G234), .A2(n1425), .A3(G221), .ZN(n1424) );
XNOR2_X1 U1147 ( .A(KEYINPUT13), .B(n1106), .ZN(n1425) );
INV_X1 U1148 ( .A(G953), .ZN(n1106) );
endmodule


