//Key = 0001010001000111101101101011111100101101001011010111110101101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292;

XNOR2_X1 U703 ( .A(G107), .B(n989), .ZN(G9) );
NOR2_X1 U704 ( .A1(n990), .A2(n991), .ZN(G75) );
NOR3_X1 U705 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
NAND3_X1 U706 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n992) );
NAND2_X1 U707 ( .A1(n998), .A2(n999), .ZN(n997) );
NAND2_X1 U708 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND3_X1 U709 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n1001) );
NAND2_X1 U710 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NAND2_X1 U711 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
OR2_X1 U712 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NAND2_X1 U713 ( .A1(n1011), .A2(n1012), .ZN(n1005) );
NAND2_X1 U714 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND2_X1 U715 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
XOR2_X1 U716 ( .A(KEYINPUT29), .B(n1017), .Z(n1013) );
NAND3_X1 U717 ( .A1(n1007), .A2(n1018), .A3(n1011), .ZN(n1000) );
NAND4_X1 U718 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NAND2_X1 U719 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
XOR2_X1 U720 ( .A(n1002), .B(KEYINPUT1), .Z(n1024) );
NAND3_X1 U721 ( .A1(n1004), .A2(n1025), .A3(n1026), .ZN(n1020) );
NAND2_X1 U722 ( .A1(n1027), .A2(n1028), .ZN(n1019) );
XNOR2_X1 U723 ( .A(n1004), .B(KEYINPUT19), .ZN(n1027) );
INV_X1 U724 ( .A(n1029), .ZN(n998) );
NOR3_X1 U725 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n990) );
INV_X1 U726 ( .A(n995), .ZN(n1030) );
NAND4_X1 U727 ( .A1(n1031), .A2(n1007), .A3(n1032), .A4(n1033), .ZN(n995) );
NOR4_X1 U728 ( .A1(n1034), .A2(n1026), .A3(n1035), .A4(n1036), .ZN(n1033) );
XOR2_X1 U729 ( .A(n1037), .B(n1038), .Z(n1036) );
XNOR2_X1 U730 ( .A(KEYINPUT36), .B(n1039), .ZN(n1037) );
NOR2_X1 U731 ( .A1(KEYINPUT0), .A2(n1040), .ZN(n1039) );
AND2_X1 U732 ( .A1(n1041), .A2(n1042), .ZN(n1035) );
NOR2_X1 U733 ( .A1(n1043), .A2(n1044), .ZN(n1032) );
XOR2_X1 U734 ( .A(n1045), .B(n1046), .Z(n1044) );
XOR2_X1 U735 ( .A(KEYINPUT26), .B(KEYINPUT22), .Z(n1046) );
XNOR2_X1 U736 ( .A(n1047), .B(n1048), .ZN(n1043) );
NOR2_X1 U737 ( .A1(KEYINPUT25), .A2(n1049), .ZN(n1048) );
XOR2_X1 U738 ( .A(n1050), .B(n1051), .Z(G72) );
NOR2_X1 U739 ( .A1(n1052), .A2(n996), .ZN(n1051) );
NOR2_X1 U740 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NOR2_X1 U741 ( .A1(KEYINPUT56), .A2(n1055), .ZN(n1050) );
NOR2_X1 U742 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XOR2_X1 U743 ( .A(n1058), .B(KEYINPUT5), .Z(n1057) );
NAND2_X1 U744 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NOR2_X1 U745 ( .A1(n1059), .A2(n1060), .ZN(n1056) );
NAND2_X1 U746 ( .A1(n994), .A2(n996), .ZN(n1060) );
AND2_X1 U747 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NAND2_X1 U748 ( .A1(n1063), .A2(G953), .ZN(n1062) );
XNOR2_X1 U749 ( .A(G900), .B(KEYINPUT20), .ZN(n1063) );
XOR2_X1 U750 ( .A(n1064), .B(n1065), .Z(n1061) );
XNOR2_X1 U751 ( .A(n1066), .B(n1067), .ZN(n1065) );
XNOR2_X1 U752 ( .A(n1068), .B(n1069), .ZN(n1064) );
XNOR2_X1 U753 ( .A(n1070), .B(n1071), .ZN(n1069) );
INV_X1 U754 ( .A(G125), .ZN(n1071) );
NAND2_X1 U755 ( .A1(KEYINPUT13), .A2(n1072), .ZN(n1070) );
NAND2_X1 U756 ( .A1(n1073), .A2(n1074), .ZN(G69) );
NAND2_X1 U757 ( .A1(n1075), .A2(n996), .ZN(n1074) );
XNOR2_X1 U758 ( .A(n1076), .B(n993), .ZN(n1075) );
NAND2_X1 U759 ( .A1(n1077), .A2(G953), .ZN(n1073) );
NAND2_X1 U760 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U761 ( .A1(n1076), .A2(n1080), .ZN(n1079) );
INV_X1 U762 ( .A(G224), .ZN(n1080) );
NAND2_X1 U763 ( .A1(G224), .A2(n1081), .ZN(n1078) );
NAND2_X1 U764 ( .A1(G898), .A2(n1076), .ZN(n1081) );
NAND2_X1 U765 ( .A1(n1082), .A2(n1083), .ZN(n1076) );
NAND2_X1 U766 ( .A1(G953), .A2(n1084), .ZN(n1083) );
XOR2_X1 U767 ( .A(n1085), .B(n1086), .Z(n1082) );
XNOR2_X1 U768 ( .A(n1087), .B(n1088), .ZN(n1086) );
NAND2_X1 U769 ( .A1(KEYINPUT42), .A2(n1089), .ZN(n1087) );
XOR2_X1 U770 ( .A(G119), .B(n1090), .Z(n1089) );
NOR2_X1 U771 ( .A1(n1091), .A2(n1092), .ZN(G66) );
XOR2_X1 U772 ( .A(n1093), .B(n1094), .Z(n1092) );
NOR2_X1 U773 ( .A1(KEYINPUT43), .A2(n1095), .ZN(n1094) );
XOR2_X1 U774 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U775 ( .A1(n1098), .A2(n1042), .ZN(n1093) );
NOR2_X1 U776 ( .A1(n1091), .A2(n1099), .ZN(G63) );
XOR2_X1 U777 ( .A(n1100), .B(n1101), .Z(n1099) );
AND2_X1 U778 ( .A1(G478), .A2(n1098), .ZN(n1100) );
NOR2_X1 U779 ( .A1(n1091), .A2(n1102), .ZN(G60) );
XNOR2_X1 U780 ( .A(n1103), .B(n1104), .ZN(n1102) );
AND2_X1 U781 ( .A1(G475), .A2(n1098), .ZN(n1104) );
XNOR2_X1 U782 ( .A(G104), .B(n1105), .ZN(G6) );
NOR2_X1 U783 ( .A1(n1091), .A2(n1106), .ZN(G57) );
XOR2_X1 U784 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U785 ( .A(n1109), .B(n1110), .Z(n1108) );
XNOR2_X1 U786 ( .A(n1111), .B(n1112), .ZN(n1110) );
XOR2_X1 U787 ( .A(n1113), .B(n1114), .Z(n1107) );
XOR2_X1 U788 ( .A(n1115), .B(n1116), .Z(n1113) );
NOR2_X1 U789 ( .A1(n1049), .A2(n1117), .ZN(n1116) );
INV_X1 U790 ( .A(G472), .ZN(n1049) );
NAND2_X1 U791 ( .A1(KEYINPUT30), .A2(n1118), .ZN(n1115) );
NOR2_X1 U792 ( .A1(n1091), .A2(n1119), .ZN(G54) );
XOR2_X1 U793 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U794 ( .A1(n1098), .A2(G469), .ZN(n1121) );
INV_X1 U795 ( .A(n1117), .ZN(n1098) );
NAND2_X1 U796 ( .A1(KEYINPUT31), .A2(n1122), .ZN(n1120) );
XNOR2_X1 U797 ( .A(G110), .B(n1123), .ZN(n1122) );
NOR2_X1 U798 ( .A1(n1091), .A2(n1124), .ZN(G51) );
XOR2_X1 U799 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U800 ( .A1(n1127), .A2(n1117), .ZN(n1126) );
NAND2_X1 U801 ( .A1(G902), .A2(n1128), .ZN(n1117) );
OR2_X1 U802 ( .A1(n994), .A2(n993), .ZN(n1128) );
NAND2_X1 U803 ( .A1(n1129), .A2(n1130), .ZN(n993) );
AND4_X1 U804 ( .A1(n1131), .A2(n989), .A3(n1132), .A4(n1133), .ZN(n1130) );
NAND3_X1 U805 ( .A1(n1010), .A2(n1004), .A3(n1134), .ZN(n989) );
AND4_X1 U806 ( .A1(n1135), .A2(n1136), .A3(n1105), .A4(n1137), .ZN(n1129) );
OR2_X1 U807 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND3_X1 U808 ( .A1(n1134), .A2(n1004), .A3(n1009), .ZN(n1105) );
NAND4_X1 U809 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n994) );
NOR4_X1 U810 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
AND2_X1 U811 ( .A1(n1148), .A2(n1149), .ZN(n1142) );
NAND4_X1 U812 ( .A1(n1150), .A2(n1017), .A3(n1009), .A4(n1151), .ZN(n1141) );
NOR2_X1 U813 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U814 ( .A1(n1154), .A2(n1155), .ZN(n1140) );
NAND2_X1 U815 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
NAND2_X1 U816 ( .A1(n1028), .A2(n1158), .ZN(n1157) );
XOR2_X1 U817 ( .A(KEYINPUT54), .B(n1159), .Z(n1158) );
NAND2_X1 U818 ( .A1(n1150), .A2(n1153), .ZN(n1156) );
INV_X1 U819 ( .A(KEYINPUT38), .ZN(n1153) );
NAND2_X1 U820 ( .A1(n1160), .A2(KEYINPUT21), .ZN(n1125) );
XOR2_X1 U821 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U822 ( .A(G125), .B(n1163), .ZN(n1162) );
XOR2_X1 U823 ( .A(n1164), .B(n1165), .Z(n1161) );
NAND2_X1 U824 ( .A1(KEYINPUT34), .A2(n1118), .ZN(n1164) );
NOR2_X1 U825 ( .A1(n996), .A2(G952), .ZN(n1091) );
XNOR2_X1 U826 ( .A(G146), .B(n1166), .ZN(G48) );
NAND3_X1 U827 ( .A1(n1159), .A2(n1028), .A3(n1154), .ZN(n1166) );
XNOR2_X1 U828 ( .A(G143), .B(n1148), .ZN(G45) );
NAND3_X1 U829 ( .A1(n1167), .A2(n1168), .A3(n1169), .ZN(n1148) );
XOR2_X1 U830 ( .A(G140), .B(n1147), .Z(G42) );
AND3_X1 U831 ( .A1(n1023), .A2(n1002), .A3(n1154), .ZN(n1147) );
XNOR2_X1 U832 ( .A(n1146), .B(n1170), .ZN(G39) );
NAND2_X1 U833 ( .A1(KEYINPUT53), .A2(G137), .ZN(n1170) );
AND4_X1 U834 ( .A1(n1011), .A2(n1159), .A3(n1168), .A4(n1002), .ZN(n1146) );
NAND2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(G36) );
NAND2_X1 U836 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
NAND2_X1 U837 ( .A1(G134), .A2(n1175), .ZN(n1171) );
NAND2_X1 U838 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND2_X1 U839 ( .A1(KEYINPUT46), .A2(n1145), .ZN(n1177) );
OR2_X1 U840 ( .A1(n1173), .A2(KEYINPUT46), .ZN(n1176) );
AND2_X1 U841 ( .A1(KEYINPUT60), .A2(n1145), .ZN(n1173) );
AND3_X1 U842 ( .A1(n1168), .A2(n1010), .A3(n1150), .ZN(n1145) );
XNOR2_X1 U843 ( .A(G131), .B(n1178), .ZN(G33) );
NAND2_X1 U844 ( .A1(n1154), .A2(n1150), .ZN(n1178) );
INV_X1 U845 ( .A(n1022), .ZN(n1150) );
NAND2_X1 U846 ( .A1(n1167), .A2(n1002), .ZN(n1022) );
NAND2_X1 U847 ( .A1(n1179), .A2(n1180), .ZN(n1002) );
OR2_X1 U848 ( .A1(n1138), .A2(KEYINPUT58), .ZN(n1180) );
NAND3_X1 U849 ( .A1(n1025), .A2(n1181), .A3(KEYINPUT58), .ZN(n1179) );
AND2_X1 U850 ( .A1(n1009), .A2(n1168), .ZN(n1154) );
XNOR2_X1 U851 ( .A(G128), .B(n1182), .ZN(G30) );
NAND2_X1 U852 ( .A1(KEYINPUT27), .A2(n1144), .ZN(n1182) );
AND4_X1 U853 ( .A1(n1159), .A2(n1168), .A3(n1010), .A4(n1028), .ZN(n1144) );
AND2_X1 U854 ( .A1(n1017), .A2(n1152), .ZN(n1168) );
XOR2_X1 U855 ( .A(n1136), .B(n1183), .Z(G3) );
NAND2_X1 U856 ( .A1(KEYINPUT50), .A2(G101), .ZN(n1183) );
NAND3_X1 U857 ( .A1(n1167), .A2(n1134), .A3(n1011), .ZN(n1136) );
XNOR2_X1 U858 ( .A(G125), .B(n1149), .ZN(G27) );
NAND4_X1 U859 ( .A1(n1023), .A2(n1009), .A3(n1184), .A4(n1007), .ZN(n1149) );
AND2_X1 U860 ( .A1(n1152), .A2(n1028), .ZN(n1184) );
NAND2_X1 U861 ( .A1(n1029), .A2(n1185), .ZN(n1152) );
NAND4_X1 U862 ( .A1(G953), .A2(G902), .A3(n1186), .A4(n1054), .ZN(n1185) );
INV_X1 U863 ( .A(G900), .ZN(n1054) );
XNOR2_X1 U864 ( .A(G122), .B(n1135), .ZN(G24) );
NAND3_X1 U865 ( .A1(n1187), .A2(n1004), .A3(n1169), .ZN(n1135) );
NOR3_X1 U866 ( .A1(n1138), .A2(n1188), .A3(n1189), .ZN(n1169) );
NOR2_X1 U867 ( .A1(n1190), .A2(n1191), .ZN(n1004) );
XOR2_X1 U868 ( .A(G119), .B(n1192), .Z(G21) );
NOR2_X1 U869 ( .A1(n1193), .A2(n1138), .ZN(n1192) );
XOR2_X1 U870 ( .A(n1139), .B(KEYINPUT41), .Z(n1193) );
NAND3_X1 U871 ( .A1(n1011), .A2(n1159), .A3(n1187), .ZN(n1139) );
AND2_X1 U872 ( .A1(n1191), .A2(n1190), .ZN(n1159) );
INV_X1 U873 ( .A(n1194), .ZN(n1190) );
NAND2_X1 U874 ( .A1(n1195), .A2(n1196), .ZN(G18) );
NAND2_X1 U875 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XOR2_X1 U876 ( .A(KEYINPUT45), .B(n1199), .Z(n1195) );
NOR2_X1 U877 ( .A1(n1197), .A2(n1198), .ZN(n1199) );
INV_X1 U878 ( .A(n1131), .ZN(n1197) );
NAND4_X1 U879 ( .A1(n1187), .A2(n1167), .A3(n1010), .A4(n1028), .ZN(n1131) );
NOR2_X1 U880 ( .A1(n1045), .A2(n1188), .ZN(n1010) );
INV_X1 U881 ( .A(n1200), .ZN(n1188) );
XNOR2_X1 U882 ( .A(G113), .B(n1133), .ZN(G15) );
NAND4_X1 U883 ( .A1(n1187), .A2(n1009), .A3(n1167), .A4(n1201), .ZN(n1133) );
AND2_X1 U884 ( .A1(n1194), .A2(n1191), .ZN(n1167) );
NOR2_X1 U885 ( .A1(n1200), .A2(n1189), .ZN(n1009) );
XNOR2_X1 U886 ( .A(n1045), .B(KEYINPUT12), .ZN(n1189) );
AND2_X1 U887 ( .A1(n1007), .A2(n1202), .ZN(n1187) );
NOR2_X1 U888 ( .A1(n1203), .A2(n1015), .ZN(n1007) );
XOR2_X1 U889 ( .A(n1132), .B(n1204), .Z(G12) );
NAND2_X1 U890 ( .A1(KEYINPUT49), .A2(G110), .ZN(n1204) );
NAND3_X1 U891 ( .A1(n1011), .A2(n1134), .A3(n1023), .ZN(n1132) );
NOR2_X1 U892 ( .A1(n1191), .A2(n1194), .ZN(n1023) );
NOR2_X1 U893 ( .A1(n1205), .A2(n1034), .ZN(n1194) );
NOR2_X1 U894 ( .A1(n1041), .A2(n1042), .ZN(n1034) );
AND2_X1 U895 ( .A1(n1206), .A2(n1041), .ZN(n1205) );
NAND2_X1 U896 ( .A1(n1207), .A2(n1208), .ZN(n1041) );
XNOR2_X1 U897 ( .A(n1096), .B(n1097), .ZN(n1207) );
XNOR2_X1 U898 ( .A(n1209), .B(n1210), .ZN(n1097) );
NAND2_X1 U899 ( .A1(n1211), .A2(G221), .ZN(n1209) );
XOR2_X1 U900 ( .A(n1212), .B(n1213), .Z(n1096) );
NOR2_X1 U901 ( .A1(KEYINPUT10), .A2(n1214), .ZN(n1213) );
XOR2_X1 U902 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND2_X1 U903 ( .A1(KEYINPUT9), .A2(n1217), .ZN(n1215) );
XNOR2_X1 U904 ( .A(G128), .B(G137), .ZN(n1212) );
XNOR2_X1 U905 ( .A(n1042), .B(KEYINPUT24), .ZN(n1206) );
AND2_X1 U906 ( .A1(G217), .A2(n1218), .ZN(n1042) );
XNOR2_X1 U907 ( .A(n1047), .B(G472), .ZN(n1191) );
NAND2_X1 U908 ( .A1(n1219), .A2(n1208), .ZN(n1047) );
XOR2_X1 U909 ( .A(n1114), .B(n1220), .Z(n1219) );
XOR2_X1 U910 ( .A(n1221), .B(n1222), .Z(n1220) );
NAND3_X1 U911 ( .A1(n1223), .A2(n1224), .A3(n1225), .ZN(n1222) );
NAND2_X1 U912 ( .A1(KEYINPUT6), .A2(n1112), .ZN(n1225) );
OR3_X1 U913 ( .A1(n1112), .A2(KEYINPUT6), .A3(n1109), .ZN(n1224) );
NAND2_X1 U914 ( .A1(n1226), .A2(n1109), .ZN(n1223) );
NAND3_X1 U915 ( .A1(n1227), .A2(n996), .A3(G210), .ZN(n1109) );
NAND2_X1 U916 ( .A1(n1228), .A2(n1229), .ZN(n1226) );
INV_X1 U917 ( .A(KEYINPUT6), .ZN(n1229) );
XNOR2_X1 U918 ( .A(G101), .B(KEYINPUT3), .ZN(n1228) );
NAND2_X1 U919 ( .A1(KEYINPUT16), .A2(n1230), .ZN(n1221) );
XNOR2_X1 U920 ( .A(n1111), .B(n1118), .ZN(n1230) );
XOR2_X1 U921 ( .A(n1231), .B(n1232), .Z(n1114) );
XNOR2_X1 U922 ( .A(G116), .B(G119), .ZN(n1231) );
AND3_X1 U923 ( .A1(n1201), .A2(n1202), .A3(n1017), .ZN(n1134) );
NOR2_X1 U924 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
AND2_X1 U925 ( .A1(G221), .A2(n1218), .ZN(n1015) );
NAND2_X1 U926 ( .A1(G234), .A2(n1208), .ZN(n1218) );
INV_X1 U927 ( .A(n1203), .ZN(n1016) );
XNOR2_X1 U928 ( .A(n1233), .B(G469), .ZN(n1203) );
NAND2_X1 U929 ( .A1(n1234), .A2(n1208), .ZN(n1233) );
XOR2_X1 U930 ( .A(n1235), .B(n1123), .Z(n1234) );
XOR2_X1 U931 ( .A(n1236), .B(n1237), .Z(n1123) );
XOR2_X1 U932 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U933 ( .A(n1111), .B(n1240), .Z(n1239) );
NOR2_X1 U934 ( .A1(G953), .A2(n1053), .ZN(n1240) );
INV_X1 U935 ( .A(G227), .ZN(n1053) );
NAND3_X1 U936 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1111) );
NAND2_X1 U937 ( .A1(KEYINPUT32), .A2(n1072), .ZN(n1243) );
OR3_X1 U938 ( .A1(n1072), .A2(KEYINPUT32), .A3(n1244), .ZN(n1242) );
NAND2_X1 U939 ( .A1(n1244), .A2(n1245), .ZN(n1241) );
NAND2_X1 U940 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
INV_X1 U941 ( .A(KEYINPUT32), .ZN(n1247) );
XNOR2_X1 U942 ( .A(KEYINPUT7), .B(n1072), .ZN(n1246) );
INV_X1 U943 ( .A(G131), .ZN(n1072) );
XOR2_X1 U944 ( .A(n1248), .B(n1068), .Z(n1244) );
XNOR2_X1 U945 ( .A(G137), .B(n1174), .ZN(n1068) );
XNOR2_X1 U946 ( .A(KEYINPUT17), .B(KEYINPUT11), .ZN(n1248) );
NAND2_X1 U947 ( .A1(KEYINPUT57), .A2(n1112), .ZN(n1238) );
INV_X1 U948 ( .A(G101), .ZN(n1112) );
XOR2_X1 U949 ( .A(n1249), .B(n1250), .Z(n1236) );
XNOR2_X1 U950 ( .A(n1066), .B(n1217), .ZN(n1249) );
INV_X1 U951 ( .A(n1067), .ZN(n1217) );
NAND2_X1 U952 ( .A1(KEYINPUT15), .A2(n1088), .ZN(n1235) );
NAND2_X1 U953 ( .A1(n1029), .A2(n1251), .ZN(n1202) );
NAND4_X1 U954 ( .A1(G953), .A2(G902), .A3(n1186), .A4(n1084), .ZN(n1251) );
INV_X1 U955 ( .A(G898), .ZN(n1084) );
NAND3_X1 U956 ( .A1(n1186), .A2(n996), .A3(G952), .ZN(n1029) );
NAND2_X1 U957 ( .A1(G237), .A2(G234), .ZN(n1186) );
XNOR2_X1 U958 ( .A(n1138), .B(KEYINPUT61), .ZN(n1201) );
INV_X1 U959 ( .A(n1028), .ZN(n1138) );
NOR2_X1 U960 ( .A1(n1025), .A2(n1026), .ZN(n1028) );
INV_X1 U961 ( .A(n1181), .ZN(n1026) );
NAND2_X1 U962 ( .A1(G214), .A2(n1252), .ZN(n1181) );
XNOR2_X1 U963 ( .A(n1031), .B(KEYINPUT63), .ZN(n1025) );
XNOR2_X1 U964 ( .A(n1253), .B(n1127), .ZN(n1031) );
NAND2_X1 U965 ( .A1(G210), .A2(n1252), .ZN(n1127) );
NAND2_X1 U966 ( .A1(n1227), .A2(n1208), .ZN(n1252) );
INV_X1 U967 ( .A(G237), .ZN(n1227) );
NAND2_X1 U968 ( .A1(n1254), .A2(n1208), .ZN(n1253) );
XOR2_X1 U969 ( .A(n1255), .B(n1165), .Z(n1254) );
XNOR2_X1 U970 ( .A(n1256), .B(n1257), .ZN(n1165) );
XOR2_X1 U971 ( .A(KEYINPUT14), .B(n1210), .Z(n1257) );
XNOR2_X1 U972 ( .A(n1088), .B(G119), .ZN(n1210) );
INV_X1 U973 ( .A(G110), .ZN(n1088) );
XOR2_X1 U974 ( .A(n1085), .B(n1090), .Z(n1256) );
XNOR2_X1 U975 ( .A(n1258), .B(n1259), .ZN(n1090) );
NOR2_X1 U976 ( .A1(KEYINPUT40), .A2(n1232), .ZN(n1259) );
XNOR2_X1 U977 ( .A(G113), .B(KEYINPUT62), .ZN(n1232) );
NAND2_X1 U978 ( .A1(KEYINPUT37), .A2(n1198), .ZN(n1258) );
XOR2_X1 U979 ( .A(n1260), .B(n1261), .Z(n1085) );
XNOR2_X1 U980 ( .A(G122), .B(n1262), .ZN(n1261) );
XNOR2_X1 U981 ( .A(KEYINPUT51), .B(KEYINPUT35), .ZN(n1262) );
XNOR2_X1 U982 ( .A(G101), .B(n1250), .ZN(n1260) );
XOR2_X1 U983 ( .A(G104), .B(G107), .Z(n1250) );
NAND2_X1 U984 ( .A1(n1263), .A2(KEYINPUT28), .ZN(n1255) );
XNOR2_X1 U985 ( .A(n1118), .B(n1264), .ZN(n1263) );
XNOR2_X1 U986 ( .A(n1163), .B(n1265), .ZN(n1264) );
NOR2_X1 U987 ( .A1(G125), .A2(KEYINPUT59), .ZN(n1265) );
NAND2_X1 U988 ( .A1(n1266), .A2(n996), .ZN(n1163) );
XNOR2_X1 U989 ( .A(G224), .B(KEYINPUT52), .ZN(n1266) );
XNOR2_X1 U990 ( .A(n1066), .B(KEYINPUT44), .ZN(n1118) );
XNOR2_X1 U991 ( .A(n1267), .B(n1268), .ZN(n1066) );
NOR2_X1 U992 ( .A1(n1200), .A2(n1045), .ZN(n1011) );
XNOR2_X1 U993 ( .A(n1269), .B(G475), .ZN(n1045) );
NAND2_X1 U994 ( .A1(n1103), .A2(n1208), .ZN(n1269) );
INV_X1 U995 ( .A(G902), .ZN(n1208) );
XNOR2_X1 U996 ( .A(n1270), .B(n1271), .ZN(n1103) );
XNOR2_X1 U997 ( .A(n1272), .B(n1273), .ZN(n1271) );
NOR2_X1 U998 ( .A1(KEYINPUT8), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U999 ( .A(n1216), .B(n1067), .ZN(n1274) );
XOR2_X1 U1000 ( .A(G140), .B(KEYINPUT2), .Z(n1067) );
XOR2_X1 U1001 ( .A(G125), .B(n1268), .Z(n1216) );
XOR2_X1 U1002 ( .A(G146), .B(KEYINPUT55), .Z(n1268) );
NAND2_X1 U1003 ( .A1(KEYINPUT39), .A2(n1275), .ZN(n1272) );
XOR2_X1 U1004 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U1005 ( .A(G122), .B(G104), .Z(n1277) );
NOR2_X1 U1006 ( .A1(KEYINPUT23), .A2(n1278), .ZN(n1276) );
INV_X1 U1007 ( .A(G113), .ZN(n1278) );
XNOR2_X1 U1008 ( .A(G131), .B(n1279), .ZN(n1270) );
NOR3_X1 U1009 ( .A1(n1280), .A2(KEYINPUT4), .A3(n1281), .ZN(n1279) );
NOR4_X1 U1010 ( .A1(G953), .A2(G237), .A3(n1282), .A4(n1283), .ZN(n1281) );
XNOR2_X1 U1011 ( .A(n1284), .B(KEYINPUT48), .ZN(n1282) );
NOR2_X1 U1012 ( .A1(n1285), .A2(n1286), .ZN(n1280) );
XNOR2_X1 U1013 ( .A(n1284), .B(KEYINPUT47), .ZN(n1286) );
NOR3_X1 U1014 ( .A1(n1283), .A2(G953), .A3(G237), .ZN(n1285) );
INV_X1 U1015 ( .A(G214), .ZN(n1283) );
XNOR2_X1 U1016 ( .A(n1040), .B(n1038), .ZN(n1200) );
XOR2_X1 U1017 ( .A(G478), .B(KEYINPUT33), .Z(n1038) );
OR2_X1 U1018 ( .A1(n1101), .A2(G902), .ZN(n1040) );
XNOR2_X1 U1019 ( .A(n1287), .B(n1288), .ZN(n1101) );
XNOR2_X1 U1020 ( .A(n1198), .B(n1289), .ZN(n1288) );
XNOR2_X1 U1021 ( .A(n1174), .B(G122), .ZN(n1289) );
INV_X1 U1022 ( .A(G134), .ZN(n1174) );
INV_X1 U1023 ( .A(G116), .ZN(n1198) );
XNOR2_X1 U1024 ( .A(n1290), .B(n1291), .ZN(n1287) );
INV_X1 U1025 ( .A(n1267), .ZN(n1291) );
XOR2_X1 U1026 ( .A(G128), .B(n1284), .Z(n1267) );
XOR2_X1 U1027 ( .A(G143), .B(KEYINPUT18), .Z(n1284) );
XOR2_X1 U1028 ( .A(n1292), .B(G107), .Z(n1290) );
NAND2_X1 U1029 ( .A1(G217), .A2(n1211), .ZN(n1292) );
AND2_X1 U1030 ( .A1(G234), .A2(n996), .ZN(n1211) );
INV_X1 U1031 ( .A(G953), .ZN(n996) );
endmodule


