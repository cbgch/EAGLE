//Key = 0001111010011010111110011000101110000101100010001111100101101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413;

NAND2_X1 U770 ( .A1(n1068), .A2(n1069), .ZN(G9) );
NAND2_X1 U771 ( .A1(G107), .A2(n1070), .ZN(n1069) );
XOR2_X1 U772 ( .A(KEYINPUT4), .B(n1071), .Z(n1068) );
NOR2_X1 U773 ( .A1(G107), .A2(n1070), .ZN(n1071) );
NAND3_X1 U774 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1070) );
NOR2_X1 U775 ( .A1(n1075), .A2(n1076), .ZN(G75) );
NOR4_X1 U776 ( .A1(G953), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1076) );
NOR2_X1 U777 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR2_X1 U778 ( .A1(n1082), .A2(n1083), .ZN(n1080) );
NOR2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
NOR2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U782 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U784 ( .A1(n1094), .A2(n1095), .ZN(n1092) );
NOR2_X1 U785 ( .A1(n1096), .A2(n1097), .ZN(n1094) );
XOR2_X1 U786 ( .A(KEYINPUT43), .B(n1098), .Z(n1097) );
NOR2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1090) );
NOR2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
AND2_X1 U789 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR3_X1 U790 ( .A1(n1093), .A2(n1105), .A3(n1100), .ZN(n1086) );
NOR2_X1 U791 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NOR4_X1 U793 ( .A1(n1110), .A2(n1100), .A3(n1093), .A4(n1089), .ZN(n1082) );
NOR2_X1 U794 ( .A1(n1072), .A2(n1111), .ZN(n1110) );
NOR3_X1 U795 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1075) );
AND4_X1 U796 ( .A1(n1112), .A2(n1096), .A3(n1113), .A4(n1114), .ZN(n1077) );
NOR4_X1 U797 ( .A1(n1115), .A2(n1116), .A3(n1089), .A4(n1117), .ZN(n1114) );
XOR2_X1 U798 ( .A(KEYINPUT33), .B(n1098), .Z(n1117) );
XOR2_X1 U799 ( .A(n1118), .B(G475), .Z(n1115) );
NAND2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U801 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n1119) );
NOR2_X1 U802 ( .A1(n1121), .A2(n1122), .ZN(n1113) );
NOR2_X1 U803 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
AND2_X1 U805 ( .A1(n1127), .A2(KEYINPUT17), .ZN(n1126) );
NOR2_X1 U806 ( .A1(G472), .A2(n1128), .ZN(n1125) );
NOR2_X1 U807 ( .A1(KEYINPUT49), .A2(n1127), .ZN(n1128) );
AND4_X1 U808 ( .A1(n1129), .A2(n1127), .A3(KEYINPUT17), .A4(KEYINPUT49), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1130), .B(n1131), .Z(G72) );
XOR2_X1 U810 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XOR2_X1 U812 ( .A(n1136), .B(n1137), .Z(n1135) );
XNOR2_X1 U813 ( .A(n1138), .B(n1139), .ZN(n1137) );
XOR2_X1 U814 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U815 ( .A1(KEYINPUT53), .A2(n1142), .ZN(n1141) );
NAND2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1140) );
NAND2_X1 U817 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND2_X1 U819 ( .A1(KEYINPUT9), .A2(n1149), .ZN(n1148) );
NAND3_X1 U820 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1143) );
INV_X1 U821 ( .A(KEYINPUT9), .ZN(n1152) );
NAND2_X1 U822 ( .A1(G137), .A2(n1149), .ZN(n1151) );
NAND2_X1 U823 ( .A1(n1153), .A2(n1147), .ZN(n1150) );
INV_X1 U824 ( .A(G137), .ZN(n1147) );
NAND2_X1 U825 ( .A1(n1154), .A2(n1149), .ZN(n1153) );
INV_X1 U826 ( .A(KEYINPUT35), .ZN(n1149) );
XOR2_X1 U827 ( .A(n1155), .B(n1156), .Z(n1136) );
NOR2_X1 U828 ( .A1(KEYINPUT15), .A2(n1157), .ZN(n1156) );
XOR2_X1 U829 ( .A(n1158), .B(G140), .Z(n1157) );
XOR2_X1 U830 ( .A(n1159), .B(KEYINPUT62), .Z(n1155) );
NOR2_X1 U831 ( .A1(KEYINPUT41), .A2(n1160), .ZN(n1132) );
NOR2_X1 U832 ( .A1(n1161), .A2(G953), .ZN(n1160) );
NOR2_X1 U833 ( .A1(n1162), .A2(n1134), .ZN(n1130) );
NOR2_X1 U834 ( .A1(G227), .A2(n1163), .ZN(n1162) );
NAND2_X1 U835 ( .A1(n1164), .A2(n1165), .ZN(G69) );
NAND2_X1 U836 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
NAND2_X1 U837 ( .A1(G953), .A2(n1168), .ZN(n1167) );
NAND2_X1 U838 ( .A1(G898), .A2(G224), .ZN(n1168) );
INV_X1 U839 ( .A(n1169), .ZN(n1166) );
NAND2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1164) );
NAND2_X1 U841 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND2_X1 U842 ( .A1(G953), .A2(n1173), .ZN(n1172) );
XOR2_X1 U843 ( .A(n1174), .B(n1175), .Z(n1169) );
NOR2_X1 U844 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U845 ( .A(n1163), .B(KEYINPUT37), .Z(n1177) );
NOR2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(n1176) );
NAND2_X1 U847 ( .A1(n1180), .A2(n1171), .ZN(n1174) );
INV_X1 U848 ( .A(n1181), .ZN(n1171) );
XOR2_X1 U849 ( .A(n1182), .B(n1183), .Z(n1180) );
NOR2_X1 U850 ( .A1(n1184), .A2(n1185), .ZN(G66) );
XOR2_X1 U851 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XNOR2_X1 U853 ( .A(G217), .B(KEYINPUT36), .ZN(n1188) );
NAND2_X1 U854 ( .A1(KEYINPUT14), .A2(n1190), .ZN(n1186) );
NOR2_X1 U855 ( .A1(n1184), .A2(n1191), .ZN(G63) );
XOR2_X1 U856 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U857 ( .A(KEYINPUT48), .B(n1194), .Z(n1193) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1189), .ZN(n1194) );
INV_X1 U859 ( .A(G478), .ZN(n1195) );
NOR2_X1 U860 ( .A1(n1196), .A2(n1197), .ZN(G60) );
XNOR2_X1 U861 ( .A(n1198), .B(n1199), .ZN(n1197) );
NOR2_X1 U862 ( .A1(n1200), .A2(n1189), .ZN(n1198) );
INV_X1 U863 ( .A(G475), .ZN(n1200) );
XNOR2_X1 U864 ( .A(n1184), .B(KEYINPUT44), .ZN(n1196) );
XOR2_X1 U865 ( .A(G104), .B(n1201), .Z(G6) );
NOR4_X1 U866 ( .A1(KEYINPUT7), .A2(n1093), .A3(n1202), .A4(n1203), .ZN(n1201) );
NOR2_X1 U867 ( .A1(n1184), .A2(n1204), .ZN(G57) );
XOR2_X1 U868 ( .A(n1205), .B(n1206), .Z(n1204) );
XOR2_X1 U869 ( .A(n1207), .B(n1208), .Z(n1206) );
NOR2_X1 U870 ( .A1(n1129), .A2(n1189), .ZN(n1208) );
INV_X1 U871 ( .A(G472), .ZN(n1129) );
NOR2_X1 U872 ( .A1(KEYINPUT42), .A2(n1209), .ZN(n1207) );
XOR2_X1 U873 ( .A(G101), .B(n1210), .Z(n1209) );
NOR2_X1 U874 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U875 ( .A(KEYINPUT47), .B(KEYINPUT21), .Z(n1212) );
NOR2_X1 U876 ( .A1(n1213), .A2(n1214), .ZN(n1205) );
NOR2_X1 U877 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
XNOR2_X1 U878 ( .A(n1217), .B(KEYINPUT54), .ZN(n1216) );
NOR2_X1 U879 ( .A1(n1218), .A2(n1217), .ZN(n1213) );
XNOR2_X1 U880 ( .A(n1219), .B(n1220), .ZN(n1217) );
NOR2_X1 U881 ( .A1(n1184), .A2(n1221), .ZN(G54) );
XOR2_X1 U882 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U883 ( .A1(n1224), .A2(n1189), .ZN(n1223) );
INV_X1 U884 ( .A(G469), .ZN(n1224) );
NOR2_X1 U885 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
XOR2_X1 U886 ( .A(KEYINPUT34), .B(n1227), .Z(n1226) );
NOR2_X1 U887 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
AND2_X1 U888 ( .A1(n1229), .A2(n1228), .ZN(n1225) );
XNOR2_X1 U889 ( .A(n1230), .B(n1231), .ZN(n1229) );
NOR2_X1 U890 ( .A1(KEYINPUT27), .A2(n1232), .ZN(n1231) );
NOR2_X1 U891 ( .A1(n1163), .A2(G952), .ZN(n1184) );
NOR2_X1 U892 ( .A1(n1233), .A2(n1234), .ZN(G51) );
XOR2_X1 U893 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U894 ( .A1(n1237), .A2(n1189), .ZN(n1236) );
NAND2_X1 U895 ( .A1(G902), .A2(n1079), .ZN(n1189) );
NAND3_X1 U896 ( .A1(n1238), .A2(n1161), .A3(n1239), .ZN(n1079) );
XOR2_X1 U897 ( .A(n1178), .B(KEYINPUT55), .Z(n1239) );
NAND4_X1 U898 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1178) );
NAND2_X1 U899 ( .A1(n1095), .A2(n1244), .ZN(n1240) );
XNOR2_X1 U900 ( .A(KEYINPUT45), .B(n1245), .ZN(n1244) );
AND4_X1 U901 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1161) );
NOR4_X1 U902 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1249) );
NOR2_X1 U903 ( .A1(n1254), .A2(n1255), .ZN(n1252) );
NOR2_X1 U904 ( .A1(n1256), .A2(n1257), .ZN(n1254) );
NOR2_X1 U905 ( .A1(n1258), .A2(n1259), .ZN(n1251) );
XOR2_X1 U906 ( .A(KEYINPUT50), .B(n1111), .Z(n1259) );
OR2_X1 U907 ( .A1(n1258), .A2(n1260), .ZN(n1248) );
INV_X1 U908 ( .A(n1179), .ZN(n1238) );
NAND3_X1 U909 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1179) );
NAND2_X1 U910 ( .A1(n1074), .A2(n1264), .ZN(n1263) );
NAND2_X1 U911 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U912 ( .A1(n1267), .A2(n1072), .ZN(n1266) );
XOR2_X1 U913 ( .A(n1093), .B(KEYINPUT40), .Z(n1267) );
INV_X1 U914 ( .A(n1073), .ZN(n1093) );
NAND2_X1 U915 ( .A1(n1111), .A2(n1073), .ZN(n1265) );
NOR2_X1 U916 ( .A1(n1268), .A2(n1269), .ZN(n1235) );
XOR2_X1 U917 ( .A(n1270), .B(KEYINPUT16), .Z(n1269) );
NAND2_X1 U918 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
NOR2_X1 U919 ( .A1(n1272), .A2(n1271), .ZN(n1268) );
XOR2_X1 U920 ( .A(n1218), .B(n1273), .Z(n1271) );
NOR2_X1 U921 ( .A1(G952), .A2(n1274), .ZN(n1233) );
XOR2_X1 U922 ( .A(n1163), .B(KEYINPUT38), .Z(n1274) );
XOR2_X1 U923 ( .A(n1275), .B(n1276), .Z(G48) );
NAND2_X1 U924 ( .A1(n1095), .A2(n1277), .ZN(n1276) );
XOR2_X1 U925 ( .A(KEYINPUT29), .B(n1256), .Z(n1277) );
NOR2_X1 U926 ( .A1(n1203), .A2(n1278), .ZN(n1256) );
XNOR2_X1 U927 ( .A(G143), .B(n1247), .ZN(G45) );
NAND4_X1 U928 ( .A1(n1279), .A2(n1095), .A3(n1102), .A4(n1280), .ZN(n1247) );
AND3_X1 U929 ( .A1(n1107), .A2(n1281), .A3(n1116), .ZN(n1280) );
XOR2_X1 U930 ( .A(n1282), .B(n1283), .Z(G42) );
XOR2_X1 U931 ( .A(n1284), .B(KEYINPUT58), .Z(n1283) );
NAND2_X1 U932 ( .A1(n1285), .A2(n1286), .ZN(n1282) );
NAND4_X1 U933 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1286) );
INV_X1 U934 ( .A(KEYINPUT51), .ZN(n1290) );
NAND2_X1 U935 ( .A1(n1250), .A2(KEYINPUT51), .ZN(n1285) );
AND3_X1 U936 ( .A1(n1107), .A2(n1287), .A3(n1289), .ZN(n1250) );
XOR2_X1 U937 ( .A(G137), .B(n1253), .Z(G39) );
NOR3_X1 U938 ( .A1(n1085), .A2(n1100), .A3(n1278), .ZN(n1253) );
INV_X1 U939 ( .A(n1287), .ZN(n1100) );
XOR2_X1 U940 ( .A(G134), .B(n1291), .Z(G36) );
NOR2_X1 U941 ( .A1(n1260), .A2(n1258), .ZN(n1291) );
XOR2_X1 U942 ( .A(G131), .B(n1292), .Z(G33) );
NOR2_X1 U943 ( .A1(n1203), .A2(n1258), .ZN(n1292) );
NAND4_X1 U944 ( .A1(n1102), .A2(n1107), .A3(n1287), .A4(n1281), .ZN(n1258) );
NAND2_X1 U945 ( .A1(n1293), .A2(n1294), .ZN(n1287) );
NAND3_X1 U946 ( .A1(n1295), .A2(n1096), .A3(n1296), .ZN(n1294) );
INV_X1 U947 ( .A(KEYINPUT43), .ZN(n1296) );
NAND2_X1 U948 ( .A1(KEYINPUT43), .A2(n1095), .ZN(n1293) );
INV_X1 U949 ( .A(n1111), .ZN(n1203) );
NAND2_X1 U950 ( .A1(n1297), .A2(n1298), .ZN(G30) );
NAND2_X1 U951 ( .A1(G128), .A2(n1246), .ZN(n1298) );
XOR2_X1 U952 ( .A(KEYINPUT28), .B(n1299), .Z(n1297) );
NOR2_X1 U953 ( .A1(G128), .A2(n1246), .ZN(n1299) );
OR3_X1 U954 ( .A1(n1260), .A2(n1255), .A3(n1278), .ZN(n1246) );
NAND4_X1 U955 ( .A1(n1107), .A2(n1300), .A3(n1281), .A4(n1103), .ZN(n1278) );
XOR2_X1 U956 ( .A(n1301), .B(n1261), .Z(G3) );
NAND3_X1 U957 ( .A1(n1074), .A2(n1302), .A3(n1102), .ZN(n1261) );
XOR2_X1 U958 ( .A(G125), .B(n1303), .Z(G27) );
NOR2_X1 U959 ( .A1(n1255), .A2(n1304), .ZN(n1303) );
XOR2_X1 U960 ( .A(KEYINPUT60), .B(n1257), .Z(n1304) );
AND2_X1 U961 ( .A1(n1289), .A2(n1305), .ZN(n1257) );
AND4_X1 U962 ( .A1(n1111), .A2(n1104), .A3(n1281), .A4(n1103), .ZN(n1289) );
NAND2_X1 U963 ( .A1(n1081), .A2(n1306), .ZN(n1281) );
NAND3_X1 U964 ( .A1(G902), .A2(n1307), .A3(n1134), .ZN(n1306) );
NOR2_X1 U965 ( .A1(G900), .A2(n1163), .ZN(n1134) );
XNOR2_X1 U966 ( .A(G122), .B(n1241), .ZN(G24) );
NAND4_X1 U967 ( .A1(n1308), .A2(n1073), .A3(n1279), .A4(n1116), .ZN(n1241) );
NOR2_X1 U968 ( .A1(n1103), .A2(n1300), .ZN(n1073) );
XOR2_X1 U969 ( .A(n1309), .B(n1310), .Z(G21) );
XOR2_X1 U970 ( .A(KEYINPUT22), .B(G119), .Z(n1310) );
NOR2_X1 U971 ( .A1(n1255), .A2(n1245), .ZN(n1309) );
NAND4_X1 U972 ( .A1(n1103), .A2(n1311), .A3(n1300), .A4(n1312), .ZN(n1245) );
NOR2_X1 U973 ( .A1(n1085), .A2(n1089), .ZN(n1312) );
INV_X1 U974 ( .A(n1302), .ZN(n1085) );
INV_X1 U975 ( .A(n1313), .ZN(n1300) );
XNOR2_X1 U976 ( .A(G116), .B(n1242), .ZN(G18) );
NAND3_X1 U977 ( .A1(n1102), .A2(n1072), .A3(n1308), .ZN(n1242) );
INV_X1 U978 ( .A(n1260), .ZN(n1072) );
NAND2_X1 U979 ( .A1(n1314), .A2(n1116), .ZN(n1260) );
XOR2_X1 U980 ( .A(KEYINPUT10), .B(n1315), .Z(n1314) );
XNOR2_X1 U981 ( .A(G113), .B(n1243), .ZN(G15) );
NAND3_X1 U982 ( .A1(n1102), .A2(n1111), .A3(n1308), .ZN(n1243) );
AND3_X1 U983 ( .A1(n1095), .A2(n1311), .A3(n1305), .ZN(n1308) );
INV_X1 U984 ( .A(n1089), .ZN(n1305) );
NAND2_X1 U985 ( .A1(n1316), .A2(n1109), .ZN(n1089) );
INV_X1 U986 ( .A(n1108), .ZN(n1316) );
NOR2_X1 U987 ( .A1(n1103), .A2(n1313), .ZN(n1102) );
XOR2_X1 U988 ( .A(n1317), .B(n1262), .Z(G12) );
NAND4_X1 U989 ( .A1(n1074), .A2(n1302), .A3(n1104), .A4(n1103), .ZN(n1262) );
NAND3_X1 U990 ( .A1(n1318), .A2(n1319), .A3(n1112), .ZN(n1103) );
NAND2_X1 U991 ( .A1(G217), .A2(n1320), .ZN(n1112) );
NAND2_X1 U992 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
OR2_X1 U993 ( .A1(n1190), .A2(G234), .ZN(n1321) );
NAND2_X1 U994 ( .A1(n1121), .A2(KEYINPUT57), .ZN(n1319) );
AND3_X1 U995 ( .A1(n1323), .A2(n1322), .A3(n1190), .ZN(n1121) );
NAND2_X1 U996 ( .A1(G217), .A2(n1324), .ZN(n1323) );
NAND2_X1 U997 ( .A1(n1325), .A2(n1326), .ZN(n1318) );
INV_X1 U998 ( .A(KEYINPUT57), .ZN(n1326) );
NAND2_X1 U999 ( .A1(n1190), .A2(n1322), .ZN(n1325) );
XNOR2_X1 U1000 ( .A(n1327), .B(n1328), .ZN(n1190) );
XOR2_X1 U1001 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1002 ( .A(n1331), .B(G110), .Z(n1330) );
NAND2_X1 U1003 ( .A1(KEYINPUT19), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1004 ( .A(n1275), .B(n1333), .Z(n1332) );
NAND3_X1 U1005 ( .A1(n1334), .A2(n1335), .A3(KEYINPUT8), .ZN(n1333) );
NAND3_X1 U1006 ( .A1(n1336), .A2(n1158), .A3(n1337), .ZN(n1335) );
INV_X1 U1007 ( .A(KEYINPUT18), .ZN(n1337) );
XOR2_X1 U1008 ( .A(KEYINPUT11), .B(n1284), .Z(n1336) );
INV_X1 U1009 ( .A(G140), .ZN(n1284) );
NAND2_X1 U1010 ( .A1(n1338), .A2(KEYINPUT18), .ZN(n1334) );
XOR2_X1 U1011 ( .A(G140), .B(n1339), .Z(n1338) );
AND2_X1 U1012 ( .A1(n1158), .A2(KEYINPUT11), .ZN(n1339) );
INV_X1 U1013 ( .A(G146), .ZN(n1275) );
NAND2_X1 U1014 ( .A1(n1340), .A2(G221), .ZN(n1329) );
XNOR2_X1 U1015 ( .A(G119), .B(n1341), .ZN(n1327) );
XOR2_X1 U1016 ( .A(G137), .B(G128), .Z(n1341) );
XNOR2_X1 U1017 ( .A(n1313), .B(KEYINPUT63), .ZN(n1104) );
XOR2_X1 U1018 ( .A(n1127), .B(G472), .Z(n1313) );
NAND2_X1 U1019 ( .A1(n1342), .A2(n1322), .ZN(n1127) );
XOR2_X1 U1020 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1021 ( .A(n1345), .B(n1219), .Z(n1344) );
XNOR2_X1 U1022 ( .A(G116), .B(n1346), .ZN(n1219) );
NAND2_X1 U1023 ( .A1(n1347), .A2(n1348), .ZN(n1345) );
NAND2_X1 U1024 ( .A1(n1218), .A2(n1220), .ZN(n1348) );
XOR2_X1 U1025 ( .A(n1349), .B(KEYINPUT13), .Z(n1347) );
NAND2_X1 U1026 ( .A1(n1230), .A2(n1215), .ZN(n1349) );
INV_X1 U1027 ( .A(n1218), .ZN(n1215) );
XOR2_X1 U1028 ( .A(G101), .B(n1350), .Z(n1343) );
NOR2_X1 U1029 ( .A1(KEYINPUT56), .A2(n1351), .ZN(n1350) );
XNOR2_X1 U1030 ( .A(KEYINPUT31), .B(n1211), .ZN(n1351) );
NAND2_X1 U1031 ( .A1(n1352), .A2(G210), .ZN(n1211) );
NAND2_X1 U1032 ( .A1(n1353), .A2(n1354), .ZN(n1302) );
OR3_X1 U1033 ( .A1(n1279), .A2(n1116), .A3(KEYINPUT10), .ZN(n1354) );
NAND2_X1 U1034 ( .A1(KEYINPUT10), .A2(n1111), .ZN(n1353) );
NOR2_X1 U1035 ( .A1(n1116), .A2(n1315), .ZN(n1111) );
INV_X1 U1036 ( .A(n1279), .ZN(n1315) );
XOR2_X1 U1037 ( .A(n1120), .B(n1355), .Z(n1279) );
XOR2_X1 U1038 ( .A(KEYINPUT6), .B(G475), .Z(n1355) );
NAND2_X1 U1039 ( .A1(n1356), .A2(n1199), .ZN(n1120) );
XOR2_X1 U1040 ( .A(n1357), .B(n1358), .Z(n1199) );
XOR2_X1 U1041 ( .A(n1359), .B(n1360), .Z(n1358) );
XOR2_X1 U1042 ( .A(G131), .B(G125), .Z(n1360) );
XOR2_X1 U1043 ( .A(KEYINPUT24), .B(G140), .Z(n1359) );
XOR2_X1 U1044 ( .A(n1361), .B(n1362), .Z(n1357) );
XOR2_X1 U1045 ( .A(G122), .B(G113), .Z(n1362) );
XOR2_X1 U1046 ( .A(n1363), .B(n1364), .Z(n1361) );
AND2_X1 U1047 ( .A1(G214), .A2(n1352), .ZN(n1364) );
NOR2_X1 U1048 ( .A1(G953), .A2(G237), .ZN(n1352) );
XOR2_X1 U1049 ( .A(n1322), .B(KEYINPUT46), .Z(n1356) );
XNOR2_X1 U1050 ( .A(n1365), .B(G478), .ZN(n1116) );
NAND2_X1 U1051 ( .A1(n1192), .A2(n1322), .ZN(n1365) );
XOR2_X1 U1052 ( .A(n1366), .B(n1367), .Z(n1192) );
XOR2_X1 U1053 ( .A(n1368), .B(n1369), .Z(n1367) );
XOR2_X1 U1054 ( .A(G143), .B(n1159), .Z(n1369) );
INV_X1 U1055 ( .A(G128), .ZN(n1159) );
NAND2_X1 U1056 ( .A1(KEYINPUT39), .A2(n1370), .ZN(n1368) );
XOR2_X1 U1057 ( .A(G107), .B(n1371), .Z(n1370) );
XOR2_X1 U1058 ( .A(G122), .B(G116), .Z(n1371) );
XOR2_X1 U1059 ( .A(n1372), .B(n1373), .Z(n1366) );
NOR2_X1 U1060 ( .A1(n1374), .A2(KEYINPUT25), .ZN(n1373) );
AND2_X1 U1061 ( .A1(n1340), .A2(G217), .ZN(n1374) );
NOR2_X1 U1062 ( .A1(n1324), .A2(G953), .ZN(n1340) );
INV_X1 U1063 ( .A(G234), .ZN(n1324) );
NAND2_X1 U1064 ( .A1(KEYINPUT12), .A2(n1154), .ZN(n1372) );
INV_X1 U1065 ( .A(n1202), .ZN(n1074) );
NAND3_X1 U1066 ( .A1(n1107), .A2(n1311), .A3(n1095), .ZN(n1202) );
INV_X1 U1067 ( .A(n1255), .ZN(n1095) );
NAND2_X1 U1068 ( .A1(n1098), .A2(n1096), .ZN(n1255) );
NAND2_X1 U1069 ( .A1(G214), .A2(n1375), .ZN(n1096) );
INV_X1 U1070 ( .A(n1295), .ZN(n1098) );
XNOR2_X1 U1071 ( .A(n1376), .B(n1237), .ZN(n1295) );
NAND2_X1 U1072 ( .A1(G210), .A2(n1375), .ZN(n1237) );
NAND2_X1 U1073 ( .A1(n1377), .A2(n1322), .ZN(n1375) );
INV_X1 U1074 ( .A(G237), .ZN(n1377) );
NAND2_X1 U1075 ( .A1(n1378), .A2(n1322), .ZN(n1376) );
XNOR2_X1 U1076 ( .A(n1272), .B(n1379), .ZN(n1378) );
XNOR2_X1 U1077 ( .A(n1380), .B(n1273), .ZN(n1379) );
XNOR2_X1 U1078 ( .A(n1158), .B(n1381), .ZN(n1273) );
NOR2_X1 U1079 ( .A1(G953), .A2(n1173), .ZN(n1381) );
INV_X1 U1080 ( .A(G224), .ZN(n1173) );
INV_X1 U1081 ( .A(G125), .ZN(n1158) );
NAND2_X1 U1082 ( .A1(KEYINPUT30), .A2(n1218), .ZN(n1380) );
XOR2_X1 U1083 ( .A(n1382), .B(G128), .Z(n1218) );
NAND2_X1 U1084 ( .A1(n1383), .A2(KEYINPUT23), .ZN(n1382) );
XNOR2_X1 U1085 ( .A(G143), .B(n1384), .ZN(n1383) );
NOR2_X1 U1086 ( .A1(KEYINPUT26), .A2(n1385), .ZN(n1384) );
XOR2_X1 U1087 ( .A(KEYINPUT61), .B(G146), .Z(n1385) );
XOR2_X1 U1088 ( .A(n1386), .B(n1182), .Z(n1272) );
NAND2_X1 U1089 ( .A1(n1387), .A2(n1388), .ZN(n1182) );
NAND2_X1 U1090 ( .A1(G122), .A2(n1317), .ZN(n1388) );
XOR2_X1 U1091 ( .A(KEYINPUT3), .B(n1389), .Z(n1387) );
NOR2_X1 U1092 ( .A1(G122), .A2(n1317), .ZN(n1389) );
NAND2_X1 U1093 ( .A1(n1390), .A2(n1391), .ZN(n1386) );
OR2_X1 U1094 ( .A1(n1183), .A2(KEYINPUT0), .ZN(n1391) );
XNOR2_X1 U1095 ( .A(n1392), .B(n1393), .ZN(n1183) );
NAND3_X1 U1096 ( .A1(n1393), .A2(n1392), .A3(KEYINPUT0), .ZN(n1390) );
XOR2_X1 U1097 ( .A(n1394), .B(n1395), .Z(n1392) );
NOR2_X1 U1098 ( .A1(G104), .A2(KEYINPUT59), .ZN(n1395) );
AND2_X1 U1099 ( .A1(n1396), .A2(n1397), .ZN(n1393) );
OR2_X1 U1100 ( .A1(n1346), .A2(G116), .ZN(n1397) );
NAND2_X1 U1101 ( .A1(G116), .A2(n1398), .ZN(n1396) );
XNOR2_X1 U1102 ( .A(n1346), .B(KEYINPUT20), .ZN(n1398) );
XOR2_X1 U1103 ( .A(G113), .B(G119), .Z(n1346) );
NAND2_X1 U1104 ( .A1(n1081), .A2(n1399), .ZN(n1311) );
NAND3_X1 U1105 ( .A1(n1181), .A2(n1400), .A3(G902), .ZN(n1399) );
XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1307), .ZN(n1400) );
NOR2_X1 U1107 ( .A1(n1163), .A2(G898), .ZN(n1181) );
NAND3_X1 U1108 ( .A1(n1307), .A2(n1163), .A3(G952), .ZN(n1081) );
NAND2_X1 U1109 ( .A1(G237), .A2(G234), .ZN(n1307) );
INV_X1 U1110 ( .A(n1288), .ZN(n1107) );
NAND2_X1 U1111 ( .A1(n1108), .A2(n1109), .ZN(n1288) );
NAND2_X1 U1112 ( .A1(G221), .A2(n1401), .ZN(n1109) );
NAND2_X1 U1113 ( .A1(G234), .A2(n1322), .ZN(n1401) );
XNOR2_X1 U1114 ( .A(n1402), .B(G469), .ZN(n1108) );
NAND2_X1 U1115 ( .A1(n1403), .A2(n1322), .ZN(n1402) );
INV_X1 U1116 ( .A(G902), .ZN(n1322) );
XNOR2_X1 U1117 ( .A(n1232), .B(n1404), .ZN(n1403) );
XOR2_X1 U1118 ( .A(n1405), .B(n1220), .Z(n1404) );
INV_X1 U1119 ( .A(n1230), .ZN(n1220) );
XOR2_X1 U1120 ( .A(n1406), .B(n1145), .Z(n1230) );
INV_X1 U1121 ( .A(n1154), .ZN(n1145) );
XNOR2_X1 U1122 ( .A(G134), .B(KEYINPUT32), .ZN(n1154) );
XOR2_X1 U1123 ( .A(n1142), .B(G137), .Z(n1406) );
INV_X1 U1124 ( .A(G131), .ZN(n1142) );
NOR2_X1 U1125 ( .A1(n1228), .A2(KEYINPUT2), .ZN(n1405) );
AND2_X1 U1126 ( .A1(n1407), .A2(n1408), .ZN(n1228) );
NAND3_X1 U1127 ( .A1(G227), .A2(n1163), .A3(n1409), .ZN(n1408) );
XOR2_X1 U1128 ( .A(n1317), .B(G140), .Z(n1409) );
NAND2_X1 U1129 ( .A1(n1410), .A2(n1411), .ZN(n1407) );
NAND2_X1 U1130 ( .A1(G227), .A2(n1163), .ZN(n1411) );
INV_X1 U1131 ( .A(G953), .ZN(n1163) );
XOR2_X1 U1132 ( .A(G140), .B(G110), .Z(n1410) );
XNOR2_X1 U1133 ( .A(n1412), .B(n1413), .ZN(n1232) );
INV_X1 U1134 ( .A(n1394), .ZN(n1413) );
XOR2_X1 U1135 ( .A(n1301), .B(G107), .Z(n1394) );
INV_X1 U1136 ( .A(G101), .ZN(n1301) );
XOR2_X1 U1137 ( .A(n1363), .B(G128), .Z(n1412) );
XNOR2_X1 U1138 ( .A(G104), .B(n1138), .ZN(n1363) );
XOR2_X1 U1139 ( .A(G143), .B(G146), .Z(n1138) );
INV_X1 U1140 ( .A(G110), .ZN(n1317) );
endmodule


