//Key = 1000001011101000111100011010101000000110101110011110001110000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
n1442, n1443;

XNOR2_X1 U794 ( .A(G107), .B(n1102), .ZN(G9) );
NOR2_X1 U795 ( .A1(n1103), .A2(n1104), .ZN(G75) );
XOR2_X1 U796 ( .A(KEYINPUT60), .B(n1105), .Z(n1104) );
AND3_X1 U797 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1105) );
NOR4_X1 U798 ( .A1(n1109), .A2(n1110), .A3(n1108), .A4(n1111), .ZN(n1103) );
INV_X1 U799 ( .A(G952), .ZN(n1108) );
XOR2_X1 U800 ( .A(KEYINPUT59), .B(n1112), .Z(n1110) );
NOR3_X1 U801 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NAND3_X1 U802 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1113) );
NAND4_X1 U803 ( .A1(n1119), .A2(n1106), .A3(n1120), .A4(n1107), .ZN(n1109) );
NAND4_X1 U804 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
NOR3_X1 U805 ( .A1(n1114), .A2(n1125), .A3(n1126), .ZN(n1124) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
INV_X1 U807 ( .A(n1129), .ZN(n1114) );
OR2_X1 U808 ( .A1(n1130), .A2(n1117), .ZN(n1122) );
OR4_X1 U809 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1121) );
NAND4_X1 U810 ( .A1(n1135), .A2(n1117), .A3(n1136), .A4(n1137), .ZN(n1106) );
NOR4_X1 U811 ( .A1(n1138), .A2(n1134), .A3(n1139), .A4(n1140), .ZN(n1137) );
XNOR2_X1 U812 ( .A(n1141), .B(KEYINPUT57), .ZN(n1140) );
XOR2_X1 U813 ( .A(n1142), .B(n1143), .Z(n1139) );
NOR2_X1 U814 ( .A1(KEYINPUT34), .A2(G478), .ZN(n1143) );
XNOR2_X1 U815 ( .A(n1144), .B(KEYINPUT27), .ZN(n1142) );
XOR2_X1 U816 ( .A(n1145), .B(KEYINPUT40), .Z(n1136) );
NAND2_X1 U817 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND4_X1 U818 ( .A1(n1148), .A2(n1118), .A3(n1117), .A4(n1149), .ZN(n1119) );
NAND2_X1 U819 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND2_X1 U820 ( .A1(n1123), .A2(n1152), .ZN(n1151) );
NAND2_X1 U821 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NAND2_X1 U822 ( .A1(n1138), .A2(n1141), .ZN(n1154) );
NAND2_X1 U823 ( .A1(n1155), .A2(n1129), .ZN(n1150) );
INV_X1 U824 ( .A(n1126), .ZN(n1118) );
XOR2_X1 U825 ( .A(n1156), .B(n1157), .Z(G72) );
XOR2_X1 U826 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U827 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XNOR2_X1 U828 ( .A(G953), .B(KEYINPUT3), .ZN(n1161) );
AND2_X1 U829 ( .A1(G227), .A2(G900), .ZN(n1160) );
NAND2_X1 U830 ( .A1(n1162), .A2(n1163), .ZN(n1158) );
NAND2_X1 U831 ( .A1(G953), .A2(n1164), .ZN(n1163) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1162) );
XOR2_X1 U833 ( .A(n1167), .B(n1168), .Z(n1166) );
NOR2_X1 U834 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U835 ( .A1(n1171), .A2(G140), .ZN(n1170) );
NOR2_X1 U836 ( .A1(KEYINPUT22), .A2(n1172), .ZN(n1171) );
NOR2_X1 U837 ( .A1(KEYINPUT22), .A2(n1173), .ZN(n1169) );
NAND2_X1 U838 ( .A1(n1174), .A2(n1175), .ZN(n1167) );
NAND2_X1 U839 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U840 ( .A(KEYINPUT44), .B(n1178), .Z(n1174) );
NOR2_X1 U841 ( .A1(n1177), .A2(n1176), .ZN(n1178) );
XNOR2_X1 U842 ( .A(KEYINPUT62), .B(n1179), .ZN(n1176) );
XNOR2_X1 U843 ( .A(n1180), .B(G131), .ZN(n1165) );
NAND2_X1 U844 ( .A1(n1107), .A2(n1181), .ZN(n1156) );
NAND2_X1 U845 ( .A1(n1182), .A2(n1183), .ZN(G69) );
NAND2_X1 U846 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
INV_X1 U847 ( .A(n1186), .ZN(n1185) );
NAND2_X1 U848 ( .A1(n1187), .A2(n1188), .ZN(n1184) );
INV_X1 U849 ( .A(n1189), .ZN(n1188) );
NAND2_X1 U850 ( .A1(n1186), .A2(n1187), .ZN(n1182) );
AND2_X1 U851 ( .A1(n1190), .A2(n1191), .ZN(n1187) );
OR2_X1 U852 ( .A1(n1107), .A2(G224), .ZN(n1191) );
NAND2_X1 U853 ( .A1(n1192), .A2(n1107), .ZN(n1190) );
NOR4_X1 U854 ( .A1(n1193), .A2(n1194), .A3(KEYINPUT2), .A4(n1189), .ZN(n1186) );
XOR2_X1 U855 ( .A(KEYINPUT7), .B(n1195), .Z(n1194) );
NOR2_X1 U856 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
AND2_X1 U857 ( .A1(n1197), .A2(n1196), .ZN(n1193) );
NOR2_X1 U858 ( .A1(n1198), .A2(n1199), .ZN(G66) );
XOR2_X1 U859 ( .A(n1200), .B(n1201), .Z(n1199) );
NAND2_X1 U860 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
XOR2_X1 U861 ( .A(KEYINPUT61), .B(G217), .Z(n1203) );
NOR2_X1 U862 ( .A1(n1198), .A2(n1204), .ZN(G63) );
NOR3_X1 U863 ( .A1(n1144), .A2(n1205), .A3(n1206), .ZN(n1204) );
AND3_X1 U864 ( .A1(n1207), .A2(G478), .A3(n1202), .ZN(n1206) );
NOR2_X1 U865 ( .A1(n1208), .A2(n1207), .ZN(n1205) );
AND2_X1 U866 ( .A1(n1111), .A2(G478), .ZN(n1208) );
INV_X1 U867 ( .A(n1209), .ZN(n1111) );
NOR2_X1 U868 ( .A1(n1198), .A2(n1210), .ZN(G60) );
XNOR2_X1 U869 ( .A(n1211), .B(n1212), .ZN(n1210) );
NAND2_X1 U870 ( .A1(KEYINPUT24), .A2(n1213), .ZN(n1211) );
NAND2_X1 U871 ( .A1(n1202), .A2(G475), .ZN(n1213) );
XNOR2_X1 U872 ( .A(G104), .B(n1214), .ZN(G6) );
NOR2_X1 U873 ( .A1(n1198), .A2(n1215), .ZN(G57) );
XOR2_X1 U874 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U875 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U876 ( .A(n1220), .B(n1221), .Z(n1216) );
XOR2_X1 U877 ( .A(n1222), .B(n1223), .Z(n1221) );
NAND2_X1 U878 ( .A1(KEYINPUT8), .A2(n1224), .ZN(n1223) );
NAND2_X1 U879 ( .A1(n1202), .A2(G472), .ZN(n1224) );
NAND2_X1 U880 ( .A1(KEYINPUT17), .A2(n1225), .ZN(n1220) );
NOR2_X1 U881 ( .A1(n1198), .A2(n1226), .ZN(G54) );
NOR3_X1 U882 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1226) );
NOR2_X1 U883 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NOR2_X1 U884 ( .A1(n1232), .A2(n1233), .ZN(n1230) );
XOR2_X1 U885 ( .A(n1234), .B(KEYINPUT58), .Z(n1232) );
NOR3_X1 U886 ( .A1(n1235), .A2(n1234), .A3(n1233), .ZN(n1228) );
INV_X1 U887 ( .A(n1231), .ZN(n1235) );
XNOR2_X1 U888 ( .A(n1236), .B(n1237), .ZN(n1231) );
XNOR2_X1 U889 ( .A(n1238), .B(n1239), .ZN(n1236) );
NAND2_X1 U890 ( .A1(KEYINPUT9), .A2(n1180), .ZN(n1239) );
NAND2_X1 U891 ( .A1(KEYINPUT47), .A2(n1240), .ZN(n1238) );
AND2_X1 U892 ( .A1(n1233), .A2(n1234), .ZN(n1227) );
NAND2_X1 U893 ( .A1(n1202), .A2(G469), .ZN(n1234) );
INV_X1 U894 ( .A(KEYINPUT54), .ZN(n1233) );
NOR2_X1 U895 ( .A1(n1198), .A2(n1241), .ZN(G51) );
XOR2_X1 U896 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR3_X1 U897 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1243) );
AND2_X1 U898 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NOR3_X1 U899 ( .A1(n1248), .A2(KEYINPUT29), .A3(n1247), .ZN(n1245) );
OR2_X1 U900 ( .A1(KEYINPUT52), .A2(n1249), .ZN(n1247) );
NOR2_X1 U901 ( .A1(n1250), .A2(n1251), .ZN(n1248) );
AND2_X1 U902 ( .A1(n1252), .A2(n1253), .ZN(n1250) );
AND2_X1 U903 ( .A1(n1249), .A2(KEYINPUT29), .ZN(n1244) );
INV_X1 U904 ( .A(n1254), .ZN(n1249) );
NAND2_X1 U905 ( .A1(n1202), .A2(n1255), .ZN(n1242) );
NOR2_X1 U906 ( .A1(n1256), .A2(n1209), .ZN(n1202) );
NOR2_X1 U907 ( .A1(n1181), .A2(n1192), .ZN(n1209) );
NAND4_X1 U908 ( .A1(n1257), .A2(n1214), .A3(n1258), .A4(n1259), .ZN(n1192) );
AND3_X1 U909 ( .A1(n1260), .A2(n1102), .A3(n1261), .ZN(n1259) );
NAND3_X1 U910 ( .A1(n1116), .A2(n1117), .A3(n1262), .ZN(n1102) );
NAND2_X1 U911 ( .A1(n1131), .A2(n1263), .ZN(n1258) );
NAND3_X1 U912 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1263) );
XOR2_X1 U913 ( .A(n1267), .B(KEYINPUT39), .Z(n1266) );
NAND3_X1 U914 ( .A1(n1268), .A2(n1123), .A3(n1269), .ZN(n1264) );
NAND3_X1 U915 ( .A1(n1262), .A2(n1117), .A3(n1155), .ZN(n1214) );
NAND3_X1 U916 ( .A1(n1123), .A2(n1262), .A3(n1133), .ZN(n1257) );
NAND4_X1 U917 ( .A1(n1270), .A2(n1271), .A3(n1272), .A4(n1273), .ZN(n1181) );
AND4_X1 U918 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1273) );
NOR3_X1 U919 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1272) );
NOR2_X1 U920 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
NAND4_X1 U921 ( .A1(n1116), .A2(n1283), .A3(n1284), .A4(n1285), .ZN(n1282) );
INV_X1 U922 ( .A(KEYINPUT11), .ZN(n1281) );
NOR2_X1 U923 ( .A1(KEYINPUT11), .A2(n1286), .ZN(n1279) );
NOR3_X1 U924 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1278) );
NOR2_X1 U925 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
INV_X1 U926 ( .A(KEYINPUT4), .ZN(n1291) );
NOR3_X1 U927 ( .A1(n1115), .A2(n1292), .A3(n1293), .ZN(n1290) );
NOR2_X1 U928 ( .A1(KEYINPUT4), .A2(n1294), .ZN(n1288) );
NOR2_X1 U929 ( .A1(n1107), .A2(G952), .ZN(n1198) );
XNOR2_X1 U930 ( .A(G146), .B(n1274), .ZN(G48) );
NAND4_X1 U931 ( .A1(n1155), .A2(n1268), .A3(n1283), .A4(n1284), .ZN(n1274) );
XNOR2_X1 U932 ( .A(G143), .B(n1270), .ZN(G45) );
NAND4_X1 U933 ( .A1(n1295), .A2(n1296), .A3(n1284), .A4(n1297), .ZN(n1270) );
NAND2_X1 U934 ( .A1(n1298), .A2(n1299), .ZN(G42) );
NAND4_X1 U935 ( .A1(n1294), .A2(n1300), .A3(n1301), .A4(n1302), .ZN(n1299) );
NAND2_X1 U936 ( .A1(KEYINPUT16), .A2(G140), .ZN(n1302) );
OR2_X1 U937 ( .A1(G140), .A2(KEYINPUT37), .ZN(n1301) );
NAND3_X1 U938 ( .A1(G140), .A2(n1303), .A3(KEYINPUT16), .ZN(n1298) );
NAND3_X1 U939 ( .A1(n1294), .A2(n1300), .A3(KEYINPUT37), .ZN(n1303) );
XNOR2_X1 U940 ( .A(G137), .B(n1271), .ZN(G39) );
NAND3_X1 U941 ( .A1(n1268), .A2(n1123), .A3(n1294), .ZN(n1271) );
XNOR2_X1 U942 ( .A(G134), .B(n1277), .ZN(G36) );
NAND3_X1 U943 ( .A1(n1294), .A2(n1116), .A3(n1133), .ZN(n1277) );
XNOR2_X1 U944 ( .A(G131), .B(n1276), .ZN(G33) );
NAND3_X1 U945 ( .A1(n1294), .A2(n1155), .A3(n1133), .ZN(n1276) );
NOR3_X1 U946 ( .A1(n1153), .A2(n1293), .A3(n1115), .ZN(n1294) );
INV_X1 U947 ( .A(n1148), .ZN(n1115) );
NOR2_X1 U948 ( .A1(n1304), .A2(n1134), .ZN(n1148) );
INV_X1 U949 ( .A(n1284), .ZN(n1293) );
XNOR2_X1 U950 ( .A(G128), .B(n1286), .ZN(G30) );
NAND4_X1 U951 ( .A1(n1268), .A2(n1116), .A3(n1283), .A4(n1284), .ZN(n1286) );
XNOR2_X1 U952 ( .A(G101), .B(n1305), .ZN(G3) );
NAND4_X1 U953 ( .A1(KEYINPUT38), .A2(n1295), .A3(n1123), .A4(n1306), .ZN(n1305) );
XNOR2_X1 U954 ( .A(KEYINPUT28), .B(n1307), .ZN(n1306) );
AND2_X1 U955 ( .A1(n1133), .A2(n1283), .ZN(n1295) );
XOR2_X1 U956 ( .A(n1275), .B(n1308), .Z(G27) );
NOR2_X1 U957 ( .A1(G125), .A2(KEYINPUT20), .ZN(n1308) );
NAND4_X1 U958 ( .A1(n1300), .A2(n1129), .A3(n1131), .A4(n1284), .ZN(n1275) );
NAND2_X1 U959 ( .A1(n1126), .A2(n1309), .ZN(n1284) );
NAND4_X1 U960 ( .A1(G953), .A2(G902), .A3(n1310), .A4(n1164), .ZN(n1309) );
INV_X1 U961 ( .A(G900), .ZN(n1164) );
INV_X1 U962 ( .A(n1287), .ZN(n1300) );
NAND2_X1 U963 ( .A1(n1132), .A2(n1155), .ZN(n1287) );
XOR2_X1 U964 ( .A(n1260), .B(n1311), .Z(G24) );
XNOR2_X1 U965 ( .A(G122), .B(KEYINPUT33), .ZN(n1311) );
NAND4_X1 U966 ( .A1(n1269), .A2(n1127), .A3(n1296), .A4(n1297), .ZN(n1260) );
AND2_X1 U967 ( .A1(n1117), .A2(n1131), .ZN(n1127) );
NOR2_X1 U968 ( .A1(n1312), .A2(n1313), .ZN(n1117) );
XNOR2_X1 U969 ( .A(G119), .B(n1314), .ZN(G21) );
NAND4_X1 U970 ( .A1(n1315), .A2(n1269), .A3(n1268), .A4(n1123), .ZN(n1314) );
INV_X1 U971 ( .A(n1285), .ZN(n1268) );
NAND2_X1 U972 ( .A1(n1313), .A2(n1312), .ZN(n1285) );
XNOR2_X1 U973 ( .A(n1131), .B(KEYINPUT10), .ZN(n1315) );
XNOR2_X1 U974 ( .A(G116), .B(n1316), .ZN(G18) );
NAND2_X1 U975 ( .A1(n1317), .A2(n1131), .ZN(n1316) );
XOR2_X1 U976 ( .A(n1265), .B(KEYINPUT56), .Z(n1317) );
NAND3_X1 U977 ( .A1(n1133), .A2(n1116), .A3(n1269), .ZN(n1265) );
AND2_X1 U978 ( .A1(n1318), .A2(n1296), .ZN(n1116) );
XNOR2_X1 U979 ( .A(n1319), .B(n1320), .ZN(G15) );
NOR2_X1 U980 ( .A1(n1321), .A2(n1267), .ZN(n1320) );
NAND3_X1 U981 ( .A1(n1133), .A2(n1155), .A3(n1269), .ZN(n1267) );
AND2_X1 U982 ( .A1(n1129), .A2(n1307), .ZN(n1269) );
NOR2_X1 U983 ( .A1(n1322), .A2(n1138), .ZN(n1129) );
INV_X1 U984 ( .A(n1141), .ZN(n1322) );
NOR2_X1 U985 ( .A1(n1323), .A2(n1318), .ZN(n1155) );
AND2_X1 U986 ( .A1(n1324), .A2(n1312), .ZN(n1133) );
XNOR2_X1 U987 ( .A(G110), .B(n1261), .ZN(G12) );
NAND3_X1 U988 ( .A1(n1123), .A2(n1262), .A3(n1132), .ZN(n1261) );
NOR2_X1 U989 ( .A1(n1312), .A2(n1324), .ZN(n1132) );
INV_X1 U990 ( .A(n1313), .ZN(n1324) );
XNOR2_X1 U991 ( .A(n1325), .B(n1326), .ZN(n1313) );
AND2_X1 U992 ( .A1(n1327), .A2(G217), .ZN(n1326) );
NAND2_X1 U993 ( .A1(n1201), .A2(n1256), .ZN(n1325) );
XOR2_X1 U994 ( .A(n1328), .B(n1329), .Z(n1201) );
XOR2_X1 U995 ( .A(G128), .B(n1330), .Z(n1329) );
XNOR2_X1 U996 ( .A(KEYINPUT1), .B(n1331), .ZN(n1330) );
XOR2_X1 U997 ( .A(n1332), .B(n1333), .Z(n1328) );
XNOR2_X1 U998 ( .A(G110), .B(n1334), .ZN(n1333) );
NAND3_X1 U999 ( .A1(n1335), .A2(n1336), .A3(n1337), .ZN(n1334) );
OR2_X1 U1000 ( .A1(n1338), .A2(n1173), .ZN(n1337) );
NAND3_X1 U1001 ( .A1(n1338), .A2(n1172), .A3(G140), .ZN(n1336) );
NAND2_X1 U1002 ( .A1(n1339), .A2(n1240), .ZN(n1335) );
XNOR2_X1 U1003 ( .A(n1340), .B(n1338), .ZN(n1339) );
XOR2_X1 U1004 ( .A(n1341), .B(n1177), .Z(n1338) );
INV_X1 U1005 ( .A(G137), .ZN(n1177) );
NAND2_X1 U1006 ( .A1(KEYINPUT6), .A2(n1342), .ZN(n1341) );
NAND3_X1 U1007 ( .A1(G234), .A2(n1107), .A3(G221), .ZN(n1342) );
NAND2_X1 U1008 ( .A1(KEYINPUT0), .A2(G119), .ZN(n1332) );
XNOR2_X1 U1009 ( .A(n1343), .B(G472), .ZN(n1312) );
NAND2_X1 U1010 ( .A1(n1344), .A2(n1256), .ZN(n1343) );
XOR2_X1 U1011 ( .A(n1345), .B(n1218), .Z(n1344) );
XOR2_X1 U1012 ( .A(n1346), .B(G101), .Z(n1218) );
NAND2_X1 U1013 ( .A1(n1347), .A2(G210), .ZN(n1346) );
NAND3_X1 U1014 ( .A1(n1348), .A2(n1349), .A3(n1350), .ZN(n1345) );
NAND2_X1 U1015 ( .A1(n1351), .A2(n1352), .ZN(n1350) );
OR3_X1 U1016 ( .A1(n1352), .A2(n1351), .A3(n1222), .ZN(n1349) );
INV_X1 U1017 ( .A(KEYINPUT19), .ZN(n1352) );
NAND2_X1 U1018 ( .A1(n1353), .A2(n1222), .ZN(n1348) );
NAND3_X1 U1019 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1222) );
INV_X1 U1020 ( .A(n1357), .ZN(n1356) );
NAND2_X1 U1021 ( .A1(n1358), .A2(n1359), .ZN(n1355) );
INV_X1 U1022 ( .A(KEYINPUT51), .ZN(n1359) );
NAND2_X1 U1023 ( .A1(n1360), .A2(KEYINPUT51), .ZN(n1354) );
XNOR2_X1 U1024 ( .A(n1319), .B(n1361), .ZN(n1360) );
NOR2_X1 U1025 ( .A1(G116), .A2(n1362), .ZN(n1361) );
NAND2_X1 U1026 ( .A1(n1363), .A2(KEYINPUT19), .ZN(n1353) );
XNOR2_X1 U1027 ( .A(n1351), .B(KEYINPUT46), .ZN(n1363) );
XNOR2_X1 U1028 ( .A(n1225), .B(n1219), .ZN(n1351) );
AND2_X1 U1029 ( .A1(n1283), .A2(n1307), .ZN(n1262) );
NAND2_X1 U1030 ( .A1(n1126), .A2(n1364), .ZN(n1307) );
NAND3_X1 U1031 ( .A1(G902), .A2(n1310), .A3(n1189), .ZN(n1364) );
NOR2_X1 U1032 ( .A1(G898), .A2(n1107), .ZN(n1189) );
NAND3_X1 U1033 ( .A1(n1310), .A2(n1107), .A3(G952), .ZN(n1126) );
NAND2_X1 U1034 ( .A1(G237), .A2(n1365), .ZN(n1310) );
NOR2_X1 U1035 ( .A1(n1321), .A2(n1153), .ZN(n1283) );
INV_X1 U1036 ( .A(n1292), .ZN(n1153) );
NOR2_X1 U1037 ( .A1(n1141), .A2(n1138), .ZN(n1292) );
AND2_X1 U1038 ( .A1(G221), .A2(n1327), .ZN(n1138) );
NAND2_X1 U1039 ( .A1(n1366), .A2(n1256), .ZN(n1327) );
XOR2_X1 U1040 ( .A(KEYINPUT5), .B(n1365), .Z(n1366) );
XOR2_X1 U1041 ( .A(G234), .B(KEYINPUT21), .Z(n1365) );
XNOR2_X1 U1042 ( .A(n1367), .B(n1368), .ZN(n1141) );
XOR2_X1 U1043 ( .A(KEYINPUT43), .B(G469), .Z(n1368) );
NAND2_X1 U1044 ( .A1(n1369), .A2(n1256), .ZN(n1367) );
XNOR2_X1 U1045 ( .A(n1237), .B(n1370), .ZN(n1369) );
XNOR2_X1 U1046 ( .A(n1180), .B(G140), .ZN(n1370) );
AND2_X1 U1047 ( .A1(n1371), .A2(n1372), .ZN(n1180) );
NAND2_X1 U1048 ( .A1(G128), .A2(n1373), .ZN(n1372) );
XOR2_X1 U1049 ( .A(KEYINPUT55), .B(n1374), .Z(n1371) );
NOR2_X1 U1050 ( .A1(G128), .A2(n1373), .ZN(n1374) );
XNOR2_X1 U1051 ( .A(n1331), .B(n1375), .ZN(n1373) );
NOR2_X1 U1052 ( .A1(KEYINPUT32), .A2(n1376), .ZN(n1375) );
XNOR2_X1 U1053 ( .A(n1377), .B(n1378), .ZN(n1237) );
XOR2_X1 U1054 ( .A(n1219), .B(n1379), .Z(n1378) );
XNOR2_X1 U1055 ( .A(n1380), .B(n1381), .ZN(n1219) );
NOR2_X1 U1056 ( .A1(KEYINPUT45), .A2(G134), .ZN(n1381) );
XNOR2_X1 U1057 ( .A(G131), .B(G137), .ZN(n1380) );
XOR2_X1 U1058 ( .A(n1382), .B(n1383), .Z(n1377) );
XNOR2_X1 U1059 ( .A(KEYINPUT18), .B(n1384), .ZN(n1383) );
INV_X1 U1060 ( .A(G110), .ZN(n1384) );
NAND2_X1 U1061 ( .A1(G227), .A2(n1107), .ZN(n1382) );
INV_X1 U1062 ( .A(n1131), .ZN(n1321) );
NOR2_X1 U1063 ( .A1(n1128), .A2(n1134), .ZN(n1131) );
INV_X1 U1064 ( .A(n1130), .ZN(n1134) );
NAND2_X1 U1065 ( .A1(G214), .A2(n1385), .ZN(n1130) );
INV_X1 U1066 ( .A(n1304), .ZN(n1128) );
XNOR2_X1 U1067 ( .A(n1135), .B(KEYINPUT36), .ZN(n1304) );
XOR2_X1 U1068 ( .A(n1386), .B(n1255), .Z(n1135) );
AND2_X1 U1069 ( .A1(G210), .A2(n1385), .ZN(n1255) );
NAND2_X1 U1070 ( .A1(n1387), .A2(n1256), .ZN(n1385) );
INV_X1 U1071 ( .A(G237), .ZN(n1387) );
NAND2_X1 U1072 ( .A1(n1388), .A2(n1389), .ZN(n1386) );
XOR2_X1 U1073 ( .A(n1390), .B(n1391), .Z(n1389) );
NOR3_X1 U1074 ( .A1(n1251), .A2(n1392), .A3(n1393), .ZN(n1391) );
NOR2_X1 U1075 ( .A1(KEYINPUT63), .A2(n1253), .ZN(n1393) );
AND3_X1 U1076 ( .A1(n1253), .A2(n1252), .A3(KEYINPUT63), .ZN(n1392) );
NOR2_X1 U1077 ( .A1(n1253), .A2(n1252), .ZN(n1251) );
XOR2_X1 U1078 ( .A(n1225), .B(n1172), .Z(n1252) );
XNOR2_X1 U1079 ( .A(G146), .B(n1394), .ZN(n1225) );
NAND2_X1 U1080 ( .A1(G224), .A2(n1107), .ZN(n1253) );
NAND2_X1 U1081 ( .A1(KEYINPUT49), .A2(n1254), .ZN(n1390) );
XNOR2_X1 U1082 ( .A(n1197), .B(n1196), .ZN(n1254) );
XNOR2_X1 U1083 ( .A(n1379), .B(n1395), .ZN(n1196) );
NOR2_X1 U1084 ( .A1(n1357), .A2(n1358), .ZN(n1395) );
NAND2_X1 U1085 ( .A1(n1396), .A2(n1397), .ZN(n1358) );
NAND3_X1 U1086 ( .A1(n1319), .A2(n1398), .A3(n1362), .ZN(n1397) );
INV_X1 U1087 ( .A(G119), .ZN(n1362) );
NAND2_X1 U1088 ( .A1(n1399), .A2(G119), .ZN(n1396) );
XNOR2_X1 U1089 ( .A(n1398), .B(G113), .ZN(n1399) );
NOR3_X1 U1090 ( .A1(n1319), .A2(G119), .A3(n1398), .ZN(n1357) );
XNOR2_X1 U1091 ( .A(n1400), .B(n1401), .ZN(n1379) );
XNOR2_X1 U1092 ( .A(G101), .B(G104), .ZN(n1400) );
XNOR2_X1 U1093 ( .A(G110), .B(n1402), .ZN(n1197) );
XNOR2_X1 U1094 ( .A(G902), .B(KEYINPUT14), .ZN(n1388) );
AND2_X1 U1095 ( .A1(n1318), .A2(n1403), .ZN(n1123) );
XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1323), .Z(n1403) );
XOR2_X1 U1097 ( .A(n1296), .B(KEYINPUT53), .Z(n1323) );
XOR2_X1 U1098 ( .A(n1144), .B(G478), .Z(n1296) );
NOR2_X1 U1099 ( .A1(n1207), .A2(G902), .ZN(n1144) );
XNOR2_X1 U1100 ( .A(n1404), .B(n1405), .ZN(n1207) );
AND3_X1 U1101 ( .A1(G217), .A2(n1107), .A3(G234), .ZN(n1405) );
INV_X1 U1102 ( .A(G953), .ZN(n1107) );
NAND2_X1 U1103 ( .A1(n1406), .A2(n1407), .ZN(n1404) );
NAND2_X1 U1104 ( .A1(n1408), .A2(n1409), .ZN(n1407) );
XOR2_X1 U1105 ( .A(KEYINPUT42), .B(n1410), .Z(n1406) );
NOR2_X1 U1106 ( .A1(n1408), .A2(n1409), .ZN(n1410) );
XNOR2_X1 U1107 ( .A(n1411), .B(n1401), .ZN(n1409) );
XOR2_X1 U1108 ( .A(G107), .B(KEYINPUT13), .Z(n1401) );
NAND2_X1 U1109 ( .A1(n1412), .A2(n1413), .ZN(n1411) );
NAND2_X1 U1110 ( .A1(G116), .A2(n1402), .ZN(n1413) );
INV_X1 U1111 ( .A(G122), .ZN(n1402) );
XOR2_X1 U1112 ( .A(n1414), .B(KEYINPUT15), .Z(n1412) );
NAND2_X1 U1113 ( .A1(G122), .A2(n1398), .ZN(n1414) );
INV_X1 U1114 ( .A(G116), .ZN(n1398) );
XOR2_X1 U1115 ( .A(n1415), .B(n1394), .Z(n1408) );
XNOR2_X1 U1116 ( .A(G128), .B(n1376), .ZN(n1394) );
INV_X1 U1117 ( .A(G143), .ZN(n1376) );
NAND2_X1 U1118 ( .A1(KEYINPUT30), .A2(n1179), .ZN(n1415) );
INV_X1 U1119 ( .A(G134), .ZN(n1179) );
INV_X1 U1120 ( .A(n1297), .ZN(n1318) );
NAND2_X1 U1121 ( .A1(n1416), .A2(n1147), .ZN(n1297) );
NAND2_X1 U1122 ( .A1(G475), .A2(n1417), .ZN(n1147) );
XOR2_X1 U1123 ( .A(n1146), .B(KEYINPUT25), .Z(n1416) );
OR2_X1 U1124 ( .A1(n1417), .A2(G475), .ZN(n1146) );
NAND2_X1 U1125 ( .A1(n1212), .A2(n1256), .ZN(n1417) );
INV_X1 U1126 ( .A(G902), .ZN(n1256) );
XNOR2_X1 U1127 ( .A(n1418), .B(n1419), .ZN(n1212) );
XOR2_X1 U1128 ( .A(n1420), .B(n1421), .Z(n1419) );
XNOR2_X1 U1129 ( .A(n1331), .B(G131), .ZN(n1421) );
INV_X1 U1130 ( .A(G146), .ZN(n1331) );
NOR2_X1 U1131 ( .A1(KEYINPUT35), .A2(G143), .ZN(n1420) );
XOR2_X1 U1132 ( .A(n1422), .B(n1423), .Z(n1418) );
AND2_X1 U1133 ( .A1(G214), .A2(n1347), .ZN(n1423) );
NOR2_X1 U1134 ( .A1(G953), .A2(G237), .ZN(n1347) );
XOR2_X1 U1135 ( .A(n1424), .B(n1425), .Z(n1422) );
NOR2_X1 U1136 ( .A1(n1426), .A2(n1427), .ZN(n1425) );
NOR2_X1 U1137 ( .A1(n1428), .A2(n1173), .ZN(n1427) );
NAND2_X1 U1138 ( .A1(G140), .A2(n1340), .ZN(n1173) );
NOR2_X1 U1139 ( .A1(n1429), .A2(n1340), .ZN(n1426) );
INV_X1 U1140 ( .A(n1172), .ZN(n1340) );
XOR2_X1 U1141 ( .A(G125), .B(KEYINPUT23), .Z(n1172) );
NOR2_X1 U1142 ( .A1(n1240), .A2(n1428), .ZN(n1429) );
INV_X1 U1143 ( .A(KEYINPUT12), .ZN(n1428) );
INV_X1 U1144 ( .A(G140), .ZN(n1240) );
NAND2_X1 U1145 ( .A1(n1430), .A2(n1431), .ZN(n1424) );
NAND2_X1 U1146 ( .A1(n1432), .A2(n1433), .ZN(n1431) );
NAND2_X1 U1147 ( .A1(KEYINPUT26), .A2(n1434), .ZN(n1433) );
NAND2_X1 U1148 ( .A1(n1435), .A2(n1436), .ZN(n1434) );
INV_X1 U1149 ( .A(n1437), .ZN(n1432) );
NAND2_X1 U1150 ( .A1(n1438), .A2(n1439), .ZN(n1430) );
NAND2_X1 U1151 ( .A1(n1436), .A2(n1440), .ZN(n1439) );
NAND2_X1 U1152 ( .A1(KEYINPUT26), .A2(n1437), .ZN(n1440) );
XOR2_X1 U1153 ( .A(G104), .B(KEYINPUT31), .Z(n1437) );
INV_X1 U1154 ( .A(KEYINPUT41), .ZN(n1436) );
INV_X1 U1155 ( .A(n1435), .ZN(n1438) );
NAND2_X1 U1156 ( .A1(n1441), .A2(n1442), .ZN(n1435) );
NAND2_X1 U1157 ( .A1(G122), .A2(n1319), .ZN(n1442) );
XOR2_X1 U1158 ( .A(KEYINPUT48), .B(n1443), .Z(n1441) );
NOR2_X1 U1159 ( .A1(G122), .A2(n1319), .ZN(n1443) );
INV_X1 U1160 ( .A(G113), .ZN(n1319) );
endmodule


