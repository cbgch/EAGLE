//Key = 0001111100010000001111110100001011010000011000000101000010100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316;

XNOR2_X1 U724 ( .A(G107), .B(n992), .ZN(G9) );
NOR2_X1 U725 ( .A1(n993), .A2(n994), .ZN(G75) );
NOR4_X1 U726 ( .A1(n995), .A2(n996), .A3(n997), .A4(n998), .ZN(n994) );
NOR2_X1 U727 ( .A1(KEYINPUT42), .A2(n999), .ZN(n997) );
NOR3_X1 U728 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n999) );
NAND3_X1 U729 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1000) );
NAND4_X1 U730 ( .A1(n1006), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n995) );
NAND2_X1 U731 ( .A1(n1010), .A2(n1011), .ZN(n1006) );
NAND2_X1 U732 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NAND3_X1 U733 ( .A1(n1004), .A2(n1014), .A3(n1015), .ZN(n1013) );
NAND2_X1 U734 ( .A1(n1016), .A2(n1017), .ZN(n1014) );
NAND2_X1 U735 ( .A1(n1005), .A2(n1018), .ZN(n1017) );
NAND2_X1 U736 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U737 ( .A1(KEYINPUT42), .A2(n1003), .ZN(n1020) );
NAND2_X1 U738 ( .A1(n1021), .A2(n1022), .ZN(n1016) );
NAND2_X1 U739 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND3_X1 U741 ( .A1(n1021), .A2(n1027), .A3(n1005), .ZN(n1012) );
NAND2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U743 ( .A1(n1015), .A2(n1030), .ZN(n1029) );
NAND2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U745 ( .A1(n1004), .A2(n1033), .ZN(n1028) );
NAND2_X1 U746 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NAND2_X1 U747 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
INV_X1 U748 ( .A(n1002), .ZN(n1010) );
AND3_X1 U749 ( .A1(n1008), .A2(n1009), .A3(n1038), .ZN(n993) );
NAND4_X1 U750 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1008) );
AND4_X1 U751 ( .A1(n1043), .A2(n1044), .A3(n1004), .A4(n1045), .ZN(n1042) );
XNOR2_X1 U752 ( .A(G469), .B(n1046), .ZN(n1041) );
NOR2_X1 U753 ( .A1(KEYINPUT15), .A2(n1047), .ZN(n1046) );
XNOR2_X1 U754 ( .A(n1048), .B(n1049), .ZN(n1040) );
XOR2_X1 U755 ( .A(n1050), .B(n1051), .Z(n1039) );
NOR2_X1 U756 ( .A1(KEYINPUT17), .A2(n1052), .ZN(n1051) );
XOR2_X1 U757 ( .A(n1053), .B(n1054), .Z(G72) );
NOR2_X1 U758 ( .A1(n1055), .A2(n1009), .ZN(n1054) );
AND2_X1 U759 ( .A1(G227), .A2(G900), .ZN(n1055) );
NAND2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1053) );
OR3_X1 U761 ( .A1(n1058), .A2(G953), .A3(n1059), .ZN(n1057) );
NAND3_X1 U762 ( .A1(n1060), .A2(n1061), .A3(n1059), .ZN(n1056) );
XOR2_X1 U763 ( .A(n1062), .B(n1063), .Z(n1059) );
NOR2_X1 U764 ( .A1(KEYINPUT24), .A2(n1064), .ZN(n1063) );
NAND2_X1 U765 ( .A1(G953), .A2(n1065), .ZN(n1061) );
XNOR2_X1 U766 ( .A(n1058), .B(KEYINPUT32), .ZN(n1060) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(G69) );
NAND2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
OR2_X1 U769 ( .A1(n1009), .A2(G224), .ZN(n1069) );
NAND3_X1 U770 ( .A1(G953), .A2(n1070), .A3(n1071), .ZN(n1066) );
INV_X1 U771 ( .A(n1068), .ZN(n1071) );
XNOR2_X1 U772 ( .A(n1072), .B(n1073), .ZN(n1068) );
NOR3_X1 U773 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1073) );
NOR2_X1 U774 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U775 ( .A(n1079), .B(KEYINPUT49), .Z(n1078) );
NOR2_X1 U776 ( .A1(n1080), .A2(n1081), .ZN(n1075) );
XOR2_X1 U777 ( .A(n1079), .B(KEYINPUT8), .Z(n1081) );
XOR2_X1 U778 ( .A(n1082), .B(n1083), .Z(n1079) );
XNOR2_X1 U779 ( .A(KEYINPUT0), .B(n1084), .ZN(n1082) );
NOR2_X1 U780 ( .A1(KEYINPUT46), .A2(n1085), .ZN(n1084) );
NOR2_X1 U781 ( .A1(G898), .A2(n1009), .ZN(n1074) );
NAND2_X1 U782 ( .A1(n1086), .A2(n1009), .ZN(n1072) );
XOR2_X1 U783 ( .A(n1087), .B(KEYINPUT57), .Z(n1086) );
NAND2_X1 U784 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U785 ( .A(n1007), .B(KEYINPUT28), .Z(n1088) );
NAND2_X1 U786 ( .A1(G898), .A2(G224), .ZN(n1070) );
NOR2_X1 U787 ( .A1(n1090), .A2(n1091), .ZN(G66) );
XOR2_X1 U788 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U789 ( .A1(n1094), .A2(G217), .ZN(n1092) );
NOR2_X1 U790 ( .A1(n1090), .A2(n1095), .ZN(G63) );
XOR2_X1 U791 ( .A(n1096), .B(n1097), .Z(n1095) );
AND2_X1 U792 ( .A1(G478), .A2(n1094), .ZN(n1096) );
NOR3_X1 U793 ( .A1(n1098), .A2(n1099), .A3(n1100), .ZN(G60) );
AND2_X1 U794 ( .A1(KEYINPUT20), .A2(n1090), .ZN(n1100) );
NOR3_X1 U795 ( .A1(KEYINPUT20), .A2(n1009), .A3(n1038), .ZN(n1099) );
INV_X1 U796 ( .A(G952), .ZN(n1038) );
XOR2_X1 U797 ( .A(n1101), .B(n1102), .Z(n1098) );
NOR2_X1 U798 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U799 ( .A(G475), .B(KEYINPUT55), .ZN(n1103) );
NAND2_X1 U800 ( .A1(KEYINPUT61), .A2(n1105), .ZN(n1101) );
XNOR2_X1 U801 ( .A(G104), .B(n1106), .ZN(G6) );
NOR2_X1 U802 ( .A1(n1090), .A2(n1107), .ZN(G57) );
XOR2_X1 U803 ( .A(n1108), .B(n1109), .Z(n1107) );
XOR2_X1 U804 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U805 ( .A1(n1094), .A2(G472), .ZN(n1110) );
XOR2_X1 U806 ( .A(n1112), .B(n1113), .Z(n1108) );
NOR2_X1 U807 ( .A1(KEYINPUT1), .A2(n1114), .ZN(n1113) );
XNOR2_X1 U808 ( .A(n1115), .B(n1116), .ZN(n1112) );
NOR2_X1 U809 ( .A1(n1090), .A2(n1117), .ZN(G54) );
XOR2_X1 U810 ( .A(n1118), .B(n1119), .Z(n1117) );
XOR2_X1 U811 ( .A(n1120), .B(n1121), .Z(n1119) );
XNOR2_X1 U812 ( .A(n1122), .B(n1123), .ZN(n1121) );
NAND3_X1 U813 ( .A1(KEYINPUT21), .A2(n1124), .A3(n1125), .ZN(n1122) );
XOR2_X1 U814 ( .A(n1126), .B(KEYINPUT48), .Z(n1125) );
NAND2_X1 U815 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
OR2_X1 U816 ( .A1(n1128), .A2(n1127), .ZN(n1124) );
XNOR2_X1 U817 ( .A(G128), .B(n1129), .ZN(n1127) );
XOR2_X1 U818 ( .A(n1130), .B(n1131), .Z(n1118) );
XOR2_X1 U819 ( .A(KEYINPUT34), .B(n1132), .Z(n1131) );
NAND3_X1 U820 ( .A1(n1094), .A2(G469), .A3(KEYINPUT23), .ZN(n1130) );
INV_X1 U821 ( .A(n1104), .ZN(n1094) );
NOR2_X1 U822 ( .A1(n1090), .A2(n1133), .ZN(G51) );
XOR2_X1 U823 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U824 ( .A1(KEYINPUT53), .A2(n1136), .ZN(n1135) );
XOR2_X1 U825 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U826 ( .A1(KEYINPUT45), .A2(n1139), .ZN(n1137) );
OR2_X1 U827 ( .A1(n1104), .A2(n1052), .ZN(n1134) );
NAND2_X1 U828 ( .A1(G902), .A2(n1140), .ZN(n1104) );
NAND3_X1 U829 ( .A1(n1058), .A2(n1007), .A3(n1089), .ZN(n1140) );
INV_X1 U830 ( .A(n996), .ZN(n1089) );
NAND4_X1 U831 ( .A1(n1141), .A2(n1142), .A3(n992), .A4(n1143), .ZN(n996) );
NOR3_X1 U832 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1143) );
NOR2_X1 U833 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND4_X1 U834 ( .A1(n1149), .A2(n1004), .A3(n1150), .A4(n1034), .ZN(n1148) );
INV_X1 U835 ( .A(KEYINPUT29), .ZN(n1147) );
NOR2_X1 U836 ( .A1(KEYINPUT29), .A2(n1106), .ZN(n1145) );
NAND4_X1 U837 ( .A1(n1149), .A2(n1151), .A3(n1004), .A4(n1150), .ZN(n1106) );
NAND3_X1 U838 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1144) );
OR2_X1 U839 ( .A1(n1155), .A2(KEYINPUT62), .ZN(n1154) );
NAND2_X1 U840 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
NAND2_X1 U841 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NAND2_X1 U842 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U843 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U844 ( .A1(KEYINPUT62), .A2(n1019), .ZN(n1163) );
NAND2_X1 U845 ( .A1(KEYINPUT58), .A2(n1164), .ZN(n1158) );
NAND3_X1 U846 ( .A1(n1164), .A2(n1165), .A3(n1031), .ZN(n1152) );
INV_X1 U847 ( .A(n1156), .ZN(n1031) );
INV_X1 U848 ( .A(KEYINPUT58), .ZN(n1165) );
NAND4_X1 U849 ( .A1(n1151), .A2(n1003), .A3(n1004), .A4(n1150), .ZN(n992) );
INV_X1 U850 ( .A(n998), .ZN(n1058) );
NAND4_X1 U851 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n998) );
NOR4_X1 U852 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
NAND2_X1 U853 ( .A1(n1151), .A2(n1174), .ZN(n1168) );
NAND2_X1 U854 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NAND3_X1 U855 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
NAND2_X1 U856 ( .A1(n1180), .A2(n1149), .ZN(n1175) );
NAND3_X1 U857 ( .A1(n1181), .A2(n1182), .A3(n1015), .ZN(n1166) );
NOR2_X1 U858 ( .A1(n1009), .A2(G952), .ZN(n1090) );
NAND2_X1 U859 ( .A1(n1183), .A2(n1184), .ZN(G48) );
NAND2_X1 U860 ( .A1(G146), .A2(n1185), .ZN(n1184) );
XOR2_X1 U861 ( .A(KEYINPUT19), .B(n1186), .Z(n1183) );
NOR2_X1 U862 ( .A1(G146), .A2(n1185), .ZN(n1186) );
NAND2_X1 U863 ( .A1(n1151), .A2(n1187), .ZN(n1185) );
XOR2_X1 U864 ( .A(KEYINPUT12), .B(n1188), .Z(n1187) );
NOR2_X1 U865 ( .A1(n1019), .A2(n1189), .ZN(n1188) );
INV_X1 U866 ( .A(n1149), .ZN(n1019) );
XNOR2_X1 U867 ( .A(G143), .B(n1190), .ZN(G45) );
NAND4_X1 U868 ( .A1(n1177), .A2(n1179), .A3(n1191), .A4(n1178), .ZN(n1190) );
XNOR2_X1 U869 ( .A(KEYINPUT31), .B(n1034), .ZN(n1191) );
XOR2_X1 U870 ( .A(G140), .B(n1192), .Z(G42) );
NOR3_X1 U871 ( .A1(n1193), .A2(n1023), .A3(n1194), .ZN(n1192) );
XNOR2_X1 U872 ( .A(KEYINPUT33), .B(n1001), .ZN(n1193) );
INV_X1 U873 ( .A(n1015), .ZN(n1001) );
XNOR2_X1 U874 ( .A(G137), .B(n1167), .ZN(G39) );
NAND3_X1 U875 ( .A1(n1180), .A2(n1021), .A3(n1015), .ZN(n1167) );
INV_X1 U876 ( .A(n1189), .ZN(n1180) );
XOR2_X1 U877 ( .A(G134), .B(n1173), .Z(G36) );
AND3_X1 U878 ( .A1(n1015), .A2(n1003), .A3(n1179), .ZN(n1173) );
XOR2_X1 U879 ( .A(G131), .B(n1172), .Z(G33) );
AND3_X1 U880 ( .A1(n1015), .A2(n1149), .A3(n1179), .ZN(n1172) );
AND3_X1 U881 ( .A1(n1182), .A2(n1195), .A3(n1156), .ZN(n1179) );
NOR2_X1 U882 ( .A1(n1196), .A2(n1036), .ZN(n1015) );
XOR2_X1 U883 ( .A(G128), .B(n1171), .Z(G30) );
NOR3_X1 U884 ( .A1(n1034), .A2(n1162), .A3(n1189), .ZN(n1171) );
NAND4_X1 U885 ( .A1(n1182), .A2(n1197), .A3(n1198), .A4(n1195), .ZN(n1189) );
INV_X1 U886 ( .A(n1003), .ZN(n1162) );
INV_X1 U887 ( .A(n1151), .ZN(n1034) );
XNOR2_X1 U888 ( .A(G101), .B(n1199), .ZN(G3) );
NAND2_X1 U889 ( .A1(n1200), .A2(n1164), .ZN(n1199) );
XNOR2_X1 U890 ( .A(n1156), .B(KEYINPUT22), .ZN(n1200) );
XOR2_X1 U891 ( .A(n1201), .B(n1170), .Z(G27) );
AND3_X1 U892 ( .A1(n1005), .A2(n1151), .A3(n1181), .ZN(n1170) );
INV_X1 U893 ( .A(n1194), .ZN(n1181) );
NAND3_X1 U894 ( .A1(n1202), .A2(n1195), .A3(n1149), .ZN(n1194) );
NAND2_X1 U895 ( .A1(n1002), .A2(n1203), .ZN(n1195) );
NAND4_X1 U896 ( .A1(G953), .A2(G902), .A3(n1065), .A4(n1204), .ZN(n1203) );
XOR2_X1 U897 ( .A(KEYINPUT41), .B(G900), .Z(n1065) );
NAND2_X1 U898 ( .A1(KEYINPUT5), .A2(n1205), .ZN(n1201) );
XNOR2_X1 U899 ( .A(G122), .B(n1007), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1177), .A2(n1160), .A3(n1004), .A4(n1178), .ZN(n1007) );
NOR2_X1 U901 ( .A1(n1198), .A2(n1197), .ZN(n1004) );
XNOR2_X1 U902 ( .A(n1141), .B(n1206), .ZN(G21) );
NOR2_X1 U903 ( .A1(KEYINPUT54), .A2(n1207), .ZN(n1206) );
NAND4_X1 U904 ( .A1(n1160), .A2(n1021), .A3(n1197), .A4(n1198), .ZN(n1141) );
XNOR2_X1 U905 ( .A(G116), .B(n1208), .ZN(G18) );
NAND4_X1 U906 ( .A1(n1156), .A2(n1005), .A3(n1209), .A4(n1003), .ZN(n1208) );
NOR2_X1 U907 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XNOR2_X1 U908 ( .A(n1151), .B(KEYINPUT26), .ZN(n1211) );
XOR2_X1 U909 ( .A(n1155), .B(n1212), .Z(G15) );
NAND2_X1 U910 ( .A1(KEYINPUT25), .A2(G113), .ZN(n1212) );
NAND3_X1 U911 ( .A1(n1149), .A2(n1160), .A3(n1156), .ZN(n1155) );
NOR2_X1 U912 ( .A1(n1197), .A2(n1213), .ZN(n1156) );
AND3_X1 U913 ( .A1(n1151), .A2(n1214), .A3(n1005), .ZN(n1160) );
NOR2_X1 U914 ( .A1(n1215), .A2(n1025), .ZN(n1005) );
NOR2_X1 U915 ( .A1(n1216), .A2(n1178), .ZN(n1149) );
XNOR2_X1 U916 ( .A(G110), .B(n1142), .ZN(G12) );
NAND2_X1 U917 ( .A1(n1164), .A2(n1202), .ZN(n1142) );
INV_X1 U918 ( .A(n1032), .ZN(n1202) );
NAND2_X1 U919 ( .A1(n1213), .A2(n1197), .ZN(n1032) );
XNOR2_X1 U920 ( .A(n1217), .B(n1218), .ZN(n1197) );
NOR2_X1 U921 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
INV_X1 U922 ( .A(G217), .ZN(n1220) );
XOR2_X1 U923 ( .A(n1221), .B(KEYINPUT4), .Z(n1219) );
NAND2_X1 U924 ( .A1(n1093), .A2(n1222), .ZN(n1217) );
XNOR2_X1 U925 ( .A(n1223), .B(n1224), .ZN(n1093) );
XOR2_X1 U926 ( .A(n1225), .B(n1226), .Z(n1224) );
XNOR2_X1 U927 ( .A(n1227), .B(n1228), .ZN(n1226) );
NOR2_X1 U928 ( .A1(KEYINPUT36), .A2(n1207), .ZN(n1228) );
NOR2_X1 U929 ( .A1(KEYINPUT38), .A2(n1229), .ZN(n1227) );
XOR2_X1 U930 ( .A(n1230), .B(n1062), .Z(n1229) );
XNOR2_X1 U931 ( .A(G146), .B(KEYINPUT43), .ZN(n1230) );
NAND2_X1 U932 ( .A1(G221), .A2(n1231), .ZN(n1225) );
XNOR2_X1 U933 ( .A(n1232), .B(n1233), .ZN(n1223) );
INV_X1 U934 ( .A(n1198), .ZN(n1213) );
XNOR2_X1 U935 ( .A(n1234), .B(G472), .ZN(n1198) );
NAND2_X1 U936 ( .A1(n1235), .A2(n1222), .ZN(n1234) );
XOR2_X1 U937 ( .A(n1236), .B(n1237), .Z(n1235) );
XOR2_X1 U938 ( .A(n1115), .B(n1238), .Z(n1237) );
NAND2_X1 U939 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
OR2_X1 U940 ( .A1(n1114), .A2(n1111), .ZN(n1240) );
XOR2_X1 U941 ( .A(n1241), .B(KEYINPUT2), .Z(n1239) );
NAND2_X1 U942 ( .A1(n1111), .A2(n1114), .ZN(n1241) );
XNOR2_X1 U943 ( .A(n1242), .B(n1120), .ZN(n1114) );
XOR2_X1 U944 ( .A(G137), .B(n1243), .Z(n1120) );
XOR2_X1 U945 ( .A(n1139), .B(KEYINPUT9), .Z(n1242) );
XNOR2_X1 U946 ( .A(n1244), .B(G113), .ZN(n1111) );
NAND2_X1 U947 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND2_X1 U948 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
XNOR2_X1 U949 ( .A(KEYINPUT3), .B(n1249), .ZN(n1248) );
XNOR2_X1 U950 ( .A(G119), .B(KEYINPUT27), .ZN(n1247) );
NAND2_X1 U951 ( .A1(n1250), .A2(n1251), .ZN(n1245) );
XNOR2_X1 U952 ( .A(KEYINPUT3), .B(G116), .ZN(n1251) );
XNOR2_X1 U953 ( .A(G119), .B(KEYINPUT56), .ZN(n1250) );
NAND2_X1 U954 ( .A1(n1252), .A2(G210), .ZN(n1115) );
NAND2_X1 U955 ( .A1(KEYINPUT11), .A2(n1116), .ZN(n1236) );
INV_X1 U956 ( .A(G101), .ZN(n1116) );
AND3_X1 U957 ( .A1(n1150), .A2(n1021), .A3(n1151), .ZN(n1164) );
NOR2_X1 U958 ( .A1(n1037), .A2(n1036), .ZN(n1151) );
INV_X1 U959 ( .A(n1044), .ZN(n1036) );
NAND2_X1 U960 ( .A1(G214), .A2(n1253), .ZN(n1044) );
INV_X1 U961 ( .A(n1196), .ZN(n1037) );
XOR2_X1 U962 ( .A(n1050), .B(n1052), .Z(n1196) );
NAND2_X1 U963 ( .A1(G210), .A2(n1253), .ZN(n1052) );
NAND2_X1 U964 ( .A1(n1254), .A2(n1222), .ZN(n1253) );
INV_X1 U965 ( .A(G237), .ZN(n1254) );
NAND2_X1 U966 ( .A1(n1255), .A2(n1222), .ZN(n1050) );
XNOR2_X1 U967 ( .A(n1138), .B(n1256), .ZN(n1255) );
XOR2_X1 U968 ( .A(n1139), .B(KEYINPUT18), .Z(n1256) );
NAND2_X1 U969 ( .A1(n1257), .A2(n1258), .ZN(n1139) );
NAND2_X1 U970 ( .A1(G128), .A2(n1259), .ZN(n1258) );
XOR2_X1 U971 ( .A(KEYINPUT30), .B(n1260), .Z(n1257) );
NOR2_X1 U972 ( .A1(G128), .A2(n1259), .ZN(n1260) );
NAND2_X1 U973 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
NAND2_X1 U974 ( .A1(G146), .A2(n1263), .ZN(n1262) );
XOR2_X1 U975 ( .A(KEYINPUT7), .B(n1264), .Z(n1261) );
NOR2_X1 U976 ( .A1(G146), .A2(n1263), .ZN(n1264) );
XNOR2_X1 U977 ( .A(n1265), .B(n1266), .ZN(n1138) );
XNOR2_X1 U978 ( .A(n1205), .B(n1267), .ZN(n1266) );
NOR2_X1 U979 ( .A1(KEYINPUT13), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U980 ( .A(n1083), .B(n1085), .ZN(n1268) );
XOR2_X1 U981 ( .A(n1269), .B(KEYINPUT44), .Z(n1085) );
NAND3_X1 U982 ( .A1(n1270), .A2(n1271), .A3(n1272), .ZN(n1269) );
NAND2_X1 U983 ( .A1(KEYINPUT40), .A2(G101), .ZN(n1272) );
OR3_X1 U984 ( .A1(G101), .A2(KEYINPUT40), .A3(n1273), .ZN(n1271) );
NAND2_X1 U985 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
NAND2_X1 U986 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
INV_X1 U987 ( .A(KEYINPUT40), .ZN(n1276) );
XNOR2_X1 U988 ( .A(G101), .B(KEYINPUT60), .ZN(n1275) );
XOR2_X1 U989 ( .A(G113), .B(n1277), .Z(n1083) );
XNOR2_X1 U990 ( .A(n1207), .B(G116), .ZN(n1277) );
INV_X1 U991 ( .A(G119), .ZN(n1207) );
INV_X1 U992 ( .A(G125), .ZN(n1205) );
XNOR2_X1 U993 ( .A(n1278), .B(n1077), .ZN(n1265) );
INV_X1 U994 ( .A(n1080), .ZN(n1077) );
XOR2_X1 U995 ( .A(n1279), .B(n1280), .Z(n1080) );
XNOR2_X1 U996 ( .A(G122), .B(KEYINPUT10), .ZN(n1279) );
NAND2_X1 U997 ( .A1(G224), .A2(n1009), .ZN(n1278) );
NAND2_X1 U998 ( .A1(n1281), .A2(n1282), .ZN(n1021) );
OR3_X1 U999 ( .A1(n1177), .A2(n1178), .A3(KEYINPUT14), .ZN(n1282) );
NAND2_X1 U1000 ( .A1(KEYINPUT14), .A2(n1003), .ZN(n1281) );
NOR2_X1 U1001 ( .A1(n1177), .A2(n1045), .ZN(n1003) );
INV_X1 U1002 ( .A(n1178), .ZN(n1045) );
XNOR2_X1 U1003 ( .A(n1283), .B(G478), .ZN(n1178) );
OR2_X1 U1004 ( .A1(n1097), .A2(G902), .ZN(n1283) );
XNOR2_X1 U1005 ( .A(n1284), .B(n1285), .ZN(n1097) );
XOR2_X1 U1006 ( .A(G128), .B(n1286), .Z(n1285) );
XNOR2_X1 U1007 ( .A(n1263), .B(G134), .ZN(n1286) );
XOR2_X1 U1008 ( .A(n1287), .B(n1288), .Z(n1284) );
XNOR2_X1 U1009 ( .A(G107), .B(n1289), .ZN(n1288) );
NAND2_X1 U1010 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U1011 ( .A1(G116), .A2(n1292), .ZN(n1291) );
INV_X1 U1012 ( .A(G122), .ZN(n1292) );
XOR2_X1 U1013 ( .A(n1293), .B(KEYINPUT39), .Z(n1290) );
NAND2_X1 U1014 ( .A1(G122), .A2(n1249), .ZN(n1293) );
INV_X1 U1015 ( .A(G116), .ZN(n1249) );
NAND2_X1 U1016 ( .A1(G217), .A2(n1231), .ZN(n1287) );
AND2_X1 U1017 ( .A1(G234), .A2(n1009), .ZN(n1231) );
INV_X1 U1018 ( .A(n1216), .ZN(n1177) );
XOR2_X1 U1019 ( .A(n1294), .B(n1048), .Z(n1216) );
NAND2_X1 U1020 ( .A1(n1105), .A2(n1222), .ZN(n1048) );
XNOR2_X1 U1021 ( .A(n1295), .B(n1296), .ZN(n1105) );
XOR2_X1 U1022 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U1023 ( .A(G131), .B(G104), .Z(n1298) );
NOR2_X1 U1024 ( .A1(KEYINPUT50), .A2(n1299), .ZN(n1297) );
XNOR2_X1 U1025 ( .A(G113), .B(G122), .ZN(n1299) );
XOR2_X1 U1026 ( .A(n1300), .B(n1062), .Z(n1295) );
XOR2_X1 U1027 ( .A(G125), .B(G140), .Z(n1062) );
XOR2_X1 U1028 ( .A(n1301), .B(n1302), .Z(n1300) );
NAND2_X1 U1029 ( .A1(n1252), .A2(G214), .ZN(n1301) );
NOR2_X1 U1030 ( .A1(G953), .A2(G237), .ZN(n1252) );
NAND2_X1 U1031 ( .A1(KEYINPUT51), .A2(n1049), .ZN(n1294) );
INV_X1 U1032 ( .A(G475), .ZN(n1049) );
NOR2_X1 U1033 ( .A1(n1023), .A2(n1210), .ZN(n1150) );
INV_X1 U1034 ( .A(n1214), .ZN(n1210) );
NAND2_X1 U1035 ( .A1(n1002), .A2(n1303), .ZN(n1214) );
NAND4_X1 U1036 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1304), .ZN(n1303) );
INV_X1 U1037 ( .A(G898), .ZN(n1304) );
NAND3_X1 U1038 ( .A1(n1204), .A2(n1009), .A3(G952), .ZN(n1002) );
NAND2_X1 U1039 ( .A1(G237), .A2(G234), .ZN(n1204) );
INV_X1 U1040 ( .A(n1182), .ZN(n1023) );
NOR2_X1 U1041 ( .A1(n1026), .A2(n1025), .ZN(n1182) );
INV_X1 U1042 ( .A(n1043), .ZN(n1025) );
NAND2_X1 U1043 ( .A1(G221), .A2(n1221), .ZN(n1043) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1222), .ZN(n1221) );
INV_X1 U1045 ( .A(n1215), .ZN(n1026) );
XNOR2_X1 U1046 ( .A(n1047), .B(G469), .ZN(n1215) );
NAND2_X1 U1047 ( .A1(n1305), .A2(n1222), .ZN(n1047) );
INV_X1 U1048 ( .A(G902), .ZN(n1222) );
XOR2_X1 U1049 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U1050 ( .A(n1064), .B(n1308), .ZN(n1307) );
NOR2_X1 U1051 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NOR2_X1 U1052 ( .A1(KEYINPUT37), .A2(n1123), .ZN(n1310) );
INV_X1 U1053 ( .A(n1311), .ZN(n1123) );
NOR2_X1 U1054 ( .A1(KEYINPUT35), .A2(n1311), .ZN(n1309) );
XOR2_X1 U1055 ( .A(G140), .B(n1280), .Z(n1311) );
INV_X1 U1056 ( .A(n1232), .ZN(n1280) );
XOR2_X1 U1057 ( .A(G110), .B(KEYINPUT16), .Z(n1232) );
XOR2_X1 U1058 ( .A(n1312), .B(n1243), .Z(n1064) );
XOR2_X1 U1059 ( .A(G131), .B(G134), .Z(n1243) );
XNOR2_X1 U1060 ( .A(n1233), .B(n1129), .ZN(n1312) );
NOR2_X1 U1061 ( .A1(KEYINPUT59), .A2(n1313), .ZN(n1129) );
XOR2_X1 U1062 ( .A(KEYINPUT63), .B(n1302), .Z(n1313) );
XNOR2_X1 U1063 ( .A(n1263), .B(G146), .ZN(n1302) );
INV_X1 U1064 ( .A(G143), .ZN(n1263) );
XOR2_X1 U1065 ( .A(G137), .B(G128), .Z(n1233) );
XNOR2_X1 U1066 ( .A(n1132), .B(n1314), .ZN(n1306) );
XNOR2_X1 U1067 ( .A(KEYINPUT47), .B(n1315), .ZN(n1314) );
NOR2_X1 U1068 ( .A1(KEYINPUT52), .A2(n1316), .ZN(n1315) );
XNOR2_X1 U1069 ( .A(n1128), .B(KEYINPUT6), .ZN(n1316) );
XOR2_X1 U1070 ( .A(G101), .B(n1273), .Z(n1128) );
XOR2_X1 U1071 ( .A(G104), .B(G107), .Z(n1273) );
AND2_X1 U1072 ( .A1(G227), .A2(n1009), .ZN(n1132) );
INV_X1 U1073 ( .A(G953), .ZN(n1009) );
endmodule


