//Key = 1011011100011001010010010101110011110100110110100001011101100011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390;

XOR2_X1 U762 ( .A(n1056), .B(G107), .Z(G9) );
NAND2_X1 U763 ( .A1(KEYINPUT5), .A2(n1057), .ZN(n1056) );
NOR2_X1 U764 ( .A1(n1058), .A2(n1059), .ZN(G75) );
NOR3_X1 U765 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NAND3_X1 U766 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1060) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND3_X1 U769 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U770 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NAND2_X1 U771 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U772 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1068) );
NAND2_X1 U773 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NAND3_X1 U774 ( .A1(n1070), .A2(n1082), .A3(n1072), .ZN(n1080) );
NAND2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND3_X1 U776 ( .A1(n1085), .A2(n1086), .A3(n1075), .ZN(n1077) );
NAND2_X1 U777 ( .A1(n1072), .A2(n1087), .ZN(n1086) );
OR2_X1 U778 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U779 ( .A1(n1070), .A2(n1090), .ZN(n1085) );
NAND2_X1 U780 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
INV_X1 U782 ( .A(n1095), .ZN(n1066) );
NOR3_X1 U783 ( .A1(n1096), .A2(G953), .A3(G952), .ZN(n1058) );
INV_X1 U784 ( .A(n1063), .ZN(n1096) );
NAND4_X1 U785 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1063) );
NOR4_X1 U786 ( .A1(n1093), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1104), .B(KEYINPUT17), .Z(n1103) );
NAND2_X1 U788 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U789 ( .A(KEYINPUT22), .B(n1107), .Z(n1105) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(n1102) );
NOR2_X1 U791 ( .A1(KEYINPUT38), .A2(n1110), .ZN(n1109) );
XNOR2_X1 U792 ( .A(KEYINPUT52), .B(n1111), .ZN(n1110) );
NOR2_X1 U793 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
XOR2_X1 U794 ( .A(G478), .B(KEYINPUT56), .Z(n1107) );
NOR3_X1 U795 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1099) );
NOR2_X1 U796 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
INV_X1 U797 ( .A(KEYINPUT18), .ZN(n1116) );
NOR3_X1 U798 ( .A1(n1117), .A2(n1118), .A3(n1083), .ZN(n1115) );
NOR2_X1 U799 ( .A1(KEYINPUT18), .A2(n1075), .ZN(n1113) );
XOR2_X1 U800 ( .A(n1119), .B(n1120), .Z(n1112) );
XOR2_X1 U801 ( .A(n1121), .B(KEYINPUT53), .Z(n1120) );
NAND2_X1 U802 ( .A1(KEYINPUT25), .A2(n1122), .ZN(n1119) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(G72) );
XOR2_X1 U804 ( .A(n1125), .B(n1126), .Z(n1124) );
AND2_X1 U805 ( .A1(n1061), .A2(n1064), .ZN(n1126) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1128) );
XNOR2_X1 U808 ( .A(G134), .B(n1131), .ZN(n1130) );
NAND2_X1 U809 ( .A1(n1132), .A2(KEYINPUT2), .ZN(n1131) );
XOR2_X1 U810 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U811 ( .A1(G140), .A2(KEYINPUT59), .ZN(n1134) );
XOR2_X1 U812 ( .A(n1135), .B(n1136), .Z(n1129) );
NOR2_X1 U813 ( .A1(G900), .A2(n1064), .ZN(n1127) );
NOR2_X1 U814 ( .A1(n1137), .A2(n1064), .ZN(n1123) );
NOR2_X1 U815 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(G69) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U818 ( .A1(n1144), .A2(n1064), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U820 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(n1148) );
NAND2_X1 U822 ( .A1(KEYINPUT40), .A2(n1151), .ZN(n1149) );
XOR2_X1 U823 ( .A(n1152), .B(KEYINPUT50), .Z(n1147) );
NAND2_X1 U824 ( .A1(G953), .A2(n1146), .ZN(n1152) );
NAND2_X1 U825 ( .A1(n1064), .A2(n1062), .ZN(n1140) );
NOR2_X1 U826 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XNOR2_X1 U827 ( .A(n1155), .B(n1156), .ZN(n1154) );
XNOR2_X1 U828 ( .A(n1157), .B(KEYINPUT4), .ZN(n1156) );
NAND3_X1 U829 ( .A1(n1158), .A2(n1159), .A3(KEYINPUT37), .ZN(n1157) );
NOR2_X1 U830 ( .A1(n1153), .A2(n1160), .ZN(G63) );
XOR2_X1 U831 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U832 ( .A1(KEYINPUT48), .A2(n1163), .ZN(n1162) );
AND2_X1 U833 ( .A1(G478), .A2(n1158), .ZN(n1161) );
NOR2_X1 U834 ( .A1(n1153), .A2(n1164), .ZN(G60) );
XOR2_X1 U835 ( .A(n1165), .B(n1166), .Z(n1164) );
AND2_X1 U836 ( .A1(G475), .A2(n1158), .ZN(n1165) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(G6) );
NOR2_X1 U838 ( .A1(n1153), .A2(n1169), .ZN(G57) );
XOR2_X1 U839 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1171) );
NAND2_X1 U841 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
INV_X1 U842 ( .A(n1176), .ZN(n1175) );
XOR2_X1 U843 ( .A(KEYINPUT44), .B(n1177), .Z(n1174) );
NAND3_X1 U844 ( .A1(n1178), .A2(n1179), .A3(n1180), .ZN(n1172) );
NAND2_X1 U845 ( .A1(KEYINPUT9), .A2(n1181), .ZN(n1180) );
NAND2_X1 U846 ( .A1(n1182), .A2(n1183), .ZN(n1179) );
OR3_X1 U847 ( .A1(n1183), .A2(KEYINPUT9), .A3(n1182), .ZN(n1178) );
OR2_X1 U848 ( .A1(KEYINPUT31), .A2(n1181), .ZN(n1183) );
NOR2_X1 U849 ( .A1(n1108), .A2(n1184), .ZN(n1170) );
INV_X1 U850 ( .A(G472), .ZN(n1108) );
NOR2_X1 U851 ( .A1(n1153), .A2(n1185), .ZN(G54) );
XOR2_X1 U852 ( .A(n1186), .B(n1187), .Z(n1185) );
NOR2_X1 U853 ( .A1(n1117), .A2(n1184), .ZN(n1187) );
INV_X1 U854 ( .A(G469), .ZN(n1117) );
NOR2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
XOR2_X1 U856 ( .A(n1190), .B(KEYINPUT15), .Z(n1189) );
NAND2_X1 U857 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U858 ( .A(KEYINPUT32), .B(n1193), .ZN(n1192) );
NOR2_X1 U859 ( .A1(n1193), .A2(n1191), .ZN(n1188) );
XOR2_X1 U860 ( .A(n1194), .B(n1195), .Z(n1191) );
XOR2_X1 U861 ( .A(n1196), .B(n1197), .Z(n1193) );
XOR2_X1 U862 ( .A(G140), .B(n1198), .Z(n1197) );
NAND2_X1 U863 ( .A1(KEYINPUT28), .A2(n1199), .ZN(n1196) );
NOR2_X1 U864 ( .A1(n1153), .A2(n1200), .ZN(G51) );
XOR2_X1 U865 ( .A(n1201), .B(n1202), .Z(n1200) );
NAND2_X1 U866 ( .A1(n1158), .A2(n1203), .ZN(n1202) );
INV_X1 U867 ( .A(n1184), .ZN(n1158) );
NAND2_X1 U868 ( .A1(G902), .A2(n1204), .ZN(n1184) );
OR2_X1 U869 ( .A1(n1062), .A2(n1061), .ZN(n1204) );
NAND4_X1 U870 ( .A1(n1205), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1061) );
AND4_X1 U871 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208) );
NAND2_X1 U872 ( .A1(n1213), .A2(n1214), .ZN(n1207) );
NAND2_X1 U873 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NAND2_X1 U874 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XNOR2_X1 U875 ( .A(n1219), .B(KEYINPUT7), .ZN(n1217) );
NAND2_X1 U876 ( .A1(n1072), .A2(n1088), .ZN(n1215) );
NAND4_X1 U877 ( .A1(n1220), .A2(n1168), .A3(n1221), .A4(n1222), .ZN(n1062) );
NOR4_X1 U878 ( .A1(n1223), .A2(n1224), .A3(n1225), .A4(n1226), .ZN(n1222) );
INV_X1 U879 ( .A(n1057), .ZN(n1223) );
NAND3_X1 U880 ( .A1(n1076), .A2(n1070), .A3(n1227), .ZN(n1057) );
NAND2_X1 U881 ( .A1(n1228), .A2(n1229), .ZN(n1221) );
NAND2_X1 U882 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND3_X1 U883 ( .A1(n1079), .A2(n1232), .A3(n1219), .ZN(n1231) );
XOR2_X1 U884 ( .A(KEYINPUT14), .B(n1075), .Z(n1232) );
NAND2_X1 U885 ( .A1(n1233), .A2(n1234), .ZN(n1230) );
XOR2_X1 U886 ( .A(KEYINPUT24), .B(n1088), .Z(n1234) );
NAND4_X1 U887 ( .A1(n1235), .A2(n1227), .A3(n1070), .A4(n1236), .ZN(n1168) );
NAND3_X1 U888 ( .A1(n1237), .A2(n1238), .A3(n1218), .ZN(n1220) );
NAND2_X1 U889 ( .A1(KEYINPUT12), .A2(n1239), .ZN(n1238) );
NAND2_X1 U890 ( .A1(n1240), .A2(n1241), .ZN(n1237) );
INV_X1 U891 ( .A(KEYINPUT12), .ZN(n1241) );
NAND2_X1 U892 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
NAND3_X1 U893 ( .A1(n1244), .A2(n1245), .A3(KEYINPUT23), .ZN(n1201) );
NAND2_X1 U894 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
NAND2_X1 U895 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
OR2_X1 U896 ( .A1(n1250), .A2(KEYINPUT58), .ZN(n1249) );
NAND3_X1 U897 ( .A1(n1251), .A2(n1252), .A3(KEYINPUT58), .ZN(n1244) );
NAND2_X1 U898 ( .A1(KEYINPUT27), .A2(n1253), .ZN(n1252) );
NAND2_X1 U899 ( .A1(n1254), .A2(n1248), .ZN(n1253) );
NAND2_X1 U900 ( .A1(n1248), .A2(n1250), .ZN(n1251) );
INV_X1 U901 ( .A(KEYINPUT27), .ZN(n1250) );
XNOR2_X1 U902 ( .A(n1255), .B(n1256), .ZN(n1248) );
NAND2_X1 U903 ( .A1(KEYINPUT46), .A2(n1257), .ZN(n1255) );
XOR2_X1 U904 ( .A(G125), .B(n1258), .Z(n1257) );
NOR2_X1 U905 ( .A1(n1064), .A2(G952), .ZN(n1153) );
XNOR2_X1 U906 ( .A(G146), .B(n1259), .ZN(G48) );
NAND2_X1 U907 ( .A1(n1213), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U908 ( .A(G143), .B(n1205), .ZN(G45) );
NAND4_X1 U909 ( .A1(n1261), .A2(n1088), .A3(n1262), .A4(n1218), .ZN(n1205) );
NOR2_X1 U910 ( .A1(n1235), .A2(n1263), .ZN(n1262) );
XOR2_X1 U911 ( .A(n1206), .B(n1264), .Z(G42) );
XOR2_X1 U912 ( .A(KEYINPUT0), .B(G140), .Z(n1264) );
NAND3_X1 U913 ( .A1(n1072), .A2(n1089), .A3(n1213), .ZN(n1206) );
XNOR2_X1 U914 ( .A(G137), .B(n1212), .ZN(G39) );
NAND4_X1 U915 ( .A1(n1072), .A2(n1261), .A3(n1219), .A4(n1079), .ZN(n1212) );
XNOR2_X1 U916 ( .A(G134), .B(n1211), .ZN(G36) );
NAND4_X1 U917 ( .A1(n1072), .A2(n1261), .A3(n1088), .A4(n1076), .ZN(n1211) );
NAND2_X1 U918 ( .A1(n1265), .A2(n1266), .ZN(G33) );
NAND2_X1 U919 ( .A1(G131), .A2(n1267), .ZN(n1266) );
XOR2_X1 U920 ( .A(n1268), .B(KEYINPUT21), .Z(n1265) );
OR2_X1 U921 ( .A1(n1267), .A2(G131), .ZN(n1268) );
NAND3_X1 U922 ( .A1(n1213), .A2(n1088), .A3(n1269), .ZN(n1267) );
XNOR2_X1 U923 ( .A(n1072), .B(KEYINPUT20), .ZN(n1269) );
NOR2_X1 U924 ( .A1(n1270), .A2(n1093), .ZN(n1072) );
INV_X1 U925 ( .A(n1094), .ZN(n1270) );
AND3_X1 U926 ( .A1(n1235), .A2(n1236), .A3(n1261), .ZN(n1213) );
XNOR2_X1 U927 ( .A(G128), .B(n1210), .ZN(G30) );
NAND3_X1 U928 ( .A1(n1260), .A2(n1076), .A3(n1261), .ZN(n1210) );
AND3_X1 U929 ( .A1(n1271), .A2(n1272), .A3(n1084), .ZN(n1261) );
INV_X1 U930 ( .A(n1273), .ZN(n1076) );
AND2_X1 U931 ( .A1(n1219), .A2(n1218), .ZN(n1260) );
XOR2_X1 U932 ( .A(G101), .B(n1226), .Z(G3) );
AND3_X1 U933 ( .A1(n1079), .A2(n1227), .A3(n1088), .ZN(n1226) );
XOR2_X1 U934 ( .A(n1133), .B(n1209), .Z(G27) );
NAND4_X1 U935 ( .A1(n1233), .A2(n1089), .A3(n1218), .A4(n1272), .ZN(n1209) );
NAND2_X1 U936 ( .A1(n1274), .A2(n1095), .ZN(n1272) );
NAND2_X1 U937 ( .A1(n1275), .A2(n1139), .ZN(n1274) );
INV_X1 U938 ( .A(G900), .ZN(n1139) );
INV_X1 U939 ( .A(n1073), .ZN(n1233) );
NAND2_X1 U940 ( .A1(n1276), .A2(n1277), .ZN(G24) );
NAND3_X1 U941 ( .A1(G122), .A2(n1278), .A3(n1279), .ZN(n1277) );
NAND2_X1 U942 ( .A1(n1280), .A2(n1281), .ZN(n1276) );
NAND2_X1 U943 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U944 ( .A1(G122), .A2(n1284), .ZN(n1283) );
INV_X1 U945 ( .A(KEYINPUT35), .ZN(n1284) );
NAND2_X1 U946 ( .A1(KEYINPUT35), .A2(n1285), .ZN(n1282) );
NAND2_X1 U947 ( .A1(G122), .A2(n1278), .ZN(n1285) );
INV_X1 U948 ( .A(KEYINPUT60), .ZN(n1278) );
INV_X1 U949 ( .A(n1279), .ZN(n1280) );
NAND2_X1 U950 ( .A1(n1286), .A2(n1218), .ZN(n1279) );
XOR2_X1 U951 ( .A(n1239), .B(KEYINPUT11), .Z(n1286) );
NAND2_X1 U952 ( .A1(n1243), .A2(n1287), .ZN(n1239) );
AND4_X1 U953 ( .A1(n1075), .A2(n1070), .A3(n1236), .A4(n1288), .ZN(n1243) );
NOR2_X1 U954 ( .A1(n1289), .A2(n1290), .ZN(n1070) );
XNOR2_X1 U955 ( .A(G119), .B(n1291), .ZN(G21) );
NAND4_X1 U956 ( .A1(n1219), .A2(n1075), .A3(n1079), .A4(n1228), .ZN(n1291) );
NOR2_X1 U957 ( .A1(n1292), .A2(n1098), .ZN(n1219) );
XOR2_X1 U958 ( .A(G116), .B(n1225), .Z(G18) );
NOR3_X1 U959 ( .A1(n1293), .A2(n1273), .A3(n1081), .ZN(n1225) );
INV_X1 U960 ( .A(n1075), .ZN(n1081) );
NAND2_X1 U961 ( .A1(n1263), .A2(n1288), .ZN(n1273) );
XOR2_X1 U962 ( .A(G113), .B(n1294), .Z(G15) );
NOR2_X1 U963 ( .A1(n1293), .A2(n1073), .ZN(n1294) );
NAND3_X1 U964 ( .A1(n1235), .A2(n1236), .A3(n1075), .ZN(n1073) );
NOR2_X1 U965 ( .A1(n1084), .A2(n1083), .ZN(n1075) );
INV_X1 U966 ( .A(n1271), .ZN(n1083) );
NAND2_X1 U967 ( .A1(n1088), .A2(n1228), .ZN(n1293) );
NOR2_X1 U968 ( .A1(n1289), .A2(n1292), .ZN(n1088) );
INV_X1 U969 ( .A(n1098), .ZN(n1289) );
NAND3_X1 U970 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(G12) );
NAND2_X1 U971 ( .A1(KEYINPUT45), .A2(n1298), .ZN(n1297) );
NAND3_X1 U972 ( .A1(n1224), .A2(n1299), .A3(n1199), .ZN(n1296) );
INV_X1 U973 ( .A(n1298), .ZN(n1224) );
NAND2_X1 U974 ( .A1(G110), .A2(n1300), .ZN(n1295) );
NAND2_X1 U975 ( .A1(n1301), .A2(n1299), .ZN(n1300) );
INV_X1 U976 ( .A(KEYINPUT45), .ZN(n1299) );
XOR2_X1 U977 ( .A(n1298), .B(KEYINPUT3), .Z(n1301) );
NAND3_X1 U978 ( .A1(n1089), .A2(n1227), .A3(n1079), .ZN(n1298) );
NOR2_X1 U979 ( .A1(n1288), .A2(n1236), .ZN(n1079) );
INV_X1 U980 ( .A(n1263), .ZN(n1236) );
XOR2_X1 U981 ( .A(n1097), .B(KEYINPUT1), .Z(n1263) );
XOR2_X1 U982 ( .A(n1302), .B(G475), .Z(n1097) );
OR2_X1 U983 ( .A1(n1166), .A2(G902), .ZN(n1302) );
XNOR2_X1 U984 ( .A(n1303), .B(n1304), .ZN(n1166) );
XOR2_X1 U985 ( .A(n1305), .B(n1306), .Z(n1304) );
XOR2_X1 U986 ( .A(n1307), .B(n1308), .Z(n1306) );
NOR2_X1 U987 ( .A1(G143), .A2(KEYINPUT10), .ZN(n1307) );
XOR2_X1 U988 ( .A(n1309), .B(n1310), .Z(n1305) );
NOR2_X1 U989 ( .A1(KEYINPUT61), .A2(n1133), .ZN(n1310) );
AND3_X1 U990 ( .A1(G214), .A2(n1064), .A3(n1311), .ZN(n1309) );
XOR2_X1 U991 ( .A(n1312), .B(n1313), .Z(n1303) );
XOR2_X1 U992 ( .A(G146), .B(G131), .Z(n1313) );
XOR2_X1 U993 ( .A(n1167), .B(n1314), .Z(n1312) );
NOR2_X1 U994 ( .A1(KEYINPUT30), .A2(n1315), .ZN(n1314) );
XOR2_X1 U995 ( .A(n1316), .B(G122), .Z(n1315) );
INV_X1 U996 ( .A(n1235), .ZN(n1288) );
XOR2_X1 U997 ( .A(n1106), .B(G478), .Z(n1235) );
NAND2_X1 U998 ( .A1(n1163), .A2(n1317), .ZN(n1106) );
XOR2_X1 U999 ( .A(n1318), .B(n1319), .Z(n1163) );
XOR2_X1 U1000 ( .A(G107), .B(n1320), .Z(n1319) );
NOR2_X1 U1001 ( .A1(KEYINPUT13), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1002 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1003 ( .A(G143), .B(G134), .Z(n1323) );
XOR2_X1 U1004 ( .A(n1324), .B(n1325), .Z(n1318) );
AND2_X1 U1005 ( .A1(n1326), .A2(G217), .ZN(n1325) );
NAND2_X1 U1006 ( .A1(KEYINPUT33), .A2(n1327), .ZN(n1324) );
XOR2_X1 U1007 ( .A(G122), .B(G116), .Z(n1327) );
AND3_X1 U1008 ( .A1(n1084), .A2(n1271), .A3(n1228), .ZN(n1227) );
NOR2_X1 U1009 ( .A1(n1091), .A2(n1242), .ZN(n1228) );
INV_X1 U1010 ( .A(n1287), .ZN(n1242) );
NAND2_X1 U1011 ( .A1(n1328), .A2(n1095), .ZN(n1287) );
NAND3_X1 U1012 ( .A1(n1329), .A2(n1064), .A3(G952), .ZN(n1095) );
NAND2_X1 U1013 ( .A1(n1275), .A2(n1146), .ZN(n1328) );
INV_X1 U1014 ( .A(G898), .ZN(n1146) );
AND3_X1 U1015 ( .A1(G953), .A2(n1329), .A3(n1330), .ZN(n1275) );
XOR2_X1 U1016 ( .A(n1317), .B(KEYINPUT54), .Z(n1330) );
NAND2_X1 U1017 ( .A1(G237), .A2(G234), .ZN(n1329) );
INV_X1 U1018 ( .A(n1218), .ZN(n1091) );
NOR2_X1 U1019 ( .A1(n1094), .A2(n1093), .ZN(n1218) );
AND2_X1 U1020 ( .A1(G214), .A2(n1331), .ZN(n1093) );
XOR2_X1 U1021 ( .A(n1122), .B(n1203), .Z(n1094) );
INV_X1 U1022 ( .A(n1121), .ZN(n1203) );
NAND2_X1 U1023 ( .A1(G210), .A2(n1331), .ZN(n1121) );
NAND2_X1 U1024 ( .A1(n1311), .A2(n1317), .ZN(n1331) );
INV_X1 U1025 ( .A(G237), .ZN(n1311) );
NAND3_X1 U1026 ( .A1(n1332), .A2(n1317), .A3(n1333), .ZN(n1122) );
XOR2_X1 U1027 ( .A(KEYINPUT43), .B(n1334), .Z(n1333) );
NOR2_X1 U1028 ( .A1(n1335), .A2(n1246), .ZN(n1334) );
NAND2_X1 U1029 ( .A1(n1335), .A2(n1246), .ZN(n1332) );
INV_X1 U1030 ( .A(n1254), .ZN(n1246) );
XNOR2_X1 U1031 ( .A(n1150), .B(n1151), .ZN(n1254) );
XOR2_X1 U1032 ( .A(n1336), .B(n1337), .Z(n1151) );
XOR2_X1 U1033 ( .A(G104), .B(G101), .Z(n1337) );
XOR2_X1 U1034 ( .A(n1338), .B(G107), .Z(n1336) );
XNOR2_X1 U1035 ( .A(KEYINPUT8), .B(KEYINPUT39), .ZN(n1338) );
XOR2_X1 U1036 ( .A(n1339), .B(n1340), .Z(n1150) );
NOR2_X1 U1037 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1038 ( .A(n1343), .B(KEYINPUT51), .Z(n1342) );
NAND2_X1 U1039 ( .A1(n1344), .A2(n1316), .ZN(n1343) );
NOR2_X1 U1040 ( .A1(n1316), .A2(n1344), .ZN(n1341) );
XOR2_X1 U1041 ( .A(KEYINPUT19), .B(n1345), .Z(n1344) );
XOR2_X1 U1042 ( .A(n1199), .B(G122), .Z(n1339) );
XNOR2_X1 U1043 ( .A(n1346), .B(n1347), .ZN(n1335) );
XOR2_X1 U1044 ( .A(G125), .B(n1256), .Z(n1347) );
NOR2_X1 U1045 ( .A1(n1145), .A2(G953), .ZN(n1256) );
INV_X1 U1046 ( .A(G224), .ZN(n1145) );
NAND2_X1 U1047 ( .A1(KEYINPUT63), .A2(n1258), .ZN(n1346) );
NAND2_X1 U1048 ( .A1(G221), .A2(n1348), .ZN(n1271) );
XOR2_X1 U1049 ( .A(n1118), .B(G469), .Z(n1084) );
AND2_X1 U1050 ( .A1(n1349), .A2(n1317), .ZN(n1118) );
NAND2_X1 U1051 ( .A1(n1350), .A2(n1351), .ZN(n1349) );
NAND3_X1 U1052 ( .A1(n1194), .A2(n1352), .A3(KEYINPUT6), .ZN(n1351) );
XOR2_X1 U1053 ( .A(n1353), .B(n1354), .Z(n1352) );
AND2_X1 U1054 ( .A1(n1195), .A2(KEYINPUT57), .ZN(n1353) );
NAND2_X1 U1055 ( .A1(n1355), .A2(n1356), .ZN(n1350) );
NAND2_X1 U1056 ( .A1(KEYINPUT6), .A2(n1194), .ZN(n1356) );
XOR2_X1 U1057 ( .A(n1357), .B(n1358), .Z(n1194) );
INV_X1 U1058 ( .A(n1135), .ZN(n1358) );
XOR2_X1 U1059 ( .A(n1359), .B(n1360), .Z(n1135) );
NOR2_X1 U1060 ( .A1(G143), .A2(KEYINPUT36), .ZN(n1360) );
XOR2_X1 U1061 ( .A(n1361), .B(G101), .Z(n1357) );
NAND3_X1 U1062 ( .A1(n1362), .A2(n1363), .A3(n1364), .ZN(n1361) );
OR2_X1 U1063 ( .A1(n1365), .A2(KEYINPUT41), .ZN(n1364) );
NAND3_X1 U1064 ( .A1(KEYINPUT41), .A2(n1365), .A3(G104), .ZN(n1363) );
NAND2_X1 U1065 ( .A1(n1366), .A2(n1167), .ZN(n1362) );
INV_X1 U1066 ( .A(G104), .ZN(n1167) );
NAND2_X1 U1067 ( .A1(n1367), .A2(KEYINPUT41), .ZN(n1366) );
XOR2_X1 U1068 ( .A(n1365), .B(KEYINPUT47), .Z(n1367) );
INV_X1 U1069 ( .A(G107), .ZN(n1365) );
XNOR2_X1 U1070 ( .A(n1368), .B(n1354), .ZN(n1355) );
XNOR2_X1 U1071 ( .A(n1369), .B(n1370), .ZN(n1354) );
XOR2_X1 U1072 ( .A(G140), .B(G110), .Z(n1370) );
NAND2_X1 U1073 ( .A1(KEYINPUT55), .A2(n1198), .ZN(n1369) );
NOR2_X1 U1074 ( .A1(n1138), .A2(G953), .ZN(n1198) );
INV_X1 U1075 ( .A(G227), .ZN(n1138) );
NAND2_X1 U1076 ( .A1(KEYINPUT57), .A2(n1371), .ZN(n1368) );
NOR2_X1 U1077 ( .A1(n1290), .A2(n1098), .ZN(n1089) );
XOR2_X1 U1078 ( .A(n1372), .B(n1159), .Z(n1098) );
AND2_X1 U1079 ( .A1(G217), .A2(n1348), .ZN(n1159) );
NAND2_X1 U1080 ( .A1(G234), .A2(n1317), .ZN(n1348) );
NAND2_X1 U1081 ( .A1(n1155), .A2(n1317), .ZN(n1372) );
XNOR2_X1 U1082 ( .A(n1373), .B(n1374), .ZN(n1155) );
XOR2_X1 U1083 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1084 ( .A(n1377), .B(G119), .Z(n1376) );
NAND2_X1 U1085 ( .A1(n1326), .A2(G221), .ZN(n1377) );
AND2_X1 U1086 ( .A1(G234), .A2(n1064), .ZN(n1326) );
XOR2_X1 U1087 ( .A(G137), .B(n1133), .Z(n1375) );
INV_X1 U1088 ( .A(G125), .ZN(n1133) );
XOR2_X1 U1089 ( .A(n1378), .B(n1308), .Z(n1373) );
XOR2_X1 U1090 ( .A(G140), .B(KEYINPUT26), .Z(n1308) );
XOR2_X1 U1091 ( .A(n1359), .B(n1379), .Z(n1378) );
NOR2_X1 U1092 ( .A1(KEYINPUT49), .A2(n1199), .ZN(n1379) );
INV_X1 U1093 ( .A(G110), .ZN(n1199) );
INV_X1 U1094 ( .A(n1292), .ZN(n1290) );
XOR2_X1 U1095 ( .A(n1111), .B(G472), .Z(n1292) );
NAND2_X1 U1096 ( .A1(n1380), .A2(n1317), .ZN(n1111) );
INV_X1 U1097 ( .A(G902), .ZN(n1317) );
XOR2_X1 U1098 ( .A(n1182), .B(n1381), .Z(n1380) );
XOR2_X1 U1099 ( .A(n1382), .B(n1383), .Z(n1381) );
NOR2_X1 U1100 ( .A1(KEYINPUT42), .A2(n1181), .ZN(n1383) );
XNOR2_X1 U1101 ( .A(n1345), .B(n1316), .ZN(n1181) );
INV_X1 U1102 ( .A(G113), .ZN(n1316) );
XNOR2_X1 U1103 ( .A(n1384), .B(n1385), .ZN(n1345) );
XOR2_X1 U1104 ( .A(KEYINPUT62), .B(G119), .Z(n1385) );
INV_X1 U1105 ( .A(G116), .ZN(n1384) );
NOR2_X1 U1106 ( .A1(n1177), .A2(n1176), .ZN(n1382) );
NOR2_X1 U1107 ( .A1(G101), .A2(n1386), .ZN(n1176) );
AND3_X1 U1108 ( .A1(n1387), .A2(n1064), .A3(G210), .ZN(n1386) );
AND4_X1 U1109 ( .A1(G210), .A2(G101), .A3(n1387), .A4(n1064), .ZN(n1177) );
INV_X1 U1110 ( .A(G953), .ZN(n1064) );
XOR2_X1 U1111 ( .A(G237), .B(KEYINPUT34), .Z(n1387) );
XOR2_X1 U1112 ( .A(n1258), .B(n1195), .Z(n1182) );
INV_X1 U1113 ( .A(n1371), .ZN(n1195) );
NAND2_X1 U1114 ( .A1(n1388), .A2(n1389), .ZN(n1371) );
OR2_X1 U1115 ( .A1(n1136), .A2(G134), .ZN(n1389) );
NAND2_X1 U1116 ( .A1(G134), .A2(n1390), .ZN(n1388) );
XNOR2_X1 U1117 ( .A(n1136), .B(KEYINPUT29), .ZN(n1390) );
XOR2_X1 U1118 ( .A(G137), .B(G131), .Z(n1136) );
XNOR2_X1 U1119 ( .A(n1359), .B(G143), .ZN(n1258) );
XNOR2_X1 U1120 ( .A(G146), .B(n1322), .ZN(n1359) );
XOR2_X1 U1121 ( .A(G128), .B(KEYINPUT16), .Z(n1322) );
endmodule


