//Key = 0110101010010100010000011100111010111011110101111000111110101111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341;

XNOR2_X1 U741 ( .A(G107), .B(n1026), .ZN(G9) );
NAND3_X1 U742 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
XNOR2_X1 U743 ( .A(n1030), .B(KEYINPUT35), .ZN(n1029) );
AND2_X1 U744 ( .A1(n1031), .A2(n1032), .ZN(G75) );
OR3_X1 U745 ( .A1(G952), .A2(G953), .A3(n1033), .ZN(n1032) );
NAND4_X1 U746 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1031) );
NOR4_X1 U747 ( .A1(KEYINPUT3), .A2(G953), .A3(n1033), .A4(n1038), .ZN(n1037) );
NOR3_X1 U748 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
INV_X1 U751 ( .A(n1046), .ZN(n1039) );
AND4_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1033) );
XOR2_X1 U753 ( .A(KEYINPUT26), .B(n1051), .Z(n1050) );
NOR3_X1 U754 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
XOR2_X1 U755 ( .A(n1055), .B(KEYINPUT11), .Z(n1054) );
NAND2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
XNOR2_X1 U757 ( .A(KEYINPUT27), .B(n1058), .ZN(n1056) );
XNOR2_X1 U758 ( .A(n1059), .B(n1060), .ZN(n1053) );
NAND2_X1 U759 ( .A1(KEYINPUT28), .A2(n1061), .ZN(n1059) );
NAND3_X1 U760 ( .A1(n1062), .A2(n1045), .A3(n1063), .ZN(n1052) );
NAND2_X1 U761 ( .A1(G469), .A2(n1058), .ZN(n1063) );
NOR2_X1 U762 ( .A1(n1064), .A2(n1065), .ZN(n1049) );
NAND3_X1 U763 ( .A1(n1066), .A2(n1045), .A3(n1067), .ZN(n1035) );
NAND2_X1 U764 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND2_X1 U765 ( .A1(n1046), .A2(n1070), .ZN(n1069) );
NAND2_X1 U766 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR3_X1 U767 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1046) );
NAND3_X1 U768 ( .A1(n1076), .A2(n1077), .A3(n1048), .ZN(n1068) );
NAND2_X1 U769 ( .A1(n1078), .A2(n1075), .ZN(n1077) );
NAND2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
INV_X1 U771 ( .A(KEYINPUT46), .ZN(n1080) );
NAND4_X1 U772 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1076) );
INV_X1 U773 ( .A(n1075), .ZN(n1084) );
NAND2_X1 U774 ( .A1(n1030), .A2(n1085), .ZN(n1083) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U777 ( .A1(n1047), .A2(n1090), .ZN(n1089) );
NAND2_X1 U778 ( .A1(KEYINPUT46), .A2(n1079), .ZN(n1081) );
NOR3_X1 U779 ( .A1(n1074), .A2(n1091), .A3(n1062), .ZN(n1079) );
XOR2_X1 U780 ( .A(n1092), .B(n1093), .Z(G72) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR3_X1 U782 ( .A1(n1096), .A2(KEYINPUT12), .A3(n1097), .ZN(n1095) );
XOR2_X1 U783 ( .A(n1098), .B(n1099), .Z(n1096) );
XOR2_X1 U784 ( .A(n1100), .B(n1101), .Z(n1099) );
XNOR2_X1 U785 ( .A(n1102), .B(n1103), .ZN(n1101) );
NAND2_X1 U786 ( .A1(KEYINPUT32), .A2(n1104), .ZN(n1102) );
INV_X1 U787 ( .A(G125), .ZN(n1104) );
NAND2_X1 U788 ( .A1(KEYINPUT48), .A2(n1105), .ZN(n1100) );
XOR2_X1 U789 ( .A(n1106), .B(n1107), .Z(n1098) );
NAND2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1094) );
XNOR2_X1 U791 ( .A(KEYINPUT1), .B(n1110), .ZN(n1108) );
NAND2_X1 U792 ( .A1(n1111), .A2(n1112), .ZN(n1092) );
NAND2_X1 U793 ( .A1(G900), .A2(G227), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(G69) );
NAND4_X1 U795 ( .A1(n1111), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1114) );
XOR2_X1 U796 ( .A(n1118), .B(KEYINPUT15), .Z(n1113) );
NAND2_X1 U797 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1115), .ZN(n1120) );
NAND2_X1 U799 ( .A1(G898), .A2(G224), .ZN(n1115) );
XNOR2_X1 U800 ( .A(n1110), .B(KEYINPUT42), .ZN(n1111) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1119) );
NAND3_X1 U802 ( .A1(n1121), .A2(n1122), .A3(n1034), .ZN(n1117) );
NAND2_X1 U803 ( .A1(G953), .A2(n1123), .ZN(n1122) );
OR3_X1 U804 ( .A1(n1034), .A2(G953), .A3(n1121), .ZN(n1116) );
NOR2_X1 U805 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XOR2_X1 U806 ( .A(n1126), .B(n1127), .Z(n1125) );
XOR2_X1 U807 ( .A(KEYINPUT17), .B(n1128), .Z(n1127) );
NOR2_X1 U808 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U809 ( .A1(n1124), .A2(n1131), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1132), .B(n1133), .ZN(n1131) );
XOR2_X1 U811 ( .A(KEYINPUT16), .B(n1134), .Z(n1133) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1130), .ZN(n1134) );
NOR2_X1 U813 ( .A1(n1124), .A2(n1136), .ZN(G60) );
XNOR2_X1 U814 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1139), .A2(n1130), .ZN(n1138) );
XNOR2_X1 U816 ( .A(G104), .B(n1140), .ZN(G6) );
NOR2_X1 U817 ( .A1(n1124), .A2(n1141), .ZN(G57) );
XOR2_X1 U818 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U819 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1142) );
NOR2_X1 U821 ( .A1(n1148), .A2(n1130), .ZN(n1147) );
NAND2_X1 U822 ( .A1(KEYINPUT40), .A2(n1149), .ZN(n1146) );
NOR2_X1 U823 ( .A1(n1124), .A2(n1150), .ZN(G54) );
XOR2_X1 U824 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND3_X1 U825 ( .A1(G469), .A2(n1153), .A3(n1154), .ZN(n1152) );
XOR2_X1 U826 ( .A(n1155), .B(KEYINPUT37), .Z(n1154) );
NAND2_X1 U827 ( .A1(n1156), .A2(n1157), .ZN(n1151) );
NAND2_X1 U828 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U829 ( .A(KEYINPUT58), .B(n1160), .Z(n1156) );
NOR2_X1 U830 ( .A1(n1158), .A2(n1159), .ZN(n1160) );
XNOR2_X1 U831 ( .A(n1161), .B(n1162), .ZN(n1159) );
XNOR2_X1 U832 ( .A(KEYINPUT53), .B(n1163), .ZN(n1162) );
XNOR2_X1 U833 ( .A(n1164), .B(n1165), .ZN(n1161) );
NAND2_X1 U834 ( .A1(n1166), .A2(n1103), .ZN(n1164) );
INV_X1 U835 ( .A(G140), .ZN(n1103) );
XNOR2_X1 U836 ( .A(KEYINPUT45), .B(KEYINPUT2), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1167), .B(n1168), .Z(n1158) );
XOR2_X1 U838 ( .A(n1169), .B(n1106), .Z(n1168) );
XNOR2_X1 U839 ( .A(KEYINPUT30), .B(n1170), .ZN(n1167) );
NOR2_X1 U840 ( .A1(KEYINPUT19), .A2(n1171), .ZN(n1170) );
XNOR2_X1 U841 ( .A(n1172), .B(n1173), .ZN(n1171) );
NOR2_X1 U842 ( .A1(n1124), .A2(n1174), .ZN(G51) );
XOR2_X1 U843 ( .A(n1121), .B(n1175), .Z(n1174) );
XOR2_X1 U844 ( .A(n1176), .B(n1177), .Z(n1175) );
NOR3_X1 U845 ( .A1(n1178), .A2(n1061), .A3(n1130), .ZN(n1177) );
NAND2_X1 U846 ( .A1(n1155), .A2(n1153), .ZN(n1130) );
NAND2_X1 U847 ( .A1(n1036), .A2(n1034), .ZN(n1153) );
AND4_X1 U848 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1034) );
NOR4_X1 U849 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1182) );
INV_X1 U850 ( .A(n1140), .ZN(n1186) );
NAND3_X1 U851 ( .A1(n1027), .A2(n1030), .A3(n1187), .ZN(n1140) );
INV_X1 U852 ( .A(n1188), .ZN(n1183) );
NOR2_X1 U853 ( .A1(n1189), .A2(n1190), .ZN(n1181) );
AND3_X1 U854 ( .A1(n1027), .A2(n1030), .A3(n1028), .ZN(n1190) );
NOR4_X1 U855 ( .A1(n1191), .A2(n1192), .A3(n1041), .A4(n1088), .ZN(n1189) );
INV_X1 U856 ( .A(n1048), .ZN(n1041) );
NOR2_X1 U857 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U858 ( .A(KEYINPUT18), .ZN(n1194) );
NOR3_X1 U859 ( .A1(n1195), .A2(n1196), .A3(n1085), .ZN(n1193) );
NOR2_X1 U860 ( .A1(KEYINPUT18), .A2(n1027), .ZN(n1191) );
INV_X1 U861 ( .A(n1109), .ZN(n1036) );
NAND4_X1 U862 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1109) );
AND4_X1 U863 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
OR2_X1 U864 ( .A1(n1205), .A2(n1073), .ZN(n1204) );
XOR2_X1 U865 ( .A(n1206), .B(KEYINPUT57), .Z(n1205) );
NAND4_X1 U866 ( .A1(n1028), .A2(n1043), .A3(n1207), .A4(n1208), .ZN(n1206) );
XNOR2_X1 U867 ( .A(KEYINPUT20), .B(n1088), .ZN(n1207) );
NOR2_X1 U868 ( .A1(n1209), .A2(n1210), .ZN(n1199) );
INV_X1 U869 ( .A(n1211), .ZN(n1209) );
NAND4_X1 U870 ( .A1(n1043), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1198) );
NOR3_X1 U871 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1214) );
XNOR2_X1 U872 ( .A(n1085), .B(KEYINPUT50), .ZN(n1215) );
XNOR2_X1 U873 ( .A(KEYINPUT6), .B(n1208), .ZN(n1212) );
INV_X1 U874 ( .A(n1218), .ZN(n1197) );
XNOR2_X1 U875 ( .A(G902), .B(KEYINPUT41), .ZN(n1155) );
XOR2_X1 U876 ( .A(KEYINPUT22), .B(KEYINPUT21), .Z(n1178) );
NOR3_X1 U877 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1176) );
NOR2_X1 U878 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
AND3_X1 U879 ( .A1(n1222), .A2(n1223), .A3(KEYINPUT34), .ZN(n1220) );
AND2_X1 U880 ( .A1(KEYINPUT55), .A2(n1224), .ZN(n1223) );
NOR2_X1 U881 ( .A1(KEYINPUT34), .A2(n1224), .ZN(n1219) );
AND2_X1 U882 ( .A1(n1225), .A2(n1226), .ZN(n1224) );
NAND2_X1 U883 ( .A1(KEYINPUT62), .A2(n1227), .ZN(n1226) );
NAND3_X1 U884 ( .A1(G125), .A2(n1228), .A3(n1229), .ZN(n1225) );
INV_X1 U885 ( .A(KEYINPUT62), .ZN(n1229) );
NOR2_X1 U886 ( .A1(n1110), .A2(G952), .ZN(n1124) );
XNOR2_X1 U887 ( .A(n1230), .B(n1210), .ZN(G48) );
AND3_X1 U888 ( .A1(n1231), .A2(n1085), .A3(n1187), .ZN(n1210) );
XOR2_X1 U889 ( .A(n1232), .B(n1233), .Z(G45) );
NAND2_X1 U890 ( .A1(KEYINPUT43), .A2(G143), .ZN(n1233) );
OR4_X1 U891 ( .A1(n1234), .A2(n1235), .A3(n1217), .A4(n1216), .ZN(n1232) );
INV_X1 U892 ( .A(n1236), .ZN(n1217) );
XNOR2_X1 U893 ( .A(G140), .B(n1203), .ZN(G42) );
NAND3_X1 U894 ( .A1(n1086), .A2(n1043), .A3(n1237), .ZN(n1203) );
XNOR2_X1 U895 ( .A(G137), .B(n1211), .ZN(G39) );
NAND3_X1 U896 ( .A1(n1086), .A2(n1048), .A3(n1231), .ZN(n1211) );
XOR2_X1 U897 ( .A(G134), .B(n1238), .Z(G36) );
NOR3_X1 U898 ( .A1(n1234), .A2(n1072), .A3(n1073), .ZN(n1238) );
NAND2_X1 U899 ( .A1(n1239), .A2(n1240), .ZN(G33) );
NAND2_X1 U900 ( .A1(G131), .A2(n1202), .ZN(n1240) );
INV_X1 U901 ( .A(n1241), .ZN(n1202) );
XOR2_X1 U902 ( .A(n1242), .B(KEYINPUT9), .Z(n1239) );
NAND2_X1 U903 ( .A1(n1241), .A2(n1105), .ZN(n1242) );
NOR3_X1 U904 ( .A1(n1071), .A2(n1073), .A3(n1234), .ZN(n1241) );
NAND3_X1 U905 ( .A1(n1043), .A2(n1208), .A3(n1213), .ZN(n1234) );
INV_X1 U906 ( .A(n1086), .ZN(n1073) );
NOR2_X1 U907 ( .A1(n1091), .A2(n1243), .ZN(n1086) );
INV_X1 U908 ( .A(n1062), .ZN(n1243) );
XOR2_X1 U909 ( .A(n1244), .B(G128), .Z(G30) );
NAND2_X1 U910 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NAND3_X1 U911 ( .A1(n1085), .A2(n1247), .A3(n1248), .ZN(n1246) );
INV_X1 U912 ( .A(KEYINPUT23), .ZN(n1248) );
NAND2_X1 U913 ( .A1(n1218), .A2(KEYINPUT23), .ZN(n1245) );
NOR2_X1 U914 ( .A1(n1247), .A2(n1235), .ZN(n1218) );
NAND2_X1 U915 ( .A1(n1231), .A2(n1028), .ZN(n1247) );
AND4_X1 U916 ( .A1(n1043), .A2(n1249), .A3(n1208), .A4(n1090), .ZN(n1231) );
XOR2_X1 U917 ( .A(n1250), .B(n1251), .Z(G3) );
NOR2_X1 U918 ( .A1(G101), .A2(KEYINPUT0), .ZN(n1251) );
NAND4_X1 U919 ( .A1(n1252), .A2(n1213), .A3(n1253), .A4(n1048), .ZN(n1250) );
NOR2_X1 U920 ( .A1(n1196), .A2(n1235), .ZN(n1253) );
XNOR2_X1 U921 ( .A(n1043), .B(KEYINPUT8), .ZN(n1252) );
INV_X1 U922 ( .A(n1195), .ZN(n1043) );
XNOR2_X1 U923 ( .A(G125), .B(n1201), .ZN(G27) );
NAND4_X1 U924 ( .A1(n1237), .A2(n1085), .A3(n1067), .A4(n1045), .ZN(n1201) );
AND4_X1 U925 ( .A1(n1047), .A2(n1187), .A3(n1208), .A4(n1090), .ZN(n1237) );
NAND2_X1 U926 ( .A1(n1075), .A2(n1254), .ZN(n1208) );
NAND3_X1 U927 ( .A1(G902), .A2(n1255), .A3(n1097), .ZN(n1254) );
NOR2_X1 U928 ( .A1(n1110), .A2(G900), .ZN(n1097) );
XNOR2_X1 U929 ( .A(G122), .B(n1179), .ZN(G24) );
NAND4_X1 U930 ( .A1(n1256), .A2(n1030), .A3(n1236), .A4(n1257), .ZN(n1179) );
INV_X1 U931 ( .A(n1074), .ZN(n1030) );
NAND2_X1 U932 ( .A1(n1258), .A2(n1047), .ZN(n1074) );
XNOR2_X1 U933 ( .A(G119), .B(n1180), .ZN(G21) );
NAND4_X1 U934 ( .A1(n1256), .A2(n1048), .A3(n1249), .A4(n1090), .ZN(n1180) );
XNOR2_X1 U935 ( .A(n1259), .B(n1185), .ZN(G18) );
AND3_X1 U936 ( .A1(n1213), .A2(n1028), .A3(n1256), .ZN(n1185) );
INV_X1 U937 ( .A(n1072), .ZN(n1028) );
NAND2_X1 U938 ( .A1(n1260), .A2(n1257), .ZN(n1072) );
XNOR2_X1 U939 ( .A(n1236), .B(KEYINPUT44), .ZN(n1260) );
XOR2_X1 U940 ( .A(G113), .B(n1184), .Z(G15) );
AND3_X1 U941 ( .A1(n1213), .A2(n1187), .A3(n1256), .ZN(n1184) );
AND4_X1 U942 ( .A1(n1085), .A2(n1067), .A3(n1261), .A4(n1045), .ZN(n1256) );
INV_X1 U943 ( .A(n1235), .ZN(n1085) );
INV_X1 U944 ( .A(n1071), .ZN(n1187) );
NAND2_X1 U945 ( .A1(n1262), .A2(n1236), .ZN(n1071) );
XNOR2_X1 U946 ( .A(KEYINPUT47), .B(n1216), .ZN(n1262) );
INV_X1 U947 ( .A(n1257), .ZN(n1216) );
INV_X1 U948 ( .A(n1088), .ZN(n1213) );
NAND2_X1 U949 ( .A1(n1258), .A2(n1249), .ZN(n1088) );
XNOR2_X1 U950 ( .A(n1047), .B(KEYINPUT14), .ZN(n1249) );
XNOR2_X1 U951 ( .A(G110), .B(n1188), .ZN(G12) );
NAND4_X1 U952 ( .A1(n1048), .A2(n1027), .A3(n1047), .A4(n1090), .ZN(n1188) );
INV_X1 U953 ( .A(n1258), .ZN(n1090) );
NOR2_X1 U954 ( .A1(n1263), .A2(n1065), .ZN(n1258) );
NOR2_X1 U955 ( .A1(n1129), .A2(n1264), .ZN(n1065) );
AND2_X1 U956 ( .A1(n1126), .A2(n1265), .ZN(n1264) );
XOR2_X1 U957 ( .A(n1064), .B(KEYINPUT5), .Z(n1263) );
AND3_X1 U958 ( .A1(n1129), .A2(n1265), .A3(n1126), .ZN(n1064) );
XOR2_X1 U959 ( .A(n1266), .B(n1267), .Z(n1126) );
XOR2_X1 U960 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U961 ( .A(G128), .B(n1163), .ZN(n1269) );
XNOR2_X1 U962 ( .A(KEYINPUT33), .B(n1270), .ZN(n1268) );
INV_X1 U963 ( .A(G137), .ZN(n1270) );
XOR2_X1 U964 ( .A(n1271), .B(n1272), .Z(n1266) );
XOR2_X1 U965 ( .A(n1273), .B(n1274), .Z(n1271) );
NAND2_X1 U966 ( .A1(n1275), .A2(G221), .ZN(n1273) );
NAND2_X1 U967 ( .A1(G217), .A2(n1276), .ZN(n1129) );
XNOR2_X1 U968 ( .A(n1277), .B(n1148), .ZN(n1047) );
INV_X1 U969 ( .A(G472), .ZN(n1148) );
NAND2_X1 U970 ( .A1(n1278), .A2(n1265), .ZN(n1277) );
XOR2_X1 U971 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U972 ( .A(n1145), .B(n1149), .Z(n1280) );
XNOR2_X1 U973 ( .A(n1281), .B(n1274), .ZN(n1149) );
XNOR2_X1 U974 ( .A(G116), .B(n1282), .ZN(n1281) );
XNOR2_X1 U975 ( .A(n1228), .B(n1283), .ZN(n1145) );
AND2_X1 U976 ( .A1(G210), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U977 ( .A(G101), .B(n1285), .ZN(n1279) );
NOR2_X1 U978 ( .A1(KEYINPUT10), .A2(n1169), .ZN(n1285) );
NOR3_X1 U979 ( .A1(n1235), .A2(n1196), .A3(n1195), .ZN(n1027) );
NAND2_X1 U980 ( .A1(n1044), .A2(n1045), .ZN(n1195) );
NAND2_X1 U981 ( .A1(G221), .A2(n1276), .ZN(n1045) );
NAND2_X1 U982 ( .A1(G234), .A2(n1265), .ZN(n1276) );
INV_X1 U983 ( .A(n1067), .ZN(n1044) );
XNOR2_X1 U984 ( .A(n1058), .B(n1286), .ZN(n1067) );
XNOR2_X1 U985 ( .A(KEYINPUT54), .B(n1057), .ZN(n1286) );
INV_X1 U986 ( .A(G469), .ZN(n1057) );
NAND2_X1 U987 ( .A1(n1287), .A2(n1265), .ZN(n1058) );
XOR2_X1 U988 ( .A(n1288), .B(n1289), .Z(n1287) );
XNOR2_X1 U989 ( .A(n1290), .B(n1291), .ZN(n1289) );
NOR2_X1 U990 ( .A1(KEYINPUT49), .A2(n1292), .ZN(n1291) );
XNOR2_X1 U991 ( .A(G110), .B(G140), .ZN(n1292) );
NAND2_X1 U992 ( .A1(n1293), .A2(KEYINPUT61), .ZN(n1290) );
XOR2_X1 U993 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U994 ( .A(n1172), .B(n1106), .Z(n1295) );
XOR2_X1 U995 ( .A(n1296), .B(n1297), .Z(n1106) );
NAND2_X1 U996 ( .A1(KEYINPUT63), .A2(n1230), .ZN(n1296) );
XNOR2_X1 U997 ( .A(G104), .B(n1298), .ZN(n1172) );
XOR2_X1 U998 ( .A(KEYINPUT38), .B(G107), .Z(n1298) );
XOR2_X1 U999 ( .A(n1144), .B(KEYINPUT7), .Z(n1294) );
XNOR2_X1 U1000 ( .A(n1169), .B(n1173), .ZN(n1144) );
INV_X1 U1001 ( .A(G101), .ZN(n1173) );
XOR2_X1 U1002 ( .A(n1299), .B(n1107), .Z(n1169) );
XOR2_X1 U1003 ( .A(G134), .B(G137), .Z(n1107) );
NAND2_X1 U1004 ( .A1(KEYINPUT13), .A2(n1105), .ZN(n1299) );
XOR2_X1 U1005 ( .A(n1165), .B(KEYINPUT4), .Z(n1288) );
NAND2_X1 U1006 ( .A1(G227), .A2(n1110), .ZN(n1165) );
INV_X1 U1007 ( .A(n1261), .ZN(n1196) );
NAND2_X1 U1008 ( .A1(n1075), .A2(n1300), .ZN(n1261) );
NAND4_X1 U1009 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1123), .ZN(n1300) );
INV_X1 U1010 ( .A(G898), .ZN(n1123) );
NAND3_X1 U1011 ( .A1(n1255), .A2(n1110), .A3(G952), .ZN(n1075) );
NAND2_X1 U1012 ( .A1(G237), .A2(G234), .ZN(n1255) );
NAND2_X1 U1013 ( .A1(n1301), .A2(n1062), .ZN(n1235) );
NAND2_X1 U1014 ( .A1(G214), .A2(n1302), .ZN(n1062) );
XOR2_X1 U1015 ( .A(n1091), .B(KEYINPUT31), .Z(n1301) );
XNOR2_X1 U1016 ( .A(n1303), .B(n1061), .ZN(n1091) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1302), .ZN(n1061) );
NAND2_X1 U1018 ( .A1(n1304), .A2(n1265), .ZN(n1302) );
INV_X1 U1019 ( .A(G237), .ZN(n1304) );
XOR2_X1 U1020 ( .A(n1060), .B(KEYINPUT24), .Z(n1303) );
NAND2_X1 U1021 ( .A1(n1305), .A2(n1265), .ZN(n1060) );
XNOR2_X1 U1022 ( .A(n1227), .B(n1306), .ZN(n1305) );
XOR2_X1 U1023 ( .A(n1222), .B(n1307), .Z(n1306) );
NOR2_X1 U1024 ( .A1(KEYINPUT51), .A2(n1121), .ZN(n1307) );
XNOR2_X1 U1025 ( .A(n1308), .B(n1309), .ZN(n1121) );
XOR2_X1 U1026 ( .A(G107), .B(n1310), .Z(n1309) );
XNOR2_X1 U1027 ( .A(G122), .B(n1163), .ZN(n1310) );
INV_X1 U1028 ( .A(G110), .ZN(n1163) );
XOR2_X1 U1029 ( .A(n1311), .B(n1312), .Z(n1308) );
XNOR2_X1 U1030 ( .A(G101), .B(n1313), .ZN(n1312) );
NAND3_X1 U1031 ( .A1(n1314), .A2(n1315), .A3(n1316), .ZN(n1313) );
NAND2_X1 U1032 ( .A1(KEYINPUT59), .A2(n1317), .ZN(n1316) );
NAND3_X1 U1033 ( .A1(n1318), .A2(n1319), .A3(n1282), .ZN(n1315) );
INV_X1 U1034 ( .A(KEYINPUT59), .ZN(n1319) );
OR2_X1 U1035 ( .A1(n1282), .A2(n1318), .ZN(n1314) );
NOR2_X1 U1036 ( .A1(n1320), .A2(n1317), .ZN(n1318) );
XOR2_X1 U1037 ( .A(n1321), .B(n1259), .Z(n1317) );
NAND2_X1 U1038 ( .A1(KEYINPUT36), .A2(n1274), .ZN(n1321) );
XOR2_X1 U1039 ( .A(G119), .B(KEYINPUT39), .Z(n1274) );
INV_X1 U1040 ( .A(KEYINPUT25), .ZN(n1320) );
XOR2_X1 U1041 ( .A(G113), .B(KEYINPUT29), .Z(n1282) );
NAND2_X1 U1042 ( .A1(KEYINPUT60), .A2(G104), .ZN(n1311) );
AND2_X1 U1043 ( .A1(G224), .A2(n1110), .ZN(n1222) );
XOR2_X1 U1044 ( .A(n1228), .B(G125), .Z(n1227) );
XNOR2_X1 U1045 ( .A(G146), .B(n1297), .ZN(n1228) );
XOR2_X1 U1046 ( .A(G128), .B(G143), .Z(n1297) );
NOR2_X1 U1047 ( .A1(n1257), .A2(n1236), .ZN(n1048) );
XOR2_X1 U1048 ( .A(n1322), .B(n1139), .Z(n1236) );
INV_X1 U1049 ( .A(G475), .ZN(n1139) );
NAND2_X1 U1050 ( .A1(n1137), .A2(n1265), .ZN(n1322) );
XNOR2_X1 U1051 ( .A(n1323), .B(n1324), .ZN(n1137) );
XOR2_X1 U1052 ( .A(G113), .B(n1325), .Z(n1324) );
XOR2_X1 U1053 ( .A(KEYINPUT52), .B(G122), .Z(n1325) );
XNOR2_X1 U1054 ( .A(n1272), .B(n1326), .ZN(n1323) );
XNOR2_X1 U1055 ( .A(n1327), .B(n1328), .ZN(n1326) );
NOR2_X1 U1056 ( .A1(n1329), .A2(n1330), .ZN(n1328) );
XOR2_X1 U1057 ( .A(n1331), .B(KEYINPUT56), .Z(n1330) );
NAND2_X1 U1058 ( .A1(n1332), .A2(n1105), .ZN(n1331) );
NOR2_X1 U1059 ( .A1(n1332), .A2(n1105), .ZN(n1329) );
INV_X1 U1060 ( .A(G131), .ZN(n1105) );
XNOR2_X1 U1061 ( .A(n1333), .B(G143), .ZN(n1332) );
NAND2_X1 U1062 ( .A1(n1284), .A2(G214), .ZN(n1333) );
NOR2_X1 U1063 ( .A1(G953), .A2(G237), .ZN(n1284) );
INV_X1 U1064 ( .A(G104), .ZN(n1327) );
XOR2_X1 U1065 ( .A(G125), .B(n1334), .Z(n1272) );
XNOR2_X1 U1066 ( .A(n1230), .B(G140), .ZN(n1334) );
INV_X1 U1067 ( .A(G146), .ZN(n1230) );
XOR2_X1 U1068 ( .A(n1335), .B(n1135), .Z(n1257) );
INV_X1 U1069 ( .A(G478), .ZN(n1135) );
NAND2_X1 U1070 ( .A1(n1132), .A2(n1265), .ZN(n1335) );
INV_X1 U1071 ( .A(G902), .ZN(n1265) );
XNOR2_X1 U1072 ( .A(n1336), .B(n1337), .ZN(n1132) );
XOR2_X1 U1073 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1074 ( .A(G128), .B(G122), .Z(n1339) );
XOR2_X1 U1075 ( .A(G143), .B(G134), .Z(n1338) );
XOR2_X1 U1076 ( .A(n1340), .B(n1341), .Z(n1336) );
XNOR2_X1 U1077 ( .A(n1259), .B(G107), .ZN(n1341) );
INV_X1 U1078 ( .A(G116), .ZN(n1259) );
NAND2_X1 U1079 ( .A1(G217), .A2(n1275), .ZN(n1340) );
AND2_X1 U1080 ( .A1(G234), .A2(n1110), .ZN(n1275) );
INV_X1 U1081 ( .A(G953), .ZN(n1110) );
endmodule


