//Key = 0001100011110101100000101101011100011100001010010111101111110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318;

NAND2_X1 U737 ( .A1(n1018), .A2(n1019), .ZN(G9) );
NAND2_X1 U738 ( .A1(G107), .A2(n1020), .ZN(n1019) );
XOR2_X1 U739 ( .A(KEYINPUT24), .B(n1021), .Z(n1018) );
NOR2_X1 U740 ( .A1(G107), .A2(n1020), .ZN(n1021) );
NOR2_X1 U741 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U742 ( .A1(n1024), .A2(n1025), .A3(G953), .A4(n1026), .ZN(n1023) );
NAND3_X1 U743 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1024) );
XOR2_X1 U744 ( .A(n1030), .B(KEYINPUT22), .Z(n1029) );
NAND2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND4_X1 U746 ( .A1(n1033), .A2(n1034), .A3(n1035), .A4(n1036), .ZN(n1032) );
NAND2_X1 U747 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1035) );
NAND2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND3_X1 U750 ( .A1(n1043), .A2(n1044), .A3(n1033), .ZN(n1031) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND3_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1046) );
NAND2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1045) );
NAND3_X1 U754 ( .A1(n1052), .A2(n1040), .A3(n1033), .ZN(n1028) );
NAND3_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1052) );
XOR2_X1 U756 ( .A(KEYINPUT47), .B(n1056), .Z(n1055) );
AND3_X1 U757 ( .A1(n1049), .A2(n1057), .A3(n1058), .ZN(n1056) );
NAND4_X1 U758 ( .A1(n1050), .A2(n1059), .A3(n1057), .A4(n1060), .ZN(n1054) );
INV_X1 U759 ( .A(n1061), .ZN(n1050) );
NAND3_X1 U760 ( .A1(n1062), .A2(n1063), .A3(n1034), .ZN(n1053) );
NAND3_X1 U761 ( .A1(n1034), .A2(n1043), .A3(n1064), .ZN(n1027) );
AND2_X1 U762 ( .A1(n1049), .A2(n1060), .ZN(n1034) );
NOR2_X1 U763 ( .A1(n1061), .A2(n1065), .ZN(n1049) );
NOR3_X1 U764 ( .A1(n1026), .A2(G953), .A3(G952), .ZN(n1022) );
AND4_X1 U765 ( .A1(n1066), .A2(n1043), .A3(n1067), .A4(n1068), .ZN(n1026) );
NOR4_X1 U766 ( .A1(n1069), .A2(n1070), .A3(n1071), .A4(n1048), .ZN(n1068) );
NOR2_X1 U767 ( .A1(n1072), .A2(n1073), .ZN(n1070) );
XOR2_X1 U768 ( .A(n1074), .B(n1075), .Z(n1067) );
XOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT1), .Z(n1075) );
XNOR2_X1 U770 ( .A(G472), .B(n1076), .ZN(n1074) );
NOR2_X1 U771 ( .A1(n1077), .A2(KEYINPUT40), .ZN(n1076) );
XOR2_X1 U772 ( .A(n1078), .B(n1079), .Z(n1066) );
XOR2_X1 U773 ( .A(KEYINPUT44), .B(n1080), .Z(n1079) );
NOR2_X1 U774 ( .A1(KEYINPUT62), .A2(n1081), .ZN(n1080) );
INV_X1 U775 ( .A(n1082), .ZN(n1081) );
XOR2_X1 U776 ( .A(n1083), .B(n1084), .Z(G72) );
XOR2_X1 U777 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NAND2_X1 U779 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XNOR2_X1 U780 ( .A(KEYINPUT54), .B(n1091), .ZN(n1090) );
NAND2_X1 U781 ( .A1(n1092), .A2(n1093), .ZN(n1085) );
NAND2_X1 U782 ( .A1(G953), .A2(n1094), .ZN(n1093) );
XOR2_X1 U783 ( .A(n1095), .B(n1096), .Z(n1092) );
XOR2_X1 U784 ( .A(n1097), .B(n1098), .Z(n1096) );
XNOR2_X1 U785 ( .A(n1099), .B(G131), .ZN(n1098) );
XOR2_X1 U786 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n1097) );
XNOR2_X1 U787 ( .A(n1100), .B(n1101), .ZN(n1095) );
XNOR2_X1 U788 ( .A(n1102), .B(n1103), .ZN(n1101) );
NOR3_X1 U789 ( .A1(n1087), .A2(KEYINPUT19), .A3(n1104), .ZN(n1083) );
AND2_X1 U790 ( .A1(G227), .A2(G900), .ZN(n1104) );
XOR2_X1 U791 ( .A(n1105), .B(n1106), .Z(G69) );
XOR2_X1 U792 ( .A(n1107), .B(n1108), .Z(n1106) );
OR2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U794 ( .A1(G953), .A2(n1111), .ZN(n1107) );
NAND2_X1 U795 ( .A1(G898), .A2(G224), .ZN(n1111) );
NOR2_X1 U796 ( .A1(n1112), .A2(G953), .ZN(n1105) );
NOR3_X1 U797 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(G66) );
NOR4_X1 U798 ( .A1(n1116), .A2(n1117), .A3(KEYINPUT7), .A4(n1118), .ZN(n1115) );
INV_X1 U799 ( .A(n1119), .ZN(n1116) );
NOR2_X1 U800 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
NOR3_X1 U801 ( .A1(n1117), .A2(n1121), .A3(n1118), .ZN(n1120) );
AND2_X1 U802 ( .A1(n1122), .A2(KEYINPUT7), .ZN(n1121) );
NOR2_X1 U803 ( .A1(KEYINPUT32), .A2(n1122), .ZN(n1119) );
NOR2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(G63) );
XOR2_X1 U805 ( .A(n1125), .B(n1126), .Z(n1124) );
NOR2_X1 U806 ( .A1(n1073), .A2(n1117), .ZN(n1125) );
INV_X1 U807 ( .A(G478), .ZN(n1073) );
NOR2_X1 U808 ( .A1(G952), .A2(n1127), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1128), .B(KEYINPUT6), .Z(n1127) );
NOR2_X1 U810 ( .A1(n1113), .A2(n1129), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1130), .B(n1131), .ZN(n1129) );
AND2_X1 U812 ( .A1(G475), .A2(n1132), .ZN(n1131) );
XNOR2_X1 U813 ( .A(G104), .B(n1133), .ZN(G6) );
NAND2_X1 U814 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
XNOR2_X1 U815 ( .A(KEYINPUT57), .B(n1136), .ZN(n1135) );
NOR2_X1 U816 ( .A1(n1113), .A2(n1137), .ZN(G57) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U818 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U819 ( .A(n1142), .B(n1143), .ZN(n1141) );
NAND2_X1 U820 ( .A1(KEYINPUT58), .A2(n1144), .ZN(n1142) );
XOR2_X1 U821 ( .A(n1145), .B(n1146), .Z(n1138) );
XNOR2_X1 U822 ( .A(KEYINPUT53), .B(n1147), .ZN(n1146) );
XNOR2_X1 U823 ( .A(n1148), .B(n1149), .ZN(n1145) );
NAND3_X1 U824 ( .A1(n1132), .A2(G472), .A3(KEYINPUT3), .ZN(n1148) );
NOR2_X1 U825 ( .A1(n1113), .A2(n1150), .ZN(G54) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U827 ( .A(n1153), .B(n1154), .ZN(n1152) );
AND2_X1 U828 ( .A1(G469), .A2(n1132), .ZN(n1154) );
INV_X1 U829 ( .A(n1117), .ZN(n1132) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1151) );
XNOR2_X1 U831 ( .A(KEYINPUT9), .B(n1157), .ZN(n1156) );
NAND2_X1 U832 ( .A1(KEYINPUT8), .A2(n1140), .ZN(n1155) );
NOR2_X1 U833 ( .A1(n1113), .A2(n1158), .ZN(G51) );
NOR2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1161), .B(n1162), .Z(n1160) );
NOR2_X1 U836 ( .A1(KEYINPUT14), .A2(n1163), .ZN(n1162) );
NOR2_X1 U837 ( .A1(n1082), .A2(n1117), .ZN(n1161) );
NAND2_X1 U838 ( .A1(G902), .A2(n1025), .ZN(n1117) );
NAND3_X1 U839 ( .A1(n1089), .A2(n1091), .A3(n1112), .ZN(n1025) );
AND4_X1 U840 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1112) );
AND4_X1 U841 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NOR2_X1 U842 ( .A1(n1172), .A2(n1173), .ZN(n1166) );
INV_X1 U843 ( .A(n1020), .ZN(n1172) );
NAND3_X1 U844 ( .A1(n1051), .A2(n1136), .A3(n1174), .ZN(n1020) );
AND3_X1 U845 ( .A1(n1175), .A2(n1176), .A3(n1060), .ZN(n1051) );
NAND2_X1 U846 ( .A1(n1134), .A2(n1136), .ZN(n1164) );
AND3_X1 U847 ( .A1(n1174), .A2(n1060), .A3(n1059), .ZN(n1134) );
AND4_X1 U848 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1089) );
AND4_X1 U849 ( .A1(n1181), .A2(n1182), .A3(n1183), .A4(n1184), .ZN(n1180) );
AND2_X1 U850 ( .A1(n1163), .A2(KEYINPUT14), .ZN(n1159) );
XNOR2_X1 U851 ( .A(n1185), .B(n1186), .ZN(n1163) );
NOR2_X1 U852 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U853 ( .A(n1189), .B(KEYINPUT52), .Z(n1188) );
NAND2_X1 U854 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U855 ( .A1(n1191), .A2(n1190), .ZN(n1187) );
XNOR2_X1 U856 ( .A(n1102), .B(n1192), .ZN(n1190) );
NAND2_X1 U857 ( .A1(KEYINPUT16), .A2(n1109), .ZN(n1185) );
NOR2_X1 U858 ( .A1(n1128), .A2(G952), .ZN(n1113) );
XNOR2_X1 U859 ( .A(G953), .B(KEYINPUT34), .ZN(n1128) );
XOR2_X1 U860 ( .A(n1179), .B(n1193), .Z(G48) );
NAND2_X1 U861 ( .A1(KEYINPUT37), .A2(G146), .ZN(n1193) );
NAND3_X1 U862 ( .A1(n1174), .A2(n1194), .A3(n1195), .ZN(n1179) );
XNOR2_X1 U863 ( .A(G143), .B(n1178), .ZN(G45) );
NAND3_X1 U864 ( .A1(n1196), .A2(n1058), .A3(n1197), .ZN(n1178) );
XNOR2_X1 U865 ( .A(G140), .B(n1184), .ZN(G42) );
NAND4_X1 U866 ( .A1(n1059), .A2(n1198), .A3(n1047), .A4(n1048), .ZN(n1184) );
XNOR2_X1 U867 ( .A(G137), .B(n1183), .ZN(G39) );
NAND4_X1 U868 ( .A1(n1199), .A2(n1198), .A3(n1194), .A4(n1048), .ZN(n1183) );
XNOR2_X1 U869 ( .A(n1200), .B(n1091), .ZN(G36) );
NAND4_X1 U870 ( .A1(n1058), .A2(n1198), .A3(n1175), .A4(n1176), .ZN(n1091) );
NAND2_X1 U871 ( .A1(KEYINPUT51), .A2(n1099), .ZN(n1200) );
XNOR2_X1 U872 ( .A(G131), .B(n1182), .ZN(G33) );
NAND3_X1 U873 ( .A1(n1058), .A2(n1198), .A3(n1059), .ZN(n1182) );
AND3_X1 U874 ( .A1(n1033), .A2(n1062), .A3(n1201), .ZN(n1198) );
AND3_X1 U875 ( .A1(n1202), .A2(n1040), .A3(n1063), .ZN(n1201) );
XOR2_X1 U876 ( .A(n1181), .B(n1203), .Z(G30) );
NAND2_X1 U877 ( .A1(KEYINPUT4), .A2(G128), .ZN(n1203) );
NAND4_X1 U878 ( .A1(n1197), .A2(n1194), .A3(n1048), .A4(n1176), .ZN(n1181) );
AND3_X1 U879 ( .A1(n1175), .A2(n1202), .A3(n1174), .ZN(n1197) );
NAND3_X1 U880 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(G3) );
NAND2_X1 U881 ( .A1(n1207), .A2(n1147), .ZN(n1206) );
NAND2_X1 U882 ( .A1(n1208), .A2(n1209), .ZN(n1205) );
INV_X1 U883 ( .A(KEYINPUT31), .ZN(n1209) );
NAND2_X1 U884 ( .A1(n1210), .A2(G101), .ZN(n1208) );
XNOR2_X1 U885 ( .A(KEYINPUT33), .B(n1207), .ZN(n1210) );
NAND2_X1 U886 ( .A1(KEYINPUT31), .A2(n1211), .ZN(n1204) );
NAND2_X1 U887 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
OR3_X1 U888 ( .A1(n1147), .A2(n1207), .A3(KEYINPUT33), .ZN(n1213) );
NAND2_X1 U889 ( .A1(KEYINPUT33), .A2(n1207), .ZN(n1212) );
INV_X1 U890 ( .A(n1171), .ZN(n1207) );
NAND4_X1 U891 ( .A1(n1199), .A2(n1058), .A3(n1174), .A4(n1136), .ZN(n1171) );
XNOR2_X1 U892 ( .A(G125), .B(n1177), .ZN(G27) );
NAND4_X1 U893 ( .A1(n1195), .A2(n1043), .A3(n1047), .A4(n1064), .ZN(n1177) );
AND3_X1 U894 ( .A1(n1048), .A2(n1202), .A3(n1059), .ZN(n1195) );
NAND2_X1 U895 ( .A1(n1061), .A2(n1214), .ZN(n1202) );
NAND4_X1 U896 ( .A1(G902), .A2(G953), .A3(n1215), .A4(n1094), .ZN(n1214) );
INV_X1 U897 ( .A(G900), .ZN(n1094) );
XNOR2_X1 U898 ( .A(G122), .B(n1170), .ZN(G24) );
NAND4_X1 U899 ( .A1(n1196), .A2(n1216), .A3(n1175), .A4(n1060), .ZN(n1170) );
NOR2_X1 U900 ( .A1(n1048), .A2(n1194), .ZN(n1060) );
NAND2_X1 U901 ( .A1(n1217), .A2(n1218), .ZN(G21) );
NAND2_X1 U902 ( .A1(G119), .A2(n1165), .ZN(n1218) );
XOR2_X1 U903 ( .A(n1219), .B(KEYINPUT48), .Z(n1217) );
OR2_X1 U904 ( .A1(n1165), .A2(G119), .ZN(n1219) );
NAND4_X1 U905 ( .A1(n1199), .A2(n1216), .A3(n1194), .A4(n1048), .ZN(n1165) );
INV_X1 U906 ( .A(n1047), .ZN(n1194) );
XNOR2_X1 U907 ( .A(G116), .B(n1169), .ZN(G18) );
NAND4_X1 U908 ( .A1(n1216), .A2(n1058), .A3(n1175), .A4(n1176), .ZN(n1169) );
XOR2_X1 U909 ( .A(n1220), .B(KEYINPUT2), .Z(n1175) );
XOR2_X1 U910 ( .A(n1168), .B(n1221), .Z(G15) );
XNOR2_X1 U911 ( .A(G113), .B(KEYINPUT23), .ZN(n1221) );
NAND3_X1 U912 ( .A1(n1216), .A2(n1058), .A3(n1059), .ZN(n1168) );
AND2_X1 U913 ( .A1(n1196), .A2(n1222), .ZN(n1059) );
INV_X1 U914 ( .A(n1176), .ZN(n1196) );
NOR2_X1 U915 ( .A1(n1048), .A2(n1047), .ZN(n1058) );
AND3_X1 U916 ( .A1(n1064), .A2(n1136), .A3(n1043), .ZN(n1216) );
NOR2_X1 U917 ( .A1(n1038), .A2(n1037), .ZN(n1043) );
INV_X1 U918 ( .A(n1057), .ZN(n1038) );
NOR2_X1 U919 ( .A1(n1062), .A2(n1041), .ZN(n1057) );
XOR2_X1 U920 ( .A(G110), .B(n1173), .Z(G12) );
AND4_X1 U921 ( .A1(n1048), .A2(n1136), .A3(n1047), .A4(n1223), .ZN(n1173) );
AND2_X1 U922 ( .A1(n1174), .A2(n1199), .ZN(n1223) );
INV_X1 U923 ( .A(n1065), .ZN(n1199) );
NAND2_X1 U924 ( .A1(n1222), .A2(n1176), .ZN(n1065) );
XNOR2_X1 U925 ( .A(n1224), .B(n1071), .ZN(n1176) );
XNOR2_X1 U926 ( .A(n1225), .B(G475), .ZN(n1071) );
NAND2_X1 U927 ( .A1(n1130), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U928 ( .A(n1227), .B(n1228), .ZN(n1130) );
XOR2_X1 U929 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U930 ( .A(G122), .B(G113), .Z(n1230) );
XOR2_X1 U931 ( .A(KEYINPUT29), .B(G131), .Z(n1229) );
XOR2_X1 U932 ( .A(n1231), .B(n1232), .Z(n1227) );
XNOR2_X1 U933 ( .A(G104), .B(n1233), .ZN(n1232) );
NAND2_X1 U934 ( .A1(n1234), .A2(G214), .ZN(n1233) );
XNOR2_X1 U935 ( .A(n1235), .B(n1236), .ZN(n1231) );
NOR2_X1 U936 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U937 ( .A(KEYINPUT0), .B(n1239), .Z(n1238) );
AND2_X1 U938 ( .A1(n1102), .A2(G140), .ZN(n1239) );
NOR2_X1 U939 ( .A1(G140), .A2(n1102), .ZN(n1237) );
XNOR2_X1 U940 ( .A(KEYINPUT41), .B(KEYINPUT10), .ZN(n1224) );
XNOR2_X1 U941 ( .A(KEYINPUT26), .B(n1220), .ZN(n1222) );
NAND2_X1 U942 ( .A1(n1240), .A2(n1241), .ZN(n1220) );
NAND2_X1 U943 ( .A1(G478), .A2(n1242), .ZN(n1241) );
XNOR2_X1 U944 ( .A(n1069), .B(KEYINPUT38), .ZN(n1240) );
NOR2_X1 U945 ( .A1(n1242), .A2(G478), .ZN(n1069) );
INV_X1 U946 ( .A(n1072), .ZN(n1242) );
NOR2_X1 U947 ( .A1(n1126), .A2(G902), .ZN(n1072) );
XNOR2_X1 U948 ( .A(n1243), .B(n1244), .ZN(n1126) );
NOR3_X1 U949 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
NOR2_X1 U950 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
INV_X1 U951 ( .A(n1250), .ZN(n1249) );
NOR2_X1 U952 ( .A1(n1251), .A2(n1252), .ZN(n1248) );
NOR4_X1 U953 ( .A1(n1250), .A2(n1252), .A3(KEYINPUT39), .A4(n1251), .ZN(n1246) );
INV_X1 U954 ( .A(KEYINPUT30), .ZN(n1252) );
XOR2_X1 U955 ( .A(G107), .B(n1253), .Z(n1250) );
NOR2_X1 U956 ( .A1(KEYINPUT61), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U957 ( .A(G116), .B(G122), .ZN(n1254) );
AND2_X1 U958 ( .A1(n1251), .A2(KEYINPUT39), .ZN(n1245) );
XNOR2_X1 U959 ( .A(n1255), .B(n1256), .ZN(n1251) );
XNOR2_X1 U960 ( .A(KEYINPUT21), .B(n1099), .ZN(n1256) );
XOR2_X1 U961 ( .A(n1257), .B(G128), .Z(n1255) );
NAND2_X1 U962 ( .A1(KEYINPUT36), .A2(n1258), .ZN(n1257) );
NAND2_X1 U963 ( .A1(KEYINPUT42), .A2(n1259), .ZN(n1243) );
NAND3_X1 U964 ( .A1(G234), .A2(n1087), .A3(G217), .ZN(n1259) );
NOR4_X1 U965 ( .A1(n1033), .A2(n1042), .A3(n1041), .A4(n1037), .ZN(n1174) );
INV_X1 U966 ( .A(n1040), .ZN(n1037) );
NAND2_X1 U967 ( .A1(G214), .A2(n1260), .ZN(n1040) );
INV_X1 U968 ( .A(n1063), .ZN(n1041) );
NAND2_X1 U969 ( .A1(G221), .A2(n1261), .ZN(n1063) );
INV_X1 U970 ( .A(n1062), .ZN(n1042) );
XNOR2_X1 U971 ( .A(n1262), .B(G469), .ZN(n1062) );
NAND2_X1 U972 ( .A1(n1263), .A2(n1226), .ZN(n1262) );
XOR2_X1 U973 ( .A(n1153), .B(n1264), .Z(n1263) );
XOR2_X1 U974 ( .A(n1265), .B(n1140), .Z(n1264) );
NOR2_X1 U975 ( .A1(KEYINPUT5), .A2(n1157), .ZN(n1265) );
NAND2_X1 U976 ( .A1(G227), .A2(n1087), .ZN(n1157) );
XNOR2_X1 U977 ( .A(n1266), .B(n1267), .ZN(n1153) );
INV_X1 U978 ( .A(n1100), .ZN(n1267) );
XOR2_X1 U979 ( .A(n1235), .B(n1268), .Z(n1100) );
XNOR2_X1 U980 ( .A(G140), .B(n1269), .ZN(n1268) );
NAND2_X1 U981 ( .A1(KEYINPUT13), .A2(G128), .ZN(n1269) );
INV_X1 U982 ( .A(n1064), .ZN(n1033) );
XOR2_X1 U983 ( .A(n1078), .B(n1082), .Z(n1064) );
NAND2_X1 U984 ( .A1(G210), .A2(n1260), .ZN(n1082) );
NAND2_X1 U985 ( .A1(n1270), .A2(n1226), .ZN(n1260) );
INV_X1 U986 ( .A(G237), .ZN(n1270) );
NAND2_X1 U987 ( .A1(n1271), .A2(n1226), .ZN(n1078) );
XOR2_X1 U988 ( .A(n1109), .B(n1272), .Z(n1271) );
XOR2_X1 U989 ( .A(n1273), .B(n1191), .Z(n1272) );
NAND2_X1 U990 ( .A1(G224), .A2(n1087), .ZN(n1191) );
NAND3_X1 U991 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
NAND2_X1 U992 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
OR3_X1 U993 ( .A1(n1278), .A2(n1277), .A3(KEYINPUT20), .ZN(n1275) );
XOR2_X1 U994 ( .A(n1144), .B(KEYINPUT50), .Z(n1277) );
OR2_X1 U995 ( .A1(G125), .A2(KEYINPUT18), .ZN(n1278) );
NAND2_X1 U996 ( .A1(KEYINPUT20), .A2(G125), .ZN(n1274) );
XNOR2_X1 U997 ( .A(n1279), .B(n1280), .ZN(n1109) );
XOR2_X1 U998 ( .A(G122), .B(n1266), .Z(n1280) );
XNOR2_X1 U999 ( .A(n1281), .B(n1282), .ZN(n1266) );
XOR2_X1 U1000 ( .A(G110), .B(G107), .Z(n1282) );
XNOR2_X1 U1001 ( .A(G104), .B(G101), .ZN(n1281) );
NAND2_X1 U1002 ( .A1(n1283), .A2(n1284), .ZN(n1279) );
NAND2_X1 U1003 ( .A1(n1285), .A2(G119), .ZN(n1284) );
NAND2_X1 U1004 ( .A1(n1286), .A2(n1287), .ZN(n1283) );
INV_X1 U1005 ( .A(G119), .ZN(n1287) );
XNOR2_X1 U1006 ( .A(KEYINPUT12), .B(n1285), .ZN(n1286) );
XNOR2_X1 U1007 ( .A(n1077), .B(G472), .ZN(n1047) );
AND2_X1 U1008 ( .A1(n1288), .A2(n1226), .ZN(n1077) );
XOR2_X1 U1009 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U1010 ( .A(n1291), .B(n1292), .Z(n1290) );
XOR2_X1 U1011 ( .A(n1149), .B(n1293), .Z(n1292) );
NOR2_X1 U1012 ( .A1(KEYINPUT17), .A2(n1143), .ZN(n1293) );
XNOR2_X1 U1013 ( .A(n1285), .B(G119), .ZN(n1143) );
XNOR2_X1 U1014 ( .A(G113), .B(n1294), .ZN(n1285) );
XNOR2_X1 U1015 ( .A(KEYINPUT11), .B(n1295), .ZN(n1294) );
INV_X1 U1016 ( .A(G116), .ZN(n1295) );
NAND2_X1 U1017 ( .A1(n1234), .A2(G210), .ZN(n1149) );
NOR2_X1 U1018 ( .A1(G953), .A2(G237), .ZN(n1234) );
NAND2_X1 U1019 ( .A1(KEYINPUT56), .A2(n1296), .ZN(n1291) );
XNOR2_X1 U1020 ( .A(KEYINPUT49), .B(n1147), .ZN(n1296) );
INV_X1 U1021 ( .A(G101), .ZN(n1147) );
XNOR2_X1 U1022 ( .A(n1192), .B(n1140), .ZN(n1289) );
XNOR2_X1 U1023 ( .A(n1297), .B(n1103), .ZN(n1140) );
XOR2_X1 U1024 ( .A(n1298), .B(G131), .Z(n1297) );
NAND2_X1 U1025 ( .A1(KEYINPUT35), .A2(n1099), .ZN(n1298) );
INV_X1 U1026 ( .A(G134), .ZN(n1099) );
INV_X1 U1027 ( .A(n1144), .ZN(n1192) );
XOR2_X1 U1028 ( .A(G128), .B(n1299), .Z(n1144) );
INV_X1 U1029 ( .A(n1235), .ZN(n1299) );
XOR2_X1 U1030 ( .A(G146), .B(n1258), .Z(n1235) );
XOR2_X1 U1031 ( .A(G143), .B(KEYINPUT28), .Z(n1258) );
NAND2_X1 U1032 ( .A1(n1061), .A2(n1300), .ZN(n1136) );
NAND3_X1 U1033 ( .A1(n1301), .A2(n1215), .A3(n1110), .ZN(n1300) );
NOR2_X1 U1034 ( .A1(n1087), .A2(G898), .ZN(n1110) );
XNOR2_X1 U1035 ( .A(KEYINPUT43), .B(n1226), .ZN(n1301) );
NAND3_X1 U1036 ( .A1(n1215), .A2(n1087), .A3(G952), .ZN(n1061) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1215) );
XNOR2_X1 U1038 ( .A(n1302), .B(n1303), .ZN(n1048) );
NOR2_X1 U1039 ( .A1(n1118), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U1040 ( .A(KEYINPUT46), .B(n1261), .ZN(n1304) );
NAND2_X1 U1041 ( .A1(G234), .A2(n1226), .ZN(n1261) );
INV_X1 U1042 ( .A(G902), .ZN(n1226) );
INV_X1 U1043 ( .A(G217), .ZN(n1118) );
OR2_X1 U1044 ( .A1(n1122), .A2(G902), .ZN(n1302) );
XNOR2_X1 U1045 ( .A(n1305), .B(n1306), .ZN(n1122) );
XOR2_X1 U1046 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1047 ( .A(G128), .B(G110), .Z(n1308) );
XOR2_X1 U1048 ( .A(KEYINPUT29), .B(G146), .Z(n1307) );
XOR2_X1 U1049 ( .A(n1309), .B(n1310), .Z(n1305) );
XOR2_X1 U1050 ( .A(n1311), .B(n1312), .Z(n1310) );
NOR2_X1 U1051 ( .A1(G119), .A2(KEYINPUT45), .ZN(n1312) );
AND3_X1 U1052 ( .A1(G221), .A2(n1087), .A3(G234), .ZN(n1311) );
INV_X1 U1053 ( .A(G953), .ZN(n1087) );
XOR2_X1 U1054 ( .A(n1313), .B(n1103), .Z(n1309) );
XOR2_X1 U1055 ( .A(G137), .B(KEYINPUT25), .Z(n1103) );
NAND2_X1 U1056 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NAND2_X1 U1057 ( .A1(n1316), .A2(n1102), .ZN(n1315) );
INV_X1 U1058 ( .A(G125), .ZN(n1102) );
XNOR2_X1 U1059 ( .A(G140), .B(n1317), .ZN(n1316) );
XNOR2_X1 U1060 ( .A(KEYINPUT63), .B(KEYINPUT55), .ZN(n1317) );
NAND2_X1 U1061 ( .A1(n1318), .A2(G125), .ZN(n1314) );
XNOR2_X1 U1062 ( .A(G140), .B(KEYINPUT15), .ZN(n1318) );
endmodule


