//Key = 1100110000110010011001101000011110001110111110011101101111100101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353;

XOR2_X1 U727 ( .A(n1013), .B(n1014), .Z(G9) );
XNOR2_X1 U728 ( .A(G107), .B(KEYINPUT15), .ZN(n1014) );
NAND2_X1 U729 ( .A1(KEYINPUT1), .A2(n1015), .ZN(n1013) );
NOR2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1018), .A2(n1019), .A3(G953), .A4(n1020), .ZN(n1017) );
NOR3_X1 U732 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1019) );
NOR2_X1 U733 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U734 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NAND3_X1 U735 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1018) );
NAND2_X1 U736 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NAND3_X1 U737 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1032) );
NAND2_X1 U738 ( .A1(KEYINPUT23), .A2(n1036), .ZN(n1035) );
NAND4_X1 U739 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
NAND3_X1 U740 ( .A1(n1039), .A2(n1041), .A3(n1037), .ZN(n1034) );
NAND2_X1 U741 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U743 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U744 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
XNOR2_X1 U745 ( .A(n1050), .B(KEYINPUT29), .ZN(n1048) );
NAND2_X1 U746 ( .A1(n1040), .A2(n1051), .ZN(n1042) );
NAND2_X1 U747 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
OR2_X1 U748 ( .A1(n1054), .A2(KEYINPUT23), .ZN(n1053) );
NAND2_X1 U749 ( .A1(n1055), .A2(n1056), .ZN(n1033) );
NAND2_X1 U750 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
INV_X1 U751 ( .A(n1021), .ZN(n1055) );
NAND3_X1 U752 ( .A1(n1044), .A2(n1040), .A3(n1037), .ZN(n1021) );
INV_X1 U753 ( .A(n1059), .ZN(n1037) );
NOR3_X1 U754 ( .A1(n1020), .A2(G953), .A3(G952), .ZN(n1016) );
AND4_X1 U755 ( .A1(n1044), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1020) );
NOR4_X1 U756 ( .A1(n1063), .A2(n1064), .A3(n1049), .A4(n1065), .ZN(n1062) );
NOR2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1061) );
AND2_X1 U758 ( .A1(n1023), .A2(KEYINPUT37), .ZN(n1067) );
INV_X1 U759 ( .A(n1039), .ZN(n1023) );
NOR2_X1 U760 ( .A1(KEYINPUT37), .A2(n1068), .ZN(n1066) );
XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n1069), .ZN(n1060) );
INV_X1 U762 ( .A(n1026), .ZN(n1069) );
XOR2_X1 U763 ( .A(n1070), .B(n1071), .Z(G72) );
NOR2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
AND4_X1 U765 ( .A1(KEYINPUT27), .A2(G900), .A3(G227), .A4(G953), .ZN(n1073) );
NOR2_X1 U766 ( .A1(KEYINPUT27), .A2(n1074), .ZN(n1072) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR2_X1 U768 ( .A1(G227), .A2(n1077), .ZN(n1075) );
XOR2_X1 U769 ( .A(n1078), .B(n1079), .Z(n1070) );
NOR2_X1 U770 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NOR2_X1 U771 ( .A1(n1082), .A2(KEYINPUT45), .ZN(n1081) );
NOR2_X1 U772 ( .A1(G953), .A2(n1028), .ZN(n1082) );
NOR3_X1 U773 ( .A1(n1028), .A2(KEYINPUT43), .A3(G953), .ZN(n1080) );
NAND2_X1 U774 ( .A1(n1083), .A2(n1084), .ZN(n1078) );
INV_X1 U775 ( .A(n1076), .ZN(n1084) );
XNOR2_X1 U776 ( .A(n1085), .B(n1086), .ZN(n1083) );
NAND2_X1 U777 ( .A1(n1087), .A2(KEYINPUT58), .ZN(n1085) );
XOR2_X1 U778 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U779 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NAND2_X1 U780 ( .A1(G131), .A2(n1092), .ZN(n1091) );
XOR2_X1 U781 ( .A(KEYINPUT57), .B(n1093), .Z(n1090) );
NOR2_X1 U782 ( .A1(G131), .A2(n1092), .ZN(n1093) );
NAND3_X1 U783 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1092) );
NAND2_X1 U784 ( .A1(KEYINPUT53), .A2(G137), .ZN(n1096) );
NAND3_X1 U785 ( .A1(n1097), .A2(n1098), .A3(G134), .ZN(n1095) );
NAND2_X1 U786 ( .A1(n1099), .A2(n1100), .ZN(n1094) );
NAND2_X1 U787 ( .A1(n1101), .A2(n1098), .ZN(n1099) );
INV_X1 U788 ( .A(KEYINPUT53), .ZN(n1098) );
XNOR2_X1 U789 ( .A(KEYINPUT21), .B(n1097), .ZN(n1101) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(G69) );
XOR2_X1 U791 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U792 ( .A1(G953), .A2(n1106), .ZN(n1105) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1106) );
NAND3_X1 U794 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1104) );
NAND2_X1 U795 ( .A1(G953), .A2(n1110), .ZN(n1109) );
NAND2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1108) );
NAND2_X1 U797 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NAND2_X1 U798 ( .A1(KEYINPUT7), .A2(n1115), .ZN(n1114) );
NAND2_X1 U799 ( .A1(n1116), .A2(n1117), .ZN(n1113) );
INV_X1 U800 ( .A(KEYINPUT7), .ZN(n1117) );
OR2_X1 U801 ( .A1(n1112), .A2(n1116), .ZN(n1107) );
NAND2_X1 U802 ( .A1(n1118), .A2(n1115), .ZN(n1116) );
NAND2_X1 U803 ( .A1(n1119), .A2(n1120), .ZN(n1115) );
NAND2_X1 U804 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U805 ( .A(n1123), .B(KEYINPUT13), .Z(n1119) );
OR2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1123) );
XNOR2_X1 U807 ( .A(KEYINPUT32), .B(KEYINPUT17), .ZN(n1118) );
NOR2_X1 U808 ( .A1(n1030), .A2(G953), .ZN(n1102) );
NOR2_X1 U809 ( .A1(n1124), .A2(n1125), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1126), .B(n1127), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NOR2_X1 U812 ( .A1(n1124), .A2(n1130), .ZN(G63) );
XOR2_X1 U813 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR2_X1 U814 ( .A1(n1133), .A2(n1129), .ZN(n1132) );
INV_X1 U815 ( .A(G478), .ZN(n1133) );
NOR2_X1 U816 ( .A1(n1124), .A2(n1134), .ZN(G60) );
XOR2_X1 U817 ( .A(n1135), .B(n1136), .Z(n1134) );
NOR2_X1 U818 ( .A1(n1137), .A2(n1129), .ZN(n1135) );
XNOR2_X1 U819 ( .A(G104), .B(n1138), .ZN(G6) );
NOR2_X1 U820 ( .A1(n1124), .A2(n1139), .ZN(G57) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U822 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U823 ( .A1(n1144), .A2(KEYINPUT9), .ZN(n1143) );
NOR2_X1 U824 ( .A1(n1145), .A2(n1129), .ZN(n1142) );
XOR2_X1 U825 ( .A(n1146), .B(n1147), .Z(n1140) );
NAND2_X1 U826 ( .A1(n1148), .A2(KEYINPUT31), .ZN(n1146) );
XNOR2_X1 U827 ( .A(n1149), .B(n1150), .ZN(n1148) );
NOR2_X1 U828 ( .A1(n1124), .A2(n1151), .ZN(G54) );
XOR2_X1 U829 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U830 ( .A(n1154), .B(n1155), .Z(n1152) );
NOR2_X1 U831 ( .A1(n1156), .A2(n1129), .ZN(n1155) );
INV_X1 U832 ( .A(G469), .ZN(n1156) );
NAND2_X1 U833 ( .A1(n1157), .A2(n1158), .ZN(n1154) );
NAND3_X1 U834 ( .A1(n1159), .A2(n1077), .A3(G227), .ZN(n1158) );
XOR2_X1 U835 ( .A(KEYINPUT49), .B(n1160), .Z(n1159) );
NAND2_X1 U836 ( .A1(n1160), .A2(n1161), .ZN(n1157) );
NAND2_X1 U837 ( .A1(G227), .A2(n1077), .ZN(n1161) );
XNOR2_X1 U838 ( .A(n1162), .B(n1163), .ZN(n1160) );
NOR2_X1 U839 ( .A1(n1077), .A2(G952), .ZN(n1124) );
NOR2_X1 U840 ( .A1(n1164), .A2(n1165), .ZN(G51) );
XOR2_X1 U841 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U842 ( .A1(n1168), .A2(n1129), .ZN(n1166) );
NAND2_X1 U843 ( .A1(G902), .A2(n1169), .ZN(n1129) );
NAND2_X1 U844 ( .A1(n1030), .A2(n1028), .ZN(n1169) );
AND4_X1 U845 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1028) );
NOR4_X1 U846 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
NOR2_X1 U847 ( .A1(n1178), .A2(n1179), .ZN(n1172) );
NOR2_X1 U848 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XNOR2_X1 U849 ( .A(KEYINPUT47), .B(n1182), .ZN(n1181) );
AND4_X1 U850 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1030) );
NOR4_X1 U851 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1186) );
NOR2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U853 ( .A(KEYINPUT4), .B(n1193), .ZN(n1192) );
INV_X1 U854 ( .A(n1138), .ZN(n1189) );
NAND4_X1 U855 ( .A1(n1194), .A2(n1195), .A3(n1044), .A4(n1196), .ZN(n1138) );
NOR4_X1 U856 ( .A1(n1197), .A2(n1198), .A3(n1058), .A4(n1052), .ZN(n1188) );
NOR2_X1 U857 ( .A1(KEYINPUT38), .A2(n1199), .ZN(n1198) );
AND3_X1 U858 ( .A1(n1040), .A2(n1182), .A3(n1200), .ZN(n1199) );
AND2_X1 U859 ( .A1(n1201), .A2(KEYINPUT38), .ZN(n1197) );
NOR3_X1 U860 ( .A1(n1202), .A2(n1052), .A3(n1203), .ZN(n1187) );
XNOR2_X1 U861 ( .A(KEYINPUT40), .B(n1046), .ZN(n1202) );
NOR2_X1 U862 ( .A1(n1015), .A2(n1204), .ZN(n1185) );
NOR3_X1 U863 ( .A1(n1054), .A2(n1205), .A3(n1203), .ZN(n1204) );
XNOR2_X1 U864 ( .A(n1195), .B(KEYINPUT20), .ZN(n1205) );
AND4_X1 U865 ( .A1(n1195), .A2(n1068), .A3(n1044), .A4(n1196), .ZN(n1015) );
NOR2_X1 U866 ( .A1(G952), .A2(n1206), .ZN(n1164) );
XNOR2_X1 U867 ( .A(G953), .B(KEYINPUT62), .ZN(n1206) );
XNOR2_X1 U868 ( .A(n1178), .B(n1207), .ZN(G48) );
NAND2_X1 U869 ( .A1(KEYINPUT18), .A2(G146), .ZN(n1207) );
AND3_X1 U870 ( .A1(n1194), .A2(n1025), .A3(n1208), .ZN(n1178) );
XOR2_X1 U871 ( .A(n1209), .B(n1210), .Z(G45) );
NAND2_X1 U872 ( .A1(KEYINPUT56), .A2(G143), .ZN(n1210) );
OR2_X1 U873 ( .A1(n1180), .A2(n1182), .ZN(n1209) );
NAND4_X1 U874 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1180) );
XOR2_X1 U875 ( .A(n1215), .B(G140), .Z(G42) );
NAND2_X1 U876 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND2_X1 U877 ( .A1(n1177), .A2(n1218), .ZN(n1217) );
INV_X1 U878 ( .A(KEYINPUT35), .ZN(n1218) );
AND3_X1 U879 ( .A1(n1031), .A2(n1038), .A3(n1219), .ZN(n1177) );
NAND4_X1 U880 ( .A1(n1038), .A2(n1220), .A3(n1219), .A4(KEYINPUT35), .ZN(n1216) );
INV_X1 U881 ( .A(n1031), .ZN(n1220) );
XNOR2_X1 U882 ( .A(n1097), .B(n1176), .ZN(G39) );
AND3_X1 U883 ( .A1(n1031), .A2(n1039), .A3(n1208), .ZN(n1176) );
XNOR2_X1 U884 ( .A(n1175), .B(n1221), .ZN(G36) );
NAND2_X1 U885 ( .A1(KEYINPUT63), .A2(G134), .ZN(n1221) );
AND4_X1 U886 ( .A1(n1031), .A2(n1211), .A3(n1212), .A4(n1068), .ZN(n1175) );
XNOR2_X1 U887 ( .A(n1174), .B(n1222), .ZN(G33) );
NAND2_X1 U888 ( .A1(KEYINPUT51), .A2(G131), .ZN(n1222) );
AND3_X1 U889 ( .A1(n1031), .A2(n1212), .A3(n1219), .ZN(n1174) );
AND2_X1 U890 ( .A1(n1211), .A2(n1194), .ZN(n1219) );
NOR2_X1 U891 ( .A1(n1026), .A2(n1065), .ZN(n1031) );
INV_X1 U892 ( .A(n1027), .ZN(n1065) );
XNOR2_X1 U893 ( .A(G128), .B(n1170), .ZN(G30) );
NAND3_X1 U894 ( .A1(n1068), .A2(n1025), .A3(n1208), .ZN(n1170) );
AND3_X1 U895 ( .A1(n1223), .A2(n1224), .A3(n1211), .ZN(n1208) );
AND2_X1 U896 ( .A1(n1195), .A2(n1225), .ZN(n1211) );
XOR2_X1 U897 ( .A(G101), .B(n1226), .Z(G3) );
AND2_X1 U898 ( .A1(n1212), .A2(n1227), .ZN(n1226) );
XNOR2_X1 U899 ( .A(G125), .B(n1171), .ZN(G27) );
NAND4_X1 U900 ( .A1(n1040), .A2(n1225), .A3(n1025), .A4(n1228), .ZN(n1171) );
NOR2_X1 U901 ( .A1(n1057), .A2(n1054), .ZN(n1228) );
INV_X1 U902 ( .A(n1038), .ZN(n1054) );
NAND2_X1 U903 ( .A1(n1229), .A2(n1059), .ZN(n1225) );
NAND3_X1 U904 ( .A1(G902), .A2(n1230), .A3(n1076), .ZN(n1229) );
NOR2_X1 U905 ( .A1(n1077), .A2(G900), .ZN(n1076) );
XOR2_X1 U906 ( .A(n1231), .B(n1232), .Z(G24) );
NOR2_X1 U907 ( .A1(n1193), .A2(n1191), .ZN(n1232) );
NAND3_X1 U908 ( .A1(n1213), .A2(n1214), .A3(n1233), .ZN(n1191) );
INV_X1 U909 ( .A(n1044), .ZN(n1193) );
NOR2_X1 U910 ( .A1(n1224), .A2(n1223), .ZN(n1044) );
NOR2_X1 U911 ( .A1(KEYINPUT39), .A2(n1234), .ZN(n1231) );
XNOR2_X1 U912 ( .A(G119), .B(n1183), .ZN(G21) );
NAND4_X1 U913 ( .A1(n1235), .A2(n1040), .A3(n1223), .A4(n1224), .ZN(n1183) );
INV_X1 U914 ( .A(n1203), .ZN(n1235) );
XOR2_X1 U915 ( .A(G116), .B(n1236), .Z(G18) );
NOR4_X1 U916 ( .A1(KEYINPUT26), .A2(n1058), .A3(n1201), .A4(n1052), .ZN(n1236) );
INV_X1 U917 ( .A(n1068), .ZN(n1058) );
NOR2_X1 U918 ( .A1(n1214), .A2(n1237), .ZN(n1068) );
XNOR2_X1 U919 ( .A(G113), .B(n1184), .ZN(G15) );
NAND3_X1 U920 ( .A1(n1194), .A2(n1233), .A3(n1212), .ZN(n1184) );
INV_X1 U921 ( .A(n1052), .ZN(n1212) );
NAND2_X1 U922 ( .A1(n1238), .A2(n1223), .ZN(n1052) );
INV_X1 U923 ( .A(n1201), .ZN(n1233) );
NAND2_X1 U924 ( .A1(n1196), .A2(n1040), .ZN(n1201) );
NAND2_X1 U925 ( .A1(n1239), .A2(n1240), .ZN(n1040) );
OR2_X1 U926 ( .A1(n1046), .A2(KEYINPUT29), .ZN(n1240) );
NAND3_X1 U927 ( .A1(n1050), .A2(n1241), .A3(KEYINPUT29), .ZN(n1239) );
INV_X1 U928 ( .A(n1057), .ZN(n1194) );
NAND2_X1 U929 ( .A1(n1237), .A2(n1214), .ZN(n1057) );
INV_X1 U930 ( .A(n1213), .ZN(n1237) );
XOR2_X1 U931 ( .A(n1242), .B(n1243), .Z(G12) );
NAND2_X1 U932 ( .A1(n1227), .A2(n1038), .ZN(n1243) );
NOR2_X1 U933 ( .A1(n1223), .A2(n1238), .ZN(n1038) );
INV_X1 U934 ( .A(n1224), .ZN(n1238) );
XOR2_X1 U935 ( .A(n1244), .B(n1128), .Z(n1224) );
NAND2_X1 U936 ( .A1(G217), .A2(n1245), .ZN(n1128) );
NAND2_X1 U937 ( .A1(n1246), .A2(n1126), .ZN(n1244) );
NAND3_X1 U938 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1126) );
NAND2_X1 U939 ( .A1(KEYINPUT50), .A2(n1250), .ZN(n1249) );
OR3_X1 U940 ( .A1(n1250), .A2(KEYINPUT50), .A3(n1251), .ZN(n1248) );
NAND2_X1 U941 ( .A1(n1251), .A2(n1252), .ZN(n1247) );
NAND2_X1 U942 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
INV_X1 U943 ( .A(KEYINPUT50), .ZN(n1254) );
XNOR2_X1 U944 ( .A(n1250), .B(KEYINPUT34), .ZN(n1253) );
XNOR2_X1 U945 ( .A(n1255), .B(n1256), .ZN(n1250) );
XOR2_X1 U946 ( .A(KEYINPUT30), .B(G146), .Z(n1256) );
XNOR2_X1 U947 ( .A(n1257), .B(n1258), .ZN(n1255) );
INV_X1 U948 ( .A(n1086), .ZN(n1258) );
NAND3_X1 U949 ( .A1(n1259), .A2(n1260), .A3(n1261), .ZN(n1257) );
NAND2_X1 U950 ( .A1(n1262), .A2(n1162), .ZN(n1261) );
NAND3_X1 U951 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1262) );
NAND2_X1 U952 ( .A1(KEYINPUT8), .A2(n1266), .ZN(n1265) );
NAND2_X1 U953 ( .A1(KEYINPUT41), .A2(n1267), .ZN(n1264) );
NAND2_X1 U954 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U955 ( .A1(KEYINPUT28), .A2(n1270), .ZN(n1269) );
NAND2_X1 U956 ( .A1(n1268), .A2(n1271), .ZN(n1263) );
INV_X1 U957 ( .A(KEYINPUT41), .ZN(n1271) );
NAND4_X1 U958 ( .A1(n1268), .A2(n1266), .A3(G110), .A4(n1270), .ZN(n1260) );
INV_X1 U959 ( .A(KEYINPUT8), .ZN(n1270) );
INV_X1 U960 ( .A(KEYINPUT28), .ZN(n1266) );
NAND2_X1 U961 ( .A1(KEYINPUT8), .A2(n1272), .ZN(n1259) );
NAND2_X1 U962 ( .A1(n1268), .A2(n1273), .ZN(n1272) );
NAND2_X1 U963 ( .A1(KEYINPUT28), .A2(G110), .ZN(n1273) );
XOR2_X1 U964 ( .A(G119), .B(G128), .Z(n1268) );
XOR2_X1 U965 ( .A(G137), .B(n1274), .Z(n1251) );
AND3_X1 U966 ( .A1(G221), .A2(n1077), .A3(G234), .ZN(n1274) );
XOR2_X1 U967 ( .A(n1275), .B(n1145), .Z(n1223) );
INV_X1 U968 ( .A(G472), .ZN(n1145) );
NAND2_X1 U969 ( .A1(n1276), .A2(n1246), .ZN(n1275) );
XOR2_X1 U970 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U971 ( .A(n1279), .B(n1280), .Z(n1278) );
NAND2_X1 U972 ( .A1(KEYINPUT0), .A2(n1150), .ZN(n1279) );
NAND3_X1 U973 ( .A1(n1281), .A2(n1077), .A3(G210), .ZN(n1150) );
XOR2_X1 U974 ( .A(KEYINPUT44), .B(n1144), .Z(n1277) );
AND2_X1 U975 ( .A1(n1282), .A2(n1283), .ZN(n1144) );
NAND2_X1 U976 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U977 ( .A(KEYINPUT22), .B(n1286), .Z(n1282) );
NOR2_X1 U978 ( .A1(n1284), .A2(n1285), .ZN(n1286) );
XNOR2_X1 U979 ( .A(n1287), .B(KEYINPUT48), .ZN(n1284) );
NOR2_X1 U980 ( .A1(n1203), .A2(n1046), .ZN(n1227) );
INV_X1 U981 ( .A(n1195), .ZN(n1046) );
NOR2_X1 U982 ( .A1(n1050), .A2(n1049), .ZN(n1195) );
INV_X1 U983 ( .A(n1241), .ZN(n1049) );
NAND2_X1 U984 ( .A1(n1288), .A2(G221), .ZN(n1241) );
XOR2_X1 U985 ( .A(n1245), .B(KEYINPUT33), .Z(n1288) );
NAND2_X1 U986 ( .A1(G234), .A2(n1246), .ZN(n1245) );
AND3_X1 U987 ( .A1(n1289), .A2(n1290), .A3(n1291), .ZN(n1050) );
INV_X1 U988 ( .A(n1063), .ZN(n1291) );
NOR2_X1 U989 ( .A1(n1292), .A2(G469), .ZN(n1063) );
OR2_X1 U990 ( .A1(G469), .A2(KEYINPUT55), .ZN(n1290) );
NAND2_X1 U991 ( .A1(n1064), .A2(KEYINPUT55), .ZN(n1289) );
AND2_X1 U992 ( .A1(G469), .A2(n1292), .ZN(n1064) );
NAND2_X1 U993 ( .A1(n1293), .A2(n1246), .ZN(n1292) );
XNOR2_X1 U994 ( .A(n1153), .B(n1294), .ZN(n1293) );
XOR2_X1 U995 ( .A(n1295), .B(n1296), .Z(n1294) );
NAND2_X1 U996 ( .A1(KEYINPUT24), .A2(G227), .ZN(n1296) );
NAND3_X1 U997 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1295) );
NAND2_X1 U998 ( .A1(n1163), .A2(n1300), .ZN(n1299) );
INV_X1 U999 ( .A(KEYINPUT36), .ZN(n1300) );
NAND3_X1 U1000 ( .A1(KEYINPUT36), .A2(n1301), .A3(n1162), .ZN(n1298) );
OR2_X1 U1001 ( .A1(n1162), .A2(n1301), .ZN(n1297) );
NOR2_X1 U1002 ( .A1(KEYINPUT59), .A2(n1163), .ZN(n1301) );
XNOR2_X1 U1003 ( .A(n1280), .B(n1302), .ZN(n1153) );
XNOR2_X1 U1004 ( .A(G107), .B(n1303), .ZN(n1302) );
NAND2_X1 U1005 ( .A1(KEYINPUT52), .A2(n1304), .ZN(n1303) );
XOR2_X1 U1006 ( .A(n1147), .B(n1149), .Z(n1280) );
XNOR2_X1 U1007 ( .A(n1305), .B(n1089), .ZN(n1147) );
NAND3_X1 U1008 ( .A1(n1306), .A2(n1307), .A3(n1308), .ZN(n1305) );
NAND2_X1 U1009 ( .A1(G131), .A2(n1309), .ZN(n1308) );
NAND2_X1 U1010 ( .A1(KEYINPUT3), .A2(n1310), .ZN(n1307) );
NAND2_X1 U1011 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
XNOR2_X1 U1012 ( .A(n1313), .B(n1309), .ZN(n1311) );
NAND2_X1 U1013 ( .A1(n1314), .A2(n1315), .ZN(n1306) );
INV_X1 U1014 ( .A(KEYINPUT3), .ZN(n1315) );
NAND2_X1 U1015 ( .A1(n1316), .A2(n1317), .ZN(n1314) );
NAND2_X1 U1016 ( .A1(n1309), .A2(n1313), .ZN(n1317) );
OR3_X1 U1017 ( .A1(n1309), .A2(G131), .A3(n1313), .ZN(n1316) );
INV_X1 U1018 ( .A(KEYINPUT11), .ZN(n1313) );
XNOR2_X1 U1019 ( .A(G134), .B(n1097), .ZN(n1309) );
INV_X1 U1020 ( .A(G137), .ZN(n1097) );
NAND2_X1 U1021 ( .A1(n1039), .A2(n1196), .ZN(n1203) );
AND2_X1 U1022 ( .A1(n1025), .A2(n1200), .ZN(n1196) );
NAND2_X1 U1023 ( .A1(n1059), .A2(n1318), .ZN(n1200) );
NAND4_X1 U1024 ( .A1(G953), .A2(G902), .A3(n1230), .A4(n1110), .ZN(n1318) );
INV_X1 U1025 ( .A(G898), .ZN(n1110) );
NAND3_X1 U1026 ( .A1(n1230), .A2(n1077), .A3(G952), .ZN(n1059) );
NAND2_X1 U1027 ( .A1(G237), .A2(G234), .ZN(n1230) );
INV_X1 U1028 ( .A(n1182), .ZN(n1025) );
NAND2_X1 U1029 ( .A1(n1026), .A2(n1027), .ZN(n1182) );
NAND2_X1 U1030 ( .A1(G214), .A2(n1319), .ZN(n1027) );
XOR2_X1 U1031 ( .A(n1320), .B(n1168), .Z(n1026) );
NAND2_X1 U1032 ( .A1(G210), .A2(n1319), .ZN(n1168) );
NAND2_X1 U1033 ( .A1(n1281), .A2(n1246), .ZN(n1319) );
INV_X1 U1034 ( .A(G237), .ZN(n1281) );
NAND2_X1 U1035 ( .A1(n1321), .A2(n1246), .ZN(n1320) );
INV_X1 U1036 ( .A(G902), .ZN(n1246) );
XOR2_X1 U1037 ( .A(n1167), .B(n1322), .Z(n1321) );
XOR2_X1 U1038 ( .A(KEYINPUT54), .B(KEYINPUT12), .Z(n1322) );
XNOR2_X1 U1039 ( .A(n1323), .B(n1324), .ZN(n1167) );
XNOR2_X1 U1040 ( .A(n1112), .B(n1325), .ZN(n1324) );
XNOR2_X1 U1041 ( .A(n1121), .B(n1089), .ZN(n1325) );
XOR2_X1 U1042 ( .A(G128), .B(n1326), .Z(n1089) );
XOR2_X1 U1043 ( .A(n1285), .B(n1287), .Z(n1121) );
XNOR2_X1 U1044 ( .A(G116), .B(G119), .ZN(n1285) );
XNOR2_X1 U1045 ( .A(n1234), .B(n1162), .ZN(n1112) );
INV_X1 U1046 ( .A(G110), .ZN(n1162) );
XOR2_X1 U1047 ( .A(n1327), .B(n1328), .Z(n1323) );
XNOR2_X1 U1048 ( .A(KEYINPUT19), .B(n1329), .ZN(n1328) );
INV_X1 U1049 ( .A(G125), .ZN(n1329) );
XOR2_X1 U1050 ( .A(n1330), .B(n1331), .Z(n1327) );
AND2_X1 U1051 ( .A1(n1077), .A2(G224), .ZN(n1331) );
NAND2_X1 U1052 ( .A1(KEYINPUT5), .A2(n1122), .ZN(n1330) );
XNOR2_X1 U1053 ( .A(n1332), .B(n1149), .ZN(n1122) );
XNOR2_X1 U1054 ( .A(G101), .B(KEYINPUT16), .ZN(n1149) );
NAND2_X1 U1055 ( .A1(n1333), .A2(KEYINPUT42), .ZN(n1332) );
XNOR2_X1 U1056 ( .A(G104), .B(n1334), .ZN(n1333) );
XNOR2_X1 U1057 ( .A(KEYINPUT46), .B(n1335), .ZN(n1334) );
INV_X1 U1058 ( .A(G107), .ZN(n1335) );
NOR2_X1 U1059 ( .A1(n1213), .A2(n1214), .ZN(n1039) );
XOR2_X1 U1060 ( .A(n1336), .B(n1137), .Z(n1214) );
INV_X1 U1061 ( .A(G475), .ZN(n1137) );
OR2_X1 U1062 ( .A1(n1136), .A2(G902), .ZN(n1336) );
XNOR2_X1 U1063 ( .A(n1337), .B(n1338), .ZN(n1136) );
XOR2_X1 U1064 ( .A(n1339), .B(n1340), .Z(n1338) );
XNOR2_X1 U1065 ( .A(n1304), .B(n1341), .ZN(n1340) );
NOR4_X1 U1066 ( .A1(KEYINPUT2), .A2(G953), .A3(G237), .A4(n1342), .ZN(n1341) );
INV_X1 U1067 ( .A(G214), .ZN(n1342) );
INV_X1 U1068 ( .A(G104), .ZN(n1304) );
XNOR2_X1 U1069 ( .A(n1312), .B(G122), .ZN(n1339) );
INV_X1 U1070 ( .A(G131), .ZN(n1312) );
XNOR2_X1 U1071 ( .A(n1086), .B(n1343), .ZN(n1337) );
XNOR2_X1 U1072 ( .A(n1344), .B(n1326), .ZN(n1343) );
XOR2_X1 U1073 ( .A(G143), .B(G146), .Z(n1326) );
INV_X1 U1074 ( .A(n1287), .ZN(n1344) );
XOR2_X1 U1075 ( .A(G113), .B(KEYINPUT14), .Z(n1287) );
XOR2_X1 U1076 ( .A(G125), .B(n1163), .Z(n1086) );
XOR2_X1 U1077 ( .A(G140), .B(KEYINPUT25), .Z(n1163) );
XOR2_X1 U1078 ( .A(G478), .B(n1345), .Z(n1213) );
NOR2_X1 U1079 ( .A1(G902), .A2(n1131), .ZN(n1345) );
XOR2_X1 U1080 ( .A(n1346), .B(n1347), .Z(n1131) );
NOR2_X1 U1081 ( .A1(KEYINPUT6), .A2(n1348), .ZN(n1347) );
XOR2_X1 U1082 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1083 ( .A(G128), .B(n1351), .Z(n1350) );
XNOR2_X1 U1084 ( .A(G143), .B(n1100), .ZN(n1351) );
INV_X1 U1085 ( .A(G134), .ZN(n1100) );
XNOR2_X1 U1086 ( .A(G107), .B(n1352), .ZN(n1349) );
XNOR2_X1 U1087 ( .A(n1234), .B(G116), .ZN(n1352) );
INV_X1 U1088 ( .A(G122), .ZN(n1234) );
NAND3_X1 U1089 ( .A1(n1353), .A2(n1077), .A3(G217), .ZN(n1346) );
INV_X1 U1090 ( .A(G953), .ZN(n1077) );
XOR2_X1 U1091 ( .A(KEYINPUT60), .B(G234), .Z(n1353) );
NAND2_X1 U1092 ( .A1(KEYINPUT10), .A2(G110), .ZN(n1242) );
endmodule


