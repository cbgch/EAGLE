//Key = 1000111001001001100011001110100101011100000110110000010100001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392;

XNOR2_X1 U772 ( .A(n1059), .B(n1060), .ZN(G9) );
NOR2_X1 U773 ( .A1(n1061), .A2(n1062), .ZN(G75) );
XOR2_X1 U774 ( .A(KEYINPUT3), .B(n1063), .Z(n1062) );
NOR3_X1 U775 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NOR2_X1 U776 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U777 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR2_X1 U778 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U779 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
NOR2_X1 U780 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NOR3_X1 U781 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1075) );
NOR3_X1 U782 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
XOR2_X1 U783 ( .A(n1083), .B(KEYINPUT38), .Z(n1082) );
NOR3_X1 U784 ( .A1(n1084), .A2(n1085), .A3(n1083), .ZN(n1078) );
NOR2_X1 U785 ( .A1(n1086), .A2(n1087), .ZN(n1077) );
NOR2_X1 U786 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR3_X1 U787 ( .A1(n1087), .A2(n1090), .A3(n1083), .ZN(n1073) );
NOR2_X1 U788 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
AND2_X1 U789 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NOR3_X1 U790 ( .A1(n1087), .A2(n1095), .A3(n1083), .ZN(n1069) );
NOR2_X1 U791 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U792 ( .A1(n1076), .A2(n1098), .ZN(n1097) );
NOR2_X1 U793 ( .A1(n1099), .A2(n1100), .ZN(n1096) );
XNOR2_X1 U794 ( .A(n1076), .B(KEYINPUT53), .ZN(n1100) );
INV_X1 U795 ( .A(n1101), .ZN(n1076) );
INV_X1 U796 ( .A(n1102), .ZN(n1087) );
NOR2_X1 U797 ( .A1(G952), .A2(n1066), .ZN(n1061) );
NAND2_X1 U798 ( .A1(n1103), .A2(n1104), .ZN(n1066) );
NAND4_X1 U799 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1104) );
NOR4_X1 U800 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
XNOR2_X1 U801 ( .A(KEYINPUT52), .B(n1113), .ZN(n1112) );
XOR2_X1 U802 ( .A(KEYINPUT9), .B(n1114), .Z(n1111) );
NOR2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U804 ( .A(KEYINPUT56), .B(n1117), .Z(n1110) );
AND2_X1 U805 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR3_X1 U806 ( .A1(n1120), .A2(n1094), .A3(n1084), .ZN(n1107) );
NOR2_X1 U807 ( .A1(n1119), .A2(n1118), .ZN(n1120) );
XNOR2_X1 U808 ( .A(n1121), .B(n1122), .ZN(n1106) );
NOR2_X1 U809 ( .A1(G469), .A2(KEYINPUT13), .ZN(n1122) );
XOR2_X1 U810 ( .A(n1123), .B(n1124), .Z(G72) );
NOR2_X1 U811 ( .A1(n1125), .A2(G953), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U813 ( .A1(n1128), .A2(n1129), .ZN(n1123) );
NAND2_X1 U814 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
OR2_X1 U815 ( .A1(n1132), .A2(G227), .ZN(n1131) );
NAND2_X1 U816 ( .A1(G953), .A2(n1133), .ZN(n1128) );
NAND2_X1 U817 ( .A1(G900), .A2(n1134), .ZN(n1133) );
OR2_X1 U818 ( .A1(n1130), .A2(G227), .ZN(n1134) );
XNOR2_X1 U819 ( .A(n1135), .B(n1136), .ZN(n1130) );
XOR2_X1 U820 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U821 ( .A(KEYINPUT58), .B(n1139), .ZN(n1138) );
XOR2_X1 U822 ( .A(n1140), .B(n1141), .Z(n1135) );
NAND2_X1 U823 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NAND2_X1 U824 ( .A1(KEYINPUT0), .A2(n1144), .ZN(n1143) );
OR3_X1 U825 ( .A1(n1145), .A2(G137), .A3(KEYINPUT0), .ZN(n1142) );
INV_X1 U826 ( .A(G134), .ZN(n1145) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(G69) );
NOR2_X1 U828 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND3_X1 U829 ( .A1(n1150), .A2(n1151), .A3(n1152), .ZN(n1146) );
INV_X1 U830 ( .A(n1148), .ZN(n1152) );
OR2_X1 U831 ( .A1(n1132), .A2(G224), .ZN(n1151) );
NAND2_X1 U832 ( .A1(n1153), .A2(n1132), .ZN(n1150) );
NOR2_X1 U833 ( .A1(n1154), .A2(n1155), .ZN(G66) );
XOR2_X1 U834 ( .A(n1156), .B(n1157), .Z(n1155) );
NAND2_X1 U835 ( .A1(n1158), .A2(n1159), .ZN(n1156) );
XOR2_X1 U836 ( .A(KEYINPUT11), .B(G217), .Z(n1159) );
NOR2_X1 U837 ( .A1(n1154), .A2(n1160), .ZN(G63) );
XOR2_X1 U838 ( .A(n1161), .B(n1162), .Z(n1160) );
NAND3_X1 U839 ( .A1(n1163), .A2(n1164), .A3(G478), .ZN(n1161) );
OR2_X1 U840 ( .A1(n1158), .A2(KEYINPUT34), .ZN(n1164) );
NAND2_X1 U841 ( .A1(KEYINPUT34), .A2(n1165), .ZN(n1163) );
NAND2_X1 U842 ( .A1(n1064), .A2(n1166), .ZN(n1165) );
NOR2_X1 U843 ( .A1(n1154), .A2(n1167), .ZN(G60) );
XOR2_X1 U844 ( .A(n1168), .B(n1169), .Z(n1167) );
AND2_X1 U845 ( .A1(G475), .A2(n1158), .ZN(n1169) );
NAND2_X1 U846 ( .A1(KEYINPUT47), .A2(n1170), .ZN(n1168) );
XNOR2_X1 U847 ( .A(n1171), .B(n1172), .ZN(G6) );
NOR2_X1 U848 ( .A1(n1154), .A2(n1173), .ZN(G57) );
XOR2_X1 U849 ( .A(n1174), .B(n1175), .Z(n1173) );
XOR2_X1 U850 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U851 ( .A(n1178), .B(n1179), .Z(n1174) );
XOR2_X1 U852 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U853 ( .A1(n1158), .A2(G472), .ZN(n1180) );
NOR2_X1 U854 ( .A1(n1154), .A2(n1182), .ZN(G54) );
XOR2_X1 U855 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U856 ( .A1(n1158), .A2(G469), .ZN(n1184) );
NAND2_X1 U857 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
NAND2_X1 U858 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U859 ( .A(n1189), .B(KEYINPUT54), .Z(n1185) );
OR2_X1 U860 ( .A1(n1188), .A2(n1187), .ZN(n1189) );
XNOR2_X1 U861 ( .A(n1190), .B(n1191), .ZN(n1187) );
NOR2_X1 U862 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
AND3_X1 U863 ( .A1(KEYINPUT40), .A2(n1194), .A3(G110), .ZN(n1193) );
INV_X1 U864 ( .A(G140), .ZN(n1194) );
NOR2_X1 U865 ( .A1(KEYINPUT40), .A2(n1195), .ZN(n1192) );
XNOR2_X1 U866 ( .A(n1181), .B(n1196), .ZN(n1188) );
XOR2_X1 U867 ( .A(n1197), .B(n1141), .Z(n1196) );
NOR2_X1 U868 ( .A1(KEYINPUT57), .A2(n1198), .ZN(n1197) );
NOR2_X1 U869 ( .A1(n1154), .A2(n1199), .ZN(G51) );
XOR2_X1 U870 ( .A(n1200), .B(n1201), .Z(n1199) );
NOR2_X1 U871 ( .A1(KEYINPUT27), .A2(n1202), .ZN(n1201) );
NOR2_X1 U872 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
XOR2_X1 U873 ( .A(n1205), .B(KEYINPUT24), .Z(n1204) );
NAND2_X1 U874 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U875 ( .A1(n1206), .A2(n1207), .ZN(n1203) );
XNOR2_X1 U876 ( .A(n1208), .B(n1209), .ZN(n1207) );
NOR2_X1 U877 ( .A1(KEYINPUT59), .A2(n1210), .ZN(n1209) );
NAND2_X1 U878 ( .A1(n1158), .A2(n1211), .ZN(n1200) );
AND2_X1 U879 ( .A1(G902), .A2(n1064), .ZN(n1158) );
OR3_X1 U880 ( .A1(n1127), .A2(n1153), .A3(n1212), .ZN(n1064) );
XOR2_X1 U881 ( .A(n1126), .B(KEYINPUT22), .Z(n1212) );
NAND2_X1 U882 ( .A1(n1213), .A2(n1214), .ZN(n1153) );
NOR4_X1 U883 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1060), .ZN(n1214) );
NOR3_X1 U884 ( .A1(n1218), .A2(n1098), .A3(n1083), .ZN(n1060) );
NOR4_X1 U885 ( .A1(n1172), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1213) );
AND2_X1 U886 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
NOR3_X1 U887 ( .A1(n1072), .A2(n1218), .A3(n1224), .ZN(n1220) );
NOR3_X1 U888 ( .A1(n1083), .A2(n1218), .A3(n1099), .ZN(n1172) );
NAND4_X1 U889 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1127) );
NOR3_X1 U890 ( .A1(n1229), .A2(n1230), .A3(n1231), .ZN(n1228) );
INV_X1 U891 ( .A(n1232), .ZN(n1230) );
NAND2_X1 U892 ( .A1(KEYINPUT63), .A2(n1233), .ZN(n1227) );
INV_X1 U893 ( .A(n1234), .ZN(n1233) );
NAND2_X1 U894 ( .A1(n1235), .A2(n1236), .ZN(n1225) );
NAND2_X1 U895 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND4_X1 U896 ( .A1(n1089), .A2(n1109), .A3(n1239), .A4(n1240), .ZN(n1238) );
NOR2_X1 U897 ( .A1(KEYINPUT63), .A2(n1092), .ZN(n1239) );
NAND3_X1 U898 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1237) );
NAND2_X1 U899 ( .A1(n1244), .A2(n1245), .ZN(n1242) );
OR2_X1 U900 ( .A1(n1099), .A2(KEYINPUT12), .ZN(n1244) );
NAND3_X1 U901 ( .A1(n1246), .A2(n1098), .A3(n1092), .ZN(n1241) );
NAND2_X1 U902 ( .A1(KEYINPUT12), .A2(n1247), .ZN(n1246) );
NOR2_X1 U903 ( .A1(n1132), .A2(G952), .ZN(n1154) );
XNOR2_X1 U904 ( .A(G146), .B(n1248), .ZN(G48) );
NAND4_X1 U905 ( .A1(n1243), .A2(n1247), .A3(n1235), .A4(n1092), .ZN(n1248) );
XNOR2_X1 U906 ( .A(G143), .B(n1234), .ZN(G45) );
NAND4_X1 U907 ( .A1(n1089), .A2(n1235), .A3(n1249), .A4(n1092), .ZN(n1234) );
NOR2_X1 U908 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
XNOR2_X1 U909 ( .A(G140), .B(n1226), .ZN(G42) );
NAND3_X1 U910 ( .A1(n1252), .A2(n1247), .A3(n1088), .ZN(n1226) );
XNOR2_X1 U911 ( .A(G137), .B(n1253), .ZN(G39) );
NAND2_X1 U912 ( .A1(KEYINPUT25), .A2(n1229), .ZN(n1253) );
AND3_X1 U913 ( .A1(n1254), .A2(n1252), .A3(n1243), .ZN(n1229) );
XNOR2_X1 U914 ( .A(G134), .B(n1255), .ZN(G36) );
NAND2_X1 U915 ( .A1(KEYINPUT36), .A2(n1231), .ZN(n1255) );
AND3_X1 U916 ( .A1(n1089), .A2(n1256), .A3(n1252), .ZN(n1231) );
XNOR2_X1 U917 ( .A(G131), .B(n1232), .ZN(G33) );
NAND2_X1 U918 ( .A1(n1252), .A2(n1222), .ZN(n1232) );
AND2_X1 U919 ( .A1(n1235), .A2(n1101), .ZN(n1252) );
NAND2_X1 U920 ( .A1(n1257), .A2(n1258), .ZN(n1101) );
OR2_X1 U921 ( .A1(n1245), .A2(KEYINPUT16), .ZN(n1258) );
NAND3_X1 U922 ( .A1(n1093), .A2(n1259), .A3(KEYINPUT16), .ZN(n1257) );
XNOR2_X1 U923 ( .A(G128), .B(n1260), .ZN(G30) );
NAND4_X1 U924 ( .A1(n1235), .A2(n1256), .A3(n1092), .A4(n1261), .ZN(n1260) );
XOR2_X1 U925 ( .A(KEYINPUT7), .B(n1243), .Z(n1261) );
INV_X1 U926 ( .A(n1098), .ZN(n1256) );
NOR3_X1 U927 ( .A1(n1262), .A2(n1084), .A3(n1085), .ZN(n1235) );
INV_X1 U928 ( .A(n1081), .ZN(n1085) );
XOR2_X1 U929 ( .A(G101), .B(n1263), .Z(G3) );
NOR3_X1 U930 ( .A1(n1224), .A2(n1264), .A3(n1218), .ZN(n1263) );
XNOR2_X1 U931 ( .A(n1254), .B(KEYINPUT45), .ZN(n1264) );
XNOR2_X1 U932 ( .A(G125), .B(n1265), .ZN(G27) );
NAND2_X1 U933 ( .A1(KEYINPUT33), .A2(n1126), .ZN(n1265) );
AND4_X1 U934 ( .A1(n1102), .A2(n1088), .A3(n1266), .A4(n1247), .ZN(n1126) );
INV_X1 U935 ( .A(n1099), .ZN(n1247) );
NOR2_X1 U936 ( .A1(n1262), .A2(n1245), .ZN(n1266) );
AND2_X1 U937 ( .A1(n1267), .A2(n1268), .ZN(n1262) );
NAND4_X1 U938 ( .A1(G953), .A2(G902), .A3(n1269), .A4(n1270), .ZN(n1268) );
INV_X1 U939 ( .A(G900), .ZN(n1270) );
XOR2_X1 U940 ( .A(n1068), .B(KEYINPUT50), .Z(n1267) );
XNOR2_X1 U941 ( .A(n1271), .B(n1219), .ZN(G24) );
NOR4_X1 U942 ( .A1(n1272), .A2(n1083), .A3(n1251), .A4(n1250), .ZN(n1219) );
NAND2_X1 U943 ( .A1(n1113), .A2(n1273), .ZN(n1083) );
XOR2_X1 U944 ( .A(G119), .B(n1217), .Z(G21) );
AND3_X1 U945 ( .A1(n1243), .A2(n1254), .A3(n1223), .ZN(n1217) );
INV_X1 U946 ( .A(n1072), .ZN(n1254) );
NOR2_X1 U947 ( .A1(n1273), .A2(n1113), .ZN(n1243) );
XOR2_X1 U948 ( .A(G116), .B(n1216), .Z(G18) );
NOR3_X1 U949 ( .A1(n1224), .A2(n1098), .A3(n1272), .ZN(n1216) );
NAND2_X1 U950 ( .A1(n1109), .A2(n1274), .ZN(n1098) );
XNOR2_X1 U951 ( .A(G113), .B(n1275), .ZN(G15) );
NAND3_X1 U952 ( .A1(n1276), .A2(n1277), .A3(n1222), .ZN(n1275) );
NOR2_X1 U953 ( .A1(n1224), .A2(n1099), .ZN(n1222) );
NAND2_X1 U954 ( .A1(n1251), .A2(n1278), .ZN(n1099) );
XNOR2_X1 U955 ( .A(KEYINPUT62), .B(n1250), .ZN(n1278) );
INV_X1 U956 ( .A(n1089), .ZN(n1224) );
NOR2_X1 U957 ( .A1(n1279), .A2(n1113), .ZN(n1089) );
INV_X1 U958 ( .A(n1280), .ZN(n1113) );
INV_X1 U959 ( .A(n1273), .ZN(n1279) );
OR2_X1 U960 ( .A1(n1223), .A2(KEYINPUT8), .ZN(n1277) );
INV_X1 U961 ( .A(n1272), .ZN(n1223) );
NAND3_X1 U962 ( .A1(n1092), .A2(n1281), .A3(n1102), .ZN(n1272) );
NAND2_X1 U963 ( .A1(KEYINPUT8), .A2(n1282), .ZN(n1276) );
NAND3_X1 U964 ( .A1(n1281), .A2(n1245), .A3(n1102), .ZN(n1282) );
NOR2_X1 U965 ( .A1(n1081), .A2(n1084), .ZN(n1102) );
INV_X1 U966 ( .A(n1080), .ZN(n1084) );
INV_X1 U967 ( .A(n1092), .ZN(n1245) );
XOR2_X1 U968 ( .A(G110), .B(n1215), .Z(G12) );
NOR3_X1 U969 ( .A1(n1072), .A2(n1218), .A3(n1283), .ZN(n1215) );
INV_X1 U970 ( .A(n1088), .ZN(n1283) );
NOR2_X1 U971 ( .A1(n1273), .A2(n1280), .ZN(n1088) );
XNOR2_X1 U972 ( .A(n1284), .B(G472), .ZN(n1280) );
NAND2_X1 U973 ( .A1(n1285), .A2(n1166), .ZN(n1284) );
XOR2_X1 U974 ( .A(n1286), .B(n1287), .Z(n1285) );
XNOR2_X1 U975 ( .A(n1181), .B(n1177), .ZN(n1287) );
NAND2_X1 U976 ( .A1(n1288), .A2(n1289), .ZN(n1177) );
NAND2_X1 U977 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
INV_X1 U978 ( .A(KEYINPUT42), .ZN(n1291) );
XNOR2_X1 U979 ( .A(G113), .B(n1292), .ZN(n1290) );
NAND2_X1 U980 ( .A1(KEYINPUT42), .A2(n1293), .ZN(n1288) );
XNOR2_X1 U981 ( .A(G113), .B(n1294), .ZN(n1293) );
NOR2_X1 U982 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U983 ( .A(n1297), .B(n1298), .ZN(n1286) );
NOR2_X1 U984 ( .A1(KEYINPUT18), .A2(n1178), .ZN(n1298) );
XNOR2_X1 U985 ( .A(n1299), .B(G146), .ZN(n1178) );
NOR2_X1 U986 ( .A1(KEYINPUT23), .A2(n1176), .ZN(n1297) );
XOR2_X1 U987 ( .A(n1300), .B(G101), .Z(n1176) );
NAND2_X1 U988 ( .A1(G210), .A2(n1301), .ZN(n1300) );
XOR2_X1 U989 ( .A(n1302), .B(n1118), .Z(n1273) );
NAND2_X1 U990 ( .A1(G217), .A2(n1303), .ZN(n1118) );
XNOR2_X1 U991 ( .A(n1119), .B(KEYINPUT55), .ZN(n1302) );
AND2_X1 U992 ( .A1(n1157), .A2(n1304), .ZN(n1119) );
XNOR2_X1 U993 ( .A(KEYINPUT6), .B(n1166), .ZN(n1304) );
XOR2_X1 U994 ( .A(n1305), .B(n1306), .Z(n1157) );
XOR2_X1 U995 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U996 ( .A(n1309), .B(n1310), .ZN(n1308) );
NAND2_X1 U997 ( .A1(KEYINPUT15), .A2(n1311), .ZN(n1309) );
XOR2_X1 U998 ( .A(n1312), .B(KEYINPUT29), .Z(n1307) );
NAND2_X1 U999 ( .A1(G221), .A2(n1313), .ZN(n1312) );
XNOR2_X1 U1000 ( .A(n1314), .B(n1315), .ZN(n1305) );
XNOR2_X1 U1001 ( .A(n1195), .B(n1295), .ZN(n1315) );
NAND4_X1 U1002 ( .A1(n1092), .A2(n1081), .A3(n1281), .A4(n1080), .ZN(n1218) );
NAND2_X1 U1003 ( .A1(G221), .A2(n1303), .ZN(n1080) );
NAND2_X1 U1004 ( .A1(G234), .A2(n1166), .ZN(n1303) );
NAND2_X1 U1005 ( .A1(n1068), .A2(n1316), .ZN(n1281) );
NAND3_X1 U1006 ( .A1(G902), .A2(n1269), .A3(n1148), .ZN(n1316) );
NOR2_X1 U1007 ( .A1(G898), .A2(n1132), .ZN(n1148) );
NAND3_X1 U1008 ( .A1(n1103), .A2(n1269), .A3(G952), .ZN(n1068) );
NAND2_X1 U1009 ( .A1(G237), .A2(G234), .ZN(n1269) );
XNOR2_X1 U1010 ( .A(n1132), .B(KEYINPUT28), .ZN(n1103) );
XNOR2_X1 U1011 ( .A(n1121), .B(G469), .ZN(n1081) );
NAND2_X1 U1012 ( .A1(n1317), .A2(n1166), .ZN(n1121) );
XOR2_X1 U1013 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1014 ( .A(n1181), .B(n1195), .ZN(n1319) );
XOR2_X1 U1015 ( .A(G110), .B(G140), .Z(n1195) );
XOR2_X1 U1016 ( .A(n1320), .B(KEYINPUT35), .Z(n1181) );
NAND3_X1 U1017 ( .A1(n1321), .A2(n1322), .A3(n1323), .ZN(n1320) );
NAND2_X1 U1018 ( .A1(n1144), .A2(n1139), .ZN(n1323) );
NAND2_X1 U1019 ( .A1(KEYINPUT32), .A2(n1324), .ZN(n1322) );
NAND2_X1 U1020 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XNOR2_X1 U1021 ( .A(KEYINPUT1), .B(n1139), .ZN(n1325) );
NAND2_X1 U1022 ( .A1(n1327), .A2(n1328), .ZN(n1321) );
INV_X1 U1023 ( .A(KEYINPUT32), .ZN(n1328) );
NAND2_X1 U1024 ( .A1(n1329), .A2(n1330), .ZN(n1327) );
OR3_X1 U1025 ( .A1(n1139), .A2(n1144), .A3(KEYINPUT1), .ZN(n1330) );
INV_X1 U1026 ( .A(n1326), .ZN(n1144) );
XNOR2_X1 U1027 ( .A(G134), .B(n1311), .ZN(n1326) );
INV_X1 U1028 ( .A(G137), .ZN(n1311) );
NAND2_X1 U1029 ( .A1(KEYINPUT1), .A2(n1139), .ZN(n1329) );
INV_X1 U1030 ( .A(G131), .ZN(n1139) );
XOR2_X1 U1031 ( .A(n1331), .B(n1190), .Z(n1318) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1132), .ZN(n1190) );
NAND2_X1 U1033 ( .A1(KEYINPUT44), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1034 ( .A(n1198), .B(n1141), .Z(n1332) );
XNOR2_X1 U1035 ( .A(n1310), .B(n1333), .ZN(n1141) );
NOR2_X1 U1036 ( .A1(KEYINPUT49), .A2(n1334), .ZN(n1333) );
XNOR2_X1 U1037 ( .A(n1335), .B(n1336), .ZN(n1334) );
NOR2_X1 U1038 ( .A1(G146), .A2(KEYINPUT19), .ZN(n1336) );
NOR2_X1 U1039 ( .A1(n1094), .A2(n1093), .ZN(n1092) );
NOR2_X1 U1040 ( .A1(n1337), .A2(n1116), .ZN(n1093) );
NOR2_X1 U1041 ( .A1(n1338), .A2(n1211), .ZN(n1116) );
XNOR2_X1 U1042 ( .A(KEYINPUT4), .B(n1115), .ZN(n1337) );
AND2_X1 U1043 ( .A1(n1211), .A2(n1338), .ZN(n1115) );
NAND4_X1 U1044 ( .A1(n1339), .A2(n1166), .A3(n1340), .A4(n1341), .ZN(n1338) );
NAND2_X1 U1045 ( .A1(KEYINPUT51), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1046 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XNOR2_X1 U1047 ( .A(KEYINPUT37), .B(n1206), .ZN(n1343) );
NAND2_X1 U1048 ( .A1(n1345), .A2(n1346), .ZN(n1340) );
INV_X1 U1049 ( .A(KEYINPUT51), .ZN(n1346) );
NAND2_X1 U1050 ( .A1(n1347), .A2(n1348), .ZN(n1345) );
NAND3_X1 U1051 ( .A1(KEYINPUT37), .A2(n1344), .A3(n1206), .ZN(n1348) );
OR2_X1 U1052 ( .A1(n1206), .A2(KEYINPUT37), .ZN(n1347) );
OR2_X1 U1053 ( .A1(n1344), .A2(n1206), .ZN(n1339) );
INV_X1 U1054 ( .A(n1149), .ZN(n1206) );
XNOR2_X1 U1055 ( .A(n1349), .B(n1350), .ZN(n1149) );
XOR2_X1 U1056 ( .A(n1351), .B(n1198), .Z(n1350) );
XOR2_X1 U1057 ( .A(G101), .B(n1352), .Z(n1198) );
XNOR2_X1 U1058 ( .A(n1059), .B(G104), .ZN(n1352) );
INV_X1 U1059 ( .A(G107), .ZN(n1059) );
NOR2_X1 U1060 ( .A1(G110), .A2(KEYINPUT2), .ZN(n1351) );
XOR2_X1 U1061 ( .A(n1353), .B(n1354), .Z(n1349) );
XNOR2_X1 U1062 ( .A(n1271), .B(G113), .ZN(n1354) );
NAND2_X1 U1063 ( .A1(KEYINPUT31), .A2(n1292), .ZN(n1353) );
XOR2_X1 U1064 ( .A(n1295), .B(n1296), .Z(n1292) );
XOR2_X1 U1065 ( .A(G116), .B(KEYINPUT46), .Z(n1296) );
XNOR2_X1 U1066 ( .A(G119), .B(KEYINPUT20), .ZN(n1295) );
XNOR2_X1 U1067 ( .A(n1208), .B(n1210), .ZN(n1344) );
XNOR2_X1 U1068 ( .A(n1299), .B(n1314), .ZN(n1210) );
XOR2_X1 U1069 ( .A(G125), .B(G146), .Z(n1314) );
XOR2_X1 U1070 ( .A(n1355), .B(n1356), .Z(n1299) );
NOR2_X1 U1071 ( .A1(KEYINPUT41), .A2(n1310), .ZN(n1356) );
XNOR2_X1 U1072 ( .A(G143), .B(KEYINPUT61), .ZN(n1355) );
NAND2_X1 U1073 ( .A1(G224), .A2(n1132), .ZN(n1208) );
AND2_X1 U1074 ( .A1(G210), .A2(n1357), .ZN(n1211) );
INV_X1 U1075 ( .A(n1259), .ZN(n1094) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1357), .ZN(n1259) );
NAND2_X1 U1077 ( .A1(n1166), .A2(n1358), .ZN(n1357) );
INV_X1 U1078 ( .A(G237), .ZN(n1358) );
NAND2_X1 U1079 ( .A1(n1251), .A2(n1274), .ZN(n1072) );
XNOR2_X1 U1080 ( .A(n1250), .B(KEYINPUT26), .ZN(n1274) );
INV_X1 U1081 ( .A(n1240), .ZN(n1250) );
XNOR2_X1 U1082 ( .A(n1105), .B(KEYINPUT14), .ZN(n1240) );
XOR2_X1 U1083 ( .A(n1359), .B(G475), .Z(n1105) );
NAND2_X1 U1084 ( .A1(n1170), .A2(n1166), .ZN(n1359) );
XNOR2_X1 U1085 ( .A(n1360), .B(n1361), .ZN(n1170) );
NOR2_X1 U1086 ( .A1(n1362), .A2(n1363), .ZN(n1361) );
NOR2_X1 U1087 ( .A1(n1364), .A2(n1365), .ZN(n1363) );
NOR2_X1 U1088 ( .A1(n1366), .A2(n1367), .ZN(n1364) );
NOR2_X1 U1089 ( .A1(G113), .A2(n1368), .ZN(n1367) );
NOR2_X1 U1090 ( .A1(n1171), .A2(n1369), .ZN(n1366) );
NOR2_X1 U1091 ( .A1(n1370), .A2(n1371), .ZN(n1362) );
NOR2_X1 U1092 ( .A1(n1372), .A2(n1373), .ZN(n1371) );
NOR2_X1 U1093 ( .A1(n1368), .A2(n1369), .ZN(n1373) );
INV_X1 U1094 ( .A(G113), .ZN(n1369) );
XNOR2_X1 U1095 ( .A(n1171), .B(KEYINPUT17), .ZN(n1368) );
NOR2_X1 U1096 ( .A1(G113), .A2(n1171), .ZN(n1372) );
INV_X1 U1097 ( .A(G104), .ZN(n1171) );
INV_X1 U1098 ( .A(n1365), .ZN(n1370) );
NAND2_X1 U1099 ( .A1(KEYINPUT5), .A2(n1271), .ZN(n1365) );
NAND2_X1 U1100 ( .A1(KEYINPUT43), .A2(n1374), .ZN(n1360) );
XOR2_X1 U1101 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1102 ( .A(n1377), .B(n1378), .Z(n1376) );
NAND2_X1 U1103 ( .A1(G214), .A2(n1301), .ZN(n1378) );
NOR2_X1 U1104 ( .A1(G953), .A2(G237), .ZN(n1301) );
NAND2_X1 U1105 ( .A1(n1379), .A2(n1380), .ZN(n1377) );
OR2_X1 U1106 ( .A1(n1381), .A2(G146), .ZN(n1380) );
XOR2_X1 U1107 ( .A(n1382), .B(KEYINPUT48), .Z(n1379) );
NAND2_X1 U1108 ( .A1(G146), .A2(n1381), .ZN(n1382) );
XOR2_X1 U1109 ( .A(n1137), .B(KEYINPUT10), .Z(n1381) );
XOR2_X1 U1110 ( .A(G125), .B(G140), .Z(n1137) );
XNOR2_X1 U1111 ( .A(n1335), .B(G131), .ZN(n1375) );
INV_X1 U1112 ( .A(n1109), .ZN(n1251) );
XNOR2_X1 U1113 ( .A(n1383), .B(G478), .ZN(n1109) );
NAND2_X1 U1114 ( .A1(n1162), .A2(n1166), .ZN(n1383) );
INV_X1 U1115 ( .A(G902), .ZN(n1166) );
XNOR2_X1 U1116 ( .A(n1384), .B(n1385), .ZN(n1162) );
XOR2_X1 U1117 ( .A(n1386), .B(n1387), .Z(n1385) );
XNOR2_X1 U1118 ( .A(n1388), .B(n1389), .ZN(n1387) );
NOR2_X1 U1119 ( .A1(KEYINPUT30), .A2(n1310), .ZN(n1389) );
XNOR2_X1 U1120 ( .A(G128), .B(KEYINPUT60), .ZN(n1310) );
NOR2_X1 U1121 ( .A1(KEYINPUT39), .A2(n1390), .ZN(n1388) );
XNOR2_X1 U1122 ( .A(G107), .B(n1391), .ZN(n1390) );
XNOR2_X1 U1123 ( .A(n1271), .B(G116), .ZN(n1391) );
INV_X1 U1124 ( .A(G122), .ZN(n1271) );
NAND2_X1 U1125 ( .A1(n1313), .A2(G217), .ZN(n1386) );
AND2_X1 U1126 ( .A1(G234), .A2(n1132), .ZN(n1313) );
INV_X1 U1127 ( .A(G953), .ZN(n1132) );
XNOR2_X1 U1128 ( .A(G134), .B(n1392), .ZN(n1384) );
XNOR2_X1 U1129 ( .A(KEYINPUT21), .B(n1335), .ZN(n1392) );
INV_X1 U1130 ( .A(G143), .ZN(n1335) );
endmodule


