//Key = 1101101010001010010011110110010001000111100011011100111101010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304;

XOR2_X1 U735 ( .A(n1001), .B(n1002), .Z(G9) );
NAND4_X1 U736 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1002) );
NOR2_X1 U737 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
XOR2_X1 U738 ( .A(KEYINPUT25), .B(n1009), .Z(n1008) );
NOR2_X1 U739 ( .A1(n1010), .A2(n1011), .ZN(G75) );
NOR4_X1 U740 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
XOR2_X1 U741 ( .A(KEYINPUT52), .B(n1016), .Z(n1013) );
NOR2_X1 U742 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR4_X1 U743 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1018) );
NOR2_X1 U744 ( .A1(n1023), .A2(n1024), .ZN(n1019) );
NOR3_X1 U745 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
XOR2_X1 U746 ( .A(KEYINPUT1), .B(n1028), .Z(n1026) );
NOR3_X1 U747 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1023) );
AND2_X1 U748 ( .A1(n1032), .A2(n1033), .ZN(n1017) );
NAND4_X1 U749 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1012) );
NAND3_X1 U750 ( .A1(n1038), .A2(n1005), .A3(n1033), .ZN(n1035) );
NOR3_X1 U751 ( .A1(n1027), .A2(n1031), .A3(n1022), .ZN(n1033) );
NAND3_X1 U752 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1034) );
INV_X1 U753 ( .A(n1022), .ZN(n1041) );
NAND2_X1 U754 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NAND3_X1 U755 ( .A1(n1005), .A2(n1003), .A3(n1044), .ZN(n1043) );
NAND2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1042) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U759 ( .A1(n1005), .A2(n1009), .ZN(n1047) );
NOR3_X1 U760 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1010) );
INV_X1 U761 ( .A(n1036), .ZN(n1051) );
NAND4_X1 U762 ( .A1(n1052), .A2(n1039), .A3(n1053), .A4(n1054), .ZN(n1036) );
NOR4_X1 U763 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
XOR2_X1 U764 ( .A(n1059), .B(n1060), .Z(n1058) );
NOR2_X1 U765 ( .A1(n1061), .A2(KEYINPUT15), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1062), .A2(n1063), .ZN(n1057) );
INV_X1 U767 ( .A(n1025), .ZN(n1055) );
NOR2_X1 U768 ( .A1(n1064), .A2(n1065), .ZN(n1053) );
XOR2_X1 U769 ( .A(n1066), .B(KEYINPUT8), .Z(n1065) );
NAND2_X1 U770 ( .A1(n1062), .A2(n1063), .ZN(n1066) );
XNOR2_X1 U771 ( .A(n1067), .B(n1068), .ZN(n1064) );
XOR2_X1 U772 ( .A(KEYINPUT54), .B(G472), .Z(n1068) );
XOR2_X1 U773 ( .A(n1069), .B(n1070), .Z(G72) );
NOR2_X1 U774 ( .A1(n1071), .A2(n1037), .ZN(n1070) );
NOR2_X1 U775 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U776 ( .A1(n1074), .A2(n1075), .ZN(n1069) );
NAND2_X1 U777 ( .A1(n1076), .A2(n1037), .ZN(n1075) );
XNOR2_X1 U778 ( .A(n1014), .B(n1077), .ZN(n1076) );
OR3_X1 U779 ( .A1(n1073), .A2(n1077), .A3(n1037), .ZN(n1074) );
XNOR2_X1 U780 ( .A(n1078), .B(n1079), .ZN(n1077) );
XOR2_X1 U781 ( .A(n1080), .B(n1081), .Z(n1079) );
XOR2_X1 U782 ( .A(n1082), .B(n1083), .Z(n1078) );
XOR2_X1 U783 ( .A(n1084), .B(n1085), .Z(n1083) );
NAND2_X1 U784 ( .A1(KEYINPUT44), .A2(G125), .ZN(n1085) );
XOR2_X1 U785 ( .A(n1086), .B(n1087), .Z(G69) );
NAND2_X1 U786 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1088) );
NAND3_X1 U788 ( .A1(KEYINPUT23), .A2(n1089), .A3(n1090), .ZN(n1086) );
XNOR2_X1 U789 ( .A(n1091), .B(n1015), .ZN(n1090) );
NAND2_X1 U790 ( .A1(KEYINPUT4), .A2(n1092), .ZN(n1091) );
XOR2_X1 U791 ( .A(n1093), .B(n1094), .Z(n1092) );
NAND2_X1 U792 ( .A1(G953), .A2(n1095), .ZN(n1089) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XOR2_X1 U794 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NOR2_X1 U796 ( .A1(n1096), .A2(n1102), .ZN(G63) );
XOR2_X1 U797 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U798 ( .A1(KEYINPUT36), .A2(n1105), .ZN(n1104) );
NAND2_X1 U799 ( .A1(n1106), .A2(G478), .ZN(n1103) );
NOR2_X1 U800 ( .A1(n1096), .A2(n1107), .ZN(G60) );
NOR2_X1 U801 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U802 ( .A(n1110), .B(n1111), .Z(n1109) );
AND2_X1 U803 ( .A1(G475), .A2(n1106), .ZN(n1111) );
NOR2_X1 U804 ( .A1(KEYINPUT35), .A2(n1112), .ZN(n1110) );
AND2_X1 U805 ( .A1(n1112), .A2(KEYINPUT35), .ZN(n1108) );
XOR2_X1 U806 ( .A(n1113), .B(n1114), .Z(G6) );
NOR2_X1 U807 ( .A1(n1096), .A2(n1115), .ZN(G57) );
NOR2_X1 U808 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
XOR2_X1 U809 ( .A(KEYINPUT16), .B(n1118), .Z(n1117) );
NOR2_X1 U810 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XNOR2_X1 U811 ( .A(n1121), .B(KEYINPUT11), .ZN(n1120) );
INV_X1 U812 ( .A(n1122), .ZN(n1119) );
NOR2_X1 U813 ( .A1(n1121), .A2(n1122), .ZN(n1116) );
NAND2_X1 U814 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XNOR2_X1 U815 ( .A(n1125), .B(n1126), .ZN(n1121) );
XOR2_X1 U816 ( .A(n1127), .B(n1128), .Z(n1125) );
NOR2_X1 U817 ( .A1(n1129), .A2(n1101), .ZN(n1128) );
NAND2_X1 U818 ( .A1(n1130), .A2(KEYINPUT12), .ZN(n1127) );
XOR2_X1 U819 ( .A(n1131), .B(KEYINPUT10), .Z(n1130) );
NOR2_X1 U820 ( .A1(n1096), .A2(n1132), .ZN(G54) );
XOR2_X1 U821 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U822 ( .A1(KEYINPUT50), .A2(n1135), .ZN(n1134) );
XOR2_X1 U823 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U824 ( .A(n1138), .B(n1139), .Z(n1137) );
XNOR2_X1 U825 ( .A(KEYINPUT9), .B(n1140), .ZN(n1139) );
NOR2_X1 U826 ( .A1(KEYINPUT61), .A2(n1141), .ZN(n1140) );
XOR2_X1 U827 ( .A(G131), .B(n1142), .Z(n1141) );
XOR2_X1 U828 ( .A(n1143), .B(n1144), .Z(n1136) );
NAND2_X1 U829 ( .A1(n1106), .A2(G469), .ZN(n1133) );
NOR2_X1 U830 ( .A1(n1096), .A2(n1145), .ZN(G51) );
XOR2_X1 U831 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U832 ( .A1(KEYINPUT60), .A2(n1148), .ZN(n1147) );
NOR2_X1 U833 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XOR2_X1 U834 ( .A(n1151), .B(KEYINPUT57), .Z(n1150) );
NAND2_X1 U835 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U836 ( .A(n1154), .B(KEYINPUT30), .Z(n1152) );
NOR2_X1 U837 ( .A1(n1154), .A2(n1153), .ZN(n1149) );
XOR2_X1 U838 ( .A(n1155), .B(n1156), .Z(n1153) );
XNOR2_X1 U839 ( .A(n1157), .B(KEYINPUT13), .ZN(n1156) );
NAND2_X1 U840 ( .A1(KEYINPUT37), .A2(n1158), .ZN(n1157) );
NAND2_X1 U841 ( .A1(n1106), .A2(n1061), .ZN(n1146) );
INV_X1 U842 ( .A(n1101), .ZN(n1106) );
NAND2_X1 U843 ( .A1(G902), .A2(n1159), .ZN(n1101) );
OR2_X1 U844 ( .A1(n1015), .A2(n1014), .ZN(n1159) );
NAND4_X1 U845 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1014) );
NOR4_X1 U846 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
NAND3_X1 U847 ( .A1(n1009), .A2(n1168), .A3(n1169), .ZN(n1162) );
OR2_X1 U848 ( .A1(n1038), .A2(n1170), .ZN(n1168) );
NAND4_X1 U849 ( .A1(n1171), .A2(n1114), .A3(n1172), .A4(n1173), .ZN(n1015) );
AND4_X1 U850 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
NAND2_X1 U851 ( .A1(n1178), .A2(n1032), .ZN(n1172) );
NAND2_X1 U852 ( .A1(n1179), .A2(n1180), .ZN(n1032) );
NAND3_X1 U853 ( .A1(n1039), .A2(n1181), .A3(n1182), .ZN(n1180) );
NAND2_X1 U854 ( .A1(n1170), .A2(n1005), .ZN(n1179) );
NAND3_X1 U855 ( .A1(n1178), .A2(n1005), .A3(n1038), .ZN(n1114) );
INV_X1 U856 ( .A(n1020), .ZN(n1005) );
NAND3_X1 U857 ( .A1(n1183), .A2(n1184), .A3(n1038), .ZN(n1171) );
XOR2_X1 U858 ( .A(KEYINPUT2), .B(n1045), .Z(n1184) );
NOR2_X1 U859 ( .A1(n1037), .A2(G952), .ZN(n1096) );
XNOR2_X1 U860 ( .A(G146), .B(n1185), .ZN(G48) );
NAND4_X1 U861 ( .A1(KEYINPUT17), .A2(n1169), .A3(n1038), .A4(n1009), .ZN(n1185) );
XOR2_X1 U862 ( .A(n1160), .B(n1186), .Z(G45) );
NOR2_X1 U863 ( .A1(G143), .A2(KEYINPUT7), .ZN(n1186) );
NAND3_X1 U864 ( .A1(n1187), .A2(n1009), .A3(n1188), .ZN(n1160) );
NOR3_X1 U865 ( .A1(n1189), .A2(n1182), .A3(n1190), .ZN(n1188) );
XNOR2_X1 U866 ( .A(G140), .B(n1161), .ZN(G42) );
NAND3_X1 U867 ( .A1(n1044), .A2(n1003), .A3(n1191), .ZN(n1161) );
XOR2_X1 U868 ( .A(n1166), .B(n1192), .Z(G39) );
NOR2_X1 U869 ( .A1(KEYINPUT34), .A2(n1193), .ZN(n1192) );
AND3_X1 U870 ( .A1(n1044), .A2(n1039), .A3(n1169), .ZN(n1166) );
XNOR2_X1 U871 ( .A(n1165), .B(n1194), .ZN(G36) );
XOR2_X1 U872 ( .A(KEYINPUT39), .B(G134), .Z(n1194) );
AND3_X1 U873 ( .A1(n1187), .A2(n1170), .A3(n1049), .ZN(n1165) );
XOR2_X1 U874 ( .A(n1195), .B(n1196), .Z(G33) );
XNOR2_X1 U875 ( .A(G131), .B(KEYINPUT27), .ZN(n1196) );
NAND2_X1 U876 ( .A1(KEYINPUT45), .A2(n1164), .ZN(n1195) );
AND3_X1 U877 ( .A1(n1187), .A2(n1038), .A3(n1049), .ZN(n1164) );
NOR2_X1 U878 ( .A1(n1027), .A2(n1182), .ZN(n1049) );
INV_X1 U879 ( .A(n1044), .ZN(n1027) );
NOR2_X1 U880 ( .A1(n1030), .A2(n1056), .ZN(n1044) );
INV_X1 U881 ( .A(n1029), .ZN(n1056) );
XNOR2_X1 U882 ( .A(n1197), .B(KEYINPUT47), .ZN(n1030) );
XOR2_X1 U883 ( .A(G128), .B(n1198), .Z(G30) );
NOR2_X1 U884 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U885 ( .A(n1201), .B(KEYINPUT24), .Z(n1199) );
NAND2_X1 U886 ( .A1(n1169), .A2(n1170), .ZN(n1201) );
AND2_X1 U887 ( .A1(n1187), .A2(n1182), .ZN(n1169) );
AND3_X1 U888 ( .A1(n1003), .A2(n1202), .A3(n1050), .ZN(n1187) );
XNOR2_X1 U889 ( .A(G101), .B(n1176), .ZN(G3) );
NAND3_X1 U890 ( .A1(n1039), .A2(n1003), .A3(n1183), .ZN(n1176) );
XOR2_X1 U891 ( .A(G125), .B(n1167), .Z(G27) );
AND3_X1 U892 ( .A1(n1045), .A2(n1009), .A3(n1191), .ZN(n1167) );
AND4_X1 U893 ( .A1(n1182), .A2(n1038), .A3(n1181), .A4(n1202), .ZN(n1191) );
NAND2_X1 U894 ( .A1(n1022), .A2(n1203), .ZN(n1202) );
NAND4_X1 U895 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1073), .ZN(n1203) );
INV_X1 U896 ( .A(G900), .ZN(n1073) );
XNOR2_X1 U897 ( .A(G122), .B(n1175), .ZN(G24) );
NAND3_X1 U898 ( .A1(n1045), .A2(n1205), .A3(n1206), .ZN(n1175) );
NOR3_X1 U899 ( .A1(n1020), .A2(n1190), .A3(n1189), .ZN(n1206) );
NAND2_X1 U900 ( .A1(n1207), .A2(n1181), .ZN(n1020) );
XNOR2_X1 U901 ( .A(G119), .B(n1174), .ZN(G21) );
NAND3_X1 U902 ( .A1(n1045), .A2(n1205), .A3(n1208), .ZN(n1174) );
NOR3_X1 U903 ( .A1(n1181), .A2(n1021), .A3(n1207), .ZN(n1208) );
XOR2_X1 U904 ( .A(n1209), .B(G116), .Z(G18) );
NAND2_X1 U905 ( .A1(KEYINPUT26), .A2(n1177), .ZN(n1209) );
NAND3_X1 U906 ( .A1(n1045), .A2(n1170), .A3(n1183), .ZN(n1177) );
INV_X1 U907 ( .A(n1007), .ZN(n1170) );
NAND2_X1 U908 ( .A1(n1190), .A2(n1210), .ZN(n1007) );
INV_X1 U909 ( .A(n1031), .ZN(n1045) );
XOR2_X1 U910 ( .A(n1211), .B(n1212), .Z(G15) );
NAND3_X1 U911 ( .A1(n1038), .A2(n1183), .A3(n1213), .ZN(n1212) );
XOR2_X1 U912 ( .A(n1031), .B(KEYINPUT29), .Z(n1213) );
NAND2_X1 U913 ( .A1(n1214), .A2(n1025), .ZN(n1031) );
XOR2_X1 U914 ( .A(KEYINPUT1), .B(n1215), .Z(n1214) );
AND3_X1 U915 ( .A1(n1050), .A2(n1207), .A3(n1205), .ZN(n1183) );
INV_X1 U916 ( .A(n1182), .ZN(n1207) );
NOR2_X1 U917 ( .A1(n1210), .A2(n1190), .ZN(n1038) );
INV_X1 U918 ( .A(n1189), .ZN(n1210) );
XNOR2_X1 U919 ( .A(G110), .B(n1216), .ZN(G12) );
NAND4_X1 U920 ( .A1(n1182), .A2(n1178), .A3(n1217), .A4(n1181), .ZN(n1216) );
INV_X1 U921 ( .A(n1050), .ZN(n1181) );
XOR2_X1 U922 ( .A(n1129), .B(n1218), .Z(n1050) );
NOR2_X1 U923 ( .A1(n1067), .A2(KEYINPUT5), .ZN(n1218) );
AND2_X1 U924 ( .A1(n1219), .A2(n1220), .ZN(n1067) );
XOR2_X1 U925 ( .A(n1221), .B(n1126), .Z(n1219) );
XNOR2_X1 U926 ( .A(n1222), .B(n1223), .ZN(n1126) );
XOR2_X1 U927 ( .A(n1224), .B(n1225), .Z(n1221) );
INV_X1 U928 ( .A(n1131), .ZN(n1225) );
NAND2_X1 U929 ( .A1(n1226), .A2(n1124), .ZN(n1224) );
NAND2_X1 U930 ( .A1(G101), .A2(n1227), .ZN(n1124) );
XOR2_X1 U931 ( .A(n1123), .B(KEYINPUT41), .Z(n1226) );
OR2_X1 U932 ( .A1(G101), .A2(n1227), .ZN(n1123) );
AND3_X1 U933 ( .A1(n1228), .A2(n1037), .A3(G210), .ZN(n1227) );
INV_X1 U934 ( .A(G472), .ZN(n1129) );
XOR2_X1 U935 ( .A(KEYINPUT42), .B(n1039), .Z(n1217) );
INV_X1 U936 ( .A(n1021), .ZN(n1039) );
NAND2_X1 U937 ( .A1(n1189), .A2(n1190), .ZN(n1021) );
XOR2_X1 U938 ( .A(n1229), .B(G475), .Z(n1190) );
OR2_X1 U939 ( .A1(n1112), .A2(G902), .ZN(n1229) );
XOR2_X1 U940 ( .A(n1230), .B(n1231), .Z(n1112) );
XOR2_X1 U941 ( .A(G113), .B(n1232), .Z(n1231) );
XOR2_X1 U942 ( .A(G131), .B(G122), .Z(n1232) );
XOR2_X1 U943 ( .A(n1233), .B(n1234), .Z(n1230) );
NOR2_X1 U944 ( .A1(KEYINPUT51), .A2(n1235), .ZN(n1234) );
XOR2_X1 U945 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND4_X1 U946 ( .A1(KEYINPUT49), .A2(G214), .A3(n1228), .A4(n1037), .ZN(n1237) );
XOR2_X1 U947 ( .A(n1113), .B(n1238), .Z(n1233) );
NOR2_X1 U948 ( .A1(KEYINPUT31), .A2(n1239), .ZN(n1238) );
XOR2_X1 U949 ( .A(n1240), .B(n1241), .Z(n1239) );
XOR2_X1 U950 ( .A(KEYINPUT58), .B(G146), .Z(n1241) );
NAND2_X1 U951 ( .A1(KEYINPUT20), .A2(n1242), .ZN(n1240) );
XOR2_X1 U952 ( .A(G125), .B(n1243), .Z(n1242) );
XOR2_X1 U953 ( .A(KEYINPUT14), .B(G140), .Z(n1243) );
INV_X1 U954 ( .A(G104), .ZN(n1113) );
XOR2_X1 U955 ( .A(n1244), .B(G478), .Z(n1189) );
OR2_X1 U956 ( .A1(n1105), .A2(G902), .ZN(n1244) );
XOR2_X1 U957 ( .A(n1245), .B(n1246), .Z(n1105) );
XOR2_X1 U958 ( .A(n1082), .B(n1247), .Z(n1246) );
XOR2_X1 U959 ( .A(n1248), .B(n1249), .Z(n1247) );
AND3_X1 U960 ( .A1(G234), .A2(n1037), .A3(G217), .ZN(n1249) );
NAND2_X1 U961 ( .A1(KEYINPUT33), .A2(n1236), .ZN(n1248) );
XOR2_X1 U962 ( .A(n1250), .B(n1251), .Z(n1245) );
XOR2_X1 U963 ( .A(G128), .B(G122), .Z(n1251) );
XOR2_X1 U964 ( .A(G116), .B(n1001), .Z(n1250) );
AND2_X1 U965 ( .A1(n1205), .A2(n1003), .ZN(n1178) );
AND2_X1 U966 ( .A1(n1252), .A2(n1025), .ZN(n1003) );
NAND2_X1 U967 ( .A1(G221), .A2(n1253), .ZN(n1025) );
XOR2_X1 U968 ( .A(KEYINPUT18), .B(n1215), .Z(n1252) );
INV_X1 U969 ( .A(n1028), .ZN(n1215) );
XNOR2_X1 U970 ( .A(n1254), .B(n1062), .ZN(n1028) );
XNOR2_X1 U971 ( .A(G469), .B(KEYINPUT59), .ZN(n1062) );
NAND2_X1 U972 ( .A1(KEYINPUT21), .A2(n1063), .ZN(n1254) );
NAND2_X1 U973 ( .A1(n1220), .A2(n1255), .ZN(n1063) );
NAND2_X1 U974 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
NAND2_X1 U975 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U976 ( .A(n1260), .B(n1261), .Z(n1259) );
INV_X1 U977 ( .A(n1138), .ZN(n1261) );
XOR2_X1 U978 ( .A(n1222), .B(n1144), .Z(n1258) );
XOR2_X1 U979 ( .A(n1262), .B(KEYINPUT56), .Z(n1256) );
NAND2_X1 U980 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U981 ( .A(n1260), .B(n1138), .Z(n1264) );
XNOR2_X1 U982 ( .A(G140), .B(n1265), .ZN(n1138) );
NOR2_X1 U983 ( .A1(G953), .A2(n1072), .ZN(n1265) );
INV_X1 U984 ( .A(G227), .ZN(n1072) );
OR2_X1 U985 ( .A1(G110), .A2(KEYINPUT43), .ZN(n1260) );
XOR2_X1 U986 ( .A(n1222), .B(n1266), .Z(n1263) );
INV_X1 U987 ( .A(n1144), .ZN(n1266) );
XNOR2_X1 U988 ( .A(n1267), .B(n1084), .ZN(n1144) );
NAND2_X1 U989 ( .A1(n1268), .A2(n1269), .ZN(n1084) );
NAND2_X1 U990 ( .A1(G146), .A2(n1236), .ZN(n1269) );
XOR2_X1 U991 ( .A(KEYINPUT63), .B(n1270), .Z(n1268) );
NOR2_X1 U992 ( .A1(G146), .A2(n1236), .ZN(n1270) );
INV_X1 U993 ( .A(G143), .ZN(n1236) );
NAND2_X1 U994 ( .A1(n1271), .A2(n1272), .ZN(n1267) );
NAND2_X1 U995 ( .A1(n1273), .A2(G101), .ZN(n1272) );
INV_X1 U996 ( .A(n1274), .ZN(n1273) );
NAND2_X1 U997 ( .A1(n1275), .A2(n1274), .ZN(n1271) );
XOR2_X1 U998 ( .A(n1276), .B(G104), .Z(n1274) );
NAND2_X1 U999 ( .A1(KEYINPUT62), .A2(n1001), .ZN(n1276) );
INV_X1 U1000 ( .A(G107), .ZN(n1001) );
XNOR2_X1 U1001 ( .A(G101), .B(KEYINPUT32), .ZN(n1275) );
XNOR2_X1 U1002 ( .A(n1080), .B(n1142), .ZN(n1222) );
XNOR2_X1 U1003 ( .A(n1277), .B(KEYINPUT28), .ZN(n1142) );
NAND2_X1 U1004 ( .A1(n1278), .A2(KEYINPUT40), .ZN(n1277) );
XOR2_X1 U1005 ( .A(n1279), .B(n1280), .Z(n1278) );
INV_X1 U1006 ( .A(n1082), .ZN(n1280) );
XNOR2_X1 U1007 ( .A(G134), .B(KEYINPUT48), .ZN(n1082) );
NAND2_X1 U1008 ( .A1(n1281), .A2(n1193), .ZN(n1279) );
INV_X1 U1009 ( .A(G137), .ZN(n1193) );
XNOR2_X1 U1010 ( .A(KEYINPUT53), .B(KEYINPUT22), .ZN(n1281) );
XOR2_X1 U1011 ( .A(G128), .B(G131), .Z(n1080) );
AND2_X1 U1012 ( .A1(n1009), .A2(n1004), .ZN(n1205) );
NAND2_X1 U1013 ( .A1(n1022), .A2(n1282), .ZN(n1004) );
NAND4_X1 U1014 ( .A1(G953), .A2(G902), .A3(n1204), .A4(n1095), .ZN(n1282) );
INV_X1 U1015 ( .A(G898), .ZN(n1095) );
NAND3_X1 U1016 ( .A1(n1204), .A2(n1037), .A3(G952), .ZN(n1022) );
NAND2_X1 U1017 ( .A1(G237), .A2(G234), .ZN(n1204) );
INV_X1 U1018 ( .A(n1200), .ZN(n1009) );
NAND2_X1 U1019 ( .A1(n1197), .A2(n1029), .ZN(n1200) );
NAND2_X1 U1020 ( .A1(G214), .A2(n1283), .ZN(n1029) );
XNOR2_X1 U1021 ( .A(n1059), .B(n1061), .ZN(n1197) );
AND2_X1 U1022 ( .A1(G210), .A2(n1283), .ZN(n1061) );
NAND2_X1 U1023 ( .A1(n1228), .A2(n1220), .ZN(n1283) );
INV_X1 U1024 ( .A(G237), .ZN(n1228) );
NAND2_X1 U1025 ( .A1(n1284), .A2(n1220), .ZN(n1059) );
XOR2_X1 U1026 ( .A(n1285), .B(n1286), .Z(n1284) );
INV_X1 U1027 ( .A(n1154), .ZN(n1286) );
XOR2_X1 U1028 ( .A(n1287), .B(n1288), .Z(n1154) );
INV_X1 U1029 ( .A(n1093), .ZN(n1288) );
XOR2_X1 U1030 ( .A(n1289), .B(n1290), .Z(n1093) );
XOR2_X1 U1031 ( .A(G104), .B(n1291), .Z(n1290) );
XOR2_X1 U1032 ( .A(KEYINPUT0), .B(G107), .Z(n1291) );
XOR2_X1 U1033 ( .A(n1131), .B(G101), .Z(n1289) );
XOR2_X1 U1034 ( .A(n1211), .B(n1292), .Z(n1131) );
XOR2_X1 U1035 ( .A(G119), .B(G116), .Z(n1292) );
INV_X1 U1036 ( .A(G113), .ZN(n1211) );
NAND2_X1 U1037 ( .A1(KEYINPUT55), .A2(n1094), .ZN(n1287) );
XNOR2_X1 U1038 ( .A(G110), .B(G122), .ZN(n1094) );
NAND2_X1 U1039 ( .A1(n1293), .A2(KEYINPUT3), .ZN(n1285) );
XNOR2_X1 U1040 ( .A(n1155), .B(n1158), .ZN(n1293) );
XNOR2_X1 U1041 ( .A(G128), .B(n1223), .ZN(n1158) );
NOR2_X1 U1042 ( .A1(KEYINPUT19), .A2(n1294), .ZN(n1223) );
XOR2_X1 U1043 ( .A(G143), .B(n1295), .Z(n1294) );
NOR2_X1 U1044 ( .A1(G146), .A2(KEYINPUT46), .ZN(n1295) );
XOR2_X1 U1045 ( .A(n1296), .B(n1297), .Z(n1155) );
AND2_X1 U1046 ( .A1(n1037), .A2(G224), .ZN(n1297) );
INV_X1 U1047 ( .A(G125), .ZN(n1296) );
XOR2_X1 U1048 ( .A(n1052), .B(KEYINPUT6), .Z(n1182) );
XNOR2_X1 U1049 ( .A(n1298), .B(n1100), .ZN(n1052) );
NAND2_X1 U1050 ( .A1(G217), .A2(n1253), .ZN(n1100) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1220), .ZN(n1253) );
INV_X1 U1052 ( .A(G902), .ZN(n1220) );
OR2_X1 U1053 ( .A1(n1099), .A2(G902), .ZN(n1298) );
XNOR2_X1 U1054 ( .A(n1299), .B(n1300), .ZN(n1099) );
XOR2_X1 U1055 ( .A(n1301), .B(n1302), .Z(n1300) );
XOR2_X1 U1056 ( .A(G125), .B(G119), .Z(n1302) );
XOR2_X1 U1057 ( .A(KEYINPUT38), .B(G146), .Z(n1301) );
XOR2_X1 U1058 ( .A(n1303), .B(n1081), .Z(n1299) );
XOR2_X1 U1059 ( .A(G137), .B(G140), .Z(n1081) );
XOR2_X1 U1060 ( .A(n1304), .B(n1143), .Z(n1303) );
XOR2_X1 U1061 ( .A(G110), .B(G128), .Z(n1143) );
NAND3_X1 U1062 ( .A1(G234), .A2(n1037), .A3(G221), .ZN(n1304) );
INV_X1 U1063 ( .A(G953), .ZN(n1037) );
endmodule


