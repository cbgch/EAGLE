//Key = 0100100011100100011110000010110001011010110011111111000011001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;

XOR2_X1 U701 ( .A(n963), .B(n964), .Z(G9) );
NOR2_X1 U702 ( .A1(G107), .A2(KEYINPUT24), .ZN(n964) );
NAND4_X1 U703 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(n963) );
XNOR2_X1 U704 ( .A(KEYINPUT19), .B(n969), .ZN(n968) );
NOR2_X1 U705 ( .A1(n970), .A2(n971), .ZN(G75) );
NOR4_X1 U706 ( .A1(G953), .A2(n972), .A3(n973), .A4(n974), .ZN(n971) );
NOR2_X1 U707 ( .A1(n975), .A2(n976), .ZN(n973) );
NOR2_X1 U708 ( .A1(n977), .A2(n978), .ZN(n975) );
NOR3_X1 U709 ( .A1(n979), .A2(n980), .A3(n981), .ZN(n978) );
NOR2_X1 U710 ( .A1(n982), .A2(n983), .ZN(n980) );
NOR2_X1 U711 ( .A1(n984), .A2(n985), .ZN(n983) );
NOR2_X1 U712 ( .A1(n986), .A2(n987), .ZN(n984) );
NOR2_X1 U713 ( .A1(n988), .A2(n989), .ZN(n986) );
NOR2_X1 U714 ( .A1(n990), .A2(n991), .ZN(n982) );
NOR2_X1 U715 ( .A1(n965), .A2(n992), .ZN(n990) );
NOR3_X1 U716 ( .A1(n985), .A2(n993), .A3(n991), .ZN(n977) );
INV_X1 U717 ( .A(n994), .ZN(n991) );
NOR2_X1 U718 ( .A1(n995), .A2(n996), .ZN(n993) );
NOR2_X1 U719 ( .A1(n997), .A2(n981), .ZN(n996) );
NOR2_X1 U720 ( .A1(n998), .A2(n999), .ZN(n997) );
NOR2_X1 U721 ( .A1(n1000), .A2(n1001), .ZN(n998) );
XOR2_X1 U722 ( .A(KEYINPUT42), .B(n1002), .Z(n1001) );
NOR2_X1 U723 ( .A1(n1003), .A2(n979), .ZN(n995) );
NOR2_X1 U724 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NOR3_X1 U725 ( .A1(n972), .A2(G953), .A3(G952), .ZN(n970) );
AND4_X1 U726 ( .A1(n1006), .A2(n994), .A3(n1007), .A4(n1008), .ZN(n972) );
NOR3_X1 U727 ( .A1(n979), .A2(n1009), .A3(n1010), .ZN(n1008) );
XNOR2_X1 U728 ( .A(n1011), .B(n1012), .ZN(n1009) );
NOR2_X1 U729 ( .A1(KEYINPUT15), .A2(n1013), .ZN(n1012) );
INV_X1 U730 ( .A(n1014), .ZN(n979) );
XNOR2_X1 U731 ( .A(n1015), .B(G472), .ZN(n1007) );
XNOR2_X1 U732 ( .A(n1016), .B(n1017), .ZN(n1006) );
XOR2_X1 U733 ( .A(n1018), .B(n1019), .Z(G72) );
XOR2_X1 U734 ( .A(n1020), .B(n1021), .Z(n1019) );
NAND2_X1 U735 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND3_X1 U736 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
XNOR2_X1 U737 ( .A(KEYINPUT10), .B(n1027), .ZN(n1024) );
NAND2_X1 U738 ( .A1(n1028), .A2(n1029), .ZN(n1020) );
NAND2_X1 U739 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
XNOR2_X1 U740 ( .A(KEYINPUT11), .B(n1022), .ZN(n1030) );
XOR2_X1 U741 ( .A(n1032), .B(n1033), .Z(n1028) );
XOR2_X1 U742 ( .A(n1034), .B(n1035), .Z(n1033) );
XNOR2_X1 U743 ( .A(n1036), .B(n1037), .ZN(n1034) );
XOR2_X1 U744 ( .A(n1038), .B(n1039), .Z(n1032) );
NOR2_X1 U745 ( .A1(G134), .A2(KEYINPUT31), .ZN(n1039) );
XNOR2_X1 U746 ( .A(KEYINPUT6), .B(KEYINPUT47), .ZN(n1038) );
NOR2_X1 U747 ( .A1(n1040), .A2(n1022), .ZN(n1018) );
AND2_X1 U748 ( .A1(G227), .A2(G900), .ZN(n1040) );
NAND2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(G69) );
NAND2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U751 ( .A1(n1045), .A2(n1046), .ZN(n1041) );
INV_X1 U752 ( .A(n1043), .ZN(n1046) );
NOR2_X1 U753 ( .A1(KEYINPUT0), .A2(n1047), .ZN(n1043) );
XOR2_X1 U754 ( .A(n1048), .B(n1049), .Z(n1047) );
NOR2_X1 U755 ( .A1(n1050), .A2(G953), .ZN(n1049) );
NAND2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1048) );
XOR2_X1 U757 ( .A(n1053), .B(KEYINPUT1), .Z(n1051) );
NAND2_X1 U758 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U759 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
XOR2_X1 U760 ( .A(KEYINPUT37), .B(n1058), .Z(n1056) );
NAND2_X1 U761 ( .A1(n1052), .A2(n1044), .ZN(n1045) );
NAND2_X1 U762 ( .A1(G953), .A2(n1059), .ZN(n1044) );
INV_X1 U763 ( .A(G224), .ZN(n1059) );
OR2_X1 U764 ( .A1(n1022), .A2(G898), .ZN(n1052) );
NOR2_X1 U765 ( .A1(n1060), .A2(n1061), .ZN(G66) );
NOR3_X1 U766 ( .A1(n1016), .A2(n1062), .A3(n1063), .ZN(n1061) );
NOR3_X1 U767 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NOR2_X1 U768 ( .A1(n1067), .A2(n1068), .ZN(n1062) );
NOR2_X1 U769 ( .A1(n1069), .A2(n1065), .ZN(n1067) );
XOR2_X1 U770 ( .A(G217), .B(KEYINPUT60), .Z(n1065) );
NOR2_X1 U771 ( .A1(n1060), .A2(n1070), .ZN(G63) );
NOR3_X1 U772 ( .A1(n1011), .A2(n1071), .A3(n1072), .ZN(n1070) );
NOR3_X1 U773 ( .A1(n1073), .A2(n1074), .A3(n1066), .ZN(n1072) );
INV_X1 U774 ( .A(n1075), .ZN(n1073) );
NOR2_X1 U775 ( .A1(n1076), .A2(n1075), .ZN(n1071) );
NOR2_X1 U776 ( .A1(n1069), .A2(n1074), .ZN(n1076) );
INV_X1 U777 ( .A(n974), .ZN(n1069) );
NOR3_X1 U778 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(G60) );
AND2_X1 U779 ( .A1(KEYINPUT56), .A2(n1060), .ZN(n1079) );
NOR3_X1 U780 ( .A1(KEYINPUT56), .A2(n1022), .A3(n1080), .ZN(n1078) );
INV_X1 U781 ( .A(G952), .ZN(n1080) );
XNOR2_X1 U782 ( .A(n1081), .B(n1082), .ZN(n1077) );
NOR2_X1 U783 ( .A1(n1083), .A2(n1066), .ZN(n1082) );
XNOR2_X1 U784 ( .A(G104), .B(n1084), .ZN(G6) );
NOR2_X1 U785 ( .A1(n1060), .A2(n1085), .ZN(G57) );
XOR2_X1 U786 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U787 ( .A1(n1088), .A2(n1066), .ZN(n1086) );
NOR2_X1 U788 ( .A1(n1060), .A2(n1089), .ZN(G54) );
XOR2_X1 U789 ( .A(n1090), .B(n1091), .Z(n1089) );
XOR2_X1 U790 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U791 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U792 ( .A1(G140), .A2(KEYINPUT25), .ZN(n1095) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1066), .ZN(n1094) );
XOR2_X1 U794 ( .A(n1097), .B(n1098), .Z(n1090) );
XNOR2_X1 U795 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND3_X1 U796 ( .A1(KEYINPUT49), .A2(n1101), .A3(n1102), .ZN(n1099) );
XOR2_X1 U797 ( .A(n1103), .B(KEYINPUT62), .Z(n1102) );
OR2_X1 U798 ( .A1(n1104), .A2(n1037), .ZN(n1103) );
NAND2_X1 U799 ( .A1(n1104), .A2(n1037), .ZN(n1101) );
XOR2_X1 U800 ( .A(n1105), .B(KEYINPUT34), .Z(n1104) );
XNOR2_X1 U801 ( .A(G110), .B(KEYINPUT18), .ZN(n1097) );
NOR2_X1 U802 ( .A1(n1060), .A2(n1106), .ZN(G51) );
XOR2_X1 U803 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U804 ( .A(KEYINPUT54), .B(n1109), .Z(n1108) );
NOR2_X1 U805 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U806 ( .A(n1112), .B(KEYINPUT41), .Z(n1111) );
NAND2_X1 U807 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
NOR2_X1 U808 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
XOR2_X1 U809 ( .A(n1115), .B(n1116), .Z(n1113) );
XNOR2_X1 U810 ( .A(KEYINPUT32), .B(n1117), .ZN(n1116) );
XNOR2_X1 U811 ( .A(n1118), .B(n1119), .ZN(n1115) );
NOR2_X1 U812 ( .A1(n1120), .A2(n1066), .ZN(n1107) );
NAND2_X1 U813 ( .A1(G902), .A2(n974), .ZN(n1066) );
NAND4_X1 U814 ( .A1(n1050), .A2(n1026), .A3(n1121), .A4(n1027), .ZN(n974) );
XNOR2_X1 U815 ( .A(KEYINPUT51), .B(n1025), .ZN(n1121) );
NAND3_X1 U816 ( .A1(n999), .A2(n1122), .A3(n1123), .ZN(n1025) );
XNOR2_X1 U817 ( .A(KEYINPUT59), .B(n1124), .ZN(n1122) );
AND4_X1 U818 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1026) );
NOR3_X1 U819 ( .A1(n1129), .A2(n1130), .A3(n1131), .ZN(n1128) );
INV_X1 U820 ( .A(n1132), .ZN(n1130) );
AND4_X1 U821 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1050) );
NOR4_X1 U822 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1136) );
NOR3_X1 U823 ( .A1(n1141), .A2(n985), .A3(n1142), .ZN(n1140) );
XNOR2_X1 U824 ( .A(KEYINPUT13), .B(n1124), .ZN(n1141) );
INV_X1 U825 ( .A(n1084), .ZN(n1139) );
NAND4_X1 U826 ( .A1(n992), .A2(n966), .A3(n967), .A4(n969), .ZN(n1084) );
NOR3_X1 U827 ( .A1(n999), .A2(KEYINPUT57), .A3(n1143), .ZN(n1138) );
NOR2_X1 U828 ( .A1(n1144), .A2(n1145), .ZN(n1137) );
NOR3_X1 U829 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1144) );
NOR2_X1 U830 ( .A1(n1143), .A2(n1149), .ZN(n1148) );
INV_X1 U831 ( .A(KEYINPUT57), .ZN(n1149) );
AND4_X1 U832 ( .A1(n969), .A2(n1150), .A3(n966), .A4(n965), .ZN(n1147) );
XNOR2_X1 U833 ( .A(KEYINPUT30), .B(n1151), .ZN(n1146) );
NOR2_X1 U834 ( .A1(n1022), .A2(G952), .ZN(n1060) );
XOR2_X1 U835 ( .A(G146), .B(n1152), .Z(G48) );
NOR3_X1 U836 ( .A1(n1153), .A2(n1145), .A3(n1124), .ZN(n1152) );
XNOR2_X1 U837 ( .A(G143), .B(n1127), .ZN(G45) );
NAND4_X1 U838 ( .A1(n1154), .A2(n999), .A3(n1155), .A4(n1156), .ZN(n1127) );
XOR2_X1 U839 ( .A(G140), .B(n1129), .Z(G42) );
AND3_X1 U840 ( .A1(n1004), .A2(n1014), .A3(n1123), .ZN(n1129) );
XNOR2_X1 U841 ( .A(G137), .B(n1157), .ZN(G39) );
NAND2_X1 U842 ( .A1(KEYINPUT40), .A2(n1158), .ZN(n1157) );
INV_X1 U843 ( .A(n1027), .ZN(n1158) );
NAND4_X1 U844 ( .A1(n987), .A2(n1159), .A3(n1014), .A4(n1160), .ZN(n1027) );
XOR2_X1 U845 ( .A(n1161), .B(G134), .Z(G36) );
NAND2_X1 U846 ( .A1(KEYINPUT45), .A2(n1125), .ZN(n1161) );
NAND3_X1 U847 ( .A1(n1014), .A2(n965), .A3(n1154), .ZN(n1125) );
AND3_X1 U848 ( .A1(n987), .A2(n1160), .A3(n1005), .ZN(n1154) );
XOR2_X1 U849 ( .A(G131), .B(n1131), .Z(G33) );
AND3_X1 U850 ( .A1(n1005), .A2(n1014), .A3(n1123), .ZN(n1131) );
INV_X1 U851 ( .A(n1153), .ZN(n1123) );
NAND3_X1 U852 ( .A1(n987), .A2(n1160), .A3(n992), .ZN(n1153) );
XNOR2_X1 U853 ( .A(n1150), .B(KEYINPUT46), .ZN(n987) );
NOR2_X1 U854 ( .A1(n1002), .A2(n1162), .ZN(n1014) );
INV_X1 U855 ( .A(n1000), .ZN(n1162) );
XNOR2_X1 U856 ( .A(G128), .B(n1132), .ZN(G30) );
NAND4_X1 U857 ( .A1(n1163), .A2(n965), .A3(n967), .A4(n1160), .ZN(n1132) );
XNOR2_X1 U858 ( .A(n1135), .B(n1164), .ZN(G3) );
NOR2_X1 U859 ( .A1(KEYINPUT53), .A2(n1165), .ZN(n1164) );
NAND4_X1 U860 ( .A1(n1005), .A2(n1166), .A3(n967), .A4(n969), .ZN(n1135) );
NOR2_X1 U861 ( .A1(n1167), .A2(n1145), .ZN(n967) );
XNOR2_X1 U862 ( .A(G125), .B(n1126), .ZN(G27) );
NAND3_X1 U863 ( .A1(n1004), .A2(n992), .A3(n1168), .ZN(n1126) );
AND3_X1 U864 ( .A1(n994), .A2(n1160), .A3(n999), .ZN(n1168) );
NAND2_X1 U865 ( .A1(n976), .A2(n1169), .ZN(n1160) );
NAND4_X1 U866 ( .A1(G953), .A2(G902), .A3(n1170), .A4(n1031), .ZN(n1169) );
INV_X1 U867 ( .A(G900), .ZN(n1031) );
NAND2_X1 U868 ( .A1(n1171), .A2(n1172), .ZN(G24) );
NAND2_X1 U869 ( .A1(G122), .A2(n1133), .ZN(n1172) );
XOR2_X1 U870 ( .A(n1173), .B(KEYINPUT3), .Z(n1171) );
OR2_X1 U871 ( .A1(n1133), .A2(G122), .ZN(n1173) );
NAND4_X1 U872 ( .A1(n1174), .A2(n966), .A3(n1155), .A4(n1156), .ZN(n1133) );
INV_X1 U873 ( .A(n981), .ZN(n966) );
NAND2_X1 U874 ( .A1(n1175), .A2(n1176), .ZN(n981) );
XOR2_X1 U875 ( .A(n1177), .B(n1178), .Z(G21) );
NAND2_X1 U876 ( .A1(n1174), .A2(n1159), .ZN(n1178) );
NOR2_X1 U877 ( .A1(n985), .A2(n1124), .ZN(n1159) );
INV_X1 U878 ( .A(n1163), .ZN(n1124) );
NOR2_X1 U879 ( .A1(n1176), .A2(n1175), .ZN(n1163) );
INV_X1 U880 ( .A(n1166), .ZN(n985) );
NAND2_X1 U881 ( .A1(KEYINPUT44), .A2(G119), .ZN(n1177) );
XOR2_X1 U882 ( .A(G116), .B(n1179), .Z(G18) );
NOR2_X1 U883 ( .A1(n1180), .A2(n1151), .ZN(n1179) );
NAND4_X1 U884 ( .A1(n1005), .A2(n994), .A3(n965), .A4(n969), .ZN(n1151) );
NOR2_X1 U885 ( .A1(n1156), .A2(n1181), .ZN(n965) );
XNOR2_X1 U886 ( .A(n999), .B(KEYINPUT23), .ZN(n1180) );
XNOR2_X1 U887 ( .A(G113), .B(n1134), .ZN(G15) );
NAND3_X1 U888 ( .A1(n992), .A2(n1174), .A3(n1005), .ZN(n1134) );
NOR2_X1 U889 ( .A1(n1175), .A2(n1182), .ZN(n1005) );
INV_X1 U890 ( .A(n1142), .ZN(n1174) );
NAND3_X1 U891 ( .A1(n999), .A2(n969), .A3(n994), .ZN(n1142) );
NOR2_X1 U892 ( .A1(n989), .A2(n1183), .ZN(n994) );
INV_X1 U893 ( .A(n988), .ZN(n1183) );
AND2_X1 U894 ( .A1(n1181), .A2(n1156), .ZN(n992) );
INV_X1 U895 ( .A(n1155), .ZN(n1181) );
XOR2_X1 U896 ( .A(n1184), .B(n1185), .Z(G12) );
NOR2_X1 U897 ( .A1(G110), .A2(KEYINPUT43), .ZN(n1185) );
NAND2_X1 U898 ( .A1(n1186), .A2(n999), .ZN(n1184) );
INV_X1 U899 ( .A(n1145), .ZN(n999) );
NAND2_X1 U900 ( .A1(n1002), .A2(n1000), .ZN(n1145) );
NAND2_X1 U901 ( .A1(G214), .A2(n1187), .ZN(n1000) );
XOR2_X1 U902 ( .A(n1188), .B(n1120), .Z(n1002) );
NAND2_X1 U903 ( .A1(G210), .A2(n1187), .ZN(n1120) );
NAND2_X1 U904 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
NAND2_X1 U905 ( .A1(n1191), .A2(n1190), .ZN(n1188) );
XOR2_X1 U906 ( .A(n1192), .B(n1193), .Z(n1191) );
XOR2_X1 U907 ( .A(n1194), .B(n1195), .Z(n1193) );
NAND2_X1 U908 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U909 ( .A1(n1198), .A2(n1117), .ZN(n1197) );
XOR2_X1 U910 ( .A(n1118), .B(KEYINPUT35), .Z(n1198) );
NAND2_X1 U911 ( .A1(G125), .A2(n1199), .ZN(n1196) );
XOR2_X1 U912 ( .A(n1118), .B(KEYINPUT27), .Z(n1199) );
NAND2_X1 U913 ( .A1(KEYINPUT63), .A2(n1119), .ZN(n1194) );
NAND2_X1 U914 ( .A1(G224), .A2(n1022), .ZN(n1119) );
XOR2_X1 U915 ( .A(n1114), .B(KEYINPUT55), .Z(n1192) );
NAND2_X1 U916 ( .A1(n1055), .A2(n1200), .ZN(n1114) );
NAND2_X1 U917 ( .A1(n1058), .A2(n1057), .ZN(n1200) );
OR2_X1 U918 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
XNOR2_X1 U919 ( .A(G122), .B(n1201), .ZN(n1058) );
XNOR2_X1 U920 ( .A(n1202), .B(n1203), .ZN(n1057) );
XOR2_X1 U921 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U922 ( .A(n1206), .B(G113), .Z(n1202) );
NAND2_X1 U923 ( .A1(KEYINPUT9), .A2(n1207), .ZN(n1206) );
XOR2_X1 U924 ( .A(n1143), .B(KEYINPUT26), .Z(n1186) );
NAND4_X1 U925 ( .A1(n1004), .A2(n1166), .A3(n1150), .A4(n969), .ZN(n1143) );
NAND2_X1 U926 ( .A1(n976), .A2(n1208), .ZN(n969) );
NAND4_X1 U927 ( .A1(G953), .A2(G902), .A3(n1209), .A4(n1170), .ZN(n1208) );
XOR2_X1 U928 ( .A(KEYINPUT4), .B(G898), .Z(n1209) );
NAND3_X1 U929 ( .A1(n1170), .A2(n1022), .A3(G952), .ZN(n976) );
NAND2_X1 U930 ( .A1(G234), .A2(G237), .ZN(n1170) );
INV_X1 U931 ( .A(n1167), .ZN(n1150) );
NAND2_X1 U932 ( .A1(n1210), .A2(n989), .ZN(n1167) );
XOR2_X1 U933 ( .A(n1211), .B(n1096), .Z(n989) );
INV_X1 U934 ( .A(G469), .ZN(n1096) );
NAND2_X1 U935 ( .A1(n1212), .A2(n1190), .ZN(n1211) );
XOR2_X1 U936 ( .A(n1092), .B(n1213), .Z(n1212) );
XOR2_X1 U937 ( .A(n1214), .B(n1215), .Z(n1213) );
NAND3_X1 U938 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
NAND2_X1 U939 ( .A1(n1219), .A2(n1100), .ZN(n1218) );
NAND2_X1 U940 ( .A1(KEYINPUT52), .A2(n1220), .ZN(n1217) );
NAND2_X1 U941 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XNOR2_X1 U942 ( .A(KEYINPUT12), .B(n1100), .ZN(n1221) );
NAND2_X1 U943 ( .A1(n1223), .A2(n1224), .ZN(n1216) );
INV_X1 U944 ( .A(KEYINPUT52), .ZN(n1224) );
NAND2_X1 U945 ( .A1(n1225), .A2(n1226), .ZN(n1223) );
NAND2_X1 U946 ( .A1(KEYINPUT12), .A2(n1100), .ZN(n1226) );
OR3_X1 U947 ( .A1(n1219), .A2(KEYINPUT12), .A3(n1100), .ZN(n1225) );
NAND2_X1 U948 ( .A1(G227), .A2(n1022), .ZN(n1100) );
INV_X1 U949 ( .A(n1222), .ZN(n1219) );
NAND3_X1 U950 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(n1222) );
NAND2_X1 U951 ( .A1(G110), .A2(n1230), .ZN(n1229) );
OR3_X1 U952 ( .A1(n1230), .A2(n1231), .A3(G140), .ZN(n1228) );
INV_X1 U953 ( .A(KEYINPUT28), .ZN(n1230) );
NAND2_X1 U954 ( .A1(G140), .A2(n1231), .ZN(n1227) );
NAND2_X1 U955 ( .A1(KEYINPUT61), .A2(n1201), .ZN(n1231) );
NAND2_X1 U956 ( .A1(KEYINPUT48), .A2(n1232), .ZN(n1214) );
XOR2_X1 U957 ( .A(n1037), .B(n1105), .Z(n1232) );
XOR2_X1 U958 ( .A(G104), .B(n1205), .Z(n1105) );
XNOR2_X1 U959 ( .A(n1165), .B(G107), .ZN(n1205) );
XNOR2_X1 U960 ( .A(n1233), .B(G128), .ZN(n1037) );
NAND2_X1 U961 ( .A1(KEYINPUT8), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U962 ( .A(n1235), .B(n1236), .ZN(n1092) );
XOR2_X1 U963 ( .A(n988), .B(KEYINPUT2), .Z(n1210) );
NAND2_X1 U964 ( .A1(G221), .A2(n1237), .ZN(n988) );
NOR2_X1 U965 ( .A1(n1155), .A2(n1156), .ZN(n1166) );
XOR2_X1 U966 ( .A(n1010), .B(KEYINPUT22), .Z(n1156) );
XOR2_X1 U967 ( .A(n1238), .B(n1083), .Z(n1010) );
INV_X1 U968 ( .A(G475), .ZN(n1083) );
NAND2_X1 U969 ( .A1(n1081), .A2(n1190), .ZN(n1238) );
XNOR2_X1 U970 ( .A(n1239), .B(n1240), .ZN(n1081) );
XOR2_X1 U971 ( .A(n1241), .B(n1242), .Z(n1240) );
XNOR2_X1 U972 ( .A(n1207), .B(n1243), .ZN(n1242) );
NOR2_X1 U973 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
INV_X1 U974 ( .A(G214), .ZN(n1245) );
INV_X1 U975 ( .A(G104), .ZN(n1207) );
XOR2_X1 U976 ( .A(KEYINPUT38), .B(G122), .Z(n1241) );
XOR2_X1 U977 ( .A(n1246), .B(n1247), .Z(n1239) );
XNOR2_X1 U978 ( .A(n1234), .B(n1248), .ZN(n1246) );
XOR2_X1 U979 ( .A(n1011), .B(n1013), .Z(n1155) );
XNOR2_X1 U980 ( .A(n1074), .B(KEYINPUT14), .ZN(n1013) );
INV_X1 U981 ( .A(G478), .ZN(n1074) );
NOR2_X1 U982 ( .A1(n1075), .A2(G902), .ZN(n1011) );
XNOR2_X1 U983 ( .A(n1249), .B(n1250), .ZN(n1075) );
XOR2_X1 U984 ( .A(G107), .B(n1251), .Z(n1250) );
XOR2_X1 U985 ( .A(G122), .B(G116), .Z(n1251) );
XOR2_X1 U986 ( .A(n1252), .B(n1253), .Z(n1249) );
NOR2_X1 U987 ( .A1(KEYINPUT5), .A2(n1254), .ZN(n1253) );
XOR2_X1 U988 ( .A(n1255), .B(n1256), .Z(n1254) );
NOR2_X1 U989 ( .A1(KEYINPUT7), .A2(G128), .ZN(n1256) );
XNOR2_X1 U990 ( .A(G143), .B(G134), .ZN(n1255) );
NAND2_X1 U991 ( .A1(G217), .A2(n1257), .ZN(n1252) );
AND2_X1 U992 ( .A1(n1182), .A2(n1175), .ZN(n1004) );
NAND2_X1 U993 ( .A1(n1258), .A2(n1259), .ZN(n1175) );
NAND2_X1 U994 ( .A1(n1260), .A2(n1088), .ZN(n1259) );
INV_X1 U995 ( .A(G472), .ZN(n1088) );
XNOR2_X1 U996 ( .A(KEYINPUT20), .B(n1261), .ZN(n1260) );
NAND2_X1 U997 ( .A1(n1262), .A2(G472), .ZN(n1258) );
XNOR2_X1 U998 ( .A(n1015), .B(KEYINPUT50), .ZN(n1262) );
INV_X1 U999 ( .A(n1261), .ZN(n1015) );
NAND2_X1 U1000 ( .A1(n1263), .A2(n1190), .ZN(n1261) );
XOR2_X1 U1001 ( .A(KEYINPUT29), .B(n1087), .Z(n1263) );
XNOR2_X1 U1002 ( .A(n1264), .B(n1265), .ZN(n1087) );
XOR2_X1 U1003 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U1004 ( .A(n1268), .B(n1204), .Z(n1267) );
XOR2_X1 U1005 ( .A(G116), .B(G119), .Z(n1204) );
NOR2_X1 U1006 ( .A1(n1244), .A2(n1269), .ZN(n1268) );
INV_X1 U1007 ( .A(G210), .ZN(n1269) );
NAND2_X1 U1008 ( .A1(n1270), .A2(n1022), .ZN(n1244) );
XNOR2_X1 U1009 ( .A(KEYINPUT33), .B(n1189), .ZN(n1270) );
INV_X1 U1010 ( .A(G237), .ZN(n1189) );
XNOR2_X1 U1011 ( .A(KEYINPUT16), .B(n1165), .ZN(n1266) );
INV_X1 U1012 ( .A(G101), .ZN(n1165) );
XOR2_X1 U1013 ( .A(n1271), .B(n1247), .Z(n1264) );
XNOR2_X1 U1014 ( .A(G113), .B(n1235), .ZN(n1247) );
INV_X1 U1015 ( .A(n1036), .ZN(n1235) );
XOR2_X1 U1016 ( .A(G131), .B(KEYINPUT17), .Z(n1036) );
XOR2_X1 U1017 ( .A(n1118), .B(n1236), .Z(n1271) );
XOR2_X1 U1018 ( .A(G134), .B(n1272), .Z(n1236) );
NOR2_X1 U1019 ( .A1(KEYINPUT21), .A2(n1273), .ZN(n1272) );
INV_X1 U1020 ( .A(G137), .ZN(n1273) );
XNOR2_X1 U1021 ( .A(G128), .B(n1234), .ZN(n1118) );
XNOR2_X1 U1022 ( .A(G143), .B(n1274), .ZN(n1234) );
INV_X1 U1023 ( .A(n1275), .ZN(n1274) );
INV_X1 U1024 ( .A(n1176), .ZN(n1182) );
XOR2_X1 U1025 ( .A(n1016), .B(n1276), .Z(n1176) );
NOR2_X1 U1026 ( .A1(KEYINPUT58), .A2(n1277), .ZN(n1276) );
XNOR2_X1 U1027 ( .A(n1017), .B(KEYINPUT36), .ZN(n1277) );
AND2_X1 U1028 ( .A1(G217), .A2(n1237), .ZN(n1017) );
NAND2_X1 U1029 ( .A1(G234), .A2(n1190), .ZN(n1237) );
INV_X1 U1030 ( .A(G902), .ZN(n1190) );
NOR2_X1 U1031 ( .A1(n1068), .A2(G902), .ZN(n1016) );
INV_X1 U1032 ( .A(n1064), .ZN(n1068) );
XNOR2_X1 U1033 ( .A(n1278), .B(n1279), .ZN(n1064) );
XNOR2_X1 U1034 ( .A(n1201), .B(n1280), .ZN(n1279) );
XNOR2_X1 U1035 ( .A(n1281), .B(G119), .ZN(n1280) );
INV_X1 U1036 ( .A(G128), .ZN(n1281) );
INV_X1 U1037 ( .A(G110), .ZN(n1201) );
XNOR2_X1 U1038 ( .A(n1035), .B(n1282), .ZN(n1278) );
XNOR2_X1 U1039 ( .A(n1283), .B(n1275), .ZN(n1282) );
XOR2_X1 U1040 ( .A(G146), .B(KEYINPUT39), .Z(n1275) );
NAND2_X1 U1041 ( .A1(G221), .A2(n1257), .ZN(n1283) );
AND2_X1 U1042 ( .A1(G234), .A2(n1022), .ZN(n1257) );
INV_X1 U1043 ( .A(G953), .ZN(n1022) );
XOR2_X1 U1044 ( .A(G137), .B(n1248), .Z(n1035) );
XNOR2_X1 U1045 ( .A(n1117), .B(G140), .ZN(n1248) );
INV_X1 U1046 ( .A(G125), .ZN(n1117) );
endmodule


