//Key = 0010011111000001100000111001110010010010010100011000001101000010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361;

XNOR2_X1 U750 ( .A(n1036), .B(n1037), .ZN(G9) );
NOR3_X1 U751 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND4_X1 U752 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(G75) );
NAND4_X1 U753 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1043) );
NOR4_X1 U754 ( .A1(n1049), .A2(n1050), .A3(n1051), .A4(n1052), .ZN(n1048) );
XNOR2_X1 U755 ( .A(KEYINPUT17), .B(n1053), .ZN(n1052) );
XNOR2_X1 U756 ( .A(G472), .B(n1054), .ZN(n1051) );
XOR2_X1 U757 ( .A(n1055), .B(n1056), .Z(n1050) );
XNOR2_X1 U758 ( .A(KEYINPUT56), .B(n1057), .ZN(n1056) );
NOR2_X1 U759 ( .A1(KEYINPUT52), .A2(n1058), .ZN(n1055) );
INV_X1 U760 ( .A(n1059), .ZN(n1058) );
NOR3_X1 U761 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1047) );
AND2_X1 U762 ( .A1(n1063), .A2(G217), .ZN(n1060) );
XNOR2_X1 U763 ( .A(n1064), .B(n1065), .ZN(n1046) );
NOR2_X1 U764 ( .A1(n1066), .A2(KEYINPUT49), .ZN(n1065) );
XNOR2_X1 U765 ( .A(n1067), .B(n1068), .ZN(n1045) );
NAND2_X1 U766 ( .A1(KEYINPUT22), .A2(n1069), .ZN(n1068) );
NAND2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1042) );
NAND2_X1 U768 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND4_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
NAND2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U772 ( .A1(n1038), .A2(n1082), .ZN(n1081) );
NAND2_X1 U773 ( .A1(n1083), .A2(n1061), .ZN(n1082) );
NAND2_X1 U774 ( .A1(n1084), .A2(n1085), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1086), .A2(n1040), .ZN(n1085) );
NAND3_X1 U776 ( .A1(n1084), .A2(n1087), .A3(n1080), .ZN(n1072) );
NAND2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NAND2_X1 U778 ( .A1(n1074), .A2(n1090), .ZN(n1089) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U780 ( .A1(n1076), .A2(n1093), .ZN(n1092) );
NAND2_X1 U781 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U782 ( .A1(n1062), .A2(n1096), .ZN(n1095) );
NAND2_X1 U783 ( .A1(n1075), .A2(n1097), .ZN(n1091) );
NAND2_X1 U784 ( .A1(n1098), .A2(n1075), .ZN(n1088) );
INV_X1 U785 ( .A(n1099), .ZN(n1070) );
NAND2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(G72) );
NAND3_X1 U787 ( .A1(n1102), .A2(n1103), .A3(G953), .ZN(n1101) );
XOR2_X1 U788 ( .A(KEYINPUT9), .B(n1104), .Z(n1100) );
NOR2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U790 ( .A(n1107), .B(n1103), .ZN(n1106) );
NAND2_X1 U791 ( .A1(n1108), .A2(n1109), .ZN(n1103) );
NAND2_X1 U792 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1108) );
XNOR2_X1 U794 ( .A(n1113), .B(n1114), .ZN(n1112) );
XOR2_X1 U795 ( .A(n1115), .B(n1116), .Z(n1111) );
XNOR2_X1 U796 ( .A(n1117), .B(n1118), .ZN(n1115) );
NAND2_X1 U797 ( .A1(KEYINPUT57), .A2(n1119), .ZN(n1117) );
NAND2_X1 U798 ( .A1(KEYINPUT5), .A2(n1120), .ZN(n1107) );
AND2_X1 U799 ( .A1(n1102), .A2(G953), .ZN(n1105) );
NAND2_X1 U800 ( .A1(G900), .A2(G227), .ZN(n1102) );
XOR2_X1 U801 ( .A(n1121), .B(n1122), .Z(G69) );
XOR2_X1 U802 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U803 ( .A1(n1125), .A2(n1044), .ZN(n1124) );
AND2_X1 U804 ( .A1(G224), .A2(G898), .ZN(n1125) );
NAND2_X1 U805 ( .A1(n1126), .A2(n1127), .ZN(n1123) );
NAND2_X1 U806 ( .A1(G953), .A2(n1128), .ZN(n1127) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1126) );
NAND2_X1 U808 ( .A1(n1044), .A2(n1131), .ZN(n1121) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1134), .B(n1135), .ZN(n1133) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
INV_X1 U812 ( .A(G217), .ZN(n1136) );
NOR2_X1 U813 ( .A1(n1132), .A2(n1138), .ZN(G63) );
NOR3_X1 U814 ( .A1(n1067), .A2(n1139), .A3(n1140), .ZN(n1138) );
NOR4_X1 U815 ( .A1(n1141), .A2(n1142), .A3(n1069), .A4(n1137), .ZN(n1140) );
NOR2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1139) );
NOR3_X1 U817 ( .A1(n1142), .A2(n1041), .A3(n1069), .ZN(n1144) );
INV_X1 U818 ( .A(G478), .ZN(n1069) );
INV_X1 U819 ( .A(KEYINPUT7), .ZN(n1142) );
NOR2_X1 U820 ( .A1(n1132), .A2(n1145), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1059), .A2(n1146), .A3(n1147), .ZN(n1145) );
NOR3_X1 U822 ( .A1(n1148), .A2(n1057), .A3(n1137), .ZN(n1147) );
NOR2_X1 U823 ( .A1(n1149), .A2(n1150), .ZN(n1146) );
NOR2_X1 U824 ( .A1(n1041), .A2(n1057), .ZN(n1149) );
XOR2_X1 U825 ( .A(G104), .B(n1151), .Z(G6) );
NOR2_X1 U826 ( .A1(n1132), .A2(n1152), .ZN(G57) );
XOR2_X1 U827 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U829 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR3_X1 U830 ( .A1(n1137), .A2(KEYINPUT60), .A3(n1159), .ZN(n1155) );
INV_X1 U831 ( .A(G472), .ZN(n1159) );
NOR2_X1 U832 ( .A1(n1132), .A2(n1160), .ZN(G54) );
XOR2_X1 U833 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U834 ( .A(n1163), .B(n1164), .ZN(n1162) );
XOR2_X1 U835 ( .A(n1116), .B(n1165), .Z(n1161) );
XOR2_X1 U836 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U837 ( .A1(n1168), .A2(n1137), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1132), .A2(n1169), .ZN(G51) );
XOR2_X1 U839 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U841 ( .A1(n1064), .A2(n1137), .ZN(n1173) );
OR2_X1 U842 ( .A1(n1174), .A2(n1041), .ZN(n1137) );
NOR2_X1 U843 ( .A1(n1131), .A2(n1120), .ZN(n1041) );
NAND4_X1 U844 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1120) );
NOR4_X1 U845 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1178) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1184), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR4_X1 U848 ( .A1(n1187), .A2(n1074), .A3(n1040), .A4(n1188), .ZN(n1183) );
NAND4_X1 U849 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1131) );
NOR4_X1 U850 ( .A1(n1193), .A2(n1194), .A3(n1151), .A4(n1195), .ZN(n1192) );
INV_X1 U851 ( .A(n1196), .ZN(n1195) );
NOR3_X1 U852 ( .A1(n1038), .A2(n1039), .A3(n1086), .ZN(n1151) );
NOR2_X1 U853 ( .A1(n1197), .A2(n1198), .ZN(n1191) );
NOR3_X1 U854 ( .A1(n1199), .A2(n1039), .A3(n1040), .ZN(n1198) );
XNOR2_X1 U855 ( .A(KEYINPUT16), .B(n1038), .ZN(n1199) );
NOR3_X1 U856 ( .A1(n1086), .A2(n1200), .A3(n1201), .ZN(n1197) );
XNOR2_X1 U857 ( .A(n1084), .B(KEYINPUT33), .ZN(n1200) );
XOR2_X1 U858 ( .A(n1202), .B(n1203), .Z(n1170) );
NOR3_X1 U859 ( .A1(KEYINPUT63), .A2(n1204), .A3(n1205), .ZN(n1203) );
NOR2_X1 U860 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XOR2_X1 U861 ( .A(KEYINPUT28), .B(n1208), .Z(n1206) );
NOR2_X1 U862 ( .A1(n1113), .A2(n1209), .ZN(n1204) );
XNOR2_X1 U863 ( .A(n1208), .B(KEYINPUT43), .ZN(n1209) );
NOR2_X1 U864 ( .A1(n1044), .A2(G952), .ZN(n1132) );
NAND2_X1 U865 ( .A1(n1210), .A2(n1211), .ZN(G48) );
NAND2_X1 U866 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U867 ( .A(n1214), .B(KEYINPUT40), .Z(n1210) );
NAND2_X1 U868 ( .A1(G146), .A2(n1175), .ZN(n1214) );
INV_X1 U869 ( .A(n1212), .ZN(n1175) );
NOR4_X1 U870 ( .A1(n1188), .A2(n1086), .A3(n1074), .A4(n1187), .ZN(n1212) );
XOR2_X1 U871 ( .A(n1176), .B(n1215), .Z(G45) );
NOR2_X1 U872 ( .A1(G143), .A2(KEYINPUT21), .ZN(n1215) );
NAND4_X1 U873 ( .A1(n1216), .A2(n1098), .A3(n1217), .A4(n1218), .ZN(n1176) );
INV_X1 U874 ( .A(n1188), .ZN(n1216) );
NAND3_X1 U875 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1188) );
XOR2_X1 U876 ( .A(G140), .B(n1182), .Z(G42) );
NOR2_X1 U877 ( .A1(n1186), .A2(n1222), .ZN(n1182) );
INV_X1 U878 ( .A(n1223), .ZN(n1222) );
XOR2_X1 U879 ( .A(n1224), .B(n1225), .Z(G39) );
XOR2_X1 U880 ( .A(KEYINPUT54), .B(G137), .Z(n1225) );
NAND4_X1 U881 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1220), .ZN(n1224) );
XOR2_X1 U882 ( .A(KEYINPUT44), .B(n1075), .Z(n1228) );
XNOR2_X1 U883 ( .A(KEYINPUT25), .B(n1038), .ZN(n1227) );
XNOR2_X1 U884 ( .A(n1119), .B(n1181), .ZN(G36) );
NOR3_X1 U885 ( .A1(n1229), .A2(n1040), .A3(n1186), .ZN(n1181) );
INV_X1 U886 ( .A(G134), .ZN(n1119) );
XOR2_X1 U887 ( .A(n1180), .B(n1230), .Z(G33) );
NOR2_X1 U888 ( .A1(KEYINPUT46), .A2(n1231), .ZN(n1230) );
NOR3_X1 U889 ( .A1(n1086), .A2(n1229), .A3(n1186), .ZN(n1180) );
NAND3_X1 U890 ( .A1(n1075), .A2(n1220), .A3(n1221), .ZN(n1186) );
NAND2_X1 U891 ( .A1(n1232), .A2(n1233), .ZN(G30) );
NAND2_X1 U892 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U893 ( .A(KEYINPUT35), .B(n1236), .Z(n1232) );
NOR2_X1 U894 ( .A1(n1234), .A2(n1235), .ZN(n1236) );
AND4_X1 U895 ( .A1(n1221), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1234) );
NOR3_X1 U896 ( .A1(n1094), .A2(n1187), .A3(n1074), .ZN(n1239) );
INV_X1 U897 ( .A(n1219), .ZN(n1094) );
XOR2_X1 U898 ( .A(n1220), .B(KEYINPUT59), .Z(n1238) );
XNOR2_X1 U899 ( .A(G101), .B(n1240), .ZN(G3) );
NAND2_X1 U900 ( .A1(KEYINPUT29), .A2(n1194), .ZN(n1240) );
NOR3_X1 U901 ( .A1(n1201), .A2(n1038), .A3(n1241), .ZN(n1194) );
INV_X1 U902 ( .A(n1221), .ZN(n1038) );
XOR2_X1 U903 ( .A(G125), .B(n1179), .Z(G27) );
AND4_X1 U904 ( .A1(n1223), .A2(n1084), .A3(n1219), .A4(n1220), .ZN(n1179) );
NAND2_X1 U905 ( .A1(n1099), .A2(n1242), .ZN(n1220) );
NAND4_X1 U906 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1110), .ZN(n1242) );
INV_X1 U907 ( .A(G900), .ZN(n1110) );
NOR3_X1 U908 ( .A1(n1244), .A2(n1187), .A3(n1086), .ZN(n1223) );
XNOR2_X1 U909 ( .A(G122), .B(n1189), .ZN(G24) );
NAND4_X1 U910 ( .A1(n1084), .A2(n1245), .A3(n1217), .A4(n1218), .ZN(n1189) );
INV_X1 U911 ( .A(n1039), .ZN(n1245) );
NAND3_X1 U912 ( .A1(n1074), .A2(n1076), .A3(n1246), .ZN(n1039) );
XNOR2_X1 U913 ( .A(G119), .B(n1190), .ZN(G21) );
NAND3_X1 U914 ( .A1(n1084), .A2(n1246), .A3(n1226), .ZN(n1190) );
INV_X1 U915 ( .A(n1185), .ZN(n1226) );
NAND2_X1 U916 ( .A1(n1247), .A2(n1244), .ZN(n1185) );
INV_X1 U917 ( .A(n1248), .ZN(n1084) );
XNOR2_X1 U918 ( .A(n1249), .B(n1193), .ZN(G18) );
NOR3_X1 U919 ( .A1(n1248), .A2(n1040), .A3(n1201), .ZN(n1193) );
INV_X1 U920 ( .A(n1237), .ZN(n1040) );
NOR2_X1 U921 ( .A1(n1250), .A2(n1218), .ZN(n1237) );
XNOR2_X1 U922 ( .A(G113), .B(n1251), .ZN(G15) );
NOR2_X1 U923 ( .A1(KEYINPUT19), .A2(n1252), .ZN(n1251) );
NOR3_X1 U924 ( .A1(n1086), .A2(n1248), .A3(n1201), .ZN(n1252) );
NAND2_X1 U925 ( .A1(n1098), .A2(n1246), .ZN(n1201) );
INV_X1 U926 ( .A(n1229), .ZN(n1098) );
NAND2_X1 U927 ( .A1(n1076), .A2(n1244), .ZN(n1229) );
XNOR2_X1 U928 ( .A(n1097), .B(KEYINPUT30), .ZN(n1076) );
NAND2_X1 U929 ( .A1(n1253), .A2(n1083), .ZN(n1248) );
XNOR2_X1 U930 ( .A(n1061), .B(KEYINPUT20), .ZN(n1253) );
NAND2_X1 U931 ( .A1(n1218), .A2(n1250), .ZN(n1086) );
XNOR2_X1 U932 ( .A(G110), .B(n1196), .ZN(G12) );
NAND4_X1 U933 ( .A1(n1247), .A2(n1221), .A3(n1074), .A4(n1246), .ZN(n1196) );
AND2_X1 U934 ( .A1(n1219), .A2(n1254), .ZN(n1246) );
NAND2_X1 U935 ( .A1(n1255), .A2(n1099), .ZN(n1254) );
NAND3_X1 U936 ( .A1(n1243), .A2(n1044), .A3(G952), .ZN(n1099) );
NAND4_X1 U937 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1128), .ZN(n1255) );
INV_X1 U938 ( .A(G898), .ZN(n1128) );
NAND2_X1 U939 ( .A1(G237), .A2(n1256), .ZN(n1243) );
NAND2_X1 U940 ( .A1(n1257), .A2(n1258), .ZN(n1219) );
OR3_X1 U941 ( .A1(n1096), .A2(n1062), .A3(KEYINPUT51), .ZN(n1258) );
INV_X1 U942 ( .A(n1259), .ZN(n1096) );
NAND2_X1 U943 ( .A1(KEYINPUT51), .A2(n1075), .ZN(n1257) );
NOR2_X1 U944 ( .A1(n1259), .A2(n1062), .ZN(n1075) );
AND2_X1 U945 ( .A1(G214), .A2(n1260), .ZN(n1062) );
NAND2_X1 U946 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
OR2_X1 U947 ( .A1(n1064), .A2(n1066), .ZN(n1262) );
XOR2_X1 U948 ( .A(n1263), .B(KEYINPUT14), .Z(n1261) );
NAND2_X1 U949 ( .A1(n1066), .A2(n1064), .ZN(n1263) );
NAND2_X1 U950 ( .A1(G210), .A2(n1260), .ZN(n1064) );
NAND2_X1 U951 ( .A1(n1174), .A2(n1264), .ZN(n1260) );
INV_X1 U952 ( .A(G237), .ZN(n1264) );
AND3_X1 U953 ( .A1(n1265), .A2(n1174), .A3(n1266), .ZN(n1066) );
XOR2_X1 U954 ( .A(n1267), .B(KEYINPUT0), .Z(n1266) );
NAND2_X1 U955 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
INV_X1 U956 ( .A(n1270), .ZN(n1269) );
XOR2_X1 U957 ( .A(n1172), .B(KEYINPUT23), .Z(n1268) );
NAND2_X1 U958 ( .A1(n1172), .A2(n1270), .ZN(n1265) );
XOR2_X1 U959 ( .A(n1208), .B(n1271), .Z(n1270) );
XNOR2_X1 U960 ( .A(n1202), .B(n1113), .ZN(n1271) );
NAND2_X1 U961 ( .A1(G224), .A2(n1044), .ZN(n1202) );
XOR2_X1 U962 ( .A(G128), .B(n1272), .Z(n1208) );
XOR2_X1 U963 ( .A(n1130), .B(n1273), .Z(n1172) );
NOR2_X1 U964 ( .A1(KEYINPUT12), .A2(n1129), .ZN(n1273) );
NAND2_X1 U965 ( .A1(n1274), .A2(n1275), .ZN(n1129) );
NAND2_X1 U966 ( .A1(n1276), .A2(G119), .ZN(n1275) );
NAND2_X1 U967 ( .A1(n1277), .A2(n1278), .ZN(n1274) );
XNOR2_X1 U968 ( .A(n1276), .B(KEYINPUT37), .ZN(n1277) );
XOR2_X1 U969 ( .A(n1279), .B(n1280), .Z(n1130) );
XNOR2_X1 U970 ( .A(n1036), .B(n1281), .ZN(n1280) );
XNOR2_X1 U971 ( .A(KEYINPUT50), .B(n1282), .ZN(n1281) );
XOR2_X1 U972 ( .A(n1283), .B(n1284), .Z(n1279) );
XNOR2_X1 U973 ( .A(G104), .B(n1285), .ZN(n1284) );
NAND2_X1 U974 ( .A1(KEYINPUT8), .A2(n1286), .ZN(n1283) );
INV_X1 U975 ( .A(n1244), .ZN(n1074) );
XNOR2_X1 U976 ( .A(n1287), .B(n1288), .ZN(n1244) );
NOR2_X1 U977 ( .A1(KEYINPUT11), .A2(n1289), .ZN(n1288) );
INV_X1 U978 ( .A(n1054), .ZN(n1289) );
NAND2_X1 U979 ( .A1(n1290), .A2(n1174), .ZN(n1054) );
XOR2_X1 U980 ( .A(n1153), .B(n1291), .Z(n1290) );
XOR2_X1 U981 ( .A(KEYINPUT38), .B(n1292), .Z(n1291) );
NOR2_X1 U982 ( .A1(n1158), .A2(n1293), .ZN(n1292) );
XOR2_X1 U983 ( .A(KEYINPUT39), .B(n1157), .Z(n1293) );
AND2_X1 U984 ( .A1(n1294), .A2(n1285), .ZN(n1157) );
INV_X1 U985 ( .A(G101), .ZN(n1285) );
NAND2_X1 U986 ( .A1(G210), .A2(n1295), .ZN(n1294) );
AND3_X1 U987 ( .A1(n1295), .A2(G101), .A3(G210), .ZN(n1158) );
XOR2_X1 U988 ( .A(n1296), .B(n1297), .Z(n1153) );
XNOR2_X1 U989 ( .A(n1278), .B(n1276), .ZN(n1297) );
XNOR2_X1 U990 ( .A(G113), .B(n1249), .ZN(n1276) );
INV_X1 U991 ( .A(G116), .ZN(n1249) );
INV_X1 U992 ( .A(G119), .ZN(n1278) );
XOR2_X1 U993 ( .A(n1298), .B(n1272), .Z(n1296) );
XNOR2_X1 U994 ( .A(n1299), .B(n1300), .ZN(n1272) );
NOR2_X1 U995 ( .A1(KEYINPUT42), .A2(G146), .ZN(n1300) );
XNOR2_X1 U996 ( .A(G143), .B(KEYINPUT34), .ZN(n1299) );
XNOR2_X1 U997 ( .A(G472), .B(KEYINPUT41), .ZN(n1287) );
NOR2_X1 U998 ( .A1(n1083), .A2(n1061), .ZN(n1221) );
AND2_X1 U999 ( .A1(G221), .A2(n1301), .ZN(n1061) );
OR2_X1 U1000 ( .A1(n1302), .A2(G902), .ZN(n1301) );
XNOR2_X1 U1001 ( .A(n1049), .B(KEYINPUT4), .ZN(n1083) );
XOR2_X1 U1002 ( .A(n1303), .B(n1168), .Z(n1049) );
INV_X1 U1003 ( .A(G469), .ZN(n1168) );
NAND2_X1 U1004 ( .A1(n1304), .A2(n1174), .ZN(n1303) );
XNOR2_X1 U1005 ( .A(n1305), .B(n1163), .ZN(n1304) );
XOR2_X1 U1006 ( .A(n1306), .B(n1307), .Z(n1163) );
XNOR2_X1 U1007 ( .A(n1118), .B(G101), .ZN(n1307) );
XOR2_X1 U1008 ( .A(n1298), .B(n1308), .Z(n1306) );
NOR3_X1 U1009 ( .A1(KEYINPUT58), .A2(n1309), .A3(n1310), .ZN(n1308) );
NOR2_X1 U1010 ( .A1(n1311), .A2(n1036), .ZN(n1310) );
INV_X1 U1011 ( .A(G107), .ZN(n1036) );
XOR2_X1 U1012 ( .A(KEYINPUT62), .B(G104), .Z(n1311) );
NOR2_X1 U1013 ( .A1(G107), .A2(n1312), .ZN(n1309) );
XOR2_X1 U1014 ( .A(KEYINPUT18), .B(G104), .Z(n1312) );
XNOR2_X1 U1015 ( .A(G134), .B(n1114), .ZN(n1298) );
XNOR2_X1 U1016 ( .A(n1313), .B(n1314), .ZN(n1114) );
XNOR2_X1 U1017 ( .A(G131), .B(G128), .ZN(n1313) );
XNOR2_X1 U1018 ( .A(G146), .B(n1315), .ZN(n1305) );
NOR2_X1 U1019 ( .A1(KEYINPUT61), .A2(n1316), .ZN(n1315) );
NOR2_X1 U1020 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
XOR2_X1 U1021 ( .A(n1319), .B(KEYINPUT27), .Z(n1318) );
NAND2_X1 U1022 ( .A1(n1320), .A2(n1166), .ZN(n1319) );
XOR2_X1 U1023 ( .A(n1321), .B(KEYINPUT31), .Z(n1320) );
NOR2_X1 U1024 ( .A1(n1166), .A2(n1321), .ZN(n1317) );
XNOR2_X1 U1025 ( .A(G140), .B(n1164), .ZN(n1321) );
XOR2_X1 U1026 ( .A(G110), .B(KEYINPUT10), .Z(n1164) );
AND2_X1 U1027 ( .A1(G227), .A2(n1044), .ZN(n1166) );
NOR2_X1 U1028 ( .A1(n1241), .A2(n1187), .ZN(n1247) );
INV_X1 U1029 ( .A(n1097), .ZN(n1187) );
NAND2_X1 U1030 ( .A1(n1053), .A2(n1322), .ZN(n1097) );
NAND2_X1 U1031 ( .A1(G217), .A2(n1063), .ZN(n1322) );
NAND2_X1 U1032 ( .A1(n1174), .A2(n1323), .ZN(n1063) );
NAND2_X1 U1033 ( .A1(n1302), .A2(n1324), .ZN(n1323) );
INV_X1 U1034 ( .A(n1134), .ZN(n1324) );
NAND3_X1 U1035 ( .A1(n1325), .A2(n1174), .A3(n1134), .ZN(n1053) );
XNOR2_X1 U1036 ( .A(n1326), .B(n1327), .ZN(n1134) );
XOR2_X1 U1037 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U1038 ( .A(n1330), .B(KEYINPUT3), .ZN(n1329) );
NAND2_X1 U1039 ( .A1(n1331), .A2(KEYINPUT2), .ZN(n1330) );
XOR2_X1 U1040 ( .A(n1332), .B(n1333), .Z(n1331) );
XNOR2_X1 U1041 ( .A(n1235), .B(G119), .ZN(n1333) );
INV_X1 U1042 ( .A(G128), .ZN(n1235) );
NAND2_X1 U1043 ( .A1(KEYINPUT48), .A2(n1282), .ZN(n1332) );
INV_X1 U1044 ( .A(G110), .ZN(n1282) );
AND3_X1 U1045 ( .A1(G221), .A2(n1044), .A3(G234), .ZN(n1328) );
XOR2_X1 U1046 ( .A(n1334), .B(n1314), .Z(n1326) );
XOR2_X1 U1047 ( .A(G137), .B(KEYINPUT32), .Z(n1314) );
XNOR2_X1 U1048 ( .A(n1116), .B(n1335), .ZN(n1334) );
XNOR2_X1 U1049 ( .A(G140), .B(n1213), .ZN(n1116) );
INV_X1 U1050 ( .A(G146), .ZN(n1213) );
INV_X1 U1051 ( .A(G902), .ZN(n1174) );
NAND2_X1 U1052 ( .A1(n1302), .A2(G217), .ZN(n1325) );
XNOR2_X1 U1053 ( .A(n1256), .B(KEYINPUT13), .ZN(n1302) );
XOR2_X1 U1054 ( .A(G234), .B(KEYINPUT36), .Z(n1256) );
INV_X1 U1055 ( .A(n1080), .ZN(n1241) );
NOR2_X1 U1056 ( .A1(n1218), .A2(n1217), .ZN(n1080) );
INV_X1 U1057 ( .A(n1250), .ZN(n1217) );
XNOR2_X1 U1058 ( .A(n1336), .B(n1337), .ZN(n1250) );
XOR2_X1 U1059 ( .A(KEYINPUT6), .B(KEYINPUT53), .Z(n1337) );
XNOR2_X1 U1060 ( .A(n1067), .B(G478), .ZN(n1336) );
NOR2_X1 U1061 ( .A1(n1143), .A2(G902), .ZN(n1067) );
INV_X1 U1062 ( .A(n1141), .ZN(n1143) );
NAND2_X1 U1063 ( .A1(n1338), .A2(n1339), .ZN(n1141) );
NAND2_X1 U1064 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
NAND3_X1 U1065 ( .A1(G234), .A2(n1044), .A3(G217), .ZN(n1341) );
XOR2_X1 U1066 ( .A(n1342), .B(KEYINPUT45), .Z(n1338) );
NAND4_X1 U1067 ( .A1(n1343), .A2(G217), .A3(G234), .A4(n1044), .ZN(n1342) );
INV_X1 U1068 ( .A(G953), .ZN(n1044) );
INV_X1 U1069 ( .A(n1340), .ZN(n1343) );
XNOR2_X1 U1070 ( .A(n1344), .B(n1345), .ZN(n1340) );
XNOR2_X1 U1071 ( .A(G107), .B(n1346), .ZN(n1345) );
NAND2_X1 U1072 ( .A1(n1347), .A2(KEYINPUT15), .ZN(n1346) );
XNOR2_X1 U1073 ( .A(G116), .B(n1348), .ZN(n1347) );
XNOR2_X1 U1074 ( .A(KEYINPUT24), .B(n1286), .ZN(n1348) );
INV_X1 U1075 ( .A(G122), .ZN(n1286) );
XNOR2_X1 U1076 ( .A(G128), .B(n1349), .ZN(n1344) );
XNOR2_X1 U1077 ( .A(n1118), .B(G134), .ZN(n1349) );
XNOR2_X1 U1078 ( .A(n1059), .B(n1057), .ZN(n1218) );
INV_X1 U1079 ( .A(G475), .ZN(n1057) );
NOR2_X1 U1080 ( .A1(n1150), .A2(G902), .ZN(n1059) );
INV_X1 U1081 ( .A(n1148), .ZN(n1150) );
XNOR2_X1 U1082 ( .A(n1350), .B(n1351), .ZN(n1148) );
XNOR2_X1 U1083 ( .A(n1352), .B(G104), .ZN(n1351) );
INV_X1 U1084 ( .A(G113), .ZN(n1352) );
XOR2_X1 U1085 ( .A(n1353), .B(n1354), .Z(n1350) );
NOR2_X1 U1086 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
XOR2_X1 U1087 ( .A(KEYINPUT47), .B(G214), .Z(n1356) );
INV_X1 U1088 ( .A(n1295), .ZN(n1355) );
NOR2_X1 U1089 ( .A1(G953), .A2(G237), .ZN(n1295) );
XOR2_X1 U1090 ( .A(n1357), .B(n1358), .Z(n1353) );
XNOR2_X1 U1091 ( .A(n1231), .B(n1359), .ZN(n1358) );
XNOR2_X1 U1092 ( .A(n1118), .B(G140), .ZN(n1359) );
INV_X1 U1093 ( .A(G143), .ZN(n1118) );
INV_X1 U1094 ( .A(G131), .ZN(n1231) );
XOR2_X1 U1095 ( .A(n1360), .B(n1335), .Z(n1357) );
XNOR2_X1 U1096 ( .A(n1207), .B(KEYINPUT26), .ZN(n1335) );
INV_X1 U1097 ( .A(n1113), .ZN(n1207) );
XOR2_X1 U1098 ( .A(G125), .B(KEYINPUT55), .Z(n1113) );
XNOR2_X1 U1099 ( .A(G122), .B(n1361), .ZN(n1360) );
NOR2_X1 U1100 ( .A1(G146), .A2(KEYINPUT1), .ZN(n1361) );
endmodule


