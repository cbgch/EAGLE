//Key = 0101001000100100000000111011010101000101111001010111010100111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421;

XOR2_X1 U782 ( .A(n1089), .B(n1090), .Z(G9) );
NAND4_X1 U783 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
NOR2_X1 U784 ( .A1(n1095), .A2(n1096), .ZN(G75) );
NOR4_X1 U785 ( .A1(G953), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1096) );
NOR2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NOR2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U788 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U791 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NOR2_X1 U792 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NOR2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1110) );
NOR2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NOR2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
NOR3_X1 U798 ( .A1(n1113), .A2(n1124), .A3(n1119), .ZN(n1106) );
NOR2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR4_X1 U800 ( .A1(n1127), .A2(n1109), .A3(n1119), .A4(n1113), .ZN(n1102) );
NOR2_X1 U801 ( .A1(n1128), .A2(n1094), .ZN(n1127) );
NOR3_X1 U802 ( .A1(n1097), .A2(G953), .A3(G952), .ZN(n1095) );
AND4_X1 U803 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1097) );
NOR4_X1 U804 ( .A1(n1133), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1132) );
XOR2_X1 U805 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U806 ( .A(KEYINPUT56), .B(KEYINPUT29), .Z(n1138) );
XOR2_X1 U807 ( .A(n1139), .B(G472), .Z(n1137) );
AND2_X1 U808 ( .A1(n1140), .A2(G475), .ZN(n1135) );
INV_X1 U809 ( .A(n1123), .ZN(n1134) );
NOR2_X1 U810 ( .A1(n1119), .A2(n1141), .ZN(n1131) );
XOR2_X1 U811 ( .A(n1142), .B(n1143), .Z(n1130) );
XOR2_X1 U812 ( .A(KEYINPUT59), .B(KEYINPUT27), .Z(n1143) );
XNOR2_X1 U813 ( .A(G478), .B(n1144), .ZN(n1142) );
XNOR2_X1 U814 ( .A(G469), .B(n1145), .ZN(n1129) );
NOR2_X1 U815 ( .A1(KEYINPUT19), .A2(n1146), .ZN(n1145) );
XOR2_X1 U816 ( .A(n1147), .B(n1148), .Z(G72) );
NOR3_X1 U817 ( .A1(n1149), .A2(KEYINPUT63), .A3(n1150), .ZN(n1148) );
NOR2_X1 U818 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND2_X1 U819 ( .A1(n1153), .A2(n1154), .ZN(n1147) );
OR2_X1 U820 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND3_X1 U821 ( .A1(n1157), .A2(n1155), .A3(n1156), .ZN(n1153) );
XNOR2_X1 U822 ( .A(n1158), .B(n1159), .ZN(n1156) );
XOR2_X1 U823 ( .A(n1160), .B(n1161), .Z(n1158) );
NAND4_X1 U824 ( .A1(KEYINPUT33), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1160) );
NAND2_X1 U825 ( .A1(KEYINPUT25), .A2(n1165), .ZN(n1164) );
NAND2_X1 U826 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U827 ( .A(KEYINPUT31), .B(n1168), .Z(n1167) );
NAND2_X1 U828 ( .A1(n1169), .A2(n1170), .ZN(n1163) );
INV_X1 U829 ( .A(KEYINPUT25), .ZN(n1170) );
NAND2_X1 U830 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
OR2_X1 U831 ( .A1(n1173), .A2(KEYINPUT31), .ZN(n1172) );
NAND3_X1 U832 ( .A1(n1173), .A2(n1166), .A3(KEYINPUT31), .ZN(n1171) );
NAND2_X1 U833 ( .A1(n1168), .A2(n1174), .ZN(n1162) );
NAND2_X1 U834 ( .A1(n1149), .A2(n1175), .ZN(n1155) );
NAND2_X1 U835 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U836 ( .A(n1178), .B(KEYINPUT39), .Z(n1176) );
NAND2_X1 U837 ( .A1(G953), .A2(n1152), .ZN(n1157) );
NAND3_X1 U838 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(G69) );
NAND3_X1 U839 ( .A1(KEYINPUT3), .A2(n1182), .A3(n1183), .ZN(n1181) );
XNOR2_X1 U840 ( .A(n1184), .B(n1185), .ZN(n1183) );
NAND2_X1 U841 ( .A1(G953), .A2(n1186), .ZN(n1182) );
NAND2_X1 U842 ( .A1(n1185), .A2(n1187), .ZN(n1186) );
NAND2_X1 U843 ( .A1(KEYINPUT1), .A2(n1188), .ZN(n1187) );
NAND4_X1 U844 ( .A1(G953), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1180) );
NAND2_X1 U845 ( .A1(KEYINPUT3), .A2(n1185), .ZN(n1190) );
OR2_X1 U846 ( .A1(n1185), .A2(KEYINPUT1), .ZN(n1189) );
AND2_X1 U847 ( .A1(n1191), .A2(n1192), .ZN(n1185) );
NAND2_X1 U848 ( .A1(G953), .A2(n1193), .ZN(n1192) );
XOR2_X1 U849 ( .A(n1194), .B(n1195), .Z(n1191) );
NOR2_X1 U850 ( .A1(KEYINPUT18), .A2(n1196), .ZN(n1195) );
XOR2_X1 U851 ( .A(G224), .B(KEYINPUT24), .Z(n1188) );
NAND3_X1 U852 ( .A1(G953), .A2(n1193), .A3(KEYINPUT1), .ZN(n1179) );
NOR2_X1 U853 ( .A1(n1197), .A2(n1198), .ZN(G66) );
XOR2_X1 U854 ( .A(n1199), .B(n1200), .Z(n1198) );
NAND2_X1 U855 ( .A1(n1201), .A2(n1202), .ZN(n1199) );
NOR2_X1 U856 ( .A1(n1197), .A2(n1203), .ZN(G63) );
NOR3_X1 U857 ( .A1(n1144), .A2(n1204), .A3(n1205), .ZN(n1203) );
AND3_X1 U858 ( .A1(n1206), .A2(G478), .A3(n1201), .ZN(n1205) );
NOR2_X1 U859 ( .A1(n1207), .A2(n1206), .ZN(n1204) );
AND2_X1 U860 ( .A1(n1099), .A2(G478), .ZN(n1207) );
NOR2_X1 U861 ( .A1(n1197), .A2(n1208), .ZN(G60) );
XOR2_X1 U862 ( .A(n1209), .B(n1210), .Z(n1208) );
NAND2_X1 U863 ( .A1(n1201), .A2(G475), .ZN(n1209) );
XOR2_X1 U864 ( .A(G104), .B(n1211), .Z(G6) );
NOR2_X1 U865 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U866 ( .A(n1214), .B(KEYINPUT7), .Z(n1212) );
NOR2_X1 U867 ( .A1(n1215), .A2(n1216), .ZN(G57) );
XOR2_X1 U868 ( .A(KEYINPUT11), .B(n1197), .Z(n1216) );
XOR2_X1 U869 ( .A(n1217), .B(n1218), .Z(n1215) );
XOR2_X1 U870 ( .A(n1219), .B(n1220), .Z(n1218) );
XOR2_X1 U871 ( .A(n1221), .B(n1222), .Z(n1217) );
XOR2_X1 U872 ( .A(n1223), .B(KEYINPUT51), .Z(n1222) );
NAND2_X1 U873 ( .A1(n1201), .A2(G472), .ZN(n1221) );
NOR2_X1 U874 ( .A1(n1197), .A2(n1224), .ZN(G54) );
XOR2_X1 U875 ( .A(n1225), .B(n1226), .Z(n1224) );
XOR2_X1 U876 ( .A(n1227), .B(n1228), .Z(n1226) );
XOR2_X1 U877 ( .A(n1223), .B(G140), .Z(n1228) );
NAND2_X1 U878 ( .A1(n1201), .A2(G469), .ZN(n1227) );
XNOR2_X1 U879 ( .A(n1229), .B(n1230), .ZN(n1225) );
NOR2_X1 U880 ( .A1(n1197), .A2(n1231), .ZN(G51) );
XOR2_X1 U881 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U882 ( .A(n1234), .B(KEYINPUT36), .Z(n1233) );
NAND2_X1 U883 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND2_X1 U884 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U885 ( .A(n1239), .B(KEYINPUT4), .Z(n1235) );
OR2_X1 U886 ( .A1(n1238), .A2(n1237), .ZN(n1239) );
XOR2_X1 U887 ( .A(n1240), .B(KEYINPUT17), .Z(n1237) );
NAND3_X1 U888 ( .A1(n1241), .A2(n1242), .A3(n1243), .ZN(n1238) );
NAND2_X1 U889 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NAND3_X1 U890 ( .A1(n1246), .A2(n1219), .A3(G125), .ZN(n1242) );
NAND2_X1 U891 ( .A1(n1247), .A2(n1248), .ZN(n1241) );
XOR2_X1 U892 ( .A(n1219), .B(n1246), .Z(n1247) );
NAND3_X1 U893 ( .A1(n1201), .A2(n1249), .A3(KEYINPUT49), .ZN(n1232) );
AND2_X1 U894 ( .A1(G902), .A2(n1099), .ZN(n1201) );
NAND3_X1 U895 ( .A1(n1177), .A2(n1250), .A3(n1184), .ZN(n1099) );
AND4_X1 U896 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1184) );
AND3_X1 U897 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(n1254) );
OR2_X1 U898 ( .A1(n1214), .A2(n1213), .ZN(n1253) );
NAND4_X1 U899 ( .A1(n1128), .A2(n1091), .A3(n1093), .A4(n1258), .ZN(n1214) );
NAND2_X1 U900 ( .A1(n1092), .A2(n1259), .ZN(n1251) );
NAND2_X1 U901 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
NAND3_X1 U902 ( .A1(n1125), .A2(n1093), .A3(n1262), .ZN(n1261) );
NAND2_X1 U903 ( .A1(n1091), .A2(n1263), .ZN(n1260) );
NAND2_X1 U904 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U905 ( .A1(n1266), .A2(n1094), .ZN(n1265) );
XNOR2_X1 U906 ( .A(n1093), .B(KEYINPUT55), .ZN(n1266) );
NAND2_X1 U907 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
XNOR2_X1 U908 ( .A(KEYINPUT62), .B(n1178), .ZN(n1250) );
NAND4_X1 U909 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1178) );
NAND4_X1 U910 ( .A1(n1126), .A2(n1094), .A3(n1273), .A4(n1274), .ZN(n1269) );
NAND2_X1 U911 ( .A1(KEYINPUT58), .A2(n1275), .ZN(n1274) );
NAND2_X1 U912 ( .A1(n1276), .A2(n1277), .ZN(n1273) );
INV_X1 U913 ( .A(KEYINPUT58), .ZN(n1277) );
NAND3_X1 U914 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1276) );
AND4_X1 U915 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1177) );
NOR2_X1 U916 ( .A1(n1149), .A2(G952), .ZN(n1197) );
XOR2_X1 U917 ( .A(n1281), .B(n1285), .Z(G48) );
XOR2_X1 U918 ( .A(n1286), .B(KEYINPUT14), .Z(n1285) );
NAND4_X1 U919 ( .A1(n1287), .A2(n1288), .A3(n1128), .A4(n1121), .ZN(n1281) );
XNOR2_X1 U920 ( .A(G143), .B(n1282), .ZN(G45) );
NAND4_X1 U921 ( .A1(n1287), .A2(n1121), .A3(n1268), .A4(n1126), .ZN(n1282) );
XOR2_X1 U922 ( .A(n1289), .B(n1283), .Z(G42) );
NAND3_X1 U923 ( .A1(n1128), .A2(n1125), .A3(n1290), .ZN(n1283) );
XNOR2_X1 U924 ( .A(G137), .B(n1284), .ZN(G39) );
NAND3_X1 U925 ( .A1(n1262), .A2(n1288), .A3(n1290), .ZN(n1284) );
XNOR2_X1 U926 ( .A(G134), .B(n1291), .ZN(G36) );
NAND2_X1 U927 ( .A1(n1292), .A2(n1094), .ZN(n1291) );
XNOR2_X1 U928 ( .A(G131), .B(n1270), .ZN(G33) );
NAND2_X1 U929 ( .A1(n1292), .A2(n1128), .ZN(n1270) );
AND2_X1 U930 ( .A1(n1290), .A2(n1126), .ZN(n1292) );
INV_X1 U931 ( .A(n1275), .ZN(n1290) );
NAND3_X1 U932 ( .A1(n1121), .A2(n1278), .A3(n1280), .ZN(n1275) );
INV_X1 U933 ( .A(n1119), .ZN(n1280) );
NAND2_X1 U934 ( .A1(n1293), .A2(n1117), .ZN(n1119) );
INV_X1 U935 ( .A(n1279), .ZN(n1121) );
XNOR2_X1 U936 ( .A(G128), .B(n1271), .ZN(G30) );
NAND4_X1 U937 ( .A1(n1287), .A2(n1288), .A3(n1093), .A4(n1094), .ZN(n1271) );
XNOR2_X1 U938 ( .A(G101), .B(n1252), .ZN(G3) );
NAND3_X1 U939 ( .A1(n1294), .A2(n1093), .A3(n1262), .ZN(n1252) );
XOR2_X1 U940 ( .A(n1248), .B(n1272), .Z(G27) );
NAND4_X1 U941 ( .A1(n1287), .A2(n1128), .A3(n1267), .A4(n1125), .ZN(n1272) );
AND2_X1 U942 ( .A1(n1115), .A2(n1278), .ZN(n1287) );
NAND2_X1 U943 ( .A1(n1295), .A2(n1296), .ZN(n1278) );
NAND4_X1 U944 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1152), .ZN(n1296) );
INV_X1 U945 ( .A(G900), .ZN(n1152) );
XNOR2_X1 U946 ( .A(KEYINPUT40), .B(n1101), .ZN(n1295) );
NAND2_X1 U947 ( .A1(n1298), .A2(n1299), .ZN(G24) );
NAND2_X1 U948 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
INV_X1 U949 ( .A(n1302), .ZN(n1301) );
XOR2_X1 U950 ( .A(n1303), .B(KEYINPUT20), .Z(n1300) );
XOR2_X1 U951 ( .A(n1304), .B(KEYINPUT43), .Z(n1298) );
NAND2_X1 U952 ( .A1(n1305), .A2(n1302), .ZN(n1304) );
NAND4_X1 U953 ( .A1(n1306), .A2(n1091), .A3(n1092), .A4(n1268), .ZN(n1302) );
XOR2_X1 U954 ( .A(n1113), .B(KEYINPUT6), .Z(n1306) );
XOR2_X1 U955 ( .A(KEYINPUT20), .B(G122), .Z(n1305) );
XNOR2_X1 U956 ( .A(n1255), .B(n1307), .ZN(G21) );
NOR2_X1 U957 ( .A1(KEYINPUT54), .A2(n1308), .ZN(n1307) );
NAND4_X1 U958 ( .A1(n1262), .A2(n1288), .A3(n1267), .A4(n1092), .ZN(n1255) );
AND2_X1 U959 ( .A1(n1309), .A2(n1141), .ZN(n1288) );
INV_X1 U960 ( .A(n1105), .ZN(n1262) );
XOR2_X1 U961 ( .A(n1310), .B(G116), .Z(G18) );
NAND2_X1 U962 ( .A1(KEYINPUT53), .A2(n1257), .ZN(n1310) );
NAND3_X1 U963 ( .A1(n1294), .A2(n1094), .A3(n1267), .ZN(n1257) );
NAND2_X1 U964 ( .A1(n1311), .A2(n1312), .ZN(n1094) );
NAND2_X1 U965 ( .A1(n1268), .A2(n1313), .ZN(n1312) );
NOR2_X1 U966 ( .A1(n1314), .A2(n1315), .ZN(n1268) );
NAND3_X1 U967 ( .A1(n1315), .A2(n1316), .A3(KEYINPUT13), .ZN(n1311) );
XOR2_X1 U968 ( .A(n1317), .B(n1256), .Z(G15) );
NAND3_X1 U969 ( .A1(n1267), .A2(n1294), .A3(n1128), .ZN(n1256) );
NOR2_X1 U970 ( .A1(n1316), .A2(n1315), .ZN(n1128) );
AND2_X1 U971 ( .A1(n1092), .A2(n1126), .ZN(n1294) );
NAND2_X1 U972 ( .A1(n1318), .A2(n1319), .ZN(n1126) );
OR3_X1 U973 ( .A1(n1141), .A2(n1320), .A3(KEYINPUT38), .ZN(n1319) );
NAND2_X1 U974 ( .A1(KEYINPUT38), .A2(n1091), .ZN(n1318) );
AND2_X1 U975 ( .A1(n1115), .A2(n1258), .ZN(n1092) );
INV_X1 U976 ( .A(n1213), .ZN(n1115) );
INV_X1 U977 ( .A(n1113), .ZN(n1267) );
NAND2_X1 U978 ( .A1(n1321), .A2(n1123), .ZN(n1113) );
XOR2_X1 U979 ( .A(n1322), .B(n1323), .Z(G12) );
NAND4_X1 U980 ( .A1(n1093), .A2(n1258), .A3(n1125), .A4(n1324), .ZN(n1323) );
NOR2_X1 U981 ( .A1(n1325), .A2(n1105), .ZN(n1324) );
NAND2_X1 U982 ( .A1(n1326), .A2(n1314), .ZN(n1105) );
INV_X1 U983 ( .A(n1316), .ZN(n1314) );
XNOR2_X1 U984 ( .A(G478), .B(n1327), .ZN(n1316) );
NOR2_X1 U985 ( .A1(n1144), .A2(KEYINPUT8), .ZN(n1327) );
NOR2_X1 U986 ( .A1(n1206), .A2(G902), .ZN(n1144) );
XOR2_X1 U987 ( .A(n1328), .B(n1329), .Z(n1206) );
XOR2_X1 U988 ( .A(n1330), .B(n1331), .Z(n1329) );
NOR2_X1 U989 ( .A1(G143), .A2(KEYINPUT32), .ZN(n1331) );
AND2_X1 U990 ( .A1(G217), .A2(n1332), .ZN(n1330) );
XOR2_X1 U991 ( .A(n1333), .B(n1334), .Z(n1328) );
NOR2_X1 U992 ( .A1(KEYINPUT2), .A2(n1335), .ZN(n1334) );
XOR2_X1 U993 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U994 ( .A(G107), .B(n1338), .Z(n1337) );
XOR2_X1 U995 ( .A(KEYINPUT22), .B(G116), .Z(n1336) );
XNOR2_X1 U996 ( .A(G134), .B(G128), .ZN(n1333) );
XOR2_X1 U997 ( .A(n1315), .B(n1313), .Z(n1326) );
INV_X1 U998 ( .A(KEYINPUT13), .ZN(n1313) );
NOR2_X1 U999 ( .A1(n1339), .A2(n1133), .ZN(n1315) );
NOR2_X1 U1000 ( .A1(n1140), .A2(G475), .ZN(n1133) );
AND2_X1 U1001 ( .A1(n1340), .A2(n1140), .ZN(n1339) );
NAND2_X1 U1002 ( .A1(n1210), .A2(n1341), .ZN(n1140) );
XOR2_X1 U1003 ( .A(n1342), .B(n1343), .Z(n1210) );
XOR2_X1 U1004 ( .A(G113), .B(n1344), .Z(n1343) );
NOR2_X1 U1005 ( .A1(KEYINPUT30), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1006 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1007 ( .A(n1348), .B(n1174), .Z(n1347) );
AND2_X1 U1008 ( .A1(n1349), .A2(G214), .ZN(n1348) );
XOR2_X1 U1009 ( .A(n1350), .B(n1351), .Z(n1346) );
XOR2_X1 U1010 ( .A(G146), .B(G143), .Z(n1351) );
NAND2_X1 U1011 ( .A1(n1352), .A2(n1353), .ZN(n1350) );
NAND2_X1 U1012 ( .A1(G125), .A2(n1289), .ZN(n1353) );
XOR2_X1 U1013 ( .A(KEYINPUT47), .B(n1354), .Z(n1352) );
NOR2_X1 U1014 ( .A1(G125), .A2(n1289), .ZN(n1354) );
INV_X1 U1015 ( .A(G140), .ZN(n1289) );
XNOR2_X1 U1016 ( .A(n1338), .B(n1355), .ZN(n1342) );
NOR2_X1 U1017 ( .A1(G104), .A2(KEYINPUT9), .ZN(n1355) );
XNOR2_X1 U1018 ( .A(G475), .B(KEYINPUT50), .ZN(n1340) );
XOR2_X1 U1019 ( .A(n1213), .B(KEYINPUT44), .Z(n1325) );
NAND2_X1 U1020 ( .A1(n1116), .A2(n1117), .ZN(n1213) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1356), .ZN(n1117) );
INV_X1 U1022 ( .A(n1293), .ZN(n1116) );
XOR2_X1 U1023 ( .A(n1357), .B(n1249), .Z(n1293) );
AND2_X1 U1024 ( .A1(G210), .A2(n1356), .ZN(n1249) );
NAND2_X1 U1025 ( .A1(n1358), .A2(n1341), .ZN(n1356) );
INV_X1 U1026 ( .A(G237), .ZN(n1358) );
NAND2_X1 U1027 ( .A1(n1359), .A2(n1341), .ZN(n1357) );
XOR2_X1 U1028 ( .A(n1360), .B(n1361), .Z(n1359) );
XOR2_X1 U1029 ( .A(KEYINPUT5), .B(n1246), .Z(n1361) );
INV_X1 U1030 ( .A(n1245), .ZN(n1246) );
NAND2_X1 U1031 ( .A1(G224), .A2(n1149), .ZN(n1245) );
XOR2_X1 U1032 ( .A(n1240), .B(n1362), .Z(n1360) );
NOR2_X1 U1033 ( .A1(n1244), .A2(n1363), .ZN(n1362) );
NOR2_X1 U1034 ( .A1(G125), .A2(n1364), .ZN(n1363) );
XOR2_X1 U1035 ( .A(KEYINPUT28), .B(n1365), .Z(n1364) );
INV_X1 U1036 ( .A(n1219), .ZN(n1365) );
NOR2_X1 U1037 ( .A1(n1248), .A2(n1219), .ZN(n1244) );
INV_X1 U1038 ( .A(G125), .ZN(n1248) );
XNOR2_X1 U1039 ( .A(n1194), .B(n1196), .ZN(n1240) );
NAND2_X1 U1040 ( .A1(n1366), .A2(n1367), .ZN(n1196) );
OR2_X1 U1041 ( .A1(n1368), .A2(n1322), .ZN(n1367) );
XOR2_X1 U1042 ( .A(n1369), .B(KEYINPUT21), .Z(n1366) );
NAND2_X1 U1043 ( .A1(n1368), .A2(n1322), .ZN(n1369) );
XOR2_X1 U1044 ( .A(n1338), .B(KEYINPUT37), .Z(n1368) );
XNOR2_X1 U1045 ( .A(n1303), .B(KEYINPUT23), .ZN(n1338) );
INV_X1 U1046 ( .A(G122), .ZN(n1303) );
XOR2_X1 U1047 ( .A(n1370), .B(n1371), .Z(n1194) );
NOR2_X1 U1048 ( .A1(KEYINPUT0), .A2(n1372), .ZN(n1371) );
NAND2_X1 U1049 ( .A1(n1373), .A2(n1374), .ZN(n1370) );
NAND2_X1 U1050 ( .A1(n1375), .A2(n1376), .ZN(n1374) );
INV_X1 U1051 ( .A(KEYINPUT35), .ZN(n1376) );
XOR2_X1 U1052 ( .A(G113), .B(n1377), .Z(n1375) );
NAND2_X1 U1053 ( .A1(n1378), .A2(KEYINPUT35), .ZN(n1373) );
XOR2_X1 U1054 ( .A(n1317), .B(n1379), .Z(n1378) );
NAND2_X1 U1055 ( .A1(G101), .A2(n1380), .ZN(n1379) );
INV_X1 U1056 ( .A(G113), .ZN(n1317) );
NAND2_X1 U1057 ( .A1(n1381), .A2(n1382), .ZN(n1125) );
OR2_X1 U1058 ( .A1(n1109), .A2(KEYINPUT42), .ZN(n1382) );
INV_X1 U1059 ( .A(n1091), .ZN(n1109) );
NOR2_X1 U1060 ( .A1(n1141), .A2(n1309), .ZN(n1091) );
NAND3_X1 U1061 ( .A1(n1320), .A2(n1141), .A3(KEYINPUT42), .ZN(n1381) );
XNOR2_X1 U1062 ( .A(n1383), .B(n1202), .ZN(n1141) );
AND2_X1 U1063 ( .A1(G217), .A2(n1384), .ZN(n1202) );
NAND2_X1 U1064 ( .A1(n1200), .A2(n1341), .ZN(n1383) );
XNOR2_X1 U1065 ( .A(n1385), .B(n1386), .ZN(n1200) );
XOR2_X1 U1066 ( .A(n1387), .B(n1388), .Z(n1386) );
XOR2_X1 U1067 ( .A(G128), .B(G119), .Z(n1388) );
XOR2_X1 U1068 ( .A(G146), .B(G137), .Z(n1387) );
XOR2_X1 U1069 ( .A(n1389), .B(n1159), .Z(n1385) );
XOR2_X1 U1070 ( .A(G140), .B(G125), .Z(n1159) );
XOR2_X1 U1071 ( .A(n1390), .B(G110), .Z(n1389) );
NAND2_X1 U1072 ( .A1(G221), .A2(n1332), .ZN(n1390) );
AND2_X1 U1073 ( .A1(G234), .A2(n1149), .ZN(n1332) );
INV_X1 U1074 ( .A(n1309), .ZN(n1320) );
XNOR2_X1 U1075 ( .A(n1391), .B(n1139), .ZN(n1309) );
NAND2_X1 U1076 ( .A1(n1392), .A2(n1341), .ZN(n1139) );
XNOR2_X1 U1077 ( .A(n1393), .B(n1220), .ZN(n1392) );
XOR2_X1 U1078 ( .A(n1394), .B(n1395), .Z(n1220) );
XOR2_X1 U1079 ( .A(G101), .B(n1396), .Z(n1395) );
XOR2_X1 U1080 ( .A(KEYINPUT34), .B(G113), .Z(n1396) );
XNOR2_X1 U1081 ( .A(n1397), .B(n1372), .ZN(n1394) );
XOR2_X1 U1082 ( .A(G116), .B(n1308), .Z(n1372) );
INV_X1 U1083 ( .A(G119), .ZN(n1308) );
NAND2_X1 U1084 ( .A1(G210), .A2(n1349), .ZN(n1397) );
NOR2_X1 U1085 ( .A1(G953), .A2(G237), .ZN(n1349) );
XOR2_X1 U1086 ( .A(n1398), .B(n1399), .Z(n1393) );
NAND2_X1 U1087 ( .A1(KEYINPUT26), .A2(n1219), .ZN(n1398) );
XOR2_X1 U1088 ( .A(n1400), .B(n1401), .Z(n1219) );
INV_X1 U1089 ( .A(n1402), .ZN(n1401) );
NAND2_X1 U1090 ( .A1(KEYINPUT10), .A2(n1286), .ZN(n1400) );
INV_X1 U1091 ( .A(G146), .ZN(n1286) );
NAND2_X1 U1092 ( .A1(KEYINPUT60), .A2(n1403), .ZN(n1391) );
INV_X1 U1093 ( .A(G472), .ZN(n1403) );
NAND2_X1 U1094 ( .A1(n1101), .A2(n1404), .ZN(n1258) );
NAND4_X1 U1095 ( .A1(G953), .A2(G902), .A3(n1297), .A4(n1193), .ZN(n1404) );
INV_X1 U1096 ( .A(G898), .ZN(n1193) );
NAND3_X1 U1097 ( .A1(n1297), .A2(n1149), .A3(G952), .ZN(n1101) );
INV_X1 U1098 ( .A(G953), .ZN(n1149) );
NAND2_X1 U1099 ( .A1(G237), .A2(G234), .ZN(n1297) );
XNOR2_X1 U1100 ( .A(n1279), .B(KEYINPUT12), .ZN(n1093) );
NAND2_X1 U1101 ( .A1(n1122), .A2(n1123), .ZN(n1279) );
NAND2_X1 U1102 ( .A1(G221), .A2(n1384), .ZN(n1123) );
NAND2_X1 U1103 ( .A1(G234), .A2(n1341), .ZN(n1384) );
INV_X1 U1104 ( .A(n1321), .ZN(n1122) );
XOR2_X1 U1105 ( .A(n1146), .B(G469), .Z(n1321) );
NAND2_X1 U1106 ( .A1(n1405), .A2(n1341), .ZN(n1146) );
INV_X1 U1107 ( .A(G902), .ZN(n1341) );
XNOR2_X1 U1108 ( .A(n1230), .B(n1406), .ZN(n1405) );
XOR2_X1 U1109 ( .A(n1407), .B(n1408), .Z(n1406) );
NOR2_X1 U1110 ( .A1(G140), .A2(KEYINPUT15), .ZN(n1408) );
NAND3_X1 U1111 ( .A1(n1409), .A2(n1410), .A3(n1411), .ZN(n1407) );
NAND2_X1 U1112 ( .A1(KEYINPUT57), .A2(n1399), .ZN(n1411) );
NAND3_X1 U1113 ( .A1(n1412), .A2(n1413), .A3(n1229), .ZN(n1410) );
INV_X1 U1114 ( .A(KEYINPUT57), .ZN(n1413) );
OR2_X1 U1115 ( .A1(n1229), .A2(n1412), .ZN(n1409) );
NOR2_X1 U1116 ( .A1(n1399), .A2(KEYINPUT48), .ZN(n1412) );
INV_X1 U1117 ( .A(n1223), .ZN(n1399) );
NAND3_X1 U1118 ( .A1(n1414), .A2(n1415), .A3(n1416), .ZN(n1223) );
NAND2_X1 U1119 ( .A1(KEYINPUT61), .A2(n1173), .ZN(n1416) );
OR3_X1 U1120 ( .A1(n1417), .A2(KEYINPUT61), .A3(n1174), .ZN(n1415) );
NAND2_X1 U1121 ( .A1(n1174), .A2(n1417), .ZN(n1414) );
NAND2_X1 U1122 ( .A1(KEYINPUT41), .A2(n1168), .ZN(n1417) );
INV_X1 U1123 ( .A(n1173), .ZN(n1168) );
XNOR2_X1 U1124 ( .A(G134), .B(G137), .ZN(n1173) );
INV_X1 U1125 ( .A(n1166), .ZN(n1174) );
XNOR2_X1 U1126 ( .A(G131), .B(KEYINPUT16), .ZN(n1166) );
XOR2_X1 U1127 ( .A(n1161), .B(n1377), .Z(n1229) );
XOR2_X1 U1128 ( .A(G101), .B(n1380), .Z(n1377) );
XNOR2_X1 U1129 ( .A(G104), .B(n1089), .ZN(n1380) );
INV_X1 U1130 ( .A(G107), .ZN(n1089) );
XNOR2_X1 U1131 ( .A(n1418), .B(n1419), .ZN(n1161) );
XOR2_X1 U1132 ( .A(KEYINPUT52), .B(KEYINPUT45), .Z(n1419) );
XOR2_X1 U1133 ( .A(n1402), .B(G146), .Z(n1418) );
XNOR2_X1 U1134 ( .A(G128), .B(n1420), .ZN(n1402) );
XOR2_X1 U1135 ( .A(KEYINPUT46), .B(G143), .Z(n1420) );
XNOR2_X1 U1136 ( .A(n1322), .B(n1421), .ZN(n1230) );
NOR2_X1 U1137 ( .A1(G953), .A2(n1151), .ZN(n1421) );
INV_X1 U1138 ( .A(G227), .ZN(n1151) );
INV_X1 U1139 ( .A(G110), .ZN(n1322) );
endmodule


