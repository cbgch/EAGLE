//Key = 1111011111101110010001101010110011001111100011010110110111010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350;

XNOR2_X1 U737 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR3_X1 U739 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
INV_X1 U740 ( .A(n1034), .ZN(n1033) );
NOR2_X1 U741 ( .A1(KEYINPUT28), .A2(n1035), .ZN(n1032) );
AND4_X1 U742 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1035) );
NAND3_X1 U743 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1031) );
NAND2_X1 U744 ( .A1(n1039), .A2(n1043), .ZN(n1042) );
NAND2_X1 U745 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U746 ( .A1(n1046), .A2(n1047), .A3(n1037), .ZN(n1045) );
NAND2_X1 U747 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U748 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
OR2_X1 U749 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U750 ( .A1(n1036), .A2(n1054), .ZN(n1048) );
NAND2_X1 U751 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U752 ( .A1(KEYINPUT28), .A2(n1057), .ZN(n1056) );
NAND2_X1 U753 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
NAND3_X1 U754 ( .A1(n1050), .A2(n1060), .A3(n1036), .ZN(n1044) );
NAND2_X1 U755 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U756 ( .A1(n1046), .A2(n1063), .ZN(n1062) );
NAND2_X1 U757 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U758 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U759 ( .A1(n1037), .A2(n1068), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U761 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
INV_X1 U762 ( .A(n1073), .ZN(n1069) );
INV_X1 U763 ( .A(n1074), .ZN(n1039) );
AND3_X1 U764 ( .A1(n1040), .A2(n1041), .A3(n1075), .ZN(n1029) );
NAND4_X1 U765 ( .A1(n1059), .A2(n1076), .A3(n1046), .A4(n1077), .ZN(n1040) );
NOR4_X1 U766 ( .A1(n1058), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1077) );
XNOR2_X1 U767 ( .A(n1081), .B(n1082), .ZN(n1080) );
NOR2_X1 U768 ( .A1(G475), .A2(KEYINPUT42), .ZN(n1082) );
XOR2_X1 U769 ( .A(n1083), .B(n1084), .Z(n1079) );
NAND2_X1 U770 ( .A1(KEYINPUT52), .A2(n1085), .ZN(n1083) );
XOR2_X1 U771 ( .A(n1086), .B(n1087), .Z(n1078) );
NAND2_X1 U772 ( .A1(KEYINPUT26), .A2(n1088), .ZN(n1086) );
XNOR2_X1 U773 ( .A(KEYINPUT59), .B(n1089), .ZN(n1088) );
INV_X1 U774 ( .A(n1067), .ZN(n1076) );
NAND2_X1 U775 ( .A1(n1090), .A2(n1091), .ZN(G72) );
NAND4_X1 U776 ( .A1(KEYINPUT9), .A2(n1092), .A3(n1093), .A4(n1041), .ZN(n1091) );
NAND2_X1 U777 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
NAND2_X1 U778 ( .A1(n1093), .A2(n1041), .ZN(n1095) );
XOR2_X1 U779 ( .A(n1096), .B(n1097), .Z(n1094) );
NOR2_X1 U780 ( .A1(n1098), .A2(n1041), .ZN(n1097) );
XOR2_X1 U781 ( .A(n1099), .B(KEYINPUT13), .Z(n1098) );
NAND2_X1 U782 ( .A1(G900), .A2(G227), .ZN(n1099) );
NAND2_X1 U783 ( .A1(KEYINPUT9), .A2(n1092), .ZN(n1096) );
NAND3_X1 U784 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1092) );
XOR2_X1 U785 ( .A(KEYINPUT24), .B(n1103), .Z(n1102) );
NOR2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U787 ( .A1(n1105), .A2(n1104), .ZN(n1101) );
NAND2_X1 U788 ( .A1(G953), .A2(n1106), .ZN(n1100) );
XOR2_X1 U789 ( .A(n1107), .B(n1108), .Z(G69) );
NAND2_X1 U790 ( .A1(G953), .A2(n1109), .ZN(n1108) );
NAND2_X1 U791 ( .A1(G898), .A2(G224), .ZN(n1109) );
NAND2_X1 U792 ( .A1(KEYINPUT0), .A2(n1110), .ZN(n1107) );
XOR2_X1 U793 ( .A(n1111), .B(n1112), .Z(n1110) );
AND2_X1 U794 ( .A1(n1113), .A2(n1041), .ZN(n1112) );
NOR3_X1 U795 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1111) );
NOR3_X1 U796 ( .A1(n1117), .A2(KEYINPUT47), .A3(n1041), .ZN(n1116) );
AND3_X1 U797 ( .A1(n1117), .A2(G953), .A3(KEYINPUT47), .ZN(n1115) );
XOR2_X1 U798 ( .A(n1118), .B(n1119), .Z(n1114) );
XOR2_X1 U799 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND2_X1 U800 ( .A1(KEYINPUT39), .A2(n1122), .ZN(n1120) );
XOR2_X1 U801 ( .A(KEYINPUT56), .B(n1123), .Z(n1118) );
NOR2_X1 U802 ( .A1(KEYINPUT35), .A2(n1124), .ZN(n1123) );
XNOR2_X1 U803 ( .A(n1125), .B(KEYINPUT29), .ZN(n1124) );
NOR3_X1 U804 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(G66) );
AND2_X1 U805 ( .A1(KEYINPUT32), .A2(n1129), .ZN(n1128) );
NOR3_X1 U806 ( .A1(KEYINPUT32), .A2(G953), .A3(G952), .ZN(n1127) );
XOR2_X1 U807 ( .A(n1130), .B(n1131), .Z(n1126) );
NOR2_X1 U808 ( .A1(n1089), .A2(n1132), .ZN(n1130) );
NOR2_X1 U809 ( .A1(n1129), .A2(n1133), .ZN(G63) );
XNOR2_X1 U810 ( .A(n1134), .B(n1135), .ZN(n1133) );
AND2_X1 U811 ( .A1(G478), .A2(n1136), .ZN(n1135) );
NOR3_X1 U812 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(G60) );
NOR3_X1 U813 ( .A1(n1140), .A2(n1041), .A3(n1075), .ZN(n1139) );
INV_X1 U814 ( .A(G952), .ZN(n1075) );
AND2_X1 U815 ( .A1(n1140), .A2(n1129), .ZN(n1138) );
INV_X1 U816 ( .A(KEYINPUT31), .ZN(n1140) );
NOR3_X1 U817 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(n1137) );
NOR3_X1 U818 ( .A1(n1144), .A2(n1081), .A3(n1145), .ZN(n1143) );
NOR2_X1 U819 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NOR2_X1 U820 ( .A1(n1034), .A2(n1148), .ZN(n1146) );
INV_X1 U821 ( .A(KEYINPUT16), .ZN(n1144) );
NOR3_X1 U822 ( .A1(KEYINPUT16), .A2(n1149), .A3(n1147), .ZN(n1142) );
AND2_X1 U823 ( .A1(n1147), .A2(n1149), .ZN(n1141) );
NOR2_X1 U824 ( .A1(n1132), .A2(n1148), .ZN(n1149) );
NAND2_X1 U825 ( .A1(n1150), .A2(n1151), .ZN(G6) );
NAND2_X1 U826 ( .A1(G104), .A2(n1152), .ZN(n1151) );
XOR2_X1 U827 ( .A(n1153), .B(KEYINPUT19), .Z(n1150) );
OR2_X1 U828 ( .A1(n1152), .A2(G104), .ZN(n1153) );
NOR2_X1 U829 ( .A1(n1129), .A2(n1154), .ZN(G57) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U831 ( .A1(n1085), .A2(n1132), .ZN(n1156) );
INV_X1 U832 ( .A(n1136), .ZN(n1132) );
INV_X1 U833 ( .A(G472), .ZN(n1085) );
NOR2_X1 U834 ( .A1(n1129), .A2(n1157), .ZN(G54) );
XOR2_X1 U835 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U836 ( .A(n1160), .B(n1161), .Z(n1159) );
AND2_X1 U837 ( .A1(G469), .A2(n1136), .ZN(n1161) );
NAND2_X1 U838 ( .A1(n1162), .A2(KEYINPUT6), .ZN(n1160) );
XOR2_X1 U839 ( .A(n1163), .B(KEYINPUT63), .Z(n1162) );
XOR2_X1 U840 ( .A(n1164), .B(n1165), .Z(n1158) );
XNOR2_X1 U841 ( .A(G140), .B(n1166), .ZN(n1165) );
INV_X1 U842 ( .A(G110), .ZN(n1166) );
NOR2_X1 U843 ( .A1(n1129), .A2(n1167), .ZN(G51) );
NOR2_X1 U844 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U845 ( .A(n1170), .B(KEYINPUT57), .Z(n1169) );
NAND2_X1 U846 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NOR2_X1 U847 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
XOR2_X1 U848 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U849 ( .A(n1175), .B(n1176), .ZN(n1174) );
NAND2_X1 U850 ( .A1(KEYINPUT10), .A2(n1177), .ZN(n1175) );
XOR2_X1 U851 ( .A(n1178), .B(n1179), .Z(n1173) );
NAND2_X1 U852 ( .A1(KEYINPUT14), .A2(n1180), .ZN(n1178) );
INV_X1 U853 ( .A(n1181), .ZN(n1180) );
AND2_X1 U854 ( .A1(n1136), .A2(G210), .ZN(n1171) );
NOR2_X1 U855 ( .A1(n1182), .A2(n1034), .ZN(n1136) );
NOR2_X1 U856 ( .A1(n1113), .A2(n1093), .ZN(n1034) );
NAND2_X1 U857 ( .A1(n1183), .A2(n1184), .ZN(n1093) );
AND4_X1 U858 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1188), .ZN(n1184) );
NOR4_X1 U859 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1183) );
NOR2_X1 U860 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
INV_X1 U861 ( .A(n1057), .ZN(n1193) );
NOR2_X1 U862 ( .A1(n1195), .A2(n1196), .ZN(n1191) );
NAND4_X1 U863 ( .A1(n1152), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1113) );
AND4_X1 U864 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1028), .ZN(n1199) );
NAND4_X1 U865 ( .A1(n1203), .A2(n1036), .A3(n1066), .A4(n1067), .ZN(n1028) );
NOR2_X1 U866 ( .A1(n1204), .A2(n1205), .ZN(n1198) );
NOR2_X1 U867 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1206) );
NOR2_X1 U869 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
INV_X1 U870 ( .A(KEYINPUT40), .ZN(n1211) );
AND2_X1 U871 ( .A1(n1212), .A2(KEYINPUT1), .ZN(n1208) );
NOR3_X1 U872 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1204) );
NOR2_X1 U873 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NOR2_X1 U874 ( .A1(KEYINPUT40), .A2(n1210), .ZN(n1217) );
NOR2_X1 U875 ( .A1(KEYINPUT1), .A2(n1195), .ZN(n1216) );
NAND3_X1 U876 ( .A1(n1203), .A2(n1036), .A3(n1218), .ZN(n1152) );
NOR2_X1 U877 ( .A1(n1041), .A2(G952), .ZN(n1129) );
NAND2_X1 U878 ( .A1(n1219), .A2(n1220), .ZN(G48) );
OR2_X1 U879 ( .A1(n1221), .A2(G146), .ZN(n1220) );
XOR2_X1 U880 ( .A(n1222), .B(KEYINPUT41), .Z(n1219) );
NAND2_X1 U881 ( .A1(G146), .A2(n1221), .ZN(n1222) );
NAND2_X1 U882 ( .A1(n1223), .A2(n1057), .ZN(n1221) );
XOR2_X1 U883 ( .A(n1194), .B(KEYINPUT55), .Z(n1223) );
NAND3_X1 U884 ( .A1(n1224), .A2(n1218), .A3(n1225), .ZN(n1194) );
XOR2_X1 U885 ( .A(G143), .B(n1190), .Z(G45) );
AND3_X1 U886 ( .A1(n1052), .A2(n1226), .A3(n1227), .ZN(n1190) );
XNOR2_X1 U887 ( .A(n1189), .B(n1228), .ZN(G42) );
NAND2_X1 U888 ( .A1(KEYINPUT17), .A2(G140), .ZN(n1228) );
NOR3_X1 U889 ( .A1(n1064), .A2(n1229), .A3(n1196), .ZN(n1189) );
INV_X1 U890 ( .A(n1218), .ZN(n1064) );
XNOR2_X1 U891 ( .A(G137), .B(n1230), .ZN(G39) );
NAND3_X1 U892 ( .A1(n1225), .A2(n1212), .A3(n1231), .ZN(n1230) );
XNOR2_X1 U893 ( .A(KEYINPUT2), .B(n1050), .ZN(n1231) );
INV_X1 U894 ( .A(n1195), .ZN(n1212) );
XOR2_X1 U895 ( .A(n1187), .B(n1232), .Z(G36) );
NAND2_X1 U896 ( .A1(KEYINPUT53), .A2(G134), .ZN(n1232) );
OR2_X1 U897 ( .A1(n1196), .A2(n1210), .ZN(n1187) );
XNOR2_X1 U898 ( .A(G131), .B(n1186), .ZN(G33) );
NAND3_X1 U899 ( .A1(n1052), .A2(n1218), .A3(n1233), .ZN(n1186) );
INV_X1 U900 ( .A(n1196), .ZN(n1233) );
NAND2_X1 U901 ( .A1(n1225), .A2(n1050), .ZN(n1196) );
NAND2_X1 U902 ( .A1(n1234), .A2(n1235), .ZN(n1050) );
OR3_X1 U903 ( .A1(n1236), .A2(n1058), .A3(KEYINPUT34), .ZN(n1235) );
NAND2_X1 U904 ( .A1(KEYINPUT34), .A2(n1057), .ZN(n1234) );
XOR2_X1 U905 ( .A(G128), .B(n1237), .Z(G30) );
NOR2_X1 U906 ( .A1(KEYINPUT62), .A2(n1188), .ZN(n1237) );
NAND3_X1 U907 ( .A1(n1066), .A2(n1224), .A3(n1227), .ZN(n1188) );
AND3_X1 U908 ( .A1(n1057), .A2(n1067), .A3(n1225), .ZN(n1227) );
AND2_X1 U909 ( .A1(n1073), .A2(n1238), .ZN(n1225) );
XOR2_X1 U910 ( .A(n1202), .B(n1239), .Z(G3) );
XNOR2_X1 U911 ( .A(G101), .B(KEYINPUT23), .ZN(n1239) );
NAND3_X1 U912 ( .A1(n1037), .A2(n1203), .A3(n1052), .ZN(n1202) );
XNOR2_X1 U913 ( .A(n1185), .B(n1240), .ZN(G27) );
NOR2_X1 U914 ( .A1(KEYINPUT54), .A2(n1177), .ZN(n1240) );
NAND4_X1 U915 ( .A1(n1218), .A2(n1038), .A3(n1053), .A4(n1238), .ZN(n1185) );
NAND2_X1 U916 ( .A1(n1074), .A2(n1241), .ZN(n1238) );
NAND4_X1 U917 ( .A1(G953), .A2(G902), .A3(n1242), .A4(n1106), .ZN(n1241) );
INV_X1 U918 ( .A(G900), .ZN(n1106) );
XNOR2_X1 U919 ( .A(G122), .B(n1197), .ZN(G24) );
NAND4_X1 U920 ( .A1(n1243), .A2(n1036), .A3(n1067), .A4(n1226), .ZN(n1197) );
NOR2_X1 U921 ( .A1(n1244), .A2(n1245), .ZN(n1036) );
XNOR2_X1 U922 ( .A(n1246), .B(n1247), .ZN(G21) );
NOR2_X1 U923 ( .A1(n1207), .A2(n1195), .ZN(n1247) );
NAND2_X1 U924 ( .A1(n1224), .A2(n1037), .ZN(n1195) );
AND2_X1 U925 ( .A1(n1245), .A2(n1244), .ZN(n1224) );
XOR2_X1 U926 ( .A(G116), .B(n1248), .Z(G18) );
NOR2_X1 U927 ( .A1(n1207), .A2(n1210), .ZN(n1248) );
NAND3_X1 U928 ( .A1(n1066), .A2(n1067), .A3(n1052), .ZN(n1210) );
XNOR2_X1 U929 ( .A(G113), .B(n1201), .ZN(G15) );
NAND3_X1 U930 ( .A1(n1243), .A2(n1218), .A3(n1052), .ZN(n1201) );
NOR2_X1 U931 ( .A1(n1244), .A2(n1249), .ZN(n1052) );
NOR2_X1 U932 ( .A1(n1067), .A2(n1066), .ZN(n1218) );
INV_X1 U933 ( .A(n1207), .ZN(n1243) );
NAND2_X1 U934 ( .A1(n1038), .A2(n1213), .ZN(n1207) );
INV_X1 U935 ( .A(n1215), .ZN(n1038) );
NAND2_X1 U936 ( .A1(n1046), .A2(n1057), .ZN(n1215) );
NOR2_X1 U937 ( .A1(n1250), .A2(n1071), .ZN(n1046) );
XNOR2_X1 U938 ( .A(G110), .B(n1200), .ZN(G12) );
NAND3_X1 U939 ( .A1(n1053), .A2(n1203), .A3(n1037), .ZN(n1200) );
NOR2_X1 U940 ( .A1(n1067), .A2(n1226), .ZN(n1037) );
INV_X1 U941 ( .A(n1066), .ZN(n1226) );
XOR2_X1 U942 ( .A(n1081), .B(n1148), .Z(n1066) );
INV_X1 U943 ( .A(G475), .ZN(n1148) );
NOR2_X1 U944 ( .A1(n1147), .A2(G902), .ZN(n1081) );
XNOR2_X1 U945 ( .A(n1251), .B(n1252), .ZN(n1147) );
XNOR2_X1 U946 ( .A(n1253), .B(n1254), .ZN(n1252) );
NAND3_X1 U947 ( .A1(n1255), .A2(n1256), .A3(KEYINPUT44), .ZN(n1253) );
NAND2_X1 U948 ( .A1(KEYINPUT38), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U949 ( .A(G104), .B(n1258), .ZN(n1257) );
NOR2_X1 U950 ( .A1(KEYINPUT20), .A2(n1259), .ZN(n1258) );
OR3_X1 U951 ( .A1(n1260), .A2(n1259), .A3(KEYINPUT38), .ZN(n1255) );
XOR2_X1 U952 ( .A(G113), .B(G122), .Z(n1259) );
XOR2_X1 U953 ( .A(KEYINPUT20), .B(G104), .Z(n1260) );
XNOR2_X1 U954 ( .A(n1261), .B(n1262), .ZN(n1251) );
NAND2_X1 U955 ( .A1(KEYINPUT36), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U956 ( .A(n1264), .B(n1265), .ZN(n1263) );
NOR2_X1 U957 ( .A1(KEYINPUT15), .A2(n1266), .ZN(n1265) );
NAND2_X1 U958 ( .A1(n1267), .A2(KEYINPUT50), .ZN(n1261) );
XOR2_X1 U959 ( .A(n1268), .B(n1269), .Z(n1267) );
NAND2_X1 U960 ( .A1(n1270), .A2(G214), .ZN(n1268) );
XNOR2_X1 U961 ( .A(n1271), .B(n1272), .ZN(n1067) );
XOR2_X1 U962 ( .A(KEYINPUT27), .B(G478), .Z(n1272) );
NAND2_X1 U963 ( .A1(n1182), .A2(n1134), .ZN(n1271) );
NAND3_X1 U964 ( .A1(n1273), .A2(n1274), .A3(n1275), .ZN(n1134) );
NAND2_X1 U965 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND2_X1 U966 ( .A1(KEYINPUT58), .A2(n1278), .ZN(n1274) );
NAND2_X1 U967 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U968 ( .A(n1276), .ZN(n1280) );
XNOR2_X1 U969 ( .A(n1277), .B(n1281), .ZN(n1279) );
NAND2_X1 U970 ( .A1(n1282), .A2(n1283), .ZN(n1273) );
INV_X1 U971 ( .A(KEYINPUT58), .ZN(n1283) );
NAND2_X1 U972 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND2_X1 U973 ( .A1(n1277), .A2(n1281), .ZN(n1285) );
OR3_X1 U974 ( .A1(n1277), .A2(n1276), .A3(n1281), .ZN(n1284) );
INV_X1 U975 ( .A(KEYINPUT7), .ZN(n1281) );
XNOR2_X1 U976 ( .A(n1286), .B(n1287), .ZN(n1276) );
XOR2_X1 U977 ( .A(G122), .B(G116), .Z(n1287) );
XNOR2_X1 U978 ( .A(G107), .B(n1288), .ZN(n1286) );
NAND3_X1 U979 ( .A1(n1289), .A2(n1041), .A3(G217), .ZN(n1277) );
AND3_X1 U980 ( .A1(n1073), .A2(n1213), .A3(n1057), .ZN(n1203) );
NOR2_X1 U981 ( .A1(n1059), .A2(n1058), .ZN(n1057) );
NOR2_X1 U982 ( .A1(n1290), .A2(n1291), .ZN(n1058) );
INV_X1 U983 ( .A(G214), .ZN(n1290) );
INV_X1 U984 ( .A(n1236), .ZN(n1059) );
XNOR2_X1 U985 ( .A(n1292), .B(n1293), .ZN(n1236) );
NOR2_X1 U986 ( .A1(n1291), .A2(n1294), .ZN(n1293) );
XNOR2_X1 U987 ( .A(G210), .B(KEYINPUT18), .ZN(n1294) );
NOR2_X1 U988 ( .A1(G902), .A2(G237), .ZN(n1291) );
NAND2_X1 U989 ( .A1(n1295), .A2(n1182), .ZN(n1292) );
XOR2_X1 U990 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U991 ( .A(n1298), .B(n1179), .Z(n1297) );
AND2_X1 U992 ( .A1(G224), .A2(n1041), .ZN(n1179) );
NOR2_X1 U993 ( .A1(KEYINPUT51), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U994 ( .A(n1177), .B(n1176), .ZN(n1299) );
XOR2_X1 U995 ( .A(G128), .B(n1300), .Z(n1176) );
INV_X1 U996 ( .A(G125), .ZN(n1177) );
NAND2_X1 U997 ( .A1(KEYINPUT21), .A2(n1181), .ZN(n1296) );
XNOR2_X1 U998 ( .A(n1301), .B(n1125), .ZN(n1181) );
XOR2_X1 U999 ( .A(G110), .B(G122), .Z(n1125) );
XNOR2_X1 U1000 ( .A(KEYINPUT4), .B(n1302), .ZN(n1301) );
NOR2_X1 U1001 ( .A1(KEYINPUT25), .A2(n1303), .ZN(n1302) );
XNOR2_X1 U1002 ( .A(n1121), .B(n1122), .ZN(n1303) );
XNOR2_X1 U1003 ( .A(n1304), .B(KEYINPUT33), .ZN(n1121) );
NAND2_X1 U1004 ( .A1(n1074), .A2(n1305), .ZN(n1213) );
NAND4_X1 U1005 ( .A1(G953), .A2(G902), .A3(n1242), .A4(n1117), .ZN(n1305) );
INV_X1 U1006 ( .A(G898), .ZN(n1117) );
NAND3_X1 U1007 ( .A1(n1242), .A2(n1041), .A3(G952), .ZN(n1074) );
NAND2_X1 U1008 ( .A1(G237), .A2(G234), .ZN(n1242) );
NOR2_X1 U1009 ( .A1(n1072), .A2(n1071), .ZN(n1073) );
AND2_X1 U1010 ( .A1(G221), .A2(n1306), .ZN(n1071) );
INV_X1 U1011 ( .A(n1250), .ZN(n1072) );
XNOR2_X1 U1012 ( .A(n1307), .B(G469), .ZN(n1250) );
NAND2_X1 U1013 ( .A1(n1308), .A2(n1182), .ZN(n1307) );
XOR2_X1 U1014 ( .A(n1309), .B(n1163), .Z(n1308) );
XNOR2_X1 U1015 ( .A(n1104), .B(n1304), .ZN(n1163) );
XOR2_X1 U1016 ( .A(G101), .B(n1310), .Z(n1304) );
XOR2_X1 U1017 ( .A(G107), .B(G104), .Z(n1310) );
XNOR2_X1 U1018 ( .A(n1311), .B(n1312), .ZN(n1104) );
XNOR2_X1 U1019 ( .A(n1313), .B(KEYINPUT12), .ZN(n1312) );
NAND2_X1 U1020 ( .A1(KEYINPUT45), .A2(n1264), .ZN(n1313) );
XOR2_X1 U1021 ( .A(n1314), .B(n1288), .Z(n1311) );
XOR2_X1 U1022 ( .A(n1269), .B(n1315), .Z(n1288) );
NAND2_X1 U1023 ( .A1(n1316), .A2(n1317), .ZN(n1309) );
NAND2_X1 U1024 ( .A1(n1318), .A2(n1164), .ZN(n1317) );
XOR2_X1 U1025 ( .A(n1319), .B(KEYINPUT43), .Z(n1316) );
OR2_X1 U1026 ( .A1(n1164), .A2(n1318), .ZN(n1319) );
XNOR2_X1 U1027 ( .A(n1320), .B(G140), .ZN(n1318) );
NAND2_X1 U1028 ( .A1(KEYINPUT49), .A2(G110), .ZN(n1320) );
NAND2_X1 U1029 ( .A1(G227), .A2(n1041), .ZN(n1164) );
INV_X1 U1030 ( .A(n1229), .ZN(n1053) );
NAND2_X1 U1031 ( .A1(n1249), .A2(n1244), .ZN(n1229) );
XNOR2_X1 U1032 ( .A(n1087), .B(n1089), .ZN(n1244) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1306), .ZN(n1089) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1182), .ZN(n1306) );
NOR2_X1 U1035 ( .A1(n1131), .A2(G902), .ZN(n1087) );
XNOR2_X1 U1036 ( .A(n1321), .B(n1322), .ZN(n1131) );
AND3_X1 U1037 ( .A1(G221), .A2(n1041), .A3(n1289), .ZN(n1322) );
XOR2_X1 U1038 ( .A(G234), .B(KEYINPUT46), .Z(n1289) );
INV_X1 U1039 ( .A(G953), .ZN(n1041) );
XNOR2_X1 U1040 ( .A(n1323), .B(n1324), .ZN(n1321) );
NAND2_X1 U1041 ( .A1(KEYINPUT37), .A2(G137), .ZN(n1324) );
NAND3_X1 U1042 ( .A1(n1325), .A2(n1326), .A3(KEYINPUT5), .ZN(n1323) );
NAND2_X1 U1043 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
XOR2_X1 U1044 ( .A(KEYINPUT3), .B(n1329), .Z(n1325) );
NOR2_X1 U1045 ( .A1(n1328), .A2(n1327), .ZN(n1329) );
XNOR2_X1 U1046 ( .A(n1330), .B(n1266), .ZN(n1327) );
INV_X1 U1047 ( .A(n1105), .ZN(n1266) );
XOR2_X1 U1048 ( .A(G125), .B(G140), .Z(n1105) );
NOR2_X1 U1049 ( .A1(G146), .A2(KEYINPUT61), .ZN(n1330) );
XNOR2_X1 U1050 ( .A(n1331), .B(n1332), .ZN(n1328) );
XOR2_X1 U1051 ( .A(KEYINPUT60), .B(G128), .Z(n1332) );
XNOR2_X1 U1052 ( .A(G119), .B(G110), .ZN(n1331) );
INV_X1 U1053 ( .A(n1245), .ZN(n1249) );
XNOR2_X1 U1054 ( .A(n1333), .B(n1084), .ZN(n1245) );
AND3_X1 U1055 ( .A1(n1334), .A2(n1335), .A3(n1182), .ZN(n1084) );
INV_X1 U1056 ( .A(G902), .ZN(n1182) );
NAND2_X1 U1057 ( .A1(n1155), .A2(n1336), .ZN(n1335) );
INV_X1 U1058 ( .A(KEYINPUT11), .ZN(n1336) );
NAND3_X1 U1059 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1155) );
NAND3_X1 U1060 ( .A1(n1340), .A2(n1341), .A3(n1122), .ZN(n1338) );
INV_X1 U1061 ( .A(n1342), .ZN(n1122) );
NAND2_X1 U1062 ( .A1(n1343), .A2(n1342), .ZN(n1337) );
XOR2_X1 U1063 ( .A(n1340), .B(n1341), .Z(n1343) );
NAND3_X1 U1064 ( .A1(n1344), .A2(n1339), .A3(KEYINPUT11), .ZN(n1334) );
OR3_X1 U1065 ( .A1(n1340), .A2(n1342), .A3(n1341), .ZN(n1339) );
NAND2_X1 U1066 ( .A1(n1340), .A2(n1345), .ZN(n1344) );
OR2_X1 U1067 ( .A1(n1341), .A2(n1342), .ZN(n1345) );
XOR2_X1 U1068 ( .A(G113), .B(n1346), .Z(n1342) );
XNOR2_X1 U1069 ( .A(n1246), .B(G116), .ZN(n1346) );
INV_X1 U1070 ( .A(G119), .ZN(n1246) );
XNOR2_X1 U1071 ( .A(n1314), .B(n1347), .ZN(n1341) );
XOR2_X1 U1072 ( .A(n1315), .B(n1300), .Z(n1347) );
XNOR2_X1 U1073 ( .A(n1264), .B(n1348), .ZN(n1300) );
NOR2_X1 U1074 ( .A1(KEYINPUT48), .A2(n1269), .ZN(n1348) );
XOR2_X1 U1075 ( .A(G143), .B(KEYINPUT30), .Z(n1269) );
INV_X1 U1076 ( .A(G146), .ZN(n1264) );
XOR2_X1 U1077 ( .A(G134), .B(G128), .Z(n1315) );
XNOR2_X1 U1078 ( .A(G137), .B(n1254), .ZN(n1314) );
XOR2_X1 U1079 ( .A(G131), .B(KEYINPUT8), .Z(n1254) );
XOR2_X1 U1080 ( .A(n1349), .B(n1350), .Z(n1340) );
INV_X1 U1081 ( .A(G101), .ZN(n1350) );
NAND2_X1 U1082 ( .A1(n1270), .A2(G210), .ZN(n1349) );
NOR2_X1 U1083 ( .A1(G953), .A2(G237), .ZN(n1270) );
NAND2_X1 U1084 ( .A1(KEYINPUT22), .A2(G472), .ZN(n1333) );
endmodule


