//Key = 0101101011110000001111010000110000011100100011100010101001001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
n1440;

XOR2_X1 U779 ( .A(G107), .B(n1080), .Z(G9) );
NOR2_X1 U780 ( .A1(KEYINPUT38), .A2(n1081), .ZN(n1080) );
NAND3_X1 U781 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(G75) );
NAND2_X1 U782 ( .A1(G952), .A2(n1085), .ZN(n1084) );
NAND4_X1 U783 ( .A1(n1086), .A2(n1087), .A3(n1088), .A4(n1089), .ZN(n1085) );
NAND4_X1 U784 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
NAND2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND3_X1 U786 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
INV_X1 U787 ( .A(KEYINPUT36), .ZN(n1097) );
INV_X1 U788 ( .A(n1099), .ZN(n1094) );
NAND3_X1 U789 ( .A1(n1100), .A2(n1101), .A3(n1099), .ZN(n1092) );
NAND2_X1 U790 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U791 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U792 ( .A1(n1096), .A2(n1106), .ZN(n1100) );
NAND2_X1 U793 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NAND2_X1 U794 ( .A1(KEYINPUT36), .A2(n1098), .ZN(n1108) );
NAND4_X1 U795 ( .A1(n1099), .A2(n1096), .A3(n1102), .A4(n1109), .ZN(n1088) );
NAND2_X1 U796 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1090), .A2(n1112), .ZN(n1111) );
NAND3_X1 U798 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
OR2_X1 U799 ( .A1(n1116), .A2(KEYINPUT63), .ZN(n1114) );
NAND3_X1 U800 ( .A1(n1116), .A2(n1117), .A3(KEYINPUT63), .ZN(n1113) );
NAND2_X1 U801 ( .A1(n1091), .A2(n1118), .ZN(n1110) );
XOR2_X1 U802 ( .A(n1119), .B(KEYINPUT34), .Z(n1086) );
NAND4_X1 U803 ( .A1(n1099), .A2(n1096), .A3(n1120), .A4(n1121), .ZN(n1119) );
NOR3_X1 U804 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1121) );
XOR2_X1 U805 ( .A(n1125), .B(KEYINPUT31), .Z(n1099) );
NAND4_X1 U806 ( .A1(n1126), .A2(n1090), .A3(n1127), .A4(n1128), .ZN(n1082) );
NOR4_X1 U807 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1122), .ZN(n1128) );
XNOR2_X1 U808 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR2_X1 U809 ( .A1(n1134), .A2(KEYINPUT16), .ZN(n1133) );
NOR2_X1 U810 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
NOR2_X1 U811 ( .A1(G902), .A2(n1137), .ZN(n1135) );
XOR2_X1 U812 ( .A(n1138), .B(n1139), .Z(n1127) );
XOR2_X1 U813 ( .A(KEYINPUT25), .B(G478), .Z(n1139) );
XOR2_X1 U814 ( .A(n1140), .B(G472), .Z(n1126) );
XOR2_X1 U815 ( .A(n1141), .B(n1142), .Z(G72) );
XOR2_X1 U816 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U817 ( .A1(n1145), .A2(n1083), .ZN(n1144) );
NOR2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND2_X1 U819 ( .A1(n1148), .A2(n1149), .ZN(n1143) );
NAND2_X1 U820 ( .A1(n1150), .A2(G953), .ZN(n1149) );
XOR2_X1 U821 ( .A(n1147), .B(KEYINPUT15), .Z(n1150) );
XOR2_X1 U822 ( .A(n1151), .B(n1152), .Z(n1148) );
XNOR2_X1 U823 ( .A(G140), .B(n1153), .ZN(n1152) );
XNOR2_X1 U824 ( .A(KEYINPUT5), .B(KEYINPUT42), .ZN(n1153) );
XOR2_X1 U825 ( .A(n1154), .B(G125), .Z(n1151) );
NAND2_X1 U826 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NAND2_X1 U827 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U828 ( .A(KEYINPUT28), .B(n1159), .Z(n1155) );
NOR2_X1 U829 ( .A1(n1157), .A2(n1158), .ZN(n1159) );
NAND2_X1 U830 ( .A1(n1160), .A2(n1161), .ZN(n1158) );
NAND2_X1 U831 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U832 ( .A1(KEYINPUT60), .A2(n1164), .ZN(n1163) );
NAND2_X1 U833 ( .A1(G131), .A2(n1165), .ZN(n1164) );
INV_X1 U834 ( .A(n1166), .ZN(n1162) );
NAND2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1160) );
NAND2_X1 U836 ( .A1(n1165), .A2(n1169), .ZN(n1167) );
NAND2_X1 U837 ( .A1(KEYINPUT60), .A2(n1166), .ZN(n1169) );
NAND2_X1 U838 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
NAND2_X1 U839 ( .A1(G134), .A2(n1172), .ZN(n1171) );
XOR2_X1 U840 ( .A(n1173), .B(KEYINPUT33), .Z(n1170) );
NAND2_X1 U841 ( .A1(G137), .A2(n1174), .ZN(n1173) );
INV_X1 U842 ( .A(KEYINPUT27), .ZN(n1165) );
NAND2_X1 U843 ( .A1(n1083), .A2(n1175), .ZN(n1141) );
NAND2_X1 U844 ( .A1(n1176), .A2(n1177), .ZN(G69) );
NAND2_X1 U845 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND2_X1 U846 ( .A1(G953), .A2(n1180), .ZN(n1179) );
NAND2_X1 U847 ( .A1(G898), .A2(G224), .ZN(n1180) );
INV_X1 U848 ( .A(n1181), .ZN(n1178) );
NAND2_X1 U849 ( .A1(n1181), .A2(n1182), .ZN(n1176) );
NAND2_X1 U850 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND2_X1 U851 ( .A1(G953), .A2(n1185), .ZN(n1184) );
XOR2_X1 U852 ( .A(n1186), .B(n1187), .Z(n1181) );
NOR2_X1 U853 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U854 ( .A(n1083), .B(KEYINPUT20), .Z(n1189) );
INV_X1 U855 ( .A(n1190), .ZN(n1188) );
NAND2_X1 U856 ( .A1(n1191), .A2(n1183), .ZN(n1186) );
INV_X1 U857 ( .A(n1192), .ZN(n1183) );
XNOR2_X1 U858 ( .A(n1193), .B(n1194), .ZN(n1191) );
NOR2_X1 U859 ( .A1(n1195), .A2(n1196), .ZN(G66) );
NOR3_X1 U860 ( .A1(n1132), .A2(n1197), .A3(n1198), .ZN(n1196) );
NOR3_X1 U861 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
AND2_X1 U862 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
NAND3_X1 U863 ( .A1(n1134), .A2(n1202), .A3(KEYINPUT10), .ZN(n1199) );
NOR2_X1 U864 ( .A1(n1195), .A2(n1203), .ZN(G63) );
NOR3_X1 U865 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1203) );
NOR3_X1 U866 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1206) );
NOR2_X1 U867 ( .A1(n1210), .A2(n1211), .ZN(n1205) );
INV_X1 U868 ( .A(n1207), .ZN(n1211) );
NOR2_X1 U869 ( .A1(n1087), .A2(n1208), .ZN(n1210) );
INV_X1 U870 ( .A(G478), .ZN(n1208) );
NOR2_X1 U871 ( .A1(n1195), .A2(n1212), .ZN(G60) );
XOR2_X1 U872 ( .A(n1213), .B(n1137), .Z(n1212) );
NOR2_X1 U873 ( .A1(n1136), .A2(n1209), .ZN(n1213) );
INV_X1 U874 ( .A(G475), .ZN(n1136) );
XOR2_X1 U875 ( .A(G104), .B(n1214), .Z(G6) );
NOR2_X1 U876 ( .A1(n1195), .A2(n1215), .ZN(G57) );
XOR2_X1 U877 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U878 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U879 ( .A(n1220), .B(n1221), .Z(n1219) );
NOR2_X1 U880 ( .A1(n1222), .A2(n1209), .ZN(n1221) );
NOR2_X1 U881 ( .A1(KEYINPUT7), .A2(n1223), .ZN(n1220) );
XOR2_X1 U882 ( .A(n1224), .B(n1225), .Z(n1216) );
XOR2_X1 U883 ( .A(n1226), .B(KEYINPUT1), .Z(n1225) );
NOR2_X1 U884 ( .A1(n1195), .A2(n1227), .ZN(G54) );
XOR2_X1 U885 ( .A(n1228), .B(n1229), .Z(n1227) );
NOR2_X1 U886 ( .A1(n1230), .A2(n1209), .ZN(n1229) );
NAND2_X1 U887 ( .A1(G902), .A2(n1202), .ZN(n1209) );
INV_X1 U888 ( .A(G469), .ZN(n1230) );
NOR2_X1 U889 ( .A1(n1231), .A2(n1232), .ZN(n1228) );
XOR2_X1 U890 ( .A(n1233), .B(KEYINPUT52), .Z(n1232) );
NAND2_X1 U891 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U892 ( .A(n1236), .B(n1237), .Z(n1234) );
NOR3_X1 U893 ( .A1(n1238), .A2(n1239), .A3(n1240), .ZN(n1231) );
NOR2_X1 U894 ( .A1(n1236), .A2(n1241), .ZN(n1240) );
INV_X1 U895 ( .A(n1242), .ZN(n1239) );
XOR2_X1 U896 ( .A(KEYINPUT61), .B(n1235), .Z(n1238) );
XNOR2_X1 U897 ( .A(n1243), .B(n1244), .ZN(n1235) );
XOR2_X1 U898 ( .A(n1245), .B(n1246), .Z(n1243) );
NOR2_X1 U899 ( .A1(n1195), .A2(n1247), .ZN(G51) );
XOR2_X1 U900 ( .A(n1248), .B(n1249), .Z(n1247) );
NOR2_X1 U901 ( .A1(KEYINPUT41), .A2(n1250), .ZN(n1249) );
XOR2_X1 U902 ( .A(n1251), .B(n1252), .Z(n1250) );
NOR2_X1 U903 ( .A1(KEYINPUT0), .A2(n1253), .ZN(n1252) );
NOR2_X1 U904 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XOR2_X1 U905 ( .A(KEYINPUT53), .B(n1256), .Z(n1255) );
NOR2_X1 U906 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
AND2_X1 U907 ( .A1(n1257), .A2(n1258), .ZN(n1254) );
XNOR2_X1 U908 ( .A(n1259), .B(n1260), .ZN(n1258) );
NAND3_X1 U909 ( .A1(G902), .A2(n1261), .A3(n1262), .ZN(n1248) );
XOR2_X1 U910 ( .A(n1202), .B(KEYINPUT32), .Z(n1262) );
INV_X1 U911 ( .A(n1087), .ZN(n1202) );
NOR2_X1 U912 ( .A1(n1190), .A2(n1175), .ZN(n1087) );
NAND4_X1 U913 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1175) );
AND4_X1 U914 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1266) );
NOR4_X1 U915 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1265) );
NOR2_X1 U916 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NAND4_X1 U917 ( .A1(n1277), .A2(n1278), .A3(n1279), .A4(n1280), .ZN(n1276) );
INV_X1 U918 ( .A(n1281), .ZN(n1277) );
INV_X1 U919 ( .A(KEYINPUT58), .ZN(n1275) );
NOR2_X1 U920 ( .A1(KEYINPUT58), .A2(n1282), .ZN(n1273) );
NOR2_X1 U921 ( .A1(n1283), .A2(n1284), .ZN(n1272) );
INV_X1 U922 ( .A(KEYINPUT35), .ZN(n1283) );
NOR4_X1 U923 ( .A1(KEYINPUT35), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1271) );
NAND3_X1 U924 ( .A1(n1288), .A2(n1289), .A3(n1290), .ZN(n1285) );
NAND2_X1 U925 ( .A1(n1291), .A2(n1292), .ZN(n1190) );
AND4_X1 U926 ( .A1(n1081), .A2(n1293), .A3(n1294), .A4(n1295), .ZN(n1292) );
NAND3_X1 U927 ( .A1(n1296), .A2(n1102), .A3(n1297), .ZN(n1081) );
NOR4_X1 U928 ( .A1(n1298), .A2(n1299), .A3(n1214), .A4(n1300), .ZN(n1291) );
NOR2_X1 U929 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NOR2_X1 U930 ( .A1(n1296), .A2(n1303), .ZN(n1301) );
XOR2_X1 U931 ( .A(n1104), .B(KEYINPUT11), .Z(n1303) );
AND3_X1 U932 ( .A1(n1297), .A2(n1102), .A3(n1278), .ZN(n1214) );
AND2_X1 U933 ( .A1(KEYINPUT3), .A2(n1304), .ZN(n1299) );
NOR3_X1 U934 ( .A1(KEYINPUT3), .A2(n1305), .A3(n1306), .ZN(n1298) );
NOR2_X1 U935 ( .A1(n1083), .A2(G952), .ZN(n1195) );
NAND2_X1 U936 ( .A1(n1307), .A2(n1308), .ZN(G48) );
NAND2_X1 U937 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
XOR2_X1 U938 ( .A(KEYINPUT29), .B(n1311), .Z(n1307) );
NOR2_X1 U939 ( .A1(n1309), .A2(n1310), .ZN(n1311) );
XOR2_X1 U940 ( .A(KEYINPUT19), .B(G146), .Z(n1310) );
INV_X1 U941 ( .A(n1282), .ZN(n1309) );
NAND3_X1 U942 ( .A1(n1278), .A2(n1279), .A3(n1312), .ZN(n1282) );
XOR2_X1 U943 ( .A(n1313), .B(n1284), .Z(G45) );
NAND3_X1 U944 ( .A1(n1314), .A2(n1098), .A3(n1312), .ZN(n1284) );
XNOR2_X1 U945 ( .A(G140), .B(n1267), .ZN(G42) );
NAND3_X1 U946 ( .A1(n1278), .A2(n1315), .A3(n1316), .ZN(n1267) );
XOR2_X1 U947 ( .A(n1263), .B(n1317), .Z(G39) );
NAND2_X1 U948 ( .A1(KEYINPUT45), .A2(G137), .ZN(n1317) );
NAND4_X1 U949 ( .A1(n1318), .A2(n1316), .A3(n1096), .A4(n1319), .ZN(n1263) );
XOR2_X1 U950 ( .A(n1174), .B(n1264), .Z(G36) );
NAND3_X1 U951 ( .A1(n1098), .A2(n1296), .A3(n1316), .ZN(n1264) );
XOR2_X1 U952 ( .A(n1168), .B(n1270), .Z(G33) );
NAND3_X1 U953 ( .A1(n1278), .A2(n1098), .A3(n1316), .ZN(n1270) );
AND2_X1 U954 ( .A1(n1312), .A2(n1090), .ZN(n1316) );
NOR2_X1 U955 ( .A1(n1124), .A2(n1120), .ZN(n1090) );
INV_X1 U956 ( .A(n1320), .ZN(n1120) );
INV_X1 U957 ( .A(n1104), .ZN(n1278) );
XOR2_X1 U958 ( .A(n1321), .B(n1269), .Z(G30) );
NAND3_X1 U959 ( .A1(n1279), .A2(n1296), .A3(n1312), .ZN(n1269) );
INV_X1 U960 ( .A(n1287), .ZN(n1312) );
NAND2_X1 U961 ( .A1(n1280), .A2(n1281), .ZN(n1287) );
INV_X1 U962 ( .A(n1105), .ZN(n1296) );
XOR2_X1 U963 ( .A(n1226), .B(n1295), .Z(G3) );
NAND3_X1 U964 ( .A1(n1096), .A2(n1297), .A3(n1098), .ZN(n1295) );
XOR2_X1 U965 ( .A(n1260), .B(n1268), .Z(G27) );
NAND4_X1 U966 ( .A1(n1118), .A2(n1281), .A3(n1091), .A4(n1322), .ZN(n1268) );
NOR2_X1 U967 ( .A1(n1107), .A2(n1104), .ZN(n1322) );
NAND2_X1 U968 ( .A1(n1323), .A2(n1324), .ZN(n1281) );
NAND4_X1 U969 ( .A1(G902), .A2(G953), .A3(n1125), .A4(n1147), .ZN(n1324) );
INV_X1 U970 ( .A(G900), .ZN(n1147) );
XOR2_X1 U971 ( .A(G122), .B(n1304), .Z(G24) );
NOR2_X1 U972 ( .A1(n1305), .A2(n1325), .ZN(n1304) );
NAND3_X1 U973 ( .A1(n1091), .A2(n1102), .A3(n1314), .ZN(n1305) );
NOR3_X1 U974 ( .A1(n1326), .A2(n1327), .A3(n1288), .ZN(n1314) );
INV_X1 U975 ( .A(n1123), .ZN(n1102) );
NAND2_X1 U976 ( .A1(n1328), .A2(n1329), .ZN(n1123) );
XOR2_X1 U977 ( .A(n1330), .B(n1294), .Z(G21) );
NAND4_X1 U978 ( .A1(n1279), .A2(n1096), .A3(n1091), .A4(n1306), .ZN(n1294) );
AND3_X1 U979 ( .A1(n1118), .A2(n1319), .A3(n1318), .ZN(n1279) );
XOR2_X1 U980 ( .A(G116), .B(n1331), .Z(G18) );
NOR2_X1 U981 ( .A1(n1105), .A2(n1302), .ZN(n1331) );
NAND2_X1 U982 ( .A1(n1327), .A2(n1290), .ZN(n1105) );
XOR2_X1 U983 ( .A(G113), .B(n1332), .Z(G15) );
NOR2_X1 U984 ( .A1(n1104), .A2(n1302), .ZN(n1332) );
NAND4_X1 U985 ( .A1(n1098), .A2(n1091), .A3(n1118), .A4(n1306), .ZN(n1302) );
INV_X1 U986 ( .A(n1288), .ZN(n1118) );
INV_X1 U987 ( .A(n1122), .ZN(n1091) );
NAND2_X1 U988 ( .A1(n1117), .A2(n1333), .ZN(n1122) );
INV_X1 U989 ( .A(n1286), .ZN(n1098) );
NAND2_X1 U990 ( .A1(n1318), .A2(n1328), .ZN(n1286) );
XOR2_X1 U991 ( .A(n1319), .B(KEYINPUT46), .Z(n1328) );
NAND2_X1 U992 ( .A1(n1326), .A2(n1289), .ZN(n1104) );
INV_X1 U993 ( .A(n1327), .ZN(n1289) );
XOR2_X1 U994 ( .A(n1334), .B(n1293), .Z(G12) );
NAND3_X1 U995 ( .A1(n1315), .A2(n1297), .A3(n1096), .ZN(n1293) );
AND2_X1 U996 ( .A1(n1327), .A2(n1335), .ZN(n1096) );
XOR2_X1 U997 ( .A(KEYINPUT37), .B(n1290), .Z(n1335) );
INV_X1 U998 ( .A(n1326), .ZN(n1290) );
XOR2_X1 U999 ( .A(n1336), .B(G478), .Z(n1326) );
NAND2_X1 U1000 ( .A1(KEYINPUT9), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1001 ( .A(KEYINPUT14), .B(n1204), .Z(n1337) );
INV_X1 U1002 ( .A(n1138), .ZN(n1204) );
NAND2_X1 U1003 ( .A1(n1207), .A2(n1201), .ZN(n1138) );
XOR2_X1 U1004 ( .A(n1338), .B(n1339), .Z(n1207) );
XNOR2_X1 U1005 ( .A(n1340), .B(n1341), .ZN(n1339) );
NAND2_X1 U1006 ( .A1(KEYINPUT40), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1007 ( .A(n1343), .B(n1344), .Z(n1342) );
XOR2_X1 U1008 ( .A(G116), .B(n1345), .Z(n1344) );
NAND2_X1 U1009 ( .A1(KEYINPUT21), .A2(n1346), .ZN(n1343) );
XOR2_X1 U1010 ( .A(n1347), .B(G143), .Z(n1338) );
NAND3_X1 U1011 ( .A1(G234), .A2(n1083), .A3(G217), .ZN(n1347) );
NOR2_X1 U1012 ( .A1(n1348), .A2(n1129), .ZN(n1327) );
NOR3_X1 U1013 ( .A1(G475), .A2(G902), .A3(n1137), .ZN(n1129) );
AND2_X1 U1014 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
OR2_X1 U1015 ( .A1(n1137), .A2(G902), .ZN(n1350) );
XNOR2_X1 U1016 ( .A(n1351), .B(n1352), .ZN(n1137) );
XOR2_X1 U1017 ( .A(G104), .B(n1353), .Z(n1352) );
NOR2_X1 U1018 ( .A1(KEYINPUT47), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1019 ( .A(n1355), .B(n1356), .Z(n1354) );
XOR2_X1 U1020 ( .A(n1357), .B(n1245), .Z(n1356) );
INV_X1 U1021 ( .A(n1358), .ZN(n1245) );
XOR2_X1 U1022 ( .A(n1359), .B(G131), .Z(n1355) );
NAND2_X1 U1023 ( .A1(n1360), .A2(G214), .ZN(n1359) );
XOR2_X1 U1024 ( .A(G113), .B(n1345), .Z(n1351) );
XOR2_X1 U1025 ( .A(KEYINPUT48), .B(G475), .Z(n1349) );
NOR3_X1 U1026 ( .A1(n1115), .A2(n1325), .A3(n1288), .ZN(n1297) );
NAND2_X1 U1027 ( .A1(n1124), .A2(n1320), .ZN(n1288) );
NAND2_X1 U1028 ( .A1(n1361), .A2(n1362), .ZN(n1320) );
XNOR2_X1 U1029 ( .A(G214), .B(KEYINPUT18), .ZN(n1361) );
XNOR2_X1 U1030 ( .A(n1363), .B(n1261), .ZN(n1124) );
AND2_X1 U1031 ( .A1(G210), .A2(n1362), .ZN(n1261) );
NAND2_X1 U1032 ( .A1(n1364), .A2(n1201), .ZN(n1362) );
INV_X1 U1033 ( .A(G237), .ZN(n1364) );
NAND2_X1 U1034 ( .A1(n1365), .A2(n1201), .ZN(n1363) );
XOR2_X1 U1035 ( .A(n1366), .B(n1367), .Z(n1365) );
NAND2_X1 U1036 ( .A1(KEYINPUT62), .A2(n1251), .ZN(n1367) );
XOR2_X1 U1037 ( .A(n1193), .B(n1368), .Z(n1251) );
NOR2_X1 U1038 ( .A1(KEYINPUT13), .A2(n1194), .ZN(n1368) );
XNOR2_X1 U1039 ( .A(n1369), .B(G113), .ZN(n1194) );
NAND3_X1 U1040 ( .A1(n1370), .A2(n1371), .A3(n1372), .ZN(n1369) );
NAND2_X1 U1041 ( .A1(G116), .A2(n1373), .ZN(n1372) );
INV_X1 U1042 ( .A(KEYINPUT57), .ZN(n1373) );
NAND3_X1 U1043 ( .A1(KEYINPUT57), .A2(n1374), .A3(n1330), .ZN(n1371) );
OR2_X1 U1044 ( .A1(n1330), .A2(n1374), .ZN(n1370) );
NOR2_X1 U1045 ( .A1(n1375), .A2(G116), .ZN(n1374) );
INV_X1 U1046 ( .A(KEYINPUT8), .ZN(n1375) );
XOR2_X1 U1047 ( .A(n1376), .B(n1377), .Z(n1193) );
XOR2_X1 U1048 ( .A(G101), .B(n1378), .Z(n1377) );
XOR2_X1 U1049 ( .A(G110), .B(G104), .Z(n1378) );
XOR2_X1 U1050 ( .A(n1379), .B(n1380), .Z(n1376) );
NAND2_X1 U1051 ( .A1(KEYINPUT4), .A2(n1345), .ZN(n1379) );
INV_X1 U1052 ( .A(G122), .ZN(n1345) );
NAND2_X1 U1053 ( .A1(n1381), .A2(n1382), .ZN(n1366) );
NAND2_X1 U1054 ( .A1(n1257), .A2(n1383), .ZN(n1382) );
XOR2_X1 U1055 ( .A(n1384), .B(KEYINPUT55), .Z(n1381) );
OR2_X1 U1056 ( .A1(n1383), .A2(n1257), .ZN(n1384) );
NOR2_X1 U1057 ( .A1(n1185), .A2(G953), .ZN(n1257) );
INV_X1 U1058 ( .A(G224), .ZN(n1185) );
XNOR2_X1 U1059 ( .A(n1385), .B(G125), .ZN(n1383) );
NAND2_X1 U1060 ( .A1(KEYINPUT54), .A2(n1259), .ZN(n1385) );
XOR2_X1 U1061 ( .A(n1386), .B(G128), .Z(n1259) );
INV_X1 U1062 ( .A(n1306), .ZN(n1325) );
NAND2_X1 U1063 ( .A1(n1323), .A2(n1387), .ZN(n1306) );
NAND3_X1 U1064 ( .A1(n1192), .A2(n1125), .A3(G902), .ZN(n1387) );
NOR2_X1 U1065 ( .A1(n1083), .A2(G898), .ZN(n1192) );
NAND3_X1 U1066 ( .A1(n1125), .A2(n1083), .A3(G952), .ZN(n1323) );
NAND2_X1 U1067 ( .A1(G237), .A2(G234), .ZN(n1125) );
INV_X1 U1068 ( .A(n1280), .ZN(n1115) );
NOR2_X1 U1069 ( .A1(n1117), .A2(n1116), .ZN(n1280) );
INV_X1 U1070 ( .A(n1333), .ZN(n1116) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1388), .ZN(n1333) );
XNOR2_X1 U1072 ( .A(KEYINPUT6), .B(n1389), .ZN(n1388) );
XOR2_X1 U1073 ( .A(n1390), .B(G469), .Z(n1117) );
NAND2_X1 U1074 ( .A1(n1391), .A2(n1201), .ZN(n1390) );
XOR2_X1 U1075 ( .A(n1392), .B(n1393), .Z(n1391) );
XOR2_X1 U1076 ( .A(n1394), .B(n1244), .Z(n1393) );
XOR2_X1 U1077 ( .A(n1395), .B(n1226), .Z(n1244) );
NAND3_X1 U1078 ( .A1(n1396), .A2(n1397), .A3(n1398), .ZN(n1395) );
NAND2_X1 U1079 ( .A1(n1346), .A2(G104), .ZN(n1398) );
NAND2_X1 U1080 ( .A1(KEYINPUT22), .A2(n1399), .ZN(n1397) );
NAND2_X1 U1081 ( .A1(n1400), .A2(n1380), .ZN(n1399) );
INV_X1 U1082 ( .A(n1346), .ZN(n1380) );
XNOR2_X1 U1083 ( .A(KEYINPUT2), .B(G104), .ZN(n1400) );
NAND2_X1 U1084 ( .A1(n1401), .A2(n1402), .ZN(n1396) );
INV_X1 U1085 ( .A(KEYINPUT22), .ZN(n1402) );
NAND2_X1 U1086 ( .A1(n1403), .A2(n1404), .ZN(n1401) );
OR3_X1 U1087 ( .A1(n1346), .A2(G104), .A3(KEYINPUT2), .ZN(n1404) );
XNOR2_X1 U1088 ( .A(G107), .B(KEYINPUT59), .ZN(n1346) );
NAND2_X1 U1089 ( .A1(KEYINPUT2), .A2(G104), .ZN(n1403) );
XOR2_X1 U1090 ( .A(n1405), .B(n1406), .Z(n1392) );
NOR2_X1 U1091 ( .A1(KEYINPUT26), .A2(n1407), .ZN(n1406) );
INV_X1 U1092 ( .A(n1157), .ZN(n1407) );
XNOR2_X1 U1093 ( .A(n1321), .B(n1358), .ZN(n1157) );
XOR2_X1 U1094 ( .A(n1408), .B(G134), .Z(n1405) );
NAND2_X1 U1095 ( .A1(n1409), .A2(n1242), .ZN(n1408) );
NAND2_X1 U1096 ( .A1(n1236), .A2(n1241), .ZN(n1242) );
XOR2_X1 U1097 ( .A(n1410), .B(KEYINPUT49), .Z(n1409) );
NAND2_X1 U1098 ( .A1(n1411), .A2(n1237), .ZN(n1410) );
INV_X1 U1099 ( .A(n1241), .ZN(n1237) );
XOR2_X1 U1100 ( .A(n1334), .B(G140), .Z(n1241) );
XNOR2_X1 U1101 ( .A(n1236), .B(KEYINPUT39), .ZN(n1411) );
NOR2_X1 U1102 ( .A1(n1146), .A2(G953), .ZN(n1236) );
INV_X1 U1103 ( .A(G227), .ZN(n1146) );
INV_X1 U1104 ( .A(n1107), .ZN(n1315) );
NAND2_X1 U1105 ( .A1(n1319), .A2(n1329), .ZN(n1107) );
INV_X1 U1106 ( .A(n1318), .ZN(n1329) );
XNOR2_X1 U1107 ( .A(n1412), .B(n1140), .ZN(n1318) );
NAND2_X1 U1108 ( .A1(n1413), .A2(n1201), .ZN(n1140) );
XOR2_X1 U1109 ( .A(n1218), .B(n1414), .Z(n1413) );
XNOR2_X1 U1110 ( .A(n1415), .B(n1223), .ZN(n1414) );
XOR2_X1 U1111 ( .A(n1416), .B(n1417), .Z(n1223) );
XOR2_X1 U1112 ( .A(KEYINPUT51), .B(G119), .Z(n1417) );
XNOR2_X1 U1113 ( .A(G113), .B(G116), .ZN(n1416) );
NOR2_X1 U1114 ( .A1(n1418), .A2(n1419), .ZN(n1415) );
XOR2_X1 U1115 ( .A(KEYINPUT56), .B(n1420), .Z(n1419) );
NOR2_X1 U1116 ( .A1(n1226), .A2(n1224), .ZN(n1420) );
AND2_X1 U1117 ( .A1(n1226), .A2(n1224), .ZN(n1418) );
NAND2_X1 U1118 ( .A1(n1360), .A2(G210), .ZN(n1224) );
NOR2_X1 U1119 ( .A1(G953), .A2(G237), .ZN(n1360) );
INV_X1 U1120 ( .A(G101), .ZN(n1226) );
XNOR2_X1 U1121 ( .A(n1386), .B(n1246), .ZN(n1218) );
XNOR2_X1 U1122 ( .A(n1394), .B(n1341), .ZN(n1246) );
XOR2_X1 U1123 ( .A(n1321), .B(n1174), .Z(n1341) );
INV_X1 U1124 ( .A(G134), .ZN(n1174) );
INV_X1 U1125 ( .A(G128), .ZN(n1321) );
XOR2_X1 U1126 ( .A(n1168), .B(G137), .Z(n1394) );
INV_X1 U1127 ( .A(G131), .ZN(n1168) );
NAND2_X1 U1128 ( .A1(KEYINPUT23), .A2(n1358), .ZN(n1386) );
XNOR2_X1 U1129 ( .A(n1313), .B(G146), .ZN(n1358) );
INV_X1 U1130 ( .A(G143), .ZN(n1313) );
NAND2_X1 U1131 ( .A1(KEYINPUT44), .A2(n1222), .ZN(n1412) );
INV_X1 U1132 ( .A(G472), .ZN(n1222) );
XOR2_X1 U1133 ( .A(n1132), .B(n1134), .Z(n1319) );
AND2_X1 U1134 ( .A1(G217), .A2(n1389), .ZN(n1134) );
NAND2_X1 U1135 ( .A1(G234), .A2(n1201), .ZN(n1389) );
AND2_X1 U1136 ( .A1(n1200), .A2(n1201), .ZN(n1132) );
INV_X1 U1137 ( .A(G902), .ZN(n1201) );
XNOR2_X1 U1138 ( .A(n1421), .B(n1422), .ZN(n1200) );
XOR2_X1 U1139 ( .A(n1423), .B(n1424), .Z(n1422) );
NAND2_X1 U1140 ( .A1(n1425), .A2(n1426), .ZN(n1424) );
OR2_X1 U1141 ( .A1(n1427), .A2(n1172), .ZN(n1426) );
XOR2_X1 U1142 ( .A(n1428), .B(KEYINPUT43), .Z(n1425) );
NAND2_X1 U1143 ( .A1(n1172), .A2(n1427), .ZN(n1428) );
NAND3_X1 U1144 ( .A1(G234), .A2(n1083), .A3(G221), .ZN(n1427) );
INV_X1 U1145 ( .A(G953), .ZN(n1083) );
INV_X1 U1146 ( .A(G137), .ZN(n1172) );
INV_X1 U1147 ( .A(G146), .ZN(n1423) );
NAND2_X1 U1148 ( .A1(n1429), .A2(n1430), .ZN(n1421) );
NAND2_X1 U1149 ( .A1(n1431), .A2(n1432), .ZN(n1430) );
INV_X1 U1150 ( .A(KEYINPUT12), .ZN(n1432) );
XOR2_X1 U1151 ( .A(n1433), .B(n1357), .Z(n1431) );
XNOR2_X1 U1152 ( .A(n1260), .B(n1434), .ZN(n1357) );
NAND2_X1 U1153 ( .A1(n1435), .A2(KEYINPUT12), .ZN(n1429) );
XOR2_X1 U1154 ( .A(n1433), .B(n1436), .Z(n1435) );
NAND2_X1 U1155 ( .A1(n1434), .A2(n1260), .ZN(n1436) );
INV_X1 U1156 ( .A(G125), .ZN(n1260) );
XOR2_X1 U1157 ( .A(G140), .B(KEYINPUT30), .Z(n1434) );
NAND2_X1 U1158 ( .A1(n1437), .A2(KEYINPUT50), .ZN(n1433) );
XOR2_X1 U1159 ( .A(n1438), .B(n1439), .Z(n1437) );
XOR2_X1 U1160 ( .A(G110), .B(n1440), .Z(n1439) );
NOR2_X1 U1161 ( .A1(G128), .A2(KEYINPUT24), .ZN(n1440) );
XOR2_X1 U1162 ( .A(n1330), .B(KEYINPUT17), .Z(n1438) );
INV_X1 U1163 ( .A(G119), .ZN(n1330) );
INV_X1 U1164 ( .A(G110), .ZN(n1334) );
endmodule


