//Key = 0000001100100110101010010101001101011010000101111000000010111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
n1468;

XNOR2_X1 U798 ( .A(G107), .B(n1108), .ZN(G9) );
NAND2_X1 U799 ( .A1(KEYINPUT61), .A2(n1109), .ZN(n1108) );
INV_X1 U800 ( .A(n1110), .ZN(n1109) );
NOR2_X1 U801 ( .A1(n1111), .A2(n1112), .ZN(G75) );
NOR4_X1 U802 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1112) );
XOR2_X1 U803 ( .A(KEYINPUT20), .B(n1117), .Z(n1114) );
NAND4_X1 U804 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1113) );
NAND3_X1 U805 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1119) );
NAND2_X1 U806 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND4_X1 U807 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1126) );
NAND2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1125) );
NAND2_X1 U809 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U810 ( .A1(n1130), .A2(n1135), .ZN(n1134) );
NAND2_X1 U811 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
NAND2_X1 U812 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XOR2_X1 U813 ( .A(KEYINPUT12), .B(n1140), .Z(n1139) );
NAND2_X1 U814 ( .A1(n1127), .A2(n1141), .ZN(n1133) );
NAND2_X1 U815 ( .A1(n1127), .A2(n1142), .ZN(n1118) );
NAND2_X1 U816 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NAND2_X1 U817 ( .A1(n1124), .A2(n1145), .ZN(n1144) );
NAND2_X1 U818 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND3_X1 U819 ( .A1(n1130), .A2(n1148), .A3(n1122), .ZN(n1147) );
NAND2_X1 U820 ( .A1(n1131), .A2(n1149), .ZN(n1146) );
NAND2_X1 U821 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND3_X1 U822 ( .A1(n1152), .A2(n1122), .A3(KEYINPUT63), .ZN(n1151) );
NAND2_X1 U823 ( .A1(n1130), .A2(n1153), .ZN(n1150) );
OR2_X1 U824 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U825 ( .A1(n1156), .A2(n1157), .ZN(n1143) );
INV_X1 U826 ( .A(KEYINPUT63), .ZN(n1157) );
NAND4_X1 U827 ( .A1(n1124), .A2(n1152), .A3(n1131), .A4(n1122), .ZN(n1156) );
INV_X1 U828 ( .A(n1158), .ZN(n1124) );
NOR3_X1 U829 ( .A1(n1159), .A2(G953), .A3(n1160), .ZN(n1111) );
INV_X1 U830 ( .A(n1120), .ZN(n1160) );
NAND4_X1 U831 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1120) );
NOR4_X1 U832 ( .A1(n1138), .A2(n1128), .A3(n1165), .A4(n1166), .ZN(n1164) );
XNOR2_X1 U833 ( .A(n1167), .B(n1168), .ZN(n1166) );
NAND2_X1 U834 ( .A1(KEYINPUT23), .A2(n1169), .ZN(n1167) );
XOR2_X1 U835 ( .A(n1170), .B(n1171), .Z(n1165) );
NOR2_X1 U836 ( .A1(G472), .A2(KEYINPUT1), .ZN(n1171) );
NOR2_X1 U837 ( .A1(n1172), .A2(n1173), .ZN(n1163) );
XNOR2_X1 U838 ( .A(G478), .B(n1174), .ZN(n1173) );
NAND2_X1 U839 ( .A1(KEYINPUT60), .A2(n1175), .ZN(n1174) );
XNOR2_X1 U840 ( .A(G475), .B(n1176), .ZN(n1172) );
NAND2_X1 U841 ( .A1(KEYINPUT16), .A2(n1177), .ZN(n1176) );
XOR2_X1 U842 ( .A(KEYINPUT42), .B(n1178), .Z(n1162) );
NOR3_X1 U843 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1178) );
NOR3_X1 U844 ( .A1(n1182), .A2(KEYINPUT24), .A3(n1183), .ZN(n1181) );
AND2_X1 U845 ( .A1(n1182), .A2(KEYINPUT24), .ZN(n1180) );
XOR2_X1 U846 ( .A(n1184), .B(G469), .Z(n1161) );
NAND2_X1 U847 ( .A1(KEYINPUT56), .A2(n1185), .ZN(n1184) );
XNOR2_X1 U848 ( .A(KEYINPUT4), .B(n1115), .ZN(n1159) );
XOR2_X1 U849 ( .A(n1186), .B(n1187), .Z(G72) );
NOR2_X1 U850 ( .A1(n1188), .A2(n1121), .ZN(n1187) );
AND2_X1 U851 ( .A1(G227), .A2(G900), .ZN(n1188) );
XOR2_X1 U852 ( .A(n1189), .B(n1190), .Z(n1186) );
NOR2_X1 U853 ( .A1(G953), .A2(n1191), .ZN(n1190) );
NOR3_X1 U854 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1191) );
NAND2_X1 U855 ( .A1(KEYINPUT13), .A2(n1195), .ZN(n1189) );
NAND2_X1 U856 ( .A1(n1196), .A2(n1197), .ZN(n1195) );
NAND2_X1 U857 ( .A1(n1198), .A2(G953), .ZN(n1197) );
XOR2_X1 U858 ( .A(n1199), .B(n1200), .Z(n1196) );
XOR2_X1 U859 ( .A(n1201), .B(n1202), .Z(n1200) );
NOR2_X1 U860 ( .A1(G125), .A2(KEYINPUT21), .ZN(n1202) );
XNOR2_X1 U861 ( .A(G140), .B(KEYINPUT25), .ZN(n1199) );
NAND2_X1 U862 ( .A1(n1203), .A2(n1204), .ZN(G69) );
NAND3_X1 U863 ( .A1(n1205), .A2(n1206), .A3(G953), .ZN(n1204) );
XOR2_X1 U864 ( .A(n1207), .B(KEYINPUT49), .Z(n1203) );
NAND3_X1 U865 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
NAND2_X1 U866 ( .A1(n1211), .A2(n1206), .ZN(n1210) );
OR3_X1 U867 ( .A1(n1206), .A2(n1211), .A3(G953), .ZN(n1209) );
NAND2_X1 U868 ( .A1(G953), .A2(n1212), .ZN(n1208) );
OR2_X1 U869 ( .A1(n1206), .A2(n1205), .ZN(n1212) );
NAND2_X1 U870 ( .A1(G898), .A2(G224), .ZN(n1205) );
NAND2_X1 U871 ( .A1(n1213), .A2(n1214), .ZN(n1206) );
NAND2_X1 U872 ( .A1(G953), .A2(n1215), .ZN(n1214) );
XOR2_X1 U873 ( .A(n1216), .B(n1217), .Z(n1213) );
NOR2_X1 U874 ( .A1(KEYINPUT29), .A2(n1218), .ZN(n1216) );
NOR2_X1 U875 ( .A1(n1219), .A2(n1220), .ZN(G66) );
NOR2_X1 U876 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
XOR2_X1 U877 ( .A(n1223), .B(n1224), .Z(n1222) );
NOR2_X1 U878 ( .A1(n1182), .A2(n1225), .ZN(n1224) );
NOR2_X1 U879 ( .A1(KEYINPUT53), .A2(n1226), .ZN(n1223) );
AND2_X1 U880 ( .A1(n1226), .A2(KEYINPUT53), .ZN(n1221) );
NOR2_X1 U881 ( .A1(n1219), .A2(n1227), .ZN(G63) );
XOR2_X1 U882 ( .A(n1228), .B(n1229), .Z(n1227) );
NOR2_X1 U883 ( .A1(n1230), .A2(n1225), .ZN(n1229) );
NOR2_X1 U884 ( .A1(n1219), .A2(n1231), .ZN(G60) );
XOR2_X1 U885 ( .A(n1232), .B(n1233), .Z(n1231) );
NOR2_X1 U886 ( .A1(n1234), .A2(n1225), .ZN(n1233) );
XNOR2_X1 U887 ( .A(G104), .B(n1235), .ZN(G6) );
NOR3_X1 U888 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(G57) );
NOR2_X1 U889 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XNOR2_X1 U890 ( .A(n1241), .B(n1242), .ZN(n1240) );
XOR2_X1 U891 ( .A(KEYINPUT6), .B(KEYINPUT27), .Z(n1242) );
XNOR2_X1 U892 ( .A(KEYINPUT0), .B(n1243), .ZN(n1239) );
NOR2_X1 U893 ( .A1(n1241), .A2(n1244), .ZN(n1237) );
XNOR2_X1 U894 ( .A(KEYINPUT0), .B(G101), .ZN(n1244) );
XOR2_X1 U895 ( .A(n1245), .B(n1246), .Z(n1241) );
XOR2_X1 U896 ( .A(n1247), .B(n1248), .Z(n1246) );
NAND3_X1 U897 ( .A1(n1249), .A2(n1250), .A3(G472), .ZN(n1247) );
NAND2_X1 U898 ( .A1(KEYINPUT38), .A2(n1225), .ZN(n1250) );
NAND2_X1 U899 ( .A1(n1251), .A2(n1252), .ZN(n1249) );
INV_X1 U900 ( .A(KEYINPUT38), .ZN(n1252) );
NAND3_X1 U901 ( .A1(n1117), .A2(G902), .A3(n1211), .ZN(n1251) );
NAND2_X1 U902 ( .A1(n1253), .A2(KEYINPUT47), .ZN(n1245) );
XOR2_X1 U903 ( .A(n1254), .B(n1255), .Z(n1253) );
XNOR2_X1 U904 ( .A(G143), .B(n1256), .ZN(n1254) );
NOR2_X1 U905 ( .A1(KEYINPUT32), .A2(n1257), .ZN(n1256) );
XNOR2_X1 U906 ( .A(G113), .B(n1258), .ZN(n1257) );
NOR2_X1 U907 ( .A1(n1121), .A2(n1259), .ZN(n1236) );
XNOR2_X1 U908 ( .A(KEYINPUT39), .B(n1115), .ZN(n1259) );
INV_X1 U909 ( .A(G952), .ZN(n1115) );
NOR3_X1 U910 ( .A1(n1219), .A2(n1260), .A3(n1261), .ZN(G54) );
NOR2_X1 U911 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NOR2_X1 U912 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
NOR2_X1 U913 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NOR2_X1 U914 ( .A1(n1268), .A2(n1269), .ZN(n1264) );
NOR2_X1 U915 ( .A1(n1270), .A2(n1271), .ZN(n1260) );
NOR2_X1 U916 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
NOR2_X1 U917 ( .A1(n1267), .A2(n1269), .ZN(n1273) );
XNOR2_X1 U918 ( .A(KEYINPUT59), .B(n1274), .ZN(n1269) );
NOR2_X1 U919 ( .A1(n1268), .A2(n1266), .ZN(n1272) );
XNOR2_X1 U920 ( .A(n1274), .B(KEYINPUT11), .ZN(n1266) );
NOR2_X1 U921 ( .A1(n1225), .A2(n1275), .ZN(n1274) );
INV_X1 U922 ( .A(G469), .ZN(n1275) );
INV_X1 U923 ( .A(n1267), .ZN(n1268) );
NAND3_X1 U924 ( .A1(n1276), .A2(n1277), .A3(n1278), .ZN(n1267) );
NAND2_X1 U925 ( .A1(KEYINPUT57), .A2(n1279), .ZN(n1278) );
INV_X1 U926 ( .A(n1280), .ZN(n1279) );
OR3_X1 U927 ( .A1(n1281), .A2(KEYINPUT57), .A3(n1282), .ZN(n1277) );
NAND2_X1 U928 ( .A1(n1281), .A2(n1282), .ZN(n1276) );
NAND2_X1 U929 ( .A1(KEYINPUT10), .A2(n1280), .ZN(n1281) );
XNOR2_X1 U930 ( .A(G110), .B(n1283), .ZN(n1280) );
INV_X1 U931 ( .A(n1263), .ZN(n1270) );
XNOR2_X1 U932 ( .A(n1284), .B(n1285), .ZN(n1263) );
NOR2_X1 U933 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
AND2_X1 U934 ( .A1(KEYINPUT44), .A2(n1288), .ZN(n1287) );
NOR2_X1 U935 ( .A1(KEYINPUT15), .A2(n1288), .ZN(n1286) );
XOR2_X1 U936 ( .A(n1289), .B(n1290), .Z(n1288) );
XOR2_X1 U937 ( .A(n1291), .B(n1292), .Z(n1289) );
XNOR2_X1 U938 ( .A(G134), .B(n1293), .ZN(n1284) );
NOR2_X1 U939 ( .A1(n1219), .A2(n1294), .ZN(G51) );
XOR2_X1 U940 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U941 ( .A(n1297), .B(n1298), .Z(n1295) );
NOR2_X1 U942 ( .A1(n1168), .A2(n1225), .ZN(n1298) );
NAND2_X1 U943 ( .A1(G902), .A2(n1299), .ZN(n1225) );
NAND2_X1 U944 ( .A1(n1211), .A2(n1117), .ZN(n1299) );
NOR3_X1 U945 ( .A1(n1300), .A2(n1193), .A3(n1192), .ZN(n1117) );
NAND3_X1 U946 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1192) );
NAND3_X1 U947 ( .A1(n1304), .A2(n1305), .A3(n1306), .ZN(n1303) );
XOR2_X1 U948 ( .A(KEYINPUT9), .B(n1122), .Z(n1305) );
INV_X1 U949 ( .A(n1307), .ZN(n1193) );
XOR2_X1 U950 ( .A(KEYINPUT41), .B(n1194), .Z(n1300) );
NAND4_X1 U951 ( .A1(n1308), .A2(n1309), .A3(n1310), .A4(n1311), .ZN(n1194) );
NAND2_X1 U952 ( .A1(n1154), .A2(n1312), .ZN(n1309) );
NAND2_X1 U953 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND4_X1 U954 ( .A1(n1315), .A2(n1136), .A3(n1141), .A4(n1316), .ZN(n1314) );
NOR2_X1 U955 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U956 ( .A1(n1306), .A2(n1152), .ZN(n1313) );
NAND2_X1 U957 ( .A1(n1319), .A2(n1318), .ZN(n1308) );
INV_X1 U958 ( .A(KEYINPUT3), .ZN(n1318) );
INV_X1 U959 ( .A(n1116), .ZN(n1211) );
NAND4_X1 U960 ( .A1(n1320), .A2(n1235), .A3(n1321), .A4(n1322), .ZN(n1116) );
AND4_X1 U961 ( .A1(n1110), .A2(n1323), .A3(n1324), .A4(n1325), .ZN(n1322) );
NAND3_X1 U962 ( .A1(n1155), .A2(n1130), .A3(n1326), .ZN(n1110) );
NAND2_X1 U963 ( .A1(n1122), .A2(n1327), .ZN(n1321) );
NAND2_X1 U964 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND3_X1 U965 ( .A1(n1330), .A2(n1331), .A3(n1152), .ZN(n1329) );
OR2_X1 U966 ( .A1(n1326), .A2(KEYINPUT5), .ZN(n1331) );
NAND2_X1 U967 ( .A1(KEYINPUT5), .A2(n1332), .ZN(n1330) );
NAND3_X1 U968 ( .A1(n1333), .A2(n1148), .A3(n1334), .ZN(n1332) );
NAND2_X1 U969 ( .A1(n1304), .A2(n1335), .ZN(n1328) );
NAND3_X1 U970 ( .A1(n1326), .A2(n1130), .A3(n1154), .ZN(n1235) );
NAND3_X1 U971 ( .A1(n1335), .A2(n1130), .A3(n1336), .ZN(n1320) );
NAND3_X1 U972 ( .A1(n1337), .A2(n1338), .A3(n1339), .ZN(n1297) );
NAND2_X1 U973 ( .A1(n1340), .A2(n1341), .ZN(n1338) );
INV_X1 U974 ( .A(KEYINPUT58), .ZN(n1341) );
NAND2_X1 U975 ( .A1(n1342), .A2(KEYINPUT58), .ZN(n1337) );
NOR2_X1 U976 ( .A1(n1121), .A2(G952), .ZN(n1219) );
XNOR2_X1 U977 ( .A(G146), .B(n1307), .ZN(G48) );
NAND3_X1 U978 ( .A1(n1304), .A2(n1154), .A3(n1343), .ZN(n1307) );
XNOR2_X1 U979 ( .A(G143), .B(n1301), .ZN(G45) );
NAND3_X1 U980 ( .A1(n1336), .A2(n1152), .A3(n1343), .ZN(n1301) );
XOR2_X1 U981 ( .A(n1302), .B(n1344), .Z(G42) );
NAND2_X1 U982 ( .A1(KEYINPUT62), .A2(G140), .ZN(n1344) );
NAND3_X1 U983 ( .A1(n1154), .A2(n1141), .A3(n1306), .ZN(n1302) );
XOR2_X1 U984 ( .A(G137), .B(n1345), .Z(G39) );
AND3_X1 U985 ( .A1(n1306), .A2(n1122), .A3(n1304), .ZN(n1345) );
XNOR2_X1 U986 ( .A(G134), .B(n1310), .ZN(G36) );
NAND3_X1 U987 ( .A1(n1152), .A2(n1155), .A3(n1306), .ZN(n1310) );
AND3_X1 U988 ( .A1(n1148), .A2(n1315), .A3(n1127), .ZN(n1306) );
NAND3_X1 U989 ( .A1(n1346), .A2(n1347), .A3(n1348), .ZN(G33) );
NAND2_X1 U990 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND3_X1 U991 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1350) );
NAND2_X1 U992 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NAND2_X1 U993 ( .A1(G131), .A2(n1356), .ZN(n1352) );
INV_X1 U994 ( .A(KEYINPUT33), .ZN(n1356) );
NAND2_X1 U995 ( .A1(KEYINPUT33), .A2(n1357), .ZN(n1351) );
NAND2_X1 U996 ( .A1(G131), .A2(n1358), .ZN(n1357) );
NAND2_X1 U997 ( .A1(KEYINPUT14), .A2(KEYINPUT52), .ZN(n1358) );
INV_X1 U998 ( .A(n1359), .ZN(n1349) );
NAND4_X1 U999 ( .A1(n1359), .A2(n1355), .A3(G131), .A4(KEYINPUT14), .ZN(n1347) );
INV_X1 U1000 ( .A(KEYINPUT52), .ZN(n1355) );
NAND2_X1 U1001 ( .A1(n1360), .A2(n1354), .ZN(n1346) );
INV_X1 U1002 ( .A(KEYINPUT14), .ZN(n1354) );
NAND2_X1 U1003 ( .A1(G131), .A2(n1361), .ZN(n1360) );
NAND2_X1 U1004 ( .A1(KEYINPUT52), .A2(n1359), .ZN(n1361) );
NAND4_X1 U1005 ( .A1(n1127), .A2(n1152), .A3(n1362), .A4(n1154), .ZN(n1359) );
NOR2_X1 U1006 ( .A1(n1363), .A2(n1364), .ZN(n1362) );
XNOR2_X1 U1007 ( .A(n1148), .B(KEYINPUT26), .ZN(n1364) );
AND2_X1 U1008 ( .A1(n1140), .A2(n1365), .ZN(n1127) );
XNOR2_X1 U1009 ( .A(G128), .B(n1311), .ZN(G30) );
NAND3_X1 U1010 ( .A1(n1304), .A2(n1155), .A3(n1343), .ZN(n1311) );
NOR3_X1 U1011 ( .A1(n1366), .A2(n1363), .A3(n1136), .ZN(n1343) );
INV_X1 U1012 ( .A(n1315), .ZN(n1363) );
XNOR2_X1 U1013 ( .A(G101), .B(n1367), .ZN(G3) );
NAND2_X1 U1014 ( .A1(n1152), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1015 ( .A(G125), .B(n1319), .Z(G27) );
AND4_X1 U1016 ( .A1(n1333), .A2(n1315), .A3(n1141), .A4(n1369), .ZN(n1319) );
NOR2_X1 U1017 ( .A1(n1317), .A2(n1370), .ZN(n1369) );
NAND2_X1 U1018 ( .A1(n1158), .A2(n1371), .ZN(n1315) );
NAND2_X1 U1019 ( .A1(n1198), .A2(n1372), .ZN(n1371) );
XNOR2_X1 U1020 ( .A(G900), .B(KEYINPUT22), .ZN(n1198) );
XNOR2_X1 U1021 ( .A(G122), .B(n1373), .ZN(G24) );
NAND3_X1 U1022 ( .A1(n1130), .A2(n1374), .A3(n1335), .ZN(n1373) );
XOR2_X1 U1023 ( .A(KEYINPUT55), .B(n1336), .Z(n1374) );
AND2_X1 U1024 ( .A1(n1375), .A2(n1376), .ZN(n1336) );
NOR2_X1 U1025 ( .A1(n1377), .A2(n1378), .ZN(n1130) );
XNOR2_X1 U1026 ( .A(G119), .B(n1379), .ZN(G21) );
NAND4_X1 U1027 ( .A1(n1304), .A2(n1122), .A3(n1380), .A4(n1381), .ZN(n1379) );
OR2_X1 U1028 ( .A1(n1382), .A2(n1335), .ZN(n1381) );
NAND2_X1 U1029 ( .A1(n1383), .A2(n1382), .ZN(n1380) );
INV_X1 U1030 ( .A(KEYINPUT31), .ZN(n1382) );
NAND3_X1 U1031 ( .A1(n1384), .A2(n1136), .A3(n1131), .ZN(n1383) );
INV_X1 U1032 ( .A(n1317), .ZN(n1131) );
NOR2_X1 U1033 ( .A1(n1385), .A2(n1386), .ZN(n1304) );
XNOR2_X1 U1034 ( .A(G116), .B(n1325), .ZN(G18) );
NAND3_X1 U1035 ( .A1(n1335), .A2(n1155), .A3(n1152), .ZN(n1325) );
NOR2_X1 U1036 ( .A1(n1376), .A2(n1387), .ZN(n1155) );
XNOR2_X1 U1037 ( .A(G113), .B(n1324), .ZN(G15) );
NAND3_X1 U1038 ( .A1(n1335), .A2(n1154), .A3(n1152), .ZN(n1324) );
NOR2_X1 U1039 ( .A1(n1377), .A2(n1385), .ZN(n1152) );
INV_X1 U1040 ( .A(n1378), .ZN(n1385) );
INV_X1 U1041 ( .A(n1386), .ZN(n1377) );
INV_X1 U1042 ( .A(n1370), .ZN(n1154) );
NAND2_X1 U1043 ( .A1(n1387), .A2(n1376), .ZN(n1370) );
NOR3_X1 U1044 ( .A1(n1136), .A2(n1334), .A3(n1317), .ZN(n1335) );
NAND2_X1 U1045 ( .A1(n1129), .A2(n1388), .ZN(n1317) );
XNOR2_X1 U1046 ( .A(G110), .B(n1323), .ZN(G12) );
NAND2_X1 U1047 ( .A1(n1368), .A2(n1141), .ZN(n1323) );
NOR2_X1 U1048 ( .A1(n1378), .A2(n1386), .ZN(n1141) );
NOR2_X1 U1049 ( .A1(n1179), .A2(n1389), .ZN(n1386) );
NOR2_X1 U1050 ( .A1(n1182), .A2(n1183), .ZN(n1389) );
AND2_X1 U1051 ( .A1(n1183), .A2(n1182), .ZN(n1179) );
NAND2_X1 U1052 ( .A1(G217), .A2(n1390), .ZN(n1182) );
NOR2_X1 U1053 ( .A1(n1226), .A2(G902), .ZN(n1183) );
XOR2_X1 U1054 ( .A(n1391), .B(n1392), .Z(n1226) );
XOR2_X1 U1055 ( .A(n1393), .B(n1394), .Z(n1392) );
XNOR2_X1 U1056 ( .A(G128), .B(n1395), .ZN(n1394) );
XOR2_X1 U1057 ( .A(KEYINPUT17), .B(G137), .Z(n1393) );
XOR2_X1 U1058 ( .A(n1396), .B(n1397), .Z(n1391) );
XOR2_X1 U1059 ( .A(n1398), .B(n1399), .Z(n1397) );
NAND2_X1 U1060 ( .A1(KEYINPUT48), .A2(n1400), .ZN(n1399) );
NAND2_X1 U1061 ( .A1(n1401), .A2(n1402), .ZN(n1398) );
NAND2_X1 U1062 ( .A1(G125), .A2(n1283), .ZN(n1402) );
XOR2_X1 U1063 ( .A(KEYINPUT35), .B(n1403), .Z(n1401) );
NOR2_X1 U1064 ( .A1(G125), .A2(n1283), .ZN(n1403) );
XNOR2_X1 U1065 ( .A(n1404), .B(n1405), .ZN(n1396) );
NAND2_X1 U1066 ( .A1(n1406), .A2(G221), .ZN(n1404) );
XNOR2_X1 U1067 ( .A(n1170), .B(G472), .ZN(n1378) );
NAND2_X1 U1068 ( .A1(n1407), .A2(n1408), .ZN(n1170) );
XOR2_X1 U1069 ( .A(n1409), .B(n1410), .Z(n1408) );
XNOR2_X1 U1070 ( .A(n1258), .B(n1411), .ZN(n1410) );
XNOR2_X1 U1071 ( .A(n1248), .B(n1243), .ZN(n1411) );
NAND2_X1 U1072 ( .A1(n1412), .A2(G210), .ZN(n1248) );
XOR2_X1 U1073 ( .A(G119), .B(n1413), .Z(n1258) );
NOR2_X1 U1074 ( .A1(G116), .A2(KEYINPUT19), .ZN(n1413) );
XNOR2_X1 U1075 ( .A(n1255), .B(n1414), .ZN(n1409) );
XNOR2_X1 U1076 ( .A(G902), .B(KEYINPUT34), .ZN(n1407) );
AND2_X1 U1077 ( .A1(n1122), .A2(n1326), .ZN(n1368) );
NOR3_X1 U1078 ( .A1(n1366), .A2(n1334), .A3(n1136), .ZN(n1326) );
INV_X1 U1079 ( .A(n1333), .ZN(n1136) );
NOR2_X1 U1080 ( .A1(n1140), .A2(n1138), .ZN(n1333) );
INV_X1 U1081 ( .A(n1365), .ZN(n1138) );
NAND2_X1 U1082 ( .A1(G214), .A2(n1415), .ZN(n1365) );
XOR2_X1 U1083 ( .A(n1416), .B(n1169), .Z(n1140) );
NAND2_X1 U1084 ( .A1(n1417), .A2(n1418), .ZN(n1169) );
XOR2_X1 U1085 ( .A(n1419), .B(n1296), .Z(n1417) );
XNOR2_X1 U1086 ( .A(n1218), .B(n1217), .ZN(n1296) );
XNOR2_X1 U1087 ( .A(n1420), .B(n1421), .ZN(n1217) );
XNOR2_X1 U1088 ( .A(n1243), .B(n1422), .ZN(n1421) );
NOR2_X1 U1089 ( .A1(KEYINPUT51), .A2(n1423), .ZN(n1422) );
XNOR2_X1 U1090 ( .A(G104), .B(n1424), .ZN(n1423) );
NAND2_X1 U1091 ( .A1(KEYINPUT18), .A2(n1425), .ZN(n1424) );
INV_X1 U1092 ( .A(G101), .ZN(n1243) );
XNOR2_X1 U1093 ( .A(G110), .B(n1426), .ZN(n1420) );
XNOR2_X1 U1094 ( .A(KEYINPUT37), .B(n1427), .ZN(n1426) );
NAND2_X1 U1095 ( .A1(n1428), .A2(n1429), .ZN(n1218) );
NAND2_X1 U1096 ( .A1(n1430), .A2(n1395), .ZN(n1429) );
INV_X1 U1097 ( .A(G119), .ZN(n1395) );
XOR2_X1 U1098 ( .A(n1431), .B(KEYINPUT43), .Z(n1430) );
NAND2_X1 U1099 ( .A1(G119), .A2(n1432), .ZN(n1428) );
XOR2_X1 U1100 ( .A(n1431), .B(KEYINPUT40), .Z(n1432) );
XNOR2_X1 U1101 ( .A(G113), .B(G116), .ZN(n1431) );
NOR2_X1 U1102 ( .A1(n1342), .A2(n1433), .ZN(n1419) );
INV_X1 U1103 ( .A(n1339), .ZN(n1433) );
NAND2_X1 U1104 ( .A1(n1340), .A2(n1434), .ZN(n1339) );
NOR2_X1 U1105 ( .A1(n1434), .A2(n1340), .ZN(n1342) );
XNOR2_X1 U1106 ( .A(n1435), .B(n1290), .ZN(n1340) );
XNOR2_X1 U1107 ( .A(G128), .B(n1400), .ZN(n1290) );
XNOR2_X1 U1108 ( .A(G125), .B(G143), .ZN(n1435) );
NAND2_X1 U1109 ( .A1(G224), .A2(n1121), .ZN(n1434) );
NAND2_X1 U1110 ( .A1(KEYINPUT36), .A2(n1168), .ZN(n1416) );
NAND2_X1 U1111 ( .A1(G210), .A2(n1415), .ZN(n1168) );
NAND2_X1 U1112 ( .A1(n1436), .A2(n1418), .ZN(n1415) );
INV_X1 U1113 ( .A(G237), .ZN(n1436) );
INV_X1 U1114 ( .A(n1384), .ZN(n1334) );
NAND2_X1 U1115 ( .A1(n1437), .A2(n1158), .ZN(n1384) );
NAND3_X1 U1116 ( .A1(n1438), .A2(n1121), .A3(G952), .ZN(n1158) );
NAND2_X1 U1117 ( .A1(n1372), .A2(n1215), .ZN(n1437) );
INV_X1 U1118 ( .A(G898), .ZN(n1215) );
AND3_X1 U1119 ( .A1(G902), .A2(n1438), .A3(G953), .ZN(n1372) );
NAND2_X1 U1120 ( .A1(G237), .A2(G234), .ZN(n1438) );
INV_X1 U1121 ( .A(n1148), .ZN(n1366) );
NOR2_X1 U1122 ( .A1(n1129), .A2(n1128), .ZN(n1148) );
INV_X1 U1123 ( .A(n1388), .ZN(n1128) );
NAND2_X1 U1124 ( .A1(G221), .A2(n1390), .ZN(n1388) );
NAND2_X1 U1125 ( .A1(G234), .A2(n1418), .ZN(n1390) );
XNOR2_X1 U1126 ( .A(n1185), .B(n1439), .ZN(n1129) );
XOR2_X1 U1127 ( .A(KEYINPUT8), .B(G469), .Z(n1439) );
AND2_X1 U1128 ( .A1(n1440), .A2(n1418), .ZN(n1185) );
INV_X1 U1129 ( .A(G902), .ZN(n1418) );
XOR2_X1 U1130 ( .A(n1441), .B(n1442), .Z(n1440) );
XNOR2_X1 U1131 ( .A(n1283), .B(n1443), .ZN(n1442) );
NOR2_X1 U1132 ( .A1(KEYINPUT54), .A2(n1444), .ZN(n1443) );
XOR2_X1 U1133 ( .A(n1201), .B(n1291), .Z(n1444) );
XNOR2_X1 U1134 ( .A(G101), .B(n1445), .ZN(n1291) );
XNOR2_X1 U1135 ( .A(n1425), .B(G104), .ZN(n1445) );
XNOR2_X1 U1136 ( .A(n1255), .B(n1292), .ZN(n1201) );
AND2_X1 U1137 ( .A1(KEYINPUT46), .A2(n1446), .ZN(n1292) );
XOR2_X1 U1138 ( .A(KEYINPUT45), .B(G143), .Z(n1446) );
XNOR2_X1 U1139 ( .A(n1447), .B(n1448), .ZN(n1255) );
XNOR2_X1 U1140 ( .A(G146), .B(n1293), .ZN(n1447) );
XOR2_X1 U1141 ( .A(G137), .B(G131), .Z(n1293) );
INV_X1 U1142 ( .A(G140), .ZN(n1283) );
XNOR2_X1 U1143 ( .A(n1449), .B(n1282), .ZN(n1441) );
NAND2_X1 U1144 ( .A1(G227), .A2(n1121), .ZN(n1282) );
NAND2_X1 U1145 ( .A1(KEYINPUT30), .A2(n1405), .ZN(n1449) );
INV_X1 U1146 ( .A(G110), .ZN(n1405) );
NOR2_X1 U1147 ( .A1(n1375), .A2(n1376), .ZN(n1122) );
XNOR2_X1 U1148 ( .A(n1177), .B(n1234), .ZN(n1376) );
INV_X1 U1149 ( .A(G475), .ZN(n1234) );
NOR2_X1 U1150 ( .A1(n1232), .A2(G902), .ZN(n1177) );
XOR2_X1 U1151 ( .A(n1450), .B(n1451), .Z(n1232) );
XOR2_X1 U1152 ( .A(n1452), .B(n1453), .Z(n1451) );
XOR2_X1 U1153 ( .A(n1454), .B(n1414), .Z(n1453) );
XOR2_X1 U1154 ( .A(G113), .B(G143), .Z(n1414) );
NAND2_X1 U1155 ( .A1(n1412), .A2(G214), .ZN(n1454) );
NOR2_X1 U1156 ( .A1(G953), .A2(G237), .ZN(n1412) );
NAND2_X1 U1157 ( .A1(n1455), .A2(n1456), .ZN(n1452) );
NAND2_X1 U1158 ( .A1(n1457), .A2(n1400), .ZN(n1456) );
INV_X1 U1159 ( .A(G146), .ZN(n1400) );
XNOR2_X1 U1160 ( .A(n1458), .B(KEYINPUT28), .ZN(n1457) );
NAND2_X1 U1161 ( .A1(n1459), .A2(G146), .ZN(n1455) );
XNOR2_X1 U1162 ( .A(KEYINPUT2), .B(n1460), .ZN(n1459) );
INV_X1 U1163 ( .A(n1458), .ZN(n1460) );
XOR2_X1 U1164 ( .A(G125), .B(n1461), .Z(n1458) );
NOR2_X1 U1165 ( .A1(G140), .A2(KEYINPUT50), .ZN(n1461) );
XOR2_X1 U1166 ( .A(n1462), .B(n1463), .Z(n1450) );
XOR2_X1 U1167 ( .A(G131), .B(G104), .Z(n1463) );
NAND2_X1 U1168 ( .A1(KEYINPUT7), .A2(n1427), .ZN(n1462) );
INV_X1 U1169 ( .A(n1387), .ZN(n1375) );
XOR2_X1 U1170 ( .A(n1175), .B(n1230), .Z(n1387) );
INV_X1 U1171 ( .A(G478), .ZN(n1230) );
NOR2_X1 U1172 ( .A1(n1228), .A2(G902), .ZN(n1175) );
XOR2_X1 U1173 ( .A(n1464), .B(n1465), .Z(n1228) );
XOR2_X1 U1174 ( .A(G116), .B(n1466), .Z(n1465) );
XNOR2_X1 U1175 ( .A(G143), .B(n1427), .ZN(n1466) );
INV_X1 U1176 ( .A(G122), .ZN(n1427) );
XOR2_X1 U1177 ( .A(n1467), .B(n1448), .Z(n1464) );
XOR2_X1 U1178 ( .A(G134), .B(G128), .Z(n1448) );
XNOR2_X1 U1179 ( .A(n1468), .B(n1425), .ZN(n1467) );
INV_X1 U1180 ( .A(G107), .ZN(n1425) );
NAND2_X1 U1181 ( .A1(G217), .A2(n1406), .ZN(n1468) );
AND2_X1 U1182 ( .A1(G234), .A2(n1121), .ZN(n1406) );
INV_X1 U1183 ( .A(G953), .ZN(n1121) );
endmodule


