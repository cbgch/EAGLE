//Key = 1101111100101010101111000100011101010101010011111101111100110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413;

XOR2_X1 U771 ( .A(n1082), .B(n1083), .Z(G9) );
NOR4_X1 U772 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1083) );
INV_X1 U773 ( .A(n1088), .ZN(n1085) );
XOR2_X1 U774 ( .A(n1089), .B(KEYINPUT17), .Z(n1084) );
NAND2_X1 U775 ( .A1(KEYINPUT51), .A2(n1090), .ZN(n1082) );
NOR2_X1 U776 ( .A1(n1091), .A2(n1092), .ZN(G75) );
XOR2_X1 U777 ( .A(n1093), .B(KEYINPUT29), .Z(n1092) );
NAND3_X1 U778 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1093) );
NOR2_X1 U779 ( .A1(n1097), .A2(n1098), .ZN(n1091) );
NAND4_X1 U780 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(G952), .ZN(n1098) );
XOR2_X1 U781 ( .A(n1102), .B(KEYINPUT59), .Z(n1099) );
NAND2_X1 U782 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U783 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND3_X1 U784 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1103) );
NAND2_X1 U785 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NAND2_X1 U786 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U787 ( .A1(n1114), .A2(n1115), .ZN(n1110) );
OR2_X1 U788 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND4_X1 U789 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1096), .ZN(n1097) );
NAND4_X1 U790 ( .A1(n1114), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1096) );
NOR4_X1 U791 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1123) );
XOR2_X1 U792 ( .A(n1128), .B(G472), .Z(n1126) );
NAND2_X1 U793 ( .A1(KEYINPUT20), .A2(n1129), .ZN(n1128) );
INV_X1 U794 ( .A(n1130), .ZN(n1125) );
INV_X1 U795 ( .A(n1131), .ZN(n1124) );
NOR4_X1 U796 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1122) );
NOR3_X1 U797 ( .A1(n1136), .A2(KEYINPUT50), .A3(n1137), .ZN(n1135) );
AND2_X1 U798 ( .A1(n1136), .A2(KEYINPUT50), .ZN(n1134) );
NOR3_X1 U799 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1133) );
INV_X1 U800 ( .A(KEYINPUT39), .ZN(n1138) );
NOR2_X1 U801 ( .A1(KEYINPUT39), .A2(G475), .ZN(n1132) );
NAND3_X1 U802 ( .A1(n1107), .A2(n1141), .A3(n1109), .ZN(n1120) );
NAND2_X1 U803 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND3_X1 U804 ( .A1(n1144), .A2(n1145), .A3(n1112), .ZN(n1143) );
NAND2_X1 U805 ( .A1(n1114), .A2(n1146), .ZN(n1142) );
NAND2_X1 U806 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
NAND3_X1 U807 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
NAND2_X1 U808 ( .A1(n1121), .A2(n1152), .ZN(n1147) );
NAND2_X1 U809 ( .A1(n1105), .A2(n1088), .ZN(n1119) );
AND3_X1 U810 ( .A1(n1112), .A2(n1114), .A3(n1109), .ZN(n1105) );
INV_X1 U811 ( .A(n1153), .ZN(n1109) );
NOR2_X1 U812 ( .A1(n1154), .A2(n1086), .ZN(n1112) );
XOR2_X1 U813 ( .A(KEYINPUT49), .B(G953), .Z(n1118) );
XOR2_X1 U814 ( .A(n1155), .B(n1156), .Z(G72) );
XOR2_X1 U815 ( .A(n1157), .B(n1158), .Z(n1156) );
NOR2_X1 U816 ( .A1(n1101), .A2(n1159), .ZN(n1158) );
XOR2_X1 U817 ( .A(KEYINPUT26), .B(G953), .Z(n1159) );
NAND3_X1 U818 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1157) );
XOR2_X1 U819 ( .A(n1163), .B(KEYINPUT43), .Z(n1162) );
OR2_X1 U820 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U821 ( .A1(n1164), .A2(n1165), .ZN(n1161) );
XNOR2_X1 U822 ( .A(n1166), .B(n1167), .ZN(n1164) );
XOR2_X1 U823 ( .A(n1168), .B(G131), .Z(n1166) );
NAND2_X1 U824 ( .A1(G953), .A2(n1169), .ZN(n1160) );
NAND2_X1 U825 ( .A1(G953), .A2(n1170), .ZN(n1155) );
NAND2_X1 U826 ( .A1(G900), .A2(G227), .ZN(n1170) );
XOR2_X1 U827 ( .A(n1171), .B(n1172), .Z(G69) );
XOR2_X1 U828 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U829 ( .A1(n1175), .A2(n1095), .ZN(n1174) );
NOR2_X1 U830 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND2_X1 U831 ( .A1(n1178), .A2(n1179), .ZN(n1173) );
NAND2_X1 U832 ( .A1(G953), .A2(n1177), .ZN(n1179) );
XOR2_X1 U833 ( .A(n1180), .B(n1181), .Z(n1178) );
XOR2_X1 U834 ( .A(n1182), .B(n1183), .Z(n1181) );
XNOR2_X1 U835 ( .A(KEYINPUT13), .B(n1184), .ZN(n1180) );
NOR2_X1 U836 ( .A1(KEYINPUT24), .A2(n1185), .ZN(n1184) );
NAND2_X1 U837 ( .A1(n1095), .A2(n1186), .ZN(n1171) );
NOR3_X1 U838 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(G66) );
AND3_X1 U839 ( .A1(KEYINPUT36), .A2(n1095), .A3(n1094), .ZN(n1189) );
NOR2_X1 U840 ( .A1(KEYINPUT36), .A2(n1190), .ZN(n1188) );
XOR2_X1 U841 ( .A(n1191), .B(n1192), .Z(n1187) );
NOR2_X1 U842 ( .A1(n1136), .A2(n1193), .ZN(n1192) );
NAND2_X1 U843 ( .A1(KEYINPUT55), .A2(n1194), .ZN(n1191) );
NOR2_X1 U844 ( .A1(n1195), .A2(n1196), .ZN(G63) );
XOR2_X1 U845 ( .A(n1197), .B(n1198), .Z(n1196) );
AND2_X1 U846 ( .A1(G478), .A2(n1199), .ZN(n1197) );
NOR2_X1 U847 ( .A1(n1195), .A2(n1200), .ZN(G60) );
XOR2_X1 U848 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U849 ( .A(KEYINPUT62), .B(n1203), .Z(n1202) );
NOR2_X1 U850 ( .A1(n1140), .A2(n1193), .ZN(n1203) );
XOR2_X1 U851 ( .A(G104), .B(n1204), .Z(G6) );
NOR2_X1 U852 ( .A1(n1205), .A2(n1206), .ZN(G57) );
XOR2_X1 U853 ( .A(n1207), .B(n1208), .Z(n1206) );
XOR2_X1 U854 ( .A(n1209), .B(G101), .Z(n1208) );
NAND2_X1 U855 ( .A1(n1210), .A2(KEYINPUT45), .ZN(n1209) );
XOR2_X1 U856 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U857 ( .A(n1213), .B(n1214), .Z(n1212) );
AND2_X1 U858 ( .A1(G472), .A2(n1199), .ZN(n1214) );
NAND2_X1 U859 ( .A1(KEYINPUT7), .A2(n1215), .ZN(n1213) );
NAND2_X1 U860 ( .A1(KEYINPUT6), .A2(n1216), .ZN(n1207) );
XOR2_X1 U861 ( .A(n1190), .B(KEYINPUT4), .Z(n1205) );
NOR3_X1 U862 ( .A1(n1195), .A2(n1217), .A3(n1218), .ZN(G54) );
NOR2_X1 U863 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NOR2_X1 U864 ( .A1(n1221), .A2(n1222), .ZN(n1219) );
NOR2_X1 U865 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
NOR2_X1 U866 ( .A1(n1225), .A2(n1226), .ZN(n1221) );
NOR2_X1 U867 ( .A1(n1227), .A2(n1228), .ZN(n1217) );
NOR2_X1 U868 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
NOR2_X1 U869 ( .A1(n1224), .A2(n1226), .ZN(n1230) );
XOR2_X1 U870 ( .A(n1231), .B(KEYINPUT48), .Z(n1226) );
NOR2_X1 U871 ( .A1(n1225), .A2(n1223), .ZN(n1229) );
XOR2_X1 U872 ( .A(n1231), .B(KEYINPUT32), .Z(n1223) );
NAND2_X1 U873 ( .A1(n1199), .A2(G469), .ZN(n1231) );
INV_X1 U874 ( .A(n1193), .ZN(n1199) );
INV_X1 U875 ( .A(n1224), .ZN(n1225) );
XOR2_X1 U876 ( .A(n1232), .B(n1233), .Z(n1224) );
XOR2_X1 U877 ( .A(KEYINPUT54), .B(n1234), .Z(n1233) );
NAND2_X1 U878 ( .A1(n1235), .A2(n1236), .ZN(n1232) );
NAND2_X1 U879 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XOR2_X1 U880 ( .A(n1239), .B(KEYINPUT42), .Z(n1235) );
OR2_X1 U881 ( .A1(n1237), .A2(n1238), .ZN(n1239) );
INV_X1 U882 ( .A(n1220), .ZN(n1227) );
XOR2_X1 U883 ( .A(n1240), .B(n1241), .Z(n1220) );
NOR2_X1 U884 ( .A1(KEYINPUT34), .A2(n1242), .ZN(n1241) );
NOR2_X1 U885 ( .A1(n1195), .A2(n1243), .ZN(G51) );
XOR2_X1 U886 ( .A(n1244), .B(n1245), .Z(n1243) );
XOR2_X1 U887 ( .A(KEYINPUT11), .B(n1246), .Z(n1245) );
NOR2_X1 U888 ( .A1(n1247), .A2(n1193), .ZN(n1246) );
NAND2_X1 U889 ( .A1(G902), .A2(n1248), .ZN(n1193) );
NAND2_X1 U890 ( .A1(n1100), .A2(n1101), .ZN(n1248) );
AND4_X1 U891 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1101) );
AND4_X1 U892 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1252) );
NAND3_X1 U893 ( .A1(n1257), .A2(n1113), .A3(n1088), .ZN(n1256) );
AND2_X1 U894 ( .A1(n1258), .A2(n1259), .ZN(n1251) );
NAND2_X1 U895 ( .A1(n1260), .A2(n1261), .ZN(n1249) );
XNOR2_X1 U896 ( .A(n1152), .B(KEYINPUT44), .ZN(n1260) );
INV_X1 U897 ( .A(n1186), .ZN(n1100) );
NAND4_X1 U898 ( .A1(n1262), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(n1186) );
AND4_X1 U899 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1269), .ZN(n1265) );
NOR2_X1 U900 ( .A1(n1270), .A2(n1204), .ZN(n1264) );
AND3_X1 U901 ( .A1(n1106), .A2(n1271), .A3(n1116), .ZN(n1204) );
NOR2_X1 U902 ( .A1(n1154), .A2(n1272), .ZN(n1270) );
NAND4_X1 U903 ( .A1(n1116), .A2(n1088), .A3(n1273), .A4(n1274), .ZN(n1262) );
NAND2_X1 U904 ( .A1(KEYINPUT19), .A2(n1087), .ZN(n1274) );
NAND2_X1 U905 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
INV_X1 U906 ( .A(KEYINPUT19), .ZN(n1276) );
NAND2_X1 U907 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
NOR2_X1 U908 ( .A1(n1086), .A2(n1089), .ZN(n1116) );
INV_X1 U909 ( .A(n1190), .ZN(n1195) );
NAND2_X1 U910 ( .A1(G953), .A2(n1094), .ZN(n1190) );
INV_X1 U911 ( .A(G952), .ZN(n1094) );
XNOR2_X1 U912 ( .A(G146), .B(n1255), .ZN(G48) );
NAND3_X1 U913 ( .A1(n1106), .A2(n1113), .A3(n1257), .ZN(n1255) );
XOR2_X1 U914 ( .A(n1279), .B(n1250), .Z(G45) );
NAND4_X1 U915 ( .A1(n1280), .A2(n1281), .A3(n1113), .A4(n1282), .ZN(n1250) );
XNOR2_X1 U916 ( .A(G140), .B(n1259), .ZN(G42) );
NAND4_X1 U917 ( .A1(n1114), .A2(n1106), .A3(n1283), .A4(n1152), .ZN(n1259) );
NOR2_X1 U918 ( .A1(n1284), .A2(n1089), .ZN(n1283) );
XNOR2_X1 U919 ( .A(G137), .B(n1254), .ZN(G39) );
NAND3_X1 U920 ( .A1(n1114), .A2(n1107), .A3(n1257), .ZN(n1254) );
XNOR2_X1 U921 ( .A(G134), .B(n1253), .ZN(G36) );
NAND3_X1 U922 ( .A1(n1114), .A2(n1088), .A3(n1281), .ZN(n1253) );
XOR2_X1 U923 ( .A(n1285), .B(n1258), .Z(G33) );
NAND3_X1 U924 ( .A1(n1114), .A2(n1106), .A3(n1281), .ZN(n1258) );
AND2_X1 U925 ( .A1(n1286), .A2(n1287), .ZN(n1281) );
NOR2_X1 U926 ( .A1(n1288), .A2(n1145), .ZN(n1114) );
INV_X1 U927 ( .A(n1144), .ZN(n1288) );
XOR2_X1 U928 ( .A(G128), .B(n1289), .Z(G30) );
NOR2_X1 U929 ( .A1(n1290), .A2(n1277), .ZN(n1289) );
INV_X1 U930 ( .A(n1113), .ZN(n1277) );
XOR2_X1 U931 ( .A(n1291), .B(KEYINPUT2), .Z(n1290) );
NAND2_X1 U932 ( .A1(n1257), .A2(n1088), .ZN(n1291) );
AND2_X1 U933 ( .A1(n1286), .A2(n1292), .ZN(n1257) );
NOR3_X1 U934 ( .A1(n1293), .A2(n1284), .A3(n1089), .ZN(n1286) );
INV_X1 U935 ( .A(n1294), .ZN(n1089) );
INV_X1 U936 ( .A(n1295), .ZN(n1284) );
NAND2_X1 U937 ( .A1(n1296), .A2(n1297), .ZN(G3) );
OR2_X1 U938 ( .A1(n1263), .A2(G101), .ZN(n1297) );
XOR2_X1 U939 ( .A(n1298), .B(KEYINPUT61), .Z(n1296) );
NAND2_X1 U940 ( .A1(G101), .A2(n1263), .ZN(n1298) );
NAND3_X1 U941 ( .A1(n1287), .A2(n1299), .A3(n1300), .ZN(n1263) );
XOR2_X1 U942 ( .A(n1301), .B(n1302), .Z(G27) );
AND2_X1 U943 ( .A1(n1152), .A2(n1261), .ZN(n1302) );
AND4_X1 U944 ( .A1(n1106), .A2(n1121), .A3(n1113), .A4(n1295), .ZN(n1261) );
NAND2_X1 U945 ( .A1(n1153), .A2(n1303), .ZN(n1295) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1304), .A4(n1169), .ZN(n1303) );
INV_X1 U947 ( .A(G900), .ZN(n1169) );
XOR2_X1 U948 ( .A(n1305), .B(KEYINPUT46), .Z(n1301) );
XOR2_X1 U949 ( .A(G122), .B(n1306), .Z(G24) );
NOR2_X1 U950 ( .A1(n1272), .A2(n1307), .ZN(n1306) );
XOR2_X1 U951 ( .A(KEYINPUT18), .B(n1121), .Z(n1307) );
NAND4_X1 U952 ( .A1(n1271), .A2(n1150), .A3(n1280), .A4(n1282), .ZN(n1272) );
INV_X1 U953 ( .A(n1086), .ZN(n1150) );
NAND2_X1 U954 ( .A1(n1287), .A2(n1293), .ZN(n1086) );
NAND3_X1 U955 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(G21) );
OR2_X1 U956 ( .A1(G119), .A2(KEYINPUT37), .ZN(n1310) );
NAND3_X1 U957 ( .A1(KEYINPUT37), .A2(G119), .A3(n1269), .ZN(n1309) );
NAND2_X1 U958 ( .A1(n1311), .A2(n1312), .ZN(n1308) );
NAND2_X1 U959 ( .A1(n1313), .A2(KEYINPUT37), .ZN(n1312) );
XOR2_X1 U960 ( .A(n1314), .B(KEYINPUT33), .Z(n1313) );
INV_X1 U961 ( .A(n1269), .ZN(n1311) );
NAND4_X1 U962 ( .A1(n1121), .A2(n1107), .A3(n1315), .A4(n1271), .ZN(n1269) );
NOR2_X1 U963 ( .A1(n1287), .A2(n1293), .ZN(n1315) );
INV_X1 U964 ( .A(n1154), .ZN(n1121) );
XOR2_X1 U965 ( .A(n1316), .B(n1268), .Z(G18) );
NAND3_X1 U966 ( .A1(n1271), .A2(n1088), .A3(n1117), .ZN(n1268) );
NOR2_X1 U967 ( .A1(n1282), .A2(n1317), .ZN(n1088) );
XOR2_X1 U968 ( .A(G113), .B(n1318), .Z(G15) );
NOR2_X1 U969 ( .A1(KEYINPUT23), .A2(n1267), .ZN(n1318) );
NAND3_X1 U970 ( .A1(n1106), .A2(n1271), .A3(n1117), .ZN(n1267) );
NOR3_X1 U971 ( .A1(n1292), .A2(n1293), .A3(n1154), .ZN(n1117) );
NAND2_X1 U972 ( .A1(n1149), .A2(n1319), .ZN(n1154) );
AND2_X1 U973 ( .A1(n1317), .A2(n1282), .ZN(n1106) );
INV_X1 U974 ( .A(n1280), .ZN(n1317) );
XOR2_X1 U975 ( .A(n1320), .B(n1266), .Z(G12) );
NAND2_X1 U976 ( .A1(n1152), .A2(n1300), .ZN(n1266) );
AND3_X1 U977 ( .A1(n1271), .A2(n1294), .A3(n1107), .ZN(n1300) );
NOR2_X1 U978 ( .A1(n1282), .A2(n1280), .ZN(n1107) );
XNOR2_X1 U979 ( .A(n1127), .B(KEYINPUT10), .ZN(n1280) );
XNOR2_X1 U980 ( .A(n1321), .B(G478), .ZN(n1127) );
OR2_X1 U981 ( .A1(n1198), .A2(G902), .ZN(n1321) );
XNOR2_X1 U982 ( .A(n1322), .B(n1323), .ZN(n1198) );
XOR2_X1 U983 ( .A(n1324), .B(n1325), .Z(n1323) );
XOR2_X1 U984 ( .A(n1090), .B(n1326), .Z(n1325) );
NOR2_X1 U985 ( .A1(G128), .A2(KEYINPUT56), .ZN(n1326) );
NAND3_X1 U986 ( .A1(G234), .A2(n1095), .A3(G217), .ZN(n1324) );
XOR2_X1 U987 ( .A(n1327), .B(n1328), .Z(n1322) );
XOR2_X1 U988 ( .A(G143), .B(G134), .Z(n1328) );
XOR2_X1 U989 ( .A(n1316), .B(G122), .Z(n1327) );
NAND2_X1 U990 ( .A1(n1329), .A2(n1131), .ZN(n1282) );
NAND2_X1 U991 ( .A1(n1139), .A2(n1140), .ZN(n1131) );
OR2_X1 U992 ( .A1(n1140), .A2(n1139), .ZN(n1329) );
NOR2_X1 U993 ( .A1(n1201), .A2(G902), .ZN(n1139) );
XOR2_X1 U994 ( .A(n1330), .B(n1331), .Z(n1201) );
XOR2_X1 U995 ( .A(n1332), .B(n1333), .Z(n1331) );
XOR2_X1 U996 ( .A(G113), .B(G104), .Z(n1333) );
XOR2_X1 U997 ( .A(G131), .B(G122), .Z(n1332) );
XNOR2_X1 U998 ( .A(n1165), .B(n1334), .ZN(n1330) );
XNOR2_X1 U999 ( .A(n1335), .B(n1336), .ZN(n1334) );
NOR2_X1 U1000 ( .A1(KEYINPUT22), .A2(n1337), .ZN(n1336) );
XOR2_X1 U1001 ( .A(n1279), .B(n1338), .Z(n1337) );
AND3_X1 U1002 ( .A1(G214), .A2(n1095), .A3(n1339), .ZN(n1338) );
INV_X1 U1003 ( .A(G143), .ZN(n1279) );
NAND2_X1 U1004 ( .A1(KEYINPUT3), .A2(G146), .ZN(n1335) );
XOR2_X1 U1005 ( .A(G125), .B(G140), .Z(n1165) );
INV_X1 U1006 ( .A(G475), .ZN(n1140) );
NOR2_X1 U1007 ( .A1(n1149), .A2(n1151), .ZN(n1294) );
INV_X1 U1008 ( .A(n1319), .ZN(n1151) );
NAND2_X1 U1009 ( .A1(G221), .A2(n1340), .ZN(n1319) );
XOR2_X1 U1010 ( .A(n1341), .B(G469), .Z(n1149) );
NAND2_X1 U1011 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1012 ( .A(n1344), .B(n1345), .Z(n1342) );
XNOR2_X1 U1013 ( .A(n1242), .B(n1237), .ZN(n1345) );
XOR2_X1 U1014 ( .A(G101), .B(n1346), .Z(n1237) );
XOR2_X1 U1015 ( .A(n1347), .B(n1238), .Z(n1344) );
INV_X1 U1016 ( .A(n1168), .ZN(n1238) );
XOR2_X1 U1017 ( .A(n1348), .B(n1349), .Z(n1168) );
XOR2_X1 U1018 ( .A(G143), .B(G128), .Z(n1349) );
NAND2_X1 U1019 ( .A1(KEYINPUT25), .A2(G146), .ZN(n1348) );
XOR2_X1 U1020 ( .A(n1350), .B(KEYINPUT58), .Z(n1347) );
NAND3_X1 U1021 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1350) );
NAND2_X1 U1022 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
INV_X1 U1023 ( .A(KEYINPUT53), .ZN(n1355) );
NAND3_X1 U1024 ( .A1(KEYINPUT53), .A2(n1234), .A3(n1356), .ZN(n1352) );
OR2_X1 U1025 ( .A1(n1356), .A2(n1234), .ZN(n1351) );
AND2_X1 U1026 ( .A1(G227), .A2(n1095), .ZN(n1234) );
NOR2_X1 U1027 ( .A1(KEYINPUT38), .A2(n1354), .ZN(n1356) );
XOR2_X1 U1028 ( .A(n1240), .B(KEYINPUT27), .Z(n1354) );
XOR2_X1 U1029 ( .A(n1320), .B(G140), .Z(n1240) );
INV_X1 U1030 ( .A(n1087), .ZN(n1271) );
NAND2_X1 U1031 ( .A1(n1113), .A2(n1278), .ZN(n1087) );
NAND2_X1 U1032 ( .A1(n1153), .A2(n1357), .ZN(n1278) );
NAND4_X1 U1033 ( .A1(G953), .A2(G902), .A3(n1304), .A4(n1177), .ZN(n1357) );
INV_X1 U1034 ( .A(G898), .ZN(n1177) );
NAND3_X1 U1035 ( .A1(n1304), .A2(n1095), .A3(G952), .ZN(n1153) );
NAND2_X1 U1036 ( .A1(n1358), .A2(G234), .ZN(n1304) );
XOR2_X1 U1037 ( .A(n1339), .B(KEYINPUT21), .Z(n1358) );
NOR2_X1 U1038 ( .A1(n1144), .A2(n1145), .ZN(n1113) );
AND2_X1 U1039 ( .A1(G214), .A2(n1359), .ZN(n1145) );
XNOR2_X1 U1040 ( .A(n1360), .B(n1247), .ZN(n1144) );
NAND2_X1 U1041 ( .A1(G210), .A2(n1359), .ZN(n1247) );
NAND2_X1 U1042 ( .A1(n1339), .A2(n1343), .ZN(n1359) );
OR2_X1 U1043 ( .A1(n1244), .A2(G902), .ZN(n1360) );
XNOR2_X1 U1044 ( .A(n1361), .B(n1362), .ZN(n1244) );
XOR2_X1 U1045 ( .A(n1363), .B(n1364), .Z(n1362) );
XOR2_X1 U1046 ( .A(n1365), .B(n1366), .Z(n1364) );
NOR2_X1 U1047 ( .A1(G953), .A2(n1176), .ZN(n1366) );
INV_X1 U1048 ( .A(G224), .ZN(n1176) );
NAND2_X1 U1049 ( .A1(KEYINPUT30), .A2(n1183), .ZN(n1365) );
XOR2_X1 U1050 ( .A(n1320), .B(G122), .Z(n1183) );
XOR2_X1 U1051 ( .A(n1305), .B(KEYINPUT40), .Z(n1363) );
XOR2_X1 U1052 ( .A(n1367), .B(n1185), .Z(n1361) );
XNOR2_X1 U1053 ( .A(n1368), .B(n1346), .ZN(n1185) );
XNOR2_X1 U1054 ( .A(G104), .B(n1090), .ZN(n1346) );
INV_X1 U1055 ( .A(G107), .ZN(n1090) );
NAND2_X1 U1056 ( .A1(KEYINPUT47), .A2(n1369), .ZN(n1368) );
XOR2_X1 U1057 ( .A(KEYINPUT9), .B(G101), .Z(n1369) );
XOR2_X1 U1058 ( .A(n1370), .B(n1182), .Z(n1367) );
XNOR2_X1 U1059 ( .A(n1314), .B(n1371), .ZN(n1182) );
NOR2_X1 U1060 ( .A1(n1299), .A2(n1287), .ZN(n1152) );
INV_X1 U1061 ( .A(n1292), .ZN(n1287) );
NAND3_X1 U1062 ( .A1(n1372), .A2(n1373), .A3(n1130), .ZN(n1292) );
NAND2_X1 U1063 ( .A1(n1137), .A2(n1136), .ZN(n1130) );
INV_X1 U1064 ( .A(n1374), .ZN(n1137) );
OR2_X1 U1065 ( .A1(n1375), .A2(KEYINPUT35), .ZN(n1373) );
NAND3_X1 U1066 ( .A1(n1375), .A2(n1374), .A3(KEYINPUT35), .ZN(n1372) );
NAND2_X1 U1067 ( .A1(n1194), .A2(n1343), .ZN(n1374) );
XNOR2_X1 U1068 ( .A(n1376), .B(n1377), .ZN(n1194) );
XOR2_X1 U1069 ( .A(n1378), .B(n1379), .Z(n1377) );
NOR2_X1 U1070 ( .A1(KEYINPUT57), .A2(n1380), .ZN(n1379) );
XOR2_X1 U1071 ( .A(n1381), .B(n1382), .Z(n1380) );
NOR2_X1 U1072 ( .A1(KEYINPUT60), .A2(n1383), .ZN(n1382) );
AND3_X1 U1073 ( .A1(G221), .A2(n1095), .A3(G234), .ZN(n1381) );
NOR2_X1 U1074 ( .A1(n1384), .A2(n1385), .ZN(n1378) );
XOR2_X1 U1075 ( .A(KEYINPUT15), .B(n1386), .Z(n1385) );
NOR2_X1 U1076 ( .A1(n1320), .A2(n1387), .ZN(n1386) );
NOR2_X1 U1077 ( .A1(G110), .A2(n1388), .ZN(n1384) );
XOR2_X1 U1078 ( .A(KEYINPUT12), .B(n1387), .Z(n1388) );
XOR2_X1 U1079 ( .A(n1389), .B(n1314), .Z(n1387) );
NAND2_X1 U1080 ( .A1(KEYINPUT14), .A2(n1390), .ZN(n1389) );
XOR2_X1 U1081 ( .A(KEYINPUT52), .B(G128), .Z(n1390) );
NAND2_X1 U1082 ( .A1(n1391), .A2(KEYINPUT31), .ZN(n1376) );
XOR2_X1 U1083 ( .A(n1392), .B(G146), .Z(n1391) );
NAND2_X1 U1084 ( .A1(n1393), .A2(n1394), .ZN(n1392) );
NAND2_X1 U1085 ( .A1(G140), .A2(n1305), .ZN(n1394) );
XOR2_X1 U1086 ( .A(KEYINPUT1), .B(n1395), .Z(n1393) );
NOR2_X1 U1087 ( .A1(G140), .A2(n1305), .ZN(n1395) );
INV_X1 U1088 ( .A(G125), .ZN(n1305) );
INV_X1 U1089 ( .A(n1136), .ZN(n1375) );
NAND2_X1 U1090 ( .A1(G217), .A2(n1340), .ZN(n1136) );
NAND2_X1 U1091 ( .A1(G234), .A2(n1343), .ZN(n1340) );
INV_X1 U1092 ( .A(n1293), .ZN(n1299) );
XOR2_X1 U1093 ( .A(n1129), .B(G472), .Z(n1293) );
NAND2_X1 U1094 ( .A1(n1396), .A2(n1343), .ZN(n1129) );
INV_X1 U1095 ( .A(G902), .ZN(n1343) );
XOR2_X1 U1096 ( .A(n1397), .B(n1398), .Z(n1396) );
XOR2_X1 U1097 ( .A(G101), .B(n1216), .Z(n1398) );
AND3_X1 U1098 ( .A1(n1339), .A2(n1095), .A3(n1399), .ZN(n1216) );
XOR2_X1 U1099 ( .A(KEYINPUT8), .B(G210), .Z(n1399) );
INV_X1 U1100 ( .A(G953), .ZN(n1095) );
INV_X1 U1101 ( .A(G237), .ZN(n1339) );
XOR2_X1 U1102 ( .A(n1215), .B(n1211), .Z(n1397) );
NAND2_X1 U1103 ( .A1(n1400), .A2(n1401), .ZN(n1211) );
NAND2_X1 U1104 ( .A1(n1371), .A2(G119), .ZN(n1401) );
NAND2_X1 U1105 ( .A1(n1402), .A2(n1314), .ZN(n1400) );
INV_X1 U1106 ( .A(G119), .ZN(n1314) );
XNOR2_X1 U1107 ( .A(n1371), .B(KEYINPUT28), .ZN(n1402) );
XOR2_X1 U1108 ( .A(n1403), .B(n1316), .Z(n1371) );
INV_X1 U1109 ( .A(G116), .ZN(n1316) );
INV_X1 U1110 ( .A(G113), .ZN(n1403) );
XOR2_X1 U1111 ( .A(n1242), .B(n1404), .Z(n1215) );
INV_X1 U1112 ( .A(n1370), .ZN(n1404) );
XOR2_X1 U1113 ( .A(n1405), .B(n1406), .Z(n1370) );
XOR2_X1 U1114 ( .A(G146), .B(G143), .Z(n1406) );
NAND2_X1 U1115 ( .A1(KEYINPUT16), .A2(G128), .ZN(n1405) );
XNOR2_X1 U1116 ( .A(n1407), .B(KEYINPUT5), .ZN(n1242) );
NAND3_X1 U1117 ( .A1(n1408), .A2(n1409), .A3(n1410), .ZN(n1407) );
OR2_X1 U1118 ( .A1(n1285), .A2(KEYINPUT0), .ZN(n1410) );
NAND3_X1 U1119 ( .A1(KEYINPUT0), .A2(n1285), .A3(n1167), .ZN(n1409) );
INV_X1 U1120 ( .A(n1411), .ZN(n1167) );
INV_X1 U1121 ( .A(G131), .ZN(n1285) );
NAND2_X1 U1122 ( .A1(n1411), .A2(n1412), .ZN(n1408) );
NAND2_X1 U1123 ( .A1(KEYINPUT0), .A2(n1413), .ZN(n1412) );
XOR2_X1 U1124 ( .A(KEYINPUT41), .B(G131), .Z(n1413) );
XOR2_X1 U1125 ( .A(G134), .B(n1383), .Z(n1411) );
XNOR2_X1 U1126 ( .A(G137), .B(KEYINPUT63), .ZN(n1383) );
INV_X1 U1127 ( .A(G110), .ZN(n1320) );
endmodule


