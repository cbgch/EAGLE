//Key = 1100010100001000011111111111111101011011000101011101011100110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300;

XNOR2_X1 U725 ( .A(G107), .B(n995), .ZN(G9) );
NOR2_X1 U726 ( .A1(n996), .A2(n997), .ZN(G75) );
NOR3_X1 U727 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
XNOR2_X1 U728 ( .A(n1001), .B(KEYINPUT41), .ZN(n999) );
NAND3_X1 U729 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n998) );
NAND2_X1 U730 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
NAND2_X1 U731 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND3_X1 U732 ( .A1(n1009), .A2(n1010), .A3(n1011), .ZN(n1008) );
NAND2_X1 U733 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NAND2_X1 U734 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
OR2_X1 U735 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NAND2_X1 U736 ( .A1(n1018), .A2(n1019), .ZN(n1012) );
NAND2_X1 U737 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NAND2_X1 U738 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND3_X1 U739 ( .A1(n1014), .A2(n1024), .A3(n1018), .ZN(n1007) );
NAND2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U741 ( .A1(n1011), .A2(n1027), .ZN(n1026) );
NAND2_X1 U742 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U743 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U744 ( .A1(n1009), .A2(n1032), .ZN(n1025) );
NAND2_X1 U745 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
XOR2_X1 U747 ( .A(n1037), .B(KEYINPUT42), .Z(n1035) );
INV_X1 U748 ( .A(n1038), .ZN(n1005) );
NOR3_X1 U749 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n996) );
INV_X1 U750 ( .A(n1002), .ZN(n1039) );
NAND4_X1 U751 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1002) );
NOR4_X1 U752 ( .A1(n1031), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1043) );
XOR2_X1 U753 ( .A(KEYINPUT56), .B(n1047), .Z(n1046) );
XNOR2_X1 U754 ( .A(KEYINPUT15), .B(n1023), .ZN(n1045) );
NOR3_X1 U755 ( .A1(n1048), .A2(n1036), .A3(n1022), .ZN(n1042) );
AND2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
XOR2_X1 U757 ( .A(KEYINPUT36), .B(n1051), .Z(n1041) );
NOR2_X1 U758 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
INV_X1 U759 ( .A(n1052), .ZN(n1050) );
XNOR2_X1 U760 ( .A(KEYINPUT22), .B(n1030), .ZN(n1040) );
XOR2_X1 U761 ( .A(n1053), .B(n1054), .Z(G72) );
NOR2_X1 U762 ( .A1(n1055), .A2(G953), .ZN(n1054) );
XOR2_X1 U763 ( .A(n1056), .B(n1057), .Z(n1053) );
NOR2_X1 U764 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U765 ( .A1(n1060), .A2(n1003), .ZN(n1058) );
XNOR2_X1 U766 ( .A(G227), .B(KEYINPUT47), .ZN(n1060) );
NAND2_X1 U767 ( .A1(n1061), .A2(n1062), .ZN(n1056) );
INV_X1 U768 ( .A(n1059), .ZN(n1062) );
XOR2_X1 U769 ( .A(n1063), .B(n1064), .Z(n1061) );
XNOR2_X1 U770 ( .A(n1065), .B(KEYINPUT10), .ZN(n1063) );
NAND2_X1 U771 ( .A1(n1066), .A2(n1067), .ZN(G69) );
NAND2_X1 U772 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
OR2_X1 U773 ( .A1(n1003), .A2(G224), .ZN(n1069) );
NAND3_X1 U774 ( .A1(G953), .A2(n1070), .A3(n1071), .ZN(n1066) );
INV_X1 U775 ( .A(n1068), .ZN(n1071) );
XNOR2_X1 U776 ( .A(n1072), .B(n1073), .ZN(n1068) );
NOR2_X1 U777 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
XOR2_X1 U778 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U779 ( .A(n1078), .B(n1079), .Z(n1077) );
XOR2_X1 U780 ( .A(n1080), .B(n1081), .Z(n1076) );
XOR2_X1 U781 ( .A(n1082), .B(n1083), .Z(n1080) );
NAND3_X1 U782 ( .A1(n1084), .A2(n1003), .A3(KEYINPUT21), .ZN(n1072) );
NAND3_X1 U783 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
XNOR2_X1 U784 ( .A(KEYINPUT45), .B(n1088), .ZN(n1085) );
NAND2_X1 U785 ( .A1(G898), .A2(G224), .ZN(n1070) );
NOR2_X1 U786 ( .A1(n1089), .A2(n1090), .ZN(G66) );
XNOR2_X1 U787 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR2_X1 U788 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR2_X1 U789 ( .A1(n1089), .A2(n1095), .ZN(G63) );
XOR2_X1 U790 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U791 ( .A1(KEYINPUT61), .A2(n1098), .ZN(n1096) );
NAND2_X1 U792 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
XNOR2_X1 U793 ( .A(G478), .B(KEYINPUT28), .ZN(n1099) );
NOR2_X1 U794 ( .A1(n1089), .A2(n1101), .ZN(G60) );
XNOR2_X1 U795 ( .A(n1102), .B(n1103), .ZN(n1101) );
AND2_X1 U796 ( .A1(G475), .A2(n1100), .ZN(n1103) );
XNOR2_X1 U797 ( .A(G104), .B(n1088), .ZN(G6) );
NOR2_X1 U798 ( .A1(n1089), .A2(n1104), .ZN(G57) );
XOR2_X1 U799 ( .A(n1105), .B(n1106), .Z(n1104) );
XOR2_X1 U800 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U801 ( .A(n1109), .B(n1110), .Z(n1105) );
NOR2_X1 U802 ( .A1(KEYINPUT44), .A2(n1111), .ZN(n1110) );
XNOR2_X1 U803 ( .A(n1112), .B(n1113), .ZN(n1109) );
AND2_X1 U804 ( .A1(G472), .A2(n1100), .ZN(n1113) );
NOR2_X1 U805 ( .A1(n1089), .A2(n1114), .ZN(G54) );
XOR2_X1 U806 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U807 ( .A(n1117), .B(n1064), .Z(n1116) );
XNOR2_X1 U808 ( .A(n1111), .B(G140), .ZN(n1064) );
XNOR2_X1 U809 ( .A(n1118), .B(n1119), .ZN(n1117) );
NAND2_X1 U810 ( .A1(KEYINPUT51), .A2(n1120), .ZN(n1119) );
NAND3_X1 U811 ( .A1(n1100), .A2(G469), .A3(KEYINPUT27), .ZN(n1118) );
INV_X1 U812 ( .A(n1094), .ZN(n1100) );
XOR2_X1 U813 ( .A(n1121), .B(n1122), .Z(n1115) );
NOR2_X1 U814 ( .A1(KEYINPUT40), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U815 ( .A(G110), .B(KEYINPUT50), .ZN(n1121) );
NOR3_X1 U816 ( .A1(n1089), .A2(n1124), .A3(n1125), .ZN(G51) );
NOR3_X1 U817 ( .A1(n1126), .A2(n1127), .A3(n1128), .ZN(n1125) );
XOR2_X1 U818 ( .A(KEYINPUT1), .B(n1129), .Z(n1128) );
NOR2_X1 U819 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
INV_X1 U820 ( .A(KEYINPUT52), .ZN(n1131) );
NOR2_X1 U821 ( .A1(n1132), .A2(n1133), .ZN(n1124) );
INV_X1 U822 ( .A(n1126), .ZN(n1133) );
XOR2_X1 U823 ( .A(n1134), .B(n1135), .Z(n1126) );
NAND2_X1 U824 ( .A1(KEYINPUT55), .A2(n1136), .ZN(n1134) );
NOR2_X1 U825 ( .A1(KEYINPUT52), .A2(n1130), .ZN(n1132) );
XNOR2_X1 U826 ( .A(n1129), .B(KEYINPUT9), .ZN(n1130) );
NOR2_X1 U827 ( .A1(n1094), .A2(n1052), .ZN(n1129) );
NAND2_X1 U828 ( .A1(G902), .A2(n1137), .ZN(n1094) );
NAND2_X1 U829 ( .A1(n1055), .A2(n1001), .ZN(n1137) );
AND3_X1 U830 ( .A1(n1138), .A2(n1088), .A3(n1087), .ZN(n1001) );
AND4_X1 U831 ( .A1(n1139), .A2(n995), .A3(n1140), .A4(n1141), .ZN(n1087) );
NOR3_X1 U832 ( .A1(n1142), .A2(n1143), .A3(n1144), .ZN(n1141) );
INV_X1 U833 ( .A(n1145), .ZN(n1143) );
AND3_X1 U834 ( .A1(n1146), .A2(n1017), .A3(n1147), .ZN(n1142) );
NAND3_X1 U835 ( .A1(n1017), .A2(n1009), .A3(n1148), .ZN(n995) );
NAND3_X1 U836 ( .A1(n1148), .A2(n1009), .A3(n1016), .ZN(n1088) );
XNOR2_X1 U837 ( .A(KEYINPUT49), .B(n1086), .ZN(n1138) );
INV_X1 U838 ( .A(n1000), .ZN(n1055) );
NAND4_X1 U839 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1000) );
NOR4_X1 U840 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1152) );
NOR3_X1 U841 ( .A1(n1157), .A2(n1158), .A3(n1159), .ZN(n1151) );
NOR2_X1 U842 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
INV_X1 U843 ( .A(KEYINPUT20), .ZN(n1160) );
NOR4_X1 U844 ( .A1(KEYINPUT20), .A2(n1162), .A3(n1163), .A4(n1028), .ZN(n1158) );
NAND3_X1 U845 ( .A1(n1164), .A2(n1020), .A3(n1016), .ZN(n1162) );
NOR2_X1 U846 ( .A1(n1003), .A2(G952), .ZN(n1089) );
XNOR2_X1 U847 ( .A(G146), .B(n1150), .ZN(G48) );
NAND3_X1 U848 ( .A1(n1016), .A2(n1165), .A3(n1166), .ZN(n1150) );
XOR2_X1 U849 ( .A(G143), .B(n1156), .Z(G45) );
AND4_X1 U850 ( .A1(n1167), .A2(n1165), .A3(n1147), .A4(n1168), .ZN(n1156) );
NOR3_X1 U851 ( .A1(n1020), .A2(n1169), .A3(n1170), .ZN(n1168) );
NAND2_X1 U852 ( .A1(n1171), .A2(n1172), .ZN(G42) );
NAND2_X1 U853 ( .A1(n1155), .A2(n1173), .ZN(n1172) );
XOR2_X1 U854 ( .A(KEYINPUT59), .B(n1174), .Z(n1171) );
NOR2_X1 U855 ( .A1(n1155), .A2(n1173), .ZN(n1174) );
AND3_X1 U856 ( .A1(n1175), .A2(n1176), .A3(n1011), .ZN(n1155) );
XNOR2_X1 U857 ( .A(n1177), .B(n1157), .ZN(G39) );
AND3_X1 U858 ( .A1(n1011), .A2(n1166), .A3(n1018), .ZN(n1157) );
INV_X1 U859 ( .A(n1163), .ZN(n1011) );
XNOR2_X1 U860 ( .A(G134), .B(n1149), .ZN(G36) );
NAND2_X1 U861 ( .A1(n1178), .A2(n1017), .ZN(n1149) );
XNOR2_X1 U862 ( .A(n1161), .B(n1179), .ZN(G33) );
NOR2_X1 U863 ( .A1(KEYINPUT4), .A2(n1180), .ZN(n1179) );
NAND2_X1 U864 ( .A1(n1178), .A2(n1016), .ZN(n1161) );
NOR4_X1 U865 ( .A1(n1028), .A2(n1163), .A3(n1020), .A4(n1169), .ZN(n1178) );
INV_X1 U866 ( .A(n1164), .ZN(n1169) );
NAND2_X1 U867 ( .A1(n1037), .A2(n1181), .ZN(n1163) );
INV_X1 U868 ( .A(n1147), .ZN(n1028) );
XOR2_X1 U869 ( .A(G128), .B(n1154), .Z(G30) );
AND3_X1 U870 ( .A1(n1017), .A2(n1165), .A3(n1166), .ZN(n1154) );
AND4_X1 U871 ( .A1(n1176), .A2(n1031), .A3(n1182), .A4(n1164), .ZN(n1166) );
NAND2_X1 U872 ( .A1(n1183), .A2(n1184), .ZN(G3) );
OR2_X1 U873 ( .A1(n1185), .A2(G101), .ZN(n1184) );
NAND2_X1 U874 ( .A1(G101), .A2(n1186), .ZN(n1183) );
NAND2_X1 U875 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
NAND2_X1 U876 ( .A1(n1144), .A2(n1189), .ZN(n1188) );
INV_X1 U877 ( .A(KEYINPUT54), .ZN(n1189) );
NAND2_X1 U878 ( .A1(KEYINPUT54), .A2(n1185), .ZN(n1187) );
NAND2_X1 U879 ( .A1(KEYINPUT38), .A2(n1144), .ZN(n1185) );
AND3_X1 U880 ( .A1(n1147), .A2(n1148), .A3(n1018), .ZN(n1144) );
XOR2_X1 U881 ( .A(G125), .B(n1153), .Z(G27) );
AND3_X1 U882 ( .A1(n1175), .A2(n1165), .A3(n1014), .ZN(n1153) );
AND4_X1 U883 ( .A1(n1030), .A2(n1016), .A3(n1031), .A4(n1164), .ZN(n1175) );
NAND2_X1 U884 ( .A1(n1038), .A2(n1190), .ZN(n1164) );
NAND3_X1 U885 ( .A1(G902), .A2(n1191), .A3(n1059), .ZN(n1190) );
NOR2_X1 U886 ( .A1(G900), .A2(n1003), .ZN(n1059) );
XNOR2_X1 U887 ( .A(G122), .B(n1145), .ZN(G24) );
NAND4_X1 U888 ( .A1(n1167), .A2(n1146), .A3(n1009), .A4(n1044), .ZN(n1145) );
NOR2_X1 U889 ( .A1(n1182), .A2(n1031), .ZN(n1009) );
XOR2_X1 U890 ( .A(n1140), .B(n1192), .Z(G21) );
NAND2_X1 U891 ( .A1(KEYINPUT39), .A2(G119), .ZN(n1192) );
NAND4_X1 U892 ( .A1(n1146), .A2(n1018), .A3(n1031), .A4(n1182), .ZN(n1140) );
XOR2_X1 U893 ( .A(n1193), .B(n1194), .Z(G18) );
NOR2_X1 U894 ( .A1(KEYINPUT16), .A2(n1195), .ZN(n1194) );
XOR2_X1 U895 ( .A(KEYINPUT13), .B(G116), .Z(n1195) );
NAND4_X1 U896 ( .A1(n1147), .A2(n1014), .A3(n1196), .A4(n1017), .ZN(n1193) );
NOR2_X1 U897 ( .A1(n1170), .A2(n1167), .ZN(n1017) );
NOR2_X1 U898 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
XNOR2_X1 U899 ( .A(n1165), .B(KEYINPUT8), .ZN(n1198) );
XNOR2_X1 U900 ( .A(G113), .B(n1139), .ZN(G15) );
NAND3_X1 U901 ( .A1(n1147), .A2(n1016), .A3(n1146), .ZN(n1139) );
AND3_X1 U902 ( .A1(n1165), .A2(n1199), .A3(n1014), .ZN(n1146) );
NOR2_X1 U903 ( .A1(n1200), .A2(n1022), .ZN(n1014) );
AND2_X1 U904 ( .A1(n1167), .A2(n1170), .ZN(n1016) );
INV_X1 U905 ( .A(n1044), .ZN(n1170) );
NOR2_X1 U906 ( .A1(n1031), .A2(n1030), .ZN(n1147) );
XOR2_X1 U907 ( .A(n1086), .B(n1201), .Z(G12) );
NAND2_X1 U908 ( .A1(n1202), .A2(G110), .ZN(n1201) );
XNOR2_X1 U909 ( .A(KEYINPUT5), .B(KEYINPUT25), .ZN(n1202) );
NAND4_X1 U910 ( .A1(n1018), .A2(n1148), .A3(n1030), .A4(n1031), .ZN(n1086) );
XOR2_X1 U911 ( .A(n1203), .B(n1093), .Z(n1031) );
NAND2_X1 U912 ( .A1(G217), .A2(n1204), .ZN(n1093) );
NAND2_X1 U913 ( .A1(n1091), .A2(n1205), .ZN(n1203) );
XNOR2_X1 U914 ( .A(n1206), .B(n1207), .ZN(n1091) );
XOR2_X1 U915 ( .A(n1208), .B(n1083), .Z(n1207) );
XOR2_X1 U916 ( .A(G119), .B(G110), .Z(n1083) );
XOR2_X1 U917 ( .A(n1209), .B(n1210), .Z(n1206) );
NOR2_X1 U918 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U919 ( .A(n1213), .B(KEYINPUT7), .Z(n1212) );
NAND3_X1 U920 ( .A1(G137), .A2(G221), .A3(n1214), .ZN(n1213) );
NOR2_X1 U921 ( .A1(n1215), .A2(n1216), .ZN(n1211) );
XNOR2_X1 U922 ( .A(G137), .B(KEYINPUT58), .ZN(n1216) );
AND2_X1 U923 ( .A1(G221), .A2(n1214), .ZN(n1215) );
XOR2_X1 U924 ( .A(n1217), .B(KEYINPUT60), .Z(n1209) );
NAND3_X1 U925 ( .A1(n1218), .A2(n1219), .A3(n1220), .ZN(n1217) );
NAND2_X1 U926 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
INV_X1 U927 ( .A(KEYINPUT18), .ZN(n1222) );
NAND3_X1 U928 ( .A1(KEYINPUT18), .A2(n1223), .A3(G125), .ZN(n1219) );
OR2_X1 U929 ( .A1(n1223), .A2(G125), .ZN(n1218) );
NOR2_X1 U930 ( .A1(KEYINPUT46), .A2(n1221), .ZN(n1223) );
XNOR2_X1 U931 ( .A(n1173), .B(KEYINPUT30), .ZN(n1221) );
INV_X1 U932 ( .A(n1182), .ZN(n1030) );
XNOR2_X1 U933 ( .A(n1224), .B(G472), .ZN(n1182) );
NAND2_X1 U934 ( .A1(n1225), .A2(n1205), .ZN(n1224) );
XOR2_X1 U935 ( .A(n1226), .B(n1227), .Z(n1225) );
XOR2_X1 U936 ( .A(n1107), .B(n1228), .Z(n1227) );
NOR2_X1 U937 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
AND2_X1 U938 ( .A1(KEYINPUT48), .A2(n1231), .ZN(n1230) );
NOR2_X1 U939 ( .A1(KEYINPUT33), .A2(n1231), .ZN(n1229) );
XOR2_X1 U940 ( .A(n1111), .B(n1108), .Z(n1231) );
XNOR2_X1 U941 ( .A(n1232), .B(n1081), .ZN(n1107) );
XOR2_X1 U942 ( .A(G101), .B(G116), .Z(n1081) );
XNOR2_X1 U943 ( .A(n1233), .B(n1234), .ZN(n1232) );
NOR2_X1 U944 ( .A1(G119), .A2(KEYINPUT37), .ZN(n1234) );
NOR2_X1 U945 ( .A1(KEYINPUT3), .A2(n1235), .ZN(n1233) );
XOR2_X1 U946 ( .A(KEYINPUT6), .B(G113), .Z(n1235) );
XOR2_X1 U947 ( .A(n1236), .B(KEYINPUT12), .Z(n1226) );
NAND2_X1 U948 ( .A1(KEYINPUT63), .A2(n1112), .ZN(n1236) );
AND3_X1 U949 ( .A1(n1237), .A2(n1003), .A3(G210), .ZN(n1112) );
NOR3_X1 U950 ( .A1(n1020), .A2(n1197), .A3(n1033), .ZN(n1148) );
INV_X1 U951 ( .A(n1165), .ZN(n1033) );
NOR2_X1 U952 ( .A1(n1037), .A2(n1036), .ZN(n1165) );
INV_X1 U953 ( .A(n1181), .ZN(n1036) );
NAND2_X1 U954 ( .A1(G214), .A2(n1238), .ZN(n1181) );
XOR2_X1 U955 ( .A(n1049), .B(n1239), .Z(n1037) );
XNOR2_X1 U956 ( .A(KEYINPUT14), .B(n1052), .ZN(n1239) );
NAND2_X1 U957 ( .A1(G210), .A2(n1238), .ZN(n1052) );
NAND2_X1 U958 ( .A1(n1240), .A2(n1237), .ZN(n1238) );
NAND2_X1 U959 ( .A1(n1241), .A2(n1205), .ZN(n1049) );
XNOR2_X1 U960 ( .A(n1242), .B(n1136), .ZN(n1241) );
XOR2_X1 U961 ( .A(n1243), .B(n1244), .Z(n1136) );
INV_X1 U962 ( .A(n1065), .ZN(n1244) );
XOR2_X1 U963 ( .A(G125), .B(n1108), .Z(n1065) );
NAND2_X1 U964 ( .A1(G224), .A2(n1003), .ZN(n1243) );
NAND2_X1 U965 ( .A1(KEYINPUT62), .A2(n1135), .ZN(n1242) );
XOR2_X1 U966 ( .A(n1245), .B(n1246), .Z(n1135) );
XNOR2_X1 U967 ( .A(n1247), .B(G110), .ZN(n1246) );
NAND4_X1 U968 ( .A1(KEYINPUT19), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1245) );
NAND3_X1 U969 ( .A1(KEYINPUT23), .A2(n1251), .A3(n1252), .ZN(n1250) );
OR2_X1 U970 ( .A1(n1252), .A2(n1251), .ZN(n1249) );
NOR2_X1 U971 ( .A1(KEYINPUT57), .A2(n1253), .ZN(n1251) );
XNOR2_X1 U972 ( .A(n1254), .B(n1079), .ZN(n1252) );
XNOR2_X1 U973 ( .A(n1255), .B(KEYINPUT43), .ZN(n1079) );
NAND2_X1 U974 ( .A1(KEYINPUT35), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U975 ( .A(G101), .B(G107), .ZN(n1254) );
NAND2_X1 U976 ( .A1(n1253), .A2(n1257), .ZN(n1248) );
INV_X1 U977 ( .A(KEYINPUT23), .ZN(n1257) );
XOR2_X1 U978 ( .A(n1082), .B(n1258), .Z(n1253) );
XOR2_X1 U979 ( .A(G119), .B(G116), .Z(n1258) );
NAND2_X1 U980 ( .A1(n1259), .A2(KEYINPUT17), .ZN(n1082) );
XNOR2_X1 U981 ( .A(KEYINPUT6), .B(G113), .ZN(n1259) );
INV_X1 U982 ( .A(n1199), .ZN(n1197) );
NAND2_X1 U983 ( .A1(n1038), .A2(n1260), .ZN(n1199) );
NAND3_X1 U984 ( .A1(G902), .A2(n1191), .A3(n1074), .ZN(n1260) );
NOR2_X1 U985 ( .A1(n1003), .A2(G898), .ZN(n1074) );
NAND3_X1 U986 ( .A1(n1191), .A2(n1003), .A3(G952), .ZN(n1038) );
NAND2_X1 U987 ( .A1(G237), .A2(G234), .ZN(n1191) );
INV_X1 U988 ( .A(n1176), .ZN(n1020) );
NOR2_X1 U989 ( .A1(n1023), .A2(n1022), .ZN(n1176) );
AND2_X1 U990 ( .A1(G221), .A2(n1204), .ZN(n1022) );
NAND2_X1 U991 ( .A1(G234), .A2(n1240), .ZN(n1204) );
XNOR2_X1 U992 ( .A(n1205), .B(KEYINPUT29), .ZN(n1240) );
INV_X1 U993 ( .A(n1200), .ZN(n1023) );
XNOR2_X1 U994 ( .A(n1261), .B(G469), .ZN(n1200) );
NAND2_X1 U995 ( .A1(n1262), .A2(n1205), .ZN(n1261) );
XOR2_X1 U996 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U997 ( .A(n1123), .B(n1265), .ZN(n1264) );
NOR2_X1 U998 ( .A1(KEYINPUT2), .A2(n1111), .ZN(n1265) );
XNOR2_X1 U999 ( .A(G131), .B(n1266), .ZN(n1111) );
XNOR2_X1 U1000 ( .A(n1177), .B(G134), .ZN(n1266) );
INV_X1 U1001 ( .A(G137), .ZN(n1177) );
XNOR2_X1 U1002 ( .A(n1267), .B(n1108), .ZN(n1123) );
XOR2_X1 U1003 ( .A(G143), .B(n1208), .Z(n1108) );
XOR2_X1 U1004 ( .A(G146), .B(n1268), .Z(n1208) );
XOR2_X1 U1005 ( .A(n1269), .B(G101), .Z(n1267) );
NAND2_X1 U1006 ( .A1(KEYINPUT53), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U1007 ( .A(n1271), .B(G104), .ZN(n1270) );
INV_X1 U1008 ( .A(G107), .ZN(n1271) );
XNOR2_X1 U1009 ( .A(n1120), .B(n1272), .ZN(n1263) );
NOR2_X1 U1010 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NOR2_X1 U1011 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NOR2_X1 U1012 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
INV_X1 U1013 ( .A(KEYINPUT0), .ZN(n1278) );
NOR2_X1 U1014 ( .A1(G110), .A2(KEYINPUT11), .ZN(n1277) );
NOR2_X1 U1015 ( .A1(n1279), .A2(n1280), .ZN(n1273) );
INV_X1 U1016 ( .A(G110), .ZN(n1280) );
NOR2_X1 U1017 ( .A1(n1281), .A2(KEYINPUT11), .ZN(n1279) );
AND2_X1 U1018 ( .A1(n1276), .A2(KEYINPUT0), .ZN(n1281) );
XNOR2_X1 U1019 ( .A(G140), .B(KEYINPUT24), .ZN(n1276) );
AND2_X1 U1020 ( .A1(G227), .A2(n1003), .ZN(n1120) );
NOR2_X1 U1021 ( .A1(n1044), .A2(n1167), .ZN(n1018) );
XNOR2_X1 U1022 ( .A(n1047), .B(KEYINPUT26), .ZN(n1167) );
XNOR2_X1 U1023 ( .A(n1282), .B(G475), .ZN(n1047) );
NAND2_X1 U1024 ( .A1(n1102), .A2(n1205), .ZN(n1282) );
INV_X1 U1025 ( .A(G902), .ZN(n1205) );
XNOR2_X1 U1026 ( .A(n1283), .B(n1284), .ZN(n1102) );
XNOR2_X1 U1027 ( .A(n1247), .B(G113), .ZN(n1284) );
XNOR2_X1 U1028 ( .A(n1285), .B(n1256), .ZN(n1283) );
INV_X1 U1029 ( .A(G104), .ZN(n1256) );
NAND2_X1 U1030 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U1031 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XOR2_X1 U1032 ( .A(KEYINPUT31), .B(n1290), .Z(n1286) );
NOR2_X1 U1033 ( .A1(n1288), .A2(n1289), .ZN(n1290) );
XOR2_X1 U1034 ( .A(n1291), .B(n1292), .Z(n1289) );
XNOR2_X1 U1035 ( .A(G143), .B(n1180), .ZN(n1292) );
INV_X1 U1036 ( .A(G131), .ZN(n1180) );
NAND3_X1 U1037 ( .A1(n1237), .A2(n1003), .A3(G214), .ZN(n1291) );
INV_X1 U1038 ( .A(G237), .ZN(n1237) );
XNOR2_X1 U1039 ( .A(G125), .B(n1293), .ZN(n1288) );
XNOR2_X1 U1040 ( .A(G146), .B(n1173), .ZN(n1293) );
INV_X1 U1041 ( .A(G140), .ZN(n1173) );
XNOR2_X1 U1042 ( .A(n1294), .B(G478), .ZN(n1044) );
OR2_X1 U1043 ( .A1(n1097), .A2(G902), .ZN(n1294) );
XNOR2_X1 U1044 ( .A(n1295), .B(n1296), .ZN(n1097) );
XNOR2_X1 U1045 ( .A(n1078), .B(n1297), .ZN(n1296) );
XOR2_X1 U1046 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U1047 ( .A1(KEYINPUT32), .A2(n1268), .ZN(n1299) );
XOR2_X1 U1048 ( .A(G128), .B(KEYINPUT34), .Z(n1268) );
NAND2_X1 U1049 ( .A1(G217), .A2(n1214), .ZN(n1298) );
AND2_X1 U1050 ( .A1(G234), .A2(n1003), .ZN(n1214) );
INV_X1 U1051 ( .A(G953), .ZN(n1003) );
XNOR2_X1 U1052 ( .A(G107), .B(n1247), .ZN(n1078) );
INV_X1 U1053 ( .A(G122), .ZN(n1247) );
XNOR2_X1 U1054 ( .A(G116), .B(n1300), .ZN(n1295) );
XOR2_X1 U1055 ( .A(G143), .B(G134), .Z(n1300) );
endmodule


