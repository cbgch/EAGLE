//Key = 0001111100000010100101101110101101101000101010011100011001100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;

NAND2_X1 U737 ( .A1(n1031), .A2(n1032), .ZN(G9) );
NAND2_X1 U738 ( .A1(G107), .A2(n1033), .ZN(n1032) );
XOR2_X1 U739 ( .A(n1034), .B(KEYINPUT17), .Z(n1031) );
OR2_X1 U740 ( .A1(n1033), .A2(G107), .ZN(n1034) );
NAND4_X1 U741 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(G75) );
NAND4_X1 U742 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1037) );
NOR4_X1 U743 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NOR3_X1 U744 ( .A1(n1047), .A2(KEYINPUT10), .A3(n1048), .ZN(n1046) );
AND2_X1 U745 ( .A1(n1047), .A2(KEYINPUT10), .ZN(n1045) );
XNOR2_X1 U746 ( .A(G469), .B(n1049), .ZN(n1044) );
NAND3_X1 U747 ( .A1(n1050), .A2(n1051), .A3(n1052), .ZN(n1043) );
XOR2_X1 U748 ( .A(n1053), .B(n1054), .Z(n1052) );
XOR2_X1 U749 ( .A(n1055), .B(KEYINPUT39), .Z(n1050) );
NOR3_X1 U750 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1041) );
INV_X1 U751 ( .A(n1059), .ZN(n1058) );
NAND2_X1 U752 ( .A1(n1060), .A2(n1061), .ZN(n1036) );
NAND2_X1 U753 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND4_X1 U754 ( .A1(n1039), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1063) );
NAND2_X1 U755 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U756 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1067) );
INV_X1 U757 ( .A(KEYINPUT4), .ZN(n1070) );
NAND3_X1 U758 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1065) );
NAND2_X1 U759 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
OR2_X1 U760 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NAND2_X1 U761 ( .A1(n1069), .A2(n1079), .ZN(n1072) );
NAND2_X1 U762 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
NAND2_X1 U763 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
INV_X1 U764 ( .A(n1040), .ZN(n1082) );
NAND2_X1 U765 ( .A1(KEYINPUT4), .A2(n1071), .ZN(n1080) );
NAND3_X1 U766 ( .A1(n1069), .A2(n1084), .A3(n1075), .ZN(n1062) );
NAND2_X1 U767 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND3_X1 U768 ( .A1(n1087), .A2(n1088), .A3(n1039), .ZN(n1086) );
NAND2_X1 U769 ( .A1(n1089), .A2(n1068), .ZN(n1088) );
NAND3_X1 U770 ( .A1(n1090), .A2(n1091), .A3(n1064), .ZN(n1087) );
NAND2_X1 U771 ( .A1(n1092), .A2(n1057), .ZN(n1090) );
NAND2_X1 U772 ( .A1(n1074), .A2(n1093), .ZN(n1085) );
INV_X1 U773 ( .A(n1068), .ZN(n1074) );
INV_X1 U774 ( .A(n1094), .ZN(n1060) );
XOR2_X1 U775 ( .A(n1095), .B(n1096), .Z(G72) );
NOR2_X1 U776 ( .A1(KEYINPUT38), .A2(n1097), .ZN(n1096) );
XOR2_X1 U777 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U778 ( .A1(n1100), .A2(G953), .ZN(n1099) );
NOR3_X1 U779 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1098) );
NOR2_X1 U780 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U781 ( .A(n1106), .B(KEYINPUT54), .Z(n1105) );
NOR2_X1 U782 ( .A1(n1107), .A2(n1106), .ZN(n1102) );
XNOR2_X1 U783 ( .A(n1108), .B(n1109), .ZN(n1106) );
NAND2_X1 U784 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
INV_X1 U785 ( .A(n1112), .ZN(n1110) );
NAND2_X1 U786 ( .A1(G953), .A2(n1113), .ZN(n1095) );
NAND2_X1 U787 ( .A1(G900), .A2(G227), .ZN(n1113) );
XOR2_X1 U788 ( .A(n1114), .B(n1115), .Z(G69) );
XOR2_X1 U789 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U790 ( .A1(G953), .A2(n1118), .ZN(n1117) );
NAND2_X1 U791 ( .A1(G898), .A2(G224), .ZN(n1118) );
NAND3_X1 U792 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1116) );
NAND2_X1 U793 ( .A1(G953), .A2(n1122), .ZN(n1121) );
NAND2_X1 U794 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
NAND2_X1 U795 ( .A1(n1125), .A2(n1126), .ZN(n1119) );
INV_X1 U796 ( .A(n1123), .ZN(n1126) );
XNOR2_X1 U797 ( .A(KEYINPUT12), .B(n1124), .ZN(n1125) );
NOR2_X1 U798 ( .A1(n1127), .A2(G953), .ZN(n1114) );
NOR2_X1 U799 ( .A1(n1128), .A2(n1129), .ZN(G66) );
NOR3_X1 U800 ( .A1(n1053), .A2(n1130), .A3(n1131), .ZN(n1129) );
AND3_X1 U801 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR2_X1 U802 ( .A1(n1135), .A2(n1132), .ZN(n1130) );
NOR2_X1 U803 ( .A1(n1035), .A2(n1054), .ZN(n1135) );
NOR2_X1 U804 ( .A1(n1128), .A2(n1136), .ZN(G63) );
XNOR2_X1 U805 ( .A(n1137), .B(n1138), .ZN(n1136) );
AND2_X1 U806 ( .A1(G478), .A2(n1134), .ZN(n1137) );
NOR2_X1 U807 ( .A1(n1128), .A2(n1139), .ZN(G60) );
NOR2_X1 U808 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
NOR2_X1 U809 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NOR2_X1 U810 ( .A1(n1144), .A2(n1145), .ZN(n1140) );
XOR2_X1 U811 ( .A(KEYINPUT22), .B(n1142), .Z(n1145) );
AND2_X1 U812 ( .A1(n1134), .A2(G475), .ZN(n1142) );
XNOR2_X1 U813 ( .A(n1143), .B(KEYINPUT0), .ZN(n1144) );
XNOR2_X1 U814 ( .A(G104), .B(n1146), .ZN(G6) );
NOR2_X1 U815 ( .A1(n1128), .A2(n1147), .ZN(G57) );
XOR2_X1 U816 ( .A(n1148), .B(n1149), .Z(n1147) );
XNOR2_X1 U817 ( .A(G101), .B(n1150), .ZN(n1149) );
NAND3_X1 U818 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NAND2_X1 U819 ( .A1(KEYINPUT20), .A2(n1154), .ZN(n1153) );
OR3_X1 U820 ( .A1(n1154), .A2(KEYINPUT20), .A3(n1155), .ZN(n1152) );
NAND2_X1 U821 ( .A1(n1155), .A2(n1156), .ZN(n1151) );
NAND2_X1 U822 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
INV_X1 U823 ( .A(KEYINPUT20), .ZN(n1158) );
XNOR2_X1 U824 ( .A(n1154), .B(KEYINPUT45), .ZN(n1157) );
XOR2_X1 U825 ( .A(n1159), .B(n1160), .Z(n1148) );
AND2_X1 U826 ( .A1(G472), .A2(n1134), .ZN(n1160) );
NOR2_X1 U827 ( .A1(n1128), .A2(n1161), .ZN(G54) );
NOR2_X1 U828 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U829 ( .A(n1164), .B(n1165), .Z(n1163) );
AND2_X1 U830 ( .A1(n1166), .A2(KEYINPUT6), .ZN(n1165) );
AND2_X1 U831 ( .A1(G469), .A2(n1134), .ZN(n1164) );
NOR2_X1 U832 ( .A1(KEYINPUT6), .A2(n1166), .ZN(n1162) );
XNOR2_X1 U833 ( .A(n1167), .B(n1168), .ZN(n1166) );
XOR2_X1 U834 ( .A(n1169), .B(n1170), .Z(n1168) );
NAND2_X1 U835 ( .A1(n1171), .A2(KEYINPUT16), .ZN(n1170) );
XOR2_X1 U836 ( .A(n1172), .B(G140), .Z(n1171) );
NAND2_X1 U837 ( .A1(KEYINPUT24), .A2(n1173), .ZN(n1172) );
XOR2_X1 U838 ( .A(n1174), .B(n1175), .Z(n1167) );
NAND2_X1 U839 ( .A1(n1176), .A2(n1177), .ZN(n1174) );
NAND2_X1 U840 ( .A1(KEYINPUT44), .A2(n1178), .ZN(n1177) );
XOR2_X1 U841 ( .A(n1179), .B(n1107), .Z(n1178) );
OR3_X1 U842 ( .A1(n1179), .A2(n1107), .A3(KEYINPUT44), .ZN(n1176) );
NOR2_X1 U843 ( .A1(n1128), .A2(n1180), .ZN(G51) );
XOR2_X1 U844 ( .A(n1181), .B(n1182), .Z(n1180) );
XNOR2_X1 U845 ( .A(n1183), .B(n1184), .ZN(n1182) );
NAND2_X1 U846 ( .A1(KEYINPUT36), .A2(n1185), .ZN(n1183) );
XOR2_X1 U847 ( .A(n1107), .B(n1186), .Z(n1185) );
XNOR2_X1 U848 ( .A(n1187), .B(KEYINPUT61), .ZN(n1186) );
NAND2_X1 U849 ( .A1(KEYINPUT5), .A2(n1188), .ZN(n1187) );
XOR2_X1 U850 ( .A(n1189), .B(n1190), .Z(n1181) );
NAND3_X1 U851 ( .A1(n1134), .A2(G210), .A3(KEYINPUT26), .ZN(n1189) );
NOR2_X1 U852 ( .A1(n1191), .A2(n1035), .ZN(n1134) );
AND2_X1 U853 ( .A1(n1127), .A2(n1100), .ZN(n1035) );
AND2_X1 U854 ( .A1(n1192), .A2(n1193), .ZN(n1100) );
NOR4_X1 U855 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1193) );
AND4_X1 U856 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1192) );
OR2_X1 U857 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XOR2_X1 U858 ( .A(n1204), .B(KEYINPUT59), .Z(n1202) );
AND2_X1 U859 ( .A1(n1205), .A2(n1206), .ZN(n1127) );
AND4_X1 U860 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
AND4_X1 U861 ( .A1(n1033), .A2(n1211), .A3(n1212), .A4(n1146), .ZN(n1205) );
NAND3_X1 U862 ( .A1(n1213), .A2(n1064), .A3(n1078), .ZN(n1146) );
NAND3_X1 U863 ( .A1(n1213), .A2(n1064), .A3(n1077), .ZN(n1033) );
NOR2_X1 U864 ( .A1(n1214), .A2(G952), .ZN(n1128) );
XOR2_X1 U865 ( .A(G953), .B(KEYINPUT34), .Z(n1214) );
XOR2_X1 U866 ( .A(G146), .B(n1197), .Z(G48) );
AND3_X1 U867 ( .A1(n1078), .A2(n1071), .A3(n1215), .ZN(n1197) );
NAND2_X1 U868 ( .A1(n1216), .A2(n1217), .ZN(G45) );
NAND2_X1 U869 ( .A1(n1196), .A2(n1218), .ZN(n1217) );
XOR2_X1 U870 ( .A(KEYINPUT57), .B(n1219), .Z(n1216) );
NOR2_X1 U871 ( .A1(n1196), .A2(n1218), .ZN(n1219) );
INV_X1 U872 ( .A(G143), .ZN(n1218) );
AND4_X1 U873 ( .A1(n1071), .A2(n1220), .A3(n1093), .A4(n1221), .ZN(n1196) );
NOR3_X1 U874 ( .A1(n1222), .A2(n1223), .A3(n1051), .ZN(n1221) );
XNOR2_X1 U875 ( .A(n1195), .B(n1224), .ZN(G42) );
NAND2_X1 U876 ( .A1(KEYINPUT42), .A2(G140), .ZN(n1224) );
AND4_X1 U877 ( .A1(n1089), .A2(n1225), .A3(n1039), .A4(n1078), .ZN(n1195) );
NAND3_X1 U878 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(G39) );
NAND2_X1 U879 ( .A1(KEYINPUT9), .A2(n1229), .ZN(n1228) );
NAND3_X1 U880 ( .A1(G137), .A2(n1230), .A3(n1200), .ZN(n1227) );
NAND2_X1 U881 ( .A1(n1231), .A2(n1232), .ZN(n1226) );
NAND2_X1 U882 ( .A1(n1233), .A2(n1230), .ZN(n1232) );
INV_X1 U883 ( .A(KEYINPUT9), .ZN(n1230) );
XOR2_X1 U884 ( .A(KEYINPUT11), .B(G137), .Z(n1233) );
INV_X1 U885 ( .A(n1200), .ZN(n1231) );
NAND4_X1 U886 ( .A1(n1089), .A2(n1225), .A3(n1069), .A4(n1234), .ZN(n1200) );
XOR2_X1 U887 ( .A(G134), .B(n1235), .Z(G36) );
NOR2_X1 U888 ( .A1(n1204), .A2(n1203), .ZN(n1235) );
NAND2_X1 U889 ( .A1(n1225), .A2(n1077), .ZN(n1203) );
XNOR2_X1 U890 ( .A(G131), .B(n1199), .ZN(G33) );
NAND3_X1 U891 ( .A1(n1093), .A2(n1078), .A3(n1225), .ZN(n1199) );
NOR3_X1 U892 ( .A1(n1236), .A2(n1223), .A3(n1068), .ZN(n1225) );
NAND2_X1 U893 ( .A1(n1092), .A2(n1237), .ZN(n1068) );
XOR2_X1 U894 ( .A(n1238), .B(KEYINPUT40), .Z(n1092) );
XOR2_X1 U895 ( .A(G128), .B(n1194), .Z(G30) );
AND3_X1 U896 ( .A1(n1077), .A2(n1239), .A3(n1215), .ZN(n1194) );
NOR4_X1 U897 ( .A1(n1064), .A2(n1091), .A3(n1039), .A4(n1223), .ZN(n1215) );
XNOR2_X1 U898 ( .A(G101), .B(n1212), .ZN(G3) );
NAND4_X1 U899 ( .A1(n1093), .A2(n1240), .A3(n1069), .A4(n1239), .ZN(n1212) );
XOR2_X1 U900 ( .A(n1188), .B(n1198), .Z(G27) );
NAND4_X1 U901 ( .A1(n1078), .A2(n1075), .A3(n1089), .A4(n1241), .ZN(n1198) );
NOR3_X1 U902 ( .A1(n1234), .A2(n1223), .A3(n1091), .ZN(n1241) );
AND2_X1 U903 ( .A1(n1242), .A2(n1094), .ZN(n1223) );
NAND3_X1 U904 ( .A1(G902), .A2(n1243), .A3(n1101), .ZN(n1242) );
NOR2_X1 U905 ( .A1(n1038), .A2(G900), .ZN(n1101) );
INV_X1 U906 ( .A(G125), .ZN(n1188) );
XOR2_X1 U907 ( .A(n1210), .B(n1244), .Z(G24) );
XNOR2_X1 U908 ( .A(G122), .B(KEYINPUT60), .ZN(n1244) );
NAND3_X1 U909 ( .A1(n1039), .A2(n1245), .A3(n1246), .ZN(n1210) );
NOR3_X1 U910 ( .A1(n1222), .A2(n1051), .A3(n1089), .ZN(n1246) );
XOR2_X1 U911 ( .A(n1247), .B(KEYINPUT33), .Z(n1222) );
XNOR2_X1 U912 ( .A(G119), .B(n1209), .ZN(G21) );
NAND4_X1 U913 ( .A1(n1089), .A2(n1245), .A3(n1069), .A4(n1234), .ZN(n1209) );
XOR2_X1 U914 ( .A(n1248), .B(n1208), .Z(G18) );
NAND3_X1 U915 ( .A1(n1245), .A2(n1077), .A3(n1093), .ZN(n1208) );
XNOR2_X1 U916 ( .A(G113), .B(n1207), .ZN(G15) );
NAND3_X1 U917 ( .A1(n1245), .A2(n1078), .A3(n1093), .ZN(n1207) );
INV_X1 U918 ( .A(n1204), .ZN(n1093) );
NAND2_X1 U919 ( .A1(n1064), .A2(n1234), .ZN(n1204) );
INV_X1 U920 ( .A(n1039), .ZN(n1234) );
INV_X1 U921 ( .A(n1089), .ZN(n1064) );
AND2_X1 U922 ( .A1(n1249), .A2(n1247), .ZN(n1078) );
XOR2_X1 U923 ( .A(KEYINPUT43), .B(n1051), .Z(n1249) );
AND2_X1 U924 ( .A1(n1075), .A2(n1240), .ZN(n1245) );
AND2_X1 U925 ( .A1(n1083), .A2(n1040), .ZN(n1075) );
XOR2_X1 U926 ( .A(n1250), .B(KEYINPUT21), .Z(n1083) );
NAND2_X1 U927 ( .A1(n1251), .A2(n1252), .ZN(G12) );
NAND2_X1 U928 ( .A1(G110), .A2(n1211), .ZN(n1252) );
XOR2_X1 U929 ( .A(n1253), .B(KEYINPUT37), .Z(n1251) );
OR2_X1 U930 ( .A1(n1211), .A2(G110), .ZN(n1253) );
NAND3_X1 U931 ( .A1(n1213), .A2(n1069), .A3(n1089), .ZN(n1211) );
XNOR2_X1 U932 ( .A(n1053), .B(n1254), .ZN(n1089) );
NOR2_X1 U933 ( .A1(n1133), .A2(KEYINPUT35), .ZN(n1254) );
INV_X1 U934 ( .A(n1054), .ZN(n1133) );
NAND2_X1 U935 ( .A1(G217), .A2(n1255), .ZN(n1054) );
NOR2_X1 U936 ( .A1(n1132), .A2(G902), .ZN(n1053) );
XNOR2_X1 U937 ( .A(n1256), .B(n1257), .ZN(n1132) );
XNOR2_X1 U938 ( .A(n1258), .B(n1259), .ZN(n1257) );
XOR2_X1 U939 ( .A(n1260), .B(n1261), .Z(n1259) );
NOR2_X1 U940 ( .A1(G110), .A2(KEYINPUT15), .ZN(n1261) );
NAND2_X1 U941 ( .A1(G221), .A2(n1262), .ZN(n1260) );
XOR2_X1 U942 ( .A(n1263), .B(n1264), .Z(n1256) );
XOR2_X1 U943 ( .A(G137), .B(G128), .Z(n1264) );
NAND2_X1 U944 ( .A1(KEYINPUT28), .A2(n1265), .ZN(n1263) );
XOR2_X1 U945 ( .A(n1266), .B(n1267), .Z(n1265) );
XOR2_X1 U946 ( .A(n1268), .B(G140), .Z(n1267) );
INV_X1 U947 ( .A(G146), .ZN(n1268) );
NAND2_X1 U948 ( .A1(KEYINPUT31), .A2(G125), .ZN(n1266) );
NAND2_X1 U949 ( .A1(n1269), .A2(n1270), .ZN(n1069) );
OR3_X1 U950 ( .A1(n1247), .A2(n1271), .A3(KEYINPUT43), .ZN(n1270) );
INV_X1 U951 ( .A(n1051), .ZN(n1271) );
NAND2_X1 U952 ( .A1(KEYINPUT43), .A2(n1077), .ZN(n1269) );
NOR2_X1 U953 ( .A1(n1247), .A2(n1051), .ZN(n1077) );
XOR2_X1 U954 ( .A(n1272), .B(G478), .Z(n1051) );
NAND2_X1 U955 ( .A1(n1138), .A2(n1273), .ZN(n1272) );
XOR2_X1 U956 ( .A(KEYINPUT30), .B(G902), .Z(n1273) );
XOR2_X1 U957 ( .A(n1274), .B(n1275), .Z(n1138) );
XOR2_X1 U958 ( .A(n1276), .B(n1277), .Z(n1275) );
NAND2_X1 U959 ( .A1(n1278), .A2(KEYINPUT48), .ZN(n1277) );
XNOR2_X1 U960 ( .A(G128), .B(n1279), .ZN(n1278) );
XOR2_X1 U961 ( .A(G143), .B(G134), .Z(n1279) );
NAND2_X1 U962 ( .A1(n1280), .A2(n1281), .ZN(n1276) );
NAND2_X1 U963 ( .A1(G122), .A2(n1248), .ZN(n1281) );
XOR2_X1 U964 ( .A(n1282), .B(KEYINPUT55), .Z(n1280) );
OR2_X1 U965 ( .A1(n1248), .A2(G122), .ZN(n1282) );
XOR2_X1 U966 ( .A(n1283), .B(n1284), .Z(n1274) );
NOR2_X1 U967 ( .A1(KEYINPUT27), .A2(G107), .ZN(n1284) );
NAND2_X1 U968 ( .A1(G217), .A2(n1262), .ZN(n1283) );
AND2_X1 U969 ( .A1(G234), .A2(n1038), .ZN(n1262) );
OR2_X1 U970 ( .A1(n1056), .A2(n1285), .ZN(n1247) );
NOR2_X1 U971 ( .A1(n1047), .A2(n1048), .ZN(n1285) );
AND2_X1 U972 ( .A1(n1048), .A2(n1047), .ZN(n1056) );
INV_X1 U973 ( .A(G475), .ZN(n1047) );
NOR2_X1 U974 ( .A1(n1143), .A2(G902), .ZN(n1048) );
XNOR2_X1 U975 ( .A(n1286), .B(n1287), .ZN(n1143) );
XOR2_X1 U976 ( .A(n1288), .B(n1289), .Z(n1287) );
XOR2_X1 U977 ( .A(n1290), .B(n1291), .Z(n1289) );
NOR2_X1 U978 ( .A1(KEYINPUT50), .A2(n1109), .ZN(n1291) );
XNOR2_X1 U979 ( .A(G125), .B(G140), .ZN(n1109) );
AND2_X1 U980 ( .A1(n1292), .A2(G214), .ZN(n1290) );
XOR2_X1 U981 ( .A(G122), .B(G113), .Z(n1288) );
XOR2_X1 U982 ( .A(n1293), .B(n1294), .Z(n1286) );
XOR2_X1 U983 ( .A(n1295), .B(n1296), .Z(n1294) );
AND3_X1 U984 ( .A1(n1039), .A2(n1239), .A3(n1240), .ZN(n1213) );
AND2_X1 U985 ( .A1(n1220), .A2(n1297), .ZN(n1240) );
NAND2_X1 U986 ( .A1(n1094), .A2(n1298), .ZN(n1297) );
NAND4_X1 U987 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1122), .ZN(n1298) );
INV_X1 U988 ( .A(G898), .ZN(n1122) );
NAND3_X1 U989 ( .A1(n1243), .A2(n1038), .A3(G952), .ZN(n1094) );
NAND2_X1 U990 ( .A1(G234), .A2(G237), .ZN(n1243) );
INV_X1 U991 ( .A(n1091), .ZN(n1220) );
NAND2_X1 U992 ( .A1(n1237), .A2(n1238), .ZN(n1091) );
NAND2_X1 U993 ( .A1(n1055), .A2(n1059), .ZN(n1238) );
NAND3_X1 U994 ( .A1(n1299), .A2(n1191), .A3(n1300), .ZN(n1059) );
NAND2_X1 U995 ( .A1(G210), .A2(G237), .ZN(n1299) );
NAND3_X1 U996 ( .A1(n1301), .A2(n1302), .A3(G210), .ZN(n1055) );
NAND2_X1 U997 ( .A1(n1300), .A2(n1191), .ZN(n1301) );
XOR2_X1 U998 ( .A(n1303), .B(n1304), .Z(n1300) );
XOR2_X1 U999 ( .A(G125), .B(n1190), .Z(n1304) );
AND2_X1 U1000 ( .A1(G224), .A2(n1038), .ZN(n1190) );
XOR2_X1 U1001 ( .A(n1104), .B(n1305), .Z(n1303) );
NOR2_X1 U1002 ( .A1(KEYINPUT29), .A2(n1184), .ZN(n1305) );
XNOR2_X1 U1003 ( .A(n1124), .B(n1123), .ZN(n1184) );
XOR2_X1 U1004 ( .A(n1306), .B(G113), .Z(n1123) );
XOR2_X1 U1005 ( .A(n1307), .B(n1308), .Z(n1124) );
XNOR2_X1 U1006 ( .A(G101), .B(n1309), .ZN(n1308) );
NAND2_X1 U1007 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NAND2_X1 U1008 ( .A1(G107), .A2(n1293), .ZN(n1311) );
XOR2_X1 U1009 ( .A(n1312), .B(KEYINPUT2), .Z(n1310) );
OR2_X1 U1010 ( .A1(n1293), .A2(G107), .ZN(n1312) );
XOR2_X1 U1011 ( .A(n1173), .B(n1313), .Z(n1307) );
XOR2_X1 U1012 ( .A(KEYINPUT51), .B(G122), .Z(n1313) );
INV_X1 U1013 ( .A(G110), .ZN(n1173) );
XOR2_X1 U1014 ( .A(n1057), .B(KEYINPUT47), .Z(n1237) );
AND2_X1 U1015 ( .A1(G214), .A2(n1314), .ZN(n1057) );
XNOR2_X1 U1016 ( .A(KEYINPUT25), .B(n1302), .ZN(n1314) );
OR2_X1 U1017 ( .A1(G902), .A2(G237), .ZN(n1302) );
XOR2_X1 U1018 ( .A(n1071), .B(KEYINPUT56), .Z(n1239) );
INV_X1 U1019 ( .A(n1236), .ZN(n1071) );
NAND2_X1 U1020 ( .A1(n1250), .A2(n1040), .ZN(n1236) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1255), .ZN(n1040) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1191), .ZN(n1255) );
XOR2_X1 U1023 ( .A(n1049), .B(n1315), .Z(n1250) );
NOR2_X1 U1024 ( .A1(G469), .A2(KEYINPUT62), .ZN(n1315) );
NAND2_X1 U1025 ( .A1(n1316), .A2(n1191), .ZN(n1049) );
XOR2_X1 U1026 ( .A(n1317), .B(n1318), .Z(n1316) );
XNOR2_X1 U1027 ( .A(n1169), .B(n1319), .ZN(n1318) );
XOR2_X1 U1028 ( .A(KEYINPUT1), .B(G110), .Z(n1319) );
NAND2_X1 U1029 ( .A1(G227), .A2(n1038), .ZN(n1169) );
XOR2_X1 U1030 ( .A(n1320), .B(n1321), .Z(n1317) );
INV_X1 U1031 ( .A(n1179), .ZN(n1321) );
XOR2_X1 U1032 ( .A(n1322), .B(n1323), .Z(n1179) );
XOR2_X1 U1033 ( .A(G107), .B(G101), .Z(n1323) );
NAND2_X1 U1034 ( .A1(n1324), .A2(KEYINPUT14), .ZN(n1322) );
XOR2_X1 U1035 ( .A(n1293), .B(KEYINPUT52), .Z(n1324) );
XNOR2_X1 U1036 ( .A(G104), .B(KEYINPUT18), .ZN(n1293) );
XNOR2_X1 U1037 ( .A(n1155), .B(n1325), .ZN(n1320) );
NOR2_X1 U1038 ( .A1(G140), .A2(KEYINPUT63), .ZN(n1325) );
XOR2_X1 U1039 ( .A(n1326), .B(G472), .Z(n1039) );
NAND2_X1 U1040 ( .A1(n1327), .A2(n1191), .ZN(n1326) );
INV_X1 U1041 ( .A(G902), .ZN(n1191) );
XOR2_X1 U1042 ( .A(KEYINPUT7), .B(n1328), .Z(n1327) );
XOR2_X1 U1043 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1044 ( .A(n1331), .B(n1332), .Z(n1330) );
XNOR2_X1 U1045 ( .A(n1159), .B(n1333), .ZN(n1332) );
NOR2_X1 U1046 ( .A1(G101), .A2(KEYINPUT46), .ZN(n1333) );
NAND2_X1 U1047 ( .A1(G210), .A2(n1292), .ZN(n1159) );
AND2_X1 U1048 ( .A1(n1334), .A2(n1038), .ZN(n1292) );
INV_X1 U1049 ( .A(G953), .ZN(n1038) );
XNOR2_X1 U1050 ( .A(G237), .B(KEYINPUT8), .ZN(n1334) );
XNOR2_X1 U1051 ( .A(n1155), .B(n1154), .ZN(n1331) );
XNOR2_X1 U1052 ( .A(n1306), .B(n1335), .ZN(n1154) );
NOR2_X1 U1053 ( .A1(G113), .A2(KEYINPUT23), .ZN(n1335) );
XOR2_X1 U1054 ( .A(n1248), .B(n1258), .Z(n1306) );
XOR2_X1 U1055 ( .A(G119), .B(KEYINPUT13), .Z(n1258) );
INV_X1 U1056 ( .A(G116), .ZN(n1248) );
XOR2_X1 U1057 ( .A(n1175), .B(n1107), .Z(n1155) );
INV_X1 U1058 ( .A(n1104), .ZN(n1107) );
XNOR2_X1 U1059 ( .A(G128), .B(n1295), .ZN(n1104) );
XOR2_X1 U1060 ( .A(G146), .B(G143), .Z(n1295) );
XNOR2_X1 U1061 ( .A(n1336), .B(KEYINPUT3), .ZN(n1175) );
NAND3_X1 U1062 ( .A1(n1337), .A2(n1338), .A3(n1111), .ZN(n1336) );
NAND3_X1 U1063 ( .A1(n1339), .A2(n1229), .A3(G134), .ZN(n1111) );
NAND2_X1 U1064 ( .A1(n1340), .A2(n1341), .ZN(n1338) );
INV_X1 U1065 ( .A(KEYINPUT58), .ZN(n1341) );
XOR2_X1 U1066 ( .A(n1342), .B(n1296), .Z(n1340) );
NAND2_X1 U1067 ( .A1(G137), .A2(n1343), .ZN(n1342) );
NAND2_X1 U1068 ( .A1(KEYINPUT58), .A2(n1112), .ZN(n1337) );
NAND2_X1 U1069 ( .A1(n1344), .A2(n1345), .ZN(n1112) );
NAND2_X1 U1070 ( .A1(n1346), .A2(G137), .ZN(n1345) );
XOR2_X1 U1071 ( .A(n1343), .B(n1296), .Z(n1346) );
NAND3_X1 U1072 ( .A1(n1296), .A2(n1343), .A3(n1229), .ZN(n1344) );
INV_X1 U1073 ( .A(G137), .ZN(n1229) );
INV_X1 U1074 ( .A(G134), .ZN(n1343) );
INV_X1 U1075 ( .A(n1339), .ZN(n1296) );
XNOR2_X1 U1076 ( .A(G131), .B(KEYINPUT19), .ZN(n1339) );
XOR2_X1 U1077 ( .A(n1347), .B(n1348), .Z(n1329) );
XOR2_X1 U1078 ( .A(KEYINPUT53), .B(KEYINPUT49), .Z(n1348) );
XNOR2_X1 U1079 ( .A(KEYINPUT41), .B(KEYINPUT32), .ZN(n1347) );
endmodule


