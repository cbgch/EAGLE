//Key = 0100111001001000000010101101110010111011000000010111100100000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343;

XNOR2_X1 U734 ( .A(n1020), .B(n1021), .ZN(G9) );
NAND2_X1 U735 ( .A1(KEYINPUT27), .A2(n1022), .ZN(n1020) );
NOR2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(G75) );
NOR4_X1 U737 ( .A1(n1025), .A2(n1026), .A3(G953), .A4(n1027), .ZN(n1024) );
NOR3_X1 U738 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1026) );
NOR4_X1 U739 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1029) );
INV_X1 U740 ( .A(n1035), .ZN(n1033) );
NAND2_X1 U741 ( .A1(n1036), .A2(n1037), .ZN(n1031) );
NAND2_X1 U742 ( .A1(n1038), .A2(n1039), .ZN(n1025) );
NAND2_X1 U743 ( .A1(n1037), .A2(n1040), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND3_X1 U745 ( .A1(n1035), .A2(n1043), .A3(n1044), .ZN(n1042) );
NAND2_X1 U746 ( .A1(n1045), .A2(n1046), .ZN(n1043) );
NAND2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U748 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND3_X1 U749 ( .A1(n1051), .A2(n1028), .A3(n1036), .ZN(n1050) );
INV_X1 U750 ( .A(KEYINPUT15), .ZN(n1028) );
NAND2_X1 U751 ( .A1(n1052), .A2(n1053), .ZN(n1045) );
NAND2_X1 U752 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U753 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NAND3_X1 U754 ( .A1(n1052), .A2(n1058), .A3(n1047), .ZN(n1041) );
INV_X1 U755 ( .A(n1030), .ZN(n1047) );
NAND3_X1 U756 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NAND2_X1 U757 ( .A1(n1035), .A2(n1062), .ZN(n1061) );
OR2_X1 U758 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND2_X1 U759 ( .A1(n1044), .A2(n1065), .ZN(n1060) );
NAND2_X1 U760 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
INV_X1 U762 ( .A(KEYINPUT3), .ZN(n1069) );
INV_X1 U763 ( .A(n1070), .ZN(n1066) );
NAND3_X1 U764 ( .A1(KEYINPUT3), .A2(n1068), .A3(n1032), .ZN(n1059) );
INV_X1 U765 ( .A(n1071), .ZN(n1037) );
NOR3_X1 U766 ( .A1(n1027), .A2(G953), .A3(G952), .ZN(n1023) );
AND4_X1 U767 ( .A1(n1052), .A2(n1035), .A3(n1072), .A4(n1073), .ZN(n1027) );
NOR4_X1 U768 ( .A1(n1074), .A2(n1056), .A3(n1075), .A4(n1076), .ZN(n1073) );
NOR2_X1 U769 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U770 ( .A1(G902), .A2(n1079), .ZN(n1077) );
NOR3_X1 U771 ( .A1(n1080), .A2(KEYINPUT40), .A3(n1081), .ZN(n1075) );
INV_X1 U772 ( .A(n1082), .ZN(n1081) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1072) );
AND2_X1 U774 ( .A1(n1085), .A2(G475), .ZN(n1084) );
NOR2_X1 U775 ( .A1(G902), .A2(n1086), .ZN(n1083) );
NOR2_X1 U776 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U777 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
XNOR2_X1 U778 ( .A(n1091), .B(n1092), .ZN(n1090) );
NOR2_X1 U779 ( .A1(KEYINPUT40), .A2(n1080), .ZN(n1089) );
NOR2_X1 U780 ( .A1(G475), .A2(n1093), .ZN(n1087) );
XOR2_X1 U781 ( .A(n1094), .B(n1095), .Z(G72) );
NOR2_X1 U782 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NOR2_X1 U783 ( .A1(n1098), .A2(n1099), .ZN(n1096) );
NAND2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1094) );
OR2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND3_X1 U786 ( .A1(n1104), .A2(n1102), .A3(n1103), .ZN(n1100) );
XNOR2_X1 U787 ( .A(n1105), .B(n1106), .ZN(n1103) );
XOR2_X1 U788 ( .A(n1107), .B(n1108), .Z(n1105) );
NAND2_X1 U789 ( .A1(KEYINPUT1), .A2(n1109), .ZN(n1107) );
NAND2_X1 U790 ( .A1(n1097), .A2(n1110), .ZN(n1102) );
NAND4_X1 U791 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1110) );
NOR2_X1 U792 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U793 ( .A(n1117), .B(KEYINPUT52), .Z(n1115) );
NAND2_X1 U794 ( .A1(G953), .A2(n1099), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1118), .B(n1119), .Z(G69) );
XOR2_X1 U796 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U797 ( .A1(n1122), .A2(G953), .ZN(n1121) );
NOR2_X1 U798 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
XNOR2_X1 U799 ( .A(KEYINPUT13), .B(n1125), .ZN(n1124) );
NAND2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1120) );
NAND2_X1 U801 ( .A1(G953), .A2(n1128), .ZN(n1127) );
XNOR2_X1 U802 ( .A(n1129), .B(n1130), .ZN(n1126) );
NOR2_X1 U803 ( .A1(KEYINPUT33), .A2(n1131), .ZN(n1130) );
XNOR2_X1 U804 ( .A(n1132), .B(n1133), .ZN(n1131) );
NOR2_X1 U805 ( .A1(KEYINPUT56), .A2(n1134), .ZN(n1132) );
NAND2_X1 U806 ( .A1(G953), .A2(n1135), .ZN(n1118) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1135) );
NOR3_X1 U808 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(G66) );
AND2_X1 U809 ( .A1(KEYINPUT12), .A2(n1139), .ZN(n1138) );
NOR3_X1 U810 ( .A1(KEYINPUT12), .A2(G953), .A3(G952), .ZN(n1137) );
XOR2_X1 U811 ( .A(n1140), .B(n1141), .Z(n1136) );
NAND2_X1 U812 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NOR2_X1 U813 ( .A1(n1144), .A2(n1145), .ZN(G63) );
XNOR2_X1 U814 ( .A(n1146), .B(n1079), .ZN(n1145) );
NAND2_X1 U815 ( .A1(n1142), .A2(G478), .ZN(n1146) );
NOR2_X1 U816 ( .A1(n1147), .A2(n1097), .ZN(n1144) );
XNOR2_X1 U817 ( .A(G952), .B(KEYINPUT55), .ZN(n1147) );
NOR3_X1 U818 ( .A1(n1148), .A2(n1139), .A3(n1149), .ZN(G60) );
NOR4_X1 U819 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1149) );
NOR2_X1 U820 ( .A1(KEYINPUT14), .A2(n1154), .ZN(n1151) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1093), .ZN(n1150) );
NOR2_X1 U822 ( .A1(KEYINPUT14), .A2(n1156), .ZN(n1155) );
NOR2_X1 U823 ( .A1(n1157), .A2(n1158), .ZN(n1148) );
NOR2_X1 U824 ( .A1(n1093), .A2(n1156), .ZN(n1158) );
INV_X1 U825 ( .A(KEYINPUT62), .ZN(n1156) );
INV_X1 U826 ( .A(n1154), .ZN(n1093) );
NOR2_X1 U827 ( .A1(n1152), .A2(n1153), .ZN(n1157) );
XOR2_X1 U828 ( .A(G104), .B(n1159), .Z(G6) );
NOR2_X1 U829 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U830 ( .A(KEYINPUT18), .B(KEYINPUT10), .Z(n1161) );
NOR2_X1 U831 ( .A1(n1139), .A2(n1162), .ZN(G57) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1162) );
XNOR2_X1 U833 ( .A(n1165), .B(n1166), .ZN(n1164) );
NAND2_X1 U834 ( .A1(KEYINPUT39), .A2(n1167), .ZN(n1165) );
XOR2_X1 U835 ( .A(n1168), .B(n1169), .Z(n1163) );
XNOR2_X1 U836 ( .A(G101), .B(n1170), .ZN(n1169) );
NAND2_X1 U837 ( .A1(n1142), .A2(G472), .ZN(n1170) );
NAND2_X1 U838 ( .A1(KEYINPUT29), .A2(n1133), .ZN(n1168) );
NOR2_X1 U839 ( .A1(n1139), .A2(n1171), .ZN(G54) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1171) );
XNOR2_X1 U841 ( .A(n1174), .B(n1134), .ZN(n1173) );
XNOR2_X1 U842 ( .A(n1175), .B(n1176), .ZN(n1174) );
XOR2_X1 U843 ( .A(n1177), .B(n1178), .Z(n1172) );
NOR2_X1 U844 ( .A1(n1179), .A2(KEYINPUT44), .ZN(n1178) );
XNOR2_X1 U845 ( .A(KEYINPUT46), .B(n1180), .ZN(n1177) );
NOR3_X1 U846 ( .A1(n1153), .A2(KEYINPUT21), .A3(n1181), .ZN(n1180) );
NOR2_X1 U847 ( .A1(n1139), .A2(n1182), .ZN(G51) );
XNOR2_X1 U848 ( .A(n1092), .B(n1183), .ZN(n1182) );
XOR2_X1 U849 ( .A(n1184), .B(n1185), .Z(n1183) );
NAND2_X1 U850 ( .A1(KEYINPUT6), .A2(n1091), .ZN(n1185) );
OR2_X1 U851 ( .A1(n1153), .A2(n1080), .ZN(n1184) );
INV_X1 U852 ( .A(n1142), .ZN(n1153) );
NOR2_X1 U853 ( .A1(n1186), .A2(n1038), .ZN(n1142) );
NOR4_X1 U854 ( .A1(n1123), .A2(n1116), .A3(n1187), .A4(n1188), .ZN(n1038) );
NAND4_X1 U855 ( .A1(n1125), .A2(n1112), .A3(n1111), .A4(n1117), .ZN(n1188) );
NAND3_X1 U856 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1117) );
XNOR2_X1 U857 ( .A(KEYINPUT42), .B(n1032), .ZN(n1189) );
INV_X1 U858 ( .A(n1044), .ZN(n1032) );
XNOR2_X1 U859 ( .A(n1113), .B(KEYINPUT60), .ZN(n1187) );
NAND2_X1 U860 ( .A1(n1192), .A2(n1193), .ZN(n1113) );
XOR2_X1 U861 ( .A(KEYINPUT8), .B(n1194), .Z(n1193) );
NOR2_X1 U862 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
NAND4_X1 U863 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1116) );
NAND3_X1 U864 ( .A1(n1063), .A2(n1070), .A3(n1191), .ZN(n1198) );
NAND2_X1 U865 ( .A1(n1201), .A2(n1192), .ZN(n1197) );
XOR2_X1 U866 ( .A(n1202), .B(KEYINPUT24), .Z(n1201) );
NAND4_X1 U867 ( .A1(n1160), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1123) );
AND4_X1 U868 ( .A1(n1021), .A2(n1206), .A3(n1207), .A4(n1208), .ZN(n1205) );
NAND3_X1 U869 ( .A1(n1064), .A2(n1035), .A3(n1209), .ZN(n1021) );
NAND4_X1 U870 ( .A1(n1210), .A2(n1211), .A3(n1052), .A4(n1212), .ZN(n1204) );
XNOR2_X1 U871 ( .A(n1192), .B(KEYINPUT61), .ZN(n1210) );
NAND3_X1 U872 ( .A1(n1209), .A2(n1035), .A3(n1063), .ZN(n1160) );
NOR2_X1 U873 ( .A1(n1097), .A2(G952), .ZN(n1139) );
XNOR2_X1 U874 ( .A(G146), .B(n1213), .ZN(G48) );
NAND3_X1 U875 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1213) );
NOR3_X1 U876 ( .A1(n1054), .A2(KEYINPUT53), .A3(n1049), .ZN(n1216) );
INV_X1 U877 ( .A(n1217), .ZN(n1049) );
INV_X1 U878 ( .A(n1196), .ZN(n1215) );
NAND2_X1 U879 ( .A1(n1063), .A2(n1190), .ZN(n1196) );
XOR2_X1 U880 ( .A(n1218), .B(KEYINPUT23), .Z(n1214) );
XNOR2_X1 U881 ( .A(G143), .B(n1111), .ZN(G45) );
NAND4_X1 U882 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1070), .ZN(n1111) );
NOR2_X1 U883 ( .A1(n1222), .A2(n1054), .ZN(n1221) );
XNOR2_X1 U884 ( .A(n1223), .B(n1112), .ZN(G42) );
NAND3_X1 U885 ( .A1(n1063), .A2(n1068), .A3(n1191), .ZN(n1112) );
NOR2_X1 U886 ( .A1(KEYINPUT16), .A2(n1224), .ZN(n1223) );
XOR2_X1 U887 ( .A(KEYINPUT25), .B(G140), .Z(n1224) );
XNOR2_X1 U888 ( .A(G137), .B(n1225), .ZN(G39) );
NAND2_X1 U889 ( .A1(n1191), .A2(n1211), .ZN(n1225) );
XNOR2_X1 U890 ( .A(G134), .B(n1199), .ZN(G36) );
NAND3_X1 U891 ( .A1(n1070), .A2(n1064), .A3(n1191), .ZN(n1199) );
XNOR2_X1 U892 ( .A(G131), .B(n1226), .ZN(G33) );
NAND4_X1 U893 ( .A1(n1063), .A2(n1070), .A3(n1227), .A4(n1228), .ZN(n1226) );
OR2_X1 U894 ( .A1(n1191), .A2(KEYINPUT41), .ZN(n1228) );
NOR2_X1 U895 ( .A1(n1195), .A2(n1030), .ZN(n1191) );
NAND2_X1 U896 ( .A1(KEYINPUT41), .A2(n1229), .ZN(n1227) );
NAND2_X1 U897 ( .A1(n1219), .A2(n1030), .ZN(n1229) );
NAND2_X1 U898 ( .A1(n1057), .A2(n1230), .ZN(n1030) );
XNOR2_X1 U899 ( .A(n1231), .B(n1232), .ZN(G30) );
NOR2_X1 U900 ( .A1(n1233), .A2(n1054), .ZN(n1232) );
INV_X1 U901 ( .A(n1192), .ZN(n1054) );
XOR2_X1 U902 ( .A(n1202), .B(KEYINPUT7), .Z(n1233) );
NAND3_X1 U903 ( .A1(n1064), .A2(n1190), .A3(n1219), .ZN(n1202) );
INV_X1 U904 ( .A(n1195), .ZN(n1219) );
NAND2_X1 U905 ( .A1(n1217), .A2(n1218), .ZN(n1195) );
NAND3_X1 U906 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(G3) );
NAND2_X1 U907 ( .A1(KEYINPUT30), .A2(n1237), .ZN(n1236) );
NAND3_X1 U908 ( .A1(n1238), .A2(n1239), .A3(n1203), .ZN(n1235) );
NAND2_X1 U909 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
NAND2_X1 U910 ( .A1(n1242), .A2(n1239), .ZN(n1241) );
INV_X1 U911 ( .A(KEYINPUT30), .ZN(n1239) );
XNOR2_X1 U912 ( .A(n1238), .B(n1243), .ZN(n1242) );
XOR2_X1 U913 ( .A(KEYINPUT45), .B(KEYINPUT36), .Z(n1243) );
INV_X1 U914 ( .A(n1237), .ZN(n1238) );
XOR2_X1 U915 ( .A(G101), .B(KEYINPUT35), .Z(n1237) );
INV_X1 U916 ( .A(n1203), .ZN(n1240) );
NAND3_X1 U917 ( .A1(n1044), .A2(n1209), .A3(n1070), .ZN(n1203) );
XNOR2_X1 U918 ( .A(G125), .B(n1200), .ZN(G27) );
NAND3_X1 U919 ( .A1(n1063), .A2(n1068), .A3(n1244), .ZN(n1200) );
AND3_X1 U920 ( .A1(n1052), .A2(n1218), .A3(n1192), .ZN(n1244) );
NAND2_X1 U921 ( .A1(n1245), .A2(n1071), .ZN(n1218) );
NAND4_X1 U922 ( .A1(G902), .A2(G953), .A3(n1246), .A4(n1099), .ZN(n1245) );
INV_X1 U923 ( .A(G900), .ZN(n1099) );
XNOR2_X1 U924 ( .A(G122), .B(n1208), .ZN(G24) );
NAND4_X1 U925 ( .A1(n1220), .A2(n1247), .A3(n1035), .A4(n1248), .ZN(n1208) );
NOR2_X1 U926 ( .A1(n1249), .A2(n1250), .ZN(n1035) );
XNOR2_X1 U927 ( .A(G119), .B(n1251), .ZN(G21) );
NAND2_X1 U928 ( .A1(n1211), .A2(n1247), .ZN(n1251) );
AND2_X1 U929 ( .A1(n1044), .A2(n1190), .ZN(n1211) );
NAND2_X1 U930 ( .A1(n1252), .A2(n1253), .ZN(n1190) );
NAND3_X1 U931 ( .A1(n1250), .A2(n1249), .A3(n1254), .ZN(n1253) );
INV_X1 U932 ( .A(KEYINPUT31), .ZN(n1254) );
NAND2_X1 U933 ( .A1(KEYINPUT31), .A2(n1070), .ZN(n1252) );
NAND2_X1 U934 ( .A1(n1255), .A2(n1256), .ZN(G18) );
NAND2_X1 U935 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U936 ( .A(KEYINPUT0), .B(n1207), .ZN(n1257) );
NAND2_X1 U937 ( .A1(G116), .A2(n1259), .ZN(n1255) );
XOR2_X1 U938 ( .A(n1207), .B(KEYINPUT63), .Z(n1259) );
NAND3_X1 U939 ( .A1(n1247), .A2(n1064), .A3(n1070), .ZN(n1207) );
NOR2_X1 U940 ( .A1(n1220), .A2(n1222), .ZN(n1064) );
XNOR2_X1 U941 ( .A(G113), .B(n1125), .ZN(G15) );
NAND3_X1 U942 ( .A1(n1070), .A2(n1247), .A3(n1063), .ZN(n1125) );
NOR2_X1 U943 ( .A1(n1260), .A2(n1248), .ZN(n1063) );
AND3_X1 U944 ( .A1(n1192), .A2(n1212), .A3(n1052), .ZN(n1247) );
NOR2_X1 U945 ( .A1(n1034), .A2(n1036), .ZN(n1052) );
NOR2_X1 U946 ( .A1(n1250), .A2(n1261), .ZN(n1070) );
XNOR2_X1 U947 ( .A(G110), .B(n1206), .ZN(G12) );
NAND3_X1 U948 ( .A1(n1068), .A2(n1209), .A3(n1044), .ZN(n1206) );
NOR2_X1 U949 ( .A1(n1248), .A2(n1220), .ZN(n1044) );
INV_X1 U950 ( .A(n1260), .ZN(n1220) );
NAND3_X1 U951 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1260) );
OR2_X1 U952 ( .A1(n1152), .A2(KEYINPUT32), .ZN(n1264) );
INV_X1 U953 ( .A(G475), .ZN(n1152) );
NAND3_X1 U954 ( .A1(KEYINPUT32), .A2(n1265), .A3(n1085), .ZN(n1263) );
OR2_X1 U955 ( .A1(n1085), .A2(n1265), .ZN(n1262) );
NOR2_X1 U956 ( .A1(G475), .A2(KEYINPUT26), .ZN(n1265) );
NAND2_X1 U957 ( .A1(n1154), .A2(n1186), .ZN(n1085) );
XNOR2_X1 U958 ( .A(n1266), .B(n1267), .ZN(n1154) );
XOR2_X1 U959 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U960 ( .A(n1270), .B(G104), .Z(n1269) );
NAND2_X1 U961 ( .A1(KEYINPUT34), .A2(n1271), .ZN(n1270) );
XOR2_X1 U962 ( .A(n1106), .B(n1272), .Z(n1271) );
XNOR2_X1 U963 ( .A(n1273), .B(KEYINPUT11), .ZN(n1272) );
NAND2_X1 U964 ( .A1(KEYINPUT50), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U965 ( .A(n1275), .B(G140), .ZN(n1106) );
XNOR2_X1 U966 ( .A(G113), .B(G143), .ZN(n1268) );
XOR2_X1 U967 ( .A(n1276), .B(n1277), .Z(n1266) );
XNOR2_X1 U968 ( .A(n1278), .B(n1279), .ZN(n1277) );
NOR2_X1 U969 ( .A1(G131), .A2(KEYINPUT19), .ZN(n1279) );
NAND2_X1 U970 ( .A1(KEYINPUT47), .A2(n1280), .ZN(n1278) );
NAND2_X1 U971 ( .A1(KEYINPUT20), .A2(n1281), .ZN(n1276) );
NAND3_X1 U972 ( .A1(G214), .A2(n1097), .A3(n1282), .ZN(n1281) );
XNOR2_X1 U973 ( .A(G237), .B(KEYINPUT43), .ZN(n1282) );
INV_X1 U974 ( .A(n1222), .ZN(n1248) );
NOR2_X1 U975 ( .A1(n1283), .A2(n1074), .ZN(n1222) );
NOR3_X1 U976 ( .A1(n1284), .A2(G902), .A3(n1079), .ZN(n1074) );
AND2_X1 U977 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
NAND2_X1 U978 ( .A1(n1287), .A2(n1186), .ZN(n1286) );
INV_X1 U979 ( .A(n1079), .ZN(n1287) );
XNOR2_X1 U980 ( .A(n1288), .B(n1289), .ZN(n1079) );
XOR2_X1 U981 ( .A(n1290), .B(n1291), .Z(n1289) );
XNOR2_X1 U982 ( .A(n1022), .B(n1292), .ZN(n1291) );
NOR2_X1 U983 ( .A1(KEYINPUT57), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U984 ( .A(n1231), .B(n1294), .ZN(n1293) );
XNOR2_X1 U985 ( .A(n1295), .B(G134), .ZN(n1294) );
INV_X1 U986 ( .A(G143), .ZN(n1295) );
INV_X1 U987 ( .A(G128), .ZN(n1231) );
AND2_X1 U988 ( .A1(n1296), .A2(G217), .ZN(n1290) );
XNOR2_X1 U989 ( .A(G116), .B(n1297), .ZN(n1288) );
XNOR2_X1 U990 ( .A(KEYINPUT17), .B(n1280), .ZN(n1297) );
XNOR2_X1 U991 ( .A(KEYINPUT54), .B(n1078), .ZN(n1285) );
INV_X1 U992 ( .A(n1284), .ZN(n1078) );
XOR2_X1 U993 ( .A(G478), .B(KEYINPUT48), .Z(n1284) );
AND3_X1 U994 ( .A1(n1217), .A2(n1212), .A3(n1192), .ZN(n1209) );
NOR2_X1 U995 ( .A1(n1057), .A2(n1056), .ZN(n1192) );
INV_X1 U996 ( .A(n1230), .ZN(n1056) );
NAND2_X1 U997 ( .A1(G214), .A2(n1298), .ZN(n1230) );
XOR2_X1 U998 ( .A(n1299), .B(n1300), .Z(n1057) );
XNOR2_X1 U999 ( .A(KEYINPUT51), .B(n1080), .ZN(n1300) );
NAND2_X1 U1000 ( .A1(G210), .A2(n1298), .ZN(n1080) );
NAND2_X1 U1001 ( .A1(n1301), .A2(n1186), .ZN(n1298) );
NAND2_X1 U1002 ( .A1(KEYINPUT38), .A2(n1082), .ZN(n1299) );
NAND2_X1 U1003 ( .A1(n1302), .A2(n1186), .ZN(n1082) );
XOR2_X1 U1004 ( .A(n1091), .B(n1092), .Z(n1302) );
XNOR2_X1 U1005 ( .A(n1303), .B(n1304), .ZN(n1092) );
XNOR2_X1 U1006 ( .A(KEYINPUT59), .B(n1275), .ZN(n1304) );
INV_X1 U1007 ( .A(G125), .ZN(n1275) );
XOR2_X1 U1008 ( .A(n1305), .B(n1306), .Z(n1303) );
NOR2_X1 U1009 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
INV_X1 U1010 ( .A(G224), .ZN(n1308) );
XNOR2_X1 U1011 ( .A(G953), .B(KEYINPUT22), .ZN(n1307) );
XNOR2_X1 U1012 ( .A(n1309), .B(n1310), .ZN(n1091) );
INV_X1 U1013 ( .A(n1129), .ZN(n1310) );
XOR2_X1 U1014 ( .A(G110), .B(n1311), .Z(n1129) );
XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n1280), .ZN(n1311) );
INV_X1 U1016 ( .A(G122), .ZN(n1280) );
NAND2_X1 U1017 ( .A1(n1312), .A2(n1313), .ZN(n1309) );
NAND2_X1 U1018 ( .A1(n1134), .A2(n1133), .ZN(n1313) );
XOR2_X1 U1019 ( .A(KEYINPUT28), .B(n1314), .Z(n1312) );
NOR2_X1 U1020 ( .A1(n1134), .A2(n1133), .ZN(n1314) );
NAND2_X1 U1021 ( .A1(n1071), .A2(n1315), .ZN(n1212) );
NAND4_X1 U1022 ( .A1(G902), .A2(G953), .A3(n1246), .A4(n1128), .ZN(n1315) );
INV_X1 U1023 ( .A(G898), .ZN(n1128) );
NAND3_X1 U1024 ( .A1(n1246), .A2(n1097), .A3(n1316), .ZN(n1071) );
XNOR2_X1 U1025 ( .A(G952), .B(KEYINPUT4), .ZN(n1316) );
NAND2_X1 U1026 ( .A1(G237), .A2(G234), .ZN(n1246) );
NOR2_X1 U1027 ( .A1(n1051), .A2(n1036), .ZN(n1217) );
AND2_X1 U1028 ( .A1(G221), .A2(n1317), .ZN(n1036) );
INV_X1 U1029 ( .A(n1034), .ZN(n1051) );
XOR2_X1 U1030 ( .A(n1318), .B(n1181), .Z(n1034) );
INV_X1 U1031 ( .A(G469), .ZN(n1181) );
NAND2_X1 U1032 ( .A1(n1319), .A2(n1186), .ZN(n1318) );
XOR2_X1 U1033 ( .A(n1320), .B(n1321), .Z(n1319) );
XOR2_X1 U1034 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1035 ( .A(n1179), .B(n1324), .ZN(n1323) );
NOR2_X1 U1036 ( .A1(KEYINPUT58), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1037 ( .A(G131), .B(n1326), .ZN(n1325) );
NOR2_X1 U1038 ( .A1(n1098), .A2(G953), .ZN(n1179) );
INV_X1 U1039 ( .A(G227), .ZN(n1098) );
XNOR2_X1 U1040 ( .A(G140), .B(KEYINPUT37), .ZN(n1322) );
XNOR2_X1 U1041 ( .A(n1327), .B(n1134), .ZN(n1320) );
XNOR2_X1 U1042 ( .A(G101), .B(n1328), .ZN(n1134) );
XNOR2_X1 U1043 ( .A(n1022), .B(G104), .ZN(n1328) );
INV_X1 U1044 ( .A(G107), .ZN(n1022) );
XOR2_X1 U1045 ( .A(n1305), .B(n1329), .Z(n1327) );
NOR2_X1 U1046 ( .A1(G110), .A2(KEYINPUT2), .ZN(n1329) );
AND2_X1 U1047 ( .A1(n1261), .A2(n1250), .ZN(n1068) );
XNOR2_X1 U1048 ( .A(n1330), .B(n1143), .ZN(n1250) );
AND2_X1 U1049 ( .A1(G217), .A2(n1317), .ZN(n1143) );
NAND2_X1 U1050 ( .A1(G234), .A2(n1186), .ZN(n1317) );
NAND2_X1 U1051 ( .A1(n1141), .A2(n1186), .ZN(n1330) );
XNOR2_X1 U1052 ( .A(n1331), .B(n1332), .ZN(n1141) );
XOR2_X1 U1053 ( .A(n1333), .B(n1334), .Z(n1332) );
XNOR2_X1 U1054 ( .A(G119), .B(G125), .ZN(n1334) );
NAND2_X1 U1055 ( .A1(KEYINPUT9), .A2(n1335), .ZN(n1333) );
XNOR2_X1 U1056 ( .A(G137), .B(n1336), .ZN(n1335) );
NAND2_X1 U1057 ( .A1(n1296), .A2(G221), .ZN(n1336) );
AND2_X1 U1058 ( .A1(G234), .A2(n1097), .ZN(n1296) );
XNOR2_X1 U1059 ( .A(n1337), .B(n1176), .ZN(n1331) );
XOR2_X1 U1060 ( .A(G110), .B(G140), .Z(n1176) );
INV_X1 U1061 ( .A(n1249), .ZN(n1261) );
XNOR2_X1 U1062 ( .A(n1338), .B(G472), .ZN(n1249) );
NAND2_X1 U1063 ( .A1(n1339), .A2(n1186), .ZN(n1338) );
INV_X1 U1064 ( .A(G902), .ZN(n1186) );
XNOR2_X1 U1065 ( .A(n1340), .B(n1133), .ZN(n1339) );
XNOR2_X1 U1066 ( .A(G113), .B(n1341), .ZN(n1133) );
XNOR2_X1 U1067 ( .A(G119), .B(n1258), .ZN(n1341) );
INV_X1 U1068 ( .A(G116), .ZN(n1258) );
XOR2_X1 U1069 ( .A(n1342), .B(n1166), .Z(n1340) );
XOR2_X1 U1070 ( .A(KEYINPUT59), .B(n1175), .Z(n1166) );
XNOR2_X1 U1071 ( .A(n1108), .B(n1109), .ZN(n1175) );
INV_X1 U1072 ( .A(G131), .ZN(n1109) );
XNOR2_X1 U1073 ( .A(n1305), .B(n1326), .ZN(n1108) );
XOR2_X1 U1074 ( .A(G134), .B(G137), .Z(n1326) );
XNOR2_X1 U1075 ( .A(G143), .B(n1337), .ZN(n1305) );
XNOR2_X1 U1076 ( .A(G128), .B(n1274), .ZN(n1337) );
INV_X1 U1077 ( .A(G146), .ZN(n1274) );
NAND2_X1 U1078 ( .A1(n1343), .A2(KEYINPUT5), .ZN(n1342) );
XOR2_X1 U1079 ( .A(n1167), .B(G101), .Z(n1343) );
NAND3_X1 U1080 ( .A1(n1301), .A2(n1097), .A3(G210), .ZN(n1167) );
INV_X1 U1081 ( .A(G953), .ZN(n1097) );
INV_X1 U1082 ( .A(G237), .ZN(n1301) );
endmodule


