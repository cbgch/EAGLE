//Key = 0111101011101011111100101010111010011100010011011010001100011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
n1416, n1417, n1418, n1419;

XOR2_X1 U766 ( .A(n1066), .B(n1067), .Z(G9) );
NOR2_X1 U767 ( .A1(G107), .A2(KEYINPUT40), .ZN(n1067) );
OR2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR2_X1 U769 ( .A1(n1070), .A2(n1071), .ZN(G75) );
XOR2_X1 U770 ( .A(KEYINPUT31), .B(n1072), .Z(n1071) );
AND3_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1072) );
NOR3_X1 U772 ( .A1(n1076), .A2(n1075), .A3(n1077), .ZN(n1070) );
NAND3_X1 U773 ( .A1(n1073), .A2(n1074), .A3(n1078), .ZN(n1076) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U776 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NAND3_X1 U777 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1084) );
NAND2_X1 U778 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1087) );
XNOR2_X1 U780 ( .A(n1089), .B(KEYINPUT28), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1093), .A2(n1094), .ZN(n1086) );
NAND2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U783 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND3_X1 U784 ( .A1(n1093), .A2(n1099), .A3(n1089), .ZN(n1081) );
NAND3_X1 U785 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
NAND2_X1 U786 ( .A1(n1103), .A2(n1083), .ZN(n1102) );
NAND3_X1 U787 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1101) );
XOR2_X1 U788 ( .A(KEYINPUT49), .B(n1083), .Z(n1105) );
NAND2_X1 U789 ( .A1(n1085), .A2(n1107), .ZN(n1100) );
NAND2_X1 U790 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND4_X1 U791 ( .A1(n1110), .A2(n1085), .A3(n1111), .A4(n1112), .ZN(n1073) );
NOR4_X1 U792 ( .A1(n1097), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1112) );
XNOR2_X1 U793 ( .A(n1116), .B(n1117), .ZN(n1115) );
NAND2_X1 U794 ( .A1(KEYINPUT8), .A2(n1118), .ZN(n1116) );
INV_X1 U795 ( .A(n1119), .ZN(n1118) );
XNOR2_X1 U796 ( .A(n1120), .B(n1121), .ZN(n1114) );
NAND2_X1 U797 ( .A1(KEYINPUT22), .A2(n1122), .ZN(n1120) );
NOR2_X1 U798 ( .A1(n1123), .A2(n1124), .ZN(n1113) );
NOR2_X1 U799 ( .A1(n1125), .A2(n1126), .ZN(n1111) );
XOR2_X1 U800 ( .A(n1127), .B(KEYINPUT6), .Z(n1126) );
XOR2_X1 U801 ( .A(n1128), .B(n1129), .Z(n1125) );
XOR2_X1 U802 ( .A(KEYINPUT14), .B(G472), .Z(n1129) );
XOR2_X1 U803 ( .A(n1130), .B(KEYINPUT7), .Z(n1110) );
XOR2_X1 U804 ( .A(n1131), .B(n1132), .Z(G72) );
XOR2_X1 U805 ( .A(n1133), .B(n1134), .Z(n1132) );
NOR2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U807 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U808 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U809 ( .A1(n1141), .A2(n1142), .ZN(n1139) );
NAND3_X1 U810 ( .A1(G131), .A2(n1143), .A3(n1144), .ZN(n1142) );
INV_X1 U811 ( .A(KEYINPUT54), .ZN(n1144) );
NAND2_X1 U812 ( .A1(KEYINPUT54), .A2(n1145), .ZN(n1141) );
XNOR2_X1 U813 ( .A(G140), .B(n1146), .ZN(n1137) );
NOR2_X1 U814 ( .A1(G900), .A2(n1147), .ZN(n1135) );
XNOR2_X1 U815 ( .A(G953), .B(KEYINPUT52), .ZN(n1147) );
NOR2_X1 U816 ( .A1(KEYINPUT58), .A2(n1148), .ZN(n1133) );
NOR2_X1 U817 ( .A1(n1149), .A2(G953), .ZN(n1148) );
NAND2_X1 U818 ( .A1(G953), .A2(n1150), .ZN(n1131) );
NAND2_X1 U819 ( .A1(G900), .A2(G227), .ZN(n1150) );
XOR2_X1 U820 ( .A(n1151), .B(n1152), .Z(G69) );
XOR2_X1 U821 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U822 ( .A1(G953), .A2(n1155), .ZN(n1154) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1155) );
NAND2_X1 U824 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
NAND2_X1 U825 ( .A1(G953), .A2(n1158), .ZN(n1157) );
XOR2_X1 U826 ( .A(n1159), .B(n1160), .Z(n1156) );
NAND2_X1 U827 ( .A1(KEYINPUT10), .A2(n1161), .ZN(n1159) );
NOR2_X1 U828 ( .A1(n1162), .A2(G953), .ZN(n1151) );
NOR2_X1 U829 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1165), .A2(n1166), .ZN(G66) );
XNOR2_X1 U831 ( .A(n1167), .B(n1168), .ZN(n1166) );
NOR2_X1 U832 ( .A1(n1121), .A2(n1169), .ZN(n1168) );
NOR2_X1 U833 ( .A1(n1165), .A2(n1170), .ZN(G63) );
XOR2_X1 U834 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U835 ( .A1(n1124), .A2(n1169), .ZN(n1171) );
NOR3_X1 U836 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(G60) );
NOR3_X1 U837 ( .A1(n1176), .A2(n1074), .A3(n1075), .ZN(n1175) );
INV_X1 U838 ( .A(G952), .ZN(n1075) );
AND2_X1 U839 ( .A1(n1176), .A2(n1165), .ZN(n1174) );
INV_X1 U840 ( .A(KEYINPUT23), .ZN(n1176) );
XNOR2_X1 U841 ( .A(n1177), .B(n1178), .ZN(n1173) );
NOR2_X1 U842 ( .A1(n1117), .A2(n1169), .ZN(n1178) );
XNOR2_X1 U843 ( .A(G104), .B(n1179), .ZN(G6) );
NOR2_X1 U844 ( .A1(n1165), .A2(n1180), .ZN(G57) );
XOR2_X1 U845 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U846 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND4_X1 U847 ( .A1(KEYINPUT26), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1184) );
NAND3_X1 U848 ( .A1(n1188), .A2(n1189), .A3(n1190), .ZN(n1187) );
INV_X1 U849 ( .A(KEYINPUT11), .ZN(n1189) );
OR2_X1 U850 ( .A1(n1190), .A2(n1188), .ZN(n1186) );
NOR2_X1 U851 ( .A1(KEYINPUT13), .A2(n1191), .ZN(n1188) );
NAND2_X1 U852 ( .A1(KEYINPUT11), .A2(n1191), .ZN(n1185) );
NAND3_X1 U853 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1183) );
NAND2_X1 U854 ( .A1(KEYINPUT56), .A2(n1195), .ZN(n1194) );
NAND3_X1 U855 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(n1193) );
INV_X1 U856 ( .A(KEYINPUT56), .ZN(n1197) );
OR2_X1 U857 ( .A1(n1198), .A2(n1196), .ZN(n1192) );
NOR2_X1 U858 ( .A1(KEYINPUT21), .A2(n1195), .ZN(n1196) );
XOR2_X1 U859 ( .A(n1199), .B(n1200), .Z(n1181) );
NAND2_X1 U860 ( .A1(KEYINPUT37), .A2(n1201), .ZN(n1199) );
NAND2_X1 U861 ( .A1(n1202), .A2(G472), .ZN(n1201) );
NOR2_X1 U862 ( .A1(n1165), .A2(n1203), .ZN(G54) );
XOR2_X1 U863 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U864 ( .A(n1206), .B(n1207), .Z(n1204) );
XOR2_X1 U865 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U866 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U867 ( .A(n1212), .B(n1213), .Z(n1208) );
AND2_X1 U868 ( .A1(G469), .A2(n1202), .ZN(n1213) );
INV_X1 U869 ( .A(n1169), .ZN(n1202) );
NOR2_X1 U870 ( .A1(KEYINPUT57), .A2(n1214), .ZN(n1212) );
XOR2_X1 U871 ( .A(n1215), .B(n1216), .Z(n1206) );
XNOR2_X1 U872 ( .A(n1217), .B(n1218), .ZN(n1216) );
XNOR2_X1 U873 ( .A(G137), .B(KEYINPUT30), .ZN(n1215) );
NOR2_X1 U874 ( .A1(n1165), .A2(n1219), .ZN(G51) );
XNOR2_X1 U875 ( .A(n1220), .B(n1221), .ZN(n1219) );
XOR2_X1 U876 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U877 ( .A1(n1224), .A2(n1169), .ZN(n1223) );
NAND2_X1 U878 ( .A1(G902), .A2(n1077), .ZN(n1169) );
NAND3_X1 U879 ( .A1(n1225), .A2(n1149), .A3(n1226), .ZN(n1077) );
XNOR2_X1 U880 ( .A(n1163), .B(KEYINPUT0), .ZN(n1226) );
AND2_X1 U881 ( .A1(n1227), .A2(n1103), .ZN(n1163) );
XOR2_X1 U882 ( .A(n1069), .B(KEYINPUT35), .Z(n1227) );
NAND4_X1 U883 ( .A1(n1228), .A2(n1083), .A3(n1090), .A4(n1229), .ZN(n1069) );
AND4_X1 U884 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1149) );
NOR4_X1 U885 ( .A1(n1234), .A2(n1235), .A3(n1236), .A4(n1237), .ZN(n1233) );
AND2_X1 U886 ( .A1(n1238), .A2(n1239), .ZN(n1232) );
NAND2_X1 U887 ( .A1(n1240), .A2(n1241), .ZN(n1231) );
NAND2_X1 U888 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND4_X1 U889 ( .A1(n1244), .A2(n1245), .A3(n1228), .A4(n1246), .ZN(n1243) );
NOR3_X1 U890 ( .A1(n1247), .A2(KEYINPUT29), .A3(n1103), .ZN(n1246) );
NAND2_X1 U891 ( .A1(n1248), .A2(n1092), .ZN(n1242) );
NAND2_X1 U892 ( .A1(KEYINPUT29), .A2(n1249), .ZN(n1230) );
INV_X1 U893 ( .A(n1164), .ZN(n1225) );
NAND4_X1 U894 ( .A1(n1250), .A2(n1251), .A3(n1179), .A4(n1252), .ZN(n1164) );
AND4_X1 U895 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1252) );
NAND4_X1 U896 ( .A1(n1092), .A2(n1257), .A3(n1083), .A4(n1229), .ZN(n1179) );
NAND2_X1 U897 ( .A1(n1258), .A2(n1259), .ZN(n1222) );
OR2_X1 U898 ( .A1(n1146), .A2(n1260), .ZN(n1259) );
NOR2_X1 U899 ( .A1(n1074), .A2(G952), .ZN(n1165) );
XOR2_X1 U900 ( .A(n1237), .B(n1261), .Z(G48) );
XOR2_X1 U901 ( .A(KEYINPUT38), .B(G146), .Z(n1261) );
AND2_X1 U902 ( .A1(n1262), .A2(n1092), .ZN(n1237) );
XOR2_X1 U903 ( .A(G143), .B(n1249), .Z(G45) );
AND3_X1 U904 ( .A1(n1257), .A2(n1240), .A3(n1263), .ZN(n1249) );
NOR3_X1 U905 ( .A1(n1264), .A2(n1247), .A3(n1265), .ZN(n1263) );
XNOR2_X1 U906 ( .A(G140), .B(n1239), .ZN(G42) );
NAND3_X1 U907 ( .A1(n1092), .A2(n1266), .A3(n1248), .ZN(n1239) );
XNOR2_X1 U908 ( .A(G137), .B(n1238), .ZN(G39) );
NAND3_X1 U909 ( .A1(n1267), .A2(n1093), .A3(n1248), .ZN(n1238) );
NAND3_X1 U910 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(G36) );
NAND2_X1 U911 ( .A1(n1236), .A2(n1271), .ZN(n1270) );
NAND2_X1 U912 ( .A1(n1272), .A2(n1273), .ZN(n1269) );
INV_X1 U913 ( .A(KEYINPUT18), .ZN(n1273) );
NAND2_X1 U914 ( .A1(n1274), .A2(n1275), .ZN(n1272) );
XNOR2_X1 U915 ( .A(KEYINPUT20), .B(n1271), .ZN(n1274) );
NAND2_X1 U916 ( .A1(KEYINPUT18), .A2(n1276), .ZN(n1268) );
NAND2_X1 U917 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NAND2_X1 U918 ( .A1(KEYINPUT20), .A2(n1271), .ZN(n1278) );
OR3_X1 U919 ( .A1(n1236), .A2(KEYINPUT20), .A3(n1271), .ZN(n1277) );
INV_X1 U920 ( .A(n1275), .ZN(n1236) );
NAND3_X1 U921 ( .A1(n1090), .A2(n1240), .A3(n1248), .ZN(n1275) );
AND3_X1 U922 ( .A1(n1228), .A2(n1244), .A3(n1085), .ZN(n1248) );
XNOR2_X1 U923 ( .A(G131), .B(n1279), .ZN(G33) );
NAND3_X1 U924 ( .A1(n1280), .A2(n1085), .A3(n1281), .ZN(n1279) );
NOR3_X1 U925 ( .A1(n1282), .A2(n1264), .A3(n1109), .ZN(n1281) );
INV_X1 U926 ( .A(n1240), .ZN(n1109) );
NOR2_X1 U927 ( .A1(n1283), .A2(n1106), .ZN(n1085) );
XNOR2_X1 U928 ( .A(n1228), .B(KEYINPUT62), .ZN(n1280) );
XOR2_X1 U929 ( .A(n1235), .B(n1284), .Z(G30) );
XNOR2_X1 U930 ( .A(KEYINPUT39), .B(n1285), .ZN(n1284) );
AND2_X1 U931 ( .A1(n1262), .A2(n1090), .ZN(n1235) );
AND3_X1 U932 ( .A1(n1257), .A2(n1244), .A3(n1267), .ZN(n1262) );
XNOR2_X1 U933 ( .A(G101), .B(n1250), .ZN(G3) );
NAND2_X1 U934 ( .A1(n1286), .A2(n1240), .ZN(n1250) );
XOR2_X1 U935 ( .A(G125), .B(n1234), .Z(G27) );
AND3_X1 U936 ( .A1(n1092), .A2(n1089), .A3(n1287), .ZN(n1234) );
NOR3_X1 U937 ( .A1(n1068), .A2(n1264), .A3(n1108), .ZN(n1287) );
INV_X1 U938 ( .A(n1266), .ZN(n1108) );
INV_X1 U939 ( .A(n1244), .ZN(n1264) );
NAND2_X1 U940 ( .A1(n1288), .A2(n1289), .ZN(n1244) );
NAND4_X1 U941 ( .A1(G953), .A2(G902), .A3(n1290), .A4(n1291), .ZN(n1289) );
INV_X1 U942 ( .A(G900), .ZN(n1291) );
XNOR2_X1 U943 ( .A(G122), .B(n1251), .ZN(G24) );
NAND4_X1 U944 ( .A1(n1292), .A2(n1083), .A3(n1245), .A4(n1293), .ZN(n1251) );
AND2_X1 U945 ( .A1(n1294), .A2(n1295), .ZN(n1083) );
XNOR2_X1 U946 ( .A(KEYINPUT59), .B(n1296), .ZN(n1294) );
NAND2_X1 U947 ( .A1(n1297), .A2(n1298), .ZN(G21) );
NAND2_X1 U948 ( .A1(n1299), .A2(n1256), .ZN(n1298) );
NAND2_X1 U949 ( .A1(n1300), .A2(n1301), .ZN(n1299) );
NAND2_X1 U950 ( .A1(KEYINPUT42), .A2(KEYINPUT4), .ZN(n1301) );
NAND3_X1 U951 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1297) );
INV_X1 U952 ( .A(KEYINPUT42), .ZN(n1304) );
OR2_X1 U953 ( .A1(G119), .A2(KEYINPUT4), .ZN(n1303) );
NAND2_X1 U954 ( .A1(KEYINPUT4), .A2(n1305), .ZN(n1302) );
OR2_X1 U955 ( .A1(n1256), .A2(G119), .ZN(n1305) );
NAND3_X1 U956 ( .A1(n1267), .A2(n1093), .A3(n1292), .ZN(n1256) );
XNOR2_X1 U957 ( .A(G116), .B(n1255), .ZN(G18) );
NAND3_X1 U958 ( .A1(n1090), .A2(n1240), .A3(n1292), .ZN(n1255) );
XNOR2_X1 U959 ( .A(G113), .B(n1254), .ZN(G15) );
NAND3_X1 U960 ( .A1(n1292), .A2(n1240), .A3(n1092), .ZN(n1254) );
INV_X1 U961 ( .A(n1282), .ZN(n1092) );
NAND2_X1 U962 ( .A1(n1306), .A2(n1293), .ZN(n1282) );
XNOR2_X1 U963 ( .A(n1265), .B(KEYINPUT41), .ZN(n1306) );
NAND2_X1 U964 ( .A1(n1307), .A2(n1308), .ZN(n1240) );
NAND2_X1 U965 ( .A1(n1267), .A2(n1309), .ZN(n1308) );
OR3_X1 U966 ( .A1(n1310), .A2(n1295), .A3(n1309), .ZN(n1307) );
INV_X1 U967 ( .A(KEYINPUT59), .ZN(n1309) );
AND3_X1 U968 ( .A1(n1103), .A2(n1229), .A3(n1089), .ZN(n1292) );
AND2_X1 U969 ( .A1(n1311), .A2(n1098), .ZN(n1089) );
XNOR2_X1 U970 ( .A(n1097), .B(KEYINPUT34), .ZN(n1311) );
XNOR2_X1 U971 ( .A(G110), .B(n1253), .ZN(G12) );
NAND2_X1 U972 ( .A1(n1286), .A2(n1266), .ZN(n1253) );
NAND2_X1 U973 ( .A1(n1312), .A2(n1313), .ZN(n1266) );
NAND2_X1 U974 ( .A1(n1267), .A2(n1314), .ZN(n1313) );
INV_X1 U975 ( .A(KEYINPUT24), .ZN(n1314) );
NOR2_X1 U976 ( .A1(n1295), .A2(n1296), .ZN(n1267) );
INV_X1 U977 ( .A(n1310), .ZN(n1296) );
NAND3_X1 U978 ( .A1(n1310), .A2(n1295), .A3(KEYINPUT24), .ZN(n1312) );
XNOR2_X1 U979 ( .A(n1128), .B(n1315), .ZN(n1295) );
NOR2_X1 U980 ( .A1(G472), .A2(KEYINPUT5), .ZN(n1315) );
NAND2_X1 U981 ( .A1(n1316), .A2(n1317), .ZN(n1128) );
XOR2_X1 U982 ( .A(n1318), .B(n1319), .Z(n1316) );
NOR2_X1 U983 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
XOR2_X1 U984 ( .A(KEYINPUT51), .B(n1322), .Z(n1321) );
NOR2_X1 U985 ( .A1(n1190), .A2(n1191), .ZN(n1322) );
AND2_X1 U986 ( .A1(n1190), .A2(n1191), .ZN(n1320) );
NAND2_X1 U987 ( .A1(n1323), .A2(G210), .ZN(n1191) );
INV_X1 U988 ( .A(G101), .ZN(n1190) );
XOR2_X1 U989 ( .A(n1324), .B(n1325), .Z(n1318) );
NOR2_X1 U990 ( .A1(KEYINPUT43), .A2(n1200), .ZN(n1325) );
XNOR2_X1 U991 ( .A(n1326), .B(n1327), .ZN(n1200) );
XNOR2_X1 U992 ( .A(G116), .B(n1328), .ZN(n1327) );
NAND2_X1 U993 ( .A1(KEYINPUT2), .A2(n1300), .ZN(n1326) );
NAND3_X1 U994 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1324) );
NAND2_X1 U995 ( .A1(KEYINPUT33), .A2(n1195), .ZN(n1331) );
INV_X1 U996 ( .A(n1145), .ZN(n1195) );
OR3_X1 U997 ( .A1(n1332), .A2(KEYINPUT33), .A3(n1333), .ZN(n1330) );
NAND2_X1 U998 ( .A1(n1333), .A2(n1332), .ZN(n1329) );
NAND2_X1 U999 ( .A1(KEYINPUT32), .A2(n1145), .ZN(n1332) );
INV_X1 U1000 ( .A(n1198), .ZN(n1333) );
XOR2_X1 U1001 ( .A(n1122), .B(n1121), .Z(n1310) );
NAND2_X1 U1002 ( .A1(G217), .A2(n1334), .ZN(n1121) );
NAND2_X1 U1003 ( .A1(n1167), .A2(n1317), .ZN(n1122) );
XNOR2_X1 U1004 ( .A(n1335), .B(n1336), .ZN(n1167) );
XOR2_X1 U1005 ( .A(n1337), .B(n1211), .Z(n1336) );
XOR2_X1 U1006 ( .A(n1338), .B(n1339), .Z(n1335) );
AND3_X1 U1007 ( .A1(G221), .A2(n1074), .A3(G234), .ZN(n1339) );
XOR2_X1 U1008 ( .A(n1340), .B(G137), .Z(n1338) );
NAND3_X1 U1009 ( .A1(n1341), .A2(n1342), .A3(n1343), .ZN(n1340) );
NAND2_X1 U1010 ( .A1(KEYINPUT63), .A2(n1344), .ZN(n1343) );
INV_X1 U1011 ( .A(n1345), .ZN(n1344) );
OR3_X1 U1012 ( .A1(n1346), .A2(KEYINPUT63), .A3(G128), .ZN(n1342) );
NAND2_X1 U1013 ( .A1(G128), .A2(n1346), .ZN(n1341) );
NAND2_X1 U1014 ( .A1(KEYINPUT12), .A2(n1345), .ZN(n1346) );
XOR2_X1 U1015 ( .A(G119), .B(KEYINPUT48), .Z(n1345) );
AND3_X1 U1016 ( .A1(n1093), .A2(n1229), .A3(n1257), .ZN(n1286) );
NOR2_X1 U1017 ( .A1(n1068), .A2(n1095), .ZN(n1257) );
INV_X1 U1018 ( .A(n1228), .ZN(n1095) );
NOR2_X1 U1019 ( .A1(n1098), .A2(n1097), .ZN(n1228) );
AND2_X1 U1020 ( .A1(G221), .A2(n1334), .ZN(n1097) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1317), .ZN(n1334) );
XNOR2_X1 U1022 ( .A(n1130), .B(KEYINPUT16), .ZN(n1098) );
XOR2_X1 U1023 ( .A(n1347), .B(G469), .Z(n1130) );
NAND2_X1 U1024 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
XOR2_X1 U1025 ( .A(n1350), .B(n1351), .Z(n1349) );
XNOR2_X1 U1026 ( .A(n1214), .B(n1211), .ZN(n1351) );
XOR2_X1 U1027 ( .A(G140), .B(n1352), .Z(n1211) );
NAND2_X1 U1028 ( .A1(G227), .A2(n1074), .ZN(n1214) );
XOR2_X1 U1029 ( .A(n1353), .B(KEYINPUT44), .Z(n1350) );
NAND3_X1 U1030 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1353) );
NAND2_X1 U1031 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
INV_X1 U1032 ( .A(KEYINPUT15), .ZN(n1358) );
NAND3_X1 U1033 ( .A1(KEYINPUT15), .A2(n1359), .A3(n1145), .ZN(n1355) );
OR2_X1 U1034 ( .A1(n1145), .A2(n1359), .ZN(n1354) );
NOR2_X1 U1035 ( .A1(n1360), .A2(n1357), .ZN(n1359) );
XOR2_X1 U1036 ( .A(n1205), .B(n1140), .Z(n1357) );
XNOR2_X1 U1037 ( .A(n1285), .B(n1218), .ZN(n1140) );
NOR2_X1 U1038 ( .A1(KEYINPUT25), .A2(n1361), .ZN(n1218) );
INV_X1 U1039 ( .A(G128), .ZN(n1285) );
XNOR2_X1 U1040 ( .A(n1362), .B(n1363), .ZN(n1205) );
XNOR2_X1 U1041 ( .A(n1364), .B(G101), .ZN(n1363) );
INV_X1 U1042 ( .A(G107), .ZN(n1364) );
NAND2_X1 U1043 ( .A1(KEYINPUT45), .A2(G104), .ZN(n1362) );
INV_X1 U1044 ( .A(KEYINPUT1), .ZN(n1360) );
XOR2_X1 U1045 ( .A(G131), .B(n1143), .Z(n1145) );
XNOR2_X1 U1046 ( .A(G137), .B(n1271), .ZN(n1143) );
XNOR2_X1 U1047 ( .A(G902), .B(KEYINPUT46), .ZN(n1348) );
INV_X1 U1048 ( .A(n1103), .ZN(n1068) );
NOR2_X1 U1049 ( .A1(n1104), .A2(n1106), .ZN(n1103) );
AND2_X1 U1050 ( .A1(G214), .A2(n1365), .ZN(n1106) );
INV_X1 U1051 ( .A(n1283), .ZN(n1104) );
XOR2_X1 U1052 ( .A(n1366), .B(n1224), .Z(n1283) );
NAND2_X1 U1053 ( .A1(G210), .A2(n1365), .ZN(n1224) );
NAND2_X1 U1054 ( .A1(n1317), .A2(n1367), .ZN(n1365) );
INV_X1 U1055 ( .A(G237), .ZN(n1367) );
NAND2_X1 U1056 ( .A1(n1368), .A2(n1317), .ZN(n1366) );
INV_X1 U1057 ( .A(G902), .ZN(n1317) );
XNOR2_X1 U1058 ( .A(n1369), .B(n1370), .ZN(n1368) );
INV_X1 U1059 ( .A(n1220), .ZN(n1370) );
XOR2_X1 U1060 ( .A(n1160), .B(n1161), .Z(n1220) );
XNOR2_X1 U1061 ( .A(n1371), .B(n1372), .ZN(n1161) );
XNOR2_X1 U1062 ( .A(n1300), .B(G116), .ZN(n1372) );
INV_X1 U1063 ( .A(G119), .ZN(n1300) );
NAND2_X1 U1064 ( .A1(KEYINPUT36), .A2(n1328), .ZN(n1371) );
INV_X1 U1065 ( .A(G113), .ZN(n1328) );
XNOR2_X1 U1066 ( .A(n1373), .B(n1374), .ZN(n1160) );
XOR2_X1 U1067 ( .A(n1375), .B(n1352), .Z(n1374) );
XOR2_X1 U1068 ( .A(G110), .B(KEYINPUT50), .Z(n1352) );
XNOR2_X1 U1069 ( .A(G107), .B(G101), .ZN(n1373) );
NAND3_X1 U1070 ( .A1(n1376), .A2(n1377), .A3(n1378), .ZN(n1369) );
NAND2_X1 U1071 ( .A1(n1379), .A2(n1380), .ZN(n1378) );
NAND2_X1 U1072 ( .A1(n1381), .A2(n1382), .ZN(n1377) );
INV_X1 U1073 ( .A(KEYINPUT19), .ZN(n1382) );
NAND3_X1 U1074 ( .A1(n1383), .A2(n1384), .A3(n1385), .ZN(n1381) );
NAND2_X1 U1075 ( .A1(n1386), .A2(n1146), .ZN(n1384) );
NAND2_X1 U1076 ( .A1(n1380), .A2(n1387), .ZN(n1383) );
NAND2_X1 U1077 ( .A1(KEYINPUT19), .A2(n1388), .ZN(n1376) );
NAND2_X1 U1078 ( .A1(n1258), .A2(n1389), .ZN(n1388) );
NAND2_X1 U1079 ( .A1(n1386), .A2(n1380), .ZN(n1389) );
NAND2_X1 U1080 ( .A1(n1260), .A2(n1146), .ZN(n1258) );
NOR2_X1 U1081 ( .A1(n1379), .A2(n1386), .ZN(n1260) );
NOR2_X1 U1082 ( .A1(n1387), .A2(n1198), .ZN(n1386) );
INV_X1 U1083 ( .A(n1385), .ZN(n1379) );
NAND2_X1 U1084 ( .A1(n1198), .A2(n1387), .ZN(n1385) );
NAND2_X1 U1085 ( .A1(G224), .A2(n1074), .ZN(n1387) );
XOR2_X1 U1086 ( .A(G128), .B(n1361), .Z(n1198) );
XOR2_X1 U1087 ( .A(G146), .B(n1390), .Z(n1361) );
NAND2_X1 U1088 ( .A1(n1391), .A2(n1392), .ZN(n1229) );
NAND4_X1 U1089 ( .A1(G953), .A2(G902), .A3(n1290), .A4(n1158), .ZN(n1392) );
INV_X1 U1090 ( .A(G898), .ZN(n1158) );
XNOR2_X1 U1091 ( .A(n1079), .B(KEYINPUT53), .ZN(n1391) );
INV_X1 U1092 ( .A(n1288), .ZN(n1079) );
NAND3_X1 U1093 ( .A1(n1290), .A2(n1074), .A3(G952), .ZN(n1288) );
NAND2_X1 U1094 ( .A1(G237), .A2(G234), .ZN(n1290) );
NAND2_X1 U1095 ( .A1(n1393), .A2(n1394), .ZN(n1093) );
NAND2_X1 U1096 ( .A1(n1090), .A2(n1395), .ZN(n1394) );
INV_X1 U1097 ( .A(KEYINPUT41), .ZN(n1395) );
NOR2_X1 U1098 ( .A1(n1293), .A2(n1265), .ZN(n1090) );
NAND3_X1 U1099 ( .A1(n1265), .A2(n1247), .A3(KEYINPUT41), .ZN(n1393) );
INV_X1 U1100 ( .A(n1293), .ZN(n1247) );
NAND2_X1 U1101 ( .A1(n1396), .A2(n1397), .ZN(n1293) );
NAND2_X1 U1102 ( .A1(n1119), .A2(n1117), .ZN(n1397) );
XOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1398), .Z(n1396) );
NOR2_X1 U1104 ( .A1(n1119), .A2(n1117), .ZN(n1398) );
INV_X1 U1105 ( .A(G475), .ZN(n1117) );
NOR2_X1 U1106 ( .A1(n1399), .A2(G902), .ZN(n1119) );
INV_X1 U1107 ( .A(n1177), .ZN(n1399) );
XNOR2_X1 U1108 ( .A(n1400), .B(n1401), .ZN(n1177) );
XNOR2_X1 U1109 ( .A(n1402), .B(n1337), .ZN(n1401) );
XNOR2_X1 U1110 ( .A(G146), .B(n1380), .ZN(n1337) );
INV_X1 U1111 ( .A(n1146), .ZN(n1380) );
XOR2_X1 U1112 ( .A(G125), .B(KEYINPUT47), .Z(n1146) );
NAND2_X1 U1113 ( .A1(n1403), .A2(KEYINPUT60), .ZN(n1402) );
XNOR2_X1 U1114 ( .A(G113), .B(n1375), .ZN(n1403) );
XNOR2_X1 U1115 ( .A(G104), .B(n1404), .ZN(n1375) );
XOR2_X1 U1116 ( .A(n1405), .B(n1406), .Z(n1400) );
XNOR2_X1 U1117 ( .A(G140), .B(n1217), .ZN(n1406) );
INV_X1 U1118 ( .A(G131), .ZN(n1217) );
NAND2_X1 U1119 ( .A1(KEYINPUT55), .A2(n1407), .ZN(n1405) );
XOR2_X1 U1120 ( .A(n1408), .B(n1390), .Z(n1407) );
NAND2_X1 U1121 ( .A1(n1323), .A2(G214), .ZN(n1408) );
NOR2_X1 U1122 ( .A1(G953), .A2(G237), .ZN(n1323) );
INV_X1 U1123 ( .A(n1245), .ZN(n1265) );
NAND2_X1 U1124 ( .A1(n1127), .A2(n1409), .ZN(n1245) );
OR2_X1 U1125 ( .A1(n1124), .A2(n1123), .ZN(n1409) );
NAND2_X1 U1126 ( .A1(n1123), .A2(n1124), .ZN(n1127) );
INV_X1 U1127 ( .A(G478), .ZN(n1124) );
NOR2_X1 U1128 ( .A1(n1172), .A2(G902), .ZN(n1123) );
XNOR2_X1 U1129 ( .A(n1410), .B(n1411), .ZN(n1172) );
XNOR2_X1 U1130 ( .A(n1210), .B(n1412), .ZN(n1411) );
XOR2_X1 U1131 ( .A(n1413), .B(n1414), .Z(n1412) );
NOR2_X1 U1132 ( .A1(n1415), .A2(n1416), .ZN(n1414) );
XOR2_X1 U1133 ( .A(n1417), .B(KEYINPUT9), .Z(n1416) );
NAND2_X1 U1134 ( .A1(G116), .A2(n1404), .ZN(n1417) );
NOR2_X1 U1135 ( .A1(G116), .A2(n1404), .ZN(n1415) );
INV_X1 U1136 ( .A(G122), .ZN(n1404) );
NAND2_X1 U1137 ( .A1(KEYINPUT3), .A2(n1390), .ZN(n1413) );
XNOR2_X1 U1138 ( .A(G143), .B(KEYINPUT27), .ZN(n1390) );
XNOR2_X1 U1139 ( .A(G128), .B(n1271), .ZN(n1210) );
INV_X1 U1140 ( .A(G134), .ZN(n1271) );
XOR2_X1 U1141 ( .A(n1418), .B(n1419), .Z(n1410) );
AND3_X1 U1142 ( .A1(G217), .A2(n1074), .A3(G234), .ZN(n1419) );
INV_X1 U1143 ( .A(G953), .ZN(n1074) );
XNOR2_X1 U1144 ( .A(G107), .B(KEYINPUT17), .ZN(n1418) );
endmodule


