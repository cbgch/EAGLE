//Key = 0100001111101111001111010101100011010000010110110110111101110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260;

XNOR2_X1 U688 ( .A(G107), .B(n951), .ZN(G9) );
NOR2_X1 U689 ( .A1(n952), .A2(n953), .ZN(G75) );
NOR3_X1 U690 ( .A1(n954), .A2(n955), .A3(n956), .ZN(n953) );
NOR2_X1 U691 ( .A1(n957), .A2(n958), .ZN(n955) );
NOR2_X1 U692 ( .A1(n959), .A2(n960), .ZN(n957) );
NOR2_X1 U693 ( .A1(n961), .A2(n962), .ZN(n960) );
INV_X1 U694 ( .A(KEYINPUT56), .ZN(n962) );
NOR4_X1 U695 ( .A1(n963), .A2(n964), .A3(n965), .A4(n966), .ZN(n961) );
NOR2_X1 U696 ( .A1(n967), .A2(n966), .ZN(n959) );
NOR2_X1 U697 ( .A1(n968), .A2(n969), .ZN(n967) );
NOR2_X1 U698 ( .A1(n970), .A2(n971), .ZN(n969) );
INV_X1 U699 ( .A(n972), .ZN(n971) );
NOR2_X1 U700 ( .A1(n973), .A2(n974), .ZN(n970) );
NOR2_X1 U701 ( .A1(n975), .A2(n965), .ZN(n974) );
NOR2_X1 U702 ( .A1(n976), .A2(n977), .ZN(n975) );
NOR2_X1 U703 ( .A1(n978), .A2(n979), .ZN(n976) );
NOR2_X1 U704 ( .A1(n980), .A2(n981), .ZN(n973) );
XNOR2_X1 U705 ( .A(KEYINPUT41), .B(n964), .ZN(n981) );
NOR4_X1 U706 ( .A1(KEYINPUT56), .A2(n963), .A3(n964), .A4(n965), .ZN(n968) );
INV_X1 U707 ( .A(n982), .ZN(n965) );
NAND3_X1 U708 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n954) );
NAND3_X1 U709 ( .A1(n986), .A2(n987), .A3(n988), .ZN(n985) );
INV_X1 U710 ( .A(n966), .ZN(n988) );
NAND2_X1 U711 ( .A1(n989), .A2(n990), .ZN(n987) );
NAND3_X1 U712 ( .A1(n982), .A2(n991), .A3(n992), .ZN(n990) );
NAND3_X1 U713 ( .A1(n993), .A2(n994), .A3(n972), .ZN(n989) );
OR2_X1 U714 ( .A1(n958), .A2(n995), .ZN(n994) );
NAND2_X1 U715 ( .A1(n996), .A2(n958), .ZN(n993) );
NAND2_X1 U716 ( .A1(n982), .A2(n997), .ZN(n996) );
NAND2_X1 U717 ( .A1(n998), .A2(n999), .ZN(n997) );
NOR3_X1 U718 ( .A1(n1000), .A2(G953), .A3(G952), .ZN(n952) );
INV_X1 U719 ( .A(n983), .ZN(n1000) );
NAND4_X1 U720 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n983) );
NOR4_X1 U721 ( .A1(n964), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1004) );
XNOR2_X1 U722 ( .A(G478), .B(n1008), .ZN(n1007) );
XOR2_X1 U723 ( .A(KEYINPUT39), .B(n1009), .Z(n1006) );
NOR2_X1 U724 ( .A1(G475), .A2(n1010), .ZN(n1009) );
NOR2_X1 U725 ( .A1(n998), .A2(n1011), .ZN(n1003) );
AND2_X1 U726 ( .A1(n1010), .A2(G475), .ZN(n1011) );
XNOR2_X1 U727 ( .A(n1012), .B(n1013), .ZN(n1002) );
NOR2_X1 U728 ( .A1(n1014), .A2(KEYINPUT45), .ZN(n1013) );
INV_X1 U729 ( .A(n1015), .ZN(n1014) );
XNOR2_X1 U730 ( .A(n1016), .B(n1017), .ZN(n1001) );
NAND2_X1 U731 ( .A1(KEYINPUT35), .A2(n1018), .ZN(n1017) );
XNOR2_X1 U732 ( .A(KEYINPUT13), .B(n1019), .ZN(n1018) );
NAND2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(G72) );
NAND2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
OR2_X1 U736 ( .A1(n984), .A2(G227), .ZN(n1025) );
INV_X1 U737 ( .A(n1026), .ZN(n1024) );
NAND2_X1 U738 ( .A1(n1027), .A2(n1028), .ZN(n1020) );
INV_X1 U739 ( .A(n1022), .ZN(n1028) );
NOR3_X1 U740 ( .A1(KEYINPUT4), .A2(n1029), .A3(n1030), .ZN(n1022) );
NOR2_X1 U741 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U742 ( .A1(n1026), .A2(n1033), .ZN(n1031) );
NOR3_X1 U743 ( .A1(n1034), .A2(n1026), .A3(n1033), .ZN(n1029) );
XOR2_X1 U744 ( .A(n1035), .B(n1036), .Z(n1033) );
XOR2_X1 U745 ( .A(n1037), .B(n1038), .Z(n1036) );
XNOR2_X1 U746 ( .A(G140), .B(n1039), .ZN(n1038) );
NOR2_X1 U747 ( .A1(KEYINPUT48), .A2(n1040), .ZN(n1039) );
XOR2_X1 U748 ( .A(KEYINPUT27), .B(n1041), .Z(n1040) );
NAND2_X1 U749 ( .A1(KEYINPUT20), .A2(n1042), .ZN(n1037) );
XNOR2_X1 U750 ( .A(n1043), .B(n1044), .ZN(n1035) );
XOR2_X1 U751 ( .A(n1032), .B(KEYINPUT12), .Z(n1034) );
NAND2_X1 U752 ( .A1(n1045), .A2(n1046), .ZN(n1032) );
NAND2_X1 U753 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
XNOR2_X1 U754 ( .A(KEYINPUT23), .B(n984), .ZN(n1045) );
NAND2_X1 U755 ( .A1(G953), .A2(n1049), .ZN(n1027) );
NAND2_X1 U756 ( .A1(G900), .A2(G227), .ZN(n1049) );
XOR2_X1 U757 ( .A(n1050), .B(n1051), .Z(G69) );
XOR2_X1 U758 ( .A(n1052), .B(n1053), .Z(n1051) );
NAND2_X1 U759 ( .A1(G953), .A2(n1054), .ZN(n1053) );
NAND2_X1 U760 ( .A1(G898), .A2(G224), .ZN(n1054) );
NAND2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1052) );
NAND2_X1 U762 ( .A1(G953), .A2(n1057), .ZN(n1056) );
XOR2_X1 U763 ( .A(n1058), .B(n1059), .Z(n1055) );
XNOR2_X1 U764 ( .A(n1060), .B(n1061), .ZN(n1058) );
NAND2_X1 U765 ( .A1(KEYINPUT44), .A2(n1062), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1063), .A2(G953), .ZN(n1050) );
NOR2_X1 U767 ( .A1(n1064), .A2(n1065), .ZN(G66) );
XOR2_X1 U768 ( .A(n1066), .B(n1067), .Z(n1065) );
NAND3_X1 U769 ( .A1(n1016), .A2(n956), .A3(n1068), .ZN(n1066) );
XNOR2_X1 U770 ( .A(G902), .B(KEYINPUT46), .ZN(n1068) );
XNOR2_X1 U771 ( .A(n1069), .B(KEYINPUT54), .ZN(n1064) );
NOR2_X1 U772 ( .A1(n1069), .A2(n1070), .ZN(G63) );
XNOR2_X1 U773 ( .A(n1071), .B(n1072), .ZN(n1070) );
AND2_X1 U774 ( .A1(G478), .A2(n1073), .ZN(n1072) );
NOR2_X1 U775 ( .A1(n1069), .A2(n1074), .ZN(G60) );
XOR2_X1 U776 ( .A(n1075), .B(n1076), .Z(n1074) );
AND2_X1 U777 ( .A1(G475), .A2(n1073), .ZN(n1076) );
NAND2_X1 U778 ( .A1(KEYINPUT1), .A2(n1077), .ZN(n1075) );
XNOR2_X1 U779 ( .A(G104), .B(n1078), .ZN(G6) );
NOR2_X1 U780 ( .A1(n1069), .A2(n1079), .ZN(G57) );
XNOR2_X1 U781 ( .A(n1080), .B(n1081), .ZN(n1079) );
AND2_X1 U782 ( .A1(G472), .A2(n1073), .ZN(n1081) );
NOR2_X1 U783 ( .A1(n1069), .A2(n1082), .ZN(G54) );
XOR2_X1 U784 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U785 ( .A(n1085), .B(n1086), .Z(n1084) );
XOR2_X1 U786 ( .A(n1087), .B(KEYINPUT49), .Z(n1086) );
NAND2_X1 U787 ( .A1(KEYINPUT7), .A2(n1061), .ZN(n1087) );
NAND3_X1 U788 ( .A1(n1073), .A2(G469), .A3(KEYINPUT9), .ZN(n1085) );
INV_X1 U789 ( .A(n1088), .ZN(n1073) );
XOR2_X1 U790 ( .A(n1089), .B(n1090), .Z(n1083) );
NOR2_X1 U791 ( .A1(n1091), .A2(n1092), .ZN(G51) );
XNOR2_X1 U792 ( .A(n1069), .B(KEYINPUT50), .ZN(n1092) );
NOR2_X1 U793 ( .A1(n984), .A2(G952), .ZN(n1069) );
XOR2_X1 U794 ( .A(n1093), .B(n1094), .Z(n1091) );
NOR2_X1 U795 ( .A1(n1015), .A2(n1088), .ZN(n1094) );
NAND2_X1 U796 ( .A1(G902), .A2(n956), .ZN(n1088) );
NAND3_X1 U797 ( .A1(n1063), .A2(n1047), .A3(n1095), .ZN(n956) );
XOR2_X1 U798 ( .A(n1048), .B(KEYINPUT61), .Z(n1095) );
AND4_X1 U799 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1047) );
AND4_X1 U800 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
NAND3_X1 U801 ( .A1(n1104), .A2(n991), .A3(n1105), .ZN(n1098) );
XNOR2_X1 U802 ( .A(KEYINPUT34), .B(n958), .ZN(n1104) );
INV_X1 U803 ( .A(n992), .ZN(n958) );
AND4_X1 U804 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1063) );
AND4_X1 U805 ( .A1(n951), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1109) );
NAND3_X1 U806 ( .A1(n972), .A2(n995), .A3(n1113), .ZN(n951) );
AND2_X1 U807 ( .A1(n1114), .A2(n1078), .ZN(n1108) );
NAND3_X1 U808 ( .A1(n1113), .A2(n972), .A3(n1115), .ZN(n1078) );
NAND2_X1 U809 ( .A1(KEYINPUT18), .A2(n1116), .ZN(n1093) );
XOR2_X1 U810 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U811 ( .A(n1119), .B(n1120), .ZN(n1118) );
NAND2_X1 U812 ( .A1(KEYINPUT19), .A2(n1121), .ZN(n1119) );
XOR2_X1 U813 ( .A(KEYINPUT3), .B(n1122), .Z(n1117) );
XNOR2_X1 U814 ( .A(G146), .B(n1096), .ZN(G48) );
NAND3_X1 U815 ( .A1(n1123), .A2(n1124), .A3(n1105), .ZN(n1096) );
XNOR2_X1 U816 ( .A(G143), .B(n1048), .ZN(G45) );
NAND3_X1 U817 ( .A1(n1125), .A2(n1124), .A3(n1126), .ZN(n1048) );
NOR3_X1 U818 ( .A1(n963), .A2(n1127), .A3(n1128), .ZN(n1126) );
INV_X1 U819 ( .A(n1129), .ZN(n963) );
XOR2_X1 U820 ( .A(n1130), .B(n1131), .Z(G42) );
XNOR2_X1 U821 ( .A(G140), .B(KEYINPUT24), .ZN(n1131) );
NAND4_X1 U822 ( .A1(KEYINPUT58), .A2(n992), .A3(n1105), .A4(n991), .ZN(n1130) );
NAND3_X1 U823 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(G39) );
NAND2_X1 U824 ( .A1(KEYINPUT60), .A2(n1097), .ZN(n1134) );
OR3_X1 U825 ( .A1(n1097), .A2(KEYINPUT60), .A3(G137), .ZN(n1133) );
NAND2_X1 U826 ( .A1(G137), .A2(n1135), .ZN(n1132) );
NAND2_X1 U827 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
INV_X1 U828 ( .A(KEYINPUT60), .ZN(n1137) );
XOR2_X1 U829 ( .A(n1097), .B(KEYINPUT8), .Z(n1136) );
NAND4_X1 U830 ( .A1(n992), .A2(n1125), .A3(n1123), .A4(n982), .ZN(n1097) );
NAND2_X1 U831 ( .A1(n1138), .A2(n1139), .ZN(G36) );
OR2_X1 U832 ( .A1(n1140), .A2(G134), .ZN(n1139) );
NAND2_X1 U833 ( .A1(G134), .A2(n1141), .ZN(n1138) );
NAND2_X1 U834 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
OR2_X1 U835 ( .A1(n1102), .A2(KEYINPUT59), .ZN(n1143) );
NAND2_X1 U836 ( .A1(KEYINPUT59), .A2(n1140), .ZN(n1142) );
NAND2_X1 U837 ( .A1(KEYINPUT25), .A2(n1144), .ZN(n1140) );
INV_X1 U838 ( .A(n1102), .ZN(n1144) );
NAND4_X1 U839 ( .A1(n992), .A2(n1125), .A3(n995), .A4(n1129), .ZN(n1102) );
XNOR2_X1 U840 ( .A(G131), .B(n1101), .ZN(G33) );
NAND3_X1 U841 ( .A1(n1105), .A2(n1129), .A3(n992), .ZN(n1101) );
NOR2_X1 U842 ( .A1(n999), .A2(n998), .ZN(n992) );
AND2_X1 U843 ( .A1(n1125), .A2(n1115), .ZN(n1105) );
AND2_X1 U844 ( .A1(n977), .A2(n1145), .ZN(n1125) );
XNOR2_X1 U845 ( .A(n1146), .B(KEYINPUT14), .ZN(n977) );
XNOR2_X1 U846 ( .A(G128), .B(n1100), .ZN(G30) );
NAND4_X1 U847 ( .A1(n1123), .A2(n995), .A3(n1147), .A4(n1146), .ZN(n1100) );
AND2_X1 U848 ( .A1(n1145), .A2(n1124), .ZN(n1147) );
NAND2_X1 U849 ( .A1(n1148), .A2(n1149), .ZN(G3) );
NAND2_X1 U850 ( .A1(G101), .A2(n1114), .ZN(n1149) );
XOR2_X1 U851 ( .A(n1150), .B(KEYINPUT22), .Z(n1148) );
OR2_X1 U852 ( .A1(n1114), .A2(G101), .ZN(n1150) );
NAND3_X1 U853 ( .A1(n1113), .A2(n1129), .A3(n982), .ZN(n1114) );
XNOR2_X1 U854 ( .A(G125), .B(n1103), .ZN(G27) );
NAND4_X1 U855 ( .A1(n991), .A2(n1145), .A3(n1124), .A4(n1151), .ZN(n1103) );
NOR2_X1 U856 ( .A1(n964), .A2(n980), .ZN(n1151) );
INV_X1 U857 ( .A(n1115), .ZN(n980) );
NAND2_X1 U858 ( .A1(n966), .A2(n1152), .ZN(n1145) );
NAND3_X1 U859 ( .A1(G902), .A2(n1153), .A3(n1026), .ZN(n1152) );
NOR2_X1 U860 ( .A1(n984), .A2(G900), .ZN(n1026) );
XNOR2_X1 U861 ( .A(G122), .B(n1106), .ZN(G24) );
NAND4_X1 U862 ( .A1(n1154), .A2(n972), .A3(n1155), .A4(n1156), .ZN(n1106) );
XNOR2_X1 U863 ( .A(G119), .B(n1107), .ZN(G21) );
NAND3_X1 U864 ( .A1(n1123), .A2(n982), .A3(n1154), .ZN(n1107) );
XNOR2_X1 U865 ( .A(G116), .B(n1112), .ZN(G18) );
NAND3_X1 U866 ( .A1(n995), .A2(n1129), .A3(n1154), .ZN(n1112) );
NOR2_X1 U867 ( .A1(n1155), .A2(n1127), .ZN(n995) );
INV_X1 U868 ( .A(n1156), .ZN(n1127) );
XNOR2_X1 U869 ( .A(G113), .B(n1111), .ZN(G15) );
NAND3_X1 U870 ( .A1(n1154), .A2(n1129), .A3(n1115), .ZN(n1111) );
NOR2_X1 U871 ( .A1(n1156), .A2(n1128), .ZN(n1115) );
NAND2_X1 U872 ( .A1(n1157), .A2(n1158), .ZN(n1129) );
NAND2_X1 U873 ( .A1(n1123), .A2(n1159), .ZN(n1158) );
INV_X1 U874 ( .A(KEYINPUT6), .ZN(n1159) );
AND2_X1 U875 ( .A1(n1160), .A2(n1005), .ZN(n1123) );
NAND3_X1 U876 ( .A1(n1161), .A2(n1005), .A3(KEYINPUT6), .ZN(n1157) );
AND2_X1 U877 ( .A1(n986), .A2(n1162), .ZN(n1154) );
INV_X1 U878 ( .A(n964), .ZN(n986) );
NAND2_X1 U879 ( .A1(n1163), .A2(n979), .ZN(n964) );
INV_X1 U880 ( .A(n978), .ZN(n1163) );
XNOR2_X1 U881 ( .A(G110), .B(n1110), .ZN(G12) );
NAND3_X1 U882 ( .A1(n1113), .A2(n991), .A3(n982), .ZN(n1110) );
NOR2_X1 U883 ( .A1(n1156), .A2(n1155), .ZN(n982) );
INV_X1 U884 ( .A(n1128), .ZN(n1155) );
XOR2_X1 U885 ( .A(n1010), .B(G475), .Z(n1128) );
NAND2_X1 U886 ( .A1(n1077), .A2(n1164), .ZN(n1010) );
XNOR2_X1 U887 ( .A(n1165), .B(n1166), .ZN(n1077) );
XOR2_X1 U888 ( .A(n1167), .B(n1168), .Z(n1165) );
XOR2_X1 U889 ( .A(n1169), .B(n1170), .Z(n1168) );
XNOR2_X1 U890 ( .A(n1042), .B(G113), .ZN(n1170) );
XNOR2_X1 U891 ( .A(n1171), .B(G140), .ZN(n1169) );
XOR2_X1 U892 ( .A(n1172), .B(n1173), .Z(n1167) );
XOR2_X1 U893 ( .A(G104), .B(n1174), .Z(n1173) );
NOR2_X1 U894 ( .A1(KEYINPUT40), .A2(n1175), .ZN(n1174) );
XOR2_X1 U895 ( .A(n1176), .B(n1177), .Z(n1172) );
NOR2_X1 U896 ( .A1(KEYINPUT2), .A2(n1178), .ZN(n1177) );
INV_X1 U897 ( .A(G131), .ZN(n1178) );
NAND2_X1 U898 ( .A1(n1179), .A2(G214), .ZN(n1176) );
XOR2_X1 U899 ( .A(n1180), .B(n1008), .Z(n1156) );
NAND2_X1 U900 ( .A1(n1071), .A2(n1164), .ZN(n1008) );
XNOR2_X1 U901 ( .A(n1181), .B(n1182), .ZN(n1071) );
XNOR2_X1 U902 ( .A(n1183), .B(n1184), .ZN(n1182) );
XOR2_X1 U903 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND2_X1 U904 ( .A1(KEYINPUT21), .A2(n1187), .ZN(n1185) );
NAND2_X1 U905 ( .A1(G217), .A2(n1188), .ZN(n1187) );
INV_X1 U906 ( .A(n1189), .ZN(n1188) );
XOR2_X1 U907 ( .A(n1190), .B(n1191), .Z(n1181) );
XNOR2_X1 U908 ( .A(n1175), .B(G128), .ZN(n1191) );
INV_X1 U909 ( .A(G143), .ZN(n1175) );
XNOR2_X1 U910 ( .A(G107), .B(G116), .ZN(n1190) );
NAND2_X1 U911 ( .A1(KEYINPUT43), .A2(G478), .ZN(n1180) );
NAND2_X1 U912 ( .A1(n1192), .A2(n1193), .ZN(n991) );
NAND2_X1 U913 ( .A1(n972), .A2(n1194), .ZN(n1193) );
NOR2_X1 U914 ( .A1(n1005), .A2(n1160), .ZN(n972) );
INV_X1 U915 ( .A(n1161), .ZN(n1160) );
OR3_X1 U916 ( .A1(n1005), .A2(n1161), .A3(n1194), .ZN(n1192) );
INV_X1 U917 ( .A(KEYINPUT32), .ZN(n1194) );
XNOR2_X1 U918 ( .A(n1019), .B(n1195), .ZN(n1161) );
XOR2_X1 U919 ( .A(KEYINPUT31), .B(n1196), .Z(n1195) );
NOR2_X1 U920 ( .A1(KEYINPUT37), .A2(n1016), .ZN(n1196) );
AND2_X1 U921 ( .A1(G217), .A2(n1197), .ZN(n1016) );
NAND2_X1 U922 ( .A1(n1067), .A2(n1164), .ZN(n1019) );
XOR2_X1 U923 ( .A(n1198), .B(n1199), .Z(n1067) );
XNOR2_X1 U924 ( .A(n1200), .B(n1201), .ZN(n1199) );
XNOR2_X1 U925 ( .A(n1202), .B(n1203), .ZN(n1201) );
NOR2_X1 U926 ( .A1(KEYINPUT42), .A2(n1204), .ZN(n1203) );
XOR2_X1 U927 ( .A(KEYINPUT17), .B(n1205), .Z(n1204) );
NOR2_X1 U928 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NOR2_X1 U929 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NOR2_X1 U930 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NOR2_X1 U931 ( .A1(KEYINPUT0), .A2(n1212), .ZN(n1210) );
NOR2_X1 U932 ( .A1(n1213), .A2(n1189), .ZN(n1208) );
NOR2_X1 U933 ( .A1(G137), .A2(n1214), .ZN(n1206) );
NOR2_X1 U934 ( .A1(n1215), .A2(KEYINPUT0), .ZN(n1214) );
NOR3_X1 U935 ( .A1(n1211), .A2(n1213), .A3(n1189), .ZN(n1215) );
NAND2_X1 U936 ( .A1(G234), .A2(n984), .ZN(n1189) );
INV_X1 U937 ( .A(G221), .ZN(n1213) );
INV_X1 U938 ( .A(KEYINPUT57), .ZN(n1211) );
NOR2_X1 U939 ( .A1(KEYINPUT38), .A2(n1216), .ZN(n1202) );
XNOR2_X1 U940 ( .A(G146), .B(KEYINPUT33), .ZN(n1216) );
XNOR2_X1 U941 ( .A(n1217), .B(n1090), .ZN(n1198) );
XOR2_X1 U942 ( .A(G110), .B(G140), .Z(n1090) );
XNOR2_X1 U943 ( .A(n1218), .B(G472), .ZN(n1005) );
NAND2_X1 U944 ( .A1(n1080), .A2(n1164), .ZN(n1218) );
XNOR2_X1 U945 ( .A(n1219), .B(n1220), .ZN(n1080) );
XOR2_X1 U946 ( .A(n1221), .B(n1222), .Z(n1220) );
XOR2_X1 U947 ( .A(n1223), .B(n1224), .Z(n1222) );
AND2_X1 U948 ( .A1(G210), .A2(n1179), .ZN(n1224) );
NOR2_X1 U949 ( .A1(G953), .A2(G237), .ZN(n1179) );
NAND2_X1 U950 ( .A1(KEYINPUT10), .A2(n1225), .ZN(n1223) );
XOR2_X1 U951 ( .A(G116), .B(n1200), .Z(n1225) );
XOR2_X1 U952 ( .A(n1226), .B(n1227), .Z(n1219) );
XOR2_X1 U953 ( .A(G113), .B(G101), .Z(n1227) );
AND2_X1 U954 ( .A1(n1162), .A2(n1146), .ZN(n1113) );
AND2_X1 U955 ( .A1(n978), .A2(n979), .ZN(n1146) );
NAND2_X1 U956 ( .A1(G221), .A2(n1197), .ZN(n979) );
NAND2_X1 U957 ( .A1(G234), .A2(n1164), .ZN(n1197) );
XNOR2_X1 U958 ( .A(n1228), .B(n1229), .ZN(n978) );
XOR2_X1 U959 ( .A(KEYINPUT11), .B(G469), .Z(n1229) );
NAND2_X1 U960 ( .A1(n1230), .A2(n1164), .ZN(n1228) );
XOR2_X1 U961 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U962 ( .A(KEYINPUT26), .B(n1233), .Z(n1232) );
NOR2_X1 U963 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
XOR2_X1 U964 ( .A(n1236), .B(KEYINPUT63), .Z(n1235) );
NAND2_X1 U965 ( .A1(G110), .A2(n1237), .ZN(n1236) );
NOR2_X1 U966 ( .A1(G110), .A2(n1237), .ZN(n1234) );
XOR2_X1 U967 ( .A(KEYINPUT55), .B(G140), .Z(n1237) );
XNOR2_X1 U968 ( .A(n1089), .B(n1061), .ZN(n1231) );
XOR2_X1 U969 ( .A(n1238), .B(n1239), .Z(n1089) );
XNOR2_X1 U970 ( .A(n1044), .B(n1221), .ZN(n1239) );
XOR2_X1 U971 ( .A(n1240), .B(n1043), .Z(n1221) );
XOR2_X1 U972 ( .A(G131), .B(G128), .Z(n1043) );
NAND2_X1 U973 ( .A1(KEYINPUT47), .A2(n1241), .ZN(n1240) );
XOR2_X1 U974 ( .A(KEYINPUT16), .B(n1041), .Z(n1241) );
XNOR2_X1 U975 ( .A(n1212), .B(n1186), .ZN(n1041) );
XOR2_X1 U976 ( .A(G134), .B(KEYINPUT51), .Z(n1186) );
INV_X1 U977 ( .A(G137), .ZN(n1212) );
XOR2_X1 U978 ( .A(n1242), .B(KEYINPUT5), .Z(n1238) );
NAND2_X1 U979 ( .A1(G227), .A2(n984), .ZN(n1242) );
AND2_X1 U980 ( .A1(n1124), .A2(n1243), .ZN(n1162) );
NAND2_X1 U981 ( .A1(n966), .A2(n1244), .ZN(n1243) );
NAND4_X1 U982 ( .A1(G953), .A2(G902), .A3(n1153), .A4(n1057), .ZN(n1244) );
INV_X1 U983 ( .A(G898), .ZN(n1057) );
NAND3_X1 U984 ( .A1(n1153), .A2(n984), .A3(G952), .ZN(n966) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1153) );
NOR2_X1 U986 ( .A1(n1245), .A2(n998), .ZN(n1124) );
AND2_X1 U987 ( .A1(G214), .A2(n1246), .ZN(n998) );
INV_X1 U988 ( .A(n999), .ZN(n1245) );
XOR2_X1 U989 ( .A(n1247), .B(n1015), .Z(n999) );
NAND2_X1 U990 ( .A1(G210), .A2(n1246), .ZN(n1015) );
NAND2_X1 U991 ( .A1(n1164), .A2(n1248), .ZN(n1246) );
INV_X1 U992 ( .A(G237), .ZN(n1248) );
XOR2_X1 U993 ( .A(n1012), .B(KEYINPUT29), .Z(n1247) );
NAND2_X1 U994 ( .A1(n1249), .A2(n1164), .ZN(n1012) );
INV_X1 U995 ( .A(G902), .ZN(n1164) );
XNOR2_X1 U996 ( .A(n1250), .B(n1251), .ZN(n1249) );
XOR2_X1 U997 ( .A(n1122), .B(n1252), .Z(n1251) );
NOR2_X1 U998 ( .A1(KEYINPUT36), .A2(n1253), .ZN(n1252) );
INV_X1 U999 ( .A(n1121), .ZN(n1253) );
XNOR2_X1 U1000 ( .A(n1226), .B(n1217), .ZN(n1121) );
XNOR2_X1 U1001 ( .A(n1042), .B(G128), .ZN(n1217) );
INV_X1 U1002 ( .A(G125), .ZN(n1042) );
NAND2_X1 U1003 ( .A1(KEYINPUT15), .A2(n1044), .ZN(n1226) );
XNOR2_X1 U1004 ( .A(G143), .B(n1171), .ZN(n1044) );
INV_X1 U1005 ( .A(G146), .ZN(n1171) );
AND2_X1 U1006 ( .A1(G224), .A2(n984), .ZN(n1122) );
INV_X1 U1007 ( .A(G953), .ZN(n984) );
INV_X1 U1008 ( .A(n1120), .ZN(n1250) );
XNOR2_X1 U1009 ( .A(n1254), .B(n1059), .ZN(n1120) );
XNOR2_X1 U1010 ( .A(G110), .B(n1166), .ZN(n1059) );
INV_X1 U1011 ( .A(n1183), .ZN(n1166) );
XOR2_X1 U1012 ( .A(G122), .B(KEYINPUT28), .Z(n1183) );
NAND2_X1 U1013 ( .A1(KEYINPUT52), .A2(n1255), .ZN(n1254) );
XNOR2_X1 U1014 ( .A(n1062), .B(n1256), .ZN(n1255) );
XNOR2_X1 U1015 ( .A(KEYINPUT53), .B(n1061), .ZN(n1256) );
XNOR2_X1 U1016 ( .A(G101), .B(n1257), .ZN(n1061) );
XNOR2_X1 U1017 ( .A(n1258), .B(G104), .ZN(n1257) );
INV_X1 U1018 ( .A(G107), .ZN(n1258) );
XNOR2_X1 U1019 ( .A(G113), .B(n1259), .ZN(n1062) );
NOR2_X1 U1020 ( .A1(KEYINPUT30), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U1021 ( .A(G116), .B(n1200), .ZN(n1260) );
XOR2_X1 U1022 ( .A(G119), .B(KEYINPUT62), .Z(n1200) );
endmodule


