//Key = 1011101000100000000100000101001100100010110100101101101000100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;

XNOR2_X1 U741 ( .A(G107), .B(n1028), .ZN(G9) );
NOR2_X1 U742 ( .A1(n1029), .A2(n1030), .ZN(G75) );
NOR4_X1 U743 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NOR2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NOR3_X1 U745 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1033) );
XOR2_X1 U746 ( .A(n1036), .B(KEYINPUT21), .Z(n1038) );
NAND4_X1 U747 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1036) );
NAND3_X1 U748 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1031) );
NAND3_X1 U749 ( .A1(n1047), .A2(n1048), .A3(n1040), .ZN(n1046) );
INV_X1 U750 ( .A(n1049), .ZN(n1040) );
NAND2_X1 U751 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND3_X1 U752 ( .A1(n1043), .A2(n1052), .A3(n1041), .ZN(n1051) );
OR2_X1 U753 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U754 ( .A1(n1042), .A2(n1055), .ZN(n1050) );
NAND3_X1 U755 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1043), .A2(n1059), .ZN(n1058) );
NAND2_X1 U757 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
INV_X1 U759 ( .A(n1064), .ZN(n1060) );
NAND3_X1 U760 ( .A1(n1065), .A2(n1066), .A3(n1041), .ZN(n1056) );
NOR3_X1 U761 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1029) );
INV_X1 U762 ( .A(n1044), .ZN(n1067) );
NAND4_X1 U763 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1044) );
NOR4_X1 U764 ( .A1(n1072), .A2(n1062), .A3(n1073), .A4(n1074), .ZN(n1071) );
XOR2_X1 U765 ( .A(n1063), .B(KEYINPUT30), .Z(n1073) );
NOR2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1070) );
XOR2_X1 U767 ( .A(n1077), .B(n1078), .Z(n1076) );
XNOR2_X1 U768 ( .A(KEYINPUT26), .B(n1079), .ZN(n1078) );
NOR3_X1 U769 ( .A1(n1080), .A2(KEYINPUT33), .A3(G902), .ZN(n1077) );
INV_X1 U770 ( .A(n1081), .ZN(n1080) );
XOR2_X1 U771 ( .A(n1082), .B(n1083), .Z(n1069) );
XNOR2_X1 U772 ( .A(n1084), .B(KEYINPUT56), .ZN(n1068) );
XOR2_X1 U773 ( .A(n1085), .B(n1086), .Z(G72) );
XOR2_X1 U774 ( .A(n1087), .B(n1088), .Z(n1086) );
NAND2_X1 U775 ( .A1(G953), .A2(n1089), .ZN(n1088) );
NAND2_X1 U776 ( .A1(G900), .A2(G227), .ZN(n1089) );
NAND2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1087) );
NAND2_X1 U778 ( .A1(G953), .A2(n1092), .ZN(n1091) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1090) );
XNOR2_X1 U780 ( .A(n1095), .B(n1096), .ZN(n1094) );
NOR2_X1 U781 ( .A1(KEYINPUT57), .A2(n1097), .ZN(n1096) );
XNOR2_X1 U782 ( .A(KEYINPUT24), .B(n1098), .ZN(n1097) );
NOR2_X1 U783 ( .A1(KEYINPUT23), .A2(n1099), .ZN(n1093) );
XOR2_X1 U784 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U785 ( .A(G131), .B(n1102), .Z(n1101) );
NOR2_X1 U786 ( .A1(KEYINPUT44), .A2(n1103), .ZN(n1102) );
XOR2_X1 U787 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U788 ( .A1(KEYINPUT61), .A2(n1106), .ZN(n1104) );
NOR2_X1 U789 ( .A1(n1107), .A2(G953), .ZN(n1085) );
XOR2_X1 U790 ( .A(n1108), .B(n1109), .Z(G69) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U792 ( .A1(G953), .A2(n1112), .ZN(n1111) );
NAND2_X1 U793 ( .A1(G898), .A2(G224), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1113), .A2(n1114), .ZN(n1110) );
NAND2_X1 U795 ( .A1(G953), .A2(n1115), .ZN(n1114) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1113) );
XOR2_X1 U797 ( .A(n1118), .B(n1119), .Z(n1117) );
NOR2_X1 U798 ( .A1(n1120), .A2(G953), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(G66) );
XNOR2_X1 U800 ( .A(n1123), .B(n1124), .ZN(n1122) );
NOR3_X1 U801 ( .A1(n1125), .A2(KEYINPUT37), .A3(n1126), .ZN(n1124) );
INV_X1 U802 ( .A(G217), .ZN(n1126) );
NOR2_X1 U803 ( .A1(n1121), .A2(n1127), .ZN(G63) );
XOR2_X1 U804 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U805 ( .A1(n1130), .A2(n1125), .ZN(n1128) );
NOR2_X1 U806 ( .A1(n1121), .A2(n1131), .ZN(G60) );
XNOR2_X1 U807 ( .A(n1081), .B(n1132), .ZN(n1131) );
NOR2_X1 U808 ( .A1(n1079), .A2(n1125), .ZN(n1132) );
XOR2_X1 U809 ( .A(G104), .B(n1133), .Z(G6) );
NOR2_X1 U810 ( .A1(n1121), .A2(n1134), .ZN(G57) );
XOR2_X1 U811 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U812 ( .A(n1137), .B(n1138), .ZN(n1136) );
XNOR2_X1 U813 ( .A(G101), .B(n1139), .ZN(n1138) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XNOR2_X1 U815 ( .A(KEYINPUT54), .B(KEYINPUT16), .ZN(n1140) );
XNOR2_X1 U816 ( .A(n1142), .B(n1143), .ZN(n1135) );
XNOR2_X1 U817 ( .A(n1144), .B(n1145), .ZN(n1142) );
NOR2_X1 U818 ( .A1(n1125), .A2(n1146), .ZN(n1145) );
XOR2_X1 U819 ( .A(KEYINPUT2), .B(G472), .Z(n1146) );
NOR3_X1 U820 ( .A1(n1121), .A2(n1147), .A3(n1148), .ZN(G54) );
NOR2_X1 U821 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
INV_X1 U822 ( .A(n1151), .ZN(n1150) );
NOR2_X1 U823 ( .A1(n1152), .A2(n1153), .ZN(n1149) );
AND2_X1 U824 ( .A1(n1154), .A2(KEYINPUT15), .ZN(n1153) );
NOR3_X1 U825 ( .A1(KEYINPUT15), .A2(n1154), .A3(n1155), .ZN(n1152) );
NOR2_X1 U826 ( .A1(n1156), .A2(n1151), .ZN(n1147) );
XNOR2_X1 U827 ( .A(n1157), .B(n1158), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U829 ( .A(KEYINPUT32), .B(n1161), .Z(n1160) );
AND2_X1 U830 ( .A1(n1162), .A2(n1143), .ZN(n1161) );
NOR2_X1 U831 ( .A1(n1143), .A2(n1162), .ZN(n1159) );
XNOR2_X1 U832 ( .A(n1163), .B(n1119), .ZN(n1162) );
NAND2_X1 U833 ( .A1(n1164), .A2(KEYINPUT51), .ZN(n1157) );
XOR2_X1 U834 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U835 ( .A(KEYINPUT3), .B(KEYINPUT20), .Z(n1166) );
XNOR2_X1 U836 ( .A(n1167), .B(n1168), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1154), .A2(n1155), .ZN(n1156) );
INV_X1 U838 ( .A(KEYINPUT40), .ZN(n1155) );
NAND3_X1 U839 ( .A1(G469), .A2(G902), .A3(n1169), .ZN(n1154) );
XOR2_X1 U840 ( .A(n1032), .B(KEYINPUT59), .Z(n1169) );
NOR2_X1 U841 ( .A1(n1121), .A2(n1170), .ZN(G51) );
XOR2_X1 U842 ( .A(n1171), .B(n1172), .Z(n1170) );
XNOR2_X1 U843 ( .A(n1098), .B(n1173), .ZN(n1172) );
NOR2_X1 U844 ( .A1(n1083), .A2(n1125), .ZN(n1173) );
NAND2_X1 U845 ( .A1(G902), .A2(n1032), .ZN(n1125) );
NAND2_X1 U846 ( .A1(n1120), .A2(n1107), .ZN(n1032) );
AND4_X1 U847 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1107) );
NOR4_X1 U848 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR2_X1 U849 ( .A1(n1182), .A2(n1183), .ZN(n1176) );
AND4_X1 U850 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1120) );
AND4_X1 U851 ( .A1(n1028), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1187) );
NAND3_X1 U852 ( .A1(n1054), .A2(n1043), .A3(n1191), .ZN(n1028) );
NOR2_X1 U853 ( .A1(n1192), .A2(n1133), .ZN(n1186) );
AND3_X1 U854 ( .A1(n1191), .A2(n1043), .A3(n1053), .ZN(n1133) );
NOR4_X1 U855 ( .A1(n1193), .A2(n1057), .A3(n1194), .A4(n1195), .ZN(n1192) );
XNOR2_X1 U856 ( .A(KEYINPUT46), .B(n1035), .ZN(n1195) );
NOR2_X1 U857 ( .A1(n1045), .A2(G952), .ZN(n1121) );
XNOR2_X1 U858 ( .A(G146), .B(n1174), .ZN(G48) );
NAND3_X1 U859 ( .A1(n1053), .A2(n1196), .A3(n1197), .ZN(n1174) );
NAND2_X1 U860 ( .A1(n1198), .A2(n1199), .ZN(G45) );
NAND2_X1 U861 ( .A1(G143), .A2(n1200), .ZN(n1199) );
NAND2_X1 U862 ( .A1(n1201), .A2(n1202), .ZN(n1200) );
NAND2_X1 U863 ( .A1(KEYINPUT62), .A2(KEYINPUT4), .ZN(n1202) );
NAND3_X1 U864 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1198) );
INV_X1 U865 ( .A(KEYINPUT62), .ZN(n1205) );
OR2_X1 U866 ( .A1(n1175), .A2(KEYINPUT4), .ZN(n1204) );
NAND2_X1 U867 ( .A1(KEYINPUT4), .A2(n1206), .ZN(n1203) );
NAND2_X1 U868 ( .A1(n1201), .A2(n1207), .ZN(n1206) );
INV_X1 U869 ( .A(n1175), .ZN(n1201) );
NAND4_X1 U870 ( .A1(n1208), .A2(n1196), .A3(n1209), .A4(n1075), .ZN(n1175) );
XNOR2_X1 U871 ( .A(G140), .B(n1210), .ZN(G42) );
NAND2_X1 U872 ( .A1(KEYINPUT38), .A2(n1183), .ZN(n1210) );
AND3_X1 U873 ( .A1(n1211), .A2(n1064), .A3(n1047), .ZN(n1183) );
XNOR2_X1 U874 ( .A(n1106), .B(n1182), .ZN(G39) );
AND3_X1 U875 ( .A1(n1197), .A2(n1042), .A3(n1047), .ZN(n1182) );
XOR2_X1 U876 ( .A(G134), .B(n1181), .Z(G36) );
AND3_X1 U877 ( .A1(n1047), .A2(n1054), .A3(n1208), .ZN(n1181) );
XOR2_X1 U878 ( .A(G131), .B(n1180), .Z(G33) );
AND3_X1 U879 ( .A1(n1047), .A2(n1053), .A3(n1208), .ZN(n1180) );
AND2_X1 U880 ( .A1(n1212), .A2(n1213), .ZN(n1208) );
NOR2_X1 U881 ( .A1(n1039), .A2(n1072), .ZN(n1047) );
INV_X1 U882 ( .A(n1037), .ZN(n1072) );
XOR2_X1 U883 ( .A(n1179), .B(n1214), .Z(G30) );
NOR2_X1 U884 ( .A1(KEYINPUT53), .A2(n1215), .ZN(n1214) );
AND3_X1 U885 ( .A1(n1054), .A2(n1196), .A3(n1197), .ZN(n1179) );
AND2_X1 U886 ( .A1(n1212), .A2(n1066), .ZN(n1197) );
AND3_X1 U887 ( .A1(n1084), .A2(n1216), .A3(n1064), .ZN(n1212) );
XOR2_X1 U888 ( .A(G101), .B(n1217), .Z(G3) );
NOR2_X1 U889 ( .A1(n1184), .A2(n1218), .ZN(n1217) );
XOR2_X1 U890 ( .A(KEYINPUT60), .B(KEYINPUT39), .Z(n1218) );
NAND4_X1 U891 ( .A1(n1042), .A2(n1191), .A3(n1084), .A4(n1213), .ZN(n1184) );
XNOR2_X1 U892 ( .A(n1098), .B(n1178), .ZN(G27) );
AND3_X1 U893 ( .A1(n1041), .A2(n1196), .A3(n1211), .ZN(n1178) );
AND4_X1 U894 ( .A1(n1066), .A2(n1053), .A3(n1065), .A4(n1216), .ZN(n1211) );
NAND2_X1 U895 ( .A1(n1049), .A2(n1219), .ZN(n1216) );
NAND4_X1 U896 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1092), .ZN(n1219) );
INV_X1 U897 ( .A(G900), .ZN(n1092) );
INV_X1 U898 ( .A(n1035), .ZN(n1196) );
XOR2_X1 U899 ( .A(G122), .B(n1221), .Z(G24) );
NOR2_X1 U900 ( .A1(KEYINPUT63), .A2(n1185), .ZN(n1221) );
NAND4_X1 U901 ( .A1(n1041), .A2(n1043), .A3(n1222), .A4(n1223), .ZN(n1185) );
AND2_X1 U902 ( .A1(n1075), .A2(n1209), .ZN(n1222) );
NOR2_X1 U903 ( .A1(n1084), .A2(n1066), .ZN(n1043) );
XNOR2_X1 U904 ( .A(G119), .B(n1190), .ZN(G21) );
NAND4_X1 U905 ( .A1(n1223), .A2(n1084), .A3(n1066), .A4(n1224), .ZN(n1190) );
AND2_X1 U906 ( .A1(n1042), .A2(n1041), .ZN(n1224) );
XNOR2_X1 U907 ( .A(G116), .B(n1189), .ZN(G18) );
NAND3_X1 U908 ( .A1(n1054), .A2(n1223), .A3(n1225), .ZN(n1189) );
NOR2_X1 U909 ( .A1(n1209), .A2(n1226), .ZN(n1054) );
INV_X1 U910 ( .A(n1075), .ZN(n1226) );
NAND3_X1 U911 ( .A1(n1227), .A2(n1228), .A3(n1229), .ZN(G15) );
NAND4_X1 U912 ( .A1(n1053), .A2(n1225), .A3(n1223), .A4(n1230), .ZN(n1229) );
NAND2_X1 U913 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
NAND2_X1 U914 ( .A1(KEYINPUT52), .A2(n1233), .ZN(n1232) );
NAND3_X1 U915 ( .A1(G113), .A2(n1234), .A3(n1231), .ZN(n1228) );
INV_X1 U916 ( .A(KEYINPUT17), .ZN(n1231) );
NAND4_X1 U917 ( .A1(KEYINPUT52), .A2(n1053), .A3(n1225), .A4(n1223), .ZN(n1234) );
INV_X1 U918 ( .A(n1057), .ZN(n1225) );
NAND3_X1 U919 ( .A1(n1084), .A2(n1213), .A3(n1041), .ZN(n1057) );
AND2_X1 U920 ( .A1(n1235), .A2(n1063), .ZN(n1041) );
XNOR2_X1 U921 ( .A(n1062), .B(KEYINPUT50), .ZN(n1235) );
INV_X1 U922 ( .A(n1194), .ZN(n1053) );
NAND2_X1 U923 ( .A1(n1236), .A2(n1209), .ZN(n1194) );
XNOR2_X1 U924 ( .A(n1075), .B(KEYINPUT18), .ZN(n1236) );
NAND2_X1 U925 ( .A1(KEYINPUT17), .A2(n1233), .ZN(n1227) );
INV_X1 U926 ( .A(G113), .ZN(n1233) );
XNOR2_X1 U927 ( .A(G110), .B(n1188), .ZN(G12) );
NAND4_X1 U928 ( .A1(n1066), .A2(n1042), .A3(n1065), .A4(n1191), .ZN(n1188) );
AND2_X1 U929 ( .A1(n1223), .A2(n1064), .ZN(n1191) );
NOR2_X1 U930 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
AND2_X1 U931 ( .A1(G221), .A2(n1237), .ZN(n1062) );
XOR2_X1 U932 ( .A(n1238), .B(G469), .Z(n1063) );
NAND2_X1 U933 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XOR2_X1 U934 ( .A(n1241), .B(n1242), .Z(n1239) );
XNOR2_X1 U935 ( .A(n1163), .B(n1168), .ZN(n1242) );
XNOR2_X1 U936 ( .A(G110), .B(n1095), .ZN(n1168) );
XOR2_X1 U937 ( .A(n1100), .B(KEYINPUT42), .Z(n1163) );
XNOR2_X1 U938 ( .A(G128), .B(n1243), .ZN(n1100) );
XNOR2_X1 U939 ( .A(n1244), .B(n1143), .ZN(n1241) );
XNOR2_X1 U940 ( .A(n1245), .B(n1246), .ZN(n1244) );
NAND2_X1 U941 ( .A1(KEYINPUT48), .A2(n1119), .ZN(n1246) );
NAND2_X1 U942 ( .A1(KEYINPUT0), .A2(n1167), .ZN(n1245) );
AND2_X1 U943 ( .A1(G227), .A2(n1045), .ZN(n1167) );
NOR2_X1 U944 ( .A1(n1035), .A2(n1193), .ZN(n1223) );
AND2_X1 U945 ( .A1(n1049), .A2(n1247), .ZN(n1193) );
NAND4_X1 U946 ( .A1(G953), .A2(G902), .A3(n1220), .A4(n1115), .ZN(n1247) );
INV_X1 U947 ( .A(G898), .ZN(n1115) );
NAND3_X1 U948 ( .A1(n1220), .A2(n1045), .A3(G952), .ZN(n1049) );
NAND2_X1 U949 ( .A1(G237), .A2(G234), .ZN(n1220) );
NAND2_X1 U950 ( .A1(n1039), .A2(n1037), .ZN(n1035) );
NAND2_X1 U951 ( .A1(G214), .A2(n1248), .ZN(n1037) );
XOR2_X1 U952 ( .A(n1249), .B(n1083), .Z(n1039) );
NAND2_X1 U953 ( .A1(G210), .A2(n1248), .ZN(n1083) );
NAND2_X1 U954 ( .A1(n1240), .A2(n1250), .ZN(n1248) );
INV_X1 U955 ( .A(G237), .ZN(n1250) );
NAND2_X1 U956 ( .A1(KEYINPUT6), .A2(n1082), .ZN(n1249) );
AND3_X1 U957 ( .A1(n1251), .A2(n1252), .A3(n1240), .ZN(n1082) );
NAND2_X1 U958 ( .A1(n1171), .A2(n1098), .ZN(n1252) );
INV_X1 U959 ( .A(G125), .ZN(n1098) );
NAND2_X1 U960 ( .A1(n1253), .A2(G125), .ZN(n1251) );
XOR2_X1 U961 ( .A(KEYINPUT49), .B(n1171), .Z(n1253) );
XNOR2_X1 U962 ( .A(n1254), .B(n1255), .ZN(n1171) );
XNOR2_X1 U963 ( .A(n1256), .B(n1257), .ZN(n1255) );
NOR2_X1 U964 ( .A1(KEYINPUT7), .A2(n1258), .ZN(n1256) );
XOR2_X1 U965 ( .A(n1259), .B(n1119), .Z(n1258) );
XNOR2_X1 U966 ( .A(n1260), .B(n1261), .ZN(n1119) );
XNOR2_X1 U967 ( .A(G101), .B(G107), .ZN(n1260) );
NOR2_X1 U968 ( .A1(KEYINPUT28), .A2(n1262), .ZN(n1259) );
XOR2_X1 U969 ( .A(n1118), .B(KEYINPUT34), .Z(n1262) );
XNOR2_X1 U970 ( .A(n1144), .B(KEYINPUT45), .ZN(n1118) );
XOR2_X1 U971 ( .A(n1116), .B(n1263), .Z(n1254) );
AND2_X1 U972 ( .A1(n1045), .A2(G224), .ZN(n1263) );
XNOR2_X1 U973 ( .A(G110), .B(n1264), .ZN(n1116) );
XOR2_X1 U974 ( .A(KEYINPUT29), .B(G122), .Z(n1264) );
INV_X1 U975 ( .A(n1084), .ZN(n1065) );
XNOR2_X1 U976 ( .A(n1265), .B(G472), .ZN(n1084) );
NAND2_X1 U977 ( .A1(n1266), .A2(n1240), .ZN(n1265) );
XOR2_X1 U978 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U979 ( .A(n1137), .B(n1269), .ZN(n1268) );
XNOR2_X1 U980 ( .A(G101), .B(KEYINPUT43), .ZN(n1269) );
INV_X1 U981 ( .A(n1257), .ZN(n1137) );
NAND2_X1 U982 ( .A1(n1270), .A2(n1271), .ZN(n1257) );
NAND2_X1 U983 ( .A1(G128), .A2(n1243), .ZN(n1271) );
XOR2_X1 U984 ( .A(n1272), .B(KEYINPUT55), .Z(n1270) );
OR2_X1 U985 ( .A1(n1243), .A2(G128), .ZN(n1272) );
XOR2_X1 U986 ( .A(G143), .B(G146), .Z(n1243) );
XNOR2_X1 U987 ( .A(n1273), .B(n1274), .ZN(n1267) );
INV_X1 U988 ( .A(n1144), .ZN(n1274) );
XOR2_X1 U989 ( .A(G113), .B(n1275), .Z(n1144) );
XOR2_X1 U990 ( .A(G119), .B(G116), .Z(n1275) );
XOR2_X1 U991 ( .A(n1141), .B(n1276), .Z(n1273) );
NOR2_X1 U992 ( .A1(KEYINPUT12), .A2(n1143), .ZN(n1276) );
XNOR2_X1 U993 ( .A(n1105), .B(n1277), .ZN(n1143) );
XOR2_X1 U994 ( .A(G131), .B(n1278), .Z(n1277) );
NOR2_X1 U995 ( .A1(G137), .A2(KEYINPUT9), .ZN(n1278) );
NAND2_X1 U996 ( .A1(n1279), .A2(G210), .ZN(n1141) );
NOR2_X1 U997 ( .A1(n1075), .A2(n1209), .ZN(n1042) );
XOR2_X1 U998 ( .A(n1280), .B(n1079), .Z(n1209) );
INV_X1 U999 ( .A(G475), .ZN(n1079) );
NAND2_X1 U1000 ( .A1(n1081), .A2(n1240), .ZN(n1280) );
XNOR2_X1 U1001 ( .A(n1281), .B(n1282), .ZN(n1081) );
XOR2_X1 U1002 ( .A(n1261), .B(n1283), .Z(n1282) );
XOR2_X1 U1003 ( .A(n1284), .B(n1285), .Z(n1283) );
NOR2_X1 U1004 ( .A1(KEYINPUT5), .A2(n1286), .ZN(n1285) );
XOR2_X1 U1005 ( .A(KEYINPUT58), .B(n1287), .Z(n1286) );
NOR2_X1 U1006 ( .A1(n1288), .A2(n1289), .ZN(n1284) );
XOR2_X1 U1007 ( .A(n1290), .B(KEYINPUT10), .Z(n1289) );
NAND2_X1 U1008 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XNOR2_X1 U1009 ( .A(G131), .B(n1293), .ZN(n1292) );
XNOR2_X1 U1010 ( .A(KEYINPUT35), .B(KEYINPUT14), .ZN(n1293) );
NOR2_X1 U1011 ( .A1(G131), .A2(n1291), .ZN(n1288) );
XNOR2_X1 U1012 ( .A(n1294), .B(n1207), .ZN(n1291) );
INV_X1 U1013 ( .A(G143), .ZN(n1207) );
NAND2_X1 U1014 ( .A1(n1279), .A2(G214), .ZN(n1294) );
NOR2_X1 U1015 ( .A1(G953), .A2(G237), .ZN(n1279) );
XOR2_X1 U1016 ( .A(G104), .B(KEYINPUT25), .Z(n1261) );
XNOR2_X1 U1017 ( .A(G113), .B(n1295), .ZN(n1281) );
XOR2_X1 U1018 ( .A(G146), .B(G122), .Z(n1295) );
XOR2_X1 U1019 ( .A(n1296), .B(n1130), .Z(n1075) );
INV_X1 U1020 ( .A(G478), .ZN(n1130) );
OR2_X1 U1021 ( .A1(n1129), .A2(G902), .ZN(n1296) );
XNOR2_X1 U1022 ( .A(n1297), .B(n1298), .ZN(n1129) );
NOR2_X1 U1023 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
XOR2_X1 U1024 ( .A(n1301), .B(KEYINPUT31), .Z(n1300) );
NAND3_X1 U1025 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1301) );
XNOR2_X1 U1026 ( .A(KEYINPUT19), .B(n1305), .ZN(n1304) );
NOR2_X1 U1027 ( .A1(n1306), .A2(n1307), .ZN(n1299) );
XOR2_X1 U1028 ( .A(KEYINPUT8), .B(n1302), .Z(n1307) );
XOR2_X1 U1029 ( .A(n1105), .B(n1308), .Z(n1302) );
NOR2_X1 U1030 ( .A1(KEYINPUT11), .A2(n1309), .ZN(n1308) );
XNOR2_X1 U1031 ( .A(G143), .B(G128), .ZN(n1309) );
XOR2_X1 U1032 ( .A(G134), .B(KEYINPUT41), .Z(n1105) );
NOR2_X1 U1033 ( .A1(n1310), .A2(n1311), .ZN(n1306) );
XOR2_X1 U1034 ( .A(n1305), .B(KEYINPUT19), .Z(n1311) );
NAND2_X1 U1035 ( .A1(n1312), .A2(n1313), .ZN(n1305) );
XNOR2_X1 U1036 ( .A(G116), .B(G122), .ZN(n1312) );
INV_X1 U1037 ( .A(n1303), .ZN(n1310) );
NAND2_X1 U1038 ( .A1(n1314), .A2(n1315), .ZN(n1303) );
XNOR2_X1 U1039 ( .A(KEYINPUT36), .B(n1313), .ZN(n1315) );
INV_X1 U1040 ( .A(G107), .ZN(n1313) );
XOR2_X1 U1041 ( .A(G122), .B(G116), .Z(n1314) );
NAND2_X1 U1042 ( .A1(G217), .A2(n1316), .ZN(n1297) );
INV_X1 U1043 ( .A(n1213), .ZN(n1066) );
XOR2_X1 U1044 ( .A(n1074), .B(KEYINPUT27), .Z(n1213) );
XNOR2_X1 U1045 ( .A(n1317), .B(n1318), .ZN(n1074) );
AND2_X1 U1046 ( .A1(n1237), .A2(G217), .ZN(n1318) );
NAND2_X1 U1047 ( .A1(G234), .A2(n1240), .ZN(n1237) );
NAND2_X1 U1048 ( .A1(n1240), .A2(n1123), .ZN(n1317) );
NAND2_X1 U1049 ( .A1(n1319), .A2(n1320), .ZN(n1123) );
OR2_X1 U1050 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
XOR2_X1 U1051 ( .A(n1323), .B(KEYINPUT22), .Z(n1319) );
NAND2_X1 U1052 ( .A1(n1322), .A2(n1321), .ZN(n1323) );
XNOR2_X1 U1053 ( .A(n1324), .B(n1325), .ZN(n1321) );
XNOR2_X1 U1054 ( .A(KEYINPUT13), .B(n1106), .ZN(n1325) );
INV_X1 U1055 ( .A(G137), .ZN(n1106) );
NAND2_X1 U1056 ( .A1(n1316), .A2(G221), .ZN(n1324) );
AND2_X1 U1057 ( .A1(G234), .A2(n1045), .ZN(n1316) );
INV_X1 U1058 ( .A(G953), .ZN(n1045) );
XNOR2_X1 U1059 ( .A(n1326), .B(n1287), .ZN(n1322) );
XNOR2_X1 U1060 ( .A(n1095), .B(G125), .ZN(n1287) );
INV_X1 U1061 ( .A(G140), .ZN(n1095) );
XOR2_X1 U1062 ( .A(n1327), .B(G146), .Z(n1326) );
NAND2_X1 U1063 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
NAND2_X1 U1064 ( .A1(n1330), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1065 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
NAND2_X1 U1066 ( .A1(G110), .A2(n1334), .ZN(n1333) );
INV_X1 U1067 ( .A(KEYINPUT1), .ZN(n1332) );
NAND2_X1 U1068 ( .A1(n1335), .A2(n1336), .ZN(n1328) );
INV_X1 U1069 ( .A(G110), .ZN(n1336) );
NAND2_X1 U1070 ( .A1(n1334), .A2(n1337), .ZN(n1335) );
OR2_X1 U1071 ( .A1(n1330), .A2(KEYINPUT1), .ZN(n1337) );
XOR2_X1 U1072 ( .A(G119), .B(n1215), .Z(n1330) );
INV_X1 U1073 ( .A(G128), .ZN(n1215) );
INV_X1 U1074 ( .A(KEYINPUT47), .ZN(n1334) );
INV_X1 U1075 ( .A(G902), .ZN(n1240) );
endmodule


