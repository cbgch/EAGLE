//Key = 1110000000000001110000111011111110100010111011011101110100101101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269;

XNOR2_X1 U693 ( .A(G107), .B(n966), .ZN(G9) );
NOR2_X1 U694 ( .A1(n967), .A2(n968), .ZN(G75) );
NOR4_X1 U695 ( .A1(G953), .A2(n969), .A3(n970), .A4(n971), .ZN(n968) );
NOR2_X1 U696 ( .A1(n972), .A2(n973), .ZN(n970) );
NOR2_X1 U697 ( .A1(n974), .A2(n975), .ZN(n972) );
NOR4_X1 U698 ( .A1(n976), .A2(n977), .A3(n978), .A4(n979), .ZN(n975) );
NOR3_X1 U699 ( .A1(n980), .A2(n981), .A3(n982), .ZN(n977) );
NOR2_X1 U700 ( .A1(n983), .A2(n984), .ZN(n982) );
NOR2_X1 U701 ( .A1(n985), .A2(n986), .ZN(n983) );
NOR2_X1 U702 ( .A1(n987), .A2(n988), .ZN(n985) );
NOR2_X1 U703 ( .A1(n989), .A2(n990), .ZN(n981) );
NOR2_X1 U704 ( .A1(n991), .A2(n992), .ZN(n989) );
NOR2_X1 U705 ( .A1(n993), .A2(n994), .ZN(n976) );
NOR2_X1 U706 ( .A1(n995), .A2(n990), .ZN(n993) );
XNOR2_X1 U707 ( .A(n996), .B(KEYINPUT3), .ZN(n995) );
NOR3_X1 U708 ( .A1(n997), .A2(n980), .A3(n984), .ZN(n974) );
INV_X1 U709 ( .A(n996), .ZN(n984) );
NAND3_X1 U710 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
NAND2_X1 U711 ( .A1(n979), .A2(n978), .ZN(n999) );
INV_X1 U712 ( .A(n1001), .ZN(n978) );
OR3_X1 U713 ( .A1(n1002), .A2(n1003), .A3(n979), .ZN(n998) );
NOR3_X1 U714 ( .A1(n969), .A2(G953), .A3(G952), .ZN(n967) );
AND4_X1 U715 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n969) );
NOR4_X1 U716 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1007) );
XNOR2_X1 U717 ( .A(n1012), .B(n1013), .ZN(n1011) );
NOR2_X1 U718 ( .A1(KEYINPUT33), .A2(n1014), .ZN(n1013) );
NOR3_X1 U719 ( .A1(n1015), .A2(n980), .A3(n1016), .ZN(n1006) );
NAND2_X1 U720 ( .A1(n1017), .A2(n1018), .ZN(n1005) );
XOR2_X1 U721 ( .A(KEYINPUT5), .B(n1019), .Z(n1017) );
XOR2_X1 U722 ( .A(n1020), .B(n1021), .Z(n1004) );
NAND2_X1 U723 ( .A1(KEYINPUT27), .A2(n1022), .ZN(n1021) );
XOR2_X1 U724 ( .A(n1023), .B(n1024), .Z(G72) );
NOR2_X1 U725 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
AND2_X1 U726 ( .A1(G227), .A2(G900), .ZN(n1025) );
NOR2_X1 U727 ( .A1(KEYINPUT50), .A2(n1027), .ZN(n1023) );
NOR2_X1 U728 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
XOR2_X1 U729 ( .A(KEYINPUT59), .B(n1030), .Z(n1029) );
AND2_X1 U730 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR3_X1 U731 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1028) );
NOR2_X1 U732 ( .A1(n1034), .A2(G953), .ZN(n1032) );
XNOR2_X1 U733 ( .A(n1035), .B(n1036), .ZN(n1031) );
XOR2_X1 U734 ( .A(n1037), .B(n1038), .Z(n1036) );
XOR2_X1 U735 ( .A(KEYINPUT30), .B(KEYINPUT21), .Z(n1038) );
XOR2_X1 U736 ( .A(n1039), .B(n1040), .Z(n1035) );
XOR2_X1 U737 ( .A(n1041), .B(n1042), .Z(G69) );
XOR2_X1 U738 ( .A(n1043), .B(n1044), .Z(n1042) );
NOR2_X1 U739 ( .A1(n1045), .A2(n1026), .ZN(n1044) );
AND2_X1 U740 ( .A1(G224), .A2(G898), .ZN(n1045) );
NAND2_X1 U741 ( .A1(n1046), .A2(n1047), .ZN(n1043) );
NAND2_X1 U742 ( .A1(G953), .A2(n1048), .ZN(n1047) );
XNOR2_X1 U743 ( .A(n1049), .B(KEYINPUT14), .ZN(n1046) );
NAND2_X1 U744 ( .A1(n1026), .A2(n1050), .ZN(n1041) );
NAND2_X1 U745 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U746 ( .A1(n1053), .A2(n1054), .ZN(G66) );
XOR2_X1 U747 ( .A(n1055), .B(n1056), .Z(n1054) );
XNOR2_X1 U748 ( .A(KEYINPUT46), .B(n1057), .ZN(n1055) );
NOR3_X1 U749 ( .A1(n1058), .A2(KEYINPUT25), .A3(n1059), .ZN(n1057) );
INV_X1 U750 ( .A(G217), .ZN(n1059) );
NOR2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(G63) );
XOR2_X1 U752 ( .A(n1062), .B(n1063), .Z(n1061) );
NOR2_X1 U753 ( .A1(n1064), .A2(n1058), .ZN(n1062) );
XNOR2_X1 U754 ( .A(n1053), .B(KEYINPUT2), .ZN(n1060) );
NOR2_X1 U755 ( .A1(n1053), .A2(n1065), .ZN(G60) );
XOR2_X1 U756 ( .A(n1066), .B(n1067), .Z(n1065) );
NOR2_X1 U757 ( .A1(n1068), .A2(n1058), .ZN(n1066) );
XNOR2_X1 U758 ( .A(G104), .B(n1069), .ZN(G6) );
NOR3_X1 U759 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(G57) );
AND2_X1 U760 ( .A1(KEYINPUT26), .A2(n1053), .ZN(n1072) );
NOR3_X1 U761 ( .A1(KEYINPUT26), .A2(n1073), .A3(n1026), .ZN(n1071) );
NOR2_X1 U762 ( .A1(n1074), .A2(n1075), .ZN(n1070) );
XOR2_X1 U763 ( .A(n1076), .B(KEYINPUT29), .Z(n1075) );
NAND2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U765 ( .A1(n1078), .A2(n1077), .ZN(n1074) );
XOR2_X1 U766 ( .A(n1079), .B(n1080), .Z(n1077) );
XNOR2_X1 U767 ( .A(n1081), .B(n1082), .ZN(n1080) );
NOR2_X1 U768 ( .A1(n1022), .A2(n1058), .ZN(n1081) );
INV_X1 U769 ( .A(G472), .ZN(n1022) );
XNOR2_X1 U770 ( .A(n1083), .B(n1084), .ZN(n1079) );
NOR2_X1 U771 ( .A1(n1053), .A2(n1085), .ZN(G54) );
XOR2_X1 U772 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U773 ( .A1(n1014), .A2(n1058), .ZN(n1087) );
NAND2_X1 U774 ( .A1(G902), .A2(n971), .ZN(n1058) );
NOR2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
XOR2_X1 U776 ( .A(KEYINPUT12), .B(n1090), .Z(n1089) );
NOR2_X1 U777 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
AND2_X1 U778 ( .A1(n1092), .A2(n1091), .ZN(n1088) );
XOR2_X1 U779 ( .A(n1093), .B(n1094), .Z(n1091) );
XNOR2_X1 U780 ( .A(KEYINPUT7), .B(n1095), .ZN(n1094) );
XOR2_X1 U781 ( .A(n1096), .B(n1082), .Z(n1092) );
NOR2_X1 U782 ( .A1(n1053), .A2(n1097), .ZN(G51) );
XOR2_X1 U783 ( .A(n1098), .B(n1099), .Z(n1097) );
XNOR2_X1 U784 ( .A(n1100), .B(n1049), .ZN(n1099) );
XNOR2_X1 U785 ( .A(n1101), .B(n1083), .ZN(n1098) );
NAND3_X1 U786 ( .A1(G902), .A2(n1102), .A3(n1103), .ZN(n1101) );
XOR2_X1 U787 ( .A(n971), .B(KEYINPUT13), .Z(n1103) );
NAND3_X1 U788 ( .A1(n1051), .A2(n1034), .A3(n1104), .ZN(n971) );
XOR2_X1 U789 ( .A(n1052), .B(KEYINPUT36), .Z(n1104) );
AND4_X1 U790 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1034) );
NOR4_X1 U791 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
INV_X1 U792 ( .A(n1113), .ZN(n1112) );
NOR3_X1 U793 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1109) );
NOR2_X1 U794 ( .A1(KEYINPUT47), .A2(n1117), .ZN(n1116) );
NOR2_X1 U795 ( .A1(n1000), .A2(n1118), .ZN(n1117) );
NOR2_X1 U796 ( .A1(n1119), .A2(n1120), .ZN(n1115) );
INV_X1 U797 ( .A(KEYINPUT47), .ZN(n1120) );
NOR3_X1 U798 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1107) );
NOR3_X1 U799 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1123) );
INV_X1 U800 ( .A(KEYINPUT6), .ZN(n1124) );
NOR2_X1 U801 ( .A1(KEYINPUT6), .A2(n1127), .ZN(n1122) );
AND3_X1 U802 ( .A1(n1128), .A2(n1001), .A3(n1119), .ZN(n1121) );
AND4_X1 U803 ( .A1(n1129), .A2(n1130), .A3(n1069), .A4(n1131), .ZN(n1051) );
AND4_X1 U804 ( .A1(n966), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1131) );
NAND3_X1 U805 ( .A1(n996), .A2(n1002), .A3(n1135), .ZN(n966) );
NAND3_X1 U806 ( .A1(n1135), .A2(n996), .A3(n1003), .ZN(n1069) );
NOR2_X1 U807 ( .A1(n1026), .A2(G952), .ZN(n1053) );
XNOR2_X1 U808 ( .A(G146), .B(n1105), .ZN(G48) );
NAND4_X1 U809 ( .A1(n1128), .A2(n1136), .A3(n1003), .A4(n986), .ZN(n1105) );
XNOR2_X1 U810 ( .A(G143), .B(n1106), .ZN(G45) );
NAND4_X1 U811 ( .A1(n1136), .A2(n1137), .A3(n992), .A4(n986), .ZN(n1106) );
XNOR2_X1 U812 ( .A(G140), .B(n1113), .ZN(G42) );
NAND3_X1 U813 ( .A1(n1003), .A2(n991), .A3(n1119), .ZN(n1113) );
XNOR2_X1 U814 ( .A(G137), .B(n1138), .ZN(G39) );
NAND3_X1 U815 ( .A1(n1001), .A2(n1139), .A3(n1119), .ZN(n1138) );
XOR2_X1 U816 ( .A(KEYINPUT57), .B(n1128), .Z(n1139) );
XNOR2_X1 U817 ( .A(G134), .B(n1140), .ZN(G36) );
NAND2_X1 U818 ( .A1(n1119), .A2(n1141), .ZN(n1140) );
NAND2_X1 U819 ( .A1(n1142), .A2(n1143), .ZN(G33) );
NAND2_X1 U820 ( .A1(n1111), .A2(n1144), .ZN(n1143) );
XOR2_X1 U821 ( .A(KEYINPUT52), .B(n1145), .Z(n1142) );
NOR2_X1 U822 ( .A1(n1111), .A2(n1144), .ZN(n1145) );
AND3_X1 U823 ( .A1(n1003), .A2(n992), .A3(n1119), .ZN(n1111) );
NOR2_X1 U824 ( .A1(n990), .A2(n1118), .ZN(n1119) );
INV_X1 U825 ( .A(n1136), .ZN(n1118) );
INV_X1 U826 ( .A(n1000), .ZN(n990) );
NOR2_X1 U827 ( .A1(n987), .A2(n1016), .ZN(n1000) );
XOR2_X1 U828 ( .A(n1127), .B(n1146), .Z(G30) );
NAND2_X1 U829 ( .A1(KEYINPUT16), .A2(G128), .ZN(n1146) );
NAND2_X1 U830 ( .A1(n1125), .A2(n986), .ZN(n1127) );
AND3_X1 U831 ( .A1(n1136), .A2(n1002), .A3(n1128), .ZN(n1125) );
NOR3_X1 U832 ( .A1(n980), .A2(n1147), .A3(n1148), .ZN(n1136) );
XNOR2_X1 U833 ( .A(G101), .B(n1129), .ZN(G3) );
NAND3_X1 U834 ( .A1(n1001), .A2(n1135), .A3(n992), .ZN(n1129) );
XNOR2_X1 U835 ( .A(n1110), .B(n1149), .ZN(G27) );
NAND2_X1 U836 ( .A1(KEYINPUT32), .A2(G125), .ZN(n1149) );
AND4_X1 U837 ( .A1(n1148), .A2(n991), .A3(n1003), .A4(n1150), .ZN(n1110) );
NOR3_X1 U838 ( .A1(n1126), .A2(n1147), .A3(n980), .ZN(n1150) );
INV_X1 U839 ( .A(n994), .ZN(n980) );
AND2_X1 U840 ( .A1(n1151), .A2(n973), .ZN(n1147) );
NAND3_X1 U841 ( .A1(n1033), .A2(G902), .A3(n1152), .ZN(n1151) );
XOR2_X1 U842 ( .A(n1153), .B(KEYINPUT9), .Z(n1152) );
NOR2_X1 U843 ( .A1(n1026), .A2(G900), .ZN(n1033) );
INV_X1 U844 ( .A(n986), .ZN(n1126) );
XNOR2_X1 U845 ( .A(G122), .B(n1130), .ZN(G24) );
NAND3_X1 U846 ( .A1(n1154), .A2(n996), .A3(n1137), .ZN(n1130) );
AND2_X1 U847 ( .A1(n1155), .A2(n1156), .ZN(n1137) );
XNOR2_X1 U848 ( .A(n1010), .B(KEYINPUT44), .ZN(n1155) );
NOR2_X1 U849 ( .A1(n1157), .A2(n1158), .ZN(n996) );
XNOR2_X1 U850 ( .A(n1052), .B(n1159), .ZN(G21) );
NOR2_X1 U851 ( .A1(KEYINPUT20), .A2(n1160), .ZN(n1159) );
NAND3_X1 U852 ( .A1(n1154), .A2(n1001), .A3(n1128), .ZN(n1052) );
AND2_X1 U853 ( .A1(n1157), .A2(n1158), .ZN(n1128) );
INV_X1 U854 ( .A(n1161), .ZN(n1158) );
XNOR2_X1 U855 ( .A(G116), .B(n1134), .ZN(G18) );
NAND2_X1 U856 ( .A1(n1141), .A2(n1154), .ZN(n1134) );
INV_X1 U857 ( .A(n1114), .ZN(n1141) );
NAND2_X1 U858 ( .A1(n992), .A2(n1002), .ZN(n1114) );
NOR2_X1 U859 ( .A1(n1008), .A2(n1162), .ZN(n1002) );
XNOR2_X1 U860 ( .A(G113), .B(n1133), .ZN(G15) );
NAND3_X1 U861 ( .A1(n1003), .A2(n992), .A3(n1154), .ZN(n1133) );
AND3_X1 U862 ( .A1(n1163), .A2(n994), .A3(n1148), .ZN(n1154) );
INV_X1 U863 ( .A(n979), .ZN(n1148) );
AND2_X1 U864 ( .A1(n1161), .A2(n1157), .ZN(n992) );
AND2_X1 U865 ( .A1(n1164), .A2(n1156), .ZN(n1003) );
XNOR2_X1 U866 ( .A(n1008), .B(KEYINPUT55), .ZN(n1156) );
XNOR2_X1 U867 ( .A(n1010), .B(KEYINPUT56), .ZN(n1164) );
XNOR2_X1 U868 ( .A(G110), .B(n1132), .ZN(G12) );
NAND3_X1 U869 ( .A1(n991), .A2(n1135), .A3(n1001), .ZN(n1132) );
NOR2_X1 U870 ( .A1(n1165), .A2(n1008), .ZN(n1001) );
XOR2_X1 U871 ( .A(n1166), .B(n1068), .Z(n1008) );
INV_X1 U872 ( .A(G475), .ZN(n1068) );
OR2_X1 U873 ( .A1(n1067), .A2(G902), .ZN(n1166) );
XOR2_X1 U874 ( .A(n1167), .B(n1168), .Z(n1067) );
XNOR2_X1 U875 ( .A(G104), .B(n1169), .ZN(n1168) );
NAND3_X1 U876 ( .A1(n1170), .A2(n1171), .A3(KEYINPUT28), .ZN(n1169) );
NAND3_X1 U877 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
INV_X1 U878 ( .A(KEYINPUT0), .ZN(n1174) );
NAND2_X1 U879 ( .A1(n1175), .A2(KEYINPUT0), .ZN(n1170) );
XNOR2_X1 U880 ( .A(n1176), .B(n1173), .ZN(n1175) );
XOR2_X1 U881 ( .A(n1177), .B(n1178), .Z(n1173) );
XNOR2_X1 U882 ( .A(n1179), .B(n1180), .ZN(n1178) );
NOR2_X1 U883 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
INV_X1 U884 ( .A(G214), .ZN(n1181) );
NAND2_X1 U885 ( .A1(KEYINPUT60), .A2(n1144), .ZN(n1177) );
INV_X1 U886 ( .A(G131), .ZN(n1144) );
NOR2_X1 U887 ( .A1(KEYINPUT19), .A2(n1172), .ZN(n1176) );
XNOR2_X1 U888 ( .A(n1183), .B(n1184), .ZN(n1172) );
NAND2_X1 U889 ( .A1(KEYINPUT41), .A2(n1185), .ZN(n1183) );
XNOR2_X1 U890 ( .A(n1162), .B(KEYINPUT56), .ZN(n1165) );
INV_X1 U891 ( .A(n1010), .ZN(n1162) );
XOR2_X1 U892 ( .A(n1186), .B(n1064), .Z(n1010) );
INV_X1 U893 ( .A(G478), .ZN(n1064) );
OR2_X1 U894 ( .A1(n1063), .A2(G902), .ZN(n1186) );
XNOR2_X1 U895 ( .A(n1187), .B(n1188), .ZN(n1063) );
XNOR2_X1 U896 ( .A(n1189), .B(n1190), .ZN(n1188) );
NOR2_X1 U897 ( .A1(G116), .A2(KEYINPUT10), .ZN(n1190) );
NAND2_X1 U898 ( .A1(n1191), .A2(KEYINPUT53), .ZN(n1189) );
XNOR2_X1 U899 ( .A(G134), .B(n1192), .ZN(n1191) );
XOR2_X1 U900 ( .A(n1193), .B(n1194), .Z(n1187) );
XOR2_X1 U901 ( .A(G122), .B(n1195), .Z(n1194) );
AND3_X1 U902 ( .A1(G217), .A2(n1026), .A3(G234), .ZN(n1195) );
NAND2_X1 U903 ( .A1(KEYINPUT49), .A2(n1196), .ZN(n1193) );
AND3_X1 U904 ( .A1(n979), .A2(n994), .A3(n1163), .ZN(n1135) );
AND2_X1 U905 ( .A1(n986), .A2(n1197), .ZN(n1163) );
NAND2_X1 U906 ( .A1(n1198), .A2(n973), .ZN(n1197) );
NAND3_X1 U907 ( .A1(n1153), .A2(n1026), .A3(n1199), .ZN(n973) );
XNOR2_X1 U908 ( .A(KEYINPUT4), .B(n1073), .ZN(n1199) );
INV_X1 U909 ( .A(G952), .ZN(n1073) );
NAND4_X1 U910 ( .A1(G953), .A2(G902), .A3(n1153), .A4(n1048), .ZN(n1198) );
INV_X1 U911 ( .A(G898), .ZN(n1048) );
NAND2_X1 U912 ( .A1(G237), .A2(G234), .ZN(n1153) );
NOR2_X1 U913 ( .A1(n1200), .A2(n1016), .ZN(n986) );
INV_X1 U914 ( .A(n988), .ZN(n1016) );
NAND2_X1 U915 ( .A1(G214), .A2(n1201), .ZN(n988) );
INV_X1 U916 ( .A(n987), .ZN(n1200) );
XOR2_X1 U917 ( .A(n1009), .B(KEYINPUT43), .Z(n987) );
XNOR2_X1 U918 ( .A(n1202), .B(n1102), .ZN(n1009) );
AND2_X1 U919 ( .A1(G210), .A2(n1201), .ZN(n1102) );
NAND2_X1 U920 ( .A1(n1203), .A2(n1204), .ZN(n1201) );
NAND2_X1 U921 ( .A1(n1205), .A2(n1204), .ZN(n1202) );
XNOR2_X1 U922 ( .A(n1049), .B(n1206), .ZN(n1205) );
NOR2_X1 U923 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR2_X1 U924 ( .A1(n1083), .A2(n1209), .ZN(n1208) );
XOR2_X1 U925 ( .A(n1100), .B(KEYINPUT1), .Z(n1209) );
NOR2_X1 U926 ( .A1(n1210), .A2(n1100), .ZN(n1207) );
XOR2_X1 U927 ( .A(n1211), .B(n1212), .Z(n1100) );
NAND2_X1 U928 ( .A1(G224), .A2(n1026), .ZN(n1211) );
XNOR2_X1 U929 ( .A(n1213), .B(n1214), .ZN(n1049) );
XOR2_X1 U930 ( .A(n1167), .B(n1215), .Z(n1214) );
XOR2_X1 U931 ( .A(G113), .B(G122), .Z(n1167) );
XOR2_X1 U932 ( .A(n1216), .B(n1217), .Z(n1213) );
NOR2_X1 U933 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
XOR2_X1 U934 ( .A(KEYINPUT18), .B(n1220), .Z(n1219) );
NOR2_X1 U935 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
AND2_X1 U936 ( .A1(n1222), .A2(n1221), .ZN(n1218) );
XOR2_X1 U937 ( .A(G101), .B(KEYINPUT37), .Z(n1222) );
XNOR2_X1 U938 ( .A(G110), .B(KEYINPUT35), .ZN(n1216) );
NAND2_X1 U939 ( .A1(G221), .A2(n1223), .ZN(n994) );
XOR2_X1 U940 ( .A(n1012), .B(n1014), .Z(n979) );
INV_X1 U941 ( .A(G469), .ZN(n1014) );
NAND2_X1 U942 ( .A1(n1224), .A2(n1204), .ZN(n1012) );
XNOR2_X1 U943 ( .A(n1225), .B(n1226), .ZN(n1224) );
XNOR2_X1 U944 ( .A(n1227), .B(n1228), .ZN(n1226) );
NAND2_X1 U945 ( .A1(KEYINPUT58), .A2(n1096), .ZN(n1228) );
XOR2_X1 U946 ( .A(n1229), .B(n1221), .Z(n1096) );
XNOR2_X1 U947 ( .A(G104), .B(n1196), .ZN(n1221) );
INV_X1 U948 ( .A(G107), .ZN(n1196) );
XOR2_X1 U949 ( .A(n1039), .B(G101), .Z(n1229) );
XNOR2_X1 U950 ( .A(G146), .B(n1192), .ZN(n1039) );
XOR2_X1 U951 ( .A(G128), .B(G143), .Z(n1192) );
NAND2_X1 U952 ( .A1(KEYINPUT38), .A2(n1230), .ZN(n1227) );
XOR2_X1 U953 ( .A(n1231), .B(n1093), .Z(n1230) );
XOR2_X1 U954 ( .A(n1232), .B(n1233), .Z(n1093) );
XNOR2_X1 U955 ( .A(KEYINPUT15), .B(n1234), .ZN(n1233) );
INV_X1 U956 ( .A(G140), .ZN(n1234) );
NAND2_X1 U957 ( .A1(G227), .A2(n1026), .ZN(n1232) );
NAND2_X1 U958 ( .A1(KEYINPUT17), .A2(n1235), .ZN(n1231) );
XNOR2_X1 U959 ( .A(KEYINPUT31), .B(n1095), .ZN(n1235) );
NOR2_X1 U960 ( .A1(n1157), .A2(n1161), .ZN(n991) );
NOR2_X1 U961 ( .A1(n1015), .A2(n1236), .ZN(n1161) );
AND2_X1 U962 ( .A1(n1019), .A2(n1018), .ZN(n1236) );
NOR2_X1 U963 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
AND2_X1 U964 ( .A1(n1237), .A2(G217), .ZN(n1019) );
XOR2_X1 U965 ( .A(n1223), .B(KEYINPUT8), .Z(n1237) );
NAND2_X1 U966 ( .A1(G234), .A2(n1204), .ZN(n1223) );
NAND2_X1 U967 ( .A1(n1056), .A2(n1204), .ZN(n1018) );
XNOR2_X1 U968 ( .A(n1238), .B(n1239), .ZN(n1056) );
XOR2_X1 U969 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U970 ( .A(n1242), .B(n1095), .ZN(n1241) );
INV_X1 U971 ( .A(G110), .ZN(n1095) );
NAND2_X1 U972 ( .A1(KEYINPUT63), .A2(n1184), .ZN(n1242) );
XNOR2_X1 U973 ( .A(G137), .B(KEYINPUT11), .ZN(n1240) );
XOR2_X1 U974 ( .A(n1185), .B(n1243), .Z(n1238) );
XOR2_X1 U975 ( .A(n1244), .B(n1245), .Z(n1243) );
NAND3_X1 U976 ( .A1(G234), .A2(n1026), .A3(G221), .ZN(n1245) );
NAND2_X1 U977 ( .A1(n1246), .A2(KEYINPUT51), .ZN(n1244) );
XNOR2_X1 U978 ( .A(G119), .B(G128), .ZN(n1246) );
XNOR2_X1 U979 ( .A(n1037), .B(KEYINPUT22), .ZN(n1185) );
XOR2_X1 U980 ( .A(G140), .B(n1212), .Z(n1037) );
XOR2_X1 U981 ( .A(G125), .B(KEYINPUT48), .Z(n1212) );
NAND3_X1 U982 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1157) );
NAND2_X1 U983 ( .A1(KEYINPUT62), .A2(n1020), .ZN(n1249) );
OR3_X1 U984 ( .A1(n1020), .A2(KEYINPUT62), .A3(n1250), .ZN(n1248) );
NAND2_X1 U985 ( .A1(n1250), .A2(n1251), .ZN(n1247) );
NAND2_X1 U986 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U987 ( .A(KEYINPUT62), .ZN(n1253) );
XNOR2_X1 U988 ( .A(KEYINPUT39), .B(n1020), .ZN(n1252) );
NAND2_X1 U989 ( .A1(n1254), .A2(n1204), .ZN(n1020) );
INV_X1 U990 ( .A(G902), .ZN(n1204) );
XOR2_X1 U991 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U992 ( .A(n1257), .B(KEYINPUT23), .ZN(n1256) );
NAND2_X1 U993 ( .A1(n1258), .A2(KEYINPUT61), .ZN(n1257) );
XNOR2_X1 U994 ( .A(n1259), .B(n1082), .ZN(n1258) );
INV_X1 U995 ( .A(n1225), .ZN(n1082) );
XOR2_X1 U996 ( .A(n1040), .B(KEYINPUT40), .Z(n1225) );
XOR2_X1 U997 ( .A(G131), .B(n1260), .Z(n1040) );
XOR2_X1 U998 ( .A(G137), .B(G134), .Z(n1260) );
NAND2_X1 U999 ( .A1(KEYINPUT45), .A2(n1210), .ZN(n1259) );
INV_X1 U1000 ( .A(n1083), .ZN(n1210) );
XOR2_X1 U1001 ( .A(G128), .B(n1261), .Z(n1083) );
NOR2_X1 U1002 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NOR3_X1 U1003 ( .A1(KEYINPUT34), .A2(G146), .A3(n1179), .ZN(n1263) );
INV_X1 U1004 ( .A(G143), .ZN(n1179) );
NOR2_X1 U1005 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
INV_X1 U1006 ( .A(KEYINPUT34), .ZN(n1265) );
XNOR2_X1 U1007 ( .A(n1184), .B(G143), .ZN(n1264) );
INV_X1 U1008 ( .A(G146), .ZN(n1184) );
XNOR2_X1 U1009 ( .A(n1084), .B(n1078), .ZN(n1255) );
XOR2_X1 U1010 ( .A(G101), .B(n1266), .Z(n1078) );
NOR2_X1 U1011 ( .A1(n1267), .A2(n1182), .ZN(n1266) );
NAND2_X1 U1012 ( .A1(n1268), .A2(n1026), .ZN(n1182) );
INV_X1 U1013 ( .A(G953), .ZN(n1026) );
XNOR2_X1 U1014 ( .A(KEYINPUT24), .B(n1203), .ZN(n1268) );
INV_X1 U1015 ( .A(G237), .ZN(n1203) );
INV_X1 U1016 ( .A(G210), .ZN(n1267) );
XNOR2_X1 U1017 ( .A(n1269), .B(n1215), .ZN(n1084) );
XNOR2_X1 U1018 ( .A(G116), .B(n1160), .ZN(n1215) );
INV_X1 U1019 ( .A(G119), .ZN(n1160) );
XNOR2_X1 U1020 ( .A(G113), .B(KEYINPUT42), .ZN(n1269) );
XOR2_X1 U1021 ( .A(G472), .B(KEYINPUT54), .Z(n1250) );
endmodule


