//Key = 0010110000100000101100100010110001011000101001001100010000001001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395;

XOR2_X1 U749 ( .A(G107), .B(n1039), .Z(G9) );
NOR3_X1 U750 ( .A1(n1040), .A2(KEYINPUT31), .A3(n1041), .ZN(n1039) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR4_X1 U752 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043) );
NAND3_X1 U753 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1044) );
XOR2_X1 U754 ( .A(KEYINPUT37), .B(n1051), .Z(n1050) );
NOR2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U757 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U758 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U761 ( .A1(n1064), .A2(n1065), .ZN(n1056) );
NOR2_X1 U762 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NOR3_X1 U763 ( .A1(n1068), .A2(KEYINPUT51), .A3(n1069), .ZN(n1066) );
NOR3_X1 U764 ( .A1(n1059), .A2(n1070), .A3(n1065), .ZN(n1052) );
NOR4_X1 U765 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1070) );
NOR2_X1 U766 ( .A1(n1055), .A2(n1075), .ZN(n1074) );
INV_X1 U767 ( .A(KEYINPUT51), .ZN(n1075) );
NAND3_X1 U768 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1055) );
NOR3_X1 U769 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1073) );
XNOR2_X1 U770 ( .A(n1078), .B(KEYINPUT38), .ZN(n1080) );
NOR4_X1 U771 ( .A1(n1078), .A2(n1082), .A3(KEYINPUT53), .A4(n1083), .ZN(n1072) );
INV_X1 U772 ( .A(n1084), .ZN(n1078) );
NOR2_X1 U773 ( .A1(n1085), .A2(n1084), .ZN(n1071) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U775 ( .A1(n1081), .A2(n1088), .ZN(n1087) );
NOR2_X1 U776 ( .A1(n1089), .A2(n1083), .ZN(n1086) );
NOR2_X1 U777 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
AND2_X1 U778 ( .A1(n1092), .A2(KEYINPUT53), .ZN(n1090) );
INV_X1 U779 ( .A(n1093), .ZN(n1059) );
NOR3_X1 U780 ( .A1(n1094), .A2(G953), .A3(G952), .ZN(n1042) );
INV_X1 U781 ( .A(n1048), .ZN(n1094) );
NAND4_X1 U782 ( .A1(n1076), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1048) );
NOR4_X1 U783 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XNOR2_X1 U784 ( .A(n1102), .B(n1103), .ZN(n1101) );
NAND2_X1 U785 ( .A1(KEYINPUT45), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U786 ( .A(n1105), .B(n1106), .ZN(n1100) );
NOR2_X1 U787 ( .A1(n1107), .A2(KEYINPUT57), .ZN(n1106) );
XNOR2_X1 U788 ( .A(n1108), .B(n1109), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1110), .B(n1111), .Z(n1095) );
XNOR2_X1 U790 ( .A(G469), .B(KEYINPUT10), .ZN(n1111) );
XOR2_X1 U791 ( .A(n1112), .B(n1113), .Z(G72) );
XOR2_X1 U792 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U793 ( .A1(n1049), .A2(n1116), .ZN(n1115) );
NAND2_X1 U794 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
XNOR2_X1 U795 ( .A(n1119), .B(KEYINPUT33), .ZN(n1117) );
NAND3_X1 U796 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1114) );
XOR2_X1 U797 ( .A(n1123), .B(KEYINPUT13), .Z(n1122) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U799 ( .A1(n1126), .A2(G953), .ZN(n1121) );
OR2_X1 U800 ( .A1(n1125), .A2(n1124), .ZN(n1120) );
XNOR2_X1 U801 ( .A(n1127), .B(n1128), .ZN(n1124) );
NOR2_X1 U802 ( .A1(KEYINPUT55), .A2(n1129), .ZN(n1128) );
XNOR2_X1 U803 ( .A(G125), .B(KEYINPUT44), .ZN(n1127) );
XNOR2_X1 U804 ( .A(n1130), .B(n1131), .ZN(n1125) );
XNOR2_X1 U805 ( .A(G137), .B(n1132), .ZN(n1131) );
NAND2_X1 U806 ( .A1(KEYINPUT22), .A2(n1133), .ZN(n1132) );
XNOR2_X1 U807 ( .A(n1134), .B(n1135), .ZN(n1130) );
NOR2_X1 U808 ( .A1(n1136), .A2(n1049), .ZN(n1112) );
AND2_X1 U809 ( .A1(G227), .A2(G900), .ZN(n1136) );
NAND2_X1 U810 ( .A1(n1137), .A2(n1138), .ZN(G69) );
NAND2_X1 U811 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U812 ( .A1(G953), .A2(n1141), .ZN(n1140) );
NAND3_X1 U813 ( .A1(G953), .A2(n1142), .A3(n1143), .ZN(n1137) );
INV_X1 U814 ( .A(n1139), .ZN(n1143) );
XNOR2_X1 U815 ( .A(n1144), .B(n1145), .ZN(n1139) );
NOR3_X1 U816 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(n1145) );
NOR2_X1 U817 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
INV_X1 U818 ( .A(KEYINPUT8), .ZN(n1150) );
NOR2_X1 U819 ( .A1(n1151), .A2(n1152), .ZN(n1149) );
NOR2_X1 U820 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
NOR2_X1 U821 ( .A1(n1155), .A2(n1156), .ZN(n1151) );
NOR2_X1 U822 ( .A1(KEYINPUT8), .A2(n1157), .ZN(n1147) );
NOR2_X1 U823 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U824 ( .A1(n1156), .A2(n1154), .ZN(n1159) );
XNOR2_X1 U825 ( .A(n1155), .B(KEYINPUT12), .ZN(n1154) );
INV_X1 U826 ( .A(n1153), .ZN(n1156) );
NOR2_X1 U827 ( .A1(n1153), .A2(n1155), .ZN(n1158) );
NOR2_X1 U828 ( .A1(G898), .A2(n1049), .ZN(n1146) );
NAND3_X1 U829 ( .A1(n1160), .A2(n1161), .A3(n1049), .ZN(n1144) );
NAND2_X1 U830 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
INV_X1 U831 ( .A(KEYINPUT18), .ZN(n1163) );
NAND2_X1 U832 ( .A1(KEYINPUT18), .A2(n1164), .ZN(n1160) );
NAND2_X1 U833 ( .A1(G898), .A2(G224), .ZN(n1142) );
NOR2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(G66) );
NOR3_X1 U835 ( .A1(n1105), .A2(n1167), .A3(n1168), .ZN(n1166) );
NOR3_X1 U836 ( .A1(n1169), .A2(n1170), .A3(n1171), .ZN(n1168) );
NOR2_X1 U837 ( .A1(n1172), .A2(n1173), .ZN(n1167) );
AND2_X1 U838 ( .A1(n1174), .A2(n1107), .ZN(n1172) );
INV_X1 U839 ( .A(n1170), .ZN(n1107) );
NOR2_X1 U840 ( .A1(n1165), .A2(n1175), .ZN(G63) );
XNOR2_X1 U841 ( .A(n1176), .B(n1177), .ZN(n1175) );
XOR2_X1 U842 ( .A(KEYINPUT17), .B(n1178), .Z(n1177) );
NOR2_X1 U843 ( .A1(n1179), .A2(n1171), .ZN(n1178) );
NOR2_X1 U844 ( .A1(n1165), .A2(n1180), .ZN(G60) );
NOR2_X1 U845 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U846 ( .A(KEYINPUT32), .B(n1183), .Z(n1182) );
AND2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1184), .ZN(n1181) );
NOR2_X1 U849 ( .A1(n1171), .A2(n1186), .ZN(n1185) );
INV_X1 U850 ( .A(G475), .ZN(n1186) );
XNOR2_X1 U851 ( .A(n1187), .B(n1188), .ZN(G6) );
NAND2_X1 U852 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
OR3_X1 U853 ( .A1(n1082), .A2(n1041), .A3(KEYINPUT14), .ZN(n1190) );
INV_X1 U854 ( .A(n1191), .ZN(n1041) );
NAND4_X1 U855 ( .A1(n1092), .A2(n1077), .A3(n1192), .A4(KEYINPUT14), .ZN(n1189) );
NOR2_X1 U856 ( .A1(n1067), .A2(n1193), .ZN(n1192) );
NOR2_X1 U857 ( .A1(n1165), .A2(n1194), .ZN(G57) );
XNOR2_X1 U858 ( .A(n1195), .B(n1196), .ZN(n1194) );
XNOR2_X1 U859 ( .A(n1197), .B(n1198), .ZN(n1196) );
NOR2_X1 U860 ( .A1(KEYINPUT56), .A2(n1199), .ZN(n1198) );
XOR2_X1 U861 ( .A(n1200), .B(n1201), .Z(n1199) );
XNOR2_X1 U862 ( .A(n1202), .B(n1203), .ZN(n1201) );
XNOR2_X1 U863 ( .A(n1204), .B(n1205), .ZN(n1200) );
NOR2_X1 U864 ( .A1(KEYINPUT61), .A2(n1206), .ZN(n1205) );
NOR2_X1 U865 ( .A1(n1103), .A2(n1171), .ZN(n1206) );
NAND2_X1 U866 ( .A1(KEYINPUT4), .A2(n1207), .ZN(n1204) );
NOR2_X1 U867 ( .A1(n1165), .A2(n1208), .ZN(G54) );
XOR2_X1 U868 ( .A(n1209), .B(n1210), .Z(n1208) );
NOR2_X1 U869 ( .A1(n1211), .A2(n1171), .ZN(n1210) );
INV_X1 U870 ( .A(G469), .ZN(n1211) );
NOR2_X1 U871 ( .A1(n1212), .A2(n1213), .ZN(n1209) );
XOR2_X1 U872 ( .A(KEYINPUT59), .B(n1214), .Z(n1213) );
NOR2_X1 U873 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NOR2_X1 U874 ( .A1(n1217), .A2(n1218), .ZN(n1212) );
XOR2_X1 U875 ( .A(n1215), .B(KEYINPUT2), .Z(n1218) );
XNOR2_X1 U876 ( .A(n1219), .B(n1220), .ZN(n1215) );
INV_X1 U877 ( .A(n1216), .ZN(n1217) );
XNOR2_X1 U878 ( .A(n1221), .B(n1222), .ZN(n1216) );
NOR2_X1 U879 ( .A1(KEYINPUT15), .A2(n1202), .ZN(n1222) );
NOR2_X1 U880 ( .A1(n1165), .A2(n1223), .ZN(G51) );
XOR2_X1 U881 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U882 ( .A(n1226), .B(n1207), .ZN(n1225) );
XNOR2_X1 U883 ( .A(n1227), .B(n1228), .ZN(n1226) );
NOR2_X1 U884 ( .A1(n1229), .A2(n1171), .ZN(n1228) );
NAND2_X1 U885 ( .A1(G902), .A2(n1174), .ZN(n1171) );
NAND3_X1 U886 ( .A1(n1119), .A2(n1230), .A3(n1118), .ZN(n1174) );
INV_X1 U887 ( .A(n1045), .ZN(n1118) );
NAND4_X1 U888 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1045) );
NOR2_X1 U889 ( .A1(n1235), .A2(n1236), .ZN(n1231) );
AND2_X1 U890 ( .A1(KEYINPUT26), .A2(n1237), .ZN(n1236) );
NOR3_X1 U891 ( .A1(KEYINPUT26), .A2(n1238), .A3(n1239), .ZN(n1235) );
XNOR2_X1 U892 ( .A(KEYINPUT3), .B(n1047), .ZN(n1230) );
INV_X1 U893 ( .A(n1164), .ZN(n1047) );
NOR4_X1 U894 ( .A1(n1162), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1164) );
INV_X1 U895 ( .A(n1243), .ZN(n1241) );
AND2_X1 U896 ( .A1(n1191), .A2(n1244), .ZN(n1240) );
NAND2_X1 U897 ( .A1(n1082), .A2(n1040), .ZN(n1244) );
INV_X1 U898 ( .A(n1091), .ZN(n1040) );
INV_X1 U899 ( .A(n1092), .ZN(n1082) );
NOR3_X1 U900 ( .A1(n1245), .A2(n1193), .A3(n1083), .ZN(n1191) );
NAND4_X1 U901 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1162) );
INV_X1 U902 ( .A(n1046), .ZN(n1119) );
NAND3_X1 U903 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1046) );
NAND2_X1 U904 ( .A1(n1061), .A2(n1253), .ZN(n1252) );
XOR2_X1 U905 ( .A(KEYINPUT0), .B(n1254), .Z(n1253) );
NAND3_X1 U906 ( .A1(n1255), .A2(n1256), .A3(n1092), .ZN(n1250) );
NAND2_X1 U907 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U908 ( .A1(KEYINPUT25), .A2(n1259), .ZN(n1258) );
NAND3_X1 U909 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1255) );
NAND3_X1 U910 ( .A1(n1263), .A2(n1061), .A3(n1093), .ZN(n1261) );
OR2_X1 U911 ( .A1(n1264), .A2(KEYINPUT25), .ZN(n1260) );
XNOR2_X1 U912 ( .A(n1265), .B(n1266), .ZN(n1224) );
XNOR2_X1 U913 ( .A(KEYINPUT60), .B(KEYINPUT29), .ZN(n1265) );
NOR2_X1 U914 ( .A1(n1049), .A2(G952), .ZN(n1165) );
XOR2_X1 U915 ( .A(n1232), .B(n1267), .Z(G48) );
XNOR2_X1 U916 ( .A(G146), .B(KEYINPUT7), .ZN(n1267) );
NAND3_X1 U917 ( .A1(n1268), .A2(n1061), .A3(n1092), .ZN(n1232) );
NAND2_X1 U918 ( .A1(n1269), .A2(n1270), .ZN(G45) );
NAND3_X1 U919 ( .A1(G143), .A2(n1271), .A3(n1272), .ZN(n1270) );
NAND2_X1 U920 ( .A1(n1273), .A2(n1237), .ZN(n1269) );
INV_X1 U921 ( .A(n1272), .ZN(n1237) );
NAND2_X1 U922 ( .A1(n1238), .A2(n1061), .ZN(n1272) );
AND4_X1 U923 ( .A1(n1274), .A2(n1262), .A3(n1275), .A4(n1276), .ZN(n1238) );
NOR2_X1 U924 ( .A1(n1245), .A2(n1079), .ZN(n1276) );
NAND2_X1 U925 ( .A1(n1277), .A2(n1278), .ZN(n1273) );
NAND2_X1 U926 ( .A1(KEYINPUT30), .A2(G143), .ZN(n1278) );
NAND2_X1 U927 ( .A1(n1279), .A2(n1280), .ZN(n1277) );
INV_X1 U928 ( .A(KEYINPUT30), .ZN(n1280) );
NAND2_X1 U929 ( .A1(G143), .A2(n1271), .ZN(n1279) );
INV_X1 U930 ( .A(KEYINPUT50), .ZN(n1271) );
XNOR2_X1 U931 ( .A(G140), .B(n1233), .ZN(G42) );
OR4_X1 U932 ( .A1(n1088), .A2(n1281), .A3(n1065), .A4(n1245), .ZN(n1233) );
NAND2_X1 U933 ( .A1(n1282), .A2(n1283), .ZN(G39) );
NAND2_X1 U934 ( .A1(n1284), .A2(n1234), .ZN(n1283) );
NAND2_X1 U935 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
OR2_X1 U936 ( .A1(KEYINPUT24), .A2(KEYINPUT28), .ZN(n1286) );
NAND3_X1 U937 ( .A1(n1287), .A2(n1288), .A3(KEYINPUT28), .ZN(n1282) );
OR2_X1 U938 ( .A1(n1285), .A2(KEYINPUT24), .ZN(n1288) );
NAND2_X1 U939 ( .A1(n1289), .A2(n1285), .ZN(n1287) );
OR2_X1 U940 ( .A1(n1234), .A2(KEYINPUT24), .ZN(n1289) );
NAND3_X1 U941 ( .A1(n1268), .A2(n1076), .A3(n1290), .ZN(n1234) );
XNOR2_X1 U942 ( .A(G134), .B(n1251), .ZN(G36) );
NAND3_X1 U943 ( .A1(n1091), .A2(n1262), .A3(n1259), .ZN(n1251) );
XNOR2_X1 U944 ( .A(n1133), .B(n1291), .ZN(G33) );
NOR2_X1 U945 ( .A1(n1281), .A2(n1264), .ZN(n1291) );
INV_X1 U946 ( .A(n1259), .ZN(n1264) );
NOR3_X1 U947 ( .A1(n1065), .A2(n1245), .A3(n1079), .ZN(n1259) );
INV_X1 U948 ( .A(n1290), .ZN(n1065) );
NOR2_X1 U949 ( .A1(n1099), .A2(n1062), .ZN(n1290) );
INV_X1 U950 ( .A(n1292), .ZN(n1062) );
XNOR2_X1 U951 ( .A(G128), .B(n1293), .ZN(G30) );
NAND2_X1 U952 ( .A1(n1254), .A2(n1061), .ZN(n1293) );
AND2_X1 U953 ( .A1(n1268), .A2(n1091), .ZN(n1254) );
NOR4_X1 U954 ( .A1(n1245), .A2(n1294), .A3(n1295), .A4(n1257), .ZN(n1268) );
INV_X1 U955 ( .A(n1262), .ZN(n1257) );
XNOR2_X1 U956 ( .A(G101), .B(n1243), .ZN(G3) );
NAND3_X1 U957 ( .A1(n1076), .A2(n1067), .A3(n1296), .ZN(n1243) );
INV_X1 U958 ( .A(n1245), .ZN(n1067) );
XNOR2_X1 U959 ( .A(G125), .B(n1297), .ZN(G27) );
NAND4_X1 U960 ( .A1(KEYINPUT48), .A2(n1093), .A3(n1298), .A4(n1263), .ZN(n1297) );
INV_X1 U961 ( .A(n1088), .ZN(n1263) );
NOR2_X1 U962 ( .A1(n1239), .A2(n1281), .ZN(n1298) );
NAND2_X1 U963 ( .A1(n1092), .A2(n1262), .ZN(n1281) );
NAND2_X1 U964 ( .A1(n1084), .A2(n1299), .ZN(n1262) );
NAND2_X1 U965 ( .A1(n1126), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U966 ( .A(G900), .B(KEYINPUT23), .ZN(n1126) );
INV_X1 U967 ( .A(n1061), .ZN(n1239) );
XNOR2_X1 U968 ( .A(G122), .B(n1246), .ZN(G24) );
NAND3_X1 U969 ( .A1(n1093), .A2(n1077), .A3(n1301), .ZN(n1246) );
NOR3_X1 U970 ( .A1(n1193), .A2(n1302), .A3(n1303), .ZN(n1301) );
INV_X1 U971 ( .A(n1083), .ZN(n1077) );
NAND2_X1 U972 ( .A1(n1295), .A2(n1294), .ZN(n1083) );
XOR2_X1 U973 ( .A(n1247), .B(n1304), .Z(G21) );
NOR2_X1 U974 ( .A1(G119), .A2(KEYINPUT39), .ZN(n1304) );
NAND3_X1 U975 ( .A1(n1093), .A2(n1076), .A3(n1305), .ZN(n1247) );
NOR3_X1 U976 ( .A1(n1193), .A2(n1295), .A3(n1294), .ZN(n1305) );
XNOR2_X1 U977 ( .A(G116), .B(n1248), .ZN(G18) );
NAND3_X1 U978 ( .A1(n1296), .A2(n1091), .A3(n1093), .ZN(n1248) );
NOR2_X1 U979 ( .A1(n1275), .A2(n1302), .ZN(n1091) );
INV_X1 U980 ( .A(n1274), .ZN(n1302) );
XNOR2_X1 U981 ( .A(G113), .B(n1249), .ZN(G15) );
NAND3_X1 U982 ( .A1(n1296), .A2(n1092), .A3(n1093), .ZN(n1249) );
NOR2_X1 U983 ( .A1(n1069), .A2(n1098), .ZN(n1093) );
INV_X1 U984 ( .A(n1068), .ZN(n1098) );
NOR2_X1 U985 ( .A1(n1274), .A2(n1303), .ZN(n1092) );
NOR2_X1 U986 ( .A1(n1079), .A2(n1193), .ZN(n1296) );
OR2_X1 U987 ( .A1(n1306), .A2(n1295), .ZN(n1079) );
XOR2_X1 U988 ( .A(G110), .B(n1242), .Z(G12) );
NOR4_X1 U989 ( .A1(n1088), .A2(n1081), .A3(n1245), .A4(n1193), .ZN(n1242) );
NAND2_X1 U990 ( .A1(n1061), .A2(n1307), .ZN(n1193) );
NAND2_X1 U991 ( .A1(n1308), .A2(n1084), .ZN(n1307) );
NAND3_X1 U992 ( .A1(n1309), .A2(n1049), .A3(G952), .ZN(n1084) );
NAND2_X1 U993 ( .A1(n1300), .A2(n1310), .ZN(n1308) );
INV_X1 U994 ( .A(G898), .ZN(n1310) );
AND3_X1 U995 ( .A1(G902), .A2(n1309), .A3(G953), .ZN(n1300) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1309) );
NOR2_X1 U997 ( .A1(n1292), .A2(n1099), .ZN(n1061) );
INV_X1 U998 ( .A(n1063), .ZN(n1099) );
NAND2_X1 U999 ( .A1(G214), .A2(n1311), .ZN(n1063) );
NAND2_X1 U1000 ( .A1(n1312), .A2(n1313), .ZN(n1292) );
NAND2_X1 U1001 ( .A1(n1314), .A2(n1229), .ZN(n1313) );
NAND2_X1 U1002 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
NAND2_X1 U1003 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U1004 ( .A1(n1108), .A2(n1319), .ZN(n1312) );
NAND2_X1 U1005 ( .A1(n1318), .A2(n1320), .ZN(n1319) );
NAND2_X1 U1006 ( .A1(n1109), .A2(n1315), .ZN(n1320) );
INV_X1 U1007 ( .A(KEYINPUT11), .ZN(n1315) );
INV_X1 U1008 ( .A(n1229), .ZN(n1109) );
NAND2_X1 U1009 ( .A1(G210), .A2(n1311), .ZN(n1229) );
NAND2_X1 U1010 ( .A1(n1321), .A2(n1322), .ZN(n1311) );
INV_X1 U1011 ( .A(G237), .ZN(n1321) );
INV_X1 U1012 ( .A(KEYINPUT20), .ZN(n1318) );
INV_X1 U1013 ( .A(n1317), .ZN(n1108) );
NAND2_X1 U1014 ( .A1(n1323), .A2(n1322), .ZN(n1317) );
XNOR2_X1 U1015 ( .A(n1324), .B(n1325), .ZN(n1323) );
INV_X1 U1016 ( .A(n1227), .ZN(n1325) );
XNOR2_X1 U1017 ( .A(n1326), .B(n1327), .ZN(n1227) );
NOR2_X1 U1018 ( .A1(G953), .A2(n1141), .ZN(n1327) );
INV_X1 U1019 ( .A(G224), .ZN(n1141) );
NAND2_X1 U1020 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
OR2_X1 U1021 ( .A1(n1155), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1022 ( .A(n1331), .B(KEYINPUT46), .Z(n1328) );
NAND2_X1 U1023 ( .A1(n1330), .A2(n1155), .ZN(n1331) );
XOR2_X1 U1024 ( .A(G110), .B(G122), .Z(n1155) );
XOR2_X1 U1025 ( .A(n1153), .B(KEYINPUT21), .Z(n1330) );
XNOR2_X1 U1026 ( .A(n1332), .B(n1333), .ZN(n1153) );
XOR2_X1 U1027 ( .A(KEYINPUT49), .B(n1334), .Z(n1333) );
XNOR2_X1 U1028 ( .A(n1335), .B(n1336), .ZN(n1332) );
INV_X1 U1029 ( .A(n1337), .ZN(n1336) );
NAND2_X1 U1030 ( .A1(n1338), .A2(KEYINPUT35), .ZN(n1324) );
XNOR2_X1 U1031 ( .A(n1339), .B(n1266), .ZN(n1338) );
NAND2_X1 U1032 ( .A1(KEYINPUT63), .A2(n1207), .ZN(n1339) );
NAND2_X1 U1033 ( .A1(n1069), .A2(n1068), .ZN(n1245) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1340), .ZN(n1068) );
NAND2_X1 U1035 ( .A1(n1341), .A2(n1342), .ZN(n1069) );
OR2_X1 U1036 ( .A1(n1110), .A2(G469), .ZN(n1342) );
XOR2_X1 U1037 ( .A(n1343), .B(KEYINPUT41), .Z(n1341) );
NAND2_X1 U1038 ( .A1(G469), .A2(n1110), .ZN(n1343) );
NAND2_X1 U1039 ( .A1(n1344), .A2(n1322), .ZN(n1110) );
XOR2_X1 U1040 ( .A(n1345), .B(n1346), .Z(n1344) );
XNOR2_X1 U1041 ( .A(n1221), .B(n1129), .ZN(n1346) );
XOR2_X1 U1042 ( .A(n1134), .B(n1334), .Z(n1221) );
XNOR2_X1 U1043 ( .A(n1347), .B(n1348), .ZN(n1334) );
XOR2_X1 U1044 ( .A(KEYINPUT40), .B(G107), .Z(n1348) );
XNOR2_X1 U1045 ( .A(G104), .B(G101), .ZN(n1347) );
XOR2_X1 U1046 ( .A(n1349), .B(KEYINPUT34), .Z(n1134) );
XNOR2_X1 U1047 ( .A(n1202), .B(n1350), .ZN(n1345) );
XNOR2_X1 U1048 ( .A(n1351), .B(n1352), .ZN(n1350) );
INV_X1 U1049 ( .A(n1219), .ZN(n1352) );
XNOR2_X1 U1050 ( .A(n1353), .B(KEYINPUT42), .ZN(n1219) );
NAND2_X1 U1051 ( .A1(G227), .A2(n1049), .ZN(n1353) );
NOR2_X1 U1052 ( .A1(KEYINPUT43), .A2(n1354), .ZN(n1351) );
XNOR2_X1 U1053 ( .A(G110), .B(KEYINPUT5), .ZN(n1354) );
INV_X1 U1054 ( .A(n1076), .ZN(n1081) );
NOR2_X1 U1055 ( .A1(n1274), .A2(n1275), .ZN(n1076) );
INV_X1 U1056 ( .A(n1303), .ZN(n1275) );
XOR2_X1 U1057 ( .A(n1355), .B(G475), .Z(n1303) );
OR2_X1 U1058 ( .A1(n1184), .A2(G902), .ZN(n1355) );
XNOR2_X1 U1059 ( .A(n1356), .B(n1357), .ZN(n1184) );
XNOR2_X1 U1060 ( .A(n1188), .B(n1358), .ZN(n1357) );
NOR2_X1 U1061 ( .A1(KEYINPUT47), .A2(n1335), .ZN(n1358) );
INV_X1 U1062 ( .A(G104), .ZN(n1188) );
XOR2_X1 U1063 ( .A(n1359), .B(n1360), .Z(n1356) );
NOR2_X1 U1064 ( .A1(KEYINPUT58), .A2(n1266), .ZN(n1360) );
XOR2_X1 U1065 ( .A(n1361), .B(n1362), .Z(n1359) );
XNOR2_X1 U1066 ( .A(n1133), .B(n1363), .ZN(n1362) );
XNOR2_X1 U1067 ( .A(n1364), .B(G143), .ZN(n1363) );
INV_X1 U1068 ( .A(G131), .ZN(n1133) );
XNOR2_X1 U1069 ( .A(n1365), .B(n1129), .ZN(n1361) );
INV_X1 U1070 ( .A(n1366), .ZN(n1129) );
XOR2_X1 U1071 ( .A(n1367), .B(G122), .Z(n1365) );
NAND2_X1 U1072 ( .A1(G214), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1073 ( .A(n1369), .B(n1179), .Z(n1274) );
INV_X1 U1074 ( .A(G478), .ZN(n1179) );
NAND2_X1 U1075 ( .A1(n1176), .A2(n1322), .ZN(n1369) );
XNOR2_X1 U1076 ( .A(n1370), .B(n1371), .ZN(n1176) );
XOR2_X1 U1077 ( .A(G107), .B(n1372), .Z(n1371) );
XOR2_X1 U1078 ( .A(G122), .B(G116), .Z(n1372) );
XNOR2_X1 U1079 ( .A(n1373), .B(n1135), .ZN(n1370) );
XOR2_X1 U1080 ( .A(n1374), .B(n1375), .Z(n1373) );
NAND2_X1 U1081 ( .A1(G217), .A2(n1376), .ZN(n1374) );
NAND2_X1 U1082 ( .A1(n1295), .A2(n1306), .ZN(n1088) );
INV_X1 U1083 ( .A(n1294), .ZN(n1306) );
XOR2_X1 U1084 ( .A(n1105), .B(n1170), .Z(n1294) );
NAND2_X1 U1085 ( .A1(G217), .A2(n1340), .ZN(n1170) );
NAND2_X1 U1086 ( .A1(G234), .A2(n1322), .ZN(n1340) );
NOR2_X1 U1087 ( .A1(n1173), .A2(G902), .ZN(n1105) );
INV_X1 U1088 ( .A(n1169), .ZN(n1173) );
XNOR2_X1 U1089 ( .A(n1377), .B(n1378), .ZN(n1169) );
XOR2_X1 U1090 ( .A(n1379), .B(n1380), .Z(n1378) );
XNOR2_X1 U1091 ( .A(G128), .B(n1266), .ZN(n1380) );
INV_X1 U1092 ( .A(G125), .ZN(n1266) );
XNOR2_X1 U1093 ( .A(n1364), .B(G137), .ZN(n1379) );
INV_X1 U1094 ( .A(G146), .ZN(n1364) );
XOR2_X1 U1095 ( .A(n1381), .B(n1220), .Z(n1377) );
XOR2_X1 U1096 ( .A(G110), .B(n1366), .Z(n1220) );
XOR2_X1 U1097 ( .A(G140), .B(KEYINPUT1), .Z(n1366) );
XOR2_X1 U1098 ( .A(n1382), .B(G119), .Z(n1381) );
NAND2_X1 U1099 ( .A1(G221), .A2(n1376), .ZN(n1382) );
AND2_X1 U1100 ( .A1(G234), .A2(n1049), .ZN(n1376) );
INV_X1 U1101 ( .A(G953), .ZN(n1049) );
XNOR2_X1 U1102 ( .A(n1104), .B(n1103), .ZN(n1295) );
INV_X1 U1103 ( .A(G472), .ZN(n1103) );
NAND2_X1 U1104 ( .A1(n1383), .A2(n1322), .ZN(n1104) );
INV_X1 U1105 ( .A(G902), .ZN(n1322) );
XOR2_X1 U1106 ( .A(n1384), .B(n1385), .Z(n1383) );
XOR2_X1 U1107 ( .A(n1386), .B(n1207), .Z(n1385) );
XOR2_X1 U1108 ( .A(n1349), .B(KEYINPUT6), .Z(n1207) );
XNOR2_X1 U1109 ( .A(G146), .B(n1375), .ZN(n1349) );
XOR2_X1 U1110 ( .A(G128), .B(G143), .Z(n1375) );
NAND2_X1 U1111 ( .A1(n1387), .A2(n1388), .ZN(n1386) );
OR2_X1 U1112 ( .A1(n1197), .A2(n1195), .ZN(n1388) );
XOR2_X1 U1113 ( .A(n1389), .B(KEYINPUT27), .Z(n1387) );
NAND2_X1 U1114 ( .A1(n1197), .A2(n1195), .ZN(n1389) );
NAND2_X1 U1115 ( .A1(G210), .A2(n1368), .ZN(n1195) );
NOR2_X1 U1116 ( .A1(G953), .A2(G237), .ZN(n1368) );
INV_X1 U1117 ( .A(G101), .ZN(n1197) );
XOR2_X1 U1118 ( .A(n1390), .B(n1391), .Z(n1384) );
XNOR2_X1 U1119 ( .A(KEYINPUT54), .B(n1392), .ZN(n1391) );
NOR2_X1 U1120 ( .A1(KEYINPUT52), .A2(n1202), .ZN(n1392) );
XNOR2_X1 U1121 ( .A(n1393), .B(n1394), .ZN(n1202) );
XNOR2_X1 U1122 ( .A(n1285), .B(G131), .ZN(n1394) );
INV_X1 U1123 ( .A(G137), .ZN(n1285) );
NAND2_X1 U1124 ( .A1(KEYINPUT36), .A2(n1135), .ZN(n1393) );
XNOR2_X1 U1125 ( .A(G134), .B(KEYINPUT62), .ZN(n1135) );
NAND2_X1 U1126 ( .A1(KEYINPUT19), .A2(n1203), .ZN(n1390) );
XNOR2_X1 U1127 ( .A(n1337), .B(n1395), .ZN(n1203) );
NOR2_X1 U1128 ( .A1(KEYINPUT9), .A2(n1335), .ZN(n1395) );
XNOR2_X1 U1129 ( .A(G113), .B(KEYINPUT16), .ZN(n1335) );
XOR2_X1 U1130 ( .A(G116), .B(G119), .Z(n1337) );
endmodule


