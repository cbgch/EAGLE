//Key = 0101101100101100011001011101011010100100001010110000000000100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;

XOR2_X1 U724 ( .A(G107), .B(n1015), .Z(G9) );
NOR2_X1 U725 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U726 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NAND3_X1 U727 ( .A1(n1022), .A2(n1023), .A3(n1024), .ZN(n1018) );
NAND2_X1 U728 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U729 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U730 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NAND3_X1 U731 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1030) );
NAND2_X1 U732 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND2_X1 U733 ( .A1(n1037), .A2(n1038), .ZN(n1032) );
NAND2_X1 U734 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U735 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
INV_X1 U736 ( .A(n1043), .ZN(n1039) );
NAND3_X1 U737 ( .A1(n1035), .A2(n1044), .A3(n1037), .ZN(n1027) );
NAND2_X1 U738 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U739 ( .A1(n1031), .A2(n1047), .ZN(n1046) );
OR2_X1 U740 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U741 ( .A1(n1029), .A2(n1050), .ZN(n1045) );
NAND2_X1 U742 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U743 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
INV_X1 U744 ( .A(n1055), .ZN(n1025) );
NOR3_X1 U745 ( .A1(n1056), .A2(G953), .A3(G952), .ZN(n1016) );
INV_X1 U746 ( .A(n1022), .ZN(n1056) );
NAND4_X1 U747 ( .A1(n1057), .A2(n1058), .A3(n1042), .A4(n1059), .ZN(n1022) );
NOR3_X1 U748 ( .A1(n1041), .A2(n1060), .A3(n1061), .ZN(n1059) );
XOR2_X1 U749 ( .A(KEYINPUT9), .B(n1062), .Z(n1057) );
NOR3_X1 U750 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NOR2_X1 U751 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U752 ( .A(n1068), .ZN(n1064) );
NAND3_X1 U753 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1063) );
INV_X1 U754 ( .A(n1072), .ZN(n1071) );
NAND2_X1 U755 ( .A1(KEYINPUT1), .A2(n1073), .ZN(n1070) );
OR2_X1 U756 ( .A1(n1049), .A2(KEYINPUT1), .ZN(n1069) );
XOR2_X1 U757 ( .A(n1074), .B(n1075), .Z(G72) );
NOR2_X1 U758 ( .A1(n1076), .A2(n1023), .ZN(n1075) );
AND2_X1 U759 ( .A1(G227), .A2(G900), .ZN(n1076) );
NAND2_X1 U760 ( .A1(n1077), .A2(n1078), .ZN(n1074) );
NAND3_X1 U761 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NAND2_X1 U762 ( .A1(G953), .A2(n1082), .ZN(n1080) );
XOR2_X1 U763 ( .A(KEYINPUT18), .B(n1083), .Z(n1079) );
NAND2_X1 U764 ( .A1(n1083), .A2(n1084), .ZN(n1077) );
INV_X1 U765 ( .A(n1081), .ZN(n1084) );
XNOR2_X1 U766 ( .A(n1085), .B(n1086), .ZN(n1081) );
AND2_X1 U767 ( .A1(n1087), .A2(n1023), .ZN(n1083) );
NAND2_X1 U768 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U769 ( .A(n1019), .B(KEYINPUT10), .Z(n1088) );
XOR2_X1 U770 ( .A(n1090), .B(n1091), .Z(G69) );
XOR2_X1 U771 ( .A(n1092), .B(n1093), .Z(n1091) );
NOR3_X1 U772 ( .A1(n1094), .A2(KEYINPUT19), .A3(G953), .ZN(n1093) );
INV_X1 U773 ( .A(n1021), .ZN(n1094) );
NOR2_X1 U774 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
XOR2_X1 U775 ( .A(KEYINPUT16), .B(n1097), .Z(n1096) );
NOR2_X1 U776 ( .A1(G898), .A2(n1023), .ZN(n1097) );
XOR2_X1 U777 ( .A(n1098), .B(KEYINPUT30), .Z(n1095) );
NOR2_X1 U778 ( .A1(n1099), .A2(n1023), .ZN(n1090) );
AND2_X1 U779 ( .A1(G224), .A2(G898), .ZN(n1099) );
NOR2_X1 U780 ( .A1(n1100), .A2(n1101), .ZN(G66) );
XOR2_X1 U781 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND3_X1 U782 ( .A1(n1104), .A2(G217), .A3(KEYINPUT7), .ZN(n1102) );
NOR2_X1 U783 ( .A1(n1100), .A2(n1105), .ZN(G63) );
XOR2_X1 U784 ( .A(n1106), .B(n1107), .Z(n1105) );
NOR2_X1 U785 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U786 ( .A(KEYINPUT13), .B(G478), .Z(n1109) );
NOR2_X1 U787 ( .A1(n1100), .A2(n1110), .ZN(G60) );
XNOR2_X1 U788 ( .A(n1111), .B(n1112), .ZN(n1110) );
AND2_X1 U789 ( .A1(G475), .A2(n1104), .ZN(n1112) );
XOR2_X1 U790 ( .A(G104), .B(n1113), .Z(G6) );
NOR2_X1 U791 ( .A1(n1100), .A2(n1114), .ZN(G57) );
XOR2_X1 U792 ( .A(n1115), .B(n1116), .Z(n1114) );
XOR2_X1 U793 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U794 ( .A(n1119), .B(n1120), .ZN(n1118) );
XOR2_X1 U795 ( .A(n1121), .B(n1122), .Z(n1115) );
AND2_X1 U796 ( .A1(G472), .A2(n1104), .ZN(n1122) );
XOR2_X1 U797 ( .A(n1123), .B(n1124), .Z(n1121) );
NOR3_X1 U798 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(G54) );
NOR3_X1 U799 ( .A1(n1128), .A2(G953), .A3(G952), .ZN(n1127) );
AND2_X1 U800 ( .A1(n1128), .A2(n1100), .ZN(n1126) );
INV_X1 U801 ( .A(KEYINPUT49), .ZN(n1128) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1125) );
XNOR2_X1 U803 ( .A(n1131), .B(n1132), .ZN(n1129) );
NAND2_X1 U804 ( .A1(KEYINPUT58), .A2(n1133), .ZN(n1132) );
NAND2_X1 U805 ( .A1(n1104), .A2(G469), .ZN(n1133) );
INV_X1 U806 ( .A(n1108), .ZN(n1104) );
NAND2_X1 U807 ( .A1(KEYINPUT17), .A2(n1134), .ZN(n1131) );
XOR2_X1 U808 ( .A(KEYINPUT12), .B(n1135), .Z(n1134) );
NOR3_X1 U809 ( .A1(n1100), .A2(n1136), .A3(n1137), .ZN(G51) );
NOR2_X1 U810 ( .A1(n1138), .A2(n1098), .ZN(n1137) );
XOR2_X1 U811 ( .A(KEYINPUT22), .B(n1139), .Z(n1138) );
NOR2_X1 U812 ( .A1(n1140), .A2(n1141), .ZN(n1136) );
XNOR2_X1 U813 ( .A(n1139), .B(KEYINPUT62), .ZN(n1141) );
XNOR2_X1 U814 ( .A(n1142), .B(n1143), .ZN(n1139) );
XOR2_X1 U815 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U816 ( .A(KEYINPUT41), .B(KEYINPUT20), .ZN(n1145) );
XNOR2_X1 U817 ( .A(n1146), .B(n1147), .ZN(n1142) );
NOR2_X1 U818 ( .A1(n1108), .A2(n1148), .ZN(n1147) );
XOR2_X1 U819 ( .A(KEYINPUT27), .B(G210), .Z(n1148) );
NAND2_X1 U820 ( .A1(G902), .A2(n1149), .ZN(n1108) );
OR3_X1 U821 ( .A1(n1021), .A2(n1020), .A3(n1019), .ZN(n1149) );
NAND4_X1 U822 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1019) );
NAND4_X1 U823 ( .A1(n1048), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1150) );
XNOR2_X1 U824 ( .A(n1089), .B(KEYINPUT40), .ZN(n1020) );
AND4_X1 U825 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1089) );
NAND4_X1 U826 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1021) );
NOR4_X1 U827 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1015), .ZN(n1164) );
AND3_X1 U828 ( .A1(n1029), .A2(n1168), .A3(n1036), .ZN(n1015) );
NOR2_X1 U829 ( .A1(n1113), .A2(n1169), .ZN(n1163) );
NOR3_X1 U830 ( .A1(n1073), .A2(n1170), .A3(n1171), .ZN(n1113) );
INV_X1 U831 ( .A(n1029), .ZN(n1073) );
NAND4_X1 U832 ( .A1(n1049), .A2(n1036), .A3(n1172), .A4(n1173), .ZN(n1162) );
OR2_X1 U833 ( .A1(n1174), .A2(KEYINPUT50), .ZN(n1173) );
NAND2_X1 U834 ( .A1(KEYINPUT50), .A2(n1175), .ZN(n1172) );
NAND2_X1 U835 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NAND3_X1 U836 ( .A1(n1048), .A2(n1168), .A3(n1037), .ZN(n1161) );
NOR2_X1 U837 ( .A1(n1023), .A2(G952), .ZN(n1100) );
XOR2_X1 U838 ( .A(n1178), .B(n1157), .Z(G48) );
NAND3_X1 U839 ( .A1(n1179), .A2(n1155), .A3(n1180), .ZN(n1157) );
XNOR2_X1 U840 ( .A(G143), .B(n1158), .ZN(G45) );
NAND4_X1 U841 ( .A1(n1181), .A2(n1182), .A3(n1072), .A4(n1155), .ZN(n1158) );
XOR2_X1 U842 ( .A(n1183), .B(KEYINPUT5), .Z(n1181) );
XNOR2_X1 U843 ( .A(G140), .B(n1159), .ZN(G42) );
NAND4_X1 U844 ( .A1(n1043), .A2(n1156), .A3(n1031), .A4(n1184), .ZN(n1159) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1185), .ZN(n1184) );
XNOR2_X1 U846 ( .A(G137), .B(n1160), .ZN(G39) );
NAND3_X1 U847 ( .A1(n1031), .A2(n1179), .A3(n1037), .ZN(n1160) );
XNOR2_X1 U848 ( .A(G134), .B(n1151), .ZN(G36) );
NAND3_X1 U849 ( .A1(n1182), .A2(n1036), .A3(n1031), .ZN(n1151) );
XNOR2_X1 U850 ( .A(G131), .B(n1152), .ZN(G33) );
NAND3_X1 U851 ( .A1(n1031), .A2(n1182), .A3(n1180), .ZN(n1152) );
AND3_X1 U852 ( .A1(n1043), .A2(n1156), .A3(n1049), .ZN(n1182) );
AND2_X1 U853 ( .A1(n1054), .A2(n1058), .ZN(n1031) );
XNOR2_X1 U854 ( .A(G128), .B(n1153), .ZN(G30) );
NAND3_X1 U855 ( .A1(n1036), .A2(n1155), .A3(n1179), .ZN(n1153) );
AND4_X1 U856 ( .A1(n1043), .A2(n1186), .A3(n1156), .A4(n1187), .ZN(n1179) );
XOR2_X1 U857 ( .A(G101), .B(n1167), .Z(G3) );
AND3_X1 U858 ( .A1(n1049), .A2(n1168), .A3(n1037), .ZN(n1167) );
INV_X1 U859 ( .A(n1170), .ZN(n1168) );
XOR2_X1 U860 ( .A(G125), .B(n1188), .Z(G27) );
NOR2_X1 U861 ( .A1(n1189), .A2(n1051), .ZN(n1188) );
INV_X1 U862 ( .A(n1155), .ZN(n1051) );
XOR2_X1 U863 ( .A(n1190), .B(KEYINPUT56), .Z(n1189) );
NAND3_X1 U864 ( .A1(n1191), .A2(n1156), .A3(n1154), .ZN(n1190) );
INV_X1 U865 ( .A(n1033), .ZN(n1154) );
NAND2_X1 U866 ( .A1(n1035), .A2(n1180), .ZN(n1033) );
NAND2_X1 U867 ( .A1(n1055), .A2(n1192), .ZN(n1156) );
NAND4_X1 U868 ( .A1(G953), .A2(n1193), .A3(n1194), .A4(n1082), .ZN(n1192) );
INV_X1 U869 ( .A(G900), .ZN(n1082) );
XOR2_X1 U870 ( .A(KEYINPUT26), .B(G902), .Z(n1193) );
XOR2_X1 U871 ( .A(KEYINPUT45), .B(n1048), .Z(n1191) );
INV_X1 U872 ( .A(n1185), .ZN(n1048) );
XOR2_X1 U873 ( .A(G122), .B(n1169), .Z(G24) );
AND4_X1 U874 ( .A1(n1174), .A2(n1029), .A3(n1195), .A4(n1196), .ZN(n1169) );
NAND2_X1 U875 ( .A1(KEYINPUT5), .A2(n1171), .ZN(n1196) );
NAND2_X1 U876 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
INV_X1 U877 ( .A(KEYINPUT5), .ZN(n1198) );
NAND2_X1 U878 ( .A1(n1072), .A2(n1183), .ZN(n1197) );
NOR2_X1 U879 ( .A1(n1187), .A2(n1186), .ZN(n1029) );
XOR2_X1 U880 ( .A(n1166), .B(n1199), .Z(G21) );
NOR2_X1 U881 ( .A1(KEYINPUT59), .A2(n1200), .ZN(n1199) );
AND4_X1 U882 ( .A1(n1037), .A2(n1174), .A3(n1186), .A4(n1187), .ZN(n1166) );
INV_X1 U883 ( .A(n1201), .ZN(n1186) );
NAND2_X1 U884 ( .A1(n1202), .A2(n1203), .ZN(G18) );
NAND2_X1 U885 ( .A1(G116), .A2(n1204), .ZN(n1203) );
XOR2_X1 U886 ( .A(KEYINPUT21), .B(n1205), .Z(n1202) );
NOR2_X1 U887 ( .A1(G116), .A2(n1204), .ZN(n1205) );
NAND3_X1 U888 ( .A1(n1049), .A2(n1036), .A3(n1174), .ZN(n1204) );
NOR2_X1 U889 ( .A1(n1072), .A2(n1206), .ZN(n1036) );
XOR2_X1 U890 ( .A(G113), .B(n1165), .Z(G15) );
AND3_X1 U891 ( .A1(n1180), .A2(n1049), .A3(n1174), .ZN(n1165) );
AND2_X1 U892 ( .A1(n1035), .A2(n1176), .ZN(n1174) );
INV_X1 U893 ( .A(n1177), .ZN(n1035) );
NAND2_X1 U894 ( .A1(n1207), .A2(n1042), .ZN(n1177) );
XNOR2_X1 U895 ( .A(n1041), .B(KEYINPUT28), .ZN(n1207) );
NOR2_X1 U896 ( .A1(n1187), .A2(n1201), .ZN(n1049) );
INV_X1 U897 ( .A(n1171), .ZN(n1180) );
NAND2_X1 U898 ( .A1(n1206), .A2(n1072), .ZN(n1171) );
INV_X1 U899 ( .A(n1183), .ZN(n1206) );
XOR2_X1 U900 ( .A(G110), .B(n1208), .Z(G12) );
NOR4_X1 U901 ( .A1(KEYINPUT60), .A2(n1209), .A3(n1170), .A4(n1185), .ZN(n1208) );
NAND2_X1 U902 ( .A1(n1201), .A2(n1187), .ZN(n1185) );
NAND3_X1 U903 ( .A1(n1210), .A2(n1211), .A3(n1212), .ZN(n1187) );
OR2_X1 U904 ( .A1(n1213), .A2(n1103), .ZN(n1212) );
NAND3_X1 U905 ( .A1(n1103), .A2(n1213), .A3(n1214), .ZN(n1211) );
NAND2_X1 U906 ( .A1(G217), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U907 ( .A(n1216), .B(n1217), .ZN(n1103) );
XOR2_X1 U908 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U909 ( .A(G137), .B(G110), .Z(n1219) );
XOR2_X1 U910 ( .A(KEYINPUT14), .B(G146), .Z(n1218) );
XOR2_X1 U911 ( .A(n1220), .B(n1221), .Z(n1216) );
XNOR2_X1 U912 ( .A(n1222), .B(n1223), .ZN(n1221) );
NOR2_X1 U913 ( .A1(KEYINPUT43), .A2(n1086), .ZN(n1223) );
XOR2_X1 U914 ( .A(G140), .B(n1144), .Z(n1086) );
NAND2_X1 U915 ( .A1(KEYINPUT24), .A2(n1224), .ZN(n1222) );
XOR2_X1 U916 ( .A(G128), .B(G119), .Z(n1224) );
NAND2_X1 U917 ( .A1(G221), .A2(n1225), .ZN(n1220) );
NAND2_X1 U918 ( .A1(G902), .A2(G217), .ZN(n1210) );
XOR2_X1 U919 ( .A(n1226), .B(G472), .Z(n1201) );
NAND2_X1 U920 ( .A1(n1214), .A2(n1227), .ZN(n1226) );
NAND2_X1 U921 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U922 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U923 ( .A(n1232), .B(KEYINPUT53), .Z(n1228) );
NAND2_X1 U924 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
XNOR2_X1 U925 ( .A(n1231), .B(KEYINPUT52), .ZN(n1234) );
AND2_X1 U926 ( .A1(n1235), .A2(n1236), .ZN(n1231) );
NAND2_X1 U927 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
XNOR2_X1 U928 ( .A(n1239), .B(n1119), .ZN(n1237) );
NAND2_X1 U929 ( .A1(n1240), .A2(n1117), .ZN(n1235) );
INV_X1 U930 ( .A(n1238), .ZN(n1117) );
XOR2_X1 U931 ( .A(n1241), .B(n1242), .Z(n1238) );
XOR2_X1 U932 ( .A(G113), .B(n1243), .Z(n1242) );
NOR2_X1 U933 ( .A1(G119), .A2(KEYINPUT15), .ZN(n1243) );
XNOR2_X1 U934 ( .A(G116), .B(KEYINPUT2), .ZN(n1241) );
XOR2_X1 U935 ( .A(n1239), .B(n1119), .Z(n1240) );
NAND2_X1 U936 ( .A1(KEYINPUT6), .A2(n1120), .ZN(n1239) );
XOR2_X1 U937 ( .A(n1230), .B(KEYINPUT37), .Z(n1233) );
XOR2_X1 U938 ( .A(n1244), .B(G101), .Z(n1230) );
NAND2_X1 U939 ( .A1(KEYINPUT3), .A2(n1123), .ZN(n1244) );
AND3_X1 U940 ( .A1(n1245), .A2(n1023), .A3(G210), .ZN(n1123) );
NAND2_X1 U941 ( .A1(n1043), .A2(n1176), .ZN(n1170) );
AND2_X1 U942 ( .A1(n1155), .A2(n1246), .ZN(n1176) );
NAND2_X1 U943 ( .A1(n1055), .A2(n1247), .ZN(n1246) );
NAND4_X1 U944 ( .A1(G953), .A2(G902), .A3(n1194), .A4(n1248), .ZN(n1247) );
INV_X1 U945 ( .A(G898), .ZN(n1248) );
NAND3_X1 U946 ( .A1(n1194), .A2(n1023), .A3(G952), .ZN(n1055) );
NAND2_X1 U947 ( .A1(G237), .A2(G234), .ZN(n1194) );
NOR2_X1 U948 ( .A1(n1053), .A2(n1054), .ZN(n1155) );
NOR2_X1 U949 ( .A1(n1249), .A2(n1061), .ZN(n1054) );
NOR2_X1 U950 ( .A1(n1250), .A2(n1251), .ZN(n1061) );
AND2_X1 U951 ( .A1(G210), .A2(n1252), .ZN(n1251) );
XOR2_X1 U952 ( .A(n1060), .B(KEYINPUT39), .Z(n1249) );
AND3_X1 U953 ( .A1(n1250), .A2(n1252), .A3(G210), .ZN(n1060) );
NAND2_X1 U954 ( .A1(n1253), .A2(n1214), .ZN(n1250) );
XOR2_X1 U955 ( .A(n1254), .B(n1255), .Z(n1253) );
XOR2_X1 U956 ( .A(n1140), .B(n1146), .Z(n1255) );
XOR2_X1 U957 ( .A(n1256), .B(n1119), .Z(n1146) );
XOR2_X1 U958 ( .A(n1257), .B(n1258), .Z(n1119) );
XOR2_X1 U959 ( .A(G146), .B(G128), .Z(n1258) );
NAND2_X1 U960 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
XNOR2_X1 U961 ( .A(KEYINPUT8), .B(KEYINPUT35), .ZN(n1259) );
NAND2_X1 U962 ( .A1(G224), .A2(n1023), .ZN(n1256) );
INV_X1 U963 ( .A(n1098), .ZN(n1140) );
XOR2_X1 U964 ( .A(n1261), .B(n1262), .Z(n1098) );
XNOR2_X1 U965 ( .A(n1263), .B(n1264), .ZN(n1262) );
NAND2_X1 U966 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
NAND2_X1 U967 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U968 ( .A1(KEYINPUT47), .A2(n1269), .ZN(n1268) );
NAND2_X1 U969 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
INV_X1 U970 ( .A(G113), .ZN(n1270) );
INV_X1 U971 ( .A(n1272), .ZN(n1267) );
NAND2_X1 U972 ( .A1(G113), .A2(n1273), .ZN(n1265) );
NAND2_X1 U973 ( .A1(n1271), .A2(n1274), .ZN(n1273) );
NAND2_X1 U974 ( .A1(n1272), .A2(KEYINPUT47), .ZN(n1274) );
XOR2_X1 U975 ( .A(n1200), .B(G116), .Z(n1272) );
INV_X1 U976 ( .A(G119), .ZN(n1200) );
INV_X1 U977 ( .A(KEYINPUT48), .ZN(n1271) );
XOR2_X1 U978 ( .A(n1275), .B(n1276), .Z(n1261) );
XOR2_X1 U979 ( .A(G110), .B(n1277), .Z(n1276) );
NOR2_X1 U980 ( .A1(KEYINPUT54), .A2(n1124), .ZN(n1277) );
INV_X1 U981 ( .A(G101), .ZN(n1124) );
NAND2_X1 U982 ( .A1(KEYINPUT25), .A2(n1278), .ZN(n1275) );
INV_X1 U983 ( .A(G107), .ZN(n1278) );
XNOR2_X1 U984 ( .A(KEYINPUT31), .B(n1279), .ZN(n1254) );
NOR2_X1 U985 ( .A1(KEYINPUT57), .A2(n1280), .ZN(n1279) );
XOR2_X1 U986 ( .A(n1144), .B(KEYINPUT11), .Z(n1280) );
INV_X1 U987 ( .A(n1058), .ZN(n1053) );
NAND2_X1 U988 ( .A1(G214), .A2(n1252), .ZN(n1058) );
NAND2_X1 U989 ( .A1(n1214), .A2(n1245), .ZN(n1252) );
NOR2_X1 U990 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
AND2_X1 U991 ( .A1(G221), .A2(n1281), .ZN(n1041) );
XOR2_X1 U992 ( .A(KEYINPUT44), .B(n1282), .Z(n1281) );
NOR2_X1 U993 ( .A1(G902), .A2(n1215), .ZN(n1282) );
XOR2_X1 U994 ( .A(n1283), .B(G469), .Z(n1042) );
NAND2_X1 U995 ( .A1(n1284), .A2(n1214), .ZN(n1283) );
XNOR2_X1 U996 ( .A(n1285), .B(n1135), .ZN(n1284) );
XNOR2_X1 U997 ( .A(n1286), .B(n1287), .ZN(n1135) );
XOR2_X1 U998 ( .A(G107), .B(G104), .Z(n1287) );
XOR2_X1 U999 ( .A(n1085), .B(G101), .Z(n1286) );
XOR2_X1 U1000 ( .A(n1288), .B(n1289), .Z(n1085) );
XNOR2_X1 U1001 ( .A(G128), .B(n1290), .ZN(n1289) );
NAND2_X1 U1002 ( .A1(KEYINPUT61), .A2(n1178), .ZN(n1290) );
INV_X1 U1003 ( .A(G146), .ZN(n1178) );
XNOR2_X1 U1004 ( .A(n1120), .B(n1260), .ZN(n1288) );
XOR2_X1 U1005 ( .A(G143), .B(KEYINPUT29), .Z(n1260) );
XOR2_X1 U1006 ( .A(G131), .B(n1291), .Z(n1120) );
XOR2_X1 U1007 ( .A(G137), .B(G134), .Z(n1291) );
NAND2_X1 U1008 ( .A1(n1292), .A2(n1293), .ZN(n1285) );
OR2_X1 U1009 ( .A1(n1130), .A2(KEYINPUT38), .ZN(n1293) );
XNOR2_X1 U1010 ( .A(n1294), .B(n1295), .ZN(n1130) );
NAND3_X1 U1011 ( .A1(n1295), .A2(n1294), .A3(KEYINPUT38), .ZN(n1292) );
NAND2_X1 U1012 ( .A1(G227), .A2(n1023), .ZN(n1294) );
XOR2_X1 U1013 ( .A(G110), .B(G140), .Z(n1295) );
XNOR2_X1 U1014 ( .A(n1037), .B(KEYINPUT63), .ZN(n1209) );
NOR2_X1 U1015 ( .A1(n1183), .A2(n1072), .ZN(n1037) );
XOR2_X1 U1016 ( .A(n1296), .B(n1297), .Z(n1072) );
XOR2_X1 U1017 ( .A(KEYINPUT32), .B(G475), .Z(n1297) );
NAND2_X1 U1018 ( .A1(n1111), .A2(n1214), .ZN(n1296) );
INV_X1 U1019 ( .A(G902), .ZN(n1214) );
XNOR2_X1 U1020 ( .A(n1298), .B(n1299), .ZN(n1111) );
XOR2_X1 U1021 ( .A(n1300), .B(n1301), .Z(n1299) );
XOR2_X1 U1022 ( .A(G140), .B(G113), .Z(n1301) );
XOR2_X1 U1023 ( .A(G146), .B(G143), .Z(n1300) );
XOR2_X1 U1024 ( .A(n1302), .B(n1303), .Z(n1298) );
XNOR2_X1 U1025 ( .A(n1304), .B(n1305), .ZN(n1303) );
NOR2_X1 U1026 ( .A1(KEYINPUT55), .A2(G131), .ZN(n1305) );
NAND4_X1 U1027 ( .A1(KEYINPUT46), .A2(G214), .A3(n1245), .A4(n1023), .ZN(n1304) );
INV_X1 U1028 ( .A(G953), .ZN(n1023) );
INV_X1 U1029 ( .A(G237), .ZN(n1245) );
NAND2_X1 U1030 ( .A1(n1306), .A2(n1307), .ZN(n1302) );
NAND2_X1 U1031 ( .A1(n1308), .A2(n1144), .ZN(n1307) );
INV_X1 U1032 ( .A(G125), .ZN(n1144) );
XOR2_X1 U1033 ( .A(KEYINPUT36), .B(n1264), .Z(n1308) );
NAND2_X1 U1034 ( .A1(n1309), .A2(G125), .ZN(n1306) );
XOR2_X1 U1035 ( .A(KEYINPUT42), .B(n1264), .Z(n1309) );
XOR2_X1 U1036 ( .A(G104), .B(G122), .Z(n1264) );
NAND3_X1 U1037 ( .A1(n1310), .A2(n1311), .A3(n1068), .ZN(n1183) );
NAND2_X1 U1038 ( .A1(n1066), .A2(n1067), .ZN(n1068) );
OR3_X1 U1039 ( .A1(n1067), .A2(n1066), .A3(KEYINPUT0), .ZN(n1311) );
NOR2_X1 U1040 ( .A1(n1106), .A2(G902), .ZN(n1066) );
XOR2_X1 U1041 ( .A(n1312), .B(n1313), .Z(n1106) );
XOR2_X1 U1042 ( .A(G107), .B(n1314), .Z(n1313) );
XOR2_X1 U1043 ( .A(KEYINPUT23), .B(G134), .Z(n1314) );
XOR2_X1 U1044 ( .A(n1315), .B(n1316), .Z(n1312) );
XOR2_X1 U1045 ( .A(n1317), .B(n1318), .Z(n1316) );
NAND2_X1 U1046 ( .A1(KEYINPUT4), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1047 ( .A(G143), .B(G128), .Z(n1319) );
NAND2_X1 U1048 ( .A1(n1320), .A2(n1321), .ZN(n1317) );
NAND2_X1 U1049 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1050 ( .A(KEYINPUT34), .B(n1324), .Z(n1320) );
NOR2_X1 U1051 ( .A1(n1323), .A2(n1322), .ZN(n1324) );
XOR2_X1 U1052 ( .A(KEYINPUT33), .B(G116), .Z(n1322) );
INV_X1 U1053 ( .A(G122), .ZN(n1323) );
NAND2_X1 U1054 ( .A1(G217), .A2(n1225), .ZN(n1315) );
NOR2_X1 U1055 ( .A1(n1215), .A2(G953), .ZN(n1225) );
INV_X1 U1056 ( .A(G234), .ZN(n1215) );
NAND2_X1 U1057 ( .A1(KEYINPUT0), .A2(n1067), .ZN(n1310) );
XNOR2_X1 U1058 ( .A(G478), .B(KEYINPUT51), .ZN(n1067) );
endmodule


