//Key = 1111010111001011000001011110101000001001110011111010111100001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
n1423, n1424, n1425, n1426, n1427;

XNOR2_X1 U790 ( .A(n1093), .B(n1094), .ZN(G9) );
NOR2_X1 U791 ( .A1(KEYINPUT13), .A2(n1095), .ZN(n1094) );
INV_X1 U792 ( .A(G107), .ZN(n1095) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(G75) );
NOR4_X1 U794 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XOR2_X1 U795 ( .A(n1102), .B(KEYINPUT4), .Z(n1100) );
NAND2_X1 U796 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND3_X1 U797 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
NAND3_X1 U798 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1106) );
NAND4_X1 U799 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1110) );
NAND4_X1 U800 ( .A1(KEYINPUT26), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1109) );
NAND3_X1 U801 ( .A1(n1113), .A2(n1118), .A3(n1119), .ZN(n1108) );
NAND2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1118) );
NAND2_X1 U803 ( .A1(n1114), .A2(n1122), .ZN(n1121) );
INV_X1 U804 ( .A(KEYINPUT26), .ZN(n1122) );
NAND2_X1 U805 ( .A1(n1123), .A2(n1124), .ZN(n1120) );
NAND2_X1 U806 ( .A1(n1125), .A2(n1126), .ZN(n1103) );
NAND4_X1 U807 ( .A1(n1127), .A2(n1128), .A3(n1129), .A4(n1130), .ZN(n1098) );
NAND3_X1 U808 ( .A1(n1105), .A2(n1131), .A3(n1107), .ZN(n1128) );
NAND3_X1 U809 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NAND2_X1 U810 ( .A1(n1119), .A2(n1135), .ZN(n1134) );
NAND3_X1 U811 ( .A1(n1114), .A2(n1136), .A3(n1113), .ZN(n1133) );
NAND2_X1 U812 ( .A1(n1117), .A2(n1137), .ZN(n1132) );
NAND2_X1 U813 ( .A1(n1125), .A2(n1138), .ZN(n1127) );
AND3_X1 U814 ( .A1(n1117), .A2(n1113), .A3(n1107), .ZN(n1125) );
INV_X1 U815 ( .A(n1139), .ZN(n1107) );
AND2_X1 U816 ( .A1(n1119), .A2(n1114), .ZN(n1117) );
NOR3_X1 U817 ( .A1(n1140), .A2(G953), .A3(n1141), .ZN(n1096) );
INV_X1 U818 ( .A(n1129), .ZN(n1141) );
NAND4_X1 U819 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1129) );
NOR4_X1 U820 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145) );
XOR2_X1 U821 ( .A(G475), .B(n1150), .Z(n1149) );
XNOR2_X1 U822 ( .A(n1151), .B(n1152), .ZN(n1148) );
XOR2_X1 U823 ( .A(n1153), .B(KEYINPUT51), .Z(n1152) );
XOR2_X1 U824 ( .A(n1154), .B(n1155), .Z(n1147) );
XNOR2_X1 U825 ( .A(KEYINPUT36), .B(KEYINPUT20), .ZN(n1154) );
XOR2_X1 U826 ( .A(n1156), .B(G472), .Z(n1146) );
NAND2_X1 U827 ( .A1(KEYINPUT14), .A2(n1157), .ZN(n1156) );
NOR2_X1 U828 ( .A1(n1115), .A2(n1112), .ZN(n1144) );
XOR2_X1 U829 ( .A(n1158), .B(n1159), .Z(n1143) );
NAND2_X1 U830 ( .A1(KEYINPUT5), .A2(n1160), .ZN(n1159) );
XOR2_X1 U831 ( .A(n1161), .B(n1162), .Z(n1142) );
NAND2_X1 U832 ( .A1(KEYINPUT47), .A2(n1163), .ZN(n1162) );
XOR2_X1 U833 ( .A(n1101), .B(KEYINPUT15), .Z(n1140) );
INV_X1 U834 ( .A(G952), .ZN(n1101) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(G72) );
NOR3_X1 U836 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U838 ( .A1(n1171), .A2(n1172), .ZN(n1169) );
NOR2_X1 U839 ( .A1(G953), .A2(n1173), .ZN(n1172) );
NOR2_X1 U840 ( .A1(n1130), .A2(n1174), .ZN(n1171) );
AND4_X1 U841 ( .A1(n1170), .A2(KEYINPUT55), .A3(n1130), .A4(n1173), .ZN(n1167) );
NAND2_X1 U842 ( .A1(n1175), .A2(n1176), .ZN(n1170) );
NAND3_X1 U843 ( .A1(KEYINPUT28), .A2(n1177), .A3(n1178), .ZN(n1176) );
XOR2_X1 U844 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U845 ( .A1(G125), .A2(n1181), .ZN(n1180) );
NAND2_X1 U846 ( .A1(n1182), .A2(n1183), .ZN(n1175) );
NAND2_X1 U847 ( .A1(KEYINPUT28), .A2(n1177), .ZN(n1183) );
XOR2_X1 U848 ( .A(n1179), .B(n1184), .Z(n1182) );
NOR2_X1 U849 ( .A1(n1185), .A2(n1181), .ZN(n1184) );
INV_X1 U850 ( .A(KEYINPUT60), .ZN(n1181) );
XOR2_X1 U851 ( .A(n1186), .B(n1187), .Z(n1179) );
XOR2_X1 U852 ( .A(n1188), .B(n1189), .Z(n1187) );
NOR2_X1 U853 ( .A1(G131), .A2(KEYINPUT22), .ZN(n1188) );
XOR2_X1 U854 ( .A(n1190), .B(n1191), .Z(n1186) );
NOR2_X1 U855 ( .A1(G134), .A2(KEYINPUT10), .ZN(n1191) );
NOR2_X1 U856 ( .A1(KEYINPUT55), .A2(n1192), .ZN(n1166) );
AND2_X1 U857 ( .A1(n1130), .A2(n1173), .ZN(n1192) );
NAND3_X1 U858 ( .A1(G953), .A2(n1193), .A3(KEYINPUT0), .ZN(n1164) );
NAND2_X1 U859 ( .A1(G900), .A2(G227), .ZN(n1193) );
NAND2_X1 U860 ( .A1(n1194), .A2(n1195), .ZN(G69) );
NAND4_X1 U861 ( .A1(KEYINPUT9), .A2(G953), .A3(n1196), .A4(n1197), .ZN(n1195) );
NAND2_X1 U862 ( .A1(n1198), .A2(n1199), .ZN(n1194) );
NAND2_X1 U863 ( .A1(n1200), .A2(n1197), .ZN(n1199) );
OR2_X1 U864 ( .A1(n1201), .A2(n1202), .ZN(n1197) );
XNOR2_X1 U865 ( .A(KEYINPUT9), .B(n1203), .ZN(n1200) );
NAND2_X1 U866 ( .A1(n1201), .A2(n1202), .ZN(n1203) );
NAND2_X1 U867 ( .A1(n1204), .A2(n1205), .ZN(n1201) );
NAND2_X1 U868 ( .A1(G953), .A2(n1206), .ZN(n1205) );
XOR2_X1 U869 ( .A(n1207), .B(n1208), .Z(n1204) );
NAND2_X1 U870 ( .A1(G953), .A2(n1196), .ZN(n1198) );
NAND2_X1 U871 ( .A1(G898), .A2(G224), .ZN(n1196) );
NOR2_X1 U872 ( .A1(n1209), .A2(n1210), .ZN(G66) );
NOR3_X1 U873 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
NOR3_X1 U874 ( .A1(n1214), .A2(n1158), .A3(n1215), .ZN(n1213) );
NOR2_X1 U875 ( .A1(n1216), .A2(n1217), .ZN(n1212) );
NOR2_X1 U876 ( .A1(n1218), .A2(n1158), .ZN(n1216) );
NOR2_X1 U877 ( .A1(n1209), .A2(n1219), .ZN(G63) );
NOR3_X1 U878 ( .A1(n1151), .A2(n1220), .A3(n1221), .ZN(n1219) );
AND3_X1 U879 ( .A1(n1222), .A2(G478), .A3(n1223), .ZN(n1221) );
NOR2_X1 U880 ( .A1(n1224), .A2(n1222), .ZN(n1220) );
NOR2_X1 U881 ( .A1(n1218), .A2(n1153), .ZN(n1224) );
NOR2_X1 U882 ( .A1(n1209), .A2(n1225), .ZN(G60) );
NOR3_X1 U883 ( .A1(n1150), .A2(n1226), .A3(n1227), .ZN(n1225) );
AND3_X1 U884 ( .A1(n1228), .A2(G475), .A3(n1223), .ZN(n1227) );
NOR2_X1 U885 ( .A1(n1229), .A2(n1228), .ZN(n1226) );
NOR2_X1 U886 ( .A1(n1218), .A2(n1230), .ZN(n1229) );
NAND2_X1 U887 ( .A1(n1231), .A2(n1232), .ZN(G6) );
NAND2_X1 U888 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
NAND2_X1 U889 ( .A1(n1235), .A2(G104), .ZN(n1231) );
NAND2_X1 U890 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U891 ( .A1(KEYINPUT32), .A2(n1238), .ZN(n1237) );
OR2_X1 U892 ( .A1(n1233), .A2(KEYINPUT32), .ZN(n1236) );
AND2_X1 U893 ( .A1(KEYINPUT3), .A2(n1238), .ZN(n1233) );
INV_X1 U894 ( .A(n1239), .ZN(n1238) );
NOR2_X1 U895 ( .A1(n1209), .A2(n1240), .ZN(G57) );
XOR2_X1 U896 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U897 ( .A(n1243), .B(n1244), .Z(n1242) );
NOR2_X1 U898 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U899 ( .A(KEYINPUT29), .B(n1247), .Z(n1246) );
NOR2_X1 U900 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
AND2_X1 U901 ( .A1(n1249), .A2(n1248), .ZN(n1245) );
XNOR2_X1 U902 ( .A(n1250), .B(KEYINPUT53), .ZN(n1249) );
NAND2_X1 U903 ( .A1(n1223), .A2(G472), .ZN(n1243) );
NOR2_X1 U904 ( .A1(n1209), .A2(n1251), .ZN(G54) );
XOR2_X1 U905 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U906 ( .A(n1254), .B(n1255), .Z(n1253) );
NAND2_X1 U907 ( .A1(KEYINPUT8), .A2(n1256), .ZN(n1254) );
XOR2_X1 U908 ( .A(n1257), .B(n1258), .Z(n1252) );
NOR2_X1 U909 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
XOR2_X1 U910 ( .A(KEYINPUT63), .B(n1261), .Z(n1260) );
NOR2_X1 U911 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XNOR2_X1 U912 ( .A(KEYINPUT2), .B(n1264), .ZN(n1263) );
XOR2_X1 U913 ( .A(n1265), .B(G110), .Z(n1262) );
NOR2_X1 U914 ( .A1(n1266), .A2(n1267), .ZN(n1259) );
XOR2_X1 U915 ( .A(n1268), .B(n1265), .Z(n1267) );
NAND2_X1 U916 ( .A1(KEYINPUT41), .A2(n1177), .ZN(n1265) );
XOR2_X1 U917 ( .A(KEYINPUT2), .B(n1264), .Z(n1266) );
NAND2_X1 U918 ( .A1(n1223), .A2(G469), .ZN(n1257) );
INV_X1 U919 ( .A(n1215), .ZN(n1223) );
NOR3_X1 U920 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(G51) );
NOR3_X1 U921 ( .A1(n1272), .A2(G953), .A3(G952), .ZN(n1271) );
AND2_X1 U922 ( .A1(n1272), .A2(n1209), .ZN(n1270) );
NOR2_X1 U923 ( .A1(n1130), .A2(G952), .ZN(n1209) );
INV_X1 U924 ( .A(KEYINPUT49), .ZN(n1272) );
XOR2_X1 U925 ( .A(n1273), .B(n1274), .Z(n1269) );
XOR2_X1 U926 ( .A(n1275), .B(n1276), .Z(n1273) );
NOR2_X1 U927 ( .A1(KEYINPUT43), .A2(n1277), .ZN(n1276) );
XOR2_X1 U928 ( .A(n1278), .B(n1248), .Z(n1277) );
OR2_X1 U929 ( .A1(n1215), .A2(n1161), .ZN(n1275) );
NAND2_X1 U930 ( .A1(G902), .A2(n1099), .ZN(n1215) );
INV_X1 U931 ( .A(n1218), .ZN(n1099) );
NOR2_X1 U932 ( .A1(n1202), .A2(n1173), .ZN(n1218) );
NAND4_X1 U933 ( .A1(n1279), .A2(n1280), .A3(n1281), .A4(n1282), .ZN(n1173) );
AND4_X1 U934 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1282) );
NOR2_X1 U935 ( .A1(n1287), .A2(n1288), .ZN(n1281) );
NAND2_X1 U936 ( .A1(n1119), .A2(n1289), .ZN(n1279) );
XOR2_X1 U937 ( .A(KEYINPUT38), .B(n1290), .Z(n1289) );
NAND4_X1 U938 ( .A1(n1291), .A2(n1093), .A3(n1292), .A4(n1293), .ZN(n1202) );
NOR4_X1 U939 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n1293) );
NOR2_X1 U940 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U941 ( .A(n1300), .ZN(n1296) );
NOR2_X1 U942 ( .A1(KEYINPUT62), .A2(n1301), .ZN(n1294) );
AND3_X1 U943 ( .A1(n1239), .A2(n1302), .A3(n1303), .ZN(n1292) );
NAND3_X1 U944 ( .A1(n1304), .A2(n1114), .A3(n1138), .ZN(n1239) );
NAND3_X1 U945 ( .A1(n1126), .A2(n1114), .A3(n1304), .ZN(n1093) );
NAND3_X1 U946 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1291) );
NAND2_X1 U947 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
NAND3_X1 U948 ( .A1(n1138), .A2(n1135), .A3(KEYINPUT62), .ZN(n1309) );
NAND2_X1 U949 ( .A1(n1310), .A2(n1299), .ZN(n1308) );
INV_X1 U950 ( .A(KEYINPUT12), .ZN(n1299) );
INV_X1 U951 ( .A(n1136), .ZN(n1305) );
XOR2_X1 U952 ( .A(n1280), .B(n1311), .Z(G48) );
NOR2_X1 U953 ( .A1(G146), .A2(KEYINPUT6), .ZN(n1311) );
NAND3_X1 U954 ( .A1(n1138), .A2(n1136), .A3(n1312), .ZN(n1280) );
XOR2_X1 U955 ( .A(n1287), .B(n1313), .Z(G45) );
NOR2_X1 U956 ( .A1(KEYINPUT16), .A2(n1314), .ZN(n1313) );
AND4_X1 U957 ( .A1(n1315), .A2(n1316), .A3(n1136), .A4(n1317), .ZN(n1287) );
XOR2_X1 U958 ( .A(n1177), .B(n1286), .Z(G42) );
NAND4_X1 U959 ( .A1(n1119), .A2(n1318), .A3(n1123), .A4(n1138), .ZN(n1286) );
INV_X1 U960 ( .A(G140), .ZN(n1177) );
XOR2_X1 U961 ( .A(n1190), .B(n1319), .Z(G39) );
NAND2_X1 U962 ( .A1(n1290), .A2(n1119), .ZN(n1319) );
AND2_X1 U963 ( .A1(n1312), .A2(n1105), .ZN(n1290) );
XNOR2_X1 U964 ( .A(n1320), .B(n1285), .ZN(G36) );
NAND3_X1 U965 ( .A1(n1315), .A2(n1126), .A3(n1119), .ZN(n1285) );
NAND2_X1 U966 ( .A1(KEYINPUT52), .A2(n1321), .ZN(n1320) );
XNOR2_X1 U967 ( .A(G131), .B(n1284), .ZN(G33) );
NAND3_X1 U968 ( .A1(n1315), .A2(n1138), .A3(n1119), .ZN(n1284) );
AND2_X1 U969 ( .A1(n1322), .A2(n1111), .ZN(n1119) );
XNOR2_X1 U970 ( .A(n1112), .B(KEYINPUT35), .ZN(n1322) );
AND3_X1 U971 ( .A1(n1137), .A2(n1323), .A3(n1324), .ZN(n1315) );
XOR2_X1 U972 ( .A(n1283), .B(n1325), .Z(G30) );
NAND2_X1 U973 ( .A1(KEYINPUT1), .A2(G128), .ZN(n1325) );
NAND3_X1 U974 ( .A1(n1126), .A2(n1136), .A3(n1312), .ZN(n1283) );
AND2_X1 U975 ( .A1(n1318), .A2(n1326), .ZN(n1312) );
AND3_X1 U976 ( .A1(n1137), .A2(n1323), .A3(n1124), .ZN(n1318) );
XNOR2_X1 U977 ( .A(G101), .B(n1303), .ZN(G3) );
NAND3_X1 U978 ( .A1(n1324), .A2(n1304), .A3(n1105), .ZN(n1303) );
NAND2_X1 U979 ( .A1(n1327), .A2(n1328), .ZN(G27) );
NAND2_X1 U980 ( .A1(n1288), .A2(n1185), .ZN(n1328) );
INV_X1 U981 ( .A(n1329), .ZN(n1288) );
XOR2_X1 U982 ( .A(n1330), .B(KEYINPUT19), .Z(n1327) );
NAND2_X1 U983 ( .A1(G125), .A2(n1329), .ZN(n1330) );
NAND4_X1 U984 ( .A1(n1123), .A2(n1113), .A3(n1138), .A4(n1331), .ZN(n1329) );
AND3_X1 U985 ( .A1(n1124), .A2(n1323), .A3(n1136), .ZN(n1331) );
NAND2_X1 U986 ( .A1(n1139), .A2(n1332), .ZN(n1323) );
NAND4_X1 U987 ( .A1(G953), .A2(G902), .A3(n1333), .A4(n1174), .ZN(n1332) );
INV_X1 U988 ( .A(G900), .ZN(n1174) );
XOR2_X1 U989 ( .A(n1334), .B(n1300), .Z(G24) );
NAND4_X1 U990 ( .A1(n1335), .A2(n1317), .A3(n1114), .A4(n1336), .ZN(n1300) );
AND2_X1 U991 ( .A1(n1113), .A2(n1316), .ZN(n1336) );
AND2_X1 U992 ( .A1(n1337), .A2(n1123), .ZN(n1114) );
XNOR2_X1 U993 ( .A(G119), .B(n1298), .ZN(G21) );
NAND2_X1 U994 ( .A1(n1310), .A2(n1335), .ZN(n1298) );
AND4_X1 U995 ( .A1(n1105), .A2(n1113), .A3(n1124), .A4(n1326), .ZN(n1310) );
XOR2_X1 U996 ( .A(n1338), .B(n1302), .Z(G18) );
NAND3_X1 U997 ( .A1(n1126), .A2(n1335), .A3(n1135), .ZN(n1302) );
AND2_X1 U998 ( .A1(n1317), .A2(n1339), .ZN(n1126) );
XNOR2_X1 U999 ( .A(G113), .B(n1301), .ZN(G15) );
NAND3_X1 U1000 ( .A1(n1135), .A2(n1335), .A3(n1138), .ZN(n1301) );
NOR2_X1 U1001 ( .A1(n1339), .A2(n1317), .ZN(n1138) );
AND2_X1 U1002 ( .A1(n1113), .A2(n1324), .ZN(n1135) );
AND2_X1 U1003 ( .A1(n1337), .A2(n1326), .ZN(n1324) );
INV_X1 U1004 ( .A(n1123), .ZN(n1326) );
XOR2_X1 U1005 ( .A(n1124), .B(KEYINPUT7), .Z(n1337) );
NOR2_X1 U1006 ( .A1(n1155), .A2(n1115), .ZN(n1113) );
INV_X1 U1007 ( .A(n1116), .ZN(n1155) );
NAND2_X1 U1008 ( .A1(n1340), .A2(n1341), .ZN(G12) );
NAND2_X1 U1009 ( .A1(G110), .A2(n1342), .ZN(n1341) );
XOR2_X1 U1010 ( .A(n1343), .B(KEYINPUT31), .Z(n1340) );
NAND2_X1 U1011 ( .A1(n1295), .A2(n1268), .ZN(n1343) );
INV_X1 U1012 ( .A(G110), .ZN(n1268) );
INV_X1 U1013 ( .A(n1342), .ZN(n1295) );
NAND4_X1 U1014 ( .A1(n1105), .A2(n1304), .A3(n1124), .A4(n1123), .ZN(n1342) );
XOR2_X1 U1015 ( .A(n1157), .B(n1344), .Z(n1123) );
NOR2_X1 U1016 ( .A1(KEYINPUT18), .A2(n1345), .ZN(n1344) );
INV_X1 U1017 ( .A(G472), .ZN(n1345) );
NAND2_X1 U1018 ( .A1(n1346), .A2(n1347), .ZN(n1157) );
XOR2_X1 U1019 ( .A(n1348), .B(n1256), .Z(n1346) );
XOR2_X1 U1020 ( .A(n1241), .B(n1349), .Z(n1348) );
XOR2_X1 U1021 ( .A(n1350), .B(n1351), .Z(n1241) );
XOR2_X1 U1022 ( .A(n1352), .B(n1353), .Z(n1351) );
NOR2_X1 U1023 ( .A1(G116), .A2(KEYINPUT37), .ZN(n1352) );
XOR2_X1 U1024 ( .A(n1354), .B(KEYINPUT23), .Z(n1350) );
NAND2_X1 U1025 ( .A1(n1355), .A2(G210), .ZN(n1354) );
XOR2_X1 U1026 ( .A(n1356), .B(n1211), .Z(n1124) );
INV_X1 U1027 ( .A(n1160), .ZN(n1211) );
NAND2_X1 U1028 ( .A1(n1214), .A2(n1347), .ZN(n1160) );
INV_X1 U1029 ( .A(n1217), .ZN(n1214) );
XOR2_X1 U1030 ( .A(n1357), .B(n1358), .Z(n1217) );
XOR2_X1 U1031 ( .A(n1359), .B(n1360), .Z(n1358) );
XOR2_X1 U1032 ( .A(G119), .B(n1361), .Z(n1360) );
NAND2_X1 U1033 ( .A1(KEYINPUT48), .A2(n1362), .ZN(n1359) );
XOR2_X1 U1034 ( .A(n1190), .B(n1363), .Z(n1362) );
NAND3_X1 U1035 ( .A1(n1364), .A2(G221), .A3(KEYINPUT21), .ZN(n1363) );
INV_X1 U1036 ( .A(G137), .ZN(n1190) );
XNOR2_X1 U1037 ( .A(n1365), .B(n1366), .ZN(n1357) );
NAND2_X1 U1038 ( .A1(KEYINPUT44), .A2(n1158), .ZN(n1356) );
NAND2_X1 U1039 ( .A1(G217), .A2(n1367), .ZN(n1158) );
AND2_X1 U1040 ( .A1(n1335), .A2(n1137), .ZN(n1304) );
NOR2_X1 U1041 ( .A1(n1116), .A2(n1115), .ZN(n1137) );
AND2_X1 U1042 ( .A1(G221), .A2(n1367), .ZN(n1115) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1347), .ZN(n1367) );
XOR2_X1 U1044 ( .A(n1368), .B(G469), .Z(n1116) );
NAND2_X1 U1045 ( .A1(n1369), .A2(n1347), .ZN(n1368) );
XOR2_X1 U1046 ( .A(n1370), .B(n1371), .Z(n1369) );
XOR2_X1 U1047 ( .A(n1255), .B(n1366), .Z(n1371) );
XOR2_X1 U1048 ( .A(G110), .B(G140), .Z(n1366) );
XOR2_X1 U1049 ( .A(n1372), .B(n1189), .Z(n1255) );
XNOR2_X1 U1050 ( .A(n1373), .B(n1374), .ZN(n1189) );
XOR2_X1 U1051 ( .A(n1361), .B(KEYINPUT42), .Z(n1373) );
XOR2_X1 U1052 ( .A(n1375), .B(n1376), .Z(n1372) );
NAND2_X1 U1053 ( .A1(KEYINPUT40), .A2(n1377), .ZN(n1375) );
XOR2_X1 U1054 ( .A(G107), .B(G104), .Z(n1377) );
XOR2_X1 U1055 ( .A(n1378), .B(n1256), .Z(n1370) );
INV_X1 U1056 ( .A(n1250), .ZN(n1256) );
XOR2_X1 U1057 ( .A(n1379), .B(n1380), .Z(n1250) );
XOR2_X1 U1058 ( .A(KEYINPUT11), .B(G137), .Z(n1380) );
XOR2_X1 U1059 ( .A(G131), .B(n1321), .Z(n1379) );
INV_X1 U1060 ( .A(G134), .ZN(n1321) );
XOR2_X1 U1061 ( .A(n1264), .B(KEYINPUT39), .Z(n1378) );
NAND2_X1 U1062 ( .A1(G227), .A2(n1130), .ZN(n1264) );
AND2_X1 U1063 ( .A1(n1136), .A2(n1306), .ZN(n1335) );
NAND2_X1 U1064 ( .A1(n1381), .A2(n1139), .ZN(n1306) );
NAND3_X1 U1065 ( .A1(n1333), .A2(n1130), .A3(G952), .ZN(n1139) );
NAND4_X1 U1066 ( .A1(G953), .A2(G902), .A3(n1333), .A4(n1206), .ZN(n1381) );
INV_X1 U1067 ( .A(G898), .ZN(n1206) );
NAND2_X1 U1068 ( .A1(G237), .A2(G234), .ZN(n1333) );
NOR2_X1 U1069 ( .A1(n1111), .A2(n1112), .ZN(n1136) );
AND2_X1 U1070 ( .A1(G214), .A2(n1382), .ZN(n1112) );
XNOR2_X1 U1071 ( .A(n1163), .B(n1161), .ZN(n1111) );
NAND2_X1 U1072 ( .A1(G210), .A2(n1382), .ZN(n1161) );
NAND2_X1 U1073 ( .A1(n1383), .A2(n1347), .ZN(n1382) );
INV_X1 U1074 ( .A(G237), .ZN(n1383) );
NAND2_X1 U1075 ( .A1(n1384), .A2(n1347), .ZN(n1163) );
INV_X1 U1076 ( .A(G902), .ZN(n1347) );
XOR2_X1 U1077 ( .A(n1385), .B(n1386), .Z(n1384) );
XOR2_X1 U1078 ( .A(KEYINPUT58), .B(n1387), .Z(n1386) );
NOR2_X1 U1079 ( .A1(KEYINPUT17), .A2(n1349), .ZN(n1387) );
INV_X1 U1080 ( .A(n1248), .ZN(n1349) );
XNOR2_X1 U1081 ( .A(n1374), .B(n1388), .ZN(n1248) );
NOR2_X1 U1082 ( .A1(KEYINPUT59), .A2(n1361), .ZN(n1388) );
INV_X1 U1083 ( .A(G128), .ZN(n1361) );
XOR2_X1 U1084 ( .A(G146), .B(G143), .Z(n1374) );
XNOR2_X1 U1085 ( .A(n1274), .B(n1278), .ZN(n1385) );
XNOR2_X1 U1086 ( .A(n1185), .B(n1389), .ZN(n1278) );
AND2_X1 U1087 ( .A1(n1130), .A2(G224), .ZN(n1389) );
INV_X1 U1088 ( .A(G125), .ZN(n1185) );
XNOR2_X1 U1089 ( .A(n1390), .B(n1391), .ZN(n1274) );
INV_X1 U1090 ( .A(n1207), .ZN(n1391) );
XOR2_X1 U1091 ( .A(n1392), .B(n1393), .Z(n1207) );
XOR2_X1 U1092 ( .A(KEYINPUT30), .B(G116), .Z(n1393) );
XOR2_X1 U1093 ( .A(n1394), .B(n1353), .Z(n1392) );
XNOR2_X1 U1094 ( .A(n1395), .B(n1376), .ZN(n1353) );
XOR2_X1 U1095 ( .A(G101), .B(KEYINPUT46), .Z(n1376) );
XNOR2_X1 U1096 ( .A(G113), .B(G119), .ZN(n1395) );
NAND3_X1 U1097 ( .A1(n1396), .A2(n1397), .A3(n1398), .ZN(n1394) );
NAND2_X1 U1098 ( .A1(KEYINPUT27), .A2(G104), .ZN(n1398) );
OR3_X1 U1099 ( .A1(n1399), .A2(KEYINPUT27), .A3(G107), .ZN(n1397) );
NAND2_X1 U1100 ( .A1(G107), .A2(n1399), .ZN(n1396) );
NAND2_X1 U1101 ( .A1(KEYINPUT25), .A2(n1234), .ZN(n1399) );
INV_X1 U1102 ( .A(G104), .ZN(n1234) );
NAND2_X1 U1103 ( .A1(KEYINPUT54), .A2(n1208), .ZN(n1390) );
XOR2_X1 U1104 ( .A(G122), .B(G110), .Z(n1208) );
NOR2_X1 U1105 ( .A1(n1317), .A2(n1316), .ZN(n1105) );
INV_X1 U1106 ( .A(n1339), .ZN(n1316) );
NAND3_X1 U1107 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n1339) );
NAND2_X1 U1108 ( .A1(KEYINPUT56), .A2(n1230), .ZN(n1402) );
NAND3_X1 U1109 ( .A1(n1403), .A2(n1404), .A3(n1405), .ZN(n1401) );
INV_X1 U1110 ( .A(KEYINPUT56), .ZN(n1404) );
OR2_X1 U1111 ( .A1(n1405), .A2(n1403), .ZN(n1400) );
NOR2_X1 U1112 ( .A1(KEYINPUT34), .A2(n1230), .ZN(n1403) );
INV_X1 U1113 ( .A(G475), .ZN(n1230) );
XNOR2_X1 U1114 ( .A(n1150), .B(KEYINPUT45), .ZN(n1405) );
NOR2_X1 U1115 ( .A1(n1228), .A2(G902), .ZN(n1150) );
XNOR2_X1 U1116 ( .A(n1406), .B(n1407), .ZN(n1228) );
XOR2_X1 U1117 ( .A(G122), .B(G113), .Z(n1407) );
XOR2_X1 U1118 ( .A(n1408), .B(G104), .Z(n1406) );
NAND2_X1 U1119 ( .A1(KEYINPUT24), .A2(n1409), .ZN(n1408) );
XOR2_X1 U1120 ( .A(n1410), .B(n1411), .Z(n1409) );
XOR2_X1 U1121 ( .A(n1412), .B(n1413), .Z(n1411) );
NOR2_X1 U1122 ( .A1(KEYINPUT61), .A2(n1414), .ZN(n1413) );
XOR2_X1 U1123 ( .A(G140), .B(n1365), .Z(n1414) );
XOR2_X1 U1124 ( .A(G146), .B(G125), .Z(n1365) );
NAND2_X1 U1125 ( .A1(n1355), .A2(G214), .ZN(n1412) );
NOR2_X1 U1126 ( .A1(G953), .A2(G237), .ZN(n1355) );
XOR2_X1 U1127 ( .A(G131), .B(n1314), .Z(n1410) );
INV_X1 U1128 ( .A(G143), .ZN(n1314) );
NAND3_X1 U1129 ( .A1(n1415), .A2(n1416), .A3(n1417), .ZN(n1317) );
NAND2_X1 U1130 ( .A1(KEYINPUT33), .A2(n1151), .ZN(n1417) );
OR3_X1 U1131 ( .A1(n1151), .A2(KEYINPUT33), .A3(n1153), .ZN(n1416) );
NAND2_X1 U1132 ( .A1(n1418), .A2(n1153), .ZN(n1415) );
INV_X1 U1133 ( .A(G478), .ZN(n1153) );
NAND2_X1 U1134 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
INV_X1 U1135 ( .A(KEYINPUT33), .ZN(n1420) );
XOR2_X1 U1136 ( .A(KEYINPUT50), .B(n1151), .Z(n1419) );
NOR2_X1 U1137 ( .A1(n1222), .A2(G902), .ZN(n1151) );
XNOR2_X1 U1138 ( .A(n1421), .B(n1422), .ZN(n1222) );
XOR2_X1 U1139 ( .A(n1423), .B(n1424), .Z(n1422) );
XOR2_X1 U1140 ( .A(n1338), .B(n1425), .Z(n1424) );
NOR2_X1 U1141 ( .A1(G107), .A2(KEYINPUT57), .ZN(n1425) );
INV_X1 U1142 ( .A(G116), .ZN(n1338) );
NAND2_X1 U1143 ( .A1(G217), .A2(n1364), .ZN(n1423) );
AND2_X1 U1144 ( .A1(G234), .A2(n1130), .ZN(n1364) );
INV_X1 U1145 ( .A(G953), .ZN(n1130) );
XOR2_X1 U1146 ( .A(n1426), .B(n1427), .Z(n1421) );
XOR2_X1 U1147 ( .A(G143), .B(G134), .Z(n1427) );
XOR2_X1 U1148 ( .A(n1334), .B(G128), .Z(n1426) );
INV_X1 U1149 ( .A(G122), .ZN(n1334) );
endmodule


