//Key = 0000100010110010001111111101010100011000110111100001110110111000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324;

XOR2_X1 U731 ( .A(n1010), .B(n1011), .Z(G9) );
NOR2_X1 U732 ( .A1(n1012), .A2(n1013), .ZN(G75) );
XOR2_X1 U733 ( .A(KEYINPUT62), .B(n1014), .Z(n1013) );
NOR3_X1 U734 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NAND3_X1 U735 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n1015) );
INV_X1 U736 ( .A(n1021), .ZN(n1020) );
NAND4_X1 U737 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1019) );
NAND2_X1 U738 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U739 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
NAND2_X1 U740 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND2_X1 U741 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1026) );
NAND2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
OR2_X1 U744 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND4_X1 U745 ( .A1(n1028), .A2(n1034), .A3(n1040), .A4(n1041), .ZN(n1018) );
NAND2_X1 U746 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U747 ( .A1(n1024), .A2(n1044), .A3(n1045), .ZN(n1042) );
INV_X1 U748 ( .A(KEYINPUT19), .ZN(n1044) );
NAND3_X1 U749 ( .A1(n1046), .A2(n1047), .A3(n1022), .ZN(n1040) );
INV_X1 U750 ( .A(n1043), .ZN(n1022) );
NAND2_X1 U751 ( .A1(n1024), .A2(n1048), .ZN(n1047) );
NAND2_X1 U752 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U753 ( .A1(KEYINPUT19), .A2(n1045), .ZN(n1050) );
NAND2_X1 U754 ( .A1(n1023), .A2(n1051), .ZN(n1046) );
NAND2_X1 U755 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U756 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XOR2_X1 U757 ( .A(KEYINPUT53), .B(n1056), .Z(n1055) );
NOR2_X1 U758 ( .A1(G952), .A2(n1021), .ZN(n1012) );
NAND2_X1 U759 ( .A1(n1057), .A2(n1058), .ZN(n1021) );
NAND4_X1 U760 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
NOR4_X1 U761 ( .A1(n1054), .A2(n1063), .A3(n1033), .A4(n1064), .ZN(n1062) );
XNOR2_X1 U762 ( .A(n1065), .B(n1066), .ZN(n1063) );
NAND2_X1 U763 ( .A1(KEYINPUT14), .A2(n1067), .ZN(n1065) );
INV_X1 U764 ( .A(n1068), .ZN(n1054) );
NOR3_X1 U765 ( .A1(n1056), .A2(n1069), .A3(n1070), .ZN(n1061) );
NOR2_X1 U766 ( .A1(KEYINPUT41), .A2(n1071), .ZN(n1070) );
NOR2_X1 U767 ( .A1(n1039), .A2(n1038), .ZN(n1071) );
AND2_X1 U768 ( .A1(n1072), .A2(KEYINPUT41), .ZN(n1069) );
NAND2_X1 U769 ( .A1(n1073), .A2(n1074), .ZN(n1060) );
INV_X1 U770 ( .A(KEYINPUT31), .ZN(n1074) );
NAND2_X1 U771 ( .A1(G478), .A2(n1075), .ZN(n1073) );
NAND2_X1 U772 ( .A1(KEYINPUT31), .A2(n1076), .ZN(n1059) );
XOR2_X1 U773 ( .A(n1077), .B(n1078), .Z(G72) );
XOR2_X1 U774 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U775 ( .A1(n1081), .A2(n1057), .ZN(n1080) );
XOR2_X1 U776 ( .A(n1082), .B(KEYINPUT21), .Z(n1081) );
NAND2_X1 U777 ( .A1(G900), .A2(G227), .ZN(n1082) );
NAND2_X1 U778 ( .A1(n1083), .A2(n1016), .ZN(n1079) );
XOR2_X1 U779 ( .A(KEYINPUT43), .B(G953), .Z(n1083) );
NAND2_X1 U780 ( .A1(n1084), .A2(n1085), .ZN(n1077) );
NAND2_X1 U781 ( .A1(G953), .A2(n1086), .ZN(n1085) );
XOR2_X1 U782 ( .A(n1087), .B(n1088), .Z(n1084) );
XNOR2_X1 U783 ( .A(n1089), .B(n1090), .ZN(n1088) );
NAND2_X1 U784 ( .A1(n1091), .A2(KEYINPUT46), .ZN(n1089) );
XOR2_X1 U785 ( .A(n1092), .B(G131), .Z(n1091) );
NAND3_X1 U786 ( .A1(n1093), .A2(n1094), .A3(n1095), .ZN(n1092) );
NAND2_X1 U787 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
INV_X1 U788 ( .A(KEYINPUT25), .ZN(n1097) );
NAND3_X1 U789 ( .A1(KEYINPUT25), .A2(n1098), .A3(n1099), .ZN(n1094) );
OR2_X1 U790 ( .A1(n1099), .A2(n1098), .ZN(n1093) );
NOR2_X1 U791 ( .A1(KEYINPUT9), .A2(n1096), .ZN(n1098) );
XNOR2_X1 U792 ( .A(KEYINPUT32), .B(n1100), .ZN(n1087) );
NOR2_X1 U793 ( .A1(KEYINPUT49), .A2(n1101), .ZN(n1100) );
XOR2_X1 U794 ( .A(KEYINPUT12), .B(n1102), .Z(n1101) );
XOR2_X1 U795 ( .A(n1103), .B(n1104), .Z(G69) );
XOR2_X1 U796 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U797 ( .A1(G953), .A2(n1107), .ZN(n1106) );
NAND2_X1 U798 ( .A1(G898), .A2(G224), .ZN(n1107) );
NAND2_X1 U799 ( .A1(n1108), .A2(n1109), .ZN(n1105) );
NAND2_X1 U800 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U801 ( .A(n1111), .B(KEYINPUT52), .Z(n1108) );
AND2_X1 U802 ( .A1(n1017), .A2(n1057), .ZN(n1103) );
NOR2_X1 U803 ( .A1(n1112), .A2(n1113), .ZN(G66) );
XOR2_X1 U804 ( .A(n1114), .B(n1115), .Z(n1113) );
NOR2_X1 U805 ( .A1(KEYINPUT7), .A2(n1116), .ZN(n1115) );
NAND2_X1 U806 ( .A1(n1117), .A2(G217), .ZN(n1114) );
NOR2_X1 U807 ( .A1(n1112), .A2(n1118), .ZN(G63) );
XNOR2_X1 U808 ( .A(n1119), .B(n1120), .ZN(n1118) );
AND2_X1 U809 ( .A1(G478), .A2(n1117), .ZN(n1119) );
NOR2_X1 U810 ( .A1(n1112), .A2(n1121), .ZN(G60) );
XOR2_X1 U811 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND3_X1 U812 ( .A1(n1117), .A2(G475), .A3(KEYINPUT24), .ZN(n1122) );
XOR2_X1 U813 ( .A(n1124), .B(n1125), .Z(G6) );
NOR2_X1 U814 ( .A1(KEYINPUT30), .A2(n1126), .ZN(n1125) );
NOR2_X1 U815 ( .A1(n1112), .A2(n1127), .ZN(G57) );
XOR2_X1 U816 ( .A(n1128), .B(n1129), .Z(n1127) );
XOR2_X1 U817 ( .A(n1130), .B(n1131), .Z(n1129) );
NAND2_X1 U818 ( .A1(KEYINPUT45), .A2(n1132), .ZN(n1130) );
XOR2_X1 U819 ( .A(n1133), .B(n1134), .Z(n1128) );
NOR2_X1 U820 ( .A1(n1067), .A2(n1135), .ZN(n1134) );
INV_X1 U821 ( .A(G472), .ZN(n1067) );
NAND2_X1 U822 ( .A1(n1136), .A2(n1137), .ZN(n1133) );
NAND2_X1 U823 ( .A1(n1138), .A2(G101), .ZN(n1137) );
XOR2_X1 U824 ( .A(KEYINPUT40), .B(n1139), .Z(n1136) );
NOR2_X1 U825 ( .A1(n1138), .A2(G101), .ZN(n1139) );
NOR2_X1 U826 ( .A1(n1112), .A2(n1140), .ZN(G54) );
XOR2_X1 U827 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U828 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U829 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
AND3_X1 U830 ( .A1(KEYINPUT38), .A2(n1147), .A3(G140), .ZN(n1146) );
NOR2_X1 U831 ( .A1(KEYINPUT38), .A2(n1148), .ZN(n1145) );
AND2_X1 U832 ( .A1(G469), .A2(n1117), .ZN(n1143) );
INV_X1 U833 ( .A(n1135), .ZN(n1117) );
XNOR2_X1 U834 ( .A(n1149), .B(n1150), .ZN(n1141) );
NOR2_X1 U835 ( .A1(KEYINPUT50), .A2(n1151), .ZN(n1150) );
XNOR2_X1 U836 ( .A(n1152), .B(n1153), .ZN(n1151) );
XNOR2_X1 U837 ( .A(n1090), .B(n1154), .ZN(n1153) );
NOR2_X1 U838 ( .A1(n1112), .A2(n1155), .ZN(G51) );
NOR3_X1 U839 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(n1155) );
NOR3_X1 U840 ( .A1(n1159), .A2(n1160), .A3(n1161), .ZN(n1158) );
NOR3_X1 U841 ( .A1(n1135), .A2(KEYINPUT6), .A3(n1162), .ZN(n1160) );
NOR2_X1 U842 ( .A1(KEYINPUT4), .A2(n1163), .ZN(n1157) );
NOR3_X1 U843 ( .A1(n1135), .A2(n1164), .A3(n1162), .ZN(n1156) );
NOR2_X1 U844 ( .A1(n1165), .A2(n1159), .ZN(n1164) );
INV_X1 U845 ( .A(KEYINPUT4), .ZN(n1159) );
NOR2_X1 U846 ( .A1(KEYINPUT6), .A2(n1163), .ZN(n1165) );
INV_X1 U847 ( .A(n1161), .ZN(n1163) );
XOR2_X1 U848 ( .A(n1166), .B(n1167), .Z(n1161) );
XOR2_X1 U849 ( .A(n1168), .B(n1169), .Z(n1166) );
NAND2_X1 U850 ( .A1(G902), .A2(n1170), .ZN(n1135) );
OR2_X1 U851 ( .A1(n1017), .A2(n1016), .ZN(n1170) );
NAND4_X1 U852 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1016) );
NOR4_X1 U853 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
INV_X1 U854 ( .A(n1179), .ZN(n1178) );
AND2_X1 U855 ( .A1(n1180), .A2(n1181), .ZN(n1173) );
NAND3_X1 U856 ( .A1(n1182), .A2(n1183), .A3(n1028), .ZN(n1172) );
NAND2_X1 U857 ( .A1(n1184), .A2(n1185), .ZN(n1171) );
XOR2_X1 U858 ( .A(n1186), .B(KEYINPUT36), .Z(n1184) );
NAND4_X1 U859 ( .A1(n1187), .A2(n1045), .A3(n1188), .A4(n1189), .ZN(n1186) );
XOR2_X1 U860 ( .A(KEYINPUT3), .B(n1190), .Z(n1188) );
NAND2_X1 U861 ( .A1(n1191), .A2(n1192), .ZN(n1017) );
NOR4_X1 U862 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1124), .ZN(n1192) );
AND3_X1 U863 ( .A1(n1196), .A2(n1034), .A3(n1183), .ZN(n1124) );
INV_X1 U864 ( .A(n1197), .ZN(n1193) );
NOR4_X1 U865 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1191) );
NOR3_X1 U866 ( .A1(n1030), .A2(n1202), .A3(n1203), .ZN(n1201) );
XOR2_X1 U867 ( .A(n1204), .B(KEYINPUT16), .Z(n1202) );
INV_X1 U868 ( .A(n1011), .ZN(n1198) );
NAND3_X1 U869 ( .A1(n1045), .A2(n1034), .A3(n1196), .ZN(n1011) );
NOR2_X1 U870 ( .A1(n1057), .A2(G952), .ZN(n1112) );
XOR2_X1 U871 ( .A(G146), .B(n1175), .Z(G48) );
NOR2_X1 U872 ( .A1(n1205), .A2(n1049), .ZN(n1175) );
XOR2_X1 U873 ( .A(n1206), .B(n1181), .Z(G45) );
NAND4_X1 U874 ( .A1(n1182), .A2(n1185), .A3(n1076), .A4(n1064), .ZN(n1181) );
INV_X1 U875 ( .A(n1207), .ZN(n1182) );
XNOR2_X1 U876 ( .A(G140), .B(n1180), .ZN(G42) );
NAND3_X1 U877 ( .A1(n1032), .A2(n1183), .A3(n1208), .ZN(n1180) );
XOR2_X1 U878 ( .A(n1099), .B(n1179), .Z(G39) );
NAND3_X1 U879 ( .A1(n1023), .A2(n1189), .A3(n1208), .ZN(n1179) );
NOR3_X1 U880 ( .A1(n1209), .A2(n1052), .A3(n1072), .ZN(n1208) );
XOR2_X1 U881 ( .A(G134), .B(n1177), .Z(G36) );
NOR3_X1 U882 ( .A1(n1207), .A2(n1210), .A3(n1072), .ZN(n1177) );
XOR2_X1 U883 ( .A(G131), .B(n1211), .Z(G33) );
NOR3_X1 U884 ( .A1(n1207), .A2(n1212), .A3(n1049), .ZN(n1211) );
XOR2_X1 U885 ( .A(n1072), .B(KEYINPUT37), .Z(n1212) );
INV_X1 U886 ( .A(n1028), .ZN(n1072) );
NOR2_X1 U887 ( .A1(n1039), .A2(n1213), .ZN(n1028) );
INV_X1 U888 ( .A(n1038), .ZN(n1213) );
NAND3_X1 U889 ( .A1(n1190), .A2(n1214), .A3(n1215), .ZN(n1207) );
XOR2_X1 U890 ( .A(G128), .B(n1216), .Z(G30) );
NOR3_X1 U891 ( .A1(n1205), .A2(KEYINPUT34), .A3(n1210), .ZN(n1216) );
NAND4_X1 U892 ( .A1(n1187), .A2(n1190), .A3(n1185), .A4(n1189), .ZN(n1205) );
INV_X1 U893 ( .A(n1209), .ZN(n1187) );
XOR2_X1 U894 ( .A(G101), .B(n1217), .Z(G3) );
NOR4_X1 U895 ( .A1(KEYINPUT48), .A2(n1203), .A3(n1204), .A4(n1030), .ZN(n1217) );
INV_X1 U896 ( .A(n1215), .ZN(n1030) );
XNOR2_X1 U897 ( .A(n1176), .B(n1218), .ZN(G27) );
XOR2_X1 U898 ( .A(n1219), .B(KEYINPUT33), .Z(n1218) );
AND4_X1 U899 ( .A1(n1185), .A2(n1024), .A3(n1032), .A4(n1220), .ZN(n1176) );
NOR2_X1 U900 ( .A1(n1049), .A2(n1209), .ZN(n1220) );
NAND2_X1 U901 ( .A1(n1033), .A2(n1214), .ZN(n1209) );
NAND2_X1 U902 ( .A1(n1221), .A2(n1043), .ZN(n1214) );
XOR2_X1 U903 ( .A(n1222), .B(KEYINPUT28), .Z(n1221) );
NAND4_X1 U904 ( .A1(G953), .A2(G902), .A3(n1223), .A4(n1086), .ZN(n1222) );
INV_X1 U905 ( .A(G900), .ZN(n1086) );
NAND2_X1 U906 ( .A1(n1224), .A2(n1225), .ZN(G24) );
OR2_X1 U907 ( .A1(n1226), .A2(G122), .ZN(n1225) );
NAND2_X1 U908 ( .A1(n1227), .A2(G122), .ZN(n1224) );
NAND2_X1 U909 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U910 ( .A1(n1195), .A2(n1230), .ZN(n1229) );
INV_X1 U911 ( .A(KEYINPUT29), .ZN(n1230) );
NAND2_X1 U912 ( .A1(KEYINPUT29), .A2(n1226), .ZN(n1228) );
NAND2_X1 U913 ( .A1(KEYINPUT35), .A2(n1195), .ZN(n1226) );
AND4_X1 U914 ( .A1(n1231), .A2(n1034), .A3(n1076), .A4(n1064), .ZN(n1195) );
NOR2_X1 U915 ( .A1(n1033), .A2(n1189), .ZN(n1034) );
NAND2_X1 U916 ( .A1(n1232), .A2(n1233), .ZN(G21) );
NAND2_X1 U917 ( .A1(n1200), .A2(n1234), .ZN(n1233) );
INV_X1 U918 ( .A(n1235), .ZN(n1200) );
XOR2_X1 U919 ( .A(n1236), .B(KEYINPUT61), .Z(n1232) );
NAND2_X1 U920 ( .A1(G119), .A2(n1235), .ZN(n1236) );
NAND4_X1 U921 ( .A1(n1231), .A2(n1023), .A3(n1189), .A4(n1033), .ZN(n1235) );
INV_X1 U922 ( .A(n1032), .ZN(n1189) );
XOR2_X1 U923 ( .A(G116), .B(n1199), .Z(G18) );
AND3_X1 U924 ( .A1(n1215), .A2(n1045), .A3(n1231), .ZN(n1199) );
INV_X1 U925 ( .A(n1210), .ZN(n1045) );
NAND2_X1 U926 ( .A1(n1076), .A2(n1237), .ZN(n1210) );
INV_X1 U927 ( .A(n1238), .ZN(n1076) );
XOR2_X1 U928 ( .A(G113), .B(n1194), .Z(G15) );
AND3_X1 U929 ( .A1(n1215), .A2(n1183), .A3(n1231), .ZN(n1194) );
AND3_X1 U930 ( .A1(n1024), .A2(n1239), .A3(n1185), .ZN(n1231) );
NAND2_X1 U931 ( .A1(n1240), .A2(n1241), .ZN(n1024) );
OR2_X1 U932 ( .A1(n1052), .A2(KEYINPUT53), .ZN(n1241) );
NAND3_X1 U933 ( .A1(n1242), .A2(n1068), .A3(KEYINPUT53), .ZN(n1240) );
INV_X1 U934 ( .A(n1049), .ZN(n1183) );
NAND2_X1 U935 ( .A1(n1238), .A2(n1064), .ZN(n1049) );
NOR2_X1 U936 ( .A1(n1033), .A2(n1032), .ZN(n1215) );
XNOR2_X1 U937 ( .A(n1243), .B(n1147), .ZN(G12) );
NAND2_X1 U938 ( .A1(KEYINPUT56), .A2(n1197), .ZN(n1243) );
NAND4_X1 U939 ( .A1(n1023), .A2(n1196), .A3(n1032), .A4(n1033), .ZN(n1197) );
XNOR2_X1 U940 ( .A(n1244), .B(n1245), .ZN(n1033) );
NOR2_X1 U941 ( .A1(n1116), .A2(n1246), .ZN(n1245) );
XOR2_X1 U942 ( .A(KEYINPUT63), .B(G902), .Z(n1246) );
XNOR2_X1 U943 ( .A(n1247), .B(n1248), .ZN(n1116) );
XNOR2_X1 U944 ( .A(n1148), .B(n1249), .ZN(n1248) );
XOR2_X1 U945 ( .A(n1250), .B(n1251), .Z(n1249) );
NAND2_X1 U946 ( .A1(KEYINPUT10), .A2(n1219), .ZN(n1250) );
XOR2_X1 U947 ( .A(n1252), .B(n1253), .Z(n1247) );
NOR2_X1 U948 ( .A1(KEYINPUT42), .A2(n1254), .ZN(n1253) );
XOR2_X1 U949 ( .A(n1255), .B(n1256), .Z(n1254) );
XOR2_X1 U950 ( .A(KEYINPUT2), .B(G137), .Z(n1256) );
NAND2_X1 U951 ( .A1(n1257), .A2(G221), .ZN(n1255) );
XOR2_X1 U952 ( .A(n1234), .B(KEYINPUT39), .Z(n1252) );
INV_X1 U953 ( .A(G119), .ZN(n1234) );
NAND2_X1 U954 ( .A1(G217), .A2(n1258), .ZN(n1244) );
XOR2_X1 U955 ( .A(n1066), .B(G472), .Z(n1032) );
NAND2_X1 U956 ( .A1(n1259), .A2(n1260), .ZN(n1066) );
XNOR2_X1 U957 ( .A(n1132), .B(n1261), .ZN(n1259) );
XOR2_X1 U958 ( .A(n1131), .B(n1262), .Z(n1261) );
NOR2_X1 U959 ( .A1(KEYINPUT15), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U960 ( .A(n1138), .B(n1264), .ZN(n1263) );
XOR2_X1 U961 ( .A(KEYINPUT54), .B(G101), .Z(n1264) );
AND3_X1 U962 ( .A1(n1265), .A2(n1057), .A3(G210), .ZN(n1138) );
XNOR2_X1 U963 ( .A(n1152), .B(n1266), .ZN(n1131) );
XOR2_X1 U964 ( .A(G116), .B(n1267), .Z(n1266) );
INV_X1 U965 ( .A(n1203), .ZN(n1196) );
NAND3_X1 U966 ( .A1(n1185), .A2(n1239), .A3(n1190), .ZN(n1203) );
INV_X1 U967 ( .A(n1052), .ZN(n1190) );
NAND2_X1 U968 ( .A1(n1056), .A2(n1068), .ZN(n1052) );
NAND2_X1 U969 ( .A1(G221), .A2(n1258), .ZN(n1068) );
NAND2_X1 U970 ( .A1(n1268), .A2(n1260), .ZN(n1258) );
INV_X1 U971 ( .A(n1242), .ZN(n1056) );
XOR2_X1 U972 ( .A(n1269), .B(G469), .Z(n1242) );
NAND2_X1 U973 ( .A1(n1270), .A2(n1260), .ZN(n1269) );
XOR2_X1 U974 ( .A(n1271), .B(n1272), .Z(n1270) );
XNOR2_X1 U975 ( .A(n1154), .B(n1148), .ZN(n1272) );
XOR2_X1 U976 ( .A(G110), .B(G140), .Z(n1148) );
XNOR2_X1 U977 ( .A(n1273), .B(n1274), .ZN(n1154) );
XOR2_X1 U978 ( .A(G107), .B(G104), .Z(n1274) );
INV_X1 U979 ( .A(G101), .ZN(n1273) );
XOR2_X1 U980 ( .A(n1275), .B(n1276), .Z(n1271) );
NOR2_X1 U981 ( .A1(n1149), .A2(KEYINPUT47), .ZN(n1276) );
AND2_X1 U982 ( .A1(G227), .A2(n1057), .ZN(n1149) );
XNOR2_X1 U983 ( .A(n1277), .B(n1278), .ZN(n1275) );
NAND2_X1 U984 ( .A1(KEYINPUT8), .A2(n1152), .ZN(n1278) );
AND2_X1 U985 ( .A1(n1279), .A2(n1280), .ZN(n1152) );
NAND2_X1 U986 ( .A1(n1281), .A2(n1099), .ZN(n1280) );
INV_X1 U987 ( .A(G137), .ZN(n1099) );
XOR2_X1 U988 ( .A(KEYINPUT60), .B(n1282), .Z(n1281) );
NAND2_X1 U989 ( .A1(G137), .A2(n1283), .ZN(n1279) );
XNOR2_X1 U990 ( .A(n1282), .B(KEYINPUT55), .ZN(n1283) );
XOR2_X1 U991 ( .A(n1284), .B(n1096), .Z(n1282) );
NAND2_X1 U992 ( .A1(KEYINPUT20), .A2(n1090), .ZN(n1277) );
XNOR2_X1 U993 ( .A(n1285), .B(n1286), .ZN(n1090) );
XOR2_X1 U994 ( .A(G146), .B(G143), .Z(n1286) );
NAND2_X1 U995 ( .A1(KEYINPUT23), .A2(G128), .ZN(n1285) );
NAND2_X1 U996 ( .A1(n1043), .A2(n1287), .ZN(n1239) );
NAND4_X1 U997 ( .A1(G953), .A2(G902), .A3(n1223), .A4(n1110), .ZN(n1287) );
INV_X1 U998 ( .A(G898), .ZN(n1110) );
NAND3_X1 U999 ( .A1(n1223), .A2(n1057), .A3(n1288), .ZN(n1043) );
XOR2_X1 U1000 ( .A(KEYINPUT26), .B(G952), .Z(n1288) );
NAND2_X1 U1001 ( .A1(G237), .A2(n1268), .ZN(n1223) );
XNOR2_X1 U1002 ( .A(G234), .B(KEYINPUT59), .ZN(n1268) );
INV_X1 U1003 ( .A(n1036), .ZN(n1185) );
NAND2_X1 U1004 ( .A1(n1039), .A2(n1038), .ZN(n1036) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1289), .ZN(n1038) );
XOR2_X1 U1006 ( .A(n1290), .B(n1162), .Z(n1039) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1289), .ZN(n1162) );
NAND2_X1 U1008 ( .A1(n1265), .A2(n1260), .ZN(n1289) );
NAND2_X1 U1009 ( .A1(n1291), .A2(n1260), .ZN(n1290) );
XOR2_X1 U1010 ( .A(n1292), .B(n1169), .Z(n1291) );
INV_X1 U1011 ( .A(n1111), .ZN(n1169) );
XOR2_X1 U1012 ( .A(n1293), .B(n1294), .Z(n1111) );
XOR2_X1 U1013 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1014 ( .A(n1297), .B(G101), .Z(n1296) );
NAND2_X1 U1015 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
OR2_X1 U1016 ( .A1(n1147), .A2(G122), .ZN(n1299) );
XOR2_X1 U1017 ( .A(n1300), .B(KEYINPUT17), .Z(n1298) );
NAND2_X1 U1018 ( .A1(G122), .A2(n1147), .ZN(n1300) );
INV_X1 U1019 ( .A(G110), .ZN(n1147) );
XOR2_X1 U1020 ( .A(n1126), .B(KEYINPUT1), .Z(n1295) );
XNOR2_X1 U1021 ( .A(n1267), .B(n1301), .ZN(n1293) );
XNOR2_X1 U1022 ( .A(n1302), .B(n1303), .ZN(n1301) );
NOR2_X1 U1023 ( .A1(G116), .A2(KEYINPUT5), .ZN(n1303) );
NAND2_X1 U1024 ( .A1(KEYINPUT44), .A2(n1010), .ZN(n1302) );
INV_X1 U1025 ( .A(G107), .ZN(n1010) );
XOR2_X1 U1026 ( .A(G113), .B(G119), .Z(n1267) );
XOR2_X1 U1027 ( .A(n1168), .B(n1304), .Z(n1292) );
NOR2_X1 U1028 ( .A1(KEYINPUT57), .A2(n1167), .ZN(n1304) );
XNOR2_X1 U1029 ( .A(n1132), .B(n1219), .ZN(n1167) );
INV_X1 U1030 ( .A(G125), .ZN(n1219) );
XNOR2_X1 U1031 ( .A(n1305), .B(n1251), .ZN(n1132) );
XOR2_X1 U1032 ( .A(G128), .B(G146), .Z(n1251) );
NAND2_X1 U1033 ( .A1(KEYINPUT11), .A2(n1206), .ZN(n1305) );
INV_X1 U1034 ( .A(G143), .ZN(n1206) );
NAND2_X1 U1035 ( .A1(G224), .A2(n1057), .ZN(n1168) );
INV_X1 U1036 ( .A(n1204), .ZN(n1023) );
NAND2_X1 U1037 ( .A1(n1238), .A2(n1237), .ZN(n1204) );
XOR2_X1 U1038 ( .A(n1064), .B(KEYINPUT18), .Z(n1237) );
XNOR2_X1 U1039 ( .A(n1306), .B(G475), .ZN(n1064) );
NAND2_X1 U1040 ( .A1(n1123), .A2(n1260), .ZN(n1306) );
XOR2_X1 U1041 ( .A(n1307), .B(n1308), .Z(n1123) );
XOR2_X1 U1042 ( .A(n1309), .B(n1310), .Z(n1308) );
XOR2_X1 U1043 ( .A(G122), .B(G113), .Z(n1310) );
XOR2_X1 U1044 ( .A(KEYINPUT22), .B(G146), .Z(n1309) );
XOR2_X1 U1045 ( .A(n1311), .B(n1102), .Z(n1307) );
XOR2_X1 U1046 ( .A(G125), .B(G140), .Z(n1102) );
XOR2_X1 U1047 ( .A(n1126), .B(n1312), .Z(n1311) );
NOR2_X1 U1048 ( .A1(KEYINPUT13), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1049 ( .A(n1314), .B(n1315), .Z(n1313) );
XOR2_X1 U1050 ( .A(n1316), .B(n1317), .Z(n1315) );
AND3_X1 U1051 ( .A1(G214), .A2(n1057), .A3(n1265), .ZN(n1317) );
INV_X1 U1052 ( .A(G237), .ZN(n1265) );
NOR2_X1 U1053 ( .A1(KEYINPUT0), .A2(n1284), .ZN(n1316) );
INV_X1 U1054 ( .A(G131), .ZN(n1284) );
XOR2_X1 U1055 ( .A(KEYINPUT27), .B(G143), .Z(n1314) );
INV_X1 U1056 ( .A(G104), .ZN(n1126) );
XOR2_X1 U1057 ( .A(n1075), .B(G478), .Z(n1238) );
NAND2_X1 U1058 ( .A1(n1120), .A2(n1260), .ZN(n1075) );
INV_X1 U1059 ( .A(G902), .ZN(n1260) );
XOR2_X1 U1060 ( .A(n1318), .B(n1319), .Z(n1120) );
XOR2_X1 U1061 ( .A(G107), .B(n1320), .Z(n1319) );
XOR2_X1 U1062 ( .A(G122), .B(G116), .Z(n1320) );
XOR2_X1 U1063 ( .A(n1096), .B(n1321), .Z(n1318) );
XOR2_X1 U1064 ( .A(n1322), .B(n1323), .Z(n1321) );
NAND2_X1 U1065 ( .A1(G217), .A2(n1257), .ZN(n1323) );
AND2_X1 U1066 ( .A1(G234), .A2(n1057), .ZN(n1257) );
INV_X1 U1067 ( .A(G953), .ZN(n1057) );
NAND2_X1 U1068 ( .A1(KEYINPUT51), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1069 ( .A(G143), .B(G128), .Z(n1324) );
XNOR2_X1 U1070 ( .A(G134), .B(KEYINPUT58), .ZN(n1096) );
endmodule


