//Key = 0001000111110101011001110001000011100000100101110000101011110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339;

XOR2_X1 U748 ( .A(G107), .B(n1023), .Z(G9) );
NAND3_X1 U749 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(G75) );
INV_X1 U750 ( .A(n1027), .ZN(n1026) );
NAND2_X1 U751 ( .A1(n1028), .A2(n1029), .ZN(n1025) );
INV_X1 U752 ( .A(G952), .ZN(n1029) );
NAND2_X1 U753 ( .A1(G952), .A2(n1030), .ZN(n1024) );
NAND4_X1 U754 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1030) );
NOR4_X1 U755 ( .A1(G953), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1034) );
NOR2_X1 U756 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U757 ( .A1(n1040), .A2(n1041), .ZN(n1036) );
NOR3_X1 U758 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1040) );
NOR2_X1 U759 ( .A1(n1045), .A2(n1039), .ZN(n1044) );
NOR4_X1 U760 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1043) );
INV_X1 U761 ( .A(KEYINPUT16), .ZN(n1049) );
XOR2_X1 U762 ( .A(KEYINPUT14), .B(n1050), .Z(n1042) );
NOR3_X1 U763 ( .A1(n1051), .A2(n1039), .A3(n1052), .ZN(n1050) );
NOR2_X1 U764 ( .A1(n1053), .A2(n1054), .ZN(n1035) );
NOR2_X1 U765 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR3_X1 U766 ( .A1(n1057), .A2(n1039), .A3(n1058), .ZN(n1056) );
OR3_X1 U767 ( .A1(n1059), .A2(n1060), .A3(n1048), .ZN(n1039) );
NOR3_X1 U768 ( .A1(n1048), .A2(n1061), .A3(n1041), .ZN(n1055) );
NOR3_X1 U769 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NOR2_X1 U770 ( .A1(KEYINPUT16), .A2(n1047), .ZN(n1064) );
INV_X1 U771 ( .A(n1065), .ZN(n1047) );
NOR2_X1 U772 ( .A1(n1066), .A2(n1060), .ZN(n1063) );
INV_X1 U773 ( .A(n1067), .ZN(n1060) );
NOR2_X1 U774 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
AND2_X1 U775 ( .A1(n1070), .A2(n1071), .ZN(n1062) );
XNOR2_X1 U776 ( .A(n1028), .B(KEYINPUT0), .ZN(n1033) );
AND4_X1 U777 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1028) );
NOR4_X1 U778 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1054), .ZN(n1075) );
XOR2_X1 U779 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U780 ( .A1(G475), .A2(KEYINPUT49), .ZN(n1080) );
XOR2_X1 U781 ( .A(n1081), .B(KEYINPUT2), .Z(n1079) );
XOR2_X1 U782 ( .A(n1082), .B(n1083), .Z(n1077) );
XOR2_X1 U783 ( .A(KEYINPUT19), .B(n1084), .Z(n1083) );
NOR2_X1 U784 ( .A1(KEYINPUT36), .A2(n1085), .ZN(n1084) );
XNOR2_X1 U785 ( .A(n1086), .B(n1087), .ZN(n1074) );
NAND2_X1 U786 ( .A1(KEYINPUT52), .A2(n1088), .ZN(n1086) );
XNOR2_X1 U787 ( .A(n1058), .B(KEYINPUT1), .ZN(n1073) );
XOR2_X1 U788 ( .A(n1089), .B(n1090), .Z(n1072) );
NOR2_X1 U789 ( .A1(KEYINPUT51), .A2(n1091), .ZN(n1090) );
XOR2_X1 U790 ( .A(n1092), .B(n1093), .Z(G72) );
NOR2_X1 U791 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
AND2_X1 U792 ( .A1(G227), .A2(G900), .ZN(n1094) );
NAND2_X1 U793 ( .A1(n1096), .A2(n1097), .ZN(n1092) );
OR2_X1 U794 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NAND2_X1 U795 ( .A1(n1100), .A2(n1098), .ZN(n1096) );
NAND2_X1 U796 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U797 ( .A1(n1103), .A2(G953), .ZN(n1102) );
XOR2_X1 U798 ( .A(n1104), .B(n1105), .Z(n1101) );
XNOR2_X1 U799 ( .A(n1106), .B(n1107), .ZN(n1105) );
XNOR2_X1 U800 ( .A(n1108), .B(n1109), .ZN(n1104) );
NOR2_X1 U801 ( .A1(KEYINPUT61), .A2(n1110), .ZN(n1109) );
XOR2_X1 U802 ( .A(n1111), .B(KEYINPUT57), .Z(n1100) );
NAND2_X1 U803 ( .A1(n1095), .A2(n1099), .ZN(n1111) );
XOR2_X1 U804 ( .A(n1112), .B(n1113), .Z(G69) );
XOR2_X1 U805 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U806 ( .A1(G953), .A2(n1116), .ZN(n1115) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1116) );
NAND2_X1 U808 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NAND2_X1 U809 ( .A1(G953), .A2(n1119), .ZN(n1118) );
XOR2_X1 U810 ( .A(n1120), .B(n1121), .Z(n1117) );
XNOR2_X1 U811 ( .A(n1122), .B(n1123), .ZN(n1121) );
NAND2_X1 U812 ( .A1(KEYINPUT11), .A2(n1124), .ZN(n1122) );
NOR2_X1 U813 ( .A1(n1032), .A2(G953), .ZN(n1112) );
NOR2_X1 U814 ( .A1(n1027), .A2(n1125), .ZN(G66) );
XOR2_X1 U815 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U816 ( .A1(n1087), .A2(n1128), .ZN(n1127) );
NAND2_X1 U817 ( .A1(KEYINPUT21), .A2(n1129), .ZN(n1126) );
NOR2_X1 U818 ( .A1(n1027), .A2(n1130), .ZN(G63) );
XOR2_X1 U819 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U820 ( .A(n1133), .B(KEYINPUT55), .Z(n1131) );
NAND2_X1 U821 ( .A1(n1134), .A2(G478), .ZN(n1133) );
NOR2_X1 U822 ( .A1(n1027), .A2(n1135), .ZN(G60) );
XOR2_X1 U823 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U824 ( .A1(n1134), .A2(G475), .ZN(n1136) );
XOR2_X1 U825 ( .A(G104), .B(n1138), .Z(G6) );
NOR2_X1 U826 ( .A1(n1027), .A2(n1139), .ZN(G57) );
XOR2_X1 U827 ( .A(n1140), .B(n1141), .Z(n1139) );
XNOR2_X1 U828 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR3_X1 U829 ( .A1(n1128), .A2(KEYINPUT35), .A3(n1144), .ZN(n1143) );
NAND2_X1 U830 ( .A1(n1145), .A2(KEYINPUT59), .ZN(n1142) );
XOR2_X1 U831 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U832 ( .A1(G101), .A2(KEYINPUT48), .ZN(n1147) );
XOR2_X1 U833 ( .A(n1148), .B(n1149), .Z(n1140) );
NOR2_X1 U834 ( .A1(n1027), .A2(n1150), .ZN(G54) );
XOR2_X1 U835 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U836 ( .A(n1153), .B(n1154), .Z(n1152) );
XOR2_X1 U837 ( .A(n1155), .B(KEYINPUT39), .Z(n1154) );
NAND2_X1 U838 ( .A1(n1134), .A2(G469), .ZN(n1155) );
NAND2_X1 U839 ( .A1(KEYINPUT54), .A2(n1106), .ZN(n1153) );
XNOR2_X1 U840 ( .A(n1156), .B(n1157), .ZN(n1151) );
NOR2_X1 U841 ( .A1(n1027), .A2(n1158), .ZN(G51) );
XOR2_X1 U842 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U843 ( .A(n1161), .B(KEYINPUT22), .Z(n1160) );
NAND2_X1 U844 ( .A1(n1134), .A2(n1162), .ZN(n1161) );
INV_X1 U845 ( .A(n1128), .ZN(n1134) );
NAND2_X1 U846 ( .A1(G902), .A2(n1163), .ZN(n1128) );
NAND2_X1 U847 ( .A1(n1031), .A2(n1032), .ZN(n1163) );
AND4_X1 U848 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1032) );
NOR4_X1 U849 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NOR4_X1 U850 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1038), .ZN(n1171) );
XNOR2_X1 U851 ( .A(n1175), .B(KEYINPUT15), .ZN(n1172) );
NOR2_X1 U852 ( .A1(n1138), .A2(n1023), .ZN(n1166) );
AND3_X1 U853 ( .A1(n1068), .A2(n1176), .A3(n1067), .ZN(n1023) );
AND3_X1 U854 ( .A1(n1067), .A2(n1176), .A3(n1069), .ZN(n1138) );
INV_X1 U855 ( .A(n1177), .ZN(n1165) );
INV_X1 U856 ( .A(n1099), .ZN(n1031) );
NAND4_X1 U857 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1099) );
NOR3_X1 U858 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1181) );
NOR2_X1 U859 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NOR2_X1 U860 ( .A1(n1187), .A2(n1188), .ZN(n1185) );
NOR2_X1 U861 ( .A1(n1045), .A2(n1041), .ZN(n1187) );
NOR2_X1 U862 ( .A1(n1189), .A2(n1190), .ZN(n1183) );
NOR2_X1 U863 ( .A1(n1191), .A2(n1192), .ZN(n1189) );
NOR2_X1 U864 ( .A1(n1193), .A2(n1174), .ZN(n1192) );
NOR2_X1 U865 ( .A1(n1194), .A2(n1195), .ZN(n1191) );
XNOR2_X1 U866 ( .A(n1193), .B(KEYINPUT3), .ZN(n1195) );
INV_X1 U867 ( .A(n1068), .ZN(n1194) );
NOR2_X1 U868 ( .A1(n1041), .A2(n1196), .ZN(n1182) );
NOR2_X1 U869 ( .A1(n1095), .A2(G952), .ZN(n1027) );
XOR2_X1 U870 ( .A(G146), .B(n1197), .Z(G48) );
NOR4_X1 U871 ( .A1(KEYINPUT42), .A2(n1193), .A3(n1190), .A4(n1174), .ZN(n1197) );
INV_X1 U872 ( .A(n1069), .ZN(n1174) );
NAND3_X1 U873 ( .A1(n1198), .A2(n1199), .A3(n1200), .ZN(G45) );
OR2_X1 U874 ( .A1(n1201), .A2(KEYINPUT62), .ZN(n1200) );
NAND3_X1 U875 ( .A1(KEYINPUT62), .A2(n1201), .A3(n1202), .ZN(n1199) );
NAND2_X1 U876 ( .A1(G143), .A2(n1203), .ZN(n1198) );
NAND2_X1 U877 ( .A1(KEYINPUT62), .A2(n1204), .ZN(n1203) );
XNOR2_X1 U878 ( .A(KEYINPUT24), .B(n1179), .ZN(n1204) );
INV_X1 U879 ( .A(n1201), .ZN(n1179) );
NOR4_X1 U880 ( .A1(n1190), .A2(n1173), .A3(n1205), .A4(n1206), .ZN(n1201) );
XOR2_X1 U881 ( .A(G140), .B(n1207), .Z(G42) );
NOR3_X1 U882 ( .A1(n1186), .A2(n1208), .A3(n1041), .ZN(n1207) );
XNOR2_X1 U883 ( .A(n1209), .B(KEYINPUT20), .ZN(n1208) );
XNOR2_X1 U884 ( .A(G137), .B(n1210), .ZN(G39) );
NAND2_X1 U885 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NAND2_X1 U886 ( .A1(KEYINPUT8), .A2(n1180), .ZN(n1212) );
NAND2_X1 U887 ( .A1(KEYINPUT60), .A2(n1213), .ZN(n1211) );
INV_X1 U888 ( .A(n1180), .ZN(n1213) );
NAND4_X1 U889 ( .A1(n1071), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1180) );
XOR2_X1 U890 ( .A(n1217), .B(n1218), .Z(G36) );
NOR2_X1 U891 ( .A1(KEYINPUT29), .A2(n1219), .ZN(n1218) );
NOR2_X1 U892 ( .A1(n1041), .A2(n1220), .ZN(n1217) );
XNOR2_X1 U893 ( .A(KEYINPUT58), .B(n1196), .ZN(n1220) );
NAND3_X1 U894 ( .A1(n1215), .A2(n1068), .A3(n1221), .ZN(n1196) );
INV_X1 U895 ( .A(n1214), .ZN(n1041) );
XNOR2_X1 U896 ( .A(G131), .B(n1178), .ZN(G33) );
NAND4_X1 U897 ( .A1(n1069), .A2(n1214), .A3(n1221), .A4(n1215), .ZN(n1178) );
NOR2_X1 U898 ( .A1(n1058), .A2(n1076), .ZN(n1214) );
XNOR2_X1 U899 ( .A(G128), .B(n1222), .ZN(G30) );
NAND3_X1 U900 ( .A1(n1223), .A2(n1068), .A3(n1224), .ZN(n1222) );
XNOR2_X1 U901 ( .A(KEYINPUT46), .B(n1216), .ZN(n1224) );
INV_X1 U902 ( .A(n1190), .ZN(n1223) );
NAND2_X1 U903 ( .A1(n1215), .A2(n1225), .ZN(n1190) );
AND2_X1 U904 ( .A1(n1209), .A2(n1226), .ZN(n1215) );
XNOR2_X1 U905 ( .A(G101), .B(n1164), .ZN(G3) );
NAND2_X1 U906 ( .A1(n1065), .A2(n1176), .ZN(n1164) );
NOR2_X1 U907 ( .A1(n1059), .A2(n1173), .ZN(n1065) );
XOR2_X1 U908 ( .A(G125), .B(n1227), .Z(G27) );
NOR2_X1 U909 ( .A1(n1186), .A2(n1038), .ZN(n1227) );
NAND3_X1 U910 ( .A1(n1070), .A2(n1226), .A3(n1069), .ZN(n1186) );
NAND2_X1 U911 ( .A1(n1048), .A2(n1228), .ZN(n1226) );
NAND4_X1 U912 ( .A1(n1103), .A2(G953), .A3(G902), .A4(n1229), .ZN(n1228) );
XNOR2_X1 U913 ( .A(G900), .B(KEYINPUT53), .ZN(n1103) );
XOR2_X1 U914 ( .A(G122), .B(n1170), .Z(G24) );
AND3_X1 U915 ( .A1(n1188), .A2(n1067), .A3(n1230), .ZN(n1170) );
NOR3_X1 U916 ( .A1(n1205), .A2(n1175), .A3(n1206), .ZN(n1230) );
INV_X1 U917 ( .A(n1038), .ZN(n1188) );
XNOR2_X1 U918 ( .A(G119), .B(n1231), .ZN(G21) );
NAND2_X1 U919 ( .A1(KEYINPUT43), .A2(n1177), .ZN(n1231) );
NOR4_X1 U920 ( .A1(n1038), .A2(n1059), .A3(n1193), .A4(n1175), .ZN(n1177) );
INV_X1 U921 ( .A(n1216), .ZN(n1193) );
NAND2_X1 U922 ( .A1(n1232), .A2(n1233), .ZN(n1216) );
NAND2_X1 U923 ( .A1(n1221), .A2(n1234), .ZN(n1233) );
NAND3_X1 U924 ( .A1(n1235), .A2(n1236), .A3(KEYINPUT32), .ZN(n1232) );
INV_X1 U925 ( .A(n1071), .ZN(n1059) );
XOR2_X1 U926 ( .A(G116), .B(n1169), .Z(G18) );
AND2_X1 U927 ( .A1(n1237), .A2(n1068), .ZN(n1169) );
NOR2_X1 U928 ( .A1(n1238), .A2(n1206), .ZN(n1068) );
INV_X1 U929 ( .A(n1239), .ZN(n1206) );
XOR2_X1 U930 ( .A(n1240), .B(n1241), .Z(G15) );
NAND2_X1 U931 ( .A1(n1237), .A2(n1069), .ZN(n1241) );
NOR2_X1 U932 ( .A1(n1239), .A2(n1205), .ZN(n1069) );
INV_X1 U933 ( .A(n1238), .ZN(n1205) );
NOR3_X1 U934 ( .A1(n1173), .A2(n1175), .A3(n1038), .ZN(n1237) );
NAND2_X1 U935 ( .A1(n1046), .A2(n1225), .ZN(n1038) );
INV_X1 U936 ( .A(n1054), .ZN(n1046) );
NAND2_X1 U937 ( .A1(n1242), .A2(n1051), .ZN(n1054) );
INV_X1 U938 ( .A(n1052), .ZN(n1242) );
INV_X1 U939 ( .A(n1243), .ZN(n1175) );
INV_X1 U940 ( .A(n1221), .ZN(n1173) );
NOR2_X1 U941 ( .A1(n1235), .A2(n1244), .ZN(n1221) );
NAND2_X1 U942 ( .A1(KEYINPUT40), .A2(G113), .ZN(n1240) );
XOR2_X1 U943 ( .A(G110), .B(n1168), .Z(G12) );
AND3_X1 U944 ( .A1(n1176), .A2(n1070), .A3(n1071), .ZN(n1168) );
NOR2_X1 U945 ( .A1(n1239), .A2(n1238), .ZN(n1071) );
XNOR2_X1 U946 ( .A(n1081), .B(G475), .ZN(n1238) );
NAND2_X1 U947 ( .A1(n1245), .A2(n1246), .ZN(n1081) );
XOR2_X1 U948 ( .A(n1137), .B(KEYINPUT12), .Z(n1245) );
XOR2_X1 U949 ( .A(n1247), .B(n1248), .Z(n1137) );
XOR2_X1 U950 ( .A(n1249), .B(n1250), .Z(n1248) );
XOR2_X1 U951 ( .A(G104), .B(n1251), .Z(n1250) );
NOR2_X1 U952 ( .A1(KEYINPUT50), .A2(n1107), .ZN(n1251) );
XOR2_X1 U953 ( .A(G125), .B(n1252), .Z(n1107) );
XNOR2_X1 U954 ( .A(n1108), .B(G122), .ZN(n1249) );
INV_X1 U955 ( .A(G131), .ZN(n1108) );
XNOR2_X1 U956 ( .A(n1253), .B(n1254), .ZN(n1247) );
XOR2_X1 U957 ( .A(n1255), .B(n1256), .Z(n1254) );
NAND2_X1 U958 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U959 ( .A1(G214), .A2(n1259), .ZN(n1255) );
XOR2_X1 U960 ( .A(n1089), .B(n1091), .Z(n1239) );
INV_X1 U961 ( .A(G478), .ZN(n1091) );
NAND2_X1 U962 ( .A1(n1132), .A2(n1246), .ZN(n1089) );
XNOR2_X1 U963 ( .A(n1260), .B(n1261), .ZN(n1132) );
XOR2_X1 U964 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U965 ( .A(G122), .B(G116), .Z(n1263) );
XNOR2_X1 U966 ( .A(KEYINPUT30), .B(n1219), .ZN(n1262) );
XOR2_X1 U967 ( .A(n1264), .B(n1265), .Z(n1260) );
AND3_X1 U968 ( .A1(G217), .A2(n1095), .A3(G234), .ZN(n1265) );
XOR2_X1 U969 ( .A(n1266), .B(G107), .Z(n1264) );
NAND2_X1 U970 ( .A1(KEYINPUT10), .A2(n1267), .ZN(n1266) );
INV_X1 U971 ( .A(n1268), .ZN(n1267) );
NAND2_X1 U972 ( .A1(n1269), .A2(n1270), .ZN(n1070) );
NAND2_X1 U973 ( .A1(n1067), .A2(n1234), .ZN(n1270) );
INV_X1 U974 ( .A(KEYINPUT32), .ZN(n1234) );
NOR2_X1 U975 ( .A1(n1236), .A2(n1235), .ZN(n1067) );
NAND3_X1 U976 ( .A1(n1235), .A2(n1244), .A3(KEYINPUT32), .ZN(n1269) );
INV_X1 U977 ( .A(n1236), .ZN(n1244) );
XNOR2_X1 U978 ( .A(n1082), .B(n1085), .ZN(n1236) );
XNOR2_X1 U979 ( .A(n1144), .B(KEYINPUT44), .ZN(n1085) );
INV_X1 U980 ( .A(G472), .ZN(n1144) );
NAND2_X1 U981 ( .A1(n1271), .A2(n1246), .ZN(n1082) );
XOR2_X1 U982 ( .A(n1272), .B(n1273), .Z(n1271) );
XNOR2_X1 U983 ( .A(n1274), .B(KEYINPUT33), .ZN(n1273) );
NAND2_X1 U984 ( .A1(n1275), .A2(KEYINPUT9), .ZN(n1274) );
XOR2_X1 U985 ( .A(n1146), .B(n1276), .Z(n1275) );
XOR2_X1 U986 ( .A(KEYINPUT28), .B(G101), .Z(n1276) );
NAND2_X1 U987 ( .A1(G210), .A2(n1259), .ZN(n1146) );
NOR2_X1 U988 ( .A1(G953), .A2(G237), .ZN(n1259) );
XOR2_X1 U989 ( .A(n1277), .B(n1149), .Z(n1272) );
XNOR2_X1 U990 ( .A(n1278), .B(G119), .ZN(n1149) );
NAND2_X1 U991 ( .A1(KEYINPUT23), .A2(n1148), .ZN(n1277) );
XNOR2_X1 U992 ( .A(n1279), .B(n1280), .ZN(n1148) );
XNOR2_X1 U993 ( .A(n1088), .B(n1087), .ZN(n1235) );
NAND2_X1 U994 ( .A1(G217), .A2(n1281), .ZN(n1087) );
AND2_X1 U995 ( .A1(n1129), .A2(n1246), .ZN(n1088) );
XOR2_X1 U996 ( .A(n1282), .B(n1283), .Z(n1129) );
XNOR2_X1 U997 ( .A(n1284), .B(n1285), .ZN(n1283) );
NOR2_X1 U998 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U999 ( .A(n1288), .B(KEYINPUT17), .Z(n1287) );
NAND2_X1 U1000 ( .A1(n1289), .A2(G137), .ZN(n1288) );
NOR2_X1 U1001 ( .A1(G137), .A2(n1289), .ZN(n1286) );
AND3_X1 U1002 ( .A1(G221), .A2(n1095), .A3(G234), .ZN(n1289) );
XNOR2_X1 U1003 ( .A(n1290), .B(n1291), .ZN(n1284) );
NOR2_X1 U1004 ( .A1(KEYINPUT38), .A2(G110), .ZN(n1291) );
NOR2_X1 U1005 ( .A1(KEYINPUT4), .A2(n1292), .ZN(n1290) );
XOR2_X1 U1006 ( .A(n1293), .B(n1294), .Z(n1292) );
NOR2_X1 U1007 ( .A1(KEYINPUT25), .A2(n1252), .ZN(n1294) );
XNOR2_X1 U1008 ( .A(G125), .B(KEYINPUT45), .ZN(n1293) );
XNOR2_X1 U1009 ( .A(n1295), .B(n1296), .ZN(n1282) );
XOR2_X1 U1010 ( .A(G146), .B(G128), .Z(n1296) );
AND3_X1 U1011 ( .A1(n1225), .A2(n1243), .A3(n1209), .ZN(n1176) );
INV_X1 U1012 ( .A(n1045), .ZN(n1209) );
NAND2_X1 U1013 ( .A1(n1052), .A2(n1051), .ZN(n1045) );
NAND2_X1 U1014 ( .A1(G221), .A2(n1281), .ZN(n1051) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1246), .ZN(n1281) );
XNOR2_X1 U1016 ( .A(n1297), .B(G469), .ZN(n1052) );
NAND2_X1 U1017 ( .A1(n1298), .A2(n1246), .ZN(n1297) );
XOR2_X1 U1018 ( .A(n1299), .B(n1156), .Z(n1298) );
XOR2_X1 U1019 ( .A(n1300), .B(n1301), .Z(n1156) );
XOR2_X1 U1020 ( .A(G110), .B(n1302), .Z(n1301) );
AND2_X1 U1021 ( .A1(n1095), .A2(G227), .ZN(n1302) );
XNOR2_X1 U1022 ( .A(n1279), .B(n1252), .ZN(n1300) );
XNOR2_X1 U1023 ( .A(G140), .B(KEYINPUT26), .ZN(n1252) );
XNOR2_X1 U1024 ( .A(G131), .B(n1303), .ZN(n1279) );
NOR2_X1 U1025 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NOR3_X1 U1026 ( .A1(KEYINPUT18), .A2(G137), .A3(n1219), .ZN(n1305) );
NOR2_X1 U1027 ( .A1(n1110), .A2(n1306), .ZN(n1304) );
INV_X1 U1028 ( .A(KEYINPUT18), .ZN(n1306) );
XNOR2_X1 U1029 ( .A(n1219), .B(G137), .ZN(n1110) );
INV_X1 U1030 ( .A(G134), .ZN(n1219) );
NAND3_X1 U1031 ( .A1(n1307), .A2(n1308), .A3(n1309), .ZN(n1299) );
OR2_X1 U1032 ( .A1(n1106), .A2(KEYINPUT56), .ZN(n1309) );
NAND3_X1 U1033 ( .A1(KEYINPUT56), .A2(n1106), .A3(n1123), .ZN(n1308) );
NAND2_X1 U1034 ( .A1(n1157), .A2(n1310), .ZN(n1307) );
NAND2_X1 U1035 ( .A1(n1311), .A2(KEYINPUT56), .ZN(n1310) );
XNOR2_X1 U1036 ( .A(KEYINPUT63), .B(n1312), .ZN(n1311) );
INV_X1 U1037 ( .A(n1106), .ZN(n1312) );
XOR2_X1 U1038 ( .A(G128), .B(n1313), .Z(n1106) );
NOR2_X1 U1039 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
NOR2_X1 U1040 ( .A1(KEYINPUT34), .A2(n1316), .ZN(n1315) );
AND2_X1 U1041 ( .A1(KEYINPUT47), .A2(n1316), .ZN(n1314) );
AND2_X1 U1042 ( .A1(n1317), .A2(n1257), .ZN(n1316) );
XOR2_X1 U1043 ( .A(n1258), .B(KEYINPUT31), .Z(n1317) );
OR2_X1 U1044 ( .A1(n1202), .A2(G146), .ZN(n1258) );
NAND2_X1 U1045 ( .A1(n1048), .A2(n1318), .ZN(n1243) );
NAND4_X1 U1046 ( .A1(G953), .A2(G902), .A3(n1229), .A4(n1119), .ZN(n1318) );
INV_X1 U1047 ( .A(G898), .ZN(n1119) );
NAND3_X1 U1048 ( .A1(n1229), .A2(n1095), .A3(G952), .ZN(n1048) );
NAND2_X1 U1049 ( .A1(G237), .A2(G234), .ZN(n1229) );
NOR2_X1 U1050 ( .A1(n1319), .A2(n1076), .ZN(n1225) );
INV_X1 U1051 ( .A(n1057), .ZN(n1076) );
NAND2_X1 U1052 ( .A1(n1320), .A2(n1321), .ZN(n1057) );
XOR2_X1 U1053 ( .A(KEYINPUT37), .B(G214), .Z(n1320) );
INV_X1 U1054 ( .A(n1058), .ZN(n1319) );
XNOR2_X1 U1055 ( .A(n1322), .B(n1162), .ZN(n1058) );
AND2_X1 U1056 ( .A1(G210), .A2(n1321), .ZN(n1162) );
NAND2_X1 U1057 ( .A1(n1323), .A2(n1246), .ZN(n1321) );
INV_X1 U1058 ( .A(G237), .ZN(n1323) );
NAND2_X1 U1059 ( .A1(n1324), .A2(n1246), .ZN(n1322) );
INV_X1 U1060 ( .A(G902), .ZN(n1246) );
XOR2_X1 U1061 ( .A(n1159), .B(KEYINPUT7), .Z(n1324) );
XOR2_X1 U1062 ( .A(n1325), .B(n1326), .Z(n1159) );
XOR2_X1 U1063 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1064 ( .A(G125), .B(n1280), .ZN(n1328) );
NAND3_X1 U1065 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1280) );
NAND2_X1 U1066 ( .A1(n1332), .A2(n1268), .ZN(n1331) );
XOR2_X1 U1067 ( .A(G128), .B(n1202), .Z(n1268) );
OR3_X1 U1068 ( .A1(n1202), .A2(n1332), .A3(G128), .ZN(n1330) );
NOR2_X1 U1069 ( .A1(KEYINPUT41), .A2(G146), .ZN(n1332) );
NAND2_X1 U1070 ( .A1(G128), .A2(n1333), .ZN(n1329) );
NAND2_X1 U1071 ( .A1(n1257), .A2(n1334), .ZN(n1333) );
NAND2_X1 U1072 ( .A1(KEYINPUT41), .A2(n1202), .ZN(n1334) );
NAND2_X1 U1073 ( .A1(G146), .A2(n1202), .ZN(n1257) );
INV_X1 U1074 ( .A(G143), .ZN(n1202) );
NOR2_X1 U1075 ( .A1(KEYINPUT6), .A2(n1157), .ZN(n1327) );
INV_X1 U1076 ( .A(n1123), .ZN(n1157) );
XOR2_X1 U1077 ( .A(G101), .B(n1335), .Z(n1123) );
XOR2_X1 U1078 ( .A(G107), .B(G104), .Z(n1335) );
XOR2_X1 U1079 ( .A(n1336), .B(n1124), .Z(n1325) );
XOR2_X1 U1080 ( .A(G110), .B(n1337), .Z(n1124) );
XOR2_X1 U1081 ( .A(KEYINPUT27), .B(G122), .Z(n1337) );
XOR2_X1 U1082 ( .A(n1120), .B(n1338), .Z(n1336) );
AND2_X1 U1083 ( .A1(n1095), .A2(G224), .ZN(n1338) );
INV_X1 U1084 ( .A(G953), .ZN(n1095) );
XNOR2_X1 U1085 ( .A(n1339), .B(n1278), .ZN(n1120) );
XNOR2_X1 U1086 ( .A(G116), .B(n1253), .ZN(n1278) );
XOR2_X1 U1087 ( .A(G113), .B(KEYINPUT5), .Z(n1253) );
NAND2_X1 U1088 ( .A1(KEYINPUT13), .A2(n1295), .ZN(n1339) );
INV_X1 U1089 ( .A(G119), .ZN(n1295) );
endmodule


