//Key = 0110111111101110011000101110100000110010001100100010000011111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;

XNOR2_X1 U738 ( .A(G107), .B(n1018), .ZN(G9) );
NAND3_X1 U739 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NOR2_X1 U740 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U741 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
NOR4_X1 U742 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1026) );
NOR2_X1 U743 ( .A1(n1032), .A2(n1033), .ZN(n1029) );
NAND4_X1 U744 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1033) );
NAND2_X1 U745 ( .A1(n1021), .A2(n1020), .ZN(n1037) );
NAND2_X1 U746 ( .A1(KEYINPUT7), .A2(n1038), .ZN(n1036) );
NAND2_X1 U747 ( .A1(n1039), .A2(n1040), .ZN(n1035) );
NAND2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1034) );
NOR3_X1 U749 ( .A1(n1043), .A2(n1044), .A3(n1045), .ZN(n1028) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1042), .ZN(n1045) );
INV_X1 U751 ( .A(KEYINPUT52), .ZN(n1042) );
NOR2_X1 U752 ( .A1(KEYINPUT7), .A2(n1047), .ZN(n1044) );
NAND3_X1 U753 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1024) );
NAND4_X1 U754 ( .A1(n1043), .A2(n1039), .A3(n1021), .A4(n1051), .ZN(n1050) );
NAND3_X1 U755 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1051) );
NAND2_X1 U756 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U757 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U758 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
XOR2_X1 U759 ( .A(n1061), .B(KEYINPUT12), .Z(n1059) );
INV_X1 U760 ( .A(n1062), .ZN(n1053) );
NAND3_X1 U761 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1052) );
INV_X1 U762 ( .A(n1032), .ZN(n1043) );
NOR3_X1 U763 ( .A1(n1066), .A2(G953), .A3(G952), .ZN(n1022) );
INV_X1 U764 ( .A(n1048), .ZN(n1066) );
NAND4_X1 U765 ( .A1(n1067), .A2(n1061), .A3(n1068), .A4(n1069), .ZN(n1048) );
NOR4_X1 U766 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
XOR2_X1 U767 ( .A(n1074), .B(n1075), .Z(n1073) );
XNOR2_X1 U768 ( .A(KEYINPUT8), .B(n1076), .ZN(n1075) );
XOR2_X1 U769 ( .A(n1077), .B(KEYINPUT49), .Z(n1072) );
NAND2_X1 U770 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
INV_X1 U771 ( .A(n1080), .ZN(n1078) );
XNOR2_X1 U772 ( .A(n1081), .B(KEYINPUT61), .ZN(n1071) );
NAND3_X1 U773 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1070) );
NAND3_X1 U774 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1083) );
INV_X1 U775 ( .A(KEYINPUT39), .ZN(n1087) );
NAND2_X1 U776 ( .A1(KEYINPUT39), .A2(n1088), .ZN(n1082) );
NOR3_X1 U777 ( .A1(n1089), .A2(n1065), .A3(n1090), .ZN(n1068) );
XOR2_X1 U778 ( .A(KEYINPUT62), .B(n1091), .Z(n1067) );
NOR2_X1 U779 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U780 ( .A(G475), .B(KEYINPUT51), .ZN(n1093) );
NOR2_X1 U781 ( .A1(G902), .A2(n1094), .ZN(n1092) );
XOR2_X1 U782 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U783 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U784 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
INV_X1 U785 ( .A(n1101), .ZN(n1100) );
XOR2_X1 U786 ( .A(n1102), .B(n1103), .Z(n1099) );
XOR2_X1 U787 ( .A(n1104), .B(n1105), .Z(n1103) );
NAND2_X1 U788 ( .A1(n1106), .A2(KEYINPUT46), .ZN(n1104) );
XNOR2_X1 U789 ( .A(G134), .B(G137), .ZN(n1106) );
NAND2_X1 U790 ( .A1(n1107), .A2(n1049), .ZN(n1097) );
XNOR2_X1 U791 ( .A(KEYINPUT5), .B(n1027), .ZN(n1107) );
NOR2_X1 U792 ( .A1(n1108), .A2(n1049), .ZN(n1095) );
AND2_X1 U793 ( .A1(G227), .A2(G900), .ZN(n1108) );
XOR2_X1 U794 ( .A(n1109), .B(n1110), .Z(G69) );
XOR2_X1 U795 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U796 ( .A1(n1113), .A2(n1049), .ZN(n1112) );
AND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1113) );
NAND2_X1 U798 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
OR2_X1 U799 ( .A1(n1049), .A2(G898), .ZN(n1115) );
XOR2_X1 U800 ( .A(n1116), .B(n1117), .Z(n1114) );
NAND2_X1 U801 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NAND2_X1 U802 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U803 ( .A(n1122), .B(KEYINPUT29), .Z(n1120) );
NAND2_X1 U804 ( .A1(n1123), .A2(n1124), .ZN(n1118) );
XOR2_X1 U805 ( .A(n1122), .B(KEYINPUT14), .Z(n1124) );
NAND2_X1 U806 ( .A1(n1049), .A2(n1025), .ZN(n1109) );
NOR2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(G66) );
XOR2_X1 U808 ( .A(n1127), .B(n1128), .Z(n1126) );
NAND2_X1 U809 ( .A1(n1129), .A2(n1130), .ZN(n1127) );
NOR2_X1 U810 ( .A1(n1125), .A2(n1131), .ZN(G63) );
XOR2_X1 U811 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U812 ( .A1(n1129), .A2(G478), .ZN(n1132) );
NOR2_X1 U813 ( .A1(n1125), .A2(n1134), .ZN(G60) );
XNOR2_X1 U814 ( .A(n1135), .B(n1094), .ZN(n1134) );
NAND2_X1 U815 ( .A1(n1129), .A2(G475), .ZN(n1135) );
XNOR2_X1 U816 ( .A(G104), .B(n1136), .ZN(G6) );
NAND3_X1 U817 ( .A1(n1038), .A2(n1019), .A3(KEYINPUT25), .ZN(n1136) );
INV_X1 U818 ( .A(n1047), .ZN(n1038) );
NOR2_X1 U819 ( .A1(n1125), .A2(n1137), .ZN(G57) );
XOR2_X1 U820 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U822 ( .A1(KEYINPUT58), .A2(n1142), .ZN(n1140) );
XOR2_X1 U823 ( .A(n1143), .B(n1144), .Z(n1138) );
NOR2_X1 U824 ( .A1(KEYINPUT30), .A2(n1145), .ZN(n1144) );
NAND2_X1 U825 ( .A1(n1129), .A2(G472), .ZN(n1143) );
NOR3_X1 U826 ( .A1(n1146), .A2(n1147), .A3(n1148), .ZN(G54) );
NOR3_X1 U827 ( .A1(n1149), .A2(G953), .A3(G952), .ZN(n1148) );
AND2_X1 U828 ( .A1(n1149), .A2(n1125), .ZN(n1147) );
INV_X1 U829 ( .A(KEYINPUT54), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1146) );
NAND2_X1 U831 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
NAND2_X1 U832 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U833 ( .A(n1156), .B(KEYINPUT53), .Z(n1152) );
OR2_X1 U834 ( .A1(n1155), .A2(n1154), .ZN(n1156) );
NOR2_X1 U835 ( .A1(n1157), .A2(n1158), .ZN(n1154) );
XNOR2_X1 U836 ( .A(n1159), .B(KEYINPUT31), .ZN(n1157) );
NAND2_X1 U837 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U838 ( .A(n1162), .B(n1163), .Z(n1155) );
XOR2_X1 U839 ( .A(KEYINPUT37), .B(KEYINPUT32), .Z(n1163) );
XNOR2_X1 U840 ( .A(n1164), .B(n1121), .ZN(n1162) );
NAND2_X1 U841 ( .A1(n1129), .A2(G469), .ZN(n1150) );
NOR2_X1 U842 ( .A1(n1125), .A2(n1165), .ZN(G51) );
XOR2_X1 U843 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND4_X1 U844 ( .A1(KEYINPUT43), .A2(KEYINPUT26), .A3(n1129), .A4(G210), .ZN(n1167) );
AND2_X1 U845 ( .A1(G902), .A2(n1168), .ZN(n1129) );
OR2_X1 U846 ( .A1(n1025), .A2(n1027), .ZN(n1168) );
NAND4_X1 U847 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1027) );
AND4_X1 U848 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172) );
NOR2_X1 U849 ( .A1(n1177), .A2(n1178), .ZN(n1171) );
NOR2_X1 U850 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
NOR2_X1 U851 ( .A1(n1031), .A2(n1181), .ZN(n1177) );
NAND2_X1 U852 ( .A1(n1182), .A2(n1183), .ZN(n1169) );
NAND2_X1 U853 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
NAND4_X1 U854 ( .A1(n1186), .A2(n1020), .A3(n1187), .A4(n1180), .ZN(n1185) );
INV_X1 U855 ( .A(KEYINPUT59), .ZN(n1180) );
NAND4_X1 U856 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1025) );
NOR4_X1 U857 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
INV_X1 U858 ( .A(n1196), .ZN(n1194) );
OR2_X1 U859 ( .A1(n1197), .A2(n1198), .ZN(n1190) );
NAND3_X1 U860 ( .A1(n1199), .A2(n1200), .A3(n1020), .ZN(n1189) );
NAND2_X1 U861 ( .A1(n1201), .A2(n1202), .ZN(n1199) );
NAND4_X1 U862 ( .A1(n1203), .A2(KEYINPUT41), .A3(n1021), .A4(n1204), .ZN(n1202) );
NAND4_X1 U863 ( .A1(n1040), .A2(n1205), .A3(n1030), .A4(n1197), .ZN(n1201) );
INV_X1 U864 ( .A(KEYINPUT38), .ZN(n1197) );
NAND2_X1 U865 ( .A1(n1019), .A2(n1206), .ZN(n1188) );
NAND3_X1 U866 ( .A1(n1047), .A2(n1046), .A3(n1207), .ZN(n1206) );
NAND3_X1 U867 ( .A1(n1020), .A2(n1208), .A3(n1021), .ZN(n1207) );
INV_X1 U868 ( .A(KEYINPUT41), .ZN(n1208) );
NAND2_X1 U869 ( .A1(n1209), .A2(n1021), .ZN(n1047) );
NAND2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(n1166) );
OR2_X1 U871 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XOR2_X1 U872 ( .A(n1214), .B(KEYINPUT19), .Z(n1210) );
NAND2_X1 U873 ( .A1(n1213), .A2(n1212), .ZN(n1214) );
XOR2_X1 U874 ( .A(n1215), .B(KEYINPUT20), .Z(n1212) );
NOR2_X1 U875 ( .A1(n1049), .A2(G952), .ZN(n1125) );
XOR2_X1 U876 ( .A(n1175), .B(n1216), .Z(G48) );
NAND2_X1 U877 ( .A1(KEYINPUT6), .A2(G146), .ZN(n1216) );
NAND2_X1 U878 ( .A1(n1217), .A2(n1186), .ZN(n1175) );
XNOR2_X1 U879 ( .A(n1218), .B(n1219), .ZN(G45) );
NOR2_X1 U880 ( .A1(n1220), .A2(n1184), .ZN(n1219) );
NAND4_X1 U881 ( .A1(n1221), .A2(n1040), .A3(n1222), .A4(n1223), .ZN(n1184) );
INV_X1 U882 ( .A(n1224), .ZN(n1223) );
NOR2_X1 U883 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
XNOR2_X1 U884 ( .A(n1227), .B(KEYINPUT60), .ZN(n1220) );
XOR2_X1 U885 ( .A(n1170), .B(n1228), .Z(G42) );
XOR2_X1 U886 ( .A(KEYINPUT2), .B(G140), .Z(n1228) );
NAND4_X1 U887 ( .A1(n1055), .A2(n1217), .A3(n1229), .A4(n1230), .ZN(n1170) );
XNOR2_X1 U888 ( .A(n1231), .B(n1232), .ZN(G39) );
NOR3_X1 U889 ( .A1(n1233), .A2(KEYINPUT33), .A3(n1031), .ZN(n1232) );
XNOR2_X1 U890 ( .A(KEYINPUT17), .B(n1181), .ZN(n1233) );
NAND3_X1 U891 ( .A1(n1221), .A2(n1039), .A3(n1234), .ZN(n1181) );
NOR3_X1 U892 ( .A1(n1229), .A2(n1235), .A3(n1227), .ZN(n1234) );
XNOR2_X1 U893 ( .A(G134), .B(n1176), .ZN(G36) );
NAND4_X1 U894 ( .A1(n1221), .A2(n1055), .A3(n1236), .A4(n1040), .ZN(n1176) );
AND2_X1 U895 ( .A1(n1183), .A2(n1020), .ZN(n1236) );
XNOR2_X1 U896 ( .A(G131), .B(n1237), .ZN(G33) );
NAND2_X1 U897 ( .A1(KEYINPUT4), .A2(n1238), .ZN(n1237) );
INV_X1 U898 ( .A(n1174), .ZN(n1238) );
NAND3_X1 U899 ( .A1(n1217), .A2(n1040), .A3(n1055), .ZN(n1174) );
INV_X1 U900 ( .A(n1031), .ZN(n1055) );
NAND2_X1 U901 ( .A1(n1063), .A2(n1239), .ZN(n1031) );
AND3_X1 U902 ( .A1(n1209), .A2(n1183), .A3(n1221), .ZN(n1217) );
INV_X1 U903 ( .A(n1057), .ZN(n1221) );
XOR2_X1 U904 ( .A(n1204), .B(KEYINPUT13), .Z(n1057) );
XNOR2_X1 U905 ( .A(G128), .B(n1179), .ZN(G30) );
NAND4_X1 U906 ( .A1(n1186), .A2(n1020), .A3(n1204), .A4(n1183), .ZN(n1179) );
XNOR2_X1 U907 ( .A(G101), .B(n1196), .ZN(G3) );
NAND3_X1 U908 ( .A1(n1040), .A2(n1019), .A3(n1039), .ZN(n1196) );
XNOR2_X1 U909 ( .A(G125), .B(n1173), .ZN(G27) );
NAND3_X1 U910 ( .A1(n1062), .A2(n1209), .A3(n1240), .ZN(n1173) );
NOR3_X1 U911 ( .A1(n1241), .A2(n1235), .A3(n1227), .ZN(n1240) );
INV_X1 U912 ( .A(n1183), .ZN(n1227) );
NAND2_X1 U913 ( .A1(n1032), .A2(n1242), .ZN(n1183) );
NAND3_X1 U914 ( .A1(G902), .A2(n1243), .A3(n1101), .ZN(n1242) );
NOR2_X1 U915 ( .A1(n1049), .A2(G900), .ZN(n1101) );
XNOR2_X1 U916 ( .A(G122), .B(n1244), .ZN(G24) );
NAND2_X1 U917 ( .A1(KEYINPUT42), .A2(n1193), .ZN(n1244) );
AND3_X1 U918 ( .A1(n1062), .A2(n1021), .A3(n1245), .ZN(n1193) );
NOR3_X1 U919 ( .A1(n1224), .A2(n1246), .A3(n1225), .ZN(n1245) );
NOR2_X1 U920 ( .A1(n1230), .A2(n1241), .ZN(n1021) );
INV_X1 U921 ( .A(n1229), .ZN(n1241) );
XOR2_X1 U922 ( .A(G119), .B(n1195), .Z(G21) );
AND4_X1 U923 ( .A1(n1186), .A2(n1039), .A3(n1064), .A4(n1200), .ZN(n1195) );
NOR3_X1 U924 ( .A1(n1226), .A2(n1235), .A3(n1229), .ZN(n1186) );
INV_X1 U925 ( .A(n1230), .ZN(n1235) );
XNOR2_X1 U926 ( .A(G116), .B(n1198), .ZN(G18) );
NAND4_X1 U927 ( .A1(n1062), .A2(n1040), .A3(n1020), .A4(n1200), .ZN(n1198) );
NOR2_X1 U928 ( .A1(n1247), .A2(n1224), .ZN(n1020) );
XNOR2_X1 U929 ( .A(n1084), .B(KEYINPUT34), .ZN(n1224) );
NOR2_X1 U930 ( .A1(n1030), .A2(n1226), .ZN(n1062) );
XOR2_X1 U931 ( .A(n1192), .B(n1248), .Z(G15) );
NOR2_X1 U932 ( .A1(KEYINPUT0), .A2(n1249), .ZN(n1248) );
AND4_X1 U933 ( .A1(n1040), .A2(n1209), .A3(n1064), .A4(n1250), .ZN(n1192) );
INV_X1 U934 ( .A(n1030), .ZN(n1064) );
NAND2_X1 U935 ( .A1(n1060), .A2(n1251), .ZN(n1030) );
INV_X1 U936 ( .A(n1081), .ZN(n1060) );
AND2_X1 U937 ( .A1(n1084), .A2(n1247), .ZN(n1209) );
INV_X1 U938 ( .A(n1225), .ZN(n1247) );
NOR2_X1 U939 ( .A1(n1229), .A2(n1230), .ZN(n1040) );
XNOR2_X1 U940 ( .A(G110), .B(n1252), .ZN(G12) );
NAND3_X1 U941 ( .A1(n1253), .A2(n1254), .A3(n1041), .ZN(n1252) );
INV_X1 U942 ( .A(n1046), .ZN(n1041) );
NAND3_X1 U943 ( .A1(n1229), .A2(n1230), .A3(n1039), .ZN(n1046) );
AND2_X1 U944 ( .A1(n1225), .A2(n1084), .ZN(n1039) );
XOR2_X1 U945 ( .A(n1255), .B(G478), .Z(n1084) );
NAND2_X1 U946 ( .A1(n1133), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U947 ( .A(n1257), .B(n1258), .ZN(n1133) );
XNOR2_X1 U948 ( .A(n1259), .B(n1260), .ZN(n1258) );
XNOR2_X1 U949 ( .A(n1218), .B(G134), .ZN(n1260) );
XOR2_X1 U950 ( .A(n1261), .B(n1262), .Z(n1257) );
NOR2_X1 U951 ( .A1(KEYINPUT11), .A2(n1263), .ZN(n1262) );
XNOR2_X1 U952 ( .A(n1264), .B(n1265), .ZN(n1263) );
XOR2_X1 U953 ( .A(KEYINPUT35), .B(G122), .Z(n1265) );
XOR2_X1 U954 ( .A(n1266), .B(G107), .Z(n1261) );
NAND3_X1 U955 ( .A1(G217), .A2(n1049), .A3(n1267), .ZN(n1266) );
NOR2_X1 U956 ( .A1(n1090), .A2(n1268), .ZN(n1225) );
AND2_X1 U957 ( .A1(G475), .A2(n1269), .ZN(n1268) );
NAND2_X1 U958 ( .A1(n1270), .A2(n1256), .ZN(n1269) );
INV_X1 U959 ( .A(n1094), .ZN(n1270) );
NOR3_X1 U960 ( .A1(G475), .A2(G902), .A3(n1094), .ZN(n1090) );
XNOR2_X1 U961 ( .A(n1271), .B(n1272), .ZN(n1094) );
XOR2_X1 U962 ( .A(n1273), .B(n1105), .Z(n1272) );
XNOR2_X1 U963 ( .A(G131), .B(n1274), .ZN(n1105) );
NAND2_X1 U964 ( .A1(KEYINPUT1), .A2(n1218), .ZN(n1273) );
INV_X1 U965 ( .A(G143), .ZN(n1218) );
XOR2_X1 U966 ( .A(n1275), .B(n1276), .Z(n1271) );
NOR2_X1 U967 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
INV_X1 U968 ( .A(G214), .ZN(n1278) );
XNOR2_X1 U969 ( .A(n1279), .B(n1280), .ZN(n1275) );
NAND2_X1 U970 ( .A1(n1281), .A2(n1282), .ZN(n1279) );
NAND2_X1 U971 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
XOR2_X1 U972 ( .A(KEYINPUT18), .B(n1285), .Z(n1281) );
NOR2_X1 U973 ( .A1(n1284), .A2(n1283), .ZN(n1285) );
XOR2_X1 U974 ( .A(KEYINPUT27), .B(G104), .Z(n1283) );
XNOR2_X1 U975 ( .A(n1249), .B(G122), .ZN(n1284) );
INV_X1 U976 ( .A(G113), .ZN(n1249) );
NAND3_X1 U977 ( .A1(n1286), .A2(n1287), .A3(n1079), .ZN(n1230) );
NAND2_X1 U978 ( .A1(n1288), .A2(n1289), .ZN(n1079) );
OR2_X1 U979 ( .A1(n1130), .A2(KEYINPUT28), .ZN(n1287) );
INV_X1 U980 ( .A(n1289), .ZN(n1130) );
NAND2_X1 U981 ( .A1(n1080), .A2(KEYINPUT28), .ZN(n1286) );
NOR2_X1 U982 ( .A1(n1289), .A2(n1288), .ZN(n1080) );
AND2_X1 U983 ( .A1(n1128), .A2(n1256), .ZN(n1288) );
XOR2_X1 U984 ( .A(n1290), .B(n1291), .Z(n1128) );
XOR2_X1 U985 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U986 ( .A(n1259), .B(G119), .ZN(n1293) );
XNOR2_X1 U987 ( .A(KEYINPUT16), .B(n1231), .ZN(n1292) );
XOR2_X1 U988 ( .A(n1294), .B(n1295), .Z(n1290) );
XOR2_X1 U989 ( .A(n1296), .B(n1274), .Z(n1295) );
XOR2_X1 U990 ( .A(G140), .B(G125), .Z(n1274) );
NOR2_X1 U991 ( .A1(G110), .A2(KEYINPUT44), .ZN(n1296) );
XOR2_X1 U992 ( .A(n1297), .B(n1298), .Z(n1294) );
NOR2_X1 U993 ( .A1(KEYINPUT47), .A2(n1280), .ZN(n1298) );
NAND3_X1 U994 ( .A1(n1267), .A2(n1049), .A3(G221), .ZN(n1297) );
XNOR2_X1 U995 ( .A(G234), .B(KEYINPUT24), .ZN(n1267) );
NAND2_X1 U996 ( .A1(G217), .A2(n1299), .ZN(n1289) );
XOR2_X1 U997 ( .A(n1300), .B(n1074), .Z(n1229) );
NAND2_X1 U998 ( .A1(n1301), .A2(n1256), .ZN(n1074) );
XNOR2_X1 U999 ( .A(n1141), .B(n1302), .ZN(n1301) );
XNOR2_X1 U1000 ( .A(n1142), .B(n1145), .ZN(n1302) );
INV_X1 U1001 ( .A(G101), .ZN(n1142) );
XNOR2_X1 U1002 ( .A(n1303), .B(n1304), .ZN(n1141) );
NOR2_X1 U1003 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
NOR2_X1 U1004 ( .A1(G119), .A2(n1307), .ZN(n1306) );
XOR2_X1 U1005 ( .A(KEYINPUT48), .B(n1308), .Z(n1307) );
AND2_X1 U1006 ( .A1(G119), .A2(n1308), .ZN(n1305) );
XOR2_X1 U1007 ( .A(n1309), .B(n1310), .Z(n1303) );
NOR2_X1 U1008 ( .A1(n1277), .A2(n1311), .ZN(n1310) );
INV_X1 U1009 ( .A(G210), .ZN(n1311) );
NAND2_X1 U1010 ( .A1(n1049), .A2(n1312), .ZN(n1277) );
NAND2_X1 U1011 ( .A1(KEYINPUT9), .A2(n1076), .ZN(n1300) );
INV_X1 U1012 ( .A(G472), .ZN(n1076) );
OR2_X1 U1013 ( .A1(n1019), .A2(KEYINPUT40), .ZN(n1254) );
AND2_X1 U1014 ( .A1(n1250), .A2(n1204), .ZN(n1019) );
INV_X1 U1015 ( .A(n1187), .ZN(n1204) );
NAND2_X1 U1016 ( .A1(KEYINPUT40), .A2(n1313), .ZN(n1253) );
NAND2_X1 U1017 ( .A1(n1250), .A2(n1187), .ZN(n1313) );
NAND2_X1 U1018 ( .A1(n1081), .A2(n1251), .ZN(n1187) );
XNOR2_X1 U1019 ( .A(n1061), .B(KEYINPUT56), .ZN(n1251) );
NAND2_X1 U1020 ( .A1(G221), .A2(n1299), .ZN(n1061) );
NAND2_X1 U1021 ( .A1(G234), .A2(n1256), .ZN(n1299) );
XNOR2_X1 U1022 ( .A(n1314), .B(G469), .ZN(n1081) );
NAND2_X1 U1023 ( .A1(n1315), .A2(n1256), .ZN(n1314) );
XOR2_X1 U1024 ( .A(n1164), .B(n1316), .Z(n1315) );
XOR2_X1 U1025 ( .A(n1317), .B(n1318), .Z(n1316) );
NOR2_X1 U1026 ( .A1(KEYINPUT21), .A2(n1123), .ZN(n1318) );
NOR2_X1 U1027 ( .A1(n1158), .A2(n1319), .ZN(n1317) );
NOR2_X1 U1028 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
XNOR2_X1 U1029 ( .A(KEYINPUT55), .B(n1161), .ZN(n1321) );
NOR2_X1 U1030 ( .A1(n1161), .A2(n1160), .ZN(n1158) );
INV_X1 U1031 ( .A(n1320), .ZN(n1160) );
NAND2_X1 U1032 ( .A1(G227), .A2(n1049), .ZN(n1320) );
XNOR2_X1 U1033 ( .A(G140), .B(G110), .ZN(n1161) );
XOR2_X1 U1034 ( .A(n1309), .B(n1322), .Z(n1164) );
XOR2_X1 U1035 ( .A(KEYINPUT15), .B(n1102), .Z(n1322) );
XOR2_X1 U1036 ( .A(n1323), .B(n1324), .Z(n1102) );
XNOR2_X1 U1037 ( .A(n1325), .B(KEYINPUT50), .ZN(n1324) );
NAND2_X1 U1038 ( .A1(KEYINPUT57), .A2(n1259), .ZN(n1325) );
INV_X1 U1039 ( .A(G128), .ZN(n1259) );
XOR2_X1 U1040 ( .A(n1326), .B(n1327), .Z(n1309) );
XOR2_X1 U1041 ( .A(KEYINPUT10), .B(G131), .Z(n1327) );
NAND3_X1 U1042 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1326) );
OR2_X1 U1043 ( .A1(n1231), .A2(n1331), .ZN(n1330) );
NAND3_X1 U1044 ( .A1(n1331), .A2(n1231), .A3(KEYINPUT22), .ZN(n1329) );
INV_X1 U1045 ( .A(G137), .ZN(n1231) );
NOR2_X1 U1046 ( .A1(G134), .A2(KEYINPUT36), .ZN(n1331) );
NAND2_X1 U1047 ( .A1(G134), .A2(n1332), .ZN(n1328) );
INV_X1 U1048 ( .A(KEYINPUT22), .ZN(n1332) );
NOR2_X1 U1049 ( .A1(n1203), .A2(n1246), .ZN(n1250) );
INV_X1 U1050 ( .A(n1200), .ZN(n1246) );
NAND2_X1 U1051 ( .A1(n1032), .A2(n1333), .ZN(n1200) );
NAND4_X1 U1052 ( .A1(n1334), .A2(G953), .A3(G902), .A4(n1243), .ZN(n1333) );
XNOR2_X1 U1053 ( .A(G898), .B(KEYINPUT63), .ZN(n1334) );
NAND3_X1 U1054 ( .A1(n1243), .A2(n1049), .A3(G952), .ZN(n1032) );
NAND2_X1 U1055 ( .A1(G237), .A2(G234), .ZN(n1243) );
XOR2_X1 U1056 ( .A(n1226), .B(KEYINPUT45), .Z(n1203) );
INV_X1 U1057 ( .A(n1205), .ZN(n1226) );
NOR2_X1 U1058 ( .A1(n1063), .A2(n1065), .ZN(n1205) );
INV_X1 U1059 ( .A(n1239), .ZN(n1065) );
NAND2_X1 U1060 ( .A1(G214), .A2(n1335), .ZN(n1239) );
NOR2_X1 U1061 ( .A1(n1089), .A2(n1336), .ZN(n1063) );
AND2_X1 U1062 ( .A1(n1085), .A2(n1086), .ZN(n1336) );
NOR2_X1 U1063 ( .A1(n1086), .A2(n1085), .ZN(n1089) );
INV_X1 U1064 ( .A(n1088), .ZN(n1085) );
NAND2_X1 U1065 ( .A1(G210), .A2(n1335), .ZN(n1088) );
NAND2_X1 U1066 ( .A1(n1256), .A2(n1312), .ZN(n1335) );
INV_X1 U1067 ( .A(G237), .ZN(n1312) );
NAND2_X1 U1068 ( .A1(n1337), .A2(n1256), .ZN(n1086) );
INV_X1 U1069 ( .A(G902), .ZN(n1256) );
XNOR2_X1 U1070 ( .A(n1338), .B(n1339), .ZN(n1337) );
INV_X1 U1071 ( .A(n1215), .ZN(n1339) );
XNOR2_X1 U1072 ( .A(n1340), .B(n1117), .ZN(n1215) );
XOR2_X1 U1073 ( .A(G110), .B(G122), .Z(n1117) );
XNOR2_X1 U1074 ( .A(n1122), .B(n1121), .ZN(n1340) );
INV_X1 U1075 ( .A(n1123), .ZN(n1121) );
XOR2_X1 U1076 ( .A(G101), .B(n1341), .Z(n1123) );
XOR2_X1 U1077 ( .A(G107), .B(G104), .Z(n1341) );
XNOR2_X1 U1078 ( .A(G119), .B(n1308), .ZN(n1122) );
XNOR2_X1 U1079 ( .A(G113), .B(n1264), .ZN(n1308) );
INV_X1 U1080 ( .A(G116), .ZN(n1264) );
XNOR2_X1 U1081 ( .A(n1213), .B(KEYINPUT23), .ZN(n1338) );
AND2_X1 U1082 ( .A1(n1342), .A2(n1343), .ZN(n1213) );
NAND3_X1 U1083 ( .A1(G224), .A2(n1049), .A3(n1344), .ZN(n1343) );
XNOR2_X1 U1084 ( .A(G125), .B(n1145), .ZN(n1344) );
NAND2_X1 U1085 ( .A1(n1345), .A2(n1346), .ZN(n1342) );
NAND2_X1 U1086 ( .A1(G224), .A2(n1049), .ZN(n1346) );
INV_X1 U1087 ( .A(G953), .ZN(n1049) );
XOR2_X1 U1088 ( .A(G125), .B(n1145), .Z(n1345) );
XNOR2_X1 U1089 ( .A(n1347), .B(n1323), .ZN(n1145) );
XNOR2_X1 U1090 ( .A(G143), .B(n1280), .ZN(n1323) );
INV_X1 U1091 ( .A(G146), .ZN(n1280) );
XNOR2_X1 U1092 ( .A(G128), .B(KEYINPUT3), .ZN(n1347) );
endmodule


