//Key = 0100100010011010111110100010001001001001110101000110011010101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
n1424;

XNOR2_X1 U789 ( .A(G107), .B(n1094), .ZN(G9) );
NOR2_X1 U790 ( .A1(n1095), .A2(n1096), .ZN(G75) );
NOR4_X1 U791 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
XOR2_X1 U792 ( .A(n1101), .B(KEYINPUT14), .Z(n1099) );
NAND2_X1 U793 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U794 ( .A(n1104), .B(KEYINPUT40), .Z(n1102) );
NAND4_X1 U795 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1104) );
INV_X1 U796 ( .A(n1109), .ZN(n1098) );
NAND4_X1 U797 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1097) );
NAND3_X1 U798 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1112) );
NAND3_X1 U799 ( .A1(n1103), .A2(n1117), .A3(n1105), .ZN(n1111) );
NAND2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U801 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
NAND2_X1 U802 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NAND2_X1 U803 ( .A1(n1108), .A2(n1124), .ZN(n1123) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NAND2_X1 U805 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U806 ( .A1(n1106), .A2(n1129), .ZN(n1122) );
OR2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U808 ( .A1(n1132), .A2(n1108), .ZN(n1118) );
NAND2_X1 U809 ( .A1(n1133), .A2(n1134), .ZN(n1110) );
XNOR2_X1 U810 ( .A(n1116), .B(KEYINPUT26), .ZN(n1133) );
AND4_X1 U811 ( .A1(n1105), .A2(n1106), .A3(n1120), .A4(n1108), .ZN(n1116) );
INV_X1 U812 ( .A(n1135), .ZN(n1105) );
AND3_X1 U813 ( .A1(n1136), .A2(n1137), .A3(n1113), .ZN(n1095) );
NAND4_X1 U814 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1113) );
NOR4_X1 U815 ( .A1(n1142), .A2(n1115), .A3(n1127), .A4(n1143), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U817 ( .A1(G902), .A2(n1146), .ZN(n1144) );
NOR2_X1 U818 ( .A1(n1147), .A2(n1148), .ZN(n1140) );
XNOR2_X1 U819 ( .A(KEYINPUT62), .B(n1114), .ZN(n1148) );
XNOR2_X1 U820 ( .A(KEYINPUT41), .B(n1128), .ZN(n1139) );
XOR2_X1 U821 ( .A(n1149), .B(n1150), .Z(G72) );
NAND2_X1 U822 ( .A1(KEYINPUT18), .A2(n1151), .ZN(n1150) );
XOR2_X1 U823 ( .A(n1152), .B(n1153), .Z(n1151) );
NAND2_X1 U824 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
NAND2_X1 U825 ( .A1(n1156), .A2(n1157), .ZN(n1152) );
NAND2_X1 U826 ( .A1(G953), .A2(n1158), .ZN(n1157) );
XOR2_X1 U827 ( .A(n1159), .B(n1160), .Z(n1156) );
XNOR2_X1 U828 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U829 ( .A1(G140), .A2(KEYINPUT13), .ZN(n1161) );
XOR2_X1 U830 ( .A(n1163), .B(n1164), .Z(n1159) );
NOR2_X1 U831 ( .A1(KEYINPUT31), .A2(n1165), .ZN(n1164) );
XNOR2_X1 U832 ( .A(n1166), .B(n1167), .ZN(n1165) );
XNOR2_X1 U833 ( .A(n1168), .B(G125), .ZN(n1163) );
INV_X1 U834 ( .A(n1169), .ZN(n1168) );
NAND2_X1 U835 ( .A1(G953), .A2(n1170), .ZN(n1149) );
XOR2_X1 U836 ( .A(KEYINPUT43), .B(n1171), .Z(n1170) );
AND2_X1 U837 ( .A1(G227), .A2(G900), .ZN(n1171) );
XOR2_X1 U838 ( .A(n1172), .B(n1173), .Z(G69) );
XOR2_X1 U839 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U840 ( .A1(G953), .A2(n1176), .ZN(n1175) );
NAND2_X1 U841 ( .A1(G898), .A2(G224), .ZN(n1176) );
NAND2_X1 U842 ( .A1(n1177), .A2(n1178), .ZN(n1174) );
NAND2_X1 U843 ( .A1(G953), .A2(n1179), .ZN(n1178) );
XOR2_X1 U844 ( .A(n1180), .B(n1181), .Z(n1177) );
AND2_X1 U845 ( .A1(n1182), .A2(n1154), .ZN(n1172) );
NOR2_X1 U846 ( .A1(n1183), .A2(n1184), .ZN(G66) );
XOR2_X1 U847 ( .A(n1185), .B(n1186), .Z(n1184) );
NAND3_X1 U848 ( .A1(n1187), .A2(G217), .A3(KEYINPUT54), .ZN(n1185) );
NOR2_X1 U849 ( .A1(n1183), .A2(n1188), .ZN(G63) );
XNOR2_X1 U850 ( .A(n1189), .B(n1146), .ZN(n1188) );
NAND3_X1 U851 ( .A1(n1187), .A2(G478), .A3(KEYINPUT49), .ZN(n1189) );
NOR2_X1 U852 ( .A1(n1183), .A2(n1190), .ZN(G60) );
XNOR2_X1 U853 ( .A(n1191), .B(n1192), .ZN(n1190) );
NOR3_X1 U854 ( .A1(n1193), .A2(n1109), .A3(n1194), .ZN(n1192) );
XNOR2_X1 U855 ( .A(G902), .B(KEYINPUT23), .ZN(n1194) );
XOR2_X1 U856 ( .A(G104), .B(n1195), .Z(G6) );
NOR2_X1 U857 ( .A1(n1183), .A2(n1196), .ZN(G57) );
XOR2_X1 U858 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U859 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
XOR2_X1 U860 ( .A(KEYINPUT27), .B(n1201), .Z(n1200) );
NOR2_X1 U861 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U862 ( .A1(n1204), .A2(n1205), .ZN(n1199) );
XNOR2_X1 U863 ( .A(n1203), .B(KEYINPUT32), .ZN(n1205) );
XOR2_X1 U864 ( .A(n1206), .B(n1207), .Z(n1203) );
XOR2_X1 U865 ( .A(n1208), .B(n1209), .Z(n1206) );
NAND2_X1 U866 ( .A1(KEYINPUT39), .A2(n1210), .ZN(n1208) );
XOR2_X1 U867 ( .A(n1202), .B(KEYINPUT50), .Z(n1204) );
NAND2_X1 U868 ( .A1(n1187), .A2(G472), .ZN(n1202) );
NOR2_X1 U869 ( .A1(n1183), .A2(n1211), .ZN(G54) );
XOR2_X1 U870 ( .A(n1212), .B(n1213), .Z(n1211) );
AND2_X1 U871 ( .A1(G469), .A2(n1187), .ZN(n1213) );
NAND2_X1 U872 ( .A1(KEYINPUT60), .A2(n1214), .ZN(n1212) );
XOR2_X1 U873 ( .A(n1215), .B(n1216), .Z(n1214) );
XNOR2_X1 U874 ( .A(n1217), .B(n1218), .ZN(n1216) );
XOR2_X1 U875 ( .A(n1219), .B(n1220), .Z(n1215) );
XNOR2_X1 U876 ( .A(n1169), .B(n1221), .ZN(n1220) );
NOR2_X1 U877 ( .A1(KEYINPUT10), .A2(n1222), .ZN(n1221) );
XNOR2_X1 U878 ( .A(G140), .B(G110), .ZN(n1222) );
NOR2_X1 U879 ( .A1(KEYINPUT0), .A2(n1223), .ZN(n1219) );
XNOR2_X1 U880 ( .A(n1224), .B(KEYINPUT1), .ZN(n1223) );
NOR4_X1 U881 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(G51) );
NOR3_X1 U882 ( .A1(n1229), .A2(n1154), .A3(n1137), .ZN(n1228) );
INV_X1 U883 ( .A(G952), .ZN(n1137) );
AND2_X1 U884 ( .A1(n1229), .A2(n1183), .ZN(n1227) );
NOR2_X1 U885 ( .A1(n1154), .A2(G952), .ZN(n1183) );
INV_X1 U886 ( .A(KEYINPUT57), .ZN(n1229) );
NOR3_X1 U887 ( .A1(KEYINPUT44), .A2(n1230), .A3(n1231), .ZN(n1226) );
NOR2_X1 U888 ( .A1(n1232), .A2(n1233), .ZN(n1230) );
XNOR2_X1 U889 ( .A(KEYINPUT30), .B(n1234), .ZN(n1233) );
NOR2_X1 U890 ( .A1(n1235), .A2(n1236), .ZN(n1225) );
INV_X1 U891 ( .A(KEYINPUT44), .ZN(n1236) );
NOR2_X1 U892 ( .A1(n1237), .A2(n1238), .ZN(n1235) );
AND2_X1 U893 ( .A1(KEYINPUT30), .A2(n1231), .ZN(n1238) );
AND2_X1 U894 ( .A1(n1234), .A2(n1232), .ZN(n1231) );
NOR2_X1 U895 ( .A1(n1239), .A2(n1234), .ZN(n1237) );
XOR2_X1 U896 ( .A(n1240), .B(n1241), .Z(n1234) );
NOR2_X1 U897 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U898 ( .A(n1244), .B(KEYINPUT33), .Z(n1243) );
NAND2_X1 U899 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
NOR2_X1 U900 ( .A1(n1245), .A2(n1246), .ZN(n1242) );
XOR2_X1 U901 ( .A(KEYINPUT8), .B(n1247), .Z(n1246) );
NAND2_X1 U902 ( .A1(n1187), .A2(n1248), .ZN(n1240) );
NOR2_X1 U903 ( .A1(n1249), .A2(n1109), .ZN(n1187) );
NOR2_X1 U904 ( .A1(n1182), .A2(n1155), .ZN(n1109) );
NAND4_X1 U905 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1155) );
AND4_X1 U906 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1253) );
NOR3_X1 U907 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1252) );
NOR2_X1 U908 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
INV_X1 U909 ( .A(KEYINPUT4), .ZN(n1261) );
NOR2_X1 U910 ( .A1(KEYINPUT4), .A2(n1263), .ZN(n1259) );
NAND4_X1 U911 ( .A1(n1132), .A2(n1130), .A3(n1264), .A4(n1265), .ZN(n1263) );
NOR2_X1 U912 ( .A1(n1266), .A2(n1267), .ZN(n1258) );
NAND4_X1 U913 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1250) );
NAND2_X1 U914 ( .A1(n1103), .A2(n1272), .ZN(n1271) );
NAND2_X1 U915 ( .A1(n1273), .A2(n1274), .ZN(n1270) );
NAND2_X1 U916 ( .A1(n1130), .A2(n1267), .ZN(n1273) );
INV_X1 U917 ( .A(KEYINPUT22), .ZN(n1267) );
NAND4_X1 U918 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1182) );
AND4_X1 U919 ( .A1(n1094), .A2(n1279), .A3(n1280), .A4(n1281), .ZN(n1278) );
NAND2_X1 U920 ( .A1(n1107), .A2(n1282), .ZN(n1094) );
NOR2_X1 U921 ( .A1(n1283), .A2(n1195), .ZN(n1277) );
AND2_X1 U922 ( .A1(n1269), .A2(n1282), .ZN(n1195) );
NOR3_X1 U923 ( .A1(n1284), .A2(n1147), .A3(n1125), .ZN(n1282) );
NOR2_X1 U924 ( .A1(n1285), .A2(n1286), .ZN(n1283) );
XNOR2_X1 U925 ( .A(KEYINPUT19), .B(n1125), .ZN(n1286) );
NAND4_X1 U926 ( .A1(n1132), .A2(n1131), .A3(n1287), .A4(n1288), .ZN(n1275) );
OR2_X1 U927 ( .A1(n1289), .A2(KEYINPUT63), .ZN(n1288) );
NAND2_X1 U928 ( .A1(KEYINPUT63), .A2(n1290), .ZN(n1287) );
NAND2_X1 U929 ( .A1(n1265), .A2(n1291), .ZN(n1290) );
AND2_X1 U930 ( .A1(n1232), .A2(KEYINPUT30), .ZN(n1239) );
XOR2_X1 U931 ( .A(n1257), .B(n1292), .Z(G48) );
XOR2_X1 U932 ( .A(KEYINPUT56), .B(G146), .Z(n1292) );
NAND3_X1 U933 ( .A1(n1269), .A2(n1134), .A3(n1293), .ZN(n1257) );
XOR2_X1 U934 ( .A(n1256), .B(n1294), .Z(G45) );
XNOR2_X1 U935 ( .A(G143), .B(KEYINPUT29), .ZN(n1294) );
NAND3_X1 U936 ( .A1(n1268), .A2(n1131), .A3(n1295), .ZN(n1256) );
NOR3_X1 U937 ( .A1(n1265), .A2(n1296), .A3(n1138), .ZN(n1295) );
INV_X1 U938 ( .A(n1134), .ZN(n1265) );
XNOR2_X1 U939 ( .A(G140), .B(n1266), .ZN(G42) );
NAND4_X1 U940 ( .A1(n1103), .A2(n1268), .A3(n1269), .A4(n1130), .ZN(n1266) );
XNOR2_X1 U941 ( .A(G137), .B(n1251), .ZN(G39) );
NAND3_X1 U942 ( .A1(n1293), .A2(n1120), .A3(n1103), .ZN(n1251) );
XNOR2_X1 U943 ( .A(G134), .B(n1255), .ZN(G36) );
NAND4_X1 U944 ( .A1(n1103), .A2(n1268), .A3(n1131), .A4(n1107), .ZN(n1255) );
XNOR2_X1 U945 ( .A(G131), .B(n1297), .ZN(G33) );
NAND4_X1 U946 ( .A1(n1131), .A2(n1298), .A3(n1269), .A4(n1299), .ZN(n1297) );
NOR2_X1 U947 ( .A1(n1274), .A2(n1300), .ZN(n1299) );
XNOR2_X1 U948 ( .A(KEYINPUT34), .B(n1264), .ZN(n1300) );
INV_X1 U949 ( .A(n1103), .ZN(n1274) );
NOR2_X1 U950 ( .A1(n1301), .A2(n1115), .ZN(n1103) );
XNOR2_X1 U951 ( .A(G128), .B(n1254), .ZN(G30) );
NAND3_X1 U952 ( .A1(n1107), .A2(n1134), .A3(n1293), .ZN(n1254) );
AND3_X1 U953 ( .A1(n1302), .A2(n1303), .A3(n1268), .ZN(n1293) );
AND2_X1 U954 ( .A1(n1298), .A2(n1264), .ZN(n1268) );
XNOR2_X1 U955 ( .A(G101), .B(n1281), .ZN(G3) );
NAND3_X1 U956 ( .A1(n1304), .A2(n1298), .A3(n1131), .ZN(n1281) );
XNOR2_X1 U957 ( .A(G125), .B(n1262), .ZN(G27) );
NAND4_X1 U958 ( .A1(n1132), .A2(n1130), .A3(n1134), .A4(n1264), .ZN(n1262) );
NAND2_X1 U959 ( .A1(n1135), .A2(n1305), .ZN(n1264) );
NAND4_X1 U960 ( .A1(G902), .A2(G953), .A3(n1306), .A4(n1158), .ZN(n1305) );
INV_X1 U961 ( .A(G900), .ZN(n1158) );
XOR2_X1 U962 ( .A(n1280), .B(n1307), .Z(G24) );
NOR2_X1 U963 ( .A1(G122), .A2(KEYINPUT2), .ZN(n1307) );
NAND3_X1 U964 ( .A1(n1106), .A2(n1289), .A3(n1308), .ZN(n1280) );
NOR3_X1 U965 ( .A1(n1147), .A2(n1296), .A3(n1138), .ZN(n1308) );
INV_X1 U966 ( .A(n1108), .ZN(n1147) );
NOR2_X1 U967 ( .A1(n1303), .A2(n1302), .ZN(n1108) );
XNOR2_X1 U968 ( .A(G119), .B(n1279), .ZN(G21) );
NAND4_X1 U969 ( .A1(n1106), .A2(n1304), .A3(n1302), .A4(n1303), .ZN(n1279) );
XNOR2_X1 U970 ( .A(G116), .B(n1309), .ZN(G18) );
NOR2_X1 U971 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
NOR2_X1 U972 ( .A1(n1312), .A2(n1276), .ZN(n1311) );
NAND4_X1 U973 ( .A1(n1131), .A2(n1106), .A3(n1107), .A4(n1289), .ZN(n1276) );
INV_X1 U974 ( .A(KEYINPUT16), .ZN(n1312) );
NOR2_X1 U975 ( .A1(KEYINPUT16), .A2(n1313), .ZN(n1310) );
NAND4_X1 U976 ( .A1(n1131), .A2(n1107), .A3(n1289), .A4(n1314), .ZN(n1313) );
INV_X1 U977 ( .A(n1106), .ZN(n1314) );
NOR2_X1 U978 ( .A1(n1315), .A2(n1296), .ZN(n1107) );
NAND2_X1 U979 ( .A1(n1316), .A2(n1317), .ZN(G15) );
NAND2_X1 U980 ( .A1(G113), .A2(n1318), .ZN(n1317) );
XOR2_X1 U981 ( .A(n1319), .B(KEYINPUT51), .Z(n1316) );
OR2_X1 U982 ( .A1(n1318), .A2(G113), .ZN(n1319) );
NAND3_X1 U983 ( .A1(n1131), .A2(n1289), .A3(n1132), .ZN(n1318) );
AND2_X1 U984 ( .A1(n1269), .A2(n1106), .ZN(n1132) );
NOR2_X1 U985 ( .A1(n1320), .A2(n1127), .ZN(n1106) );
AND2_X1 U986 ( .A1(n1296), .A2(n1315), .ZN(n1269) );
INV_X1 U987 ( .A(n1272), .ZN(n1131) );
NAND2_X1 U988 ( .A1(n1321), .A2(n1302), .ZN(n1272) );
XOR2_X1 U989 ( .A(G110), .B(n1322), .Z(G12) );
NOR2_X1 U990 ( .A1(n1125), .A2(n1285), .ZN(n1322) );
NAND2_X1 U991 ( .A1(n1130), .A2(n1304), .ZN(n1285) );
AND2_X1 U992 ( .A1(n1120), .A2(n1289), .ZN(n1304) );
INV_X1 U993 ( .A(n1284), .ZN(n1289) );
NAND2_X1 U994 ( .A1(n1134), .A2(n1291), .ZN(n1284) );
NAND2_X1 U995 ( .A1(n1323), .A2(n1135), .ZN(n1291) );
NAND3_X1 U996 ( .A1(n1136), .A2(n1306), .A3(G952), .ZN(n1135) );
INV_X1 U997 ( .A(n1100), .ZN(n1136) );
XOR2_X1 U998 ( .A(G953), .B(KEYINPUT37), .Z(n1100) );
NAND4_X1 U999 ( .A1(G902), .A2(G953), .A3(n1306), .A4(n1179), .ZN(n1323) );
INV_X1 U1000 ( .A(G898), .ZN(n1179) );
NAND2_X1 U1001 ( .A1(G237), .A2(G234), .ZN(n1306) );
NOR2_X1 U1002 ( .A1(n1114), .A2(n1115), .ZN(n1134) );
AND2_X1 U1003 ( .A1(G214), .A2(n1324), .ZN(n1115) );
INV_X1 U1004 ( .A(n1301), .ZN(n1114) );
XNOR2_X1 U1005 ( .A(n1325), .B(n1248), .ZN(n1301) );
AND2_X1 U1006 ( .A1(G210), .A2(n1324), .ZN(n1248) );
NAND2_X1 U1007 ( .A1(n1326), .A2(n1249), .ZN(n1324) );
XNOR2_X1 U1008 ( .A(G237), .B(KEYINPUT47), .ZN(n1326) );
NAND2_X1 U1009 ( .A1(n1327), .A2(n1249), .ZN(n1325) );
XNOR2_X1 U1010 ( .A(n1247), .B(n1328), .ZN(n1327) );
XOR2_X1 U1011 ( .A(n1245), .B(n1232), .Z(n1328) );
XNOR2_X1 U1012 ( .A(n1329), .B(n1180), .ZN(n1232) );
NAND2_X1 U1013 ( .A1(n1330), .A2(n1331), .ZN(n1180) );
NAND2_X1 U1014 ( .A1(G110), .A2(n1332), .ZN(n1331) );
XOR2_X1 U1015 ( .A(n1333), .B(KEYINPUT28), .Z(n1330) );
OR2_X1 U1016 ( .A1(n1332), .A2(G110), .ZN(n1333) );
NAND2_X1 U1017 ( .A1(KEYINPUT36), .A2(n1181), .ZN(n1329) );
XOR2_X1 U1018 ( .A(n1334), .B(n1335), .Z(n1181) );
XNOR2_X1 U1019 ( .A(n1336), .B(n1337), .ZN(n1335) );
INV_X1 U1020 ( .A(n1338), .ZN(n1336) );
XOR2_X1 U1021 ( .A(n1339), .B(n1340), .Z(n1334) );
XNOR2_X1 U1022 ( .A(n1341), .B(G104), .ZN(n1340) );
NAND2_X1 U1023 ( .A1(n1342), .A2(KEYINPUT61), .ZN(n1339) );
XNOR2_X1 U1024 ( .A(G113), .B(KEYINPUT55), .ZN(n1342) );
AND2_X1 U1025 ( .A1(G224), .A2(n1154), .ZN(n1245) );
XOR2_X1 U1026 ( .A(G125), .B(n1210), .Z(n1247) );
AND2_X1 U1027 ( .A1(n1296), .A2(n1138), .ZN(n1120) );
INV_X1 U1028 ( .A(n1315), .ZN(n1138) );
XOR2_X1 U1029 ( .A(n1343), .B(n1193), .Z(n1315) );
INV_X1 U1030 ( .A(G475), .ZN(n1193) );
NAND2_X1 U1031 ( .A1(n1191), .A2(n1249), .ZN(n1343) );
XNOR2_X1 U1032 ( .A(n1344), .B(n1345), .ZN(n1191) );
XOR2_X1 U1033 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1034 ( .A(G113), .B(G104), .Z(n1347) );
XNOR2_X1 U1035 ( .A(n1348), .B(G122), .ZN(n1346) );
XNOR2_X1 U1036 ( .A(n1349), .B(n1350), .ZN(n1344) );
INV_X1 U1037 ( .A(n1351), .ZN(n1350) );
XNOR2_X1 U1038 ( .A(n1352), .B(n1162), .ZN(n1349) );
INV_X1 U1039 ( .A(n1353), .ZN(n1162) );
NAND2_X1 U1040 ( .A1(G214), .A2(n1354), .ZN(n1352) );
NOR2_X1 U1041 ( .A1(n1355), .A2(n1142), .ZN(n1296) );
NOR3_X1 U1042 ( .A1(G478), .A2(G902), .A3(n1146), .ZN(n1142) );
AND2_X1 U1043 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
OR2_X1 U1044 ( .A1(n1146), .A2(G902), .ZN(n1357) );
XOR2_X1 U1045 ( .A(n1358), .B(n1359), .Z(n1146) );
XNOR2_X1 U1046 ( .A(n1360), .B(n1337), .ZN(n1359) );
XNOR2_X1 U1047 ( .A(G116), .B(n1361), .ZN(n1337) );
NAND2_X1 U1048 ( .A1(G217), .A2(n1362), .ZN(n1360) );
XOR2_X1 U1049 ( .A(n1363), .B(n1364), .Z(n1358) );
XNOR2_X1 U1050 ( .A(G134), .B(n1332), .ZN(n1364) );
INV_X1 U1051 ( .A(G122), .ZN(n1332) );
NAND3_X1 U1052 ( .A1(n1365), .A2(n1366), .A3(n1367), .ZN(n1363) );
NAND2_X1 U1053 ( .A1(n1368), .A2(n1348), .ZN(n1367) );
OR3_X1 U1054 ( .A1(n1348), .A2(n1368), .A3(KEYINPUT35), .ZN(n1366) );
OR2_X1 U1055 ( .A1(KEYINPUT21), .A2(n1369), .ZN(n1368) );
NAND2_X1 U1056 ( .A1(KEYINPUT35), .A2(n1369), .ZN(n1365) );
XNOR2_X1 U1057 ( .A(KEYINPUT42), .B(n1145), .ZN(n1356) );
INV_X1 U1058 ( .A(G478), .ZN(n1145) );
NOR2_X1 U1059 ( .A1(n1302), .A2(n1321), .ZN(n1130) );
INV_X1 U1060 ( .A(n1303), .ZN(n1321) );
NAND3_X1 U1061 ( .A1(n1370), .A2(n1371), .A3(n1372), .ZN(n1303) );
OR2_X1 U1062 ( .A1(n1373), .A2(n1186), .ZN(n1372) );
NAND3_X1 U1063 ( .A1(n1186), .A2(n1373), .A3(n1249), .ZN(n1371) );
NAND2_X1 U1064 ( .A1(G217), .A2(n1374), .ZN(n1373) );
XOR2_X1 U1065 ( .A(n1375), .B(n1376), .Z(n1186) );
XNOR2_X1 U1066 ( .A(n1377), .B(n1351), .ZN(n1376) );
XOR2_X1 U1067 ( .A(G125), .B(n1378), .Z(n1351) );
XOR2_X1 U1068 ( .A(G146), .B(G140), .Z(n1378) );
NAND2_X1 U1069 ( .A1(n1379), .A2(n1380), .ZN(n1377) );
NAND2_X1 U1070 ( .A1(n1166), .A2(n1381), .ZN(n1380) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1362), .ZN(n1381) );
XOR2_X1 U1072 ( .A(n1382), .B(KEYINPUT5), .Z(n1379) );
NAND3_X1 U1073 ( .A1(G221), .A2(n1362), .A3(G137), .ZN(n1382) );
NOR2_X1 U1074 ( .A1(n1374), .A2(G953), .ZN(n1362) );
INV_X1 U1075 ( .A(G234), .ZN(n1374) );
XOR2_X1 U1076 ( .A(n1383), .B(n1384), .Z(n1375) );
NOR2_X1 U1077 ( .A1(KEYINPUT46), .A2(G110), .ZN(n1384) );
XNOR2_X1 U1078 ( .A(G119), .B(G128), .ZN(n1383) );
NAND2_X1 U1079 ( .A1(G902), .A2(G217), .ZN(n1370) );
XNOR2_X1 U1080 ( .A(n1385), .B(G472), .ZN(n1302) );
NAND2_X1 U1081 ( .A1(n1386), .A2(n1249), .ZN(n1385) );
XNOR2_X1 U1082 ( .A(n1209), .B(n1387), .ZN(n1386) );
XNOR2_X1 U1083 ( .A(n1388), .B(n1389), .ZN(n1387) );
NOR2_X1 U1084 ( .A1(KEYINPUT59), .A2(n1198), .ZN(n1389) );
XNOR2_X1 U1085 ( .A(n1390), .B(n1338), .ZN(n1198) );
NAND2_X1 U1086 ( .A1(G210), .A2(n1354), .ZN(n1390) );
NOR2_X1 U1087 ( .A1(G953), .A2(G237), .ZN(n1354) );
NAND2_X1 U1088 ( .A1(KEYINPUT17), .A2(n1391), .ZN(n1388) );
XNOR2_X1 U1089 ( .A(n1210), .B(n1207), .ZN(n1391) );
INV_X1 U1090 ( .A(n1224), .ZN(n1207) );
XNOR2_X1 U1091 ( .A(n1369), .B(n1392), .ZN(n1210) );
NOR2_X1 U1092 ( .A1(KEYINPUT9), .A2(n1393), .ZN(n1392) );
XNOR2_X1 U1093 ( .A(n1348), .B(n1394), .ZN(n1393) );
NOR2_X1 U1094 ( .A1(G146), .A2(KEYINPUT6), .ZN(n1394) );
XNOR2_X1 U1095 ( .A(n1395), .B(n1396), .ZN(n1209) );
XNOR2_X1 U1096 ( .A(n1341), .B(G113), .ZN(n1396) );
INV_X1 U1097 ( .A(G119), .ZN(n1341) );
NAND2_X1 U1098 ( .A1(KEYINPUT45), .A2(G116), .ZN(n1395) );
INV_X1 U1099 ( .A(n1298), .ZN(n1125) );
NOR2_X1 U1100 ( .A1(n1128), .A2(n1127), .ZN(n1298) );
AND2_X1 U1101 ( .A1(G221), .A2(n1397), .ZN(n1127) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1249), .ZN(n1397) );
INV_X1 U1103 ( .A(n1320), .ZN(n1128) );
XNOR2_X1 U1104 ( .A(n1398), .B(G469), .ZN(n1320) );
NAND2_X1 U1105 ( .A1(n1399), .A2(n1249), .ZN(n1398) );
INV_X1 U1106 ( .A(G902), .ZN(n1249) );
XOR2_X1 U1107 ( .A(n1400), .B(n1401), .Z(n1399) );
XNOR2_X1 U1108 ( .A(n1217), .B(n1224), .ZN(n1401) );
XOR2_X1 U1109 ( .A(n1353), .B(n1402), .Z(n1224) );
XNOR2_X1 U1110 ( .A(n1166), .B(n1403), .ZN(n1402) );
NOR2_X1 U1111 ( .A1(KEYINPUT52), .A2(n1167), .ZN(n1403) );
XOR2_X1 U1112 ( .A(G134), .B(KEYINPUT24), .Z(n1167) );
INV_X1 U1113 ( .A(G137), .ZN(n1166) );
XOR2_X1 U1114 ( .A(G131), .B(KEYINPUT25), .Z(n1353) );
NAND2_X1 U1115 ( .A1(G227), .A2(n1154), .ZN(n1217) );
INV_X1 U1116 ( .A(G953), .ZN(n1154) );
XOR2_X1 U1117 ( .A(n1404), .B(n1405), .Z(n1400) );
NOR2_X1 U1118 ( .A1(G110), .A2(n1406), .ZN(n1405) );
XNOR2_X1 U1119 ( .A(KEYINPUT38), .B(KEYINPUT20), .ZN(n1406) );
XNOR2_X1 U1120 ( .A(G140), .B(n1407), .ZN(n1404) );
NOR2_X1 U1121 ( .A1(KEYINPUT48), .A2(n1408), .ZN(n1407) );
XNOR2_X1 U1122 ( .A(n1409), .B(n1169), .ZN(n1408) );
NAND2_X1 U1123 ( .A1(n1410), .A2(n1411), .ZN(n1169) );
OR2_X1 U1124 ( .A1(n1369), .A2(KEYINPUT11), .ZN(n1411) );
XOR2_X1 U1125 ( .A(n1412), .B(n1413), .Z(n1410) );
XNOR2_X1 U1126 ( .A(G146), .B(n1348), .ZN(n1413) );
INV_X1 U1127 ( .A(G143), .ZN(n1348) );
NAND2_X1 U1128 ( .A1(KEYINPUT11), .A2(n1369), .ZN(n1412) );
INV_X1 U1129 ( .A(G128), .ZN(n1369) );
NAND2_X1 U1130 ( .A1(n1414), .A2(n1415), .ZN(n1409) );
NAND2_X1 U1131 ( .A1(KEYINPUT15), .A2(n1416), .ZN(n1415) );
NAND2_X1 U1132 ( .A1(KEYINPUT53), .A2(n1218), .ZN(n1414) );
INV_X1 U1133 ( .A(n1416), .ZN(n1218) );
NAND2_X1 U1134 ( .A1(n1417), .A2(n1418), .ZN(n1416) );
NAND2_X1 U1135 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
XOR2_X1 U1136 ( .A(n1421), .B(KEYINPUT3), .Z(n1417) );
OR2_X1 U1137 ( .A1(n1420), .A2(n1419), .ZN(n1421) );
XOR2_X1 U1138 ( .A(n1338), .B(KEYINPUT58), .Z(n1419) );
XOR2_X1 U1139 ( .A(G101), .B(KEYINPUT12), .Z(n1338) );
NAND2_X1 U1140 ( .A1(n1422), .A2(n1423), .ZN(n1420) );
NAND2_X1 U1141 ( .A1(G104), .A2(n1361), .ZN(n1423) );
XOR2_X1 U1142 ( .A(n1424), .B(KEYINPUT7), .Z(n1422) );
OR2_X1 U1143 ( .A1(n1361), .A2(G104), .ZN(n1424) );
INV_X1 U1144 ( .A(G107), .ZN(n1361) );
endmodule


