//Key = 0110110100011110011100011101111100100111001101001010010001110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327;

XNOR2_X1 U732 ( .A(G107), .B(n1010), .ZN(G9) );
NAND4_X1 U733 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
NOR3_X1 U734 ( .A1(n1015), .A2(KEYINPUT22), .A3(n1016), .ZN(n1014) );
INV_X1 U735 ( .A(n1017), .ZN(n1016) );
XNOR2_X1 U736 ( .A(n1018), .B(KEYINPUT7), .ZN(n1013) );
NOR2_X1 U737 ( .A1(n1019), .A2(n1020), .ZN(G75) );
NOR4_X1 U738 ( .A1(G953), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1020) );
XOR2_X1 U739 ( .A(KEYINPUT38), .B(n1024), .Z(n1023) );
NOR4_X1 U740 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
NOR3_X1 U741 ( .A1(n1029), .A2(n1015), .A3(n1030), .ZN(n1028) );
NOR3_X1 U742 ( .A1(n1031), .A2(n1032), .A3(n1030), .ZN(n1027) );
NAND3_X1 U743 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1031) );
NAND2_X1 U744 ( .A1(n1036), .A2(n1037), .ZN(n1033) );
NAND3_X1 U745 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND2_X1 U746 ( .A1(n1041), .A2(n1042), .ZN(n1038) );
NAND2_X1 U747 ( .A1(n1011), .A2(n1012), .ZN(n1036) );
NOR2_X1 U748 ( .A1(n1043), .A2(n1032), .ZN(n1026) );
NOR2_X1 U749 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR3_X1 U750 ( .A1(n1046), .A2(n1047), .A3(n1029), .ZN(n1045) );
NOR4_X1 U751 ( .A1(n1048), .A2(n1039), .A3(n1030), .A4(n1049), .ZN(n1044) );
NAND3_X1 U752 ( .A1(n1035), .A2(n1034), .A3(n1012), .ZN(n1048) );
INV_X1 U753 ( .A(KEYINPUT16), .ZN(n1034) );
NOR2_X1 U754 ( .A1(n1050), .A2(n1029), .ZN(n1025) );
NAND3_X1 U755 ( .A1(n1040), .A2(n1012), .A3(n1051), .ZN(n1029) );
NOR3_X1 U756 ( .A1(n1052), .A2(KEYINPUT16), .A3(n1053), .ZN(n1051) );
NOR2_X1 U757 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
AND2_X1 U758 ( .A1(n1018), .A2(n1056), .ZN(n1055) );
NOR2_X1 U759 ( .A1(n1057), .A2(n1030), .ZN(n1054) );
INV_X1 U760 ( .A(n1058), .ZN(n1030) );
NOR3_X1 U761 ( .A1(n1021), .A2(G953), .A3(G952), .ZN(n1019) );
AND4_X1 U762 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1021) );
NOR4_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1049), .ZN(n1062) );
NOR3_X1 U764 ( .A1(n1053), .A2(n1066), .A3(n1067), .ZN(n1061) );
XNOR2_X1 U765 ( .A(n1068), .B(n1069), .ZN(n1059) );
NAND2_X1 U766 ( .A1(n1070), .A2(KEYINPUT12), .ZN(n1069) );
XOR2_X1 U767 ( .A(n1071), .B(KEYINPUT33), .Z(n1070) );
XOR2_X1 U768 ( .A(n1072), .B(n1073), .Z(G72) );
NOR2_X1 U769 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U771 ( .A1(KEYINPUT3), .A2(n1078), .ZN(n1072) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(n1078) );
NOR2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U774 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U775 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U776 ( .A1(KEYINPUT30), .A2(n1087), .ZN(n1086) );
NAND2_X1 U777 ( .A1(KEYINPUT24), .A2(n1088), .ZN(n1085) );
XOR2_X1 U778 ( .A(G137), .B(G134), .Z(n1088) );
XOR2_X1 U779 ( .A(n1089), .B(n1090), .Z(n1083) );
NOR2_X1 U780 ( .A1(G900), .A2(n1075), .ZN(n1081) );
NAND2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1079) );
XNOR2_X1 U782 ( .A(G953), .B(KEYINPUT10), .ZN(n1091) );
XOR2_X1 U783 ( .A(n1093), .B(n1094), .Z(G69) );
NOR3_X1 U784 ( .A1(n1095), .A2(KEYINPUT41), .A3(n1096), .ZN(n1094) );
NOR2_X1 U785 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1099), .B(KEYINPUT53), .Z(n1095) );
NAND2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1099) );
NAND2_X1 U788 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NAND2_X1 U789 ( .A1(G953), .A2(n1102), .ZN(n1101) );
XNOR2_X1 U790 ( .A(n1103), .B(n1104), .ZN(n1100) );
NOR2_X1 U791 ( .A1(KEYINPUT60), .A2(n1105), .ZN(n1104) );
XNOR2_X1 U792 ( .A(n1106), .B(n1107), .ZN(n1105) );
AND2_X1 U793 ( .A1(n1075), .A2(n1108), .ZN(n1097) );
NAND2_X1 U794 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U795 ( .A1(G953), .A2(n1111), .ZN(n1093) );
NAND2_X1 U796 ( .A1(G898), .A2(G224), .ZN(n1111) );
NOR2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(G66) );
NOR3_X1 U798 ( .A1(n1068), .A2(n1114), .A3(n1115), .ZN(n1113) );
NOR3_X1 U799 ( .A1(n1116), .A2(n1071), .A3(n1117), .ZN(n1115) );
NOR2_X1 U800 ( .A1(n1118), .A2(n1119), .ZN(n1114) );
NOR2_X1 U801 ( .A1(n1120), .A2(n1071), .ZN(n1118) );
NOR2_X1 U802 ( .A1(n1112), .A2(n1121), .ZN(G63) );
XOR2_X1 U803 ( .A(n1122), .B(n1123), .Z(n1121) );
AND2_X1 U804 ( .A1(G478), .A2(n1124), .ZN(n1123) );
NOR2_X1 U805 ( .A1(n1112), .A2(n1125), .ZN(G60) );
NOR2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U807 ( .A(n1128), .B(KEYINPUT34), .Z(n1127) );
NAND2_X1 U808 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U809 ( .A1(n1124), .A2(G475), .ZN(n1130) );
XNOR2_X1 U810 ( .A(KEYINPUT37), .B(n1131), .ZN(n1129) );
NOR3_X1 U811 ( .A1(n1117), .A2(n1131), .A3(n1132), .ZN(n1126) );
XNOR2_X1 U812 ( .A(G104), .B(n1133), .ZN(G6) );
NAND2_X1 U813 ( .A1(KEYINPUT17), .A2(n1134), .ZN(n1133) );
NOR2_X1 U814 ( .A1(n1112), .A2(n1135), .ZN(G57) );
XOR2_X1 U815 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U816 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U817 ( .A1(n1140), .A2(KEYINPUT55), .ZN(n1139) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
XOR2_X1 U819 ( .A(n1143), .B(KEYINPUT5), .Z(n1142) );
NOR2_X1 U820 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
AND2_X1 U821 ( .A1(G472), .A2(n1124), .ZN(n1138) );
NOR3_X1 U822 ( .A1(n1112), .A2(n1146), .A3(n1147), .ZN(G54) );
NOR2_X1 U823 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U824 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U825 ( .A1(KEYINPUT58), .A2(n1152), .ZN(n1150) );
NOR2_X1 U826 ( .A1(n1153), .A2(n1154), .ZN(n1146) );
XOR2_X1 U827 ( .A(n1155), .B(n1151), .Z(n1154) );
XOR2_X1 U828 ( .A(n1156), .B(n1157), .Z(n1151) );
AND2_X1 U829 ( .A1(G469), .A2(n1124), .ZN(n1157) );
NAND2_X1 U830 ( .A1(n1158), .A2(KEYINPUT58), .ZN(n1155) );
INV_X1 U831 ( .A(n1152), .ZN(n1158) );
XNOR2_X1 U832 ( .A(n1089), .B(n1159), .ZN(n1152) );
NOR2_X1 U833 ( .A1(KEYINPUT6), .A2(n1160), .ZN(n1159) );
NOR2_X1 U834 ( .A1(n1112), .A2(n1161), .ZN(G51) );
XOR2_X1 U835 ( .A(n1162), .B(n1163), .Z(n1161) );
NOR2_X1 U836 ( .A1(n1164), .A2(n1117), .ZN(n1163) );
INV_X1 U837 ( .A(n1124), .ZN(n1117) );
NOR2_X1 U838 ( .A1(n1165), .A2(n1120), .ZN(n1124) );
INV_X1 U839 ( .A(n1022), .ZN(n1120) );
NAND3_X1 U840 ( .A1(n1166), .A2(n1109), .A3(n1167), .ZN(n1022) );
XOR2_X1 U841 ( .A(n1110), .B(KEYINPUT63), .Z(n1167) );
NAND3_X1 U842 ( .A1(n1012), .A2(n1168), .A3(n1169), .ZN(n1110) );
AND4_X1 U843 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1109) );
NOR4_X1 U844 ( .A1(n1174), .A2(n1175), .A3(n1134), .A4(n1176), .ZN(n1173) );
AND3_X1 U845 ( .A1(n1177), .A2(n1012), .A3(n1169), .ZN(n1134) );
INV_X1 U846 ( .A(n1178), .ZN(n1169) );
NOR2_X1 U847 ( .A1(n1179), .A2(n1180), .ZN(n1172) );
AND4_X1 U848 ( .A1(KEYINPUT47), .A2(n1181), .A3(n1182), .A4(n1012), .ZN(n1180) );
NAND2_X1 U849 ( .A1(n1183), .A2(n1063), .ZN(n1182) );
NOR2_X1 U850 ( .A1(KEYINPUT47), .A2(n1184), .ZN(n1179) );
NAND4_X1 U851 ( .A1(n1185), .A2(n1186), .A3(n1187), .A4(n1017), .ZN(n1170) );
XOR2_X1 U852 ( .A(KEYINPUT8), .B(n1011), .Z(n1187) );
XNOR2_X1 U853 ( .A(n1058), .B(KEYINPUT29), .ZN(n1185) );
INV_X1 U854 ( .A(n1092), .ZN(n1166) );
NAND2_X1 U855 ( .A1(n1188), .A2(n1189), .ZN(n1092) );
NOR4_X1 U856 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
INV_X1 U857 ( .A(n1194), .ZN(n1193) );
NOR4_X1 U858 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1188) );
NOR2_X1 U859 ( .A1(n1057), .A2(n1199), .ZN(n1198) );
NOR3_X1 U860 ( .A1(n1041), .A2(n1015), .A3(n1200), .ZN(n1197) );
NOR2_X1 U861 ( .A1(n1201), .A2(n1202), .ZN(n1162) );
XOR2_X1 U862 ( .A(n1203), .B(KEYINPUT19), .Z(n1202) );
NAND2_X1 U863 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NOR2_X1 U864 ( .A1(n1205), .A2(n1204), .ZN(n1201) );
XOR2_X1 U865 ( .A(n1206), .B(n1207), .Z(n1204) );
XOR2_X1 U866 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U867 ( .A1(KEYINPUT51), .A2(G125), .ZN(n1208) );
NOR2_X1 U868 ( .A1(n1075), .A2(G952), .ZN(n1112) );
XNOR2_X1 U869 ( .A(G146), .B(n1210), .ZN(G48) );
NAND3_X1 U870 ( .A1(n1211), .A2(n1177), .A3(KEYINPUT50), .ZN(n1210) );
INV_X1 U871 ( .A(n1199), .ZN(n1211) );
XOR2_X1 U872 ( .A(G143), .B(n1196), .Z(G45) );
AND4_X1 U873 ( .A1(n1011), .A2(n1018), .A3(n1212), .A4(n1213), .ZN(n1196) );
AND3_X1 U874 ( .A1(n1063), .A2(n1214), .A3(n1183), .ZN(n1213) );
XOR2_X1 U875 ( .A(G140), .B(n1192), .Z(G42) );
NOR3_X1 U876 ( .A1(n1057), .A2(n1200), .A3(n1042), .ZN(n1192) );
XOR2_X1 U877 ( .A(G137), .B(n1191), .Z(G39) );
AND2_X1 U878 ( .A1(n1186), .A2(n1215), .ZN(n1191) );
XNOR2_X1 U879 ( .A(G134), .B(n1216), .ZN(G36) );
NAND4_X1 U880 ( .A1(KEYINPUT18), .A2(n1212), .A3(n1215), .A4(n1168), .ZN(n1216) );
INV_X1 U881 ( .A(n1015), .ZN(n1168) );
INV_X1 U882 ( .A(n1200), .ZN(n1215) );
XOR2_X1 U883 ( .A(G131), .B(n1190), .Z(G33) );
NOR3_X1 U884 ( .A1(n1057), .A2(n1200), .A3(n1041), .ZN(n1190) );
NAND4_X1 U885 ( .A1(n1040), .A2(n1018), .A3(n1039), .A4(n1214), .ZN(n1200) );
XNOR2_X1 U886 ( .A(n1049), .B(KEYINPUT46), .ZN(n1040) );
XOR2_X1 U887 ( .A(G128), .B(n1195), .Z(G30) );
NOR2_X1 U888 ( .A1(n1199), .A2(n1015), .ZN(n1195) );
NAND3_X1 U889 ( .A1(n1018), .A2(n1064), .A3(n1217), .ZN(n1199) );
XOR2_X1 U890 ( .A(n1218), .B(G101), .Z(G3) );
NAND2_X1 U891 ( .A1(KEYINPUT31), .A2(n1219), .ZN(n1218) );
INV_X1 U892 ( .A(n1176), .ZN(n1219) );
NOR3_X1 U893 ( .A1(n1032), .A2(n1041), .A3(n1178), .ZN(n1176) );
XNOR2_X1 U894 ( .A(G125), .B(n1194), .ZN(G27) );
NAND4_X1 U895 ( .A1(n1058), .A2(n1217), .A3(n1220), .A4(n1177), .ZN(n1194) );
AND3_X1 U896 ( .A1(n1221), .A2(n1214), .A3(n1011), .ZN(n1217) );
NAND2_X1 U897 ( .A1(n1222), .A2(n1223), .ZN(n1214) );
NAND4_X1 U898 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1077), .ZN(n1222) );
INV_X1 U899 ( .A(G900), .ZN(n1077) );
XNOR2_X1 U900 ( .A(G122), .B(n1184), .ZN(G24) );
NAND4_X1 U901 ( .A1(n1181), .A2(n1012), .A3(n1063), .A4(n1183), .ZN(n1184) );
NOR2_X1 U902 ( .A1(n1064), .A2(n1221), .ZN(n1012) );
XNOR2_X1 U903 ( .A(G119), .B(n1225), .ZN(G21) );
NAND2_X1 U904 ( .A1(n1181), .A2(n1186), .ZN(n1225) );
AND3_X1 U905 ( .A1(n1221), .A2(n1064), .A3(n1056), .ZN(n1186) );
XOR2_X1 U906 ( .A(G116), .B(n1175), .Z(G18) );
NOR3_X1 U907 ( .A1(n1041), .A2(n1015), .A3(n1226), .ZN(n1175) );
NAND2_X1 U908 ( .A1(n1227), .A2(n1183), .ZN(n1015) );
XNOR2_X1 U909 ( .A(n1063), .B(KEYINPUT15), .ZN(n1227) );
INV_X1 U910 ( .A(n1212), .ZN(n1041) );
XNOR2_X1 U911 ( .A(G113), .B(n1171), .ZN(G15) );
NAND3_X1 U912 ( .A1(n1212), .A2(n1177), .A3(n1181), .ZN(n1171) );
INV_X1 U913 ( .A(n1226), .ZN(n1181) );
NAND3_X1 U914 ( .A1(n1011), .A2(n1017), .A3(n1058), .ZN(n1226) );
NOR2_X1 U915 ( .A1(n1047), .A2(n1067), .ZN(n1058) );
INV_X1 U916 ( .A(n1046), .ZN(n1067) );
INV_X1 U917 ( .A(n1057), .ZN(n1177) );
NAND2_X1 U918 ( .A1(n1228), .A2(n1063), .ZN(n1057) );
XNOR2_X1 U919 ( .A(KEYINPUT9), .B(n1183), .ZN(n1228) );
NOR2_X1 U920 ( .A1(n1221), .A2(n1220), .ZN(n1212) );
NAND2_X1 U921 ( .A1(n1229), .A2(n1230), .ZN(G12) );
NAND2_X1 U922 ( .A1(n1174), .A2(n1231), .ZN(n1230) );
XOR2_X1 U923 ( .A(KEYINPUT57), .B(n1232), .Z(n1229) );
NOR2_X1 U924 ( .A1(n1174), .A2(n1231), .ZN(n1232) );
NOR3_X1 U925 ( .A1(n1042), .A2(n1032), .A3(n1178), .ZN(n1174) );
NAND3_X1 U926 ( .A1(n1018), .A2(n1017), .A3(n1011), .ZN(n1178) );
NOR2_X1 U927 ( .A1(n1233), .A2(n1053), .ZN(n1011) );
INV_X1 U928 ( .A(n1039), .ZN(n1053) );
NAND2_X1 U929 ( .A1(G214), .A2(n1234), .ZN(n1039) );
INV_X1 U930 ( .A(n1049), .ZN(n1233) );
XOR2_X1 U931 ( .A(n1235), .B(n1164), .Z(n1049) );
NAND2_X1 U932 ( .A1(G210), .A2(n1234), .ZN(n1164) );
NAND2_X1 U933 ( .A1(n1236), .A2(n1165), .ZN(n1234) );
NAND2_X1 U934 ( .A1(n1237), .A2(n1165), .ZN(n1235) );
XOR2_X1 U935 ( .A(n1238), .B(n1239), .Z(n1237) );
XOR2_X1 U936 ( .A(KEYINPUT1), .B(n1240), .Z(n1239) );
NOR2_X1 U937 ( .A1(KEYINPUT26), .A2(n1241), .ZN(n1240) );
XNOR2_X1 U938 ( .A(n1206), .B(n1087), .ZN(n1241) );
XOR2_X1 U939 ( .A(n1242), .B(n1209), .Z(n1238) );
AND2_X1 U940 ( .A1(G224), .A2(n1075), .ZN(n1209) );
NAND2_X1 U941 ( .A1(KEYINPUT39), .A2(n1243), .ZN(n1242) );
INV_X1 U942 ( .A(n1205), .ZN(n1243) );
XOR2_X1 U943 ( .A(n1244), .B(n1245), .Z(n1205) );
INV_X1 U944 ( .A(n1103), .ZN(n1245) );
XNOR2_X1 U945 ( .A(n1246), .B(n1247), .ZN(n1103) );
XNOR2_X1 U946 ( .A(G122), .B(KEYINPUT52), .ZN(n1246) );
XNOR2_X1 U947 ( .A(n1248), .B(n1107), .ZN(n1244) );
INV_X1 U948 ( .A(n1160), .ZN(n1107) );
NAND2_X1 U949 ( .A1(KEYINPUT11), .A2(n1106), .ZN(n1248) );
XNOR2_X1 U950 ( .A(n1249), .B(n1250), .ZN(n1106) );
XNOR2_X1 U951 ( .A(G113), .B(KEYINPUT32), .ZN(n1249) );
NAND2_X1 U952 ( .A1(n1223), .A2(n1251), .ZN(n1017) );
NAND4_X1 U953 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1102), .ZN(n1251) );
INV_X1 U954 ( .A(G898), .ZN(n1102) );
NAND2_X1 U955 ( .A1(n1035), .A2(n1075), .ZN(n1223) );
INV_X1 U956 ( .A(n1052), .ZN(n1035) );
NAND2_X1 U957 ( .A1(n1252), .A2(n1224), .ZN(n1052) );
NAND2_X1 U958 ( .A1(G237), .A2(G234), .ZN(n1224) );
XNOR2_X1 U959 ( .A(G952), .B(KEYINPUT28), .ZN(n1252) );
AND2_X1 U960 ( .A1(n1047), .A2(n1046), .ZN(n1018) );
NAND2_X1 U961 ( .A1(G221), .A2(n1253), .ZN(n1046) );
XNOR2_X1 U962 ( .A(n1065), .B(KEYINPUT45), .ZN(n1047) );
XOR2_X1 U963 ( .A(G469), .B(n1254), .Z(n1065) );
NOR2_X1 U964 ( .A1(G902), .A2(n1255), .ZN(n1254) );
NOR2_X1 U965 ( .A1(n1256), .A2(n1257), .ZN(n1255) );
XOR2_X1 U966 ( .A(KEYINPUT61), .B(n1258), .Z(n1257) );
NOR2_X1 U967 ( .A1(n1156), .A2(n1259), .ZN(n1258) );
AND2_X1 U968 ( .A1(n1259), .A2(n1156), .ZN(n1256) );
XOR2_X1 U969 ( .A(n1260), .B(n1261), .Z(n1156) );
NOR2_X1 U970 ( .A1(G953), .A2(n1076), .ZN(n1261) );
INV_X1 U971 ( .A(G227), .ZN(n1076) );
NAND2_X1 U972 ( .A1(n1262), .A2(n1263), .ZN(n1259) );
OR2_X1 U973 ( .A1(n1264), .A2(n1148), .ZN(n1263) );
XOR2_X1 U974 ( .A(n1265), .B(KEYINPUT0), .Z(n1262) );
NAND2_X1 U975 ( .A1(n1266), .A2(n1264), .ZN(n1265) );
XOR2_X1 U976 ( .A(n1160), .B(n1267), .Z(n1264) );
NOR2_X1 U977 ( .A1(KEYINPUT56), .A2(n1089), .ZN(n1267) );
XNOR2_X1 U978 ( .A(G146), .B(n1268), .ZN(n1089) );
XNOR2_X1 U979 ( .A(n1269), .B(n1270), .ZN(n1160) );
XOR2_X1 U980 ( .A(KEYINPUT42), .B(G107), .Z(n1270) );
XNOR2_X1 U981 ( .A(G101), .B(G104), .ZN(n1269) );
XNOR2_X1 U982 ( .A(n1153), .B(KEYINPUT40), .ZN(n1266) );
INV_X1 U983 ( .A(n1056), .ZN(n1032) );
NOR2_X1 U984 ( .A1(n1183), .A2(n1063), .ZN(n1056) );
XOR2_X1 U985 ( .A(n1271), .B(n1132), .Z(n1063) );
INV_X1 U986 ( .A(G475), .ZN(n1132) );
NAND2_X1 U987 ( .A1(n1131), .A2(n1165), .ZN(n1271) );
XOR2_X1 U988 ( .A(n1272), .B(n1273), .Z(n1131) );
XNOR2_X1 U989 ( .A(n1274), .B(G113), .ZN(n1273) );
XNOR2_X1 U990 ( .A(n1275), .B(n1276), .ZN(n1272) );
INV_X1 U991 ( .A(G104), .ZN(n1276) );
NAND2_X1 U992 ( .A1(n1277), .A2(KEYINPUT27), .ZN(n1275) );
XOR2_X1 U993 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U994 ( .A(G143), .B(n1280), .Z(n1279) );
AND3_X1 U995 ( .A1(n1281), .A2(n1075), .A3(G214), .ZN(n1280) );
XNOR2_X1 U996 ( .A(n1090), .B(n1282), .ZN(n1278) );
XOR2_X1 U997 ( .A(G131), .B(G140), .Z(n1090) );
NAND2_X1 U998 ( .A1(n1283), .A2(n1060), .ZN(n1183) );
NAND2_X1 U999 ( .A1(n1284), .A2(n1285), .ZN(n1060) );
XNOR2_X1 U1000 ( .A(n1066), .B(KEYINPUT36), .ZN(n1283) );
NOR2_X1 U1001 ( .A1(n1285), .A2(n1284), .ZN(n1066) );
NOR2_X1 U1002 ( .A1(n1122), .A2(G902), .ZN(n1284) );
XOR2_X1 U1003 ( .A(n1286), .B(n1287), .Z(n1122) );
XNOR2_X1 U1004 ( .A(n1288), .B(n1268), .ZN(n1287) );
NAND2_X1 U1005 ( .A1(KEYINPUT4), .A2(n1289), .ZN(n1288) );
XOR2_X1 U1006 ( .A(G107), .B(n1290), .Z(n1289) );
XNOR2_X1 U1007 ( .A(n1274), .B(G116), .ZN(n1290) );
INV_X1 U1008 ( .A(G122), .ZN(n1274) );
XOR2_X1 U1009 ( .A(n1291), .B(G134), .Z(n1286) );
NAND3_X1 U1010 ( .A1(G234), .A2(n1292), .A3(G217), .ZN(n1291) );
XNOR2_X1 U1011 ( .A(KEYINPUT25), .B(n1075), .ZN(n1292) );
XOR2_X1 U1012 ( .A(G478), .B(KEYINPUT59), .Z(n1285) );
NAND2_X1 U1013 ( .A1(n1220), .A2(n1221), .ZN(n1042) );
XNOR2_X1 U1014 ( .A(n1068), .B(n1071), .ZN(n1221) );
NAND2_X1 U1015 ( .A1(G217), .A2(n1253), .ZN(n1071) );
NAND2_X1 U1016 ( .A1(G234), .A2(n1165), .ZN(n1253) );
NOR2_X1 U1017 ( .A1(n1119), .A2(G902), .ZN(n1068) );
INV_X1 U1018 ( .A(n1116), .ZN(n1119) );
XNOR2_X1 U1019 ( .A(n1293), .B(n1294), .ZN(n1116) );
XOR2_X1 U1020 ( .A(n1295), .B(n1296), .Z(n1294) );
XOR2_X1 U1021 ( .A(G137), .B(G119), .Z(n1296) );
XOR2_X1 U1022 ( .A(KEYINPUT54), .B(KEYINPUT21), .Z(n1295) );
XOR2_X1 U1023 ( .A(n1297), .B(n1298), .Z(n1293) );
XOR2_X1 U1024 ( .A(n1299), .B(n1300), .Z(n1298) );
AND3_X1 U1025 ( .A1(G221), .A2(n1075), .A3(G234), .ZN(n1300) );
NOR2_X1 U1026 ( .A1(KEYINPUT49), .A2(G128), .ZN(n1299) );
XOR2_X1 U1027 ( .A(n1260), .B(n1282), .Z(n1297) );
XNOR2_X1 U1028 ( .A(n1087), .B(G146), .ZN(n1282) );
INV_X1 U1029 ( .A(G125), .ZN(n1087) );
XNOR2_X1 U1030 ( .A(G140), .B(n1247), .ZN(n1260) );
XNOR2_X1 U1031 ( .A(n1231), .B(KEYINPUT14), .ZN(n1247) );
INV_X1 U1032 ( .A(G110), .ZN(n1231) );
INV_X1 U1033 ( .A(n1064), .ZN(n1220) );
XNOR2_X1 U1034 ( .A(n1301), .B(G472), .ZN(n1064) );
NAND2_X1 U1035 ( .A1(n1302), .A2(n1165), .ZN(n1301) );
INV_X1 U1036 ( .A(G902), .ZN(n1165) );
XNOR2_X1 U1037 ( .A(n1303), .B(n1136), .ZN(n1302) );
XNOR2_X1 U1038 ( .A(n1304), .B(G101), .ZN(n1136) );
NAND3_X1 U1039 ( .A1(G210), .A2(n1075), .A3(n1281), .ZN(n1304) );
XOR2_X1 U1040 ( .A(n1236), .B(KEYINPUT35), .Z(n1281) );
INV_X1 U1041 ( .A(G237), .ZN(n1236) );
INV_X1 U1042 ( .A(G953), .ZN(n1075) );
NAND2_X1 U1043 ( .A1(n1305), .A2(n1306), .ZN(n1303) );
NAND2_X1 U1044 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
INV_X1 U1045 ( .A(n1145), .ZN(n1308) );
XOR2_X1 U1046 ( .A(KEYINPUT23), .B(n1144), .Z(n1307) );
XNOR2_X1 U1047 ( .A(KEYINPUT2), .B(n1143), .ZN(n1305) );
NAND2_X1 U1048 ( .A1(n1145), .A2(n1144), .ZN(n1143) );
AND3_X1 U1049 ( .A1(n1309), .A2(n1310), .A3(n1311), .ZN(n1144) );
NAND2_X1 U1050 ( .A1(n1250), .A2(n1312), .ZN(n1311) );
INV_X1 U1051 ( .A(G113), .ZN(n1312) );
NAND2_X1 U1052 ( .A1(KEYINPUT20), .A2(n1313), .ZN(n1310) );
NAND2_X1 U1053 ( .A1(n1314), .A2(G113), .ZN(n1313) );
XNOR2_X1 U1054 ( .A(KEYINPUT43), .B(n1315), .ZN(n1314) );
NAND2_X1 U1055 ( .A1(n1316), .A2(n1317), .ZN(n1309) );
INV_X1 U1056 ( .A(KEYINPUT20), .ZN(n1317) );
NAND2_X1 U1057 ( .A1(n1318), .A2(n1319), .ZN(n1316) );
OR2_X1 U1058 ( .A1(n1315), .A2(KEYINPUT43), .ZN(n1319) );
NAND3_X1 U1059 ( .A1(G113), .A2(n1315), .A3(KEYINPUT43), .ZN(n1318) );
INV_X1 U1060 ( .A(n1250), .ZN(n1315) );
XNOR2_X1 U1061 ( .A(G116), .B(G119), .ZN(n1250) );
XNOR2_X1 U1062 ( .A(n1206), .B(n1320), .ZN(n1145) );
XNOR2_X1 U1063 ( .A(KEYINPUT62), .B(n1148), .ZN(n1320) );
INV_X1 U1064 ( .A(n1153), .ZN(n1148) );
XOR2_X1 U1065 ( .A(G131), .B(n1321), .Z(n1153) );
NOR2_X1 U1066 ( .A1(KEYINPUT44), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1067 ( .A(n1323), .B(G137), .Z(n1322) );
NAND2_X1 U1068 ( .A1(KEYINPUT13), .A2(G134), .ZN(n1323) );
NAND2_X1 U1069 ( .A1(n1324), .A2(n1325), .ZN(n1206) );
NAND2_X1 U1070 ( .A1(n1326), .A2(n1327), .ZN(n1325) );
INV_X1 U1071 ( .A(G146), .ZN(n1327) );
XOR2_X1 U1072 ( .A(KEYINPUT48), .B(n1268), .Z(n1326) );
NAND2_X1 U1073 ( .A1(n1268), .A2(G146), .ZN(n1324) );
XOR2_X1 U1074 ( .A(G128), .B(G143), .Z(n1268) );
endmodule


