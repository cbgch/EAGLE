//Key = 0101000110110111000111101011101000110000010111101110001110110100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;

XNOR2_X1 U670 ( .A(G107), .B(n919), .ZN(G9) );
NOR2_X1 U671 ( .A1(n920), .A2(n921), .ZN(G75) );
NOR3_X1 U672 ( .A1(n922), .A2(G953), .A3(n923), .ZN(n921) );
NAND3_X1 U673 ( .A1(n924), .A2(n925), .A3(n926), .ZN(n922) );
NAND2_X1 U674 ( .A1(n927), .A2(n928), .ZN(n925) );
NAND2_X1 U675 ( .A1(n929), .A2(n930), .ZN(n927) );
NAND3_X1 U676 ( .A1(n931), .A2(n932), .A3(n933), .ZN(n930) );
NAND2_X1 U677 ( .A1(n934), .A2(n935), .ZN(n932) );
NAND3_X1 U678 ( .A1(n936), .A2(n937), .A3(n938), .ZN(n935) );
NAND2_X1 U679 ( .A1(n939), .A2(n940), .ZN(n937) );
OR2_X1 U680 ( .A1(n941), .A2(KEYINPUT58), .ZN(n939) );
NAND3_X1 U681 ( .A1(n942), .A2(n943), .A3(n944), .ZN(n936) );
NAND2_X1 U682 ( .A1(KEYINPUT58), .A2(n945), .ZN(n942) );
NAND3_X1 U683 ( .A1(n946), .A2(n947), .A3(n948), .ZN(n934) );
NAND2_X1 U684 ( .A1(n949), .A2(n940), .ZN(n947) );
NAND2_X1 U685 ( .A1(n938), .A2(n950), .ZN(n949) );
NAND2_X1 U686 ( .A1(n951), .A2(n952), .ZN(n950) );
OR3_X1 U687 ( .A1(n953), .A2(n954), .A3(n940), .ZN(n946) );
NAND2_X1 U688 ( .A1(n955), .A2(n956), .ZN(n929) );
NAND3_X1 U689 ( .A1(n957), .A2(n933), .A3(n958), .ZN(n924) );
XNOR2_X1 U690 ( .A(n955), .B(KEYINPUT34), .ZN(n957) );
AND4_X1 U691 ( .A1(n931), .A2(n944), .A3(n948), .A4(n938), .ZN(n955) );
INV_X1 U692 ( .A(n959), .ZN(n931) );
NOR3_X1 U693 ( .A1(n923), .A2(G953), .A3(G952), .ZN(n920) );
AND4_X1 U694 ( .A1(n960), .A2(n961), .A3(n962), .A4(n963), .ZN(n923) );
AND2_X1 U695 ( .A1(n948), .A2(n964), .ZN(n963) );
XOR2_X1 U696 ( .A(KEYINPUT30), .B(n965), .Z(n961) );
XOR2_X1 U697 ( .A(KEYINPUT37), .B(n966), .Z(n960) );
NOR2_X1 U698 ( .A1(n967), .A2(n968), .ZN(n966) );
INV_X1 U699 ( .A(n969), .ZN(n967) );
XOR2_X1 U700 ( .A(n970), .B(n971), .Z(G72) );
NOR2_X1 U701 ( .A1(KEYINPUT31), .A2(n972), .ZN(n971) );
XOR2_X1 U702 ( .A(n973), .B(n974), .Z(n972) );
NAND3_X1 U703 ( .A1(n975), .A2(n976), .A3(KEYINPUT26), .ZN(n974) );
NAND2_X1 U704 ( .A1(n977), .A2(n978), .ZN(n973) );
NAND2_X1 U705 ( .A1(G953), .A2(n979), .ZN(n978) );
XOR2_X1 U706 ( .A(n980), .B(n981), .Z(n977) );
XOR2_X1 U707 ( .A(n982), .B(n983), .Z(n981) );
NAND2_X1 U708 ( .A1(n984), .A2(n985), .ZN(n982) );
XNOR2_X1 U709 ( .A(n986), .B(KEYINPUT16), .ZN(n984) );
XOR2_X1 U710 ( .A(n987), .B(n988), .Z(n980) );
XOR2_X1 U711 ( .A(KEYINPUT53), .B(KEYINPUT45), .Z(n988) );
NAND2_X1 U712 ( .A1(KEYINPUT50), .A2(n989), .ZN(n987) );
NAND2_X1 U713 ( .A1(n990), .A2(n991), .ZN(n970) );
NAND2_X1 U714 ( .A1(G900), .A2(G227), .ZN(n991) );
INV_X1 U715 ( .A(n992), .ZN(n990) );
XOR2_X1 U716 ( .A(n993), .B(n994), .Z(G69) );
XOR2_X1 U717 ( .A(n995), .B(n996), .Z(n994) );
NOR2_X1 U718 ( .A1(n997), .A2(n992), .ZN(n996) );
XOR2_X1 U719 ( .A(G953), .B(KEYINPUT24), .Z(n992) );
AND2_X1 U720 ( .A1(G224), .A2(G898), .ZN(n997) );
NAND2_X1 U721 ( .A1(n998), .A2(n999), .ZN(n995) );
NAND2_X1 U722 ( .A1(G953), .A2(n1000), .ZN(n999) );
XNOR2_X1 U723 ( .A(n1001), .B(n1002), .ZN(n998) );
XOR2_X1 U724 ( .A(n1003), .B(KEYINPUT25), .Z(n1001) );
NAND2_X1 U725 ( .A1(n976), .A2(n1004), .ZN(n993) );
NOR3_X1 U726 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(G66) );
AND3_X1 U727 ( .A1(KEYINPUT6), .A2(n1008), .A3(n1009), .ZN(n1007) );
NOR2_X1 U728 ( .A1(KEYINPUT6), .A2(n1010), .ZN(n1006) );
XOR2_X1 U729 ( .A(n1011), .B(n1012), .Z(n1005) );
NAND2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR2_X1 U731 ( .A1(n1015), .A2(n1016), .ZN(G63) );
XOR2_X1 U732 ( .A(n1017), .B(n1018), .Z(n1016) );
NAND2_X1 U733 ( .A1(n1013), .A2(G478), .ZN(n1017) );
NOR3_X1 U734 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(G60) );
NOR3_X1 U735 ( .A1(n1022), .A2(n1009), .A3(n1008), .ZN(n1021) );
INV_X1 U736 ( .A(G952), .ZN(n1008) );
INV_X1 U737 ( .A(KEYINPUT9), .ZN(n1022) );
NOR2_X1 U738 ( .A1(KEYINPUT9), .A2(n1010), .ZN(n1020) );
INV_X1 U739 ( .A(n1015), .ZN(n1010) );
XOR2_X1 U740 ( .A(n1023), .B(n1024), .Z(n1019) );
NAND2_X1 U741 ( .A1(n1013), .A2(G475), .ZN(n1023) );
XOR2_X1 U742 ( .A(n1025), .B(n1026), .Z(G6) );
XNOR2_X1 U743 ( .A(G104), .B(KEYINPUT4), .ZN(n1026) );
NOR2_X1 U744 ( .A1(n1015), .A2(n1027), .ZN(G57) );
XOR2_X1 U745 ( .A(n1028), .B(n1029), .Z(n1027) );
XNOR2_X1 U746 ( .A(n1030), .B(n1031), .ZN(n1029) );
NOR2_X1 U747 ( .A1(KEYINPUT40), .A2(n1032), .ZN(n1031) );
NAND2_X1 U748 ( .A1(KEYINPUT56), .A2(n1033), .ZN(n1030) );
XOR2_X1 U749 ( .A(n1034), .B(n1035), .Z(n1028) );
XNOR2_X1 U750 ( .A(n1036), .B(KEYINPUT27), .ZN(n1035) );
NAND2_X1 U751 ( .A1(n1013), .A2(G472), .ZN(n1034) );
NOR2_X1 U752 ( .A1(n1015), .A2(n1037), .ZN(G54) );
NOR2_X1 U753 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
XOR2_X1 U754 ( .A(n1040), .B(n1041), .Z(n1039) );
NAND2_X1 U755 ( .A1(KEYINPUT13), .A2(n1042), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1013), .A2(G469), .ZN(n1040) );
NOR2_X1 U757 ( .A1(KEYINPUT13), .A2(n1042), .ZN(n1038) );
XOR2_X1 U758 ( .A(n1043), .B(n1044), .Z(n1042) );
XNOR2_X1 U759 ( .A(n1045), .B(KEYINPUT42), .ZN(n1044) );
NAND2_X1 U760 ( .A1(n1046), .A2(KEYINPUT59), .ZN(n1045) );
XNOR2_X1 U761 ( .A(n989), .B(n1047), .ZN(n1046) );
INV_X1 U762 ( .A(n1048), .ZN(n989) );
XNOR2_X1 U763 ( .A(n1049), .B(n1050), .ZN(n1043) );
NOR2_X1 U764 ( .A1(n1015), .A2(n1051), .ZN(G51) );
XOR2_X1 U765 ( .A(n1052), .B(n1053), .Z(n1051) );
XOR2_X1 U766 ( .A(n1054), .B(n1055), .Z(n1053) );
XOR2_X1 U767 ( .A(n1056), .B(n1057), .Z(n1052) );
NAND2_X1 U768 ( .A1(KEYINPUT7), .A2(n1058), .ZN(n1057) );
NAND2_X1 U769 ( .A1(n1013), .A2(n1059), .ZN(n1056) );
NOR2_X1 U770 ( .A1(n1060), .A2(n926), .ZN(n1013) );
NOR2_X1 U771 ( .A1(n975), .A2(n1004), .ZN(n926) );
NAND4_X1 U772 ( .A1(n1061), .A2(n1025), .A3(n1062), .A4(n1063), .ZN(n1004) );
AND4_X1 U773 ( .A1(n1064), .A2(n919), .A3(n1065), .A4(n1066), .ZN(n1063) );
NAND3_X1 U774 ( .A1(n938), .A2(n1067), .A3(n1068), .ZN(n919) );
NAND2_X1 U775 ( .A1(n1069), .A2(n1070), .ZN(n1062) );
NAND2_X1 U776 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND2_X1 U777 ( .A1(n1073), .A2(n945), .ZN(n1072) );
XNOR2_X1 U778 ( .A(KEYINPUT41), .B(n953), .ZN(n1073) );
NAND2_X1 U779 ( .A1(n1068), .A2(n953), .ZN(n1071) );
NAND3_X1 U780 ( .A1(n938), .A2(n1067), .A3(n945), .ZN(n1025) );
NAND3_X1 U781 ( .A1(n1067), .A2(n1074), .A3(n954), .ZN(n1061) );
XOR2_X1 U782 ( .A(KEYINPUT23), .B(n948), .Z(n1074) );
NAND2_X1 U783 ( .A1(n1075), .A2(n1076), .ZN(n975) );
AND4_X1 U784 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
AND4_X1 U785 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1075) );
NAND3_X1 U786 ( .A1(n1085), .A2(n953), .A3(n945), .ZN(n1084) );
NOR2_X1 U787 ( .A1(n1009), .A2(G952), .ZN(n1015) );
XOR2_X1 U788 ( .A(G953), .B(KEYINPUT11), .Z(n1009) );
XNOR2_X1 U789 ( .A(G146), .B(n1083), .ZN(G48) );
NAND3_X1 U790 ( .A1(n945), .A2(n1086), .A3(n1087), .ZN(n1083) );
XNOR2_X1 U791 ( .A(G143), .B(n1082), .ZN(G45) );
NAND4_X1 U792 ( .A1(n1087), .A2(n953), .A3(n1088), .A4(n1089), .ZN(n1082) );
XNOR2_X1 U793 ( .A(G140), .B(n1081), .ZN(G42) );
NAND3_X1 U794 ( .A1(n945), .A2(n954), .A3(n1085), .ZN(n1081) );
XNOR2_X1 U795 ( .A(G137), .B(n1080), .ZN(G39) );
NAND3_X1 U796 ( .A1(n948), .A2(n1086), .A3(n1085), .ZN(n1080) );
XOR2_X1 U797 ( .A(n1079), .B(n1090), .Z(G36) );
XNOR2_X1 U798 ( .A(G134), .B(KEYINPUT0), .ZN(n1090) );
NAND3_X1 U799 ( .A1(n1068), .A2(n953), .A3(n1085), .ZN(n1079) );
XNOR2_X1 U800 ( .A(n1091), .B(n1092), .ZN(G33) );
NAND2_X1 U801 ( .A1(KEYINPUT3), .A2(n1093), .ZN(n1091) );
NAND3_X1 U802 ( .A1(n1085), .A2(n953), .A3(n1094), .ZN(n1093) );
XNOR2_X1 U803 ( .A(n945), .B(KEYINPUT20), .ZN(n1094) );
AND3_X1 U804 ( .A1(n952), .A2(n1095), .A3(n964), .ZN(n1085) );
NOR3_X1 U805 ( .A1(n956), .A2(n951), .A3(n958), .ZN(n964) );
XNOR2_X1 U806 ( .A(G128), .B(n1078), .ZN(G30) );
NAND3_X1 U807 ( .A1(n1068), .A2(n1086), .A3(n1087), .ZN(n1078) );
AND2_X1 U808 ( .A1(n1096), .A2(n1095), .ZN(n1087) );
XNOR2_X1 U809 ( .A(G101), .B(n1097), .ZN(G3) );
NOR2_X1 U810 ( .A1(n1098), .A2(KEYINPUT32), .ZN(n1097) );
INV_X1 U811 ( .A(n1064), .ZN(n1098) );
NAND3_X1 U812 ( .A1(n1067), .A2(n953), .A3(n948), .ZN(n1064) );
XOR2_X1 U813 ( .A(n1077), .B(n1099), .Z(G27) );
NAND2_X1 U814 ( .A1(n1100), .A2(G125), .ZN(n1099) );
XNOR2_X1 U815 ( .A(KEYINPUT33), .B(KEYINPUT18), .ZN(n1100) );
NAND4_X1 U816 ( .A1(n945), .A2(n954), .A3(n1101), .A4(n1095), .ZN(n1077) );
NAND2_X1 U817 ( .A1(n959), .A2(n1102), .ZN(n1095) );
NAND2_X1 U818 ( .A1(n1103), .A2(n979), .ZN(n1102) );
INV_X1 U819 ( .A(G900), .ZN(n979) );
XNOR2_X1 U820 ( .A(G122), .B(n1066), .ZN(G24) );
NAND4_X1 U821 ( .A1(n1069), .A2(n938), .A3(n1088), .A4(n1089), .ZN(n1066) );
AND2_X1 U822 ( .A1(n962), .A2(n1104), .ZN(n938) );
XOR2_X1 U823 ( .A(KEYINPUT63), .B(n1105), .Z(n1104) );
XOR2_X1 U824 ( .A(G119), .B(n1106), .Z(G21) );
NOR2_X1 U825 ( .A1(KEYINPUT38), .A2(n1065), .ZN(n1106) );
NAND3_X1 U826 ( .A1(n948), .A2(n1086), .A3(n1069), .ZN(n1065) );
INV_X1 U827 ( .A(n1107), .ZN(n1069) );
XOR2_X1 U828 ( .A(G116), .B(n1108), .Z(G18) );
NOR4_X1 U829 ( .A1(KEYINPUT62), .A2(n1109), .A3(n943), .A4(n1107), .ZN(n1108) );
NAND2_X1 U830 ( .A1(n1101), .A2(n1110), .ZN(n1107) );
INV_X1 U831 ( .A(n1068), .ZN(n943) );
NOR2_X1 U832 ( .A1(n1089), .A2(n1111), .ZN(n1068) );
INV_X1 U833 ( .A(n953), .ZN(n1109) );
XNOR2_X1 U834 ( .A(G113), .B(n1112), .ZN(G15) );
NAND4_X1 U835 ( .A1(n945), .A2(n1101), .A3(n1113), .A4(n953), .ZN(n1112) );
NAND2_X1 U836 ( .A1(n1114), .A2(n1115), .ZN(n953) );
NAND2_X1 U837 ( .A1(n1086), .A2(n1116), .ZN(n1115) );
INV_X1 U838 ( .A(KEYINPUT10), .ZN(n1116) );
NAND2_X1 U839 ( .A1(n1117), .A2(n1118), .ZN(n1086) );
OR3_X1 U840 ( .A1(n962), .A2(n1105), .A3(KEYINPUT36), .ZN(n1118) );
NAND2_X1 U841 ( .A1(KEYINPUT36), .A2(n954), .ZN(n1117) );
NAND3_X1 U842 ( .A1(n1105), .A2(n1119), .A3(KEYINPUT10), .ZN(n1114) );
XNOR2_X1 U843 ( .A(KEYINPUT36), .B(n962), .ZN(n1119) );
INV_X1 U844 ( .A(n1120), .ZN(n962) );
XNOR2_X1 U845 ( .A(KEYINPUT19), .B(n1110), .ZN(n1113) );
NOR3_X1 U846 ( .A1(n928), .A2(n956), .A3(n940), .ZN(n1101) );
INV_X1 U847 ( .A(n944), .ZN(n940) );
NOR2_X1 U848 ( .A1(n952), .A2(n951), .ZN(n944) );
INV_X1 U849 ( .A(n1121), .ZN(n952) );
INV_X1 U850 ( .A(n941), .ZN(n945) );
NAND2_X1 U851 ( .A1(n1111), .A2(n1089), .ZN(n941) );
INV_X1 U852 ( .A(n1088), .ZN(n1111) );
XNOR2_X1 U853 ( .A(G110), .B(n1122), .ZN(G12) );
NAND3_X1 U854 ( .A1(n948), .A2(n1067), .A3(n954), .ZN(n1122) );
NOR2_X1 U855 ( .A1(n1120), .A2(n1105), .ZN(n954) );
AND2_X1 U856 ( .A1(n1123), .A2(n969), .ZN(n1105) );
NAND3_X1 U857 ( .A1(n1124), .A2(n1060), .A3(n1012), .ZN(n969) );
OR2_X1 U858 ( .A1(n1125), .A2(G234), .ZN(n1124) );
XOR2_X1 U859 ( .A(KEYINPUT46), .B(n968), .Z(n1123) );
AND2_X1 U860 ( .A1(n1014), .A2(n1126), .ZN(n968) );
NAND2_X1 U861 ( .A1(n1012), .A2(n1060), .ZN(n1126) );
XNOR2_X1 U862 ( .A(n1127), .B(n1128), .ZN(n1012) );
XOR2_X1 U863 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U864 ( .A1(G221), .A2(n1131), .ZN(n1130) );
INV_X1 U865 ( .A(n1132), .ZN(n1131) );
NAND2_X1 U866 ( .A1(KEYINPUT1), .A2(n1133), .ZN(n1129) );
XOR2_X1 U867 ( .A(G110), .B(n1134), .Z(n1133) );
XOR2_X1 U868 ( .A(G128), .B(G119), .Z(n1134) );
XOR2_X1 U869 ( .A(n1135), .B(n1136), .Z(n1127) );
NOR2_X1 U870 ( .A1(G137), .A2(KEYINPUT2), .ZN(n1136) );
XNOR2_X1 U871 ( .A(n1137), .B(n1138), .ZN(n1135) );
NAND3_X1 U872 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1137) );
XNOR2_X1 U873 ( .A(KEYINPUT28), .B(n985), .ZN(n1141) );
OR3_X1 U874 ( .A1(n1142), .A2(n1058), .A3(KEYINPUT44), .ZN(n1140) );
NAND2_X1 U875 ( .A1(n986), .A2(KEYINPUT44), .ZN(n1139) );
AND2_X1 U876 ( .A1(G217), .A2(n1143), .ZN(n1014) );
XNOR2_X1 U877 ( .A(n1144), .B(G472), .ZN(n1120) );
NAND2_X1 U878 ( .A1(n1145), .A2(n1060), .ZN(n1144) );
XOR2_X1 U879 ( .A(n1146), .B(n1147), .Z(n1145) );
XNOR2_X1 U880 ( .A(n1148), .B(n1032), .ZN(n1147) );
XOR2_X1 U881 ( .A(n1149), .B(n1150), .Z(n1032) );
XNOR2_X1 U882 ( .A(n1151), .B(n1152), .ZN(n1150) );
INV_X1 U883 ( .A(n1049), .ZN(n1152) );
XNOR2_X1 U884 ( .A(G113), .B(n1153), .ZN(n1149) );
NAND2_X1 U885 ( .A1(KEYINPUT49), .A2(n1036), .ZN(n1148) );
AND3_X1 U886 ( .A1(n1154), .A2(n976), .A3(G210), .ZN(n1036) );
XNOR2_X1 U887 ( .A(n1155), .B(n1033), .ZN(n1146) );
INV_X1 U888 ( .A(G101), .ZN(n1033) );
XNOR2_X1 U889 ( .A(KEYINPUT61), .B(KEYINPUT29), .ZN(n1155) );
AND2_X1 U890 ( .A1(n1096), .A2(n1110), .ZN(n1067) );
NAND2_X1 U891 ( .A1(n959), .A2(n1156), .ZN(n1110) );
NAND2_X1 U892 ( .A1(n1103), .A2(n1000), .ZN(n1156) );
INV_X1 U893 ( .A(G898), .ZN(n1000) );
AND3_X1 U894 ( .A1(n1157), .A2(n1158), .A3(G953), .ZN(n1103) );
XNOR2_X1 U895 ( .A(KEYINPUT60), .B(n1060), .ZN(n1157) );
NAND3_X1 U896 ( .A1(n1158), .A2(n976), .A3(G952), .ZN(n959) );
NAND2_X1 U897 ( .A1(G237), .A2(G234), .ZN(n1158) );
NOR4_X1 U898 ( .A1(n1121), .A2(n928), .A3(n956), .A4(n951), .ZN(n1096) );
AND2_X1 U899 ( .A1(G221), .A2(n1143), .ZN(n951) );
NAND2_X1 U900 ( .A1(G234), .A2(n1060), .ZN(n1143) );
INV_X1 U901 ( .A(n933), .ZN(n956) );
NAND2_X1 U902 ( .A1(G214), .A2(n1159), .ZN(n933) );
INV_X1 U903 ( .A(n958), .ZN(n928) );
XNOR2_X1 U904 ( .A(n1160), .B(n1059), .ZN(n958) );
AND2_X1 U905 ( .A1(G210), .A2(n1159), .ZN(n1059) );
NAND2_X1 U906 ( .A1(n1154), .A2(n1060), .ZN(n1159) );
NAND2_X1 U907 ( .A1(n1161), .A2(n1060), .ZN(n1160) );
XNOR2_X1 U908 ( .A(n1054), .B(n1162), .ZN(n1161) );
NOR2_X1 U909 ( .A1(KEYINPUT12), .A2(n1163), .ZN(n1162) );
XNOR2_X1 U910 ( .A(n1058), .B(n1055), .ZN(n1163) );
XNOR2_X1 U911 ( .A(n1164), .B(n1151), .ZN(n1055) );
XNOR2_X1 U912 ( .A(n1048), .B(KEYINPUT57), .ZN(n1151) );
NAND2_X1 U913 ( .A1(G224), .A2(n976), .ZN(n1164) );
XNOR2_X1 U914 ( .A(n1003), .B(n1165), .ZN(n1054) );
NOR2_X1 U915 ( .A1(KEYINPUT39), .A2(n1002), .ZN(n1165) );
XNOR2_X1 U916 ( .A(G110), .B(G122), .ZN(n1002) );
XOR2_X1 U917 ( .A(n1166), .B(n1047), .Z(n1003) );
XNOR2_X1 U918 ( .A(n1153), .B(n1167), .ZN(n1166) );
NOR2_X1 U919 ( .A1(G113), .A2(KEYINPUT47), .ZN(n1167) );
XOR2_X1 U920 ( .A(G116), .B(G119), .Z(n1153) );
XOR2_X1 U921 ( .A(n965), .B(KEYINPUT54), .Z(n1121) );
XNOR2_X1 U922 ( .A(n1168), .B(G469), .ZN(n965) );
NAND2_X1 U923 ( .A1(n1169), .A2(n1060), .ZN(n1168) );
XNOR2_X1 U924 ( .A(n1170), .B(n1050), .ZN(n1169) );
XNOR2_X1 U925 ( .A(n1171), .B(n1172), .ZN(n1050) );
XNOR2_X1 U926 ( .A(n1142), .B(G110), .ZN(n1172) );
INV_X1 U927 ( .A(G140), .ZN(n1142) );
NAND2_X1 U928 ( .A1(G227), .A2(n976), .ZN(n1171) );
NAND2_X1 U929 ( .A1(KEYINPUT43), .A2(n1173), .ZN(n1170) );
XNOR2_X1 U930 ( .A(n1049), .B(n1174), .ZN(n1173) );
XNOR2_X1 U931 ( .A(n1047), .B(n1175), .ZN(n1174) );
NOR2_X1 U932 ( .A1(KEYINPUT17), .A2(n1048), .ZN(n1175) );
XOR2_X1 U933 ( .A(G146), .B(n1176), .Z(n1048) );
XNOR2_X1 U934 ( .A(n1177), .B(n1178), .ZN(n1047) );
XOR2_X1 U935 ( .A(KEYINPUT14), .B(G107), .Z(n1178) );
XNOR2_X1 U936 ( .A(G104), .B(G101), .ZN(n1177) );
XNOR2_X1 U937 ( .A(n983), .B(KEYINPUT35), .ZN(n1049) );
XNOR2_X1 U938 ( .A(G131), .B(n1179), .ZN(n983) );
XOR2_X1 U939 ( .A(G137), .B(G134), .Z(n1179) );
NOR2_X1 U940 ( .A1(n1088), .A2(n1089), .ZN(n948) );
XNOR2_X1 U941 ( .A(n1180), .B(G475), .ZN(n1089) );
NAND2_X1 U942 ( .A1(n1024), .A2(n1060), .ZN(n1180) );
XOR2_X1 U943 ( .A(n1181), .B(n1182), .Z(n1024) );
XOR2_X1 U944 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U945 ( .A(n1185), .B(n1186), .Z(n1184) );
AND3_X1 U946 ( .A1(G214), .A2(n976), .A3(n1154), .ZN(n1186) );
INV_X1 U947 ( .A(G237), .ZN(n1154) );
NAND2_X1 U948 ( .A1(KEYINPUT15), .A2(n1187), .ZN(n1185) );
NAND2_X1 U949 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
INV_X1 U950 ( .A(n986), .ZN(n1189) );
NOR2_X1 U951 ( .A1(n1058), .A2(G140), .ZN(n986) );
XNOR2_X1 U952 ( .A(KEYINPUT8), .B(n985), .ZN(n1188) );
NAND2_X1 U953 ( .A1(G140), .A2(n1058), .ZN(n985) );
INV_X1 U954 ( .A(G125), .ZN(n1058) );
XNOR2_X1 U955 ( .A(n1190), .B(n1191), .ZN(n1183) );
NOR2_X1 U956 ( .A1(KEYINPUT52), .A2(n1092), .ZN(n1191) );
INV_X1 U957 ( .A(G131), .ZN(n1092) );
NOR2_X1 U958 ( .A1(KEYINPUT5), .A2(n1192), .ZN(n1190) );
XNOR2_X1 U959 ( .A(G113), .B(G122), .ZN(n1192) );
XOR2_X1 U960 ( .A(n1193), .B(n1194), .Z(n1181) );
XNOR2_X1 U961 ( .A(KEYINPUT21), .B(n1138), .ZN(n1194) );
INV_X1 U962 ( .A(G146), .ZN(n1138) );
XNOR2_X1 U963 ( .A(G104), .B(G143), .ZN(n1193) );
XNOR2_X1 U964 ( .A(n1195), .B(G478), .ZN(n1088) );
NAND2_X1 U965 ( .A1(n1018), .A2(n1196), .ZN(n1195) );
XNOR2_X1 U966 ( .A(KEYINPUT22), .B(n1060), .ZN(n1196) );
INV_X1 U967 ( .A(G902), .ZN(n1060) );
XOR2_X1 U968 ( .A(n1197), .B(n1198), .Z(n1018) );
XOR2_X1 U969 ( .A(G116), .B(n1199), .Z(n1198) );
XOR2_X1 U970 ( .A(G134), .B(G122), .Z(n1199) );
XOR2_X1 U971 ( .A(n1200), .B(n1201), .Z(n1197) );
NOR3_X1 U972 ( .A1(n1125), .A2(KEYINPUT51), .A3(n1132), .ZN(n1201) );
NAND2_X1 U973 ( .A1(n1202), .A2(n976), .ZN(n1132) );
INV_X1 U974 ( .A(G953), .ZN(n976) );
XNOR2_X1 U975 ( .A(G234), .B(KEYINPUT48), .ZN(n1202) );
INV_X1 U976 ( .A(G217), .ZN(n1125) );
XOR2_X1 U977 ( .A(n1203), .B(G107), .Z(n1200) );
NAND2_X1 U978 ( .A1(KEYINPUT55), .A2(n1176), .ZN(n1203) );
XNOR2_X1 U979 ( .A(G128), .B(G143), .ZN(n1176) );
endmodule


