//Key = 1110110110100000110100100101010010111111010110000101010000010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;

XOR2_X1 U728 ( .A(G107), .B(n1009), .Z(G9) );
NOR2_X1 U729 ( .A1(KEYINPUT61), .A2(n1010), .ZN(n1009) );
NOR2_X1 U730 ( .A1(n1011), .A2(n1012), .ZN(G75) );
NOR2_X1 U731 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NAND4_X1 U732 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1014) );
NAND3_X1 U733 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1018) );
NAND2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NAND4_X1 U735 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
INV_X1 U736 ( .A(KEYINPUT43), .ZN(n1027) );
NAND2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(n1022) );
NAND2_X1 U738 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NAND4_X1 U739 ( .A1(KEYINPUT22), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n1031) );
INV_X1 U740 ( .A(n1026), .ZN(n1030) );
NAND3_X1 U741 ( .A1(n1035), .A2(n1036), .A3(n1028), .ZN(n1026) );
NAND2_X1 U742 ( .A1(n1024), .A2(n1037), .ZN(n1036) );
NAND2_X1 U743 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND2_X1 U744 ( .A1(KEYINPUT43), .A2(n1025), .ZN(n1039) );
INV_X1 U745 ( .A(n1040), .ZN(n1038) );
NAND2_X1 U746 ( .A1(n1033), .A2(n1041), .ZN(n1035) );
NAND2_X1 U747 ( .A1(KEYINPUT9), .A2(n1042), .ZN(n1017) );
NAND4_X1 U748 ( .A1(n1028), .A2(n1043), .A3(n1044), .A4(n1024), .ZN(n1042) );
NOR2_X1 U749 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND4_X1 U750 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1013) );
NAND4_X1 U751 ( .A1(n1028), .A2(n1024), .A3(n1033), .A4(n1051), .ZN(n1047) );
NAND2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U753 ( .A1(n1021), .A2(n1054), .ZN(n1053) );
NAND2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U755 ( .A1(n1043), .A2(n1057), .ZN(n1056) );
INV_X1 U756 ( .A(KEYINPUT9), .ZN(n1057) );
NAND2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1019), .A2(n1060), .ZN(n1052) );
NAND3_X1 U759 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
OR2_X1 U761 ( .A1(n1045), .A2(KEYINPUT22), .ZN(n1061) );
INV_X1 U762 ( .A(n1066), .ZN(n1028) );
NOR3_X1 U763 ( .A1(n1067), .A2(G953), .A3(G952), .ZN(n1011) );
INV_X1 U764 ( .A(n1049), .ZN(n1067) );
NAND4_X1 U765 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1049) );
NOR4_X1 U766 ( .A1(n1072), .A2(n1032), .A3(n1045), .A4(n1073), .ZN(n1071) );
NOR3_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1070) );
AND3_X1 U768 ( .A1(KEYINPUT51), .A2(n1077), .A3(G475), .ZN(n1076) );
NOR2_X1 U769 ( .A1(KEYINPUT51), .A2(G475), .ZN(n1075) );
XOR2_X1 U770 ( .A(G472), .B(n1078), .Z(n1074) );
XNOR2_X1 U771 ( .A(n1079), .B(n1080), .ZN(n1069) );
XOR2_X1 U772 ( .A(KEYINPUT18), .B(G469), .Z(n1080) );
XNOR2_X1 U773 ( .A(n1081), .B(n1082), .ZN(n1068) );
XNOR2_X1 U774 ( .A(n1083), .B(KEYINPUT47), .ZN(n1081) );
XOR2_X1 U775 ( .A(n1084), .B(n1085), .Z(G72) );
NOR2_X1 U776 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U777 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1050), .ZN(n1089) );
NOR2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
INV_X1 U780 ( .A(n1093), .ZN(n1088) );
NOR2_X1 U781 ( .A1(KEYINPUT44), .A2(n1093), .ZN(n1086) );
NAND2_X1 U782 ( .A1(n1050), .A2(n1094), .ZN(n1093) );
NAND2_X1 U783 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U784 ( .A1(n1097), .A2(n1098), .ZN(n1084) );
XOR2_X1 U785 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U786 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U787 ( .A(n1103), .B(n1104), .Z(n1099) );
XNOR2_X1 U788 ( .A(G140), .B(KEYINPUT16), .ZN(n1104) );
NAND4_X1 U789 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1103) );
NAND3_X1 U790 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1108) );
INV_X1 U791 ( .A(KEYINPUT38), .ZN(n1111) );
OR2_X1 U792 ( .A1(KEYINPUT17), .A2(G137), .ZN(n1109) );
NAND3_X1 U793 ( .A1(G134), .A2(n1112), .A3(KEYINPUT38), .ZN(n1107) );
NAND2_X1 U794 ( .A1(KEYINPUT17), .A2(n1113), .ZN(n1112) );
NAND3_X1 U795 ( .A1(n1114), .A2(n1113), .A3(n1115), .ZN(n1106) );
INV_X1 U796 ( .A(KEYINPUT54), .ZN(n1115) );
XNOR2_X1 U797 ( .A(KEYINPUT17), .B(n1110), .ZN(n1114) );
NAND2_X1 U798 ( .A1(G137), .A2(KEYINPUT54), .ZN(n1105) );
AND2_X1 U799 ( .A1(n1092), .A2(n1116), .ZN(n1097) );
XOR2_X1 U800 ( .A(n1117), .B(n1118), .Z(G69) );
NOR2_X1 U801 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NOR2_X1 U802 ( .A1(G953), .A2(n1121), .ZN(n1120) );
NOR2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XOR2_X1 U804 ( .A(n1048), .B(KEYINPUT39), .Z(n1122) );
NOR2_X1 U805 ( .A1(n1124), .A2(n1050), .ZN(n1119) );
AND2_X1 U806 ( .A1(G224), .A2(G898), .ZN(n1124) );
NAND2_X1 U807 ( .A1(n1125), .A2(n1126), .ZN(n1117) );
NAND2_X1 U808 ( .A1(n1116), .A2(n1127), .ZN(n1126) );
NOR2_X1 U809 ( .A1(n1128), .A2(n1129), .ZN(G66) );
NOR3_X1 U810 ( .A1(n1083), .A2(n1130), .A3(n1131), .ZN(n1129) );
AND3_X1 U811 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1131) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1132), .ZN(n1130) );
AND2_X1 U813 ( .A1(n1136), .A2(n1133), .ZN(n1135) );
NOR2_X1 U814 ( .A1(n1128), .A2(n1137), .ZN(G63) );
XNOR2_X1 U815 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR3_X1 U816 ( .A1(n1140), .A2(KEYINPUT14), .A3(n1141), .ZN(n1139) );
XOR2_X1 U817 ( .A(KEYINPUT27), .B(G478), .Z(n1140) );
NOR2_X1 U818 ( .A1(n1128), .A2(n1142), .ZN(G60) );
XNOR2_X1 U819 ( .A(n1143), .B(n1144), .ZN(n1142) );
AND2_X1 U820 ( .A1(G475), .A2(n1134), .ZN(n1144) );
XOR2_X1 U821 ( .A(n1048), .B(n1145), .Z(G6) );
NOR2_X1 U822 ( .A1(KEYINPUT56), .A2(n1146), .ZN(n1145) );
XNOR2_X1 U823 ( .A(KEYINPUT33), .B(n1147), .ZN(n1146) );
NOR2_X1 U824 ( .A1(n1128), .A2(n1148), .ZN(G57) );
XOR2_X1 U825 ( .A(n1149), .B(n1150), .Z(n1148) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1150) );
AND2_X1 U827 ( .A1(G472), .A2(n1134), .ZN(n1151) );
NOR2_X1 U828 ( .A1(n1128), .A2(n1153), .ZN(G54) );
XOR2_X1 U829 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U830 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U831 ( .A(n1158), .B(n1159), .Z(n1154) );
XNOR2_X1 U832 ( .A(G140), .B(n1160), .ZN(n1159) );
NAND2_X1 U833 ( .A1(KEYINPUT37), .A2(n1161), .ZN(n1158) );
NAND2_X1 U834 ( .A1(n1134), .A2(G469), .ZN(n1161) );
INV_X1 U835 ( .A(n1141), .ZN(n1134) );
NOR2_X1 U836 ( .A1(n1128), .A2(n1162), .ZN(G51) );
XOR2_X1 U837 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U838 ( .A(n1165), .B(n1166), .Z(n1163) );
NOR2_X1 U839 ( .A1(n1167), .A2(n1141), .ZN(n1166) );
NAND2_X1 U840 ( .A1(G902), .A2(n1136), .ZN(n1141) );
NAND3_X1 U841 ( .A1(n1015), .A2(n1048), .A3(n1168), .ZN(n1136) );
XNOR2_X1 U842 ( .A(n1016), .B(KEYINPUT34), .ZN(n1168) );
AND2_X1 U843 ( .A1(n1095), .A2(n1169), .ZN(n1016) );
XOR2_X1 U844 ( .A(KEYINPUT42), .B(n1096), .Z(n1169) );
AND4_X1 U845 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1096) );
NOR2_X1 U846 ( .A1(n1174), .A2(n1175), .ZN(n1170) );
AND2_X1 U847 ( .A1(n1176), .A2(KEYINPUT19), .ZN(n1175) );
NOR3_X1 U848 ( .A1(KEYINPUT19), .A2(n1177), .A3(n1045), .ZN(n1174) );
NOR2_X1 U849 ( .A1(n1046), .A2(n1178), .ZN(n1177) );
AND4_X1 U850 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1095) );
NAND3_X1 U851 ( .A1(n1183), .A2(n1019), .A3(n1040), .ZN(n1048) );
INV_X1 U852 ( .A(n1123), .ZN(n1015) );
NAND4_X1 U853 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1123) );
AND4_X1 U854 ( .A1(n1010), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1187) );
NAND3_X1 U855 ( .A1(n1025), .A2(n1019), .A3(n1183), .ZN(n1010) );
NAND3_X1 U856 ( .A1(n1183), .A2(n1191), .A3(n1033), .ZN(n1186) );
XOR2_X1 U857 ( .A(KEYINPUT50), .B(n1043), .Z(n1191) );
NAND4_X1 U858 ( .A1(n1192), .A2(n1019), .A3(n1193), .A4(n1194), .ZN(n1184) );
NAND2_X1 U859 ( .A1(KEYINPUT4), .A2(n1195), .ZN(n1165) );
INV_X1 U860 ( .A(G125), .ZN(n1195) );
NOR2_X1 U861 ( .A1(n1050), .A2(G952), .ZN(n1128) );
XNOR2_X1 U862 ( .A(G146), .B(n1172), .ZN(G48) );
NAND3_X1 U863 ( .A1(n1040), .A2(n1196), .A3(n1197), .ZN(n1172) );
XNOR2_X1 U864 ( .A(G143), .B(n1198), .ZN(G45) );
NAND2_X1 U865 ( .A1(KEYINPUT59), .A2(n1199), .ZN(n1198) );
INV_X1 U866 ( .A(n1171), .ZN(n1199) );
NAND4_X1 U867 ( .A1(n1200), .A2(n1196), .A3(n1193), .A4(n1194), .ZN(n1171) );
XOR2_X1 U868 ( .A(n1201), .B(n1202), .Z(G42) );
XNOR2_X1 U869 ( .A(G140), .B(KEYINPUT3), .ZN(n1202) );
NAND2_X1 U870 ( .A1(KEYINPUT0), .A2(n1203), .ZN(n1201) );
INV_X1 U871 ( .A(n1173), .ZN(n1203) );
NAND4_X1 U872 ( .A1(n1204), .A2(n1040), .A3(n1021), .A4(n1058), .ZN(n1173) );
NAND3_X1 U873 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(G39) );
NAND2_X1 U874 ( .A1(KEYINPUT28), .A2(n1208), .ZN(n1207) );
NAND3_X1 U875 ( .A1(n1176), .A2(n1209), .A3(n1113), .ZN(n1206) );
INV_X1 U876 ( .A(G137), .ZN(n1113) );
NAND2_X1 U877 ( .A1(G137), .A2(n1210), .ZN(n1205) );
NAND2_X1 U878 ( .A1(n1211), .A2(n1209), .ZN(n1210) );
INV_X1 U879 ( .A(KEYINPUT28), .ZN(n1209) );
XNOR2_X1 U880 ( .A(KEYINPUT6), .B(n1208), .ZN(n1211) );
INV_X1 U881 ( .A(n1176), .ZN(n1208) );
NOR3_X1 U882 ( .A1(n1046), .A2(n1045), .A3(n1178), .ZN(n1176) );
INV_X1 U883 ( .A(n1033), .ZN(n1046) );
NAND2_X1 U884 ( .A1(n1212), .A2(n1213), .ZN(G36) );
NAND2_X1 U885 ( .A1(n1214), .A2(n1110), .ZN(n1213) );
XOR2_X1 U886 ( .A(KEYINPUT36), .B(n1215), .Z(n1212) );
NOR2_X1 U887 ( .A1(n1214), .A2(n1110), .ZN(n1215) );
INV_X1 U888 ( .A(G134), .ZN(n1110) );
INV_X1 U889 ( .A(n1179), .ZN(n1214) );
NAND3_X1 U890 ( .A1(n1021), .A2(n1025), .A3(n1200), .ZN(n1179) );
XNOR2_X1 U891 ( .A(G131), .B(n1182), .ZN(G33) );
NAND3_X1 U892 ( .A1(n1040), .A2(n1021), .A3(n1200), .ZN(n1182) );
AND3_X1 U893 ( .A1(n1041), .A2(n1216), .A3(n1043), .ZN(n1200) );
INV_X1 U894 ( .A(n1045), .ZN(n1021) );
NAND2_X1 U895 ( .A1(n1065), .A2(n1217), .ZN(n1045) );
XOR2_X1 U896 ( .A(G128), .B(n1218), .Z(G30) );
NOR2_X1 U897 ( .A1(KEYINPUT46), .A2(n1180), .ZN(n1218) );
NAND3_X1 U898 ( .A1(n1025), .A2(n1196), .A3(n1197), .ZN(n1180) );
INV_X1 U899 ( .A(n1178), .ZN(n1197) );
NAND2_X1 U900 ( .A1(n1204), .A2(n1219), .ZN(n1178) );
AND3_X1 U901 ( .A1(n1216), .A2(n1059), .A3(n1041), .ZN(n1204) );
XNOR2_X1 U902 ( .A(G101), .B(n1220), .ZN(G3) );
NAND4_X1 U903 ( .A1(KEYINPUT2), .A2(n1043), .A3(n1033), .A4(n1183), .ZN(n1220) );
XNOR2_X1 U904 ( .A(G125), .B(n1181), .ZN(G27) );
NAND4_X1 U905 ( .A1(n1024), .A2(n1196), .A3(n1040), .A4(n1221), .ZN(n1181) );
AND3_X1 U906 ( .A1(n1058), .A2(n1059), .A3(n1216), .ZN(n1221) );
NAND2_X1 U907 ( .A1(n1066), .A2(n1222), .ZN(n1216) );
NAND2_X1 U908 ( .A1(n1223), .A2(n1092), .ZN(n1222) );
INV_X1 U909 ( .A(G900), .ZN(n1092) );
XNOR2_X1 U910 ( .A(G122), .B(n1224), .ZN(G24) );
NAND4_X1 U911 ( .A1(n1225), .A2(n1226), .A3(n1019), .A4(n1227), .ZN(n1224) );
NOR2_X1 U912 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
AND2_X1 U913 ( .A1(n1230), .A2(n1231), .ZN(n1019) );
NAND2_X1 U914 ( .A1(KEYINPUT1), .A2(n1232), .ZN(n1226) );
NAND2_X1 U915 ( .A1(n1233), .A2(n1234), .ZN(n1225) );
INV_X1 U916 ( .A(KEYINPUT1), .ZN(n1234) );
NAND3_X1 U917 ( .A1(n1235), .A2(n1062), .A3(n1024), .ZN(n1233) );
INV_X1 U918 ( .A(n1196), .ZN(n1062) );
XOR2_X1 U919 ( .A(n1236), .B(G119), .Z(G21) );
NAND2_X1 U920 ( .A1(KEYINPUT53), .A2(n1185), .ZN(n1236) );
NAND4_X1 U921 ( .A1(n1192), .A2(n1033), .A3(n1219), .A4(n1059), .ZN(n1185) );
XNOR2_X1 U922 ( .A(G116), .B(n1190), .ZN(G18) );
NAND3_X1 U923 ( .A1(n1192), .A2(n1025), .A3(n1043), .ZN(n1190) );
NOR2_X1 U924 ( .A1(n1194), .A2(n1229), .ZN(n1025) );
INV_X1 U925 ( .A(n1193), .ZN(n1229) );
XOR2_X1 U926 ( .A(n1189), .B(n1237), .Z(G15) );
NOR2_X1 U927 ( .A1(G113), .A2(KEYINPUT23), .ZN(n1237) );
NAND3_X1 U928 ( .A1(n1192), .A2(n1040), .A3(n1043), .ZN(n1189) );
AND2_X1 U929 ( .A1(n1219), .A2(n1230), .ZN(n1043) );
XNOR2_X1 U930 ( .A(n1059), .B(KEYINPUT40), .ZN(n1230) );
INV_X1 U931 ( .A(n1231), .ZN(n1219) );
NOR2_X1 U932 ( .A1(n1193), .A2(n1228), .ZN(n1040) );
INV_X1 U933 ( .A(n1232), .ZN(n1192) );
NAND3_X1 U934 ( .A1(n1196), .A2(n1235), .A3(n1024), .ZN(n1232) );
AND2_X1 U935 ( .A1(n1034), .A2(n1238), .ZN(n1024) );
XNOR2_X1 U936 ( .A(G110), .B(n1188), .ZN(G12) );
NAND4_X1 U937 ( .A1(n1033), .A2(n1183), .A3(n1058), .A4(n1059), .ZN(n1188) );
NAND3_X1 U938 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1059) );
NAND2_X1 U939 ( .A1(n1083), .A2(n1082), .ZN(n1241) );
NAND2_X1 U940 ( .A1(KEYINPUT12), .A2(n1242), .ZN(n1240) );
NAND2_X1 U941 ( .A1(n1133), .A2(n1243), .ZN(n1242) );
XNOR2_X1 U942 ( .A(KEYINPUT41), .B(n1244), .ZN(n1243) );
NAND2_X1 U943 ( .A1(n1245), .A2(n1246), .ZN(n1239) );
INV_X1 U944 ( .A(KEYINPUT12), .ZN(n1246) );
NAND2_X1 U945 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
OR2_X1 U946 ( .A1(n1244), .A2(KEYINPUT41), .ZN(n1248) );
NAND3_X1 U947 ( .A1(n1133), .A2(n1244), .A3(KEYINPUT41), .ZN(n1247) );
INV_X1 U948 ( .A(n1083), .ZN(n1244) );
NOR2_X1 U949 ( .A1(n1132), .A2(G902), .ZN(n1083) );
XNOR2_X1 U950 ( .A(n1249), .B(n1250), .ZN(n1132) );
XOR2_X1 U951 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U952 ( .A(n1253), .B(n1254), .Z(n1249) );
XOR2_X1 U953 ( .A(n1255), .B(G128), .Z(n1253) );
NAND2_X1 U954 ( .A1(KEYINPUT8), .A2(n1256), .ZN(n1255) );
XNOR2_X1 U955 ( .A(G137), .B(n1257), .ZN(n1256) );
NAND3_X1 U956 ( .A1(G234), .A2(n1258), .A3(G221), .ZN(n1257) );
XNOR2_X1 U957 ( .A(KEYINPUT25), .B(n1050), .ZN(n1258) );
INV_X1 U958 ( .A(n1082), .ZN(n1133) );
NAND2_X1 U959 ( .A1(G217), .A2(n1259), .ZN(n1082) );
XOR2_X1 U960 ( .A(n1231), .B(KEYINPUT31), .Z(n1058) );
XOR2_X1 U961 ( .A(G472), .B(n1260), .Z(n1231) );
NOR2_X1 U962 ( .A1(n1078), .A2(KEYINPUT45), .ZN(n1260) );
AND2_X1 U963 ( .A1(n1261), .A2(n1262), .ZN(n1078) );
XNOR2_X1 U964 ( .A(n1152), .B(n1263), .ZN(n1261) );
XOR2_X1 U965 ( .A(n1264), .B(KEYINPUT10), .Z(n1263) );
NAND2_X1 U966 ( .A1(KEYINPUT7), .A2(n1149), .ZN(n1264) );
XNOR2_X1 U967 ( .A(n1265), .B(G101), .ZN(n1149) );
NAND3_X1 U968 ( .A1(n1266), .A2(n1050), .A3(G210), .ZN(n1265) );
XNOR2_X1 U969 ( .A(n1267), .B(n1268), .ZN(n1152) );
XNOR2_X1 U970 ( .A(n1269), .B(n1270), .ZN(n1268) );
INV_X1 U971 ( .A(n1271), .ZN(n1269) );
XNOR2_X1 U972 ( .A(n1272), .B(n1273), .ZN(n1267) );
INV_X1 U973 ( .A(n1274), .ZN(n1273) );
NAND2_X1 U974 ( .A1(n1275), .A2(n1276), .ZN(n1272) );
NAND3_X1 U975 ( .A1(G116), .A2(n1254), .A3(n1277), .ZN(n1276) );
INV_X1 U976 ( .A(KEYINPUT32), .ZN(n1277) );
NAND2_X1 U977 ( .A1(KEYINPUT32), .A2(n1278), .ZN(n1275) );
AND3_X1 U978 ( .A1(n1041), .A2(n1235), .A3(n1196), .ZN(n1183) );
NOR2_X1 U979 ( .A1(n1065), .A2(n1064), .ZN(n1196) );
INV_X1 U980 ( .A(n1217), .ZN(n1064) );
NAND2_X1 U981 ( .A1(G214), .A2(n1279), .ZN(n1217) );
XNOR2_X1 U982 ( .A(n1280), .B(n1167), .ZN(n1065) );
NAND2_X1 U983 ( .A1(G210), .A2(n1279), .ZN(n1167) );
NAND2_X1 U984 ( .A1(n1266), .A2(n1262), .ZN(n1279) );
INV_X1 U985 ( .A(G237), .ZN(n1266) );
NAND2_X1 U986 ( .A1(n1281), .A2(n1262), .ZN(n1280) );
XNOR2_X1 U987 ( .A(n1164), .B(G125), .ZN(n1281) );
XOR2_X1 U988 ( .A(n1125), .B(n1282), .Z(n1164) );
XNOR2_X1 U989 ( .A(n1283), .B(n1271), .ZN(n1282) );
XOR2_X1 U990 ( .A(n1284), .B(n1285), .Z(n1271) );
XOR2_X1 U991 ( .A(KEYINPUT15), .B(n1286), .Z(n1285) );
NOR2_X1 U992 ( .A1(KEYINPUT24), .A2(n1287), .ZN(n1286) );
INV_X1 U993 ( .A(G146), .ZN(n1287) );
NAND2_X1 U994 ( .A1(G224), .A2(n1050), .ZN(n1283) );
XNOR2_X1 U995 ( .A(n1288), .B(n1157), .ZN(n1125) );
XNOR2_X1 U996 ( .A(n1289), .B(n1290), .ZN(n1157) );
INV_X1 U997 ( .A(G110), .ZN(n1289) );
XOR2_X1 U998 ( .A(n1291), .B(n1292), .Z(n1288) );
NAND3_X1 U999 ( .A1(n1293), .A2(n1294), .A3(n1295), .ZN(n1291) );
NAND2_X1 U1000 ( .A1(KEYINPUT60), .A2(n1278), .ZN(n1295) );
NAND3_X1 U1001 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1294) );
INV_X1 U1002 ( .A(KEYINPUT60), .ZN(n1297) );
OR2_X1 U1003 ( .A1(n1298), .A2(n1296), .ZN(n1293) );
NOR2_X1 U1004 ( .A1(n1299), .A2(n1278), .ZN(n1296) );
XOR2_X1 U1005 ( .A(G116), .B(n1254), .Z(n1278) );
XOR2_X1 U1006 ( .A(G119), .B(KEYINPUT35), .Z(n1254) );
INV_X1 U1007 ( .A(KEYINPUT29), .ZN(n1299) );
NAND2_X1 U1008 ( .A1(n1066), .A2(n1300), .ZN(n1235) );
NAND2_X1 U1009 ( .A1(n1223), .A2(n1127), .ZN(n1300) );
INV_X1 U1010 ( .A(G898), .ZN(n1127) );
AND3_X1 U1011 ( .A1(n1116), .A2(n1301), .A3(n1302), .ZN(n1223) );
XNOR2_X1 U1012 ( .A(G902), .B(KEYINPUT5), .ZN(n1302) );
XOR2_X1 U1013 ( .A(G953), .B(KEYINPUT13), .Z(n1116) );
NAND3_X1 U1014 ( .A1(n1301), .A2(n1050), .A3(G952), .ZN(n1066) );
NAND2_X1 U1015 ( .A1(G237), .A2(G234), .ZN(n1301) );
NOR2_X1 U1016 ( .A1(n1034), .A2(n1032), .ZN(n1041) );
INV_X1 U1017 ( .A(n1238), .ZN(n1032) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1259), .ZN(n1238) );
NAND2_X1 U1019 ( .A1(G234), .A2(n1262), .ZN(n1259) );
XOR2_X1 U1020 ( .A(G469), .B(n1303), .Z(n1034) );
NOR2_X1 U1021 ( .A1(n1079), .A2(KEYINPUT20), .ZN(n1303) );
AND2_X1 U1022 ( .A1(n1304), .A2(n1262), .ZN(n1079) );
XNOR2_X1 U1023 ( .A(n1156), .B(n1305), .ZN(n1304) );
XNOR2_X1 U1024 ( .A(n1306), .B(n1290), .ZN(n1305) );
XOR2_X1 U1025 ( .A(G101), .B(G107), .Z(n1290) );
NAND2_X1 U1026 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
NAND2_X1 U1027 ( .A1(n1160), .A2(n1309), .ZN(n1308) );
XOR2_X1 U1028 ( .A(n1310), .B(KEYINPUT58), .Z(n1307) );
OR2_X1 U1029 ( .A1(n1309), .A2(n1160), .ZN(n1310) );
NOR2_X1 U1030 ( .A1(n1091), .A2(G953), .ZN(n1160) );
INV_X1 U1031 ( .A(G227), .ZN(n1091) );
XOR2_X1 U1032 ( .A(n1251), .B(KEYINPUT62), .Z(n1309) );
XOR2_X1 U1033 ( .A(G110), .B(G140), .Z(n1251) );
XNOR2_X1 U1034 ( .A(n1311), .B(n1312), .ZN(n1156) );
XNOR2_X1 U1035 ( .A(n1274), .B(n1102), .ZN(n1312) );
XOR2_X1 U1036 ( .A(n1313), .B(n1314), .Z(n1102) );
NOR2_X1 U1037 ( .A1(KEYINPUT55), .A2(n1315), .ZN(n1314) );
XNOR2_X1 U1038 ( .A(KEYINPUT15), .B(n1316), .ZN(n1315) );
XNOR2_X1 U1039 ( .A(G131), .B(G128), .ZN(n1313) );
XNOR2_X1 U1040 ( .A(n1317), .B(n1318), .ZN(n1274) );
NOR2_X1 U1041 ( .A1(KEYINPUT52), .A2(G134), .ZN(n1318) );
XNOR2_X1 U1042 ( .A(G137), .B(KEYINPUT48), .ZN(n1317) );
XNOR2_X1 U1043 ( .A(G104), .B(G146), .ZN(n1311) );
NOR2_X1 U1044 ( .A1(n1193), .A2(n1194), .ZN(n1033) );
INV_X1 U1045 ( .A(n1228), .ZN(n1194) );
NOR2_X1 U1046 ( .A1(n1072), .A2(n1319), .ZN(n1228) );
AND2_X1 U1047 ( .A1(G475), .A2(n1077), .ZN(n1319) );
NOR2_X1 U1048 ( .A1(n1077), .A2(G475), .ZN(n1072) );
NAND2_X1 U1049 ( .A1(n1143), .A2(n1262), .ZN(n1077) );
XNOR2_X1 U1050 ( .A(n1320), .B(n1321), .ZN(n1143) );
XOR2_X1 U1051 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1052 ( .A(n1324), .B(n1325), .ZN(n1323) );
NOR2_X1 U1053 ( .A1(G140), .A2(KEYINPUT11), .ZN(n1325) );
NAND2_X1 U1054 ( .A1(KEYINPUT49), .A2(n1316), .ZN(n1324) );
XOR2_X1 U1055 ( .A(KEYINPUT26), .B(n1326), .Z(n1322) );
NOR3_X1 U1056 ( .A1(n1327), .A2(G237), .A3(n1328), .ZN(n1326) );
INV_X1 U1057 ( .A(G214), .ZN(n1328) );
XNOR2_X1 U1058 ( .A(KEYINPUT57), .B(n1050), .ZN(n1327) );
XOR2_X1 U1059 ( .A(n1329), .B(n1292), .Z(n1320) );
XNOR2_X1 U1060 ( .A(n1147), .B(G122), .ZN(n1292) );
INV_X1 U1061 ( .A(G104), .ZN(n1147) );
XNOR2_X1 U1062 ( .A(n1270), .B(n1252), .ZN(n1329) );
XNOR2_X1 U1063 ( .A(n1101), .B(KEYINPUT30), .ZN(n1252) );
XNOR2_X1 U1064 ( .A(G125), .B(G146), .ZN(n1101) );
XNOR2_X1 U1065 ( .A(G131), .B(n1298), .ZN(n1270) );
INV_X1 U1066 ( .A(G113), .ZN(n1298) );
XOR2_X1 U1067 ( .A(n1073), .B(KEYINPUT21), .Z(n1193) );
XNOR2_X1 U1068 ( .A(n1330), .B(G478), .ZN(n1073) );
NAND2_X1 U1069 ( .A1(n1138), .A2(n1262), .ZN(n1330) );
INV_X1 U1070 ( .A(G902), .ZN(n1262) );
XNOR2_X1 U1071 ( .A(n1331), .B(n1332), .ZN(n1138) );
XOR2_X1 U1072 ( .A(n1333), .B(n1284), .Z(n1332) );
XNOR2_X1 U1073 ( .A(G128), .B(n1316), .ZN(n1284) );
INV_X1 U1074 ( .A(G143), .ZN(n1316) );
AND3_X1 U1075 ( .A1(G217), .A2(n1050), .A3(G234), .ZN(n1333) );
INV_X1 U1076 ( .A(G953), .ZN(n1050) );
XOR2_X1 U1077 ( .A(n1334), .B(n1335), .Z(n1331) );
NOR2_X1 U1078 ( .A1(KEYINPUT63), .A2(n1336), .ZN(n1335) );
XNOR2_X1 U1079 ( .A(G122), .B(G116), .ZN(n1336) );
XNOR2_X1 U1080 ( .A(G107), .B(G134), .ZN(n1334) );
endmodule


