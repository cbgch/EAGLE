//Key = 1000101100100011001101111100111011110010101110111011111100111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393;

XNOR2_X1 U760 ( .A(n1059), .B(n1060), .ZN(G9) );
XOR2_X1 U761 ( .A(KEYINPUT60), .B(G107), .Z(n1060) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(G75) );
NOR4_X1 U763 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
NOR4_X1 U764 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1065) );
NOR3_X1 U765 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1068) );
NOR2_X1 U766 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR2_X1 U767 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR4_X1 U768 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1072) );
INV_X1 U769 ( .A(KEYINPUT18), .ZN(n1081) );
NOR2_X1 U770 ( .A1(n1082), .A2(n1083), .ZN(n1067) );
NOR4_X1 U771 ( .A1(KEYINPUT18), .A2(n1079), .A3(n1078), .A4(n1080), .ZN(n1083) );
XOR2_X1 U772 ( .A(KEYINPUT41), .B(n1084), .Z(n1064) );
NOR3_X1 U773 ( .A1(n1085), .A2(n1078), .A3(n1071), .ZN(n1084) );
NAND3_X1 U774 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
NAND3_X1 U775 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1063) );
NAND4_X1 U776 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091) );
NAND3_X1 U777 ( .A1(n1096), .A2(n1097), .A3(n1071), .ZN(n1095) );
NAND3_X1 U778 ( .A1(n1098), .A2(n1099), .A3(n1088), .ZN(n1097) );
INV_X1 U779 ( .A(KEYINPUT58), .ZN(n1099) );
NAND2_X1 U780 ( .A1(n1100), .A2(n1101), .ZN(n1096) );
INV_X1 U781 ( .A(KEYINPUT53), .ZN(n1101) );
NAND4_X1 U782 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1082), .ZN(n1094) );
INV_X1 U783 ( .A(n1071), .ZN(n1082) );
NAND2_X1 U784 ( .A1(KEYINPUT53), .A2(n1100), .ZN(n1104) );
NAND3_X1 U785 ( .A1(n1105), .A2(n1087), .A3(n1106), .ZN(n1103) );
NAND2_X1 U786 ( .A1(n1088), .A2(n1107), .ZN(n1102) );
NAND2_X1 U787 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U788 ( .A1(KEYINPUT58), .A2(n1098), .ZN(n1109) );
INV_X1 U789 ( .A(n1110), .ZN(n1108) );
NOR3_X1 U790 ( .A1(n1111), .A2(G953), .A3(G952), .ZN(n1061) );
INV_X1 U791 ( .A(n1089), .ZN(n1111) );
NAND4_X1 U792 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1089) );
NOR4_X1 U793 ( .A1(n1116), .A2(n1117), .A3(n1070), .A4(n1075), .ZN(n1115) );
XOR2_X1 U794 ( .A(n1118), .B(KEYINPUT30), .Z(n1117) );
NOR2_X1 U795 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
NOR3_X1 U796 ( .A1(n1121), .A2(KEYINPUT5), .A3(n1122), .ZN(n1120) );
AND2_X1 U797 ( .A1(n1121), .A2(KEYINPUT5), .ZN(n1119) );
XOR2_X1 U798 ( .A(n1123), .B(n1124), .Z(n1113) );
XOR2_X1 U799 ( .A(KEYINPUT33), .B(n1125), .Z(n1124) );
NAND2_X1 U800 ( .A1(KEYINPUT10), .A2(n1126), .ZN(n1123) );
XOR2_X1 U801 ( .A(n1127), .B(KEYINPUT38), .Z(n1112) );
XOR2_X1 U802 ( .A(n1128), .B(n1129), .Z(G72) );
NOR2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U804 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U805 ( .A1(KEYINPUT43), .A2(n1134), .ZN(n1133) );
NAND2_X1 U806 ( .A1(n1135), .A2(n1136), .ZN(n1132) );
NAND3_X1 U807 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
XOR2_X1 U808 ( .A(KEYINPUT34), .B(n1140), .Z(n1135) );
NOR2_X1 U809 ( .A1(n1141), .A2(n1137), .ZN(n1140) );
XNOR2_X1 U810 ( .A(n1142), .B(n1143), .ZN(n1137) );
AND2_X1 U811 ( .A1(n1138), .A2(n1139), .ZN(n1141) );
INV_X1 U812 ( .A(n1144), .ZN(n1139) );
NAND2_X1 U813 ( .A1(n1145), .A2(n1146), .ZN(n1128) );
NAND2_X1 U814 ( .A1(n1147), .A2(n1090), .ZN(n1146) );
NAND2_X1 U815 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U816 ( .A1(G953), .A2(n1150), .ZN(n1145) );
NAND2_X1 U817 ( .A1(n1151), .A2(G227), .ZN(n1150) );
XNOR2_X1 U818 ( .A(G900), .B(KEYINPUT46), .ZN(n1151) );
XOR2_X1 U819 ( .A(n1152), .B(n1153), .Z(G69) );
XOR2_X1 U820 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U821 ( .A1(G953), .A2(n1156), .ZN(n1155) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1156) );
NAND2_X1 U823 ( .A1(n1157), .A2(n1158), .ZN(n1154) );
NAND2_X1 U824 ( .A1(G953), .A2(n1159), .ZN(n1158) );
XOR2_X1 U825 ( .A(n1160), .B(n1161), .Z(n1157) );
NOR2_X1 U826 ( .A1(n1162), .A2(G953), .ZN(n1152) );
NOR3_X1 U827 ( .A1(n1163), .A2(n1164), .A3(n1165), .ZN(G66) );
NOR3_X1 U828 ( .A1(n1166), .A2(G953), .A3(n1167), .ZN(n1165) );
AND2_X1 U829 ( .A1(n1166), .A2(n1168), .ZN(n1164) );
INV_X1 U830 ( .A(KEYINPUT3), .ZN(n1166) );
XOR2_X1 U831 ( .A(n1169), .B(n1170), .Z(n1163) );
NAND2_X1 U832 ( .A1(KEYINPUT22), .A2(n1171), .ZN(n1170) );
NAND2_X1 U833 ( .A1(n1172), .A2(n1125), .ZN(n1169) );
NOR2_X1 U834 ( .A1(n1168), .A2(n1173), .ZN(G63) );
XOR2_X1 U835 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND3_X1 U836 ( .A1(G478), .A2(G902), .A3(n1176), .ZN(n1174) );
XOR2_X1 U837 ( .A(n1066), .B(KEYINPUT8), .Z(n1176) );
NOR2_X1 U838 ( .A1(n1168), .A2(n1177), .ZN(G60) );
XOR2_X1 U839 ( .A(n1178), .B(n1179), .Z(n1177) );
NOR2_X1 U840 ( .A1(n1121), .A2(n1180), .ZN(n1178) );
NAND2_X1 U841 ( .A1(n1181), .A2(n1182), .ZN(G6) );
NAND2_X1 U842 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND2_X1 U843 ( .A1(G104), .A2(n1185), .ZN(n1181) );
NAND2_X1 U844 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U845 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
OR2_X1 U846 ( .A1(n1189), .A2(n1183), .ZN(n1186) );
NOR2_X1 U847 ( .A1(KEYINPUT17), .A2(n1190), .ZN(n1183) );
INV_X1 U848 ( .A(KEYINPUT23), .ZN(n1189) );
NOR2_X1 U849 ( .A1(n1168), .A2(n1191), .ZN(G57) );
XOR2_X1 U850 ( .A(n1192), .B(n1193), .Z(n1191) );
NAND2_X1 U851 ( .A1(n1194), .A2(KEYINPUT28), .ZN(n1192) );
XOR2_X1 U852 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U853 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U854 ( .A(n1199), .B(KEYINPUT63), .Z(n1195) );
NAND3_X1 U855 ( .A1(n1200), .A2(n1201), .A3(G472), .ZN(n1199) );
NAND2_X1 U856 ( .A1(KEYINPUT14), .A2(n1180), .ZN(n1201) );
NAND2_X1 U857 ( .A1(n1202), .A2(n1203), .ZN(n1200) );
INV_X1 U858 ( .A(KEYINPUT14), .ZN(n1203) );
OR2_X1 U859 ( .A1(n1066), .A2(n1204), .ZN(n1202) );
NOR2_X1 U860 ( .A1(n1168), .A2(n1205), .ZN(G54) );
NOR2_X1 U861 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
XOR2_X1 U862 ( .A(n1208), .B(n1209), .Z(n1207) );
NOR2_X1 U863 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
AND2_X1 U864 ( .A1(G469), .A2(n1172), .ZN(n1208) );
INV_X1 U865 ( .A(n1180), .ZN(n1172) );
AND2_X1 U866 ( .A1(n1211), .A2(n1210), .ZN(n1206) );
XNOR2_X1 U867 ( .A(n1212), .B(n1213), .ZN(n1210) );
XNOR2_X1 U868 ( .A(n1214), .B(KEYINPUT4), .ZN(n1213) );
NAND2_X1 U869 ( .A1(n1215), .A2(KEYINPUT21), .ZN(n1214) );
XOR2_X1 U870 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U871 ( .A(n1218), .B(KEYINPUT57), .Z(n1216) );
NAND2_X1 U872 ( .A1(KEYINPUT54), .A2(n1219), .ZN(n1218) );
INV_X1 U873 ( .A(G140), .ZN(n1219) );
INV_X1 U874 ( .A(KEYINPUT19), .ZN(n1211) );
NOR2_X1 U875 ( .A1(n1168), .A2(n1220), .ZN(G51) );
XOR2_X1 U876 ( .A(n1221), .B(n1222), .Z(n1220) );
XNOR2_X1 U877 ( .A(n1223), .B(n1224), .ZN(n1222) );
XOR2_X1 U878 ( .A(n1225), .B(n1226), .Z(n1221) );
XNOR2_X1 U879 ( .A(KEYINPUT45), .B(n1227), .ZN(n1226) );
NOR2_X1 U880 ( .A1(n1228), .A2(n1180), .ZN(n1225) );
NAND2_X1 U881 ( .A1(G902), .A2(n1066), .ZN(n1180) );
NAND3_X1 U882 ( .A1(n1162), .A2(n1148), .A3(n1229), .ZN(n1066) );
XOR2_X1 U883 ( .A(n1149), .B(KEYINPUT36), .Z(n1229) );
NAND2_X1 U884 ( .A1(n1230), .A2(n1076), .ZN(n1149) );
AND4_X1 U885 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1148) );
AND4_X1 U886 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1234) );
NAND2_X1 U887 ( .A1(n1239), .A2(n1098), .ZN(n1233) );
NAND3_X1 U888 ( .A1(n1077), .A2(n1240), .A3(n1241), .ZN(n1232) );
NOR3_X1 U889 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1241) );
XOR2_X1 U890 ( .A(n1245), .B(KEYINPUT32), .Z(n1243) );
NAND4_X1 U891 ( .A1(n1246), .A2(n1247), .A3(n1092), .A4(n1093), .ZN(n1231) );
XOR2_X1 U892 ( .A(n1248), .B(KEYINPUT51), .Z(n1246) );
AND4_X1 U893 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1162) );
NOR4_X1 U894 ( .A1(n1059), .A2(n1253), .A3(n1254), .A4(n1255), .ZN(n1252) );
AND3_X1 U895 ( .A1(n1100), .A2(n1076), .A3(n1256), .ZN(n1059) );
NOR2_X1 U896 ( .A1(n1257), .A2(n1188), .ZN(n1251) );
INV_X1 U897 ( .A(n1190), .ZN(n1188) );
NAND3_X1 U898 ( .A1(n1256), .A2(n1100), .A3(n1077), .ZN(n1190) );
NOR2_X1 U899 ( .A1(n1242), .A2(n1069), .ZN(n1100) );
INV_X1 U900 ( .A(n1087), .ZN(n1069) );
INV_X1 U901 ( .A(n1258), .ZN(n1256) );
NOR3_X1 U902 ( .A1(n1259), .A2(n1260), .A3(n1258), .ZN(n1257) );
XOR2_X1 U903 ( .A(n1070), .B(KEYINPUT16), .Z(n1260) );
NOR2_X1 U904 ( .A1(n1090), .A2(n1167), .ZN(n1168) );
XNOR2_X1 U905 ( .A(G952), .B(KEYINPUT55), .ZN(n1167) );
XNOR2_X1 U906 ( .A(G146), .B(n1261), .ZN(G48) );
NAND4_X1 U907 ( .A1(n1247), .A2(n1077), .A3(n1262), .A4(n1240), .ZN(n1261) );
NOR2_X1 U908 ( .A1(KEYINPUT37), .A2(n1244), .ZN(n1262) );
XOR2_X1 U909 ( .A(n1263), .B(G143), .Z(G45) );
NAND2_X1 U910 ( .A1(KEYINPUT61), .A2(n1238), .ZN(n1263) );
NAND3_X1 U911 ( .A1(n1247), .A2(n1110), .A3(n1264), .ZN(n1238) );
NOR3_X1 U912 ( .A1(n1244), .A2(n1265), .A3(n1118), .ZN(n1264) );
XOR2_X1 U913 ( .A(n1237), .B(n1266), .Z(G42) );
NAND2_X1 U914 ( .A1(KEYINPUT52), .A2(G140), .ZN(n1266) );
NAND4_X1 U915 ( .A1(n1247), .A2(n1077), .A3(n1093), .A4(n1098), .ZN(n1237) );
XOR2_X1 U916 ( .A(n1267), .B(n1268), .Z(G39) );
NAND2_X1 U917 ( .A1(n1093), .A2(n1269), .ZN(n1268) );
XOR2_X1 U918 ( .A(KEYINPUT1), .B(n1270), .Z(n1269) );
NOR2_X1 U919 ( .A1(n1259), .A2(n1271), .ZN(n1270) );
XOR2_X1 U920 ( .A(G134), .B(n1272), .Z(G36) );
NOR2_X1 U921 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XOR2_X1 U922 ( .A(KEYINPUT7), .B(n1076), .Z(n1274) );
NAND3_X1 U923 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(G33) );
NAND2_X1 U924 ( .A1(n1236), .A2(n1278), .ZN(n1277) );
OR3_X1 U925 ( .A1(n1278), .A2(n1236), .A3(G131), .ZN(n1276) );
INV_X1 U926 ( .A(KEYINPUT6), .ZN(n1278) );
NAND2_X1 U927 ( .A1(G131), .A2(n1279), .ZN(n1275) );
NAND2_X1 U928 ( .A1(KEYINPUT6), .A2(n1280), .ZN(n1279) );
XNOR2_X1 U929 ( .A(KEYINPUT56), .B(n1236), .ZN(n1280) );
NAND2_X1 U930 ( .A1(n1230), .A2(n1077), .ZN(n1236) );
INV_X1 U931 ( .A(n1273), .ZN(n1230) );
NAND3_X1 U932 ( .A1(n1093), .A2(n1110), .A3(n1247), .ZN(n1273) );
INV_X1 U933 ( .A(n1075), .ZN(n1093) );
NAND2_X1 U934 ( .A1(n1281), .A2(n1080), .ZN(n1075) );
XNOR2_X1 U935 ( .A(G128), .B(n1235), .ZN(G30) );
NAND4_X1 U936 ( .A1(n1247), .A2(n1240), .A3(n1076), .A4(n1086), .ZN(n1235) );
INV_X1 U937 ( .A(n1271), .ZN(n1247) );
NAND2_X1 U938 ( .A1(n1282), .A2(n1245), .ZN(n1271) );
XNOR2_X1 U939 ( .A(G101), .B(n1249), .ZN(G3) );
NAND2_X1 U940 ( .A1(n1283), .A2(n1110), .ZN(n1249) );
XNOR2_X1 U941 ( .A(G125), .B(n1284), .ZN(G27) );
NAND2_X1 U942 ( .A1(n1285), .A2(n1239), .ZN(n1284) );
AND4_X1 U943 ( .A1(n1077), .A2(n1088), .A3(n1086), .A4(n1245), .ZN(n1239) );
NAND2_X1 U944 ( .A1(n1071), .A2(n1286), .ZN(n1245) );
NAND3_X1 U945 ( .A1(G902), .A2(n1287), .A3(n1130), .ZN(n1286) );
NOR2_X1 U946 ( .A1(n1090), .A2(G900), .ZN(n1130) );
INV_X1 U947 ( .A(n1070), .ZN(n1088) );
XNOR2_X1 U948 ( .A(KEYINPUT40), .B(n1098), .ZN(n1285) );
XNOR2_X1 U949 ( .A(n1250), .B(n1288), .ZN(G24) );
NOR2_X1 U950 ( .A1(KEYINPUT27), .A2(n1289), .ZN(n1288) );
NAND4_X1 U951 ( .A1(n1290), .A2(n1291), .A3(n1087), .A4(n1292), .ZN(n1250) );
NAND2_X1 U952 ( .A1(n1293), .A2(n1294), .ZN(n1087) );
OR3_X1 U953 ( .A1(n1127), .A2(n1295), .A3(KEYINPUT12), .ZN(n1294) );
NAND2_X1 U954 ( .A1(KEYINPUT12), .A2(n1110), .ZN(n1293) );
XOR2_X1 U955 ( .A(n1296), .B(n1297), .Z(G21) );
NOR2_X1 U956 ( .A1(KEYINPUT39), .A2(G119), .ZN(n1297) );
NAND2_X1 U957 ( .A1(n1298), .A2(n1290), .ZN(n1296) );
INV_X1 U958 ( .A(n1259), .ZN(n1298) );
NAND2_X1 U959 ( .A1(n1240), .A2(n1092), .ZN(n1259) );
INV_X1 U960 ( .A(n1078), .ZN(n1092) );
XOR2_X1 U961 ( .A(G116), .B(n1255), .Z(G18) );
AND3_X1 U962 ( .A1(n1076), .A2(n1110), .A3(n1290), .ZN(n1255) );
NOR2_X1 U963 ( .A1(n1292), .A2(n1118), .ZN(n1076) );
INV_X1 U964 ( .A(n1265), .ZN(n1292) );
NAND2_X1 U965 ( .A1(n1299), .A2(n1300), .ZN(G15) );
NAND2_X1 U966 ( .A1(n1254), .A2(n1301), .ZN(n1300) );
NAND2_X1 U967 ( .A1(G113), .A2(n1302), .ZN(n1301) );
OR2_X1 U968 ( .A1(n1303), .A2(KEYINPUT29), .ZN(n1302) );
INV_X1 U969 ( .A(n1304), .ZN(n1254) );
NAND3_X1 U970 ( .A1(n1305), .A2(n1306), .A3(KEYINPUT29), .ZN(n1299) );
NAND2_X1 U971 ( .A1(G113), .A2(n1303), .ZN(n1306) );
INV_X1 U972 ( .A(KEYINPUT15), .ZN(n1303) );
NAND2_X1 U973 ( .A1(KEYINPUT15), .A2(n1307), .ZN(n1305) );
NAND2_X1 U974 ( .A1(G113), .A2(n1304), .ZN(n1307) );
NAND3_X1 U975 ( .A1(n1290), .A2(n1110), .A3(n1077), .ZN(n1304) );
NOR2_X1 U976 ( .A1(n1291), .A2(n1265), .ZN(n1077) );
INV_X1 U977 ( .A(n1118), .ZN(n1291) );
NOR2_X1 U978 ( .A1(n1295), .A2(n1308), .ZN(n1110) );
NOR2_X1 U979 ( .A1(n1070), .A2(n1258), .ZN(n1290) );
NAND2_X1 U980 ( .A1(n1105), .A2(n1309), .ZN(n1070) );
XOR2_X1 U981 ( .A(G110), .B(n1253), .Z(G12) );
AND2_X1 U982 ( .A1(n1283), .A2(n1098), .ZN(n1253) );
NAND2_X1 U983 ( .A1(n1310), .A2(n1311), .ZN(n1098) );
NAND3_X1 U984 ( .A1(n1308), .A2(n1295), .A3(n1312), .ZN(n1311) );
INV_X1 U985 ( .A(KEYINPUT12), .ZN(n1312) );
INV_X1 U986 ( .A(n1127), .ZN(n1308) );
NAND2_X1 U987 ( .A1(KEYINPUT12), .A2(n1240), .ZN(n1310) );
INV_X1 U988 ( .A(n1248), .ZN(n1240) );
NAND2_X1 U989 ( .A1(n1127), .A2(n1295), .ZN(n1248) );
XNOR2_X1 U990 ( .A(n1126), .B(n1125), .ZN(n1295) );
AND2_X1 U991 ( .A1(G217), .A2(n1313), .ZN(n1125) );
OR2_X1 U992 ( .A1(n1171), .A2(G902), .ZN(n1126) );
XOR2_X1 U993 ( .A(n1314), .B(n1315), .Z(n1171) );
XOR2_X1 U994 ( .A(n1316), .B(n1317), .Z(n1315) );
XOR2_X1 U995 ( .A(G128), .B(n1318), .Z(n1317) );
AND3_X1 U996 ( .A1(G221), .A2(n1090), .A3(G234), .ZN(n1318) );
XOR2_X1 U997 ( .A(KEYINPUT42), .B(G137), .Z(n1316) );
XNOR2_X1 U998 ( .A(n1319), .B(n1320), .ZN(n1314) );
XNOR2_X1 U999 ( .A(n1321), .B(n1322), .ZN(n1320) );
NOR2_X1 U1000 ( .A1(KEYINPUT2), .A2(n1323), .ZN(n1322) );
NAND2_X1 U1001 ( .A1(KEYINPUT44), .A2(n1324), .ZN(n1321) );
XOR2_X1 U1002 ( .A(n1325), .B(n1326), .Z(n1127) );
XOR2_X1 U1003 ( .A(KEYINPUT47), .B(G472), .Z(n1326) );
NAND2_X1 U1004 ( .A1(n1327), .A2(n1204), .ZN(n1325) );
XOR2_X1 U1005 ( .A(n1328), .B(n1193), .Z(n1327) );
XOR2_X1 U1006 ( .A(n1329), .B(G101), .Z(n1193) );
NAND2_X1 U1007 ( .A1(n1330), .A2(G210), .ZN(n1329) );
NAND2_X1 U1008 ( .A1(n1331), .A2(n1332), .ZN(n1328) );
NAND2_X1 U1009 ( .A1(n1198), .A2(n1197), .ZN(n1332) );
XOR2_X1 U1010 ( .A(KEYINPUT35), .B(n1333), .Z(n1331) );
NOR2_X1 U1011 ( .A1(n1198), .A2(n1197), .ZN(n1333) );
XNOR2_X1 U1012 ( .A(G119), .B(n1334), .ZN(n1197) );
XNOR2_X1 U1013 ( .A(G128), .B(n1335), .ZN(n1198) );
NOR3_X1 U1014 ( .A1(n1258), .A2(n1242), .A3(n1078), .ZN(n1283) );
NAND2_X1 U1015 ( .A1(n1118), .A2(n1265), .ZN(n1078) );
NOR2_X1 U1016 ( .A1(n1116), .A2(n1336), .ZN(n1265) );
NOR2_X1 U1017 ( .A1(n1121), .A2(n1122), .ZN(n1336) );
AND2_X1 U1018 ( .A1(n1122), .A2(n1121), .ZN(n1116) );
INV_X1 U1019 ( .A(G475), .ZN(n1121) );
NOR2_X1 U1020 ( .A1(n1179), .A2(G902), .ZN(n1122) );
XNOR2_X1 U1021 ( .A(n1337), .B(n1338), .ZN(n1179) );
XOR2_X1 U1022 ( .A(G131), .B(n1339), .Z(n1338) );
NOR2_X1 U1023 ( .A1(KEYINPUT49), .A2(n1340), .ZN(n1339) );
XOR2_X1 U1024 ( .A(G104), .B(n1341), .Z(n1340) );
XOR2_X1 U1025 ( .A(G122), .B(G113), .Z(n1341) );
XOR2_X1 U1026 ( .A(n1342), .B(n1319), .Z(n1337) );
XOR2_X1 U1027 ( .A(G146), .B(n1134), .Z(n1319) );
XOR2_X1 U1028 ( .A(G125), .B(G140), .Z(n1134) );
NAND2_X1 U1029 ( .A1(KEYINPUT25), .A2(n1343), .ZN(n1342) );
XNOR2_X1 U1030 ( .A(G143), .B(n1344), .ZN(n1343) );
NAND2_X1 U1031 ( .A1(n1330), .A2(G214), .ZN(n1344) );
NOR2_X1 U1032 ( .A1(G953), .A2(G237), .ZN(n1330) );
XOR2_X1 U1033 ( .A(n1345), .B(G478), .Z(n1118) );
NAND2_X1 U1034 ( .A1(n1175), .A2(n1204), .ZN(n1345) );
XNOR2_X1 U1035 ( .A(n1346), .B(n1347), .ZN(n1175) );
XOR2_X1 U1036 ( .A(n1348), .B(n1349), .Z(n1347) );
XOR2_X1 U1037 ( .A(n1350), .B(n1351), .Z(n1349) );
AND3_X1 U1038 ( .A1(G217), .A2(n1090), .A3(G234), .ZN(n1351) );
NAND2_X1 U1039 ( .A1(KEYINPUT24), .A2(G134), .ZN(n1350) );
XOR2_X1 U1040 ( .A(n1352), .B(n1353), .Z(n1346) );
XOR2_X1 U1041 ( .A(G143), .B(G128), .Z(n1353) );
XOR2_X1 U1042 ( .A(G116), .B(n1289), .Z(n1352) );
INV_X1 U1043 ( .A(G122), .ZN(n1289) );
INV_X1 U1044 ( .A(n1282), .ZN(n1242) );
NOR2_X1 U1045 ( .A1(n1105), .A2(n1106), .ZN(n1282) );
INV_X1 U1046 ( .A(n1309), .ZN(n1106) );
NAND2_X1 U1047 ( .A1(G221), .A2(n1313), .ZN(n1309) );
NAND2_X1 U1048 ( .A1(G234), .A2(n1204), .ZN(n1313) );
XOR2_X1 U1049 ( .A(n1354), .B(G469), .Z(n1105) );
NAND2_X1 U1050 ( .A1(n1355), .A2(n1204), .ZN(n1354) );
XOR2_X1 U1051 ( .A(n1212), .B(n1356), .Z(n1355) );
XOR2_X1 U1052 ( .A(KEYINPUT31), .B(n1357), .Z(n1356) );
NOR2_X1 U1053 ( .A1(KEYINPUT11), .A2(n1358), .ZN(n1357) );
XOR2_X1 U1054 ( .A(G140), .B(n1217), .Z(n1358) );
XNOR2_X1 U1055 ( .A(n1324), .B(n1359), .ZN(n1217) );
AND2_X1 U1056 ( .A1(n1090), .A2(G227), .ZN(n1359) );
INV_X1 U1057 ( .A(G110), .ZN(n1324) );
XNOR2_X1 U1058 ( .A(n1161), .B(n1360), .ZN(n1212) );
XOR2_X1 U1059 ( .A(n1335), .B(n1143), .Z(n1360) );
XNOR2_X1 U1060 ( .A(n1361), .B(n1362), .ZN(n1143) );
XOR2_X1 U1061 ( .A(KEYINPUT48), .B(KEYINPUT26), .Z(n1362) );
NAND2_X1 U1062 ( .A1(KEYINPUT0), .A2(n1363), .ZN(n1361) );
XOR2_X1 U1063 ( .A(KEYINPUT59), .B(G128), .Z(n1363) );
XOR2_X1 U1064 ( .A(n1364), .B(n1142), .Z(n1335) );
NAND3_X1 U1065 ( .A1(n1365), .A2(n1366), .A3(n1138), .ZN(n1364) );
NAND3_X1 U1066 ( .A1(G131), .A2(n1267), .A3(G134), .ZN(n1138) );
NAND2_X1 U1067 ( .A1(n1367), .A2(n1368), .ZN(n1366) );
INV_X1 U1068 ( .A(KEYINPUT50), .ZN(n1368) );
XOR2_X1 U1069 ( .A(G131), .B(n1369), .Z(n1367) );
NOR2_X1 U1070 ( .A1(G134), .A2(n1267), .ZN(n1369) );
INV_X1 U1071 ( .A(G137), .ZN(n1267) );
NAND2_X1 U1072 ( .A1(KEYINPUT50), .A2(n1144), .ZN(n1365) );
NAND2_X1 U1073 ( .A1(n1370), .A2(n1371), .ZN(n1144) );
OR3_X1 U1074 ( .A1(G131), .A2(G134), .A3(G137), .ZN(n1371) );
NAND2_X1 U1075 ( .A1(n1372), .A2(G137), .ZN(n1370) );
XOR2_X1 U1076 ( .A(G134), .B(G131), .Z(n1372) );
NAND2_X1 U1077 ( .A1(n1086), .A2(n1373), .ZN(n1258) );
NAND2_X1 U1078 ( .A1(n1071), .A2(n1374), .ZN(n1373) );
NAND4_X1 U1079 ( .A1(G953), .A2(G902), .A3(n1287), .A4(n1159), .ZN(n1374) );
INV_X1 U1080 ( .A(G898), .ZN(n1159) );
NAND3_X1 U1081 ( .A1(n1287), .A2(n1090), .A3(G952), .ZN(n1071) );
NAND2_X1 U1082 ( .A1(G237), .A2(G234), .ZN(n1287) );
INV_X1 U1083 ( .A(n1244), .ZN(n1086) );
NAND2_X1 U1084 ( .A1(n1079), .A2(n1080), .ZN(n1244) );
NAND2_X1 U1085 ( .A1(G214), .A2(n1375), .ZN(n1080) );
INV_X1 U1086 ( .A(n1281), .ZN(n1079) );
XNOR2_X1 U1087 ( .A(n1376), .B(n1228), .ZN(n1281) );
NAND2_X1 U1088 ( .A1(G210), .A2(n1375), .ZN(n1228) );
NAND2_X1 U1089 ( .A1(n1204), .A2(n1377), .ZN(n1375) );
INV_X1 U1090 ( .A(G237), .ZN(n1377) );
NAND2_X1 U1091 ( .A1(n1378), .A2(n1204), .ZN(n1376) );
INV_X1 U1092 ( .A(G902), .ZN(n1204) );
XOR2_X1 U1093 ( .A(n1379), .B(n1224), .Z(n1378) );
NAND2_X1 U1094 ( .A1(n1380), .A2(n1381), .ZN(n1224) );
OR2_X1 U1095 ( .A1(n1160), .A2(n1161), .ZN(n1381) );
NAND2_X1 U1096 ( .A1(n1382), .A2(n1161), .ZN(n1380) );
XNOR2_X1 U1097 ( .A(n1383), .B(n1384), .ZN(n1161) );
INV_X1 U1098 ( .A(n1348), .ZN(n1384) );
XNOR2_X1 U1099 ( .A(G107), .B(KEYINPUT20), .ZN(n1348) );
XOR2_X1 U1100 ( .A(G101), .B(n1184), .Z(n1383) );
INV_X1 U1101 ( .A(G104), .ZN(n1184) );
XOR2_X1 U1102 ( .A(n1160), .B(KEYINPUT9), .Z(n1382) );
XOR2_X1 U1103 ( .A(n1385), .B(n1386), .Z(n1160) );
XOR2_X1 U1104 ( .A(G122), .B(G110), .Z(n1386) );
NAND2_X1 U1105 ( .A1(n1387), .A2(n1388), .ZN(n1385) );
NAND2_X1 U1106 ( .A1(n1389), .A2(n1323), .ZN(n1388) );
INV_X1 U1107 ( .A(G119), .ZN(n1323) );
XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1334), .Z(n1389) );
NAND2_X1 U1109 ( .A1(n1334), .A2(G119), .ZN(n1387) );
XOR2_X1 U1110 ( .A(G116), .B(G113), .Z(n1334) );
NAND2_X1 U1111 ( .A1(n1390), .A2(n1391), .ZN(n1379) );
NAND2_X1 U1112 ( .A1(n1223), .A2(n1227), .ZN(n1391) );
XOR2_X1 U1113 ( .A(n1392), .B(KEYINPUT13), .Z(n1390) );
OR2_X1 U1114 ( .A1(n1227), .A2(n1223), .ZN(n1392) );
XOR2_X1 U1115 ( .A(n1393), .B(n1142), .Z(n1223) );
XNOR2_X1 U1116 ( .A(G146), .B(G143), .ZN(n1142) );
XNOR2_X1 U1117 ( .A(G125), .B(G128), .ZN(n1393) );
NAND2_X1 U1118 ( .A1(G224), .A2(n1090), .ZN(n1227) );
INV_X1 U1119 ( .A(G953), .ZN(n1090) );
endmodule


