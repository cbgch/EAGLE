//Key = 0101101001000011101010000100100111101011101001101101110001100010


module b04_C ( RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN, U344,
U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333, U332,
U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321, U320,
U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309, U308,
U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297, U296,
U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285, U284,
U283, U282, U281, U280, U375, KEYINPUT0, KEYINPUT1, KEYINPUT2,
KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63 );
input RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21,
KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63;
output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323,
U322, U321, U320, U319, U318, U317, U316, U315, U314, U313, U312,
U311, U310, U309, U308, U307, U306, U305, U304, U303, U302, U301,
U300, U299, U298, U297, U296, U295, U294, U293, U292, U291, U290,
U289, U288, U287, U286, U285, U284, U283, U282, U281, U280, U375;
wire   n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
n2335;

INV_X2 U1305 ( .A(n1910), .ZN(n1901) );
INV_X2 U1306 ( .A(U280), .ZN(n1902) );
NAND2_X1 U1307 ( .A1(n1755), .A2(n1756), .ZN(U344) );
NAND2_X1 U1308 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1757), .ZN(n1756) );
NAND2_X1 U1309 ( .A1(DATA_IN_7_), .A2(n1758), .ZN(n1755) );
NAND2_X1 U1310 ( .A1(n1759), .A2(n1760), .ZN(U343) );
NAND2_X1 U1311 ( .A1(n1761), .A2(n1757), .ZN(n1760) );
XOR2_X1 U1312 ( .A(RMAX_REG_6__SCAN_IN), .B(KEYINPUT24), .Z(n1761) );
NAND2_X1 U1313 ( .A1(DATA_IN_6_), .A2(n1758), .ZN(n1759) );
NAND2_X1 U1314 ( .A1(n1762), .A2(n1763), .ZN(U342) );
NAND2_X1 U1315 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1757), .ZN(n1763) );
NAND2_X1 U1316 ( .A1(DATA_IN_5_), .A2(n1758), .ZN(n1762) );
NAND2_X1 U1317 ( .A1(n1764), .A2(n1765), .ZN(U341) );
NAND2_X1 U1318 ( .A1(n1766), .A2(n1757), .ZN(n1765) );
XOR2_X1 U1319 ( .A(n1767), .B(KEYINPUT39), .Z(n1766) );
NAND2_X1 U1320 ( .A1(DATA_IN_4_), .A2(n1758), .ZN(n1764) );
NAND2_X1 U1321 ( .A1(n1768), .A2(n1769), .ZN(U340) );
NAND2_X1 U1322 ( .A1(n1770), .A2(n1757), .ZN(n1769) );
XOR2_X1 U1323 ( .A(n1771), .B(KEYINPUT42), .Z(n1770) );
NAND2_X1 U1324 ( .A1(DATA_IN_3_), .A2(n1758), .ZN(n1768) );
NAND2_X1 U1325 ( .A1(n1772), .A2(n1773), .ZN(U339) );
NAND2_X1 U1326 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1757), .ZN(n1773) );
NAND2_X1 U1327 ( .A1(DATA_IN_2_), .A2(n1758), .ZN(n1772) );
NAND2_X1 U1328 ( .A1(n1774), .A2(n1775), .ZN(U338) );
NAND2_X1 U1329 ( .A1(RMAX_REG_1__SCAN_IN), .A2(n1776), .ZN(n1775) );
XNOR2_X1 U1330 ( .A(KEYINPUT25), .B(n1757), .ZN(n1776) );
NAND2_X1 U1331 ( .A1(DATA_IN_1_), .A2(n1758), .ZN(n1774) );
NAND2_X1 U1332 ( .A1(n1777), .A2(n1778), .ZN(U337) );
NAND2_X1 U1333 ( .A1(RMAX_REG_0__SCAN_IN), .A2(n1757), .ZN(n1778) );
NAND2_X1 U1334 ( .A1(n1779), .A2(n1780), .ZN(n1757) );
NAND2_X1 U1335 ( .A1(n1781), .A2(n1782), .ZN(n1780) );
NAND2_X1 U1336 ( .A1(DATA_IN_0_), .A2(n1758), .ZN(n1777) );
NAND2_X1 U1337 ( .A1(n1782), .A2(n1783), .ZN(n1758) );
NAND2_X1 U1338 ( .A1(n1784), .A2(n1785), .ZN(n1783) );
XNOR2_X1 U1339 ( .A(STATO_REG_1__SCAN_IN), .B(KEYINPUT33), .ZN(n1784) );
NAND2_X1 U1340 ( .A1(n1786), .A2(n1787), .ZN(U336) );
NAND2_X1 U1341 ( .A1(n1788), .A2(DATA_IN_7_), .ZN(n1787) );
NAND2_X1 U1342 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1789), .ZN(n1786) );
NAND2_X1 U1343 ( .A1(n1790), .A2(n1791), .ZN(U335) );
NAND2_X1 U1344 ( .A1(n1788), .A2(DATA_IN_6_), .ZN(n1791) );
NAND2_X1 U1345 ( .A1(RMIN_REG_6__SCAN_IN), .A2(n1789), .ZN(n1790) );
NAND2_X1 U1346 ( .A1(n1792), .A2(n1793), .ZN(U334) );
NAND2_X1 U1347 ( .A1(n1788), .A2(DATA_IN_5_), .ZN(n1793) );
NAND2_X1 U1348 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1789), .ZN(n1792) );
NAND2_X1 U1349 ( .A1(n1794), .A2(n1795), .ZN(U333) );
NAND2_X1 U1350 ( .A1(n1788), .A2(DATA_IN_4_), .ZN(n1795) );
NAND2_X1 U1351 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1789), .ZN(n1794) );
NAND2_X1 U1352 ( .A1(n1796), .A2(n1797), .ZN(U332) );
NAND2_X1 U1353 ( .A1(n1788), .A2(DATA_IN_3_), .ZN(n1797) );
NAND2_X1 U1354 ( .A1(RMIN_REG_3__SCAN_IN), .A2(n1789), .ZN(n1796) );
NAND2_X1 U1355 ( .A1(n1798), .A2(n1799), .ZN(U331) );
NAND2_X1 U1356 ( .A1(n1788), .A2(DATA_IN_2_), .ZN(n1799) );
NAND2_X1 U1357 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1789), .ZN(n1798) );
NAND2_X1 U1358 ( .A1(n1800), .A2(n1801), .ZN(U330) );
NAND2_X1 U1359 ( .A1(n1788), .A2(DATA_IN_1_), .ZN(n1801) );
NAND2_X1 U1360 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1789), .ZN(n1800) );
NAND2_X1 U1361 ( .A1(n1802), .A2(n1803), .ZN(U329) );
NAND2_X1 U1362 ( .A1(n1788), .A2(DATA_IN_0_), .ZN(n1803) );
AND2_X1 U1363 ( .A1(n1804), .A2(n1779), .ZN(n1788) );
NAND2_X1 U1364 ( .A1(n1782), .A2(n1805), .ZN(n1804) );
NAND2_X1 U1365 ( .A1(RMIN_REG_0__SCAN_IN), .A2(n1789), .ZN(n1802) );
NAND2_X1 U1366 ( .A1(n1779), .A2(n1806), .ZN(n1789) );
NAND2_X1 U1367 ( .A1(n1807), .A2(n1805), .ZN(n1806) );
NAND2_X1 U1368 ( .A1(n1781), .A2(n1808), .ZN(n1805) );
NAND2_X1 U1369 ( .A1(n1809), .A2(n1810), .ZN(n1808) );
NAND3_X1 U1370 ( .A1(n1811), .A2(n1812), .A3(n1813), .ZN(n1810) );
NAND2_X1 U1371 ( .A1(RMIN_REG_7__SCAN_IN), .A2(n1814), .ZN(n1813) );
NAND3_X1 U1372 ( .A1(n1815), .A2(n1816), .A3(n1817), .ZN(n1812) );
NAND2_X1 U1373 ( .A1(RMIN_REG_5__SCAN_IN), .A2(n1818), .ZN(n1817) );
NAND3_X1 U1374 ( .A1(n1819), .A2(n1820), .A3(n1821), .ZN(n1816) );
NAND2_X1 U1375 ( .A1(DATA_IN_4_), .A2(n1822), .ZN(n1821) );
NAND3_X1 U1376 ( .A1(n1823), .A2(n1824), .A3(n1825), .ZN(n1820) );
NAND2_X1 U1377 ( .A1(RMIN_REG_4__SCAN_IN), .A2(n1826), .ZN(n1825) );
NAND3_X1 U1378 ( .A1(n1827), .A2(n1828), .A3(n1829), .ZN(n1824) );
NAND2_X1 U1379 ( .A1(DATA_IN_3_), .A2(n1830), .ZN(n1829) );
NAND3_X1 U1380 ( .A1(n1831), .A2(n1832), .A3(n1833), .ZN(n1828) );
NAND2_X1 U1381 ( .A1(RMIN_REG_2__SCAN_IN), .A2(n1834), .ZN(n1833) );
NAND3_X1 U1382 ( .A1(n1835), .A2(n1836), .A3(RMIN_REG_0__SCAN_IN), .ZN(n1832) );
INV_X1 U1383 ( .A(DATA_IN_0_), .ZN(n1836) );
NAND2_X1 U1384 ( .A1(DATA_IN_1_), .A2(n1837), .ZN(n1835) );
NAND2_X1 U1385 ( .A1(RMIN_REG_1__SCAN_IN), .A2(n1838), .ZN(n1831) );
NAND2_X1 U1386 ( .A1(DATA_IN_2_), .A2(n1839), .ZN(n1827) );
NAND2_X1 U1387 ( .A1(n1840), .A2(RMIN_REG_3__SCAN_IN), .ZN(n1823) );
XOR2_X1 U1388 ( .A(n1841), .B(KEYINPUT26), .Z(n1840) );
NAND2_X1 U1389 ( .A1(n1842), .A2(DATA_IN_5_), .ZN(n1819) );
XOR2_X1 U1390 ( .A(n1843), .B(KEYINPUT59), .Z(n1842) );
NAND2_X1 U1391 ( .A1(n1844), .A2(RMIN_REG_6__SCAN_IN), .ZN(n1815) );
XOR2_X1 U1392 ( .A(n1845), .B(KEYINPUT10), .Z(n1844) );
NAND2_X1 U1393 ( .A1(DATA_IN_6_), .A2(n1846), .ZN(n1811) );
NAND2_X1 U1394 ( .A1(DATA_IN_7_), .A2(n1847), .ZN(n1809) );
INV_X1 U1395 ( .A(n1785), .ZN(n1781) );
NAND2_X1 U1396 ( .A1(n1848), .A2(n1849), .ZN(n1785) );
NAND2_X1 U1397 ( .A1(RMAX_REG_7__SCAN_IN), .A2(n1814), .ZN(n1849) );
INV_X1 U1398 ( .A(DATA_IN_7_), .ZN(n1814) );
NAND3_X1 U1399 ( .A1(n1850), .A2(n1851), .A3(n1852), .ZN(n1848) );
NAND2_X1 U1400 ( .A1(DATA_IN_7_), .A2(n1853), .ZN(n1852) );
NAND3_X1 U1401 ( .A1(n1854), .A2(n1855), .A3(n1856), .ZN(n1851) );
NAND2_X1 U1402 ( .A1(DATA_IN_6_), .A2(n1857), .ZN(n1856) );
NAND3_X1 U1403 ( .A1(n1858), .A2(n1859), .A3(n1860), .ZN(n1855) );
NAND2_X1 U1404 ( .A1(RMAX_REG_5__SCAN_IN), .A2(n1818), .ZN(n1860) );
NAND3_X1 U1405 ( .A1(n1861), .A2(n1862), .A3(n1863), .ZN(n1859) );
NAND2_X1 U1406 ( .A1(DATA_IN_4_), .A2(n1767), .ZN(n1863) );
NAND3_X1 U1407 ( .A1(n1864), .A2(n1865), .A3(n1866), .ZN(n1862) );
NAND2_X1 U1408 ( .A1(RMAX_REG_2__SCAN_IN), .A2(n1834), .ZN(n1866) );
NAND3_X1 U1409 ( .A1(n1867), .A2(n1868), .A3(n1869), .ZN(n1865) );
NAND2_X1 U1410 ( .A1(DATA_IN_2_), .A2(n1870), .ZN(n1869) );
NAND3_X1 U1411 ( .A1(n1871), .A2(n1872), .A3(DATA_IN_0_), .ZN(n1868) );
NAND2_X1 U1412 ( .A1(n1873), .A2(RMAX_REG_1__SCAN_IN), .ZN(n1871) );
XOR2_X1 U1413 ( .A(n1838), .B(KEYINPUT43), .Z(n1873) );
NAND2_X1 U1414 ( .A1(DATA_IN_1_), .A2(n1874), .ZN(n1867) );
NAND2_X1 U1415 ( .A1(n1875), .A2(n1841), .ZN(n1864) );
XOR2_X1 U1416 ( .A(RMAX_REG_3__SCAN_IN), .B(KEYINPUT47), .Z(n1875) );
NAND2_X1 U1417 ( .A1(DATA_IN_3_), .A2(n1771), .ZN(n1861) );
NAND2_X1 U1418 ( .A1(RMAX_REG_4__SCAN_IN), .A2(n1826), .ZN(n1858) );
NAND2_X1 U1419 ( .A1(DATA_IN_5_), .A2(n1876), .ZN(n1854) );
NAND2_X1 U1420 ( .A1(RMAX_REG_6__SCAN_IN), .A2(n1845), .ZN(n1850) );
XOR2_X1 U1421 ( .A(n1782), .B(KEYINPUT44), .Z(n1807) );
NAND2_X1 U1422 ( .A1(n1877), .A2(n1878), .ZN(U328) );
NAND2_X1 U1423 ( .A1(n1879), .A2(DATA_IN_7_), .ZN(n1878) );
NAND2_X1 U1424 ( .A1(RLAST_REG_7__SCAN_IN), .A2(n1880), .ZN(n1877) );
NAND2_X1 U1425 ( .A1(n1881), .A2(n1882), .ZN(U327) );
NAND2_X1 U1426 ( .A1(n1879), .A2(DATA_IN_6_), .ZN(n1882) );
NAND2_X1 U1427 ( .A1(RLAST_REG_6__SCAN_IN), .A2(n1880), .ZN(n1881) );
NAND2_X1 U1428 ( .A1(n1883), .A2(n1884), .ZN(U326) );
NAND2_X1 U1429 ( .A1(n1879), .A2(DATA_IN_5_), .ZN(n1884) );
NAND2_X1 U1430 ( .A1(RLAST_REG_5__SCAN_IN), .A2(n1880), .ZN(n1883) );
NAND2_X1 U1431 ( .A1(n1885), .A2(n1886), .ZN(U325) );
NAND2_X1 U1432 ( .A1(n1879), .A2(DATA_IN_4_), .ZN(n1886) );
NAND2_X1 U1433 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n1880), .ZN(n1885) );
NAND2_X1 U1434 ( .A1(n1887), .A2(n1888), .ZN(U324) );
NAND2_X1 U1435 ( .A1(n1879), .A2(DATA_IN_3_), .ZN(n1888) );
NAND2_X1 U1436 ( .A1(RLAST_REG_3__SCAN_IN), .A2(n1880), .ZN(n1887) );
NAND2_X1 U1437 ( .A1(n1889), .A2(n1890), .ZN(U323) );
NAND2_X1 U1438 ( .A1(RLAST_REG_2__SCAN_IN), .A2(n1880), .ZN(n1890) );
XOR2_X1 U1439 ( .A(KEYINPUT18), .B(n1891), .Z(n1889) );
NOR2_X1 U1440 ( .A1(n1834), .A2(n1892), .ZN(n1891) );
NAND2_X1 U1441 ( .A1(n1893), .A2(n1894), .ZN(U322) );
NAND2_X1 U1442 ( .A1(n1879), .A2(DATA_IN_1_), .ZN(n1894) );
NAND2_X1 U1443 ( .A1(RLAST_REG_1__SCAN_IN), .A2(n1880), .ZN(n1893) );
NAND2_X1 U1444 ( .A1(n1895), .A2(n1896), .ZN(U321) );
NAND2_X1 U1445 ( .A1(n1879), .A2(DATA_IN_0_), .ZN(n1896) );
INV_X1 U1446 ( .A(n1892), .ZN(n1879) );
NAND2_X1 U1447 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1897), .ZN(n1892) );
NAND2_X1 U1448 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n1880), .ZN(n1895) );
NAND2_X1 U1449 ( .A1(n1779), .A2(n1897), .ZN(n1880) );
NAND2_X1 U1450 ( .A1(n1898), .A2(n1782), .ZN(n1897) );
INV_X1 U1451 ( .A(U375), .ZN(n1779) );
NOR2_X1 U1452 ( .A1(STATO_REG_0__SCAN_IN), .A2(STATO_REG_1__SCAN_IN), .ZN(U375) );
NAND2_X1 U1453 ( .A1(n1899), .A2(n1900), .ZN(U320) );
NAND2_X1 U1454 ( .A1(n1901), .A2(DATA_IN_7_), .ZN(n1900) );
NAND2_X1 U1455 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1902), .ZN(n1899) );
NAND2_X1 U1456 ( .A1(n1903), .A2(n1904), .ZN(U319) );
NAND2_X1 U1457 ( .A1(n1901), .A2(DATA_IN_6_), .ZN(n1904) );
NAND2_X1 U1458 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1902), .ZN(n1903) );
NAND2_X1 U1459 ( .A1(n1905), .A2(n1906), .ZN(U318) );
NAND2_X1 U1460 ( .A1(n1901), .A2(DATA_IN_5_), .ZN(n1906) );
NAND2_X1 U1461 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1902), .ZN(n1905) );
NAND2_X1 U1462 ( .A1(n1907), .A2(n1908), .ZN(U317) );
NAND2_X1 U1463 ( .A1(n1909), .A2(DATA_IN_4_), .ZN(n1908) );
XOR2_X1 U1464 ( .A(n1910), .B(KEYINPUT1), .Z(n1909) );
NAND2_X1 U1465 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1902), .ZN(n1907) );
NAND2_X1 U1466 ( .A1(n1911), .A2(n1912), .ZN(U316) );
NAND2_X1 U1467 ( .A1(n1901), .A2(DATA_IN_3_), .ZN(n1912) );
NAND2_X1 U1468 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1902), .ZN(n1911) );
NAND2_X1 U1469 ( .A1(n1913), .A2(n1914), .ZN(U315) );
NAND2_X1 U1470 ( .A1(n1901), .A2(n1915), .ZN(n1914) );
XOR2_X1 U1471 ( .A(KEYINPUT41), .B(DATA_IN_2_), .Z(n1915) );
NAND2_X1 U1472 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1902), .ZN(n1913) );
NAND2_X1 U1473 ( .A1(n1916), .A2(n1917), .ZN(U314) );
NAND2_X1 U1474 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1902), .ZN(n1917) );
XOR2_X1 U1475 ( .A(KEYINPUT57), .B(n1918), .Z(n1916) );
NOR2_X1 U1476 ( .A1(n1838), .A2(n1910), .ZN(n1918) );
NAND2_X1 U1477 ( .A1(n1919), .A2(n1920), .ZN(U313) );
NAND2_X1 U1478 ( .A1(n1901), .A2(DATA_IN_0_), .ZN(n1920) );
NAND2_X1 U1479 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1902), .ZN(n1919) );
NAND2_X1 U1480 ( .A1(n1921), .A2(n1922), .ZN(U312) );
NAND2_X1 U1481 ( .A1(REG1_REG_7__SCAN_IN), .A2(n1901), .ZN(n1922) );
NAND2_X1 U1482 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1902), .ZN(n1921) );
NAND2_X1 U1483 ( .A1(n1923), .A2(n1924), .ZN(U311) );
NAND2_X1 U1484 ( .A1(REG1_REG_6__SCAN_IN), .A2(n1901), .ZN(n1924) );
NAND2_X1 U1485 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1902), .ZN(n1923) );
NAND2_X1 U1486 ( .A1(n1925), .A2(n1926), .ZN(U310) );
NAND2_X1 U1487 ( .A1(REG1_REG_5__SCAN_IN), .A2(n1901), .ZN(n1926) );
NAND2_X1 U1488 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1902), .ZN(n1925) );
NAND2_X1 U1489 ( .A1(n1927), .A2(n1928), .ZN(U309) );
NAND2_X1 U1490 ( .A1(REG1_REG_4__SCAN_IN), .A2(n1901), .ZN(n1928) );
NAND2_X1 U1491 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1902), .ZN(n1927) );
NAND2_X1 U1492 ( .A1(n1929), .A2(n1930), .ZN(U308) );
NAND2_X1 U1493 ( .A1(REG1_REG_3__SCAN_IN), .A2(n1901), .ZN(n1930) );
NAND2_X1 U1494 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1902), .ZN(n1929) );
NAND2_X1 U1495 ( .A1(n1931), .A2(n1932), .ZN(U307) );
NAND2_X1 U1496 ( .A1(REG1_REG_2__SCAN_IN), .A2(n1901), .ZN(n1932) );
XOR2_X1 U1497 ( .A(KEYINPUT49), .B(n1933), .Z(n1931) );
AND2_X1 U1498 ( .A1(n1902), .A2(REG2_REG_2__SCAN_IN), .ZN(n1933) );
NAND2_X1 U1499 ( .A1(n1934), .A2(n1935), .ZN(U306) );
NAND2_X1 U1500 ( .A1(REG1_REG_1__SCAN_IN), .A2(n1901), .ZN(n1935) );
NAND2_X1 U1501 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1902), .ZN(n1934) );
NAND2_X1 U1502 ( .A1(n1936), .A2(n1937), .ZN(U305) );
NAND2_X1 U1503 ( .A1(REG1_REG_0__SCAN_IN), .A2(n1901), .ZN(n1937) );
NAND2_X1 U1504 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1902), .ZN(n1936) );
NAND2_X1 U1505 ( .A1(n1938), .A2(n1939), .ZN(U304) );
NAND2_X1 U1506 ( .A1(REG2_REG_7__SCAN_IN), .A2(n1901), .ZN(n1939) );
NAND2_X1 U1507 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1902), .ZN(n1938) );
NAND2_X1 U1508 ( .A1(n1940), .A2(n1941), .ZN(U303) );
NAND2_X1 U1509 ( .A1(REG2_REG_6__SCAN_IN), .A2(n1901), .ZN(n1941) );
NAND2_X1 U1510 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1902), .ZN(n1940) );
NAND2_X1 U1511 ( .A1(n1942), .A2(n1943), .ZN(U302) );
NAND2_X1 U1512 ( .A1(REG2_REG_5__SCAN_IN), .A2(n1901), .ZN(n1943) );
NAND2_X1 U1513 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1902), .ZN(n1942) );
NAND2_X1 U1514 ( .A1(n1944), .A2(n1945), .ZN(U301) );
NAND2_X1 U1515 ( .A1(REG2_REG_4__SCAN_IN), .A2(n1901), .ZN(n1945) );
NAND2_X1 U1516 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1902), .ZN(n1944) );
NAND2_X1 U1517 ( .A1(n1946), .A2(n1947), .ZN(U300) );
NAND2_X1 U1518 ( .A1(REG2_REG_3__SCAN_IN), .A2(n1901), .ZN(n1947) );
NAND2_X1 U1519 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1902), .ZN(n1946) );
NAND2_X1 U1520 ( .A1(n1948), .A2(n1949), .ZN(U299) );
NAND2_X1 U1521 ( .A1(REG2_REG_2__SCAN_IN), .A2(n1901), .ZN(n1949) );
NAND2_X1 U1522 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1902), .ZN(n1948) );
NAND2_X1 U1523 ( .A1(n1950), .A2(n1951), .ZN(U298) );
NAND2_X1 U1524 ( .A1(REG2_REG_1__SCAN_IN), .A2(n1901), .ZN(n1951) );
NAND2_X1 U1525 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1902), .ZN(n1950) );
NAND2_X1 U1526 ( .A1(n1952), .A2(n1953), .ZN(U297) );
NAND2_X1 U1527 ( .A1(REG2_REG_0__SCAN_IN), .A2(n1901), .ZN(n1953) );
NAND2_X1 U1528 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1902), .ZN(n1952) );
NAND2_X1 U1529 ( .A1(n1954), .A2(n1955), .ZN(U296) );
NAND2_X1 U1530 ( .A1(REG3_REG_7__SCAN_IN), .A2(n1901), .ZN(n1955) );
NAND2_X1 U1531 ( .A1(REG4_REG_7__SCAN_IN), .A2(n1902), .ZN(n1954) );
NAND2_X1 U1532 ( .A1(n1956), .A2(n1957), .ZN(U295) );
NAND2_X1 U1533 ( .A1(REG3_REG_6__SCAN_IN), .A2(n1901), .ZN(n1957) );
NAND2_X1 U1534 ( .A1(REG4_REG_6__SCAN_IN), .A2(n1902), .ZN(n1956) );
NAND2_X1 U1535 ( .A1(n1958), .A2(n1959), .ZN(U294) );
NAND2_X1 U1536 ( .A1(REG3_REG_5__SCAN_IN), .A2(n1901), .ZN(n1959) );
NAND2_X1 U1537 ( .A1(REG4_REG_5__SCAN_IN), .A2(n1902), .ZN(n1958) );
NAND2_X1 U1538 ( .A1(n1960), .A2(n1961), .ZN(U293) );
NAND2_X1 U1539 ( .A1(n1962), .A2(n1902), .ZN(n1961) );
XOR2_X1 U1540 ( .A(n1963), .B(KEYINPUT34), .Z(n1962) );
NAND2_X1 U1541 ( .A1(REG3_REG_4__SCAN_IN), .A2(n1901), .ZN(n1960) );
NAND2_X1 U1542 ( .A1(n1964), .A2(n1965), .ZN(U292) );
NAND2_X1 U1543 ( .A1(REG3_REG_3__SCAN_IN), .A2(n1901), .ZN(n1965) );
NAND2_X1 U1544 ( .A1(REG4_REG_3__SCAN_IN), .A2(n1902), .ZN(n1964) );
NAND2_X1 U1545 ( .A1(n1966), .A2(n1967), .ZN(U291) );
NAND2_X1 U1546 ( .A1(REG3_REG_2__SCAN_IN), .A2(n1901), .ZN(n1967) );
NAND2_X1 U1547 ( .A1(REG4_REG_2__SCAN_IN), .A2(n1902), .ZN(n1966) );
NAND2_X1 U1548 ( .A1(n1968), .A2(n1969), .ZN(U290) );
NAND2_X1 U1549 ( .A1(REG3_REG_1__SCAN_IN), .A2(n1901), .ZN(n1969) );
NAND2_X1 U1550 ( .A1(REG4_REG_1__SCAN_IN), .A2(n1902), .ZN(n1968) );
NAND2_X1 U1551 ( .A1(n1970), .A2(n1971), .ZN(U289) );
NAND2_X1 U1552 ( .A1(REG3_REG_0__SCAN_IN), .A2(n1901), .ZN(n1971) );
NAND2_X1 U1553 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1902), .ZN(n1970) );
NAND4_X1 U1554 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .ZN(U288));
NAND2_X1 U1555 ( .A1(n1976), .A2(n1977), .ZN(n1975) );
XOR2_X1 U1556 ( .A(KEYINPUT55), .B(n1978), .Z(n1977) );
NOR2_X1 U1557 ( .A1(n1979), .A2(n1980), .ZN(n1974) );
NOR2_X1 U1558 ( .A1(n1981), .A2(n1982), .ZN(n1980) );
XNOR2_X1 U1559 ( .A(RLAST_REG_7__SCAN_IN), .B(KEYINPUT27), .ZN(n1981) );
NAND2_X1 U1560 ( .A1(n1983), .A2(REG4_REG_7__SCAN_IN), .ZN(n1973) );
NAND2_X1 U1561 ( .A1(DATA_OUT_REG_7__SCAN_IN), .A2(n1902), .ZN(n1972) );
NAND4_X1 U1562 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .ZN(U287));
NOR3_X1 U1563 ( .A1(n1988), .A2(n1979), .A3(n1989), .ZN(n1987) );
NOR3_X1 U1564 ( .A1(n1990), .A2(n1991), .A3(n1992), .ZN(n1989) );
AND3_X1 U1565 ( .A1(n1991), .A2(n1990), .A3(n1993), .ZN(n1979) );
NAND2_X1 U1566 ( .A1(n1994), .A2(n1995), .ZN(n1990) );
AND2_X1 U1567 ( .A1(n1996), .A2(n1997), .ZN(n1991) );
NOR2_X1 U1568 ( .A1(n1998), .A2(n1999), .ZN(n1988) );
NOR2_X1 U1569 ( .A1(n2000), .A2(n1978), .ZN(n1998) );
AND3_X1 U1570 ( .A1(n2001), .A2(n1997), .A3(n2002), .ZN(n1978) );
NOR2_X1 U1571 ( .A1(n1997), .A2(n2001), .ZN(n2000) );
NAND2_X1 U1572 ( .A1(n2003), .A2(n2004), .ZN(n2001) );
NAND2_X1 U1573 ( .A1(n1983), .A2(REG4_REG_6__SCAN_IN), .ZN(n1986) );
NAND2_X1 U1574 ( .A1(DATA_OUT_REG_6__SCAN_IN), .A2(n2005), .ZN(n1985) );
XOR2_X1 U1575 ( .A(KEYINPUT19), .B(n1902), .Z(n2005) );
NAND2_X1 U1576 ( .A1(n2006), .A2(RLAST_REG_6__SCAN_IN), .ZN(n1984) );
NAND4_X1 U1577 ( .A1(n2007), .A2(n2008), .A3(n2009), .A4(n2010), .ZN(U286));
NOR3_X1 U1578 ( .A1(n2011), .A2(n2012), .A3(n2013), .ZN(n2010) );
NOR2_X1 U1579 ( .A1(n1999), .A2(n2014), .ZN(n2013) );
XNOR2_X1 U1580 ( .A(n2015), .B(n2004), .ZN(n2014) );
XNOR2_X1 U1581 ( .A(n1997), .B(n2016), .ZN(n2004) );
NOR2_X1 U1582 ( .A1(KEYINPUT13), .A2(n2017), .ZN(n2016) );
NAND2_X1 U1583 ( .A1(KEYINPUT20), .A2(n2018), .ZN(n2015) );
NOR2_X1 U1584 ( .A1(n1992), .A2(n2019), .ZN(n2012) );
XNOR2_X1 U1585 ( .A(n2020), .B(n1995), .ZN(n2019) );
XNOR2_X1 U1586 ( .A(n1997), .B(n1996), .ZN(n1995) );
NAND2_X1 U1587 ( .A1(KEYINPUT53), .A2(n2021), .ZN(n2020) );
INV_X1 U1588 ( .A(n1994), .ZN(n2021) );
NOR2_X1 U1589 ( .A1(n1997), .A2(n2022), .ZN(n2011) );
NAND2_X1 U1590 ( .A1(n2023), .A2(n2024), .ZN(n1997) );
NAND4_X1 U1591 ( .A1(n2025), .A2(n2026), .A3(n2027), .A4(n2028), .ZN(n2024));
NAND2_X1 U1592 ( .A1(n2029), .A2(n2030), .ZN(n2028) );
XOR2_X1 U1593 ( .A(REG4_REG_6__SCAN_IN), .B(DATA_IN_6_), .Z(n2029) );
NAND2_X1 U1594 ( .A1(n2031), .A2(RESTART), .ZN(n2027) );
XOR2_X1 U1595 ( .A(RMIN_REG_6__SCAN_IN), .B(RMAX_REG_6__SCAN_IN), .Z(n2031));
NAND2_X1 U1596 ( .A1(n2032), .A2(n2033), .ZN(n2026) );
XOR2_X1 U1597 ( .A(KEYINPUT7), .B(n2034), .Z(n2032) );
NAND4_X1 U1598 ( .A1(n2035), .A2(n2033), .A3(n2036), .A4(n2037), .ZN(n2023));
NAND2_X1 U1599 ( .A1(n2038), .A2(n2030), .ZN(n2037) );
XOR2_X1 U1600 ( .A(n2039), .B(DATA_IN_6_), .Z(n2038) );
NAND2_X1 U1601 ( .A1(n2040), .A2(RESTART), .ZN(n2036) );
XOR2_X1 U1602 ( .A(n1857), .B(RMIN_REG_6__SCAN_IN), .Z(n2040) );
INV_X1 U1603 ( .A(RMAX_REG_6__SCAN_IN), .ZN(n1857) );
NAND2_X1 U1604 ( .A1(n2041), .A2(n2042), .ZN(n2033) );
NAND2_X1 U1605 ( .A1(n2025), .A2(n2043), .ZN(n2035) );
NAND2_X1 U1606 ( .A1(n2044), .A2(n2045), .ZN(n2025) );
XOR2_X1 U1607 ( .A(KEYINPUT51), .B(n2046), .Z(n2009) );
NOR2_X1 U1608 ( .A1(n2047), .A2(n2048), .ZN(n2046) );
INV_X1 U1609 ( .A(RLAST_REG_5__SCAN_IN), .ZN(n2048) );
XOR2_X1 U1610 ( .A(n1982), .B(KEYINPUT22), .Z(n2047) );
NAND2_X1 U1611 ( .A1(n1983), .A2(REG4_REG_5__SCAN_IN), .ZN(n2008) );
NAND2_X1 U1612 ( .A1(DATA_OUT_REG_5__SCAN_IN), .A2(n1902), .ZN(n2007) );
NAND4_X1 U1613 ( .A1(n2049), .A2(n2050), .A3(n2051), .A4(n2052), .ZN(U285));
NOR3_X1 U1614 ( .A1(n2053), .A2(n2054), .A3(n2055), .ZN(n2052) );
NOR2_X1 U1615 ( .A1(n2056), .A2(n2022), .ZN(n2055) );
NOR3_X1 U1616 ( .A1(n1999), .A2(n2003), .A3(n2057), .ZN(n2054) );
NOR2_X1 U1617 ( .A1(n2058), .A2(n2059), .ZN(n2057) );
NOR2_X1 U1618 ( .A1(n2060), .A2(n2061), .ZN(n2058) );
XNOR2_X1 U1619 ( .A(n2062), .B(KEYINPUT29), .ZN(n2061) );
INV_X1 U1620 ( .A(n2063), .ZN(n2060) );
INV_X1 U1621 ( .A(n2018), .ZN(n2003) );
NAND3_X1 U1622 ( .A1(n2062), .A2(n2063), .A3(n2064), .ZN(n2018) );
XOR2_X1 U1623 ( .A(n2059), .B(KEYINPUT12), .Z(n2064) );
NAND2_X1 U1624 ( .A1(n2017), .A2(n2065), .ZN(n2059) );
NAND2_X1 U1625 ( .A1(n2066), .A2(n2067), .ZN(n2065) );
INV_X1 U1626 ( .A(n2002), .ZN(n2017) );
NOR2_X1 U1627 ( .A1(n2067), .A2(n2066), .ZN(n2002) );
AND2_X1 U1628 ( .A1(RLAST_REG_4__SCAN_IN), .A2(n2006), .ZN(n2053) );
XOR2_X1 U1629 ( .A(KEYINPUT9), .B(n2068), .Z(n2051) );
NOR3_X1 U1630 ( .A1(n1992), .A2(n1994), .A3(n2069), .ZN(n2068) );
NOR3_X1 U1631 ( .A1(n2070), .A2(n1996), .A3(n2071), .ZN(n2069) );
AND2_X1 U1632 ( .A1(n2072), .A2(n2066), .ZN(n2071) );
INV_X1 U1633 ( .A(n2073), .ZN(n1996) );
NOR2_X1 U1634 ( .A1(n2074), .A2(n2075), .ZN(n2070) );
NOR3_X1 U1635 ( .A1(n2074), .A2(n2076), .A3(n2075), .ZN(n1994) );
AND2_X1 U1636 ( .A1(n2077), .A2(n2073), .ZN(n2076) );
NAND2_X1 U1637 ( .A1(n2056), .A2(n2078), .ZN(n2073) );
XNOR2_X1 U1638 ( .A(KEYINPUT11), .B(n2072), .ZN(n2078) );
INV_X1 U1639 ( .A(n2066), .ZN(n2056) );
NAND2_X1 U1640 ( .A1(n2066), .A2(n2072), .ZN(n2077) );
NAND2_X1 U1641 ( .A1(n2079), .A2(n2080), .ZN(n2066) );
NAND2_X1 U1642 ( .A1(n2081), .A2(n2043), .ZN(n2080) );
NAND2_X1 U1643 ( .A1(n2082), .A2(n2083), .ZN(n2081) );
NAND2_X1 U1644 ( .A1(n2045), .A2(n2041), .ZN(n2083) );
INV_X1 U1645 ( .A(n2042), .ZN(n2045) );
XOR2_X1 U1646 ( .A(n2084), .B(KEYINPUT21), .Z(n2082) );
NAND2_X1 U1647 ( .A1(n2034), .A2(n2085), .ZN(n2079) );
NAND3_X1 U1648 ( .A1(n2086), .A2(n2087), .A3(n2088), .ZN(n2085) );
NAND2_X1 U1649 ( .A1(n2042), .A2(n2084), .ZN(n2088) );
NAND2_X1 U1650 ( .A1(n2044), .A2(n2089), .ZN(n2084) );
INV_X1 U1651 ( .A(n2041), .ZN(n2044) );
OR3_X1 U1652 ( .A1(n2041), .A2(n2089), .A3(KEYINPUT56), .ZN(n2087) );
XNOR2_X1 U1653 ( .A(n2042), .B(KEYINPUT14), .ZN(n2089) );
NAND2_X1 U1654 ( .A1(n2090), .A2(n2091), .ZN(n2042) );
NAND2_X1 U1655 ( .A1(RESTART), .A2(n1876), .ZN(n2091) );
NAND2_X1 U1656 ( .A1(n1818), .A2(n2030), .ZN(n2090) );
NAND2_X1 U1657 ( .A1(KEYINPUT56), .A2(n2041), .ZN(n2086) );
NAND2_X1 U1658 ( .A1(n2092), .A2(n2093), .ZN(n2041) );
NAND2_X1 U1659 ( .A1(RESTART), .A2(n1843), .ZN(n2093) );
NAND2_X1 U1660 ( .A1(n2094), .A2(n2030), .ZN(n2092) );
INV_X1 U1661 ( .A(n2043), .ZN(n2034) );
NAND2_X1 U1662 ( .A1(n2095), .A2(n2096), .ZN(n2043) );
NAND2_X1 U1663 ( .A1(n2097), .A2(n2098), .ZN(n2096) );
OR2_X1 U1664 ( .A1(n2099), .A2(n2100), .ZN(n2098) );
NAND2_X1 U1665 ( .A1(n2100), .A2(n2099), .ZN(n2095) );
NAND2_X1 U1666 ( .A1(n1983), .A2(REG4_REG_4__SCAN_IN), .ZN(n2050) );
NAND2_X1 U1667 ( .A1(DATA_OUT_REG_4__SCAN_IN), .A2(n1902), .ZN(n2049) );
NAND4_X1 U1668 ( .A1(n2101), .A2(n2102), .A3(n2103), .A4(n2104), .ZN(U284));
NAND3_X1 U1669 ( .A1(n2105), .A2(n2106), .A3(n1993), .ZN(n2104) );
NAND2_X1 U1670 ( .A1(n2107), .A2(n2108), .ZN(n2106) );
INV_X1 U1671 ( .A(KEYINPUT58), .ZN(n2108) );
NAND2_X1 U1672 ( .A1(n2109), .A2(n2110), .ZN(n2107) );
NAND2_X1 U1673 ( .A1(n2075), .A2(n2111), .ZN(n2110) );
NAND2_X1 U1674 ( .A1(n2074), .A2(n2112), .ZN(n2109) );
XNOR2_X1 U1675 ( .A(n2111), .B(KEYINPUT37), .ZN(n2074) );
NAND2_X1 U1676 ( .A1(n2113), .A2(KEYINPUT58), .ZN(n2105) );
XOR2_X1 U1677 ( .A(n2111), .B(n2114), .Z(n2113) );
OR2_X1 U1678 ( .A1(n2075), .A2(KEYINPUT37), .ZN(n2114) );
NAND2_X1 U1679 ( .A1(n2115), .A2(n2072), .ZN(n2111) );
NAND3_X1 U1680 ( .A1(n2116), .A2(n2117), .A3(n2118), .ZN(n2072) );
XOR2_X1 U1681 ( .A(n2119), .B(KEYINPUT16), .Z(n2116) );
NAND2_X1 U1682 ( .A1(n2119), .A2(n2120), .ZN(n2115) );
NAND2_X1 U1683 ( .A1(n2118), .A2(n2121), .ZN(n2120) );
XOR2_X1 U1684 ( .A(KEYINPUT54), .B(n2117), .Z(n2121) );
NAND2_X1 U1685 ( .A1(n2122), .A2(n1976), .ZN(n2103) );
XOR2_X1 U1686 ( .A(n2063), .B(n2062), .Z(n2122) );
NAND2_X1 U1687 ( .A1(n2067), .A2(n2123), .ZN(n2063) );
NAND2_X1 U1688 ( .A1(n2119), .A2(n2124), .ZN(n2123) );
NAND2_X1 U1689 ( .A1(n2125), .A2(n2126), .ZN(n2067) );
XOR2_X1 U1690 ( .A(KEYINPUT60), .B(n2127), .Z(n2125) );
NAND2_X1 U1691 ( .A1(DATA_OUT_REG_3__SCAN_IN), .A2(n1902), .ZN(n2102) );
XOR2_X1 U1692 ( .A(n2128), .B(KEYINPUT45), .Z(n2101) );
NAND3_X1 U1693 ( .A1(n2129), .A2(n2130), .A3(n2131), .ZN(n2128) );
NAND2_X1 U1694 ( .A1(n1983), .A2(REG4_REG_3__SCAN_IN), .ZN(n2131) );
OR2_X1 U1695 ( .A1(n2022), .A2(n2127), .ZN(n2130) );
INV_X1 U1696 ( .A(n2119), .ZN(n2127) );
NAND2_X1 U1697 ( .A1(n2132), .A2(n2133), .ZN(n2119) );
NAND2_X1 U1698 ( .A1(n2134), .A2(n2135), .ZN(n2133) );
INV_X1 U1699 ( .A(n2100), .ZN(n2135) );
XOR2_X1 U1700 ( .A(n2097), .B(n2136), .Z(n2134) );
XOR2_X1 U1701 ( .A(KEYINPUT63), .B(n2137), .Z(n2136) );
NAND2_X1 U1702 ( .A1(n2138), .A2(n2100), .ZN(n2132) );
NAND2_X1 U1703 ( .A1(n2139), .A2(n2140), .ZN(n2100) );
NAND2_X1 U1704 ( .A1(RESTART), .A2(n1767), .ZN(n2140) );
NAND2_X1 U1705 ( .A1(n1826), .A2(n2030), .ZN(n2139) );
NAND2_X1 U1706 ( .A1(n2141), .A2(n2142), .ZN(n2138) );
NAND2_X1 U1707 ( .A1(n2137), .A2(n2097), .ZN(n2142) );
NOR2_X1 U1708 ( .A1(KEYINPUT50), .A2(n2099), .ZN(n2137) );
NAND2_X1 U1709 ( .A1(n2143), .A2(n2099), .ZN(n2141) );
NAND2_X1 U1710 ( .A1(n2144), .A2(n2145), .ZN(n2099) );
NAND2_X1 U1711 ( .A1(n2146), .A2(n2147), .ZN(n2145) );
OR2_X1 U1712 ( .A1(n2148), .A2(n2149), .ZN(n2146) );
NAND2_X1 U1713 ( .A1(n2149), .A2(n2148), .ZN(n2144) );
INV_X1 U1714 ( .A(n2097), .ZN(n2143) );
NAND2_X1 U1715 ( .A1(n2150), .A2(n2151), .ZN(n2097) );
NAND2_X1 U1716 ( .A1(RESTART), .A2(n1822), .ZN(n2151) );
NAND2_X1 U1717 ( .A1(n1963), .A2(n2030), .ZN(n2150) );
NAND2_X1 U1718 ( .A1(n2006), .A2(RLAST_REG_3__SCAN_IN), .ZN(n2129) );
NAND4_X1 U1719 ( .A1(n2152), .A2(n2153), .A3(n2154), .A4(n2155), .ZN(U283));
NOR3_X1 U1720 ( .A1(n2156), .A2(n2157), .A3(n2158), .ZN(n2155) );
NOR3_X1 U1721 ( .A1(n1992), .A2(n2112), .A3(n2159), .ZN(n2158) );
NOR3_X1 U1722 ( .A1(n2117), .A2(n2160), .A3(n2161), .ZN(n2159) );
NOR2_X1 U1723 ( .A1(n2162), .A2(n2163), .ZN(n2160) );
INV_X1 U1724 ( .A(n2164), .ZN(n2117) );
INV_X1 U1725 ( .A(n2075), .ZN(n2112) );
NAND4_X1 U1726 ( .A1(n2165), .A2(n2166), .A3(n2167), .A4(n2168), .ZN(n2075));
OR2_X1 U1727 ( .A1(n2169), .A2(n2118), .ZN(n2168) );
NAND2_X1 U1728 ( .A1(n2118), .A2(n2164), .ZN(n2167) );
XOR2_X1 U1729 ( .A(n2169), .B(KEYINPUT5), .Z(n2164) );
INV_X1 U1730 ( .A(n2163), .ZN(n2165) );
NOR3_X1 U1731 ( .A1(n1999), .A2(n2062), .A3(n2170), .ZN(n2157) );
NOR2_X1 U1732 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
NOR2_X1 U1733 ( .A1(n2162), .A2(n2173), .ZN(n2171) );
NOR3_X1 U1734 ( .A1(n2174), .A2(n2162), .A3(n2173), .ZN(n2062) );
INV_X1 U1735 ( .A(n2172), .ZN(n2174) );
NAND2_X1 U1736 ( .A1(n2124), .A2(n2175), .ZN(n2172) );
NAND2_X1 U1737 ( .A1(n2161), .A2(n2169), .ZN(n2175) );
INV_X1 U1738 ( .A(n2126), .ZN(n2124) );
NOR2_X1 U1739 ( .A1(n2161), .A2(n2169), .ZN(n2126) );
INV_X1 U1740 ( .A(n2118), .ZN(n2161) );
NOR2_X1 U1741 ( .A1(n2118), .A2(n2022), .ZN(n2156) );
XOR2_X1 U1742 ( .A(n2148), .B(n2176), .Z(n2118) );
XOR2_X1 U1743 ( .A(n2147), .B(n2149), .Z(n2176) );
NAND2_X1 U1744 ( .A1(n2177), .A2(n2178), .ZN(n2149) );
NAND2_X1 U1745 ( .A1(RESTART), .A2(n1830), .ZN(n2178) );
NAND2_X1 U1746 ( .A1(n2179), .A2(n2030), .ZN(n2177) );
NAND2_X1 U1747 ( .A1(n2180), .A2(n2181), .ZN(n2147) );
NAND2_X1 U1748 ( .A1(n2182), .A2(n2183), .ZN(n2181) );
OR2_X1 U1749 ( .A1(n2184), .A2(n2185), .ZN(n2182) );
NAND2_X1 U1750 ( .A1(n2185), .A2(n2184), .ZN(n2180) );
NAND2_X1 U1751 ( .A1(n2186), .A2(n2187), .ZN(n2148) );
NAND2_X1 U1752 ( .A1(RESTART), .A2(n1771), .ZN(n2187) );
NAND2_X1 U1753 ( .A1(n1841), .A2(n2030), .ZN(n2186) );
NAND2_X1 U1754 ( .A1(DATA_OUT_REG_2__SCAN_IN), .A2(n1902), .ZN(n2154) );
NAND2_X1 U1755 ( .A1(n2006), .A2(RLAST_REG_2__SCAN_IN), .ZN(n2153) );
NAND2_X1 U1756 ( .A1(n1983), .A2(REG4_REG_2__SCAN_IN), .ZN(n2152) );
NAND4_X1 U1757 ( .A1(n2188), .A2(n2189), .A3(n2190), .A4(n2191), .ZN(U282));
NOR3_X1 U1758 ( .A1(n2192), .A2(n2193), .A3(n2194), .ZN(n2191) );
NOR2_X1 U1759 ( .A1(n1999), .A2(n2195), .ZN(n2194) );
XNOR2_X1 U1760 ( .A(n2173), .B(n2196), .ZN(n2195) );
NOR2_X1 U1761 ( .A1(KEYINPUT17), .A2(n2166), .ZN(n2196) );
NOR2_X1 U1762 ( .A1(n2197), .A2(n1992), .ZN(n2193) );
XOR2_X1 U1763 ( .A(n2198), .B(n2162), .Z(n2197) );
INV_X1 U1764 ( .A(n2166), .ZN(n2162) );
NAND2_X1 U1765 ( .A1(n2169), .A2(n2199), .ZN(n2166) );
NAND2_X1 U1766 ( .A1(n2200), .A2(n2201), .ZN(n2199) );
NAND2_X1 U1767 ( .A1(n2202), .A2(n2203), .ZN(n2201) );
NAND3_X1 U1768 ( .A1(n2204), .A2(n2203), .A3(n2202), .ZN(n2169) );
NAND2_X1 U1769 ( .A1(KEYINPUT36), .A2(n2163), .ZN(n2198) );
NOR2_X1 U1770 ( .A1(n2204), .A2(n2022), .ZN(n2192) );
INV_X1 U1771 ( .A(n2200), .ZN(n2204) );
NAND2_X1 U1772 ( .A1(n2205), .A2(n2206), .ZN(n2200) );
NAND2_X1 U1773 ( .A1(n2207), .A2(n2208), .ZN(n2206) );
NAND3_X1 U1774 ( .A1(n2209), .A2(n2210), .A3(n2211), .ZN(n2208) );
NAND2_X1 U1775 ( .A1(KEYINPUT8), .A2(n2212), .ZN(n2211) );
OR2_X1 U1776 ( .A1(n2212), .A2(KEYINPUT61), .ZN(n2210) );
NAND3_X1 U1777 ( .A1(n2184), .A2(n2213), .A3(KEYINPUT61), .ZN(n2209) );
INV_X1 U1778 ( .A(n2185), .ZN(n2213) );
INV_X1 U1779 ( .A(n2183), .ZN(n2207) );
NAND3_X1 U1780 ( .A1(n2212), .A2(n2214), .A3(n2183), .ZN(n2205) );
NAND2_X1 U1781 ( .A1(n2215), .A2(n2216), .ZN(n2183) );
NAND2_X1 U1782 ( .A1(n2217), .A2(n2218), .ZN(n2216) );
NAND2_X1 U1783 ( .A1(n2219), .A2(n2220), .ZN(n2217) );
XOR2_X1 U1784 ( .A(n2221), .B(KEYINPUT3), .Z(n2219) );
OR2_X1 U1785 ( .A1(n2220), .A2(n2222), .ZN(n2215) );
INV_X1 U1786 ( .A(KEYINPUT8), .ZN(n2214) );
XOR2_X1 U1787 ( .A(n2185), .B(n2184), .Z(n2212) );
NAND2_X1 U1788 ( .A1(n2223), .A2(n2224), .ZN(n2184) );
NAND2_X1 U1789 ( .A1(RESTART), .A2(n1870), .ZN(n2224) );
NAND2_X1 U1790 ( .A1(n1834), .A2(n2030), .ZN(n2223) );
NAND2_X1 U1791 ( .A1(n2225), .A2(n2226), .ZN(n2185) );
NAND2_X1 U1792 ( .A1(RESTART), .A2(n1839), .ZN(n2226) );
NAND2_X1 U1793 ( .A1(n2227), .A2(n2030), .ZN(n2225) );
XOR2_X1 U1794 ( .A(n2228), .B(KEYINPUT2), .Z(n2190) );
NAND2_X1 U1795 ( .A1(n2229), .A2(RLAST_REG_1__SCAN_IN), .ZN(n2228) );
XOR2_X1 U1796 ( .A(n1982), .B(KEYINPUT31), .Z(n2229) );
NAND2_X1 U1797 ( .A1(n1983), .A2(REG4_REG_1__SCAN_IN), .ZN(n2189) );
NAND2_X1 U1798 ( .A1(DATA_OUT_REG_1__SCAN_IN), .A2(n1902), .ZN(n2188) );
NAND4_X1 U1799 ( .A1(n2230), .A2(n2231), .A3(n2232), .A4(n2233), .ZN(U281));
NOR3_X1 U1800 ( .A1(n2234), .A2(n2235), .A3(n2236), .ZN(n2233) );
NOR2_X1 U1801 ( .A1(n2203), .A2(n2022), .ZN(n2236) );
NAND3_X1 U1802 ( .A1(n2237), .A2(n2238), .A3(n2239), .ZN(n2022) );
NAND2_X1 U1803 ( .A1(n2240), .A2(n2030), .ZN(n2238) );
NAND4_X1 U1804 ( .A1(ENABLE), .A2(n2241), .A3(n2242), .A4(n2243), .ZN(n2240));
INV_X1 U1805 ( .A(AVERAGE), .ZN(n2243) );
NAND2_X1 U1806 ( .A1(REG4_REG_7__SCAN_IN), .A2(DATA_IN_7_), .ZN(n2241) );
NAND2_X1 U1807 ( .A1(n2244), .A2(RESTART), .ZN(n2237) );
AND2_X1 U1808 ( .A1(RLAST_REG_0__SCAN_IN), .A2(n2006), .ZN(n2235) );
INV_X1 U1809 ( .A(n1982), .ZN(n2006) );
NAND3_X1 U1810 ( .A1(n1898), .A2(n2030), .A3(n2239), .ZN(n1982) );
INV_X1 U1811 ( .A(ENABLE), .ZN(n1898) );
AND2_X1 U1812 ( .A1(REG4_REG_0__SCAN_IN), .A2(n1983), .ZN(n2234) );
AND4_X1 U1813 ( .A1(ENABLE), .A2(AVERAGE), .A3(n2239), .A4(n2030), .ZN(n1983) );
NAND2_X1 U1814 ( .A1(DATA_OUT_REG_0__SCAN_IN), .A2(n1902), .ZN(n2232) );
NAND2_X1 U1815 ( .A1(n2163), .A2(n1993), .ZN(n2231) );
INV_X1 U1816 ( .A(n1992), .ZN(n1993) );
NAND3_X1 U1817 ( .A1(RESTART), .A2(n2239), .A3(n2244), .ZN(n1992) );
XOR2_X1 U1818 ( .A(n2245), .B(KEYINPUT46), .Z(n2244) );
NAND2_X1 U1819 ( .A1(n2246), .A2(n2247), .ZN(n2245) );
NAND2_X1 U1820 ( .A1(n2248), .A2(n2249), .ZN(n2247) );
NAND2_X1 U1821 ( .A1(RMIN_REG_7__SCAN_IN), .A2(RMAX_REG_7__SCAN_IN), .ZN(n2249) );
NAND2_X1 U1822 ( .A1(n2250), .A2(n2251), .ZN(n2248) );
NAND2_X1 U1823 ( .A1(RMIN_REG_6__SCAN_IN), .A2(RMAX_REG_6__SCAN_IN), .ZN(n2251) );
NAND3_X1 U1824 ( .A1(n2252), .A2(n2253), .A3(n2254), .ZN(n2250) );
NAND2_X1 U1825 ( .A1(n1876), .A2(n1843), .ZN(n2254) );
INV_X1 U1826 ( .A(RMIN_REG_5__SCAN_IN), .ZN(n1843) );
NAND3_X1 U1827 ( .A1(n2255), .A2(n2256), .A3(n2257), .ZN(n2253) );
NAND2_X1 U1828 ( .A1(RMIN_REG_4__SCAN_IN), .A2(RMAX_REG_4__SCAN_IN), .ZN(n2257) );
NAND3_X1 U1829 ( .A1(n2258), .A2(n2259), .A3(n2260), .ZN(n2256) );
NAND2_X1 U1830 ( .A1(n1767), .A2(n1822), .ZN(n2260) );
INV_X1 U1831 ( .A(RMIN_REG_4__SCAN_IN), .ZN(n1822) );
INV_X1 U1832 ( .A(RMAX_REG_4__SCAN_IN), .ZN(n1767) );
NAND3_X1 U1833 ( .A1(n2261), .A2(n2262), .A3(n2263), .ZN(n2259) );
NAND2_X1 U1834 ( .A1(RMIN_REG_3__SCAN_IN), .A2(RMAX_REG_3__SCAN_IN), .ZN(n2263) );
NAND3_X1 U1835 ( .A1(n2264), .A2(n2265), .A3(n2266), .ZN(n2262) );
NAND2_X1 U1836 ( .A1(n1874), .A2(n1837), .ZN(n2266) );
NAND2_X1 U1837 ( .A1(n2267), .A2(n2268), .ZN(n2265) );
NAND2_X1 U1838 ( .A1(RMIN_REG_1__SCAN_IN), .A2(RMAX_REG_1__SCAN_IN), .ZN(n2268) );
NAND2_X1 U1839 ( .A1(RMIN_REG_0__SCAN_IN), .A2(RMAX_REG_0__SCAN_IN), .ZN(n2267) );
NAND2_X1 U1840 ( .A1(n2269), .A2(n1870), .ZN(n2264) );
INV_X1 U1841 ( .A(RMAX_REG_2__SCAN_IN), .ZN(n1870) );
XOR2_X1 U1842 ( .A(RMIN_REG_2__SCAN_IN), .B(KEYINPUT62), .Z(n2269) );
NAND2_X1 U1843 ( .A1(n2270), .A2(RMAX_REG_2__SCAN_IN), .ZN(n2261) );
XOR2_X1 U1844 ( .A(n1839), .B(KEYINPUT6), .Z(n2270) );
INV_X1 U1845 ( .A(RMIN_REG_2__SCAN_IN), .ZN(n1839) );
NAND2_X1 U1846 ( .A1(n1771), .A2(n1830), .ZN(n2258) );
INV_X1 U1847 ( .A(RMIN_REG_3__SCAN_IN), .ZN(n1830) );
INV_X1 U1848 ( .A(RMAX_REG_3__SCAN_IN), .ZN(n1771) );
NAND2_X1 U1849 ( .A1(n2271), .A2(RMIN_REG_5__SCAN_IN), .ZN(n2255) );
XOR2_X1 U1850 ( .A(n1876), .B(KEYINPUT40), .Z(n2271) );
INV_X1 U1851 ( .A(RMAX_REG_5__SCAN_IN), .ZN(n1876) );
NAND2_X1 U1852 ( .A1(n2272), .A2(n1846), .ZN(n2252) );
INV_X1 U1853 ( .A(RMIN_REG_6__SCAN_IN), .ZN(n1846) );
XOR2_X1 U1854 ( .A(RMAX_REG_6__SCAN_IN), .B(KEYINPUT28), .Z(n2272) );
NAND2_X1 U1855 ( .A1(n1853), .A2(n1847), .ZN(n2246) );
INV_X1 U1856 ( .A(RMIN_REG_7__SCAN_IN), .ZN(n1847) );
INV_X1 U1857 ( .A(RMAX_REG_7__SCAN_IN), .ZN(n1853) );
XNOR2_X1 U1858 ( .A(n2273), .B(n2203), .ZN(n2163) );
NAND2_X1 U1859 ( .A1(n1976), .A2(n2173), .ZN(n2230) );
NAND2_X1 U1860 ( .A1(n2274), .A2(n2275), .ZN(n2173) );
NAND2_X1 U1861 ( .A1(n2203), .A2(n2273), .ZN(n2275) );
INV_X1 U1862 ( .A(n2276), .ZN(n2203) );
XOR2_X1 U1863 ( .A(n2277), .B(KEYINPUT35), .Z(n2274) );
NAND2_X1 U1864 ( .A1(n2202), .A2(n2276), .ZN(n2277) );
XOR2_X1 U1865 ( .A(n2278), .B(n2222), .Z(n2276) );
INV_X1 U1866 ( .A(n2221), .ZN(n2222) );
NAND2_X1 U1867 ( .A1(n2279), .A2(n2280), .ZN(n2221) );
NAND2_X1 U1868 ( .A1(n2281), .A2(n2282), .ZN(n2278) );
NAND2_X1 U1869 ( .A1(n2218), .A2(n2220), .ZN(n2282) );
NAND2_X1 U1870 ( .A1(n2283), .A2(n2284), .ZN(n2281) );
NAND2_X1 U1871 ( .A1(KEYINPUT3), .A2(n2220), .ZN(n2284) );
NAND3_X1 U1872 ( .A1(n2285), .A2(n2286), .A3(n2287), .ZN(n2220) );
NAND2_X1 U1873 ( .A1(KEYINPUT0), .A2(n1838), .ZN(n2287) );
INV_X1 U1874 ( .A(DATA_IN_1_), .ZN(n1838) );
NAND3_X1 U1875 ( .A1(DATA_IN_1_), .A2(n2288), .A3(n2030), .ZN(n2286) );
NAND2_X1 U1876 ( .A1(RESTART), .A2(n2289), .ZN(n2285) );
NAND2_X1 U1877 ( .A1(n1874), .A2(n2288), .ZN(n2289) );
INV_X1 U1878 ( .A(KEYINPUT0), .ZN(n2288) );
INV_X1 U1879 ( .A(RMAX_REG_1__SCAN_IN), .ZN(n1874) );
INV_X1 U1880 ( .A(n2218), .ZN(n2283) );
NAND2_X1 U1881 ( .A1(n2290), .A2(n2291), .ZN(n2218) );
NAND2_X1 U1882 ( .A1(n2292), .A2(n2030), .ZN(n2291) );
NAND2_X1 U1883 ( .A1(REG4_REG_1__SCAN_IN), .A2(n2293), .ZN(n2292) );
NAND2_X1 U1884 ( .A1(n2294), .A2(n1837), .ZN(n2290) );
INV_X1 U1885 ( .A(RMIN_REG_1__SCAN_IN), .ZN(n1837) );
NAND2_X1 U1886 ( .A1(REG4_REG_1__SCAN_IN), .A2(n2295), .ZN(n2294) );
NAND2_X1 U1887 ( .A1(RESTART), .A2(n2293), .ZN(n2295) );
INV_X1 U1888 ( .A(KEYINPUT30), .ZN(n2293) );
INV_X1 U1889 ( .A(n2273), .ZN(n2202) );
NAND2_X1 U1890 ( .A1(n2296), .A2(n2297), .ZN(n2273) );
NAND2_X1 U1891 ( .A1(n2298), .A2(n2279), .ZN(n2297) );
XOR2_X1 U1892 ( .A(KEYINPUT52), .B(n2299), .Z(n2296) );
NOR2_X1 U1893 ( .A1(n2298), .A2(n2279), .ZN(n2299) );
NAND2_X1 U1894 ( .A1(n2300), .A2(n2301), .ZN(n2279) );
NAND2_X1 U1895 ( .A1(REG4_REG_0__SCAN_IN), .A2(n2030), .ZN(n2301) );
NAND2_X1 U1896 ( .A1(RESTART), .A2(RMIN_REG_0__SCAN_IN), .ZN(n2300) );
INV_X1 U1897 ( .A(n2280), .ZN(n2298) );
NAND3_X1 U1898 ( .A1(n2302), .A2(n2303), .A3(n2304), .ZN(n2280) );
OR2_X1 U1899 ( .A1(DATA_IN_0_), .A2(KEYINPUT15), .ZN(n2304) );
NAND3_X1 U1900 ( .A1(KEYINPUT15), .A2(DATA_IN_0_), .A3(n2030), .ZN(n2303) );
INV_X1 U1901 ( .A(RESTART), .ZN(n2030) );
NAND2_X1 U1902 ( .A1(RESTART), .A2(n2305), .ZN(n2302) );
NAND2_X1 U1903 ( .A1(KEYINPUT15), .A2(n1872), .ZN(n2305) );
INV_X1 U1904 ( .A(RMAX_REG_0__SCAN_IN), .ZN(n1872) );
INV_X1 U1905 ( .A(n1999), .ZN(n1976) );
NAND4_X1 U1906 ( .A1(ENABLE), .A2(n2239), .A3(n2306), .A4(n2307), .ZN(n1999));
XOR2_X1 U1907 ( .A(KEYINPUT32), .B(AVERAGE), .Z(n2307) );
NOR2_X1 U1908 ( .A1(RESTART), .A2(n2308), .ZN(n2306) );
NOR2_X1 U1909 ( .A1(n2309), .A2(n2310), .ZN(n2308) );
AND2_X1 U1910 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2310) );
INV_X1 U1911 ( .A(n2242), .ZN(n2309) );
NAND3_X1 U1912 ( .A1(n2311), .A2(n2312), .A3(n2313), .ZN(n2242) );
XOR2_X1 U1913 ( .A(KEYINPUT38), .B(n2314), .Z(n2313) );
NOR2_X1 U1914 ( .A1(DATA_IN_7_), .A2(REG4_REG_7__SCAN_IN), .ZN(n2314) );
NAND3_X1 U1915 ( .A1(n2315), .A2(n2316), .A3(n2317), .ZN(n2312) );
NAND2_X1 U1916 ( .A1(n1845), .A2(n2039), .ZN(n2317) );
INV_X1 U1917 ( .A(REG4_REG_6__SCAN_IN), .ZN(n2039) );
INV_X1 U1918 ( .A(DATA_IN_6_), .ZN(n1845) );
NAND3_X1 U1919 ( .A1(n2318), .A2(n2319), .A3(n2320), .ZN(n2316) );
NAND2_X1 U1920 ( .A1(REG4_REG_5__SCAN_IN), .A2(DATA_IN_5_), .ZN(n2320) );
NAND3_X1 U1921 ( .A1(n2321), .A2(n2322), .A3(n2323), .ZN(n2319) );
NAND2_X1 U1922 ( .A1(n1826), .A2(n1963), .ZN(n2323) );
INV_X1 U1923 ( .A(REG4_REG_4__SCAN_IN), .ZN(n1963) );
INV_X1 U1924 ( .A(DATA_IN_4_), .ZN(n1826) );
NAND3_X1 U1925 ( .A1(n2324), .A2(n2325), .A3(n2326), .ZN(n2322) );
NAND2_X1 U1926 ( .A1(REG4_REG_2__SCAN_IN), .A2(DATA_IN_2_), .ZN(n2326) );
NAND3_X1 U1927 ( .A1(n2327), .A2(n2328), .A3(n2329), .ZN(n2325) );
NAND2_X1 U1928 ( .A1(n1834), .A2(n2227), .ZN(n2329) );
INV_X1 U1929 ( .A(REG4_REG_2__SCAN_IN), .ZN(n2227) );
INV_X1 U1930 ( .A(DATA_IN_2_), .ZN(n1834) );
NAND2_X1 U1931 ( .A1(n2330), .A2(n2331), .ZN(n2328) );
NAND2_X1 U1932 ( .A1(REG4_REG_1__SCAN_IN), .A2(DATA_IN_1_), .ZN(n2331) );
NAND2_X1 U1933 ( .A1(REG4_REG_0__SCAN_IN), .A2(DATA_IN_0_), .ZN(n2330) );
OR2_X1 U1934 ( .A1(DATA_IN_1_), .A2(REG4_REG_1__SCAN_IN), .ZN(n2327) );
NAND2_X1 U1935 ( .A1(n2332), .A2(REG4_REG_3__SCAN_IN), .ZN(n2324) );
XOR2_X1 U1936 ( .A(n1841), .B(KEYINPUT4), .Z(n2332) );
NAND2_X1 U1937 ( .A1(n1841), .A2(n2179), .ZN(n2321) );
INV_X1 U1938 ( .A(REG4_REG_3__SCAN_IN), .ZN(n2179) );
INV_X1 U1939 ( .A(DATA_IN_3_), .ZN(n1841) );
NAND2_X1 U1940 ( .A1(REG4_REG_4__SCAN_IN), .A2(DATA_IN_4_), .ZN(n2318) );
NAND2_X1 U1941 ( .A1(n1818), .A2(n2094), .ZN(n2315) );
INV_X1 U1942 ( .A(REG4_REG_5__SCAN_IN), .ZN(n2094) );
INV_X1 U1943 ( .A(DATA_IN_5_), .ZN(n1818) );
NAND2_X1 U1944 ( .A1(REG4_REG_6__SCAN_IN), .A2(DATA_IN_6_), .ZN(n2311) );
AND2_X1 U1945 ( .A1(STATO_REG_1__SCAN_IN), .A2(n2333), .ZN(n2239) );
XOR2_X1 U1946 ( .A(KEYINPUT48), .B(n1902), .Z(n2333) );
NAND2_X1 U1947 ( .A1(n2334), .A2(n1910), .ZN(U280) );
NAND2_X1 U1948 ( .A1(STATO_REG_1__SCAN_IN), .A2(n1782), .ZN(n1910) );
XOR2_X1 U1949 ( .A(n2335), .B(KEYINPUT23), .Z(n2334) );
OR2_X1 U1950 ( .A1(n1782), .A2(STATO_REG_1__SCAN_IN), .ZN(n2335) );
INV_X1 U1951 ( .A(STATO_REG_0__SCAN_IN), .ZN(n1782) );
endmodule


