//Key = 1111111000101111011000101010011001011000101111110100101001000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293;

XNOR2_X1 U716 ( .A(G107), .B(n982), .ZN(G9) );
NOR2_X1 U717 ( .A1(n983), .A2(n984), .ZN(G75) );
NOR3_X1 U718 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n984) );
NOR3_X1 U719 ( .A1(n988), .A2(n989), .A3(n990), .ZN(n986) );
INV_X1 U720 ( .A(n991), .ZN(n990) );
NOR2_X1 U721 ( .A1(n992), .A2(n993), .ZN(n989) );
NOR2_X1 U722 ( .A1(n994), .A2(n995), .ZN(n993) );
INV_X1 U723 ( .A(n996), .ZN(n995) );
NOR2_X1 U724 ( .A1(n997), .A2(n998), .ZN(n994) );
NOR2_X1 U725 ( .A1(n999), .A2(n1000), .ZN(n998) );
NOR2_X1 U726 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NOR2_X1 U727 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U728 ( .A1(n1005), .A2(n1006), .ZN(n997) );
NOR2_X1 U729 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR3_X1 U730 ( .A1(n1000), .A2(n1009), .A3(n1006), .ZN(n992) );
NOR2_X1 U731 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR2_X1 U732 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
NAND3_X1 U733 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n985) );
NAND3_X1 U734 ( .A1(n1017), .A2(n1018), .A3(n996), .ZN(n1016) );
NAND2_X1 U735 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
INV_X1 U736 ( .A(KEYINPUT59), .ZN(n1020) );
NAND2_X1 U737 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
OR2_X1 U738 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND3_X1 U739 ( .A1(n1021), .A2(n1023), .A3(KEYINPUT59), .ZN(n1017) );
NOR3_X1 U740 ( .A1(n1000), .A2(n1006), .A3(n988), .ZN(n1021) );
NOR3_X1 U741 ( .A1(n1025), .A2(G953), .A3(G952), .ZN(n983) );
INV_X1 U742 ( .A(n1014), .ZN(n1025) );
NAND4_X1 U743 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1014) );
NOR3_X1 U744 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NOR2_X1 U745 ( .A1(KEYINPUT1), .A2(n1033), .ZN(n1032) );
XOR2_X1 U746 ( .A(n1034), .B(G478), .Z(n1031) );
NAND2_X1 U747 ( .A1(KEYINPUT6), .A2(n1035), .ZN(n1034) );
XOR2_X1 U748 ( .A(KEYINPUT14), .B(n1036), .Z(n1035) );
NAND3_X1 U749 ( .A1(n1013), .A2(n1037), .A3(n1038), .ZN(n1030) );
NOR3_X1 U750 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1028) );
NOR2_X1 U751 ( .A1(G472), .A2(n1042), .ZN(n1041) );
NOR2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
XNOR2_X1 U753 ( .A(n1045), .B(KEYINPUT62), .ZN(n1043) );
NOR3_X1 U754 ( .A1(n1046), .A2(n1045), .A3(n1044), .ZN(n1040) );
INV_X1 U755 ( .A(KEYINPUT1), .ZN(n1044) );
XOR2_X1 U756 ( .A(n1047), .B(n1048), .Z(n1039) );
XNOR2_X1 U757 ( .A(n1049), .B(KEYINPUT48), .ZN(n1048) );
XOR2_X1 U758 ( .A(n1050), .B(n1051), .Z(G72) );
XOR2_X1 U759 ( .A(n1052), .B(n1053), .Z(n1051) );
NOR2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
XNOR2_X1 U761 ( .A(KEYINPUT28), .B(n1015), .ZN(n1055) );
NOR2_X1 U762 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
XNOR2_X1 U763 ( .A(KEYINPUT46), .B(n1015), .ZN(n1057) );
AND2_X1 U764 ( .A1(G227), .A2(G900), .ZN(n1056) );
NOR2_X1 U765 ( .A1(n1058), .A2(n1059), .ZN(n1050) );
XOR2_X1 U766 ( .A(n1060), .B(n1061), .Z(n1059) );
XOR2_X1 U767 ( .A(n1062), .B(n1063), .Z(n1061) );
XOR2_X1 U768 ( .A(n1064), .B(KEYINPUT33), .Z(n1063) );
NAND2_X1 U769 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U770 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U771 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NAND2_X1 U772 ( .A1(KEYINPUT52), .A2(G140), .ZN(n1070) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1072), .ZN(n1065) );
NAND2_X1 U774 ( .A1(KEYINPUT52), .A2(n1073), .ZN(n1071) );
NAND2_X1 U775 ( .A1(n1074), .A2(n1069), .ZN(n1073) );
INV_X1 U776 ( .A(KEYINPUT21), .ZN(n1069) );
NAND2_X1 U777 ( .A1(KEYINPUT40), .A2(G131), .ZN(n1062) );
XNOR2_X1 U778 ( .A(n1075), .B(n1076), .ZN(n1060) );
XOR2_X1 U779 ( .A(n1077), .B(n1078), .Z(G69) );
NOR3_X1 U780 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NOR2_X1 U781 ( .A1(G953), .A2(n1082), .ZN(n1081) );
NOR2_X1 U782 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
XOR2_X1 U783 ( .A(n982), .B(KEYINPUT26), .Z(n1083) );
NOR2_X1 U784 ( .A1(G224), .A2(n1015), .ZN(n1080) );
NAND2_X1 U785 ( .A1(n1085), .A2(n1086), .ZN(n1077) );
INV_X1 U786 ( .A(n1079), .ZN(n1086) );
NOR2_X1 U787 ( .A1(n1087), .A2(n1088), .ZN(G66) );
XNOR2_X1 U788 ( .A(n1089), .B(n1090), .ZN(n1088) );
XOR2_X1 U789 ( .A(KEYINPUT37), .B(n1091), .Z(n1090) );
NOR2_X1 U790 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR2_X1 U791 ( .A1(n1094), .A2(n1095), .ZN(n1087) );
XNOR2_X1 U792 ( .A(KEYINPUT3), .B(n1015), .ZN(n1095) );
XNOR2_X1 U793 ( .A(KEYINPUT47), .B(G952), .ZN(n1094) );
NOR2_X1 U794 ( .A1(n1096), .A2(n1097), .ZN(G63) );
NOR3_X1 U795 ( .A1(n1036), .A2(n1098), .A3(n1099), .ZN(n1097) );
AND3_X1 U796 ( .A1(n1100), .A2(G478), .A3(n1101), .ZN(n1099) );
NOR2_X1 U797 ( .A1(n1102), .A2(n1100), .ZN(n1098) );
AND2_X1 U798 ( .A1(n987), .A2(G478), .ZN(n1102) );
NOR2_X1 U799 ( .A1(n1096), .A2(n1103), .ZN(G60) );
XOR2_X1 U800 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U801 ( .A1(KEYINPUT27), .A2(n1106), .ZN(n1105) );
NAND2_X1 U802 ( .A1(n1101), .A2(G475), .ZN(n1104) );
XOR2_X1 U803 ( .A(n1107), .B(n1108), .Z(G6) );
NOR2_X1 U804 ( .A1(KEYINPUT39), .A2(G104), .ZN(n1108) );
NAND3_X1 U805 ( .A1(n1109), .A2(n991), .A3(n1008), .ZN(n1107) );
NOR2_X1 U806 ( .A1(n1096), .A2(n1110), .ZN(G57) );
XOR2_X1 U807 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U808 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR3_X1 U809 ( .A1(n1093), .A2(KEYINPUT8), .A3(n1046), .ZN(n1113) );
INV_X1 U810 ( .A(G472), .ZN(n1046) );
XOR2_X1 U811 ( .A(n1115), .B(n1116), .Z(n1111) );
XOR2_X1 U812 ( .A(n1117), .B(G101), .Z(n1116) );
NAND2_X1 U813 ( .A1(KEYINPUT17), .A2(n1118), .ZN(n1115) );
NOR2_X1 U814 ( .A1(n1096), .A2(n1119), .ZN(G54) );
XOR2_X1 U815 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U816 ( .A1(KEYINPUT53), .A2(n1122), .ZN(n1121) );
XOR2_X1 U817 ( .A(n1123), .B(n1124), .Z(n1122) );
XNOR2_X1 U818 ( .A(n1125), .B(n1126), .ZN(n1124) );
NAND2_X1 U819 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NAND2_X1 U820 ( .A1(n1129), .A2(n1072), .ZN(n1128) );
NAND2_X1 U821 ( .A1(n1130), .A2(G140), .ZN(n1127) );
XOR2_X1 U822 ( .A(KEYINPUT54), .B(n1129), .Z(n1130) );
XOR2_X1 U823 ( .A(G110), .B(n1131), .Z(n1129) );
XNOR2_X1 U824 ( .A(n1076), .B(n1132), .ZN(n1123) );
XNOR2_X1 U825 ( .A(n1133), .B(KEYINPUT22), .ZN(n1132) );
NAND2_X1 U826 ( .A1(KEYINPUT49), .A2(n1134), .ZN(n1133) );
NAND2_X1 U827 ( .A1(n1101), .A2(G469), .ZN(n1120) );
NOR2_X1 U828 ( .A1(n1096), .A2(n1135), .ZN(G51) );
XOR2_X1 U829 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U830 ( .A(n1138), .B(n1139), .Z(n1137) );
AND2_X1 U831 ( .A1(G210), .A2(n1101), .ZN(n1138) );
INV_X1 U832 ( .A(n1093), .ZN(n1101) );
NAND2_X1 U833 ( .A1(G902), .A2(n987), .ZN(n1093) );
NAND3_X1 U834 ( .A1(n1054), .A2(n982), .A3(n1140), .ZN(n987) );
INV_X1 U835 ( .A(n1084), .ZN(n1140) );
NAND4_X1 U836 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1084) );
NOR4_X1 U837 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1144) );
NAND3_X1 U838 ( .A1(n1008), .A2(n1109), .A3(n1149), .ZN(n1143) );
XNOR2_X1 U839 ( .A(KEYINPUT18), .B(n991), .ZN(n1149) );
NAND3_X1 U840 ( .A1(n1007), .A2(n991), .A3(n1109), .ZN(n982) );
AND2_X1 U841 ( .A1(n1150), .A2(n1151), .ZN(n1054) );
NOR4_X1 U842 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1151) );
NOR4_X1 U843 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1150) );
NOR2_X1 U844 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XNOR2_X1 U845 ( .A(n1002), .B(KEYINPUT19), .ZN(n1160) );
INV_X1 U846 ( .A(n1162), .ZN(n1158) );
NOR2_X1 U847 ( .A1(n1163), .A2(n1164), .ZN(n1136) );
NOR3_X1 U848 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1164) );
INV_X1 U849 ( .A(KEYINPUT55), .ZN(n1165) );
NOR2_X1 U850 ( .A1(KEYINPUT55), .A2(n1168), .ZN(n1163) );
AND2_X1 U851 ( .A1(G953), .A2(n1169), .ZN(n1096) );
XOR2_X1 U852 ( .A(KEYINPUT47), .B(G952), .Z(n1169) );
XNOR2_X1 U853 ( .A(G146), .B(n1170), .ZN(G48) );
OR2_X1 U854 ( .A1(n1161), .A2(n1171), .ZN(n1170) );
NAND3_X1 U855 ( .A1(n1008), .A2(n1172), .A3(n1173), .ZN(n1161) );
NAND2_X1 U856 ( .A1(n1174), .A2(n1175), .ZN(G45) );
OR2_X1 U857 ( .A1(n1162), .A2(G143), .ZN(n1175) );
XOR2_X1 U858 ( .A(n1176), .B(KEYINPUT31), .Z(n1174) );
NAND2_X1 U859 ( .A1(G143), .A2(n1162), .ZN(n1176) );
NAND3_X1 U860 ( .A1(n1173), .A2(n1024), .A3(n1177), .ZN(n1162) );
NOR3_X1 U861 ( .A1(n1171), .A2(n1178), .A3(n1026), .ZN(n1177) );
XNOR2_X1 U862 ( .A(n1072), .B(n1157), .ZN(G42) );
AND3_X1 U863 ( .A1(n1008), .A2(n1023), .A3(n1179), .ZN(n1157) );
XOR2_X1 U864 ( .A(G137), .B(n1156), .Z(G39) );
AND3_X1 U865 ( .A1(n1180), .A2(n1172), .A3(n1179), .ZN(n1156) );
XNOR2_X1 U866 ( .A(n1181), .B(n1155), .ZN(G36) );
AND3_X1 U867 ( .A1(n1007), .A2(n1024), .A3(n1179), .ZN(n1155) );
XOR2_X1 U868 ( .A(G131), .B(n1154), .Z(G33) );
AND3_X1 U869 ( .A1(n1008), .A2(n1024), .A3(n1179), .ZN(n1154) );
AND3_X1 U870 ( .A1(n1002), .A2(n1182), .A3(n996), .ZN(n1179) );
NOR2_X1 U871 ( .A1(n1183), .A2(n1012), .ZN(n996) );
XOR2_X1 U872 ( .A(n1184), .B(KEYINPUT20), .Z(n1012) );
XNOR2_X1 U873 ( .A(n1013), .B(KEYINPUT34), .ZN(n1183) );
XNOR2_X1 U874 ( .A(G128), .B(n1185), .ZN(G30) );
NOR2_X1 U875 ( .A1(n1153), .A2(KEYINPUT25), .ZN(n1185) );
AND4_X1 U876 ( .A1(n1173), .A2(n1172), .A3(n1007), .A4(n1002), .ZN(n1153) );
XNOR2_X1 U877 ( .A(G101), .B(n1141), .ZN(G3) );
NAND3_X1 U878 ( .A1(n1109), .A2(n1024), .A3(n1180), .ZN(n1141) );
XOR2_X1 U879 ( .A(G125), .B(n1152), .Z(G27) );
AND4_X1 U880 ( .A1(n1173), .A2(n1008), .A3(n1027), .A4(n1023), .ZN(n1152) );
AND2_X1 U881 ( .A1(n1011), .A2(n1182), .ZN(n1173) );
NAND2_X1 U882 ( .A1(n988), .A2(n1186), .ZN(n1182) );
NAND3_X1 U883 ( .A1(G902), .A2(n1187), .A3(n1058), .ZN(n1186) );
NOR2_X1 U884 ( .A1(n1015), .A2(G900), .ZN(n1058) );
XNOR2_X1 U885 ( .A(G122), .B(n1142), .ZN(G24) );
NAND4_X1 U886 ( .A1(n1188), .A2(n991), .A3(n1189), .A4(n1190), .ZN(n1142) );
NAND2_X1 U887 ( .A1(n1191), .A2(n1192), .ZN(n991) );
NAND2_X1 U888 ( .A1(n1024), .A2(n1193), .ZN(n1192) );
NAND3_X1 U889 ( .A1(n1194), .A2(n1195), .A3(KEYINPUT43), .ZN(n1191) );
XOR2_X1 U890 ( .A(n1148), .B(n1196), .Z(G21) );
NOR2_X1 U891 ( .A1(KEYINPUT58), .A2(n1197), .ZN(n1196) );
AND3_X1 U892 ( .A1(n1180), .A2(n1172), .A3(n1188), .ZN(n1148) );
XOR2_X1 U893 ( .A(G116), .B(n1147), .Z(G18) );
AND3_X1 U894 ( .A1(n1007), .A2(n1024), .A3(n1188), .ZN(n1147) );
NOR2_X1 U895 ( .A1(n1189), .A2(n1178), .ZN(n1007) );
XNOR2_X1 U896 ( .A(n1198), .B(n1146), .ZN(G15) );
AND3_X1 U897 ( .A1(n1008), .A2(n1024), .A3(n1188), .ZN(n1146) );
AND3_X1 U898 ( .A1(n1011), .A2(n1199), .A3(n1027), .ZN(n1188) );
INV_X1 U899 ( .A(n1006), .ZN(n1027) );
NAND2_X1 U900 ( .A1(n1200), .A2(n1004), .ZN(n1006) );
INV_X1 U901 ( .A(n1003), .ZN(n1200) );
NOR2_X1 U902 ( .A1(n1195), .A2(n1201), .ZN(n1024) );
AND2_X1 U903 ( .A1(n1202), .A2(n1189), .ZN(n1008) );
XOR2_X1 U904 ( .A(G110), .B(n1145), .Z(G12) );
AND3_X1 U905 ( .A1(n1109), .A2(n1023), .A3(n1180), .ZN(n1145) );
INV_X1 U906 ( .A(n1000), .ZN(n1180) );
NAND2_X1 U907 ( .A1(n1202), .A2(n1026), .ZN(n1000) );
INV_X1 U908 ( .A(n1189), .ZN(n1026) );
XNOR2_X1 U909 ( .A(n1203), .B(G475), .ZN(n1189) );
OR2_X1 U910 ( .A1(n1106), .A2(G902), .ZN(n1203) );
XNOR2_X1 U911 ( .A(n1204), .B(n1205), .ZN(n1106) );
XNOR2_X1 U912 ( .A(n1198), .B(n1206), .ZN(n1205) );
XOR2_X1 U913 ( .A(KEYINPUT15), .B(G122), .Z(n1206) );
XOR2_X1 U914 ( .A(n1207), .B(G104), .Z(n1204) );
NAND2_X1 U915 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U916 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U917 ( .A(KEYINPUT5), .B(n1212), .Z(n1208) );
NOR2_X1 U918 ( .A1(n1210), .A2(n1211), .ZN(n1212) );
XNOR2_X1 U919 ( .A(n1213), .B(n1214), .ZN(n1211) );
XOR2_X1 U920 ( .A(n1215), .B(KEYINPUT23), .Z(n1213) );
NAND2_X1 U921 ( .A1(n1216), .A2(n1072), .ZN(n1215) );
XNOR2_X1 U922 ( .A(KEYINPUT30), .B(KEYINPUT10), .ZN(n1216) );
XOR2_X1 U923 ( .A(n1217), .B(n1218), .Z(n1210) );
XOR2_X1 U924 ( .A(G143), .B(G131), .Z(n1218) );
NAND2_X1 U925 ( .A1(n1219), .A2(G214), .ZN(n1217) );
XNOR2_X1 U926 ( .A(n1190), .B(KEYINPUT41), .ZN(n1202) );
INV_X1 U927 ( .A(n1178), .ZN(n1190) );
XNOR2_X1 U928 ( .A(n1036), .B(G478), .ZN(n1178) );
NOR2_X1 U929 ( .A1(n1100), .A2(G902), .ZN(n1036) );
XOR2_X1 U930 ( .A(n1220), .B(n1221), .Z(n1100) );
XNOR2_X1 U931 ( .A(n1222), .B(n1223), .ZN(n1221) );
NAND2_X1 U932 ( .A1(G217), .A2(n1224), .ZN(n1222) );
XOR2_X1 U933 ( .A(n1225), .B(n1226), .Z(n1220) );
XNOR2_X1 U934 ( .A(n1181), .B(G107), .ZN(n1226) );
INV_X1 U935 ( .A(G134), .ZN(n1181) );
NAND2_X1 U936 ( .A1(KEYINPUT36), .A2(n1227), .ZN(n1225) );
NAND2_X1 U937 ( .A1(n1228), .A2(n1229), .ZN(n1023) );
NAND2_X1 U938 ( .A1(n1172), .A2(n1193), .ZN(n1229) );
INV_X1 U939 ( .A(KEYINPUT43), .ZN(n1193) );
NOR2_X1 U940 ( .A1(n1195), .A2(n1194), .ZN(n1172) );
INV_X1 U941 ( .A(n1201), .ZN(n1194) );
NAND3_X1 U942 ( .A1(n1195), .A2(n1201), .A3(KEYINPUT43), .ZN(n1228) );
NAND2_X1 U943 ( .A1(n1230), .A2(n1231), .ZN(n1201) );
NAND2_X1 U944 ( .A1(n1049), .A2(n1047), .ZN(n1231) );
XOR2_X1 U945 ( .A(KEYINPUT44), .B(n1232), .Z(n1230) );
NOR2_X1 U946 ( .A1(n1049), .A2(n1047), .ZN(n1232) );
NAND2_X1 U947 ( .A1(n1089), .A2(n1233), .ZN(n1047) );
XNOR2_X1 U948 ( .A(n1234), .B(n1235), .ZN(n1089) );
XNOR2_X1 U949 ( .A(n1214), .B(n1236), .ZN(n1235) );
XOR2_X1 U950 ( .A(n1237), .B(n1238), .Z(n1236) );
NOR2_X1 U951 ( .A1(KEYINPUT32), .A2(n1239), .ZN(n1238) );
XOR2_X1 U952 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U953 ( .A(G128), .B(G110), .ZN(n1240) );
NAND2_X1 U954 ( .A1(n1224), .A2(G221), .ZN(n1237) );
AND2_X1 U955 ( .A1(G234), .A2(n1015), .ZN(n1224) );
XNOR2_X1 U956 ( .A(G146), .B(n1074), .ZN(n1214) );
INV_X1 U957 ( .A(n1067), .ZN(n1074) );
XNOR2_X1 U958 ( .A(G137), .B(n1242), .ZN(n1234) );
XNOR2_X1 U959 ( .A(KEYINPUT9), .B(n1072), .ZN(n1242) );
INV_X1 U960 ( .A(G140), .ZN(n1072) );
INV_X1 U961 ( .A(n1092), .ZN(n1049) );
NAND2_X1 U962 ( .A1(G217), .A2(n1243), .ZN(n1092) );
XOR2_X1 U963 ( .A(n1045), .B(n1244), .Z(n1195) );
NOR2_X1 U964 ( .A1(G472), .A2(KEYINPUT7), .ZN(n1244) );
INV_X1 U965 ( .A(n1033), .ZN(n1045) );
NAND2_X1 U966 ( .A1(n1245), .A2(n1233), .ZN(n1033) );
XOR2_X1 U967 ( .A(n1246), .B(n1247), .Z(n1245) );
XNOR2_X1 U968 ( .A(n1117), .B(n1248), .ZN(n1247) );
NOR2_X1 U969 ( .A1(G101), .A2(KEYINPUT11), .ZN(n1248) );
NAND2_X1 U970 ( .A1(n1219), .A2(G210), .ZN(n1117) );
NOR2_X1 U971 ( .A1(G953), .A2(G237), .ZN(n1219) );
XOR2_X1 U972 ( .A(n1114), .B(n1118), .Z(n1246) );
XOR2_X1 U973 ( .A(n1249), .B(n1250), .Z(n1118) );
XOR2_X1 U974 ( .A(KEYINPUT29), .B(G116), .Z(n1250) );
XNOR2_X1 U975 ( .A(G113), .B(n1241), .ZN(n1249) );
XOR2_X1 U976 ( .A(n1251), .B(n1166), .Z(n1114) );
XNOR2_X1 U977 ( .A(n1134), .B(KEYINPUT0), .ZN(n1251) );
AND3_X1 U978 ( .A1(n1011), .A2(n1199), .A3(n1002), .ZN(n1109) );
INV_X1 U979 ( .A(n1171), .ZN(n1002) );
NAND2_X1 U980 ( .A1(n1003), .A2(n1004), .ZN(n1171) );
NAND2_X1 U981 ( .A1(G221), .A2(n1243), .ZN(n1004) );
NAND2_X1 U982 ( .A1(G234), .A2(n1233), .ZN(n1243) );
XNOR2_X1 U983 ( .A(n1252), .B(G469), .ZN(n1003) );
NAND2_X1 U984 ( .A1(n1253), .A2(n1233), .ZN(n1252) );
XOR2_X1 U985 ( .A(n1254), .B(n1255), .Z(n1253) );
XNOR2_X1 U986 ( .A(n1256), .B(n1131), .ZN(n1255) );
AND2_X1 U987 ( .A1(G227), .A2(n1015), .ZN(n1131) );
NAND3_X1 U988 ( .A1(n1257), .A2(n1258), .A3(n1259), .ZN(n1256) );
NAND2_X1 U989 ( .A1(n1166), .A2(n1260), .ZN(n1259) );
OR3_X1 U990 ( .A1(n1260), .A2(n1261), .A3(n1125), .ZN(n1258) );
INV_X1 U991 ( .A(KEYINPUT24), .ZN(n1260) );
NAND2_X1 U992 ( .A1(n1125), .A2(n1261), .ZN(n1257) );
NAND2_X1 U993 ( .A1(KEYINPUT2), .A2(n1076), .ZN(n1261) );
XNOR2_X1 U994 ( .A(n1262), .B(n1263), .ZN(n1254) );
NAND2_X1 U995 ( .A1(KEYINPUT61), .A2(n1134), .ZN(n1263) );
AND3_X1 U996 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1134) );
OR2_X1 U997 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NAND2_X1 U998 ( .A1(KEYINPUT38), .A2(n1269), .ZN(n1265) );
NAND2_X1 U999 ( .A1(n1270), .A2(n1267), .ZN(n1269) );
XNOR2_X1 U1000 ( .A(KEYINPUT56), .B(n1075), .ZN(n1270) );
NAND2_X1 U1001 ( .A1(n1271), .A2(n1272), .ZN(n1264) );
INV_X1 U1002 ( .A(KEYINPUT38), .ZN(n1272) );
NAND2_X1 U1003 ( .A1(n1273), .A2(n1274), .ZN(n1271) );
NAND3_X1 U1004 ( .A1(n1267), .A2(n1268), .A3(n1275), .ZN(n1274) );
INV_X1 U1005 ( .A(KEYINPUT56), .ZN(n1275) );
INV_X1 U1006 ( .A(n1075), .ZN(n1268) );
XOR2_X1 U1007 ( .A(G131), .B(KEYINPUT4), .Z(n1267) );
NAND2_X1 U1008 ( .A1(KEYINPUT56), .A2(n1075), .ZN(n1273) );
XOR2_X1 U1009 ( .A(G134), .B(G137), .Z(n1075) );
NAND2_X1 U1010 ( .A1(n1276), .A2(KEYINPUT35), .ZN(n1262) );
XNOR2_X1 U1011 ( .A(G140), .B(n1277), .ZN(n1276) );
NOR2_X1 U1012 ( .A1(G110), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U1013 ( .A(KEYINPUT63), .B(KEYINPUT42), .ZN(n1278) );
NAND2_X1 U1014 ( .A1(n1279), .A2(n988), .ZN(n1199) );
NAND3_X1 U1015 ( .A1(n1187), .A2(n1015), .A3(G952), .ZN(n988) );
XOR2_X1 U1016 ( .A(n1280), .B(KEYINPUT50), .Z(n1279) );
NAND3_X1 U1017 ( .A1(n1079), .A2(n1187), .A3(G902), .ZN(n1280) );
NAND2_X1 U1018 ( .A1(G237), .A2(G234), .ZN(n1187) );
NOR2_X1 U1019 ( .A1(G898), .A2(n1015), .ZN(n1079) );
AND2_X1 U1020 ( .A1(n1184), .A2(n1013), .ZN(n1011) );
NAND2_X1 U1021 ( .A1(G214), .A2(n1281), .ZN(n1013) );
NAND2_X1 U1022 ( .A1(n1282), .A2(n1038), .ZN(n1184) );
NAND2_X1 U1023 ( .A1(n1283), .A2(n1284), .ZN(n1038) );
XNOR2_X1 U1024 ( .A(KEYINPUT45), .B(n1037), .ZN(n1282) );
OR2_X1 U1025 ( .A1(n1284), .A2(n1283), .ZN(n1037) );
AND2_X1 U1026 ( .A1(n1285), .A2(n1233), .ZN(n1283) );
INV_X1 U1027 ( .A(G902), .ZN(n1233) );
XNOR2_X1 U1028 ( .A(n1139), .B(n1168), .ZN(n1285) );
XNOR2_X1 U1029 ( .A(n1166), .B(n1167), .ZN(n1168) );
XNOR2_X1 U1030 ( .A(n1067), .B(KEYINPUT13), .ZN(n1167) );
XOR2_X1 U1031 ( .A(G125), .B(KEYINPUT60), .Z(n1067) );
INV_X1 U1032 ( .A(n1076), .ZN(n1166) );
XOR2_X1 U1033 ( .A(G146), .B(n1223), .Z(n1076) );
XOR2_X1 U1034 ( .A(G128), .B(G143), .Z(n1223) );
XNOR2_X1 U1035 ( .A(n1286), .B(n1085), .ZN(n1139) );
XNOR2_X1 U1036 ( .A(n1287), .B(n1288), .ZN(n1085) );
XNOR2_X1 U1037 ( .A(n1125), .B(n1289), .ZN(n1288) );
XNOR2_X1 U1038 ( .A(n1227), .B(n1290), .ZN(n1289) );
NOR2_X1 U1039 ( .A1(KEYINPUT51), .A2(n1241), .ZN(n1290) );
XNOR2_X1 U1040 ( .A(n1197), .B(KEYINPUT16), .ZN(n1241) );
INV_X1 U1041 ( .A(G119), .ZN(n1197) );
XOR2_X1 U1042 ( .A(G116), .B(G122), .Z(n1227) );
XOR2_X1 U1043 ( .A(G101), .B(n1291), .Z(n1125) );
XOR2_X1 U1044 ( .A(G107), .B(G104), .Z(n1291) );
XOR2_X1 U1045 ( .A(n1292), .B(n1293), .Z(n1287) );
XOR2_X1 U1046 ( .A(KEYINPUT57), .B(G110), .Z(n1293) );
NAND2_X1 U1047 ( .A1(KEYINPUT12), .A2(n1198), .ZN(n1292) );
INV_X1 U1048 ( .A(G113), .ZN(n1198) );
NAND2_X1 U1049 ( .A1(G224), .A2(n1015), .ZN(n1286) );
INV_X1 U1050 ( .A(G953), .ZN(n1015) );
NAND2_X1 U1051 ( .A1(G210), .A2(n1281), .ZN(n1284) );
OR2_X1 U1052 ( .A1(G902), .A2(G237), .ZN(n1281) );
endmodule


