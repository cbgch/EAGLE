//Key = 1010111101101100101110100111110110001100111110100101001011001110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417;

XOR2_X1 U781 ( .A(G107), .B(n1094), .Z(G9) );
NOR2_X1 U782 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
XOR2_X1 U783 ( .A(n1097), .B(KEYINPUT52), .Z(n1095) );
NOR2_X1 U784 ( .A1(n1098), .A2(n1099), .ZN(G75) );
NOR4_X1 U785 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1099) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1104), .ZN(n1102) );
NAND3_X1 U787 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1101) );
NAND2_X1 U788 ( .A1(n1108), .A2(n1109), .ZN(n1106) );
NAND2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NAND3_X1 U790 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NAND2_X1 U791 ( .A1(n1115), .A2(n1116), .ZN(n1110) );
NAND2_X1 U792 ( .A1(n1117), .A2(n1118), .ZN(n1116) );
NAND3_X1 U793 ( .A1(n1113), .A2(n1119), .A3(n1120), .ZN(n1118) );
OR2_X1 U794 ( .A1(n1121), .A2(n1122), .ZN(n1119) );
NAND2_X1 U795 ( .A1(n1114), .A2(n1123), .ZN(n1117) );
NAND2_X1 U796 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NAND2_X1 U797 ( .A1(KEYINPUT25), .A2(n1126), .ZN(n1125) );
NAND2_X1 U798 ( .A1(n1127), .A2(n1128), .ZN(n1124) );
INV_X1 U799 ( .A(KEYINPUT59), .ZN(n1128) );
NAND4_X1 U800 ( .A1(n1115), .A2(n1129), .A3(n1114), .A4(n1130), .ZN(n1105) );
NAND2_X1 U801 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NAND2_X1 U802 ( .A1(n1126), .A2(n1133), .ZN(n1132) );
INV_X1 U803 ( .A(KEYINPUT25), .ZN(n1133) );
NAND2_X1 U804 ( .A1(KEYINPUT59), .A2(n1127), .ZN(n1131) );
NAND4_X1 U805 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1100) );
NAND3_X1 U806 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(n1135) );
XNOR2_X1 U807 ( .A(KEYINPUT39), .B(n1104), .ZN(n1139) );
NAND4_X1 U808 ( .A1(n1115), .A2(n1113), .A3(n1141), .A4(n1109), .ZN(n1104) );
NAND2_X1 U809 ( .A1(n1120), .A2(n1142), .ZN(n1134) );
XOR2_X1 U810 ( .A(KEYINPUT33), .B(n1143), .Z(n1142) );
NOR3_X1 U811 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(n1143) );
NAND3_X1 U812 ( .A1(n1147), .A2(n1109), .A3(n1113), .ZN(n1144) );
XOR2_X1 U813 ( .A(n1141), .B(KEYINPUT17), .Z(n1147) );
NOR3_X1 U814 ( .A1(n1148), .A2(G953), .A3(G952), .ZN(n1098) );
INV_X1 U815 ( .A(n1136), .ZN(n1148) );
NAND4_X1 U816 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1136) );
NOR4_X1 U817 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1152) );
XOR2_X1 U818 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U819 ( .A(n1159), .B(KEYINPUT34), .Z(n1158) );
NAND2_X1 U820 ( .A1(KEYINPUT31), .A2(n1160), .ZN(n1157) );
XOR2_X1 U821 ( .A(KEYINPUT50), .B(G472), .Z(n1160) );
XOR2_X1 U822 ( .A(KEYINPUT21), .B(n1161), .Z(n1154) );
NOR2_X1 U823 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NOR2_X1 U824 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
XNOR2_X1 U825 ( .A(n1166), .B(KEYINPUT15), .ZN(n1165) );
NOR2_X1 U826 ( .A1(n1167), .A2(n1168), .ZN(n1162) );
XNOR2_X1 U827 ( .A(KEYINPUT14), .B(n1169), .ZN(n1168) );
XOR2_X1 U828 ( .A(n1170), .B(G469), .Z(n1153) );
NAND2_X1 U829 ( .A1(KEYINPUT10), .A2(n1171), .ZN(n1170) );
NOR3_X1 U830 ( .A1(n1172), .A2(n1173), .A3(n1140), .ZN(n1151) );
INV_X1 U831 ( .A(n1174), .ZN(n1140) );
XOR2_X1 U832 ( .A(n1175), .B(n1176), .Z(n1149) );
NAND2_X1 U833 ( .A1(KEYINPUT2), .A2(n1177), .ZN(n1176) );
NAND2_X1 U834 ( .A1(n1178), .A2(n1179), .ZN(G72) );
NAND2_X1 U835 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
NAND2_X1 U836 ( .A1(n1182), .A2(n1183), .ZN(n1180) );
NAND2_X1 U837 ( .A1(KEYINPUT26), .A2(n1184), .ZN(n1183) );
NAND2_X1 U838 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
NAND2_X1 U839 ( .A1(KEYINPUT26), .A2(KEYINPUT44), .ZN(n1186) );
NAND3_X1 U840 ( .A1(KEYINPUT44), .A2(n1185), .A3(n1187), .ZN(n1178) );
INV_X1 U841 ( .A(n1181), .ZN(n1187) );
NAND2_X1 U842 ( .A1(n1188), .A2(n1189), .ZN(n1181) );
NAND3_X1 U843 ( .A1(n1190), .A2(n1191), .A3(n1192), .ZN(n1189) );
NAND2_X1 U844 ( .A1(G953), .A2(n1193), .ZN(n1191) );
NAND2_X1 U845 ( .A1(n1103), .A2(n1137), .ZN(n1190) );
XOR2_X1 U846 ( .A(KEYINPUT18), .B(n1194), .Z(n1188) );
NOR3_X1 U847 ( .A1(n1192), .A2(G953), .A3(n1195), .ZN(n1194) );
XNOR2_X1 U848 ( .A(n1196), .B(n1197), .ZN(n1192) );
XOR2_X1 U849 ( .A(n1198), .B(n1199), .Z(n1197) );
XOR2_X1 U850 ( .A(G140), .B(G125), .Z(n1199) );
NOR2_X1 U851 ( .A1(KEYINPUT55), .A2(n1200), .ZN(n1198) );
XOR2_X1 U852 ( .A(n1201), .B(n1202), .Z(n1196) );
INV_X1 U853 ( .A(n1184), .ZN(n1185) );
NAND2_X1 U854 ( .A1(G953), .A2(n1203), .ZN(n1184) );
NAND2_X1 U855 ( .A1(G900), .A2(G227), .ZN(n1203) );
NAND2_X1 U856 ( .A1(n1204), .A2(n1205), .ZN(G69) );
NAND2_X1 U857 ( .A1(n1206), .A2(n1137), .ZN(n1205) );
XOR2_X1 U858 ( .A(n1107), .B(n1207), .Z(n1206) );
NAND2_X1 U859 ( .A1(n1208), .A2(G953), .ZN(n1204) );
NAND2_X1 U860 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U861 ( .A1(n1207), .A2(n1211), .ZN(n1210) );
NAND2_X1 U862 ( .A1(G224), .A2(n1212), .ZN(n1209) );
NAND2_X1 U863 ( .A1(G898), .A2(n1207), .ZN(n1212) );
NAND2_X1 U864 ( .A1(n1213), .A2(n1214), .ZN(n1207) );
NAND2_X1 U865 ( .A1(G953), .A2(n1215), .ZN(n1214) );
XOR2_X1 U866 ( .A(n1216), .B(n1217), .Z(n1213) );
NOR2_X1 U867 ( .A1(n1218), .A2(n1219), .ZN(G66) );
XOR2_X1 U868 ( .A(n1220), .B(n1221), .Z(n1219) );
NAND2_X1 U869 ( .A1(n1222), .A2(n1223), .ZN(n1220) );
NOR2_X1 U870 ( .A1(n1218), .A2(n1224), .ZN(G63) );
XNOR2_X1 U871 ( .A(n1225), .B(n1226), .ZN(n1224) );
NOR3_X1 U872 ( .A1(n1227), .A2(KEYINPUT45), .A3(n1177), .ZN(n1226) );
NOR2_X1 U873 ( .A1(n1218), .A2(n1228), .ZN(G60) );
XOR2_X1 U874 ( .A(n1229), .B(n1230), .Z(n1228) );
NAND2_X1 U875 ( .A1(n1222), .A2(G475), .ZN(n1229) );
XOR2_X1 U876 ( .A(G104), .B(n1231), .Z(G6) );
NOR2_X1 U877 ( .A1(n1218), .A2(n1232), .ZN(G57) );
XNOR2_X1 U878 ( .A(n1233), .B(n1234), .ZN(n1232) );
XOR2_X1 U879 ( .A(n1235), .B(KEYINPUT58), .Z(n1234) );
NAND2_X1 U880 ( .A1(n1222), .A2(G472), .ZN(n1235) );
NOR2_X1 U881 ( .A1(n1218), .A2(n1236), .ZN(G54) );
XOR2_X1 U882 ( .A(n1237), .B(n1238), .Z(n1236) );
XOR2_X1 U883 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U884 ( .A1(n1222), .A2(G469), .ZN(n1240) );
NAND2_X1 U885 ( .A1(n1241), .A2(KEYINPUT19), .ZN(n1239) );
XOR2_X1 U886 ( .A(n1242), .B(n1243), .Z(n1241) );
NAND2_X1 U887 ( .A1(n1244), .A2(n1245), .ZN(n1237) );
NAND2_X1 U888 ( .A1(n1246), .A2(G110), .ZN(n1245) );
NAND2_X1 U889 ( .A1(n1247), .A2(n1248), .ZN(n1244) );
XOR2_X1 U890 ( .A(n1246), .B(KEYINPUT36), .Z(n1247) );
NOR2_X1 U891 ( .A1(n1137), .A2(G952), .ZN(n1218) );
NOR2_X1 U892 ( .A1(n1249), .A2(n1250), .ZN(G51) );
XOR2_X1 U893 ( .A(n1251), .B(n1252), .Z(n1250) );
XOR2_X1 U894 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U895 ( .A1(KEYINPUT30), .A2(n1255), .ZN(n1253) );
XOR2_X1 U896 ( .A(n1256), .B(n1257), .Z(n1251) );
XOR2_X1 U897 ( .A(G125), .B(n1258), .Z(n1257) );
NAND2_X1 U898 ( .A1(n1222), .A2(n1166), .ZN(n1256) );
INV_X1 U899 ( .A(n1169), .ZN(n1166) );
INV_X1 U900 ( .A(n1227), .ZN(n1222) );
NAND2_X1 U901 ( .A1(G902), .A2(n1259), .ZN(n1227) );
NAND2_X1 U902 ( .A1(n1107), .A2(n1195), .ZN(n1259) );
INV_X1 U903 ( .A(n1103), .ZN(n1195) );
NAND4_X1 U904 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1103) );
NOR4_X1 U905 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1263) );
NOR2_X1 U906 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NOR2_X1 U907 ( .A1(n1270), .A2(n1271), .ZN(n1266) );
NOR2_X1 U908 ( .A1(n1272), .A2(n1273), .ZN(n1265) );
AND2_X1 U909 ( .A1(n1274), .A2(KEYINPUT42), .ZN(n1264) );
AND3_X1 U910 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1262) );
NAND3_X1 U911 ( .A1(n1120), .A2(n1112), .A3(n1278), .ZN(n1261) );
NAND2_X1 U912 ( .A1(n1279), .A2(n1096), .ZN(n1260) );
NAND3_X1 U913 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1279) );
NAND3_X1 U914 ( .A1(n1115), .A2(n1269), .A3(n1278), .ZN(n1282) );
INV_X1 U915 ( .A(KEYINPUT49), .ZN(n1269) );
NAND3_X1 U916 ( .A1(n1283), .A2(n1273), .A3(n1284), .ZN(n1281) );
INV_X1 U917 ( .A(KEYINPUT56), .ZN(n1273) );
OR3_X1 U918 ( .A1(n1285), .A2(KEYINPUT42), .A3(n1270), .ZN(n1280) );
AND4_X1 U919 ( .A1(n1286), .A2(n1287), .A3(n1288), .A4(n1289), .ZN(n1107) );
NOR4_X1 U920 ( .A1(n1290), .A2(n1231), .A3(n1291), .A4(n1292), .ZN(n1289) );
NOR2_X1 U921 ( .A1(n1097), .A2(n1096), .ZN(n1292) );
NAND4_X1 U922 ( .A1(n1112), .A2(n1113), .A3(n1121), .A4(n1293), .ZN(n1097) );
NOR3_X1 U923 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(n1291) );
AND3_X1 U924 ( .A1(n1297), .A2(n1113), .A3(n1122), .ZN(n1231) );
NOR2_X1 U925 ( .A1(n1298), .A2(n1299), .ZN(n1288) );
NOR2_X1 U926 ( .A1(G952), .A2(n1300), .ZN(n1249) );
XNOR2_X1 U927 ( .A(G953), .B(KEYINPUT3), .ZN(n1300) );
XOR2_X1 U928 ( .A(G146), .B(n1274), .Z(G48) );
NOR3_X1 U929 ( .A1(n1285), .A2(n1096), .A3(n1270), .ZN(n1274) );
XNOR2_X1 U930 ( .A(G143), .B(n1272), .ZN(G45) );
NAND3_X1 U931 ( .A1(n1283), .A2(n1301), .A3(n1284), .ZN(n1272) );
INV_X1 U932 ( .A(n1294), .ZN(n1283) );
XOR2_X1 U933 ( .A(G140), .B(n1302), .Z(G42) );
NOR4_X1 U934 ( .A1(KEYINPUT24), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1302) );
XNOR2_X1 U935 ( .A(G137), .B(n1306), .ZN(G39) );
NAND4_X1 U936 ( .A1(KEYINPUT46), .A2(n1114), .A3(n1307), .A4(n1308), .ZN(n1306) );
AND3_X1 U937 ( .A1(n1155), .A2(n1309), .A3(n1310), .ZN(n1308) );
XNOR2_X1 U938 ( .A(n1112), .B(KEYINPUT20), .ZN(n1307) );
INV_X1 U939 ( .A(n1271), .ZN(n1114) );
NAND2_X1 U940 ( .A1(n1120), .A2(n1141), .ZN(n1271) );
XNOR2_X1 U941 ( .A(G134), .B(n1275), .ZN(G36) );
NAND3_X1 U942 ( .A1(n1120), .A2(n1121), .A3(n1284), .ZN(n1275) );
XNOR2_X1 U943 ( .A(G131), .B(n1277), .ZN(G33) );
NAND3_X1 U944 ( .A1(n1120), .A2(n1122), .A3(n1284), .ZN(n1277) );
AND3_X1 U945 ( .A1(n1112), .A2(n1310), .A3(n1127), .ZN(n1284) );
INV_X1 U946 ( .A(n1304), .ZN(n1120) );
NAND2_X1 U947 ( .A1(n1138), .A2(n1174), .ZN(n1304) );
XOR2_X1 U948 ( .A(n1311), .B(KEYINPUT22), .Z(n1138) );
NAND2_X1 U949 ( .A1(n1312), .A2(n1313), .ZN(G30) );
OR2_X1 U950 ( .A1(n1276), .A2(G128), .ZN(n1313) );
XOR2_X1 U951 ( .A(n1314), .B(KEYINPUT38), .Z(n1312) );
NAND2_X1 U952 ( .A1(G128), .A2(n1276), .ZN(n1314) );
NAND3_X1 U953 ( .A1(n1301), .A2(n1121), .A3(n1315), .ZN(n1276) );
INV_X1 U954 ( .A(n1270), .ZN(n1315) );
NAND4_X1 U955 ( .A1(n1112), .A2(n1155), .A3(n1310), .A4(n1309), .ZN(n1270) );
XNOR2_X1 U956 ( .A(n1316), .B(n1290), .ZN(G3) );
AND3_X1 U957 ( .A1(n1297), .A2(n1141), .A3(n1127), .ZN(n1290) );
XNOR2_X1 U958 ( .A(G125), .B(n1268), .ZN(G27) );
NAND3_X1 U959 ( .A1(n1115), .A2(n1301), .A3(n1278), .ZN(n1268) );
INV_X1 U960 ( .A(n1305), .ZN(n1278) );
NAND3_X1 U961 ( .A1(n1126), .A2(n1310), .A3(n1122), .ZN(n1305) );
NAND2_X1 U962 ( .A1(n1317), .A2(n1318), .ZN(n1310) );
NAND2_X1 U963 ( .A1(n1319), .A2(n1193), .ZN(n1318) );
INV_X1 U964 ( .A(G900), .ZN(n1193) );
XOR2_X1 U965 ( .A(G122), .B(n1320), .Z(G24) );
NOR3_X1 U966 ( .A1(n1321), .A2(n1295), .A3(n1296), .ZN(n1320) );
INV_X1 U967 ( .A(n1113), .ZN(n1295) );
NOR2_X1 U968 ( .A1(n1309), .A2(n1155), .ZN(n1113) );
XNOR2_X1 U969 ( .A(KEYINPUT43), .B(n1294), .ZN(n1321) );
NAND2_X1 U970 ( .A1(n1322), .A2(n1323), .ZN(n1294) );
XNOR2_X1 U971 ( .A(G119), .B(n1286), .ZN(G21) );
NAND4_X1 U972 ( .A1(n1324), .A2(n1141), .A3(n1155), .A4(n1309), .ZN(n1286) );
XNOR2_X1 U973 ( .A(G116), .B(n1287), .ZN(G18) );
NAND3_X1 U974 ( .A1(n1324), .A2(n1121), .A3(n1127), .ZN(n1287) );
XOR2_X1 U975 ( .A(G113), .B(n1299), .Z(G15) );
AND3_X1 U976 ( .A1(n1122), .A2(n1324), .A3(n1127), .ZN(n1299) );
AND2_X1 U977 ( .A1(n1325), .A2(n1309), .ZN(n1127) );
INV_X1 U978 ( .A(n1296), .ZN(n1324) );
NAND3_X1 U979 ( .A1(n1301), .A2(n1293), .A3(n1115), .ZN(n1296) );
NOR2_X1 U980 ( .A1(n1146), .A2(n1172), .ZN(n1115) );
INV_X1 U981 ( .A(n1145), .ZN(n1172) );
INV_X1 U982 ( .A(n1285), .ZN(n1122) );
NAND2_X1 U983 ( .A1(n1326), .A2(n1323), .ZN(n1285) );
XNOR2_X1 U984 ( .A(n1248), .B(n1298), .ZN(G12) );
AND3_X1 U985 ( .A1(n1126), .A2(n1141), .A3(n1297), .ZN(n1298) );
AND3_X1 U986 ( .A1(n1112), .A2(n1293), .A3(n1301), .ZN(n1297) );
INV_X1 U987 ( .A(n1096), .ZN(n1301) );
NAND2_X1 U988 ( .A1(n1311), .A2(n1174), .ZN(n1096) );
NAND2_X1 U989 ( .A1(G214), .A2(n1327), .ZN(n1174) );
NAND2_X1 U990 ( .A1(n1328), .A2(n1329), .ZN(n1311) );
NAND2_X1 U991 ( .A1(n1167), .A2(n1169), .ZN(n1329) );
XOR2_X1 U992 ( .A(KEYINPUT9), .B(n1330), .Z(n1328) );
NOR2_X1 U993 ( .A1(n1167), .A2(n1169), .ZN(n1330) );
NAND2_X1 U994 ( .A1(G210), .A2(n1327), .ZN(n1169) );
NAND2_X1 U995 ( .A1(n1331), .A2(n1332), .ZN(n1327) );
INV_X1 U996 ( .A(G237), .ZN(n1331) );
INV_X1 U997 ( .A(n1164), .ZN(n1167) );
NAND3_X1 U998 ( .A1(n1333), .A2(n1334), .A3(n1335), .ZN(n1164) );
NAND2_X1 U999 ( .A1(n1336), .A2(n1337), .ZN(n1334) );
XOR2_X1 U1000 ( .A(KEYINPUT63), .B(n1338), .Z(n1336) );
NAND2_X1 U1001 ( .A1(n1339), .A2(n1340), .ZN(n1333) );
INV_X1 U1002 ( .A(n1337), .ZN(n1340) );
XNOR2_X1 U1003 ( .A(n1341), .B(n1255), .ZN(n1337) );
XNOR2_X1 U1004 ( .A(G125), .B(KEYINPUT6), .ZN(n1341) );
XOR2_X1 U1005 ( .A(KEYINPUT51), .B(n1338), .Z(n1339) );
XOR2_X1 U1006 ( .A(n1258), .B(n1254), .Z(n1338) );
XNOR2_X1 U1007 ( .A(n1216), .B(n1342), .ZN(n1254) );
XNOR2_X1 U1008 ( .A(n1343), .B(KEYINPUT5), .ZN(n1342) );
NAND2_X1 U1009 ( .A1(KEYINPUT7), .A2(n1217), .ZN(n1343) );
XOR2_X1 U1010 ( .A(n1344), .B(n1345), .Z(n1216) );
XOR2_X1 U1011 ( .A(G122), .B(G113), .Z(n1345) );
XNOR2_X1 U1012 ( .A(n1346), .B(n1248), .ZN(n1344) );
NAND2_X1 U1013 ( .A1(KEYINPUT12), .A2(n1347), .ZN(n1346) );
NOR2_X1 U1014 ( .A1(n1211), .A2(G953), .ZN(n1258) );
INV_X1 U1015 ( .A(G224), .ZN(n1211) );
NAND2_X1 U1016 ( .A1(n1317), .A2(n1348), .ZN(n1293) );
NAND2_X1 U1017 ( .A1(n1319), .A2(n1215), .ZN(n1348) );
INV_X1 U1018 ( .A(G898), .ZN(n1215) );
NOR3_X1 U1019 ( .A1(n1332), .A2(n1130), .A3(n1137), .ZN(n1319) );
INV_X1 U1020 ( .A(n1109), .ZN(n1130) );
NAND3_X1 U1021 ( .A1(n1349), .A2(n1109), .A3(G952), .ZN(n1317) );
NAND2_X1 U1022 ( .A1(G237), .A2(G234), .ZN(n1109) );
XNOR2_X1 U1023 ( .A(KEYINPUT57), .B(n1137), .ZN(n1349) );
INV_X1 U1024 ( .A(n1303), .ZN(n1112) );
NAND2_X1 U1025 ( .A1(n1146), .A2(n1145), .ZN(n1303) );
NAND2_X1 U1026 ( .A1(G221), .A2(n1350), .ZN(n1145) );
XOR2_X1 U1027 ( .A(n1351), .B(n1171), .Z(n1146) );
NAND2_X1 U1028 ( .A1(n1335), .A2(n1352), .ZN(n1171) );
XOR2_X1 U1029 ( .A(n1353), .B(n1354), .Z(n1352) );
XOR2_X1 U1030 ( .A(n1246), .B(n1355), .Z(n1354) );
NOR2_X1 U1031 ( .A1(KEYINPUT11), .A2(n1356), .ZN(n1355) );
XOR2_X1 U1032 ( .A(n1242), .B(n1357), .Z(n1356) );
XNOR2_X1 U1033 ( .A(n1358), .B(KEYINPUT37), .ZN(n1357) );
NAND2_X1 U1034 ( .A1(KEYINPUT62), .A2(n1243), .ZN(n1358) );
XOR2_X1 U1035 ( .A(n1201), .B(n1217), .Z(n1242) );
XNOR2_X1 U1036 ( .A(n1316), .B(n1359), .ZN(n1217) );
XOR2_X1 U1037 ( .A(G107), .B(G104), .Z(n1359) );
INV_X1 U1038 ( .A(G101), .ZN(n1316) );
XNOR2_X1 U1039 ( .A(n1360), .B(n1361), .ZN(n1201) );
NAND2_X1 U1040 ( .A1(n1362), .A2(KEYINPUT61), .ZN(n1360) );
XNOR2_X1 U1041 ( .A(G146), .B(G143), .ZN(n1362) );
XNOR2_X1 U1042 ( .A(G140), .B(n1363), .ZN(n1246) );
AND2_X1 U1043 ( .A1(n1137), .A2(G227), .ZN(n1363) );
XNOR2_X1 U1044 ( .A(G110), .B(KEYINPUT4), .ZN(n1353) );
NAND2_X1 U1045 ( .A1(KEYINPUT60), .A2(G469), .ZN(n1351) );
NAND2_X1 U1046 ( .A1(n1364), .A2(n1365), .ZN(n1141) );
NAND2_X1 U1047 ( .A1(n1121), .A2(n1366), .ZN(n1365) );
NOR2_X1 U1048 ( .A1(n1323), .A2(n1326), .ZN(n1121) );
OR3_X1 U1049 ( .A1(n1323), .A2(n1322), .A3(n1366), .ZN(n1364) );
INV_X1 U1050 ( .A(KEYINPUT28), .ZN(n1366) );
INV_X1 U1051 ( .A(n1326), .ZN(n1322) );
XOR2_X1 U1052 ( .A(n1367), .B(n1177), .Z(n1326) );
INV_X1 U1053 ( .A(G478), .ZN(n1177) );
NAND2_X1 U1054 ( .A1(KEYINPUT41), .A2(n1175), .ZN(n1367) );
NAND2_X1 U1055 ( .A1(n1335), .A2(n1225), .ZN(n1175) );
XNOR2_X1 U1056 ( .A(n1368), .B(n1369), .ZN(n1225) );
XOR2_X1 U1057 ( .A(n1370), .B(n1371), .Z(n1369) );
NAND2_X1 U1058 ( .A1(KEYINPUT13), .A2(n1372), .ZN(n1371) );
XOR2_X1 U1059 ( .A(n1373), .B(n1374), .Z(n1372) );
XNOR2_X1 U1060 ( .A(n1375), .B(G128), .ZN(n1374) );
NOR2_X1 U1061 ( .A1(G134), .A2(KEYINPUT48), .ZN(n1373) );
NAND3_X1 U1062 ( .A1(G234), .A2(n1137), .A3(G217), .ZN(n1370) );
XOR2_X1 U1063 ( .A(n1376), .B(G107), .Z(n1368) );
NAND2_X1 U1064 ( .A1(n1377), .A2(KEYINPUT29), .ZN(n1376) );
XNOR2_X1 U1065 ( .A(G116), .B(G122), .ZN(n1377) );
NAND2_X1 U1066 ( .A1(n1378), .A2(n1150), .ZN(n1323) );
NAND2_X1 U1067 ( .A1(G475), .A2(n1379), .ZN(n1150) );
NAND2_X1 U1068 ( .A1(n1230), .A2(n1335), .ZN(n1379) );
XNOR2_X1 U1069 ( .A(n1173), .B(KEYINPUT1), .ZN(n1378) );
AND3_X1 U1070 ( .A1(n1335), .A2(n1380), .A3(n1230), .ZN(n1173) );
XOR2_X1 U1071 ( .A(n1381), .B(n1382), .Z(n1230) );
XOR2_X1 U1072 ( .A(n1383), .B(n1384), .Z(n1382) );
XNOR2_X1 U1073 ( .A(G113), .B(n1385), .ZN(n1384) );
NAND2_X1 U1074 ( .A1(n1386), .A2(KEYINPUT16), .ZN(n1385) );
XOR2_X1 U1075 ( .A(n1387), .B(n1202), .Z(n1386) );
XNOR2_X1 U1076 ( .A(n1388), .B(n1375), .ZN(n1387) );
NAND2_X1 U1077 ( .A1(n1389), .A2(G214), .ZN(n1388) );
XOR2_X1 U1078 ( .A(KEYINPUT32), .B(G122), .Z(n1383) );
XOR2_X1 U1079 ( .A(n1390), .B(n1391), .Z(n1381) );
XNOR2_X1 U1080 ( .A(n1392), .B(n1393), .ZN(n1390) );
NOR2_X1 U1081 ( .A1(G104), .A2(KEYINPUT35), .ZN(n1393) );
NOR2_X1 U1082 ( .A1(G140), .A2(KEYINPUT8), .ZN(n1392) );
INV_X1 U1083 ( .A(G475), .ZN(n1380) );
NOR2_X1 U1084 ( .A1(n1309), .A2(n1325), .ZN(n1126) );
INV_X1 U1085 ( .A(n1155), .ZN(n1325) );
XNOR2_X1 U1086 ( .A(n1394), .B(n1223), .ZN(n1155) );
AND2_X1 U1087 ( .A1(G217), .A2(n1350), .ZN(n1223) );
NAND2_X1 U1088 ( .A1(G234), .A2(n1332), .ZN(n1350) );
INV_X1 U1089 ( .A(G902), .ZN(n1332) );
NAND2_X1 U1090 ( .A1(n1221), .A2(n1335), .ZN(n1394) );
XOR2_X1 U1091 ( .A(n1395), .B(n1396), .Z(n1221) );
XOR2_X1 U1092 ( .A(n1397), .B(n1398), .Z(n1396) );
XOR2_X1 U1093 ( .A(G119), .B(n1399), .Z(n1398) );
AND3_X1 U1094 ( .A1(G221), .A2(n1137), .A3(G234), .ZN(n1399) );
INV_X1 U1095 ( .A(G953), .ZN(n1137) );
XNOR2_X1 U1096 ( .A(G140), .B(n1361), .ZN(n1397) );
INV_X1 U1097 ( .A(G128), .ZN(n1361) );
XNOR2_X1 U1098 ( .A(n1391), .B(n1400), .ZN(n1395) );
XNOR2_X1 U1099 ( .A(n1401), .B(n1402), .ZN(n1400) );
NOR2_X1 U1100 ( .A1(KEYINPUT23), .A2(n1248), .ZN(n1402) );
NAND2_X1 U1101 ( .A1(KEYINPUT54), .A2(n1403), .ZN(n1401) );
XOR2_X1 U1102 ( .A(G125), .B(G146), .Z(n1391) );
NAND2_X1 U1103 ( .A1(n1404), .A2(n1405), .ZN(n1309) );
OR2_X1 U1104 ( .A1(n1159), .A2(G472), .ZN(n1405) );
XOR2_X1 U1105 ( .A(n1406), .B(KEYINPUT53), .Z(n1404) );
NAND2_X1 U1106 ( .A1(G472), .A2(n1159), .ZN(n1406) );
NAND2_X1 U1107 ( .A1(n1407), .A2(n1335), .ZN(n1159) );
XNOR2_X1 U1108 ( .A(G902), .B(KEYINPUT47), .ZN(n1335) );
XNOR2_X1 U1109 ( .A(KEYINPUT0), .B(n1408), .ZN(n1407) );
INV_X1 U1110 ( .A(n1233), .ZN(n1408) );
XNOR2_X1 U1111 ( .A(n1409), .B(n1410), .ZN(n1233) );
XOR2_X1 U1112 ( .A(n1411), .B(n1412), .Z(n1410) );
XNOR2_X1 U1113 ( .A(G101), .B(G113), .ZN(n1412) );
NAND2_X1 U1114 ( .A1(n1389), .A2(G210), .ZN(n1411) );
NOR2_X1 U1115 ( .A1(G953), .A2(G237), .ZN(n1389) );
XOR2_X1 U1116 ( .A(n1413), .B(n1255), .Z(n1409) );
AND2_X1 U1117 ( .A1(n1414), .A2(n1415), .ZN(n1255) );
NAND2_X1 U1118 ( .A1(n1416), .A2(n1375), .ZN(n1415) );
INV_X1 U1119 ( .A(G143), .ZN(n1375) );
NAND2_X1 U1120 ( .A1(G143), .A2(n1417), .ZN(n1414) );
XOR2_X1 U1121 ( .A(n1416), .B(KEYINPUT40), .Z(n1417) );
XNOR2_X1 U1122 ( .A(G146), .B(G128), .ZN(n1416) );
XNOR2_X1 U1123 ( .A(n1347), .B(n1243), .ZN(n1413) );
XOR2_X1 U1124 ( .A(n1200), .B(n1202), .Z(n1243) );
XOR2_X1 U1125 ( .A(G131), .B(KEYINPUT27), .Z(n1202) );
XNOR2_X1 U1126 ( .A(G134), .B(n1403), .ZN(n1200) );
INV_X1 U1127 ( .A(G137), .ZN(n1403) );
XOR2_X1 U1128 ( .A(G116), .B(G119), .Z(n1347) );
INV_X1 U1129 ( .A(G110), .ZN(n1248) );
endmodule


