//Key = 0001111110111000111001100000001111110000100011101001010101111010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373;

NAND2_X1 U744 ( .A1(n1033), .A2(n1034), .ZN(G9) );
NAND2_X1 U745 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
XOR2_X1 U746 ( .A(n1037), .B(KEYINPUT14), .Z(n1033) );
NAND2_X1 U747 ( .A1(G107), .A2(n1038), .ZN(n1037) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(G75) );
NOR4_X1 U749 ( .A1(G953), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1040) );
NOR2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U752 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U757 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U758 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U759 ( .A1(n1062), .A2(n1063), .ZN(n1054) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
NOR3_X1 U761 ( .A1(n1063), .A2(n1066), .A3(n1057), .ZN(n1050) );
NOR2_X1 U762 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NOR2_X1 U763 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NOR4_X1 U764 ( .A1(n1071), .A2(n1057), .A3(n1053), .A4(n1063), .ZN(n1046) );
NOR2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR3_X1 U766 ( .A1(n1041), .A2(G953), .A3(G952), .ZN(n1039) );
AND4_X1 U767 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1041) );
NOR4_X1 U768 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
XNOR2_X1 U769 ( .A(n1082), .B(n1083), .ZN(n1081) );
NAND2_X1 U770 ( .A1(KEYINPUT35), .A2(n1084), .ZN(n1082) );
XNOR2_X1 U771 ( .A(n1085), .B(n1086), .ZN(n1080) );
NAND2_X1 U772 ( .A1(KEYINPUT60), .A2(n1087), .ZN(n1085) );
NOR3_X1 U773 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1076) );
NOR2_X1 U774 ( .A1(KEYINPUT18), .A2(n1091), .ZN(n1090) );
NOR3_X1 U775 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
AND2_X1 U776 ( .A1(n1053), .A2(KEYINPUT18), .ZN(n1089) );
INV_X1 U777 ( .A(n1095), .ZN(n1053) );
XOR2_X1 U778 ( .A(KEYINPUT42), .B(n1096), .Z(n1088) );
AND2_X1 U779 ( .A1(n1097), .A2(G475), .ZN(n1096) );
NAND2_X1 U780 ( .A1(n1098), .A2(n1099), .ZN(G72) );
NAND2_X1 U781 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
INV_X1 U783 ( .A(n1100), .ZN(n1103) );
NOR2_X1 U784 ( .A1(KEYINPUT28), .A2(n1104), .ZN(n1100) );
XOR2_X1 U785 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U786 ( .A1(n1107), .A2(G953), .ZN(n1106) );
NOR2_X1 U787 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1105) );
XOR2_X1 U789 ( .A(n1112), .B(n1113), .Z(n1110) );
XOR2_X1 U790 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U791 ( .A1(KEYINPUT55), .A2(n1116), .ZN(n1114) );
XOR2_X1 U792 ( .A(G125), .B(n1117), .Z(n1112) );
XOR2_X1 U793 ( .A(G140), .B(G137), .Z(n1117) );
NAND2_X1 U794 ( .A1(n1111), .A2(n1101), .ZN(n1102) );
NAND2_X1 U795 ( .A1(G953), .A2(n1118), .ZN(n1101) );
INV_X1 U796 ( .A(G227), .ZN(n1118) );
INV_X1 U797 ( .A(n1119), .ZN(n1111) );
XOR2_X1 U798 ( .A(n1120), .B(n1121), .Z(G69) );
XOR2_X1 U799 ( .A(n1122), .B(n1123), .Z(n1121) );
NOR2_X1 U800 ( .A1(G953), .A2(n1124), .ZN(n1123) );
NAND2_X1 U801 ( .A1(KEYINPUT3), .A2(n1125), .ZN(n1122) );
NAND2_X1 U802 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U803 ( .A(n1128), .B(n1129), .Z(n1126) );
NAND2_X1 U804 ( .A1(n1130), .A2(KEYINPUT10), .ZN(n1128) );
XOR2_X1 U805 ( .A(n1131), .B(n1132), .Z(n1130) );
XOR2_X1 U806 ( .A(n1133), .B(KEYINPUT13), .Z(n1131) );
NAND2_X1 U807 ( .A1(n1127), .A2(n1134), .ZN(n1120) );
NAND2_X1 U808 ( .A1(G953), .A2(n1135), .ZN(n1134) );
INV_X1 U809 ( .A(n1136), .ZN(n1127) );
NOR2_X1 U810 ( .A1(n1137), .A2(n1138), .ZN(G66) );
XOR2_X1 U811 ( .A(n1139), .B(n1140), .Z(n1138) );
NOR2_X1 U812 ( .A1(n1083), .A2(n1141), .ZN(n1140) );
NAND2_X1 U813 ( .A1(n1142), .A2(n1143), .ZN(n1139) );
XNOR2_X1 U814 ( .A(KEYINPUT50), .B(KEYINPUT25), .ZN(n1142) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1144), .ZN(G63) );
XOR2_X1 U816 ( .A(n1145), .B(n1146), .Z(n1144) );
AND2_X1 U817 ( .A1(G478), .A2(n1147), .ZN(n1145) );
NOR2_X1 U818 ( .A1(n1137), .A2(n1148), .ZN(G60) );
XNOR2_X1 U819 ( .A(n1149), .B(n1150), .ZN(n1148) );
NAND2_X1 U820 ( .A1(KEYINPUT45), .A2(n1151), .ZN(n1149) );
NAND2_X1 U821 ( .A1(n1147), .A2(G475), .ZN(n1151) );
XOR2_X1 U822 ( .A(G104), .B(n1152), .Z(G6) );
NOR2_X1 U823 ( .A1(n1137), .A2(n1153), .ZN(G57) );
NOR2_X1 U824 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U825 ( .A(n1156), .B(KEYINPUT16), .Z(n1155) );
NAND2_X1 U826 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XOR2_X1 U827 ( .A(KEYINPUT9), .B(n1159), .Z(n1158) );
NOR2_X1 U828 ( .A1(n1157), .A2(n1159), .ZN(n1154) );
XNOR2_X1 U829 ( .A(n1160), .B(n1161), .ZN(n1159) );
AND2_X1 U830 ( .A1(G472), .A2(n1147), .ZN(n1161) );
INV_X1 U831 ( .A(n1141), .ZN(n1147) );
NAND3_X1 U832 ( .A1(n1162), .A2(n1163), .A3(KEYINPUT32), .ZN(n1160) );
NAND3_X1 U833 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1163) );
INV_X1 U834 ( .A(KEYINPUT48), .ZN(n1166) );
NAND2_X1 U835 ( .A1(n1167), .A2(KEYINPUT48), .ZN(n1162) );
NOR2_X1 U836 ( .A1(n1137), .A2(n1168), .ZN(G54) );
XOR2_X1 U837 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U838 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U839 ( .A1(n1092), .A2(n1141), .ZN(n1172) );
INV_X1 U840 ( .A(G469), .ZN(n1092) );
NAND2_X1 U841 ( .A1(KEYINPUT53), .A2(n1173), .ZN(n1171) );
XOR2_X1 U842 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U843 ( .A1(KEYINPUT5), .A2(n1176), .ZN(n1175) );
NOR2_X1 U844 ( .A1(n1137), .A2(n1177), .ZN(G51) );
XOR2_X1 U845 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U846 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U847 ( .A1(n1087), .A2(n1141), .ZN(n1181) );
NAND2_X1 U848 ( .A1(G902), .A2(n1043), .ZN(n1141) );
NAND3_X1 U849 ( .A1(n1182), .A2(n1124), .A3(n1183), .ZN(n1043) );
XNOR2_X1 U850 ( .A(n1108), .B(KEYINPUT37), .ZN(n1183) );
AND2_X1 U851 ( .A1(n1184), .A2(n1185), .ZN(n1124) );
NOR4_X1 U852 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1035), .ZN(n1185) );
INV_X1 U853 ( .A(n1038), .ZN(n1035) );
NAND3_X1 U854 ( .A1(n1072), .A2(n1189), .A3(n1190), .ZN(n1038) );
NOR4_X1 U855 ( .A1(n1191), .A2(n1192), .A3(n1152), .A4(n1193), .ZN(n1184) );
NOR3_X1 U856 ( .A1(n1049), .A2(n1194), .A3(n1195), .ZN(n1193) );
AND3_X1 U857 ( .A1(n1190), .A2(n1189), .A3(n1073), .ZN(n1152) );
INV_X1 U858 ( .A(n1196), .ZN(n1192) );
INV_X1 U859 ( .A(n1109), .ZN(n1182) );
NAND4_X1 U860 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1109) );
NOR3_X1 U861 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
NAND2_X1 U862 ( .A1(n1204), .A2(n1205), .ZN(n1199) );
NAND2_X1 U863 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U864 ( .A1(n1068), .A2(n1208), .ZN(n1207) );
XNOR2_X1 U865 ( .A(KEYINPUT33), .B(n1209), .ZN(n1206) );
NAND2_X1 U866 ( .A1(KEYINPUT62), .A2(n1210), .ZN(n1180) );
INV_X1 U867 ( .A(G125), .ZN(n1210) );
NOR2_X1 U868 ( .A1(n1211), .A2(G952), .ZN(n1137) );
XOR2_X1 U869 ( .A(G953), .B(KEYINPUT21), .Z(n1211) );
XOR2_X1 U870 ( .A(n1212), .B(n1197), .Z(G48) );
NAND4_X1 U871 ( .A1(n1068), .A2(n1213), .A3(n1073), .A4(n1059), .ZN(n1197) );
XOR2_X1 U872 ( .A(n1214), .B(n1198), .Z(G45) );
NAND4_X1 U873 ( .A1(n1215), .A2(n1059), .A3(n1216), .A4(n1217), .ZN(n1198) );
XOR2_X1 U874 ( .A(n1218), .B(n1219), .Z(G42) );
NOR3_X1 U875 ( .A1(n1220), .A2(n1221), .A3(n1063), .ZN(n1219) );
XNOR2_X1 U876 ( .A(KEYINPUT20), .B(n1068), .ZN(n1220) );
NAND2_X1 U877 ( .A1(KEYINPUT59), .A2(n1222), .ZN(n1218) );
XOR2_X1 U878 ( .A(G137), .B(n1201), .Z(G39) );
AND4_X1 U879 ( .A1(n1213), .A2(n1223), .A3(n1068), .A4(n1204), .ZN(n1201) );
XNOR2_X1 U880 ( .A(n1203), .B(n1224), .ZN(G36) );
NOR2_X1 U881 ( .A1(G134), .A2(KEYINPUT43), .ZN(n1224) );
AND3_X1 U882 ( .A1(n1215), .A2(n1072), .A3(n1204), .ZN(n1203) );
XOR2_X1 U883 ( .A(G131), .B(n1225), .Z(G33) );
NOR2_X1 U884 ( .A1(n1063), .A2(n1209), .ZN(n1225) );
NAND2_X1 U885 ( .A1(n1215), .A2(n1073), .ZN(n1209) );
AND3_X1 U886 ( .A1(n1068), .A2(n1226), .A3(n1064), .ZN(n1215) );
XNOR2_X1 U887 ( .A(n1227), .B(KEYINPUT12), .ZN(n1068) );
INV_X1 U888 ( .A(n1204), .ZN(n1063) );
NOR2_X1 U889 ( .A1(n1060), .A2(n1079), .ZN(n1204) );
INV_X1 U890 ( .A(n1061), .ZN(n1079) );
XOR2_X1 U891 ( .A(n1228), .B(n1229), .Z(G30) );
NOR2_X1 U892 ( .A1(n1108), .A2(KEYINPUT15), .ZN(n1229) );
AND4_X1 U893 ( .A1(n1213), .A2(n1072), .A3(n1227), .A4(n1059), .ZN(n1108) );
AND3_X1 U894 ( .A1(n1230), .A2(n1226), .A3(n1231), .ZN(n1213) );
XOR2_X1 U895 ( .A(G101), .B(n1232), .Z(G3) );
NOR4_X1 U896 ( .A1(KEYINPUT1), .A2(n1194), .A3(n1195), .A4(n1049), .ZN(n1232) );
XOR2_X1 U897 ( .A(G125), .B(n1202), .Z(G27) );
AND3_X1 U898 ( .A1(n1208), .A2(n1059), .A3(n1095), .ZN(n1202) );
INV_X1 U899 ( .A(n1221), .ZN(n1208) );
NAND3_X1 U900 ( .A1(n1073), .A2(n1226), .A3(n1065), .ZN(n1221) );
NAND2_X1 U901 ( .A1(n1045), .A2(n1233), .ZN(n1226) );
NAND3_X1 U902 ( .A1(G902), .A2(n1234), .A3(n1119), .ZN(n1233) );
NOR2_X1 U903 ( .A1(G900), .A2(n1235), .ZN(n1119) );
XOR2_X1 U904 ( .A(G122), .B(n1188), .Z(G24) );
AND4_X1 U905 ( .A1(n1236), .A2(n1189), .A3(n1216), .A4(n1217), .ZN(n1188) );
INV_X1 U906 ( .A(n1057), .ZN(n1189) );
NAND2_X1 U907 ( .A1(n1237), .A2(n1238), .ZN(n1057) );
NAND2_X1 U908 ( .A1(n1239), .A2(n1240), .ZN(G21) );
NAND2_X1 U909 ( .A1(G119), .A2(n1196), .ZN(n1240) );
XOR2_X1 U910 ( .A(KEYINPUT31), .B(n1241), .Z(n1239) );
NOR2_X1 U911 ( .A1(G119), .A2(n1196), .ZN(n1241) );
NAND4_X1 U912 ( .A1(n1236), .A2(n1223), .A3(n1231), .A4(n1230), .ZN(n1196) );
XOR2_X1 U913 ( .A(G116), .B(n1187), .Z(G18) );
AND3_X1 U914 ( .A1(n1064), .A2(n1072), .A3(n1236), .ZN(n1187) );
NOR2_X1 U915 ( .A1(n1217), .A2(n1074), .ZN(n1072) );
INV_X1 U916 ( .A(n1242), .ZN(n1217) );
XOR2_X1 U917 ( .A(n1186), .B(n1243), .Z(G15) );
NOR2_X1 U918 ( .A1(KEYINPUT0), .A2(n1244), .ZN(n1243) );
AND3_X1 U919 ( .A1(n1064), .A2(n1073), .A3(n1236), .ZN(n1186) );
AND2_X1 U920 ( .A1(n1095), .A2(n1245), .ZN(n1236) );
NOR2_X1 U921 ( .A1(n1069), .A2(n1094), .ZN(n1095) );
INV_X1 U922 ( .A(n1070), .ZN(n1094) );
NOR2_X1 U923 ( .A1(n1216), .A2(n1242), .ZN(n1073) );
INV_X1 U924 ( .A(n1074), .ZN(n1216) );
INV_X1 U925 ( .A(n1195), .ZN(n1064) );
NAND2_X1 U926 ( .A1(n1237), .A2(n1231), .ZN(n1195) );
NAND3_X1 U927 ( .A1(n1246), .A2(n1247), .A3(n1248), .ZN(G12) );
NAND2_X1 U928 ( .A1(G110), .A2(n1249), .ZN(n1248) );
NAND2_X1 U929 ( .A1(KEYINPUT38), .A2(n1250), .ZN(n1247) );
NAND2_X1 U930 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
INV_X1 U931 ( .A(G110), .ZN(n1252) );
XOR2_X1 U932 ( .A(KEYINPUT19), .B(n1191), .Z(n1251) );
INV_X1 U933 ( .A(n1249), .ZN(n1191) );
NAND2_X1 U934 ( .A1(n1253), .A2(n1254), .ZN(n1246) );
INV_X1 U935 ( .A(KEYINPUT38), .ZN(n1254) );
NAND2_X1 U936 ( .A1(n1255), .A2(n1256), .ZN(n1253) );
OR3_X1 U937 ( .A1(n1249), .A2(G110), .A3(KEYINPUT19), .ZN(n1256) );
NAND2_X1 U938 ( .A1(KEYINPUT19), .A2(n1249), .ZN(n1255) );
NAND3_X1 U939 ( .A1(n1065), .A2(n1190), .A3(n1223), .ZN(n1249) );
INV_X1 U940 ( .A(n1049), .ZN(n1223) );
NAND2_X1 U941 ( .A1(n1074), .A2(n1242), .ZN(n1049) );
NOR2_X1 U942 ( .A1(n1257), .A2(n1078), .ZN(n1242) );
NOR2_X1 U943 ( .A1(n1097), .A2(G475), .ZN(n1078) );
AND2_X1 U944 ( .A1(n1258), .A2(n1097), .ZN(n1257) );
NAND2_X1 U945 ( .A1(n1150), .A2(n1259), .ZN(n1097) );
XNOR2_X1 U946 ( .A(n1260), .B(n1261), .ZN(n1150) );
XOR2_X1 U947 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U948 ( .A(G122), .B(G113), .Z(n1263) );
XOR2_X1 U949 ( .A(G143), .B(G125), .Z(n1262) );
XOR2_X1 U950 ( .A(n1264), .B(n1265), .Z(n1260) );
XNOR2_X1 U951 ( .A(G104), .B(n1266), .ZN(n1265) );
NAND2_X1 U952 ( .A1(n1267), .A2(G214), .ZN(n1266) );
XOR2_X1 U953 ( .A(n1268), .B(n1269), .Z(n1264) );
INV_X1 U954 ( .A(n1270), .ZN(n1269) );
NAND2_X1 U955 ( .A1(KEYINPUT7), .A2(G140), .ZN(n1268) );
XOR2_X1 U956 ( .A(KEYINPUT56), .B(G475), .Z(n1258) );
XOR2_X1 U957 ( .A(n1271), .B(G478), .Z(n1074) );
OR2_X1 U958 ( .A1(n1146), .A2(G902), .ZN(n1271) );
XNOR2_X1 U959 ( .A(n1272), .B(n1273), .ZN(n1146) );
XOR2_X1 U960 ( .A(G107), .B(n1274), .Z(n1273) );
XOR2_X1 U961 ( .A(G122), .B(G116), .Z(n1274) );
XOR2_X1 U962 ( .A(n1275), .B(n1276), .Z(n1272) );
AND3_X1 U963 ( .A1(G217), .A2(n1235), .A3(G234), .ZN(n1276) );
NAND2_X1 U964 ( .A1(KEYINPUT57), .A2(n1277), .ZN(n1275) );
XOR2_X1 U965 ( .A(n1116), .B(n1278), .Z(n1277) );
NAND2_X1 U966 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
XNOR2_X1 U967 ( .A(n1281), .B(KEYINPUT52), .ZN(n1279) );
INV_X1 U968 ( .A(G134), .ZN(n1116) );
INV_X1 U969 ( .A(n1194), .ZN(n1190) );
NAND2_X1 U970 ( .A1(n1245), .A2(n1227), .ZN(n1194) );
AND2_X1 U971 ( .A1(n1069), .A2(n1070), .ZN(n1227) );
NAND2_X1 U972 ( .A1(G221), .A2(n1282), .ZN(n1070) );
XOR2_X1 U973 ( .A(n1093), .B(G469), .Z(n1069) );
AND2_X1 U974 ( .A1(n1283), .A2(n1259), .ZN(n1093) );
NAND2_X1 U975 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
OR2_X1 U976 ( .A1(n1286), .A2(n1169), .ZN(n1285) );
XOR2_X1 U977 ( .A(n1287), .B(KEYINPUT49), .Z(n1284) );
NAND2_X1 U978 ( .A1(n1169), .A2(n1286), .ZN(n1287) );
XOR2_X1 U979 ( .A(n1174), .B(n1176), .Z(n1286) );
NAND2_X1 U980 ( .A1(G227), .A2(n1235), .ZN(n1174) );
XOR2_X1 U981 ( .A(n1288), .B(n1289), .Z(n1169) );
XOR2_X1 U982 ( .A(KEYINPUT39), .B(n1290), .Z(n1289) );
NOR2_X1 U983 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U984 ( .A(KEYINPUT54), .B(n1293), .Z(n1292) );
AND2_X1 U985 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
NOR2_X1 U986 ( .A1(n1294), .A2(n1295), .ZN(n1291) );
XNOR2_X1 U987 ( .A(n1296), .B(G104), .ZN(n1295) );
NAND2_X1 U988 ( .A1(KEYINPUT40), .A2(n1036), .ZN(n1296) );
XOR2_X1 U989 ( .A(n1115), .B(n1297), .Z(n1288) );
XOR2_X1 U990 ( .A(n1298), .B(n1299), .Z(n1115) );
NAND3_X1 U991 ( .A1(n1300), .A2(n1301), .A3(n1302), .ZN(n1298) );
XOR2_X1 U992 ( .A(n1303), .B(KEYINPUT30), .Z(n1302) );
NAND2_X1 U993 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND3_X1 U994 ( .A1(n1228), .A2(n1214), .A3(n1212), .ZN(n1305) );
NAND2_X1 U995 ( .A1(n1281), .A2(G146), .ZN(n1304) );
NAND3_X1 U996 ( .A1(G128), .A2(G143), .A3(n1212), .ZN(n1301) );
NAND2_X1 U997 ( .A1(n1306), .A2(G146), .ZN(n1300) );
AND2_X1 U998 ( .A1(n1059), .A2(n1307), .ZN(n1245) );
NAND2_X1 U999 ( .A1(n1045), .A2(n1308), .ZN(n1307) );
NAND3_X1 U1000 ( .A1(n1136), .A2(n1234), .A3(G902), .ZN(n1308) );
NOR2_X1 U1001 ( .A1(G898), .A2(n1235), .ZN(n1136) );
NAND3_X1 U1002 ( .A1(n1234), .A2(n1235), .A3(G952), .ZN(n1045) );
NAND2_X1 U1003 ( .A1(G237), .A2(G234), .ZN(n1234) );
AND2_X1 U1004 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1309), .ZN(n1061) );
XNOR2_X1 U1006 ( .A(n1310), .B(n1087), .ZN(n1060) );
NAND2_X1 U1007 ( .A1(G210), .A2(n1309), .ZN(n1087) );
NAND2_X1 U1008 ( .A1(n1311), .A2(n1259), .ZN(n1309) );
INV_X1 U1009 ( .A(G237), .ZN(n1311) );
XOR2_X1 U1010 ( .A(n1086), .B(KEYINPUT34), .Z(n1310) );
NAND2_X1 U1011 ( .A1(n1312), .A2(n1259), .ZN(n1086) );
XOR2_X1 U1012 ( .A(n1313), .B(n1314), .Z(n1312) );
XOR2_X1 U1013 ( .A(KEYINPUT6), .B(KEYINPUT24), .Z(n1314) );
XOR2_X1 U1014 ( .A(n1178), .B(G125), .Z(n1313) );
XOR2_X1 U1015 ( .A(n1315), .B(n1316), .Z(n1178) );
XOR2_X1 U1016 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1017 ( .A(n1212), .B(n1319), .Z(n1318) );
NOR2_X1 U1018 ( .A1(G953), .A2(n1135), .ZN(n1319) );
INV_X1 U1019 ( .A(G224), .ZN(n1135) );
NAND3_X1 U1020 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1317) );
NAND2_X1 U1021 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND2_X1 U1022 ( .A1(KEYINPUT58), .A2(n1325), .ZN(n1324) );
XOR2_X1 U1023 ( .A(KEYINPUT63), .B(n1326), .Z(n1325) );
NAND3_X1 U1024 ( .A1(KEYINPUT58), .A2(n1327), .A3(n1326), .ZN(n1321) );
INV_X1 U1025 ( .A(n1323), .ZN(n1327) );
XNOR2_X1 U1026 ( .A(n1132), .B(KEYINPUT8), .ZN(n1323) );
XNOR2_X1 U1027 ( .A(n1328), .B(n1329), .ZN(n1132) );
NOR2_X1 U1028 ( .A1(KEYINPUT47), .A2(n1330), .ZN(n1329) );
OR2_X1 U1029 ( .A1(n1326), .A2(KEYINPUT58), .ZN(n1320) );
INV_X1 U1030 ( .A(n1133), .ZN(n1326) );
XOR2_X1 U1031 ( .A(n1331), .B(n1332), .Z(n1133) );
XOR2_X1 U1032 ( .A(n1036), .B(n1333), .Z(n1332) );
XNOR2_X1 U1033 ( .A(KEYINPUT46), .B(KEYINPUT23), .ZN(n1333) );
INV_X1 U1034 ( .A(G107), .ZN(n1036) );
XNOR2_X1 U1035 ( .A(G104), .B(n1294), .ZN(n1331) );
XNOR2_X1 U1036 ( .A(n1334), .B(KEYINPUT22), .ZN(n1294) );
XOR2_X1 U1037 ( .A(n1335), .B(n1129), .Z(n1315) );
XOR2_X1 U1038 ( .A(G110), .B(G122), .Z(n1129) );
AND2_X1 U1039 ( .A1(n1238), .A2(n1230), .ZN(n1065) );
INV_X1 U1040 ( .A(n1237), .ZN(n1230) );
XOR2_X1 U1041 ( .A(n1083), .B(n1336), .Z(n1237) );
NOR2_X1 U1042 ( .A1(KEYINPUT29), .A2(n1084), .ZN(n1336) );
NAND2_X1 U1043 ( .A1(n1143), .A2(n1259), .ZN(n1084) );
XOR2_X1 U1044 ( .A(n1337), .B(n1338), .Z(n1143) );
XNOR2_X1 U1045 ( .A(n1176), .B(n1339), .ZN(n1338) );
XOR2_X1 U1046 ( .A(n1340), .B(n1341), .Z(n1339) );
NAND2_X1 U1047 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U1048 ( .A1(n1344), .A2(n1345), .ZN(n1343) );
INV_X1 U1049 ( .A(G137), .ZN(n1345) );
NAND2_X1 U1050 ( .A1(n1346), .A2(n1347), .ZN(n1344) );
NAND4_X1 U1051 ( .A1(KEYINPUT51), .A2(G221), .A3(G234), .A4(n1235), .ZN(n1347) );
NAND2_X1 U1052 ( .A1(n1348), .A2(n1349), .ZN(n1342) );
NAND3_X1 U1053 ( .A1(G234), .A2(n1235), .A3(G221), .ZN(n1349) );
INV_X1 U1054 ( .A(G953), .ZN(n1235) );
NAND2_X1 U1055 ( .A1(KEYINPUT51), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1056 ( .A1(G137), .A2(n1346), .ZN(n1350) );
INV_X1 U1057 ( .A(KEYINPUT27), .ZN(n1346) );
NAND2_X1 U1058 ( .A1(n1351), .A2(KEYINPUT11), .ZN(n1340) );
XOR2_X1 U1059 ( .A(G119), .B(n1228), .Z(n1351) );
XOR2_X1 U1060 ( .A(G110), .B(n1222), .Z(n1176) );
INV_X1 U1061 ( .A(G140), .ZN(n1222) );
XOR2_X1 U1062 ( .A(n1352), .B(n1353), .Z(n1337) );
NOR2_X1 U1063 ( .A1(KEYINPUT41), .A2(G125), .ZN(n1353) );
XOR2_X1 U1064 ( .A(n1212), .B(KEYINPUT61), .Z(n1352) );
NAND2_X1 U1065 ( .A1(G217), .A2(n1282), .ZN(n1083) );
NAND2_X1 U1066 ( .A1(G234), .A2(n1259), .ZN(n1282) );
XOR2_X1 U1067 ( .A(KEYINPUT17), .B(n1231), .Z(n1238) );
INV_X1 U1068 ( .A(n1075), .ZN(n1231) );
XOR2_X1 U1069 ( .A(n1354), .B(G472), .Z(n1075) );
NAND3_X1 U1070 ( .A1(n1355), .A2(n1356), .A3(n1259), .ZN(n1354) );
INV_X1 U1071 ( .A(G902), .ZN(n1259) );
NAND2_X1 U1072 ( .A1(n1357), .A2(n1358), .ZN(n1356) );
INV_X1 U1073 ( .A(KEYINPUT36), .ZN(n1358) );
XOR2_X1 U1074 ( .A(n1359), .B(n1157), .Z(n1357) );
AND2_X1 U1075 ( .A1(n1360), .A2(n1361), .ZN(n1157) );
NAND3_X1 U1076 ( .A1(G101), .A2(G210), .A3(n1267), .ZN(n1360) );
NAND2_X1 U1077 ( .A1(KEYINPUT36), .A2(n1362), .ZN(n1355) );
XOR2_X1 U1078 ( .A(n1167), .B(n1361), .Z(n1362) );
NAND2_X1 U1079 ( .A1(n1334), .A2(n1363), .ZN(n1361) );
NAND2_X1 U1080 ( .A1(n1267), .A2(G210), .ZN(n1363) );
NOR2_X1 U1081 ( .A1(G953), .A2(G237), .ZN(n1267) );
INV_X1 U1082 ( .A(G101), .ZN(n1334) );
INV_X1 U1083 ( .A(n1359), .ZN(n1167) );
XNOR2_X1 U1084 ( .A(n1164), .B(n1165), .ZN(n1359) );
XNOR2_X1 U1085 ( .A(n1330), .B(n1364), .ZN(n1165) );
NOR2_X1 U1086 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NOR3_X1 U1087 ( .A1(KEYINPUT44), .A2(G119), .A3(n1367), .ZN(n1366) );
AND2_X1 U1088 ( .A1(n1328), .A2(KEYINPUT44), .ZN(n1365) );
XOR2_X1 U1089 ( .A(n1367), .B(G119), .Z(n1328) );
INV_X1 U1090 ( .A(G116), .ZN(n1367) );
XNOR2_X1 U1091 ( .A(n1244), .B(KEYINPUT26), .ZN(n1330) );
INV_X1 U1092 ( .A(G113), .ZN(n1244) );
XNOR2_X1 U1093 ( .A(n1368), .B(n1335), .ZN(n1164) );
NAND2_X1 U1094 ( .A1(n1369), .A2(n1370), .ZN(n1335) );
NAND2_X1 U1095 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
INV_X1 U1096 ( .A(KEYINPUT4), .ZN(n1372) );
OR2_X1 U1097 ( .A1(n1281), .A2(n1306), .ZN(n1371) );
INV_X1 U1098 ( .A(n1280), .ZN(n1306) );
NAND2_X1 U1099 ( .A1(G128), .A2(n1214), .ZN(n1280) );
NOR2_X1 U1100 ( .A1(n1214), .A2(G128), .ZN(n1281) );
INV_X1 U1101 ( .A(G143), .ZN(n1214) );
NAND2_X1 U1102 ( .A1(KEYINPUT4), .A2(n1373), .ZN(n1369) );
XOR2_X1 U1103 ( .A(n1228), .B(G143), .Z(n1373) );
INV_X1 U1104 ( .A(G128), .ZN(n1228) );
XOR2_X1 U1105 ( .A(n1270), .B(n1297), .Z(n1368) );
XOR2_X1 U1106 ( .A(G134), .B(G137), .Z(n1297) );
XOR2_X1 U1107 ( .A(n1212), .B(n1299), .Z(n1270) );
XOR2_X1 U1108 ( .A(G131), .B(KEYINPUT2), .Z(n1299) );
INV_X1 U1109 ( .A(G146), .ZN(n1212) );
endmodule


