//Key = 0011100001001001111000011110111000000101011000000000010000011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
n1419, n1420, n1421, n1422, n1423, n1424;

XNOR2_X1 U778 ( .A(G107), .B(n1079), .ZN(G9) );
NOR2_X1 U779 ( .A1(n1080), .A2(n1081), .ZN(G75) );
NOR4_X1 U780 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1081) );
NOR2_X1 U781 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
XOR2_X1 U783 ( .A(KEYINPUT48), .B(n1090), .Z(n1089) );
NOR4_X1 U784 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
NAND2_X1 U785 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
NOR2_X1 U786 ( .A1(n1097), .A2(n1093), .ZN(n1088) );
NOR2_X1 U787 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U788 ( .A1(n1100), .A2(n1091), .ZN(n1099) );
NOR2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR3_X1 U791 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1103) );
NOR2_X1 U792 ( .A1(KEYINPUT17), .A2(n1108), .ZN(n1105) );
NOR2_X1 U793 ( .A1(n1109), .A2(n1108), .ZN(n1101) );
XNOR2_X1 U794 ( .A(n1110), .B(KEYINPUT35), .ZN(n1109) );
NOR3_X1 U795 ( .A1(n1104), .A2(n1111), .A3(n1108), .ZN(n1098) );
INV_X1 U796 ( .A(n1096), .ZN(n1108) );
NOR2_X1 U797 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND4_X1 U798 ( .A1(n1114), .A2(n1115), .A3(n1116), .A4(n1117), .ZN(n1082) );
NAND4_X1 U799 ( .A1(n1096), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1114) );
NOR2_X1 U800 ( .A1(n1091), .A2(n1093), .ZN(n1120) );
NAND2_X1 U801 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
NAND3_X1 U802 ( .A1(n1123), .A2(n1124), .A3(KEYINPUT17), .ZN(n1122) );
NOR3_X1 U803 ( .A1(n1125), .A2(G953), .A3(G952), .ZN(n1080) );
INV_X1 U804 ( .A(n1116), .ZN(n1125) );
NAND4_X1 U805 ( .A1(n1126), .A2(n1127), .A3(n1128), .A4(n1129), .ZN(n1116) );
NOR4_X1 U806 ( .A1(n1130), .A2(n1124), .A3(n1131), .A4(n1132), .ZN(n1129) );
XOR2_X1 U807 ( .A(n1123), .B(KEYINPUT3), .Z(n1131) );
NOR2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1128) );
XOR2_X1 U809 ( .A(n1135), .B(n1136), .Z(n1134) );
XNOR2_X1 U810 ( .A(KEYINPUT15), .B(n1137), .ZN(n1136) );
NOR2_X1 U811 ( .A1(n1138), .A2(KEYINPUT6), .ZN(n1135) );
XNOR2_X1 U812 ( .A(n1139), .B(n1140), .ZN(n1127) );
NAND2_X1 U813 ( .A1(KEYINPUT59), .A2(n1141), .ZN(n1139) );
XNOR2_X1 U814 ( .A(n1142), .B(n1143), .ZN(n1126) );
XNOR2_X1 U815 ( .A(KEYINPUT19), .B(n1144), .ZN(n1143) );
XOR2_X1 U816 ( .A(n1145), .B(n1146), .Z(G72) );
NOR2_X1 U817 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
XOR2_X1 U818 ( .A(n1149), .B(n1150), .Z(n1148) );
XNOR2_X1 U819 ( .A(n1151), .B(n1152), .ZN(n1150) );
XOR2_X1 U820 ( .A(n1153), .B(n1154), .Z(n1149) );
NOR2_X1 U821 ( .A1(KEYINPUT49), .A2(n1155), .ZN(n1154) );
XNOR2_X1 U822 ( .A(n1156), .B(KEYINPUT18), .ZN(n1155) );
XNOR2_X1 U823 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n1153) );
NOR2_X1 U824 ( .A1(n1157), .A2(n1117), .ZN(n1147) );
XNOR2_X1 U825 ( .A(G900), .B(KEYINPUT2), .ZN(n1157) );
NAND2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1145) );
NAND2_X1 U827 ( .A1(n1160), .A2(n1117), .ZN(n1159) );
NAND2_X1 U828 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
XOR2_X1 U829 ( .A(n1115), .B(KEYINPUT5), .Z(n1161) );
NAND2_X1 U830 ( .A1(G953), .A2(n1163), .ZN(n1158) );
NAND2_X1 U831 ( .A1(n1164), .A2(G227), .ZN(n1163) );
XNOR2_X1 U832 ( .A(G900), .B(KEYINPUT12), .ZN(n1164) );
XOR2_X1 U833 ( .A(n1165), .B(n1166), .Z(G69) );
NOR2_X1 U834 ( .A1(n1167), .A2(n1083), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1168), .A2(n1117), .ZN(n1167) );
NOR2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U837 ( .A1(KEYINPUT0), .A2(n1171), .ZN(n1165) );
NOR3_X1 U838 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1171) );
NOR2_X1 U839 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U840 ( .A(n1177), .B(n1178), .Z(n1176) );
XNOR2_X1 U841 ( .A(n1179), .B(n1180), .ZN(n1177) );
NOR2_X1 U842 ( .A1(n1181), .A2(n1182), .ZN(n1173) );
XNOR2_X1 U843 ( .A(n1183), .B(n1184), .ZN(n1182) );
NOR2_X1 U844 ( .A1(G898), .A2(n1117), .ZN(n1172) );
NOR2_X1 U845 ( .A1(n1185), .A2(n1186), .ZN(G66) );
XOR2_X1 U846 ( .A(n1187), .B(n1188), .Z(n1186) );
XOR2_X1 U847 ( .A(KEYINPUT21), .B(n1189), .Z(n1188) );
NOR2_X1 U848 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
NOR2_X1 U849 ( .A1(n1185), .A2(n1192), .ZN(G63) );
XOR2_X1 U850 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U851 ( .A(KEYINPUT4), .B(n1195), .Z(n1194) );
NOR2_X1 U852 ( .A1(n1144), .A2(n1191), .ZN(n1195) );
INV_X1 U853 ( .A(G478), .ZN(n1144) );
NOR2_X1 U854 ( .A1(n1185), .A2(n1196), .ZN(G60) );
XOR2_X1 U855 ( .A(n1197), .B(n1198), .Z(n1196) );
NOR2_X1 U856 ( .A1(n1199), .A2(n1191), .ZN(n1197) );
XNOR2_X1 U857 ( .A(G104), .B(n1200), .ZN(G6) );
NOR2_X1 U858 ( .A1(n1185), .A2(n1201), .ZN(G57) );
NOR2_X1 U859 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XOR2_X1 U860 ( .A(n1204), .B(KEYINPUT60), .Z(n1203) );
NAND2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
OR2_X1 U862 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NOR3_X1 U863 ( .A1(n1205), .A2(n1208), .A3(n1207), .ZN(n1202) );
AND2_X1 U864 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U865 ( .A(n1211), .B(KEYINPUT20), .Z(n1209) );
XOR2_X1 U866 ( .A(n1212), .B(n1213), .Z(n1205) );
XOR2_X1 U867 ( .A(n1214), .B(n1215), .Z(n1212) );
NOR2_X1 U868 ( .A1(n1137), .A2(n1191), .ZN(n1215) );
NAND2_X1 U869 ( .A1(n1216), .A2(KEYINPUT23), .ZN(n1214) );
XNOR2_X1 U870 ( .A(n1181), .B(KEYINPUT29), .ZN(n1216) );
NOR2_X1 U871 ( .A1(n1185), .A2(n1217), .ZN(G54) );
XOR2_X1 U872 ( .A(n1151), .B(n1218), .Z(n1217) );
XOR2_X1 U873 ( .A(n1219), .B(n1220), .Z(n1218) );
NOR2_X1 U874 ( .A1(n1140), .A2(n1191), .ZN(n1219) );
NOR2_X1 U875 ( .A1(n1185), .A2(n1221), .ZN(G51) );
XNOR2_X1 U876 ( .A(n1222), .B(n1223), .ZN(n1221) );
NOR2_X1 U877 ( .A1(n1224), .A2(n1191), .ZN(n1223) );
NAND2_X1 U878 ( .A1(G902), .A2(n1225), .ZN(n1191) );
NAND3_X1 U879 ( .A1(n1162), .A2(n1115), .A3(n1226), .ZN(n1225) );
INV_X1 U880 ( .A(n1083), .ZN(n1226) );
NAND4_X1 U881 ( .A1(n1200), .A2(n1227), .A3(n1079), .A4(n1228), .ZN(n1083) );
NOR4_X1 U882 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
INV_X1 U883 ( .A(n1233), .ZN(n1232) );
NOR3_X1 U884 ( .A1(n1234), .A2(KEYINPUT28), .A3(n1235), .ZN(n1230) );
NOR2_X1 U885 ( .A1(n1236), .A2(n1091), .ZN(n1229) );
NOR3_X1 U886 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1236) );
NOR2_X1 U887 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NOR3_X1 U888 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1238) );
NOR2_X1 U889 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
INV_X1 U890 ( .A(KEYINPUT27), .ZN(n1246) );
NOR3_X1 U891 ( .A1(n1247), .A2(n1248), .A3(n1249), .ZN(n1245) );
INV_X1 U892 ( .A(n1110), .ZN(n1249) );
NOR2_X1 U893 ( .A1(KEYINPUT27), .A2(n1250), .ZN(n1243) );
NOR2_X1 U894 ( .A1(n1235), .A2(n1251), .ZN(n1237) );
INV_X1 U895 ( .A(KEYINPUT28), .ZN(n1251) );
NAND3_X1 U896 ( .A1(n1250), .A2(n1112), .A3(n1096), .ZN(n1079) );
NAND3_X1 U897 ( .A1(n1096), .A2(n1250), .A3(n1113), .ZN(n1200) );
NAND2_X1 U898 ( .A1(n1252), .A2(n1253), .ZN(n1115) );
XOR2_X1 U899 ( .A(KEYINPUT46), .B(n1254), .Z(n1253) );
INV_X1 U900 ( .A(n1085), .ZN(n1162) );
NAND4_X1 U901 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1085) );
AND4_X1 U902 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1258) );
NAND3_X1 U903 ( .A1(n1252), .A2(n1263), .A3(n1264), .ZN(n1257) );
NOR2_X1 U904 ( .A1(n1117), .A2(G952), .ZN(n1185) );
XOR2_X1 U905 ( .A(n1265), .B(n1266), .Z(G48) );
NAND2_X1 U906 ( .A1(n1254), .A2(n1252), .ZN(n1266) );
AND2_X1 U907 ( .A1(n1267), .A2(n1113), .ZN(n1254) );
NAND2_X1 U908 ( .A1(KEYINPUT24), .A2(G146), .ZN(n1265) );
NAND3_X1 U909 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(G45) );
NAND2_X1 U910 ( .A1(G143), .A2(n1271), .ZN(n1270) );
NAND2_X1 U911 ( .A1(KEYINPUT57), .A2(n1272), .ZN(n1269) );
NAND2_X1 U912 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
XNOR2_X1 U913 ( .A(n1275), .B(G143), .ZN(n1274) );
INV_X1 U914 ( .A(n1271), .ZN(n1273) );
NAND2_X1 U915 ( .A1(n1276), .A2(n1277), .ZN(n1268) );
INV_X1 U916 ( .A(KEYINPUT57), .ZN(n1277) );
NAND2_X1 U917 ( .A1(n1278), .A2(n1279), .ZN(n1276) );
NAND2_X1 U918 ( .A1(G143), .A2(n1275), .ZN(n1279) );
OR3_X1 U919 ( .A1(n1271), .A2(G143), .A3(n1275), .ZN(n1278) );
INV_X1 U920 ( .A(KEYINPUT42), .ZN(n1275) );
NAND3_X1 U921 ( .A1(n1280), .A2(n1252), .A3(n1264), .ZN(n1271) );
XOR2_X1 U922 ( .A(n1263), .B(KEYINPUT43), .Z(n1280) );
XNOR2_X1 U923 ( .A(G140), .B(n1255), .ZN(G42) );
NAND3_X1 U924 ( .A1(n1281), .A2(n1110), .A3(n1282), .ZN(n1255) );
XNOR2_X1 U925 ( .A(G137), .B(n1256), .ZN(G39) );
NAND3_X1 U926 ( .A1(n1267), .A2(n1234), .A3(n1282), .ZN(n1256) );
NAND2_X1 U927 ( .A1(n1283), .A2(n1284), .ZN(G36) );
NAND2_X1 U928 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U929 ( .A1(G134), .A2(n1287), .ZN(n1283) );
NAND2_X1 U930 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U931 ( .A1(KEYINPUT58), .A2(n1290), .ZN(n1289) );
INV_X1 U932 ( .A(n1262), .ZN(n1290) );
OR2_X1 U933 ( .A1(n1285), .A2(KEYINPUT58), .ZN(n1288) );
NOR2_X1 U934 ( .A1(KEYINPUT55), .A2(n1262), .ZN(n1285) );
NAND3_X1 U935 ( .A1(n1282), .A2(n1112), .A3(n1264), .ZN(n1262) );
XNOR2_X1 U936 ( .A(G131), .B(n1261), .ZN(G33) );
NAND3_X1 U937 ( .A1(n1282), .A2(n1113), .A3(n1264), .ZN(n1261) );
AND3_X1 U938 ( .A1(n1110), .A2(n1291), .A3(n1106), .ZN(n1264) );
INV_X1 U939 ( .A(n1087), .ZN(n1282) );
NAND2_X1 U940 ( .A1(n1123), .A2(n1292), .ZN(n1087) );
XNOR2_X1 U941 ( .A(G128), .B(n1260), .ZN(G30) );
NAND3_X1 U942 ( .A1(n1112), .A2(n1252), .A3(n1267), .ZN(n1260) );
AND4_X1 U943 ( .A1(n1110), .A2(n1132), .A3(n1293), .A4(n1291), .ZN(n1267) );
NAND2_X1 U944 ( .A1(n1294), .A2(n1295), .ZN(G3) );
NAND2_X1 U945 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U946 ( .A(n1298), .B(n1299), .Z(n1294) );
NOR2_X1 U947 ( .A1(n1296), .A2(n1297), .ZN(n1299) );
INV_X1 U948 ( .A(KEYINPUT16), .ZN(n1297) );
XNOR2_X1 U949 ( .A(KEYINPUT13), .B(G101), .ZN(n1296) );
NAND3_X1 U950 ( .A1(n1106), .A2(n1250), .A3(n1234), .ZN(n1298) );
INV_X1 U951 ( .A(n1240), .ZN(n1250) );
XOR2_X1 U952 ( .A(n1259), .B(n1300), .Z(G27) );
NAND2_X1 U953 ( .A1(KEYINPUT9), .A2(G125), .ZN(n1300) );
NAND3_X1 U954 ( .A1(n1119), .A2(n1252), .A3(n1281), .ZN(n1259) );
AND3_X1 U955 ( .A1(n1113), .A2(n1291), .A3(n1107), .ZN(n1281) );
NAND2_X1 U956 ( .A1(n1093), .A2(n1301), .ZN(n1291) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1302), .A4(n1303), .ZN(n1301) );
INV_X1 U958 ( .A(G900), .ZN(n1303) );
INV_X1 U959 ( .A(n1304), .ZN(n1113) );
XNOR2_X1 U960 ( .A(G122), .B(n1233), .ZN(G24) );
NAND3_X1 U961 ( .A1(n1096), .A2(n1263), .A3(n1305), .ZN(n1233) );
NAND2_X1 U962 ( .A1(n1306), .A2(n1307), .ZN(n1263) );
NAND2_X1 U963 ( .A1(n1112), .A2(n1308), .ZN(n1307) );
INV_X1 U964 ( .A(KEYINPUT25), .ZN(n1308) );
NAND3_X1 U965 ( .A1(n1133), .A2(n1309), .A3(KEYINPUT25), .ZN(n1306) );
NOR2_X1 U966 ( .A1(n1293), .A2(n1132), .ZN(n1096) );
XNOR2_X1 U967 ( .A(n1310), .B(n1311), .ZN(G21) );
NOR2_X1 U968 ( .A1(n1235), .A2(n1091), .ZN(n1311) );
INV_X1 U969 ( .A(n1234), .ZN(n1091) );
NAND3_X1 U970 ( .A1(n1132), .A2(n1293), .A3(n1305), .ZN(n1235) );
INV_X1 U971 ( .A(n1312), .ZN(n1293) );
XNOR2_X1 U972 ( .A(G116), .B(n1227), .ZN(G18) );
NAND3_X1 U973 ( .A1(n1305), .A2(n1112), .A3(n1106), .ZN(n1227) );
NOR2_X1 U974 ( .A1(n1313), .A2(n1133), .ZN(n1112) );
NOR3_X1 U975 ( .A1(n1121), .A2(n1248), .A3(n1104), .ZN(n1305) );
XOR2_X1 U976 ( .A(G113), .B(n1231), .Z(G15) );
AND4_X1 U977 ( .A1(n1247), .A2(n1314), .A3(n1119), .A4(n1315), .ZN(n1231) );
NOR2_X1 U978 ( .A1(n1242), .A2(n1304), .ZN(n1315) );
NAND2_X1 U979 ( .A1(n1316), .A2(n1317), .ZN(n1304) );
XNOR2_X1 U980 ( .A(KEYINPUT40), .B(n1309), .ZN(n1317) );
XNOR2_X1 U981 ( .A(n1133), .B(KEYINPUT25), .ZN(n1316) );
INV_X1 U982 ( .A(n1106), .ZN(n1242) );
NOR2_X1 U983 ( .A1(n1132), .A2(n1312), .ZN(n1106) );
INV_X1 U984 ( .A(n1104), .ZN(n1119) );
NAND2_X1 U985 ( .A1(n1095), .A2(n1094), .ZN(n1104) );
NAND2_X1 U986 ( .A1(n1318), .A2(n1319), .ZN(G12) );
NAND4_X1 U987 ( .A1(n1234), .A2(n1107), .A3(n1320), .A4(n1321), .ZN(n1319) );
XOR2_X1 U988 ( .A(n1322), .B(KEYINPUT50), .Z(n1318) );
NAND2_X1 U989 ( .A1(G110), .A2(n1323), .ZN(n1322) );
NAND3_X1 U990 ( .A1(n1107), .A2(n1320), .A3(n1234), .ZN(n1323) );
NOR2_X1 U991 ( .A1(n1133), .A2(n1309), .ZN(n1234) );
INV_X1 U992 ( .A(n1313), .ZN(n1309) );
XOR2_X1 U993 ( .A(G478), .B(n1324), .Z(n1313) );
NOR2_X1 U994 ( .A1(n1142), .A2(KEYINPUT51), .ZN(n1324) );
AND2_X1 U995 ( .A1(n1193), .A2(n1325), .ZN(n1142) );
XNOR2_X1 U996 ( .A(n1326), .B(n1327), .ZN(n1193) );
XOR2_X1 U997 ( .A(n1328), .B(n1329), .Z(n1327) );
XNOR2_X1 U998 ( .A(n1286), .B(G128), .ZN(n1329) );
NOR2_X1 U999 ( .A1(KEYINPUT38), .A2(G143), .ZN(n1328) );
XOR2_X1 U1000 ( .A(n1330), .B(n1331), .Z(n1326) );
NOR2_X1 U1001 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
INV_X1 U1002 ( .A(G217), .ZN(n1332) );
NAND3_X1 U1003 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1330) );
NAND2_X1 U1004 ( .A1(G107), .A2(n1337), .ZN(n1336) );
NAND2_X1 U1005 ( .A1(n1338), .A2(KEYINPUT37), .ZN(n1337) );
XNOR2_X1 U1006 ( .A(KEYINPUT41), .B(n1339), .ZN(n1338) );
NAND3_X1 U1007 ( .A1(KEYINPUT45), .A2(n1340), .A3(n1341), .ZN(n1335) );
NAND2_X1 U1008 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
INV_X1 U1009 ( .A(KEYINPUT41), .ZN(n1342) );
NAND3_X1 U1010 ( .A1(n1344), .A2(n1345), .A3(n1339), .ZN(n1334) );
INV_X1 U1011 ( .A(n1341), .ZN(n1339) );
XOR2_X1 U1012 ( .A(G116), .B(n1346), .Z(n1341) );
INV_X1 U1013 ( .A(KEYINPUT45), .ZN(n1345) );
NAND2_X1 U1014 ( .A1(KEYINPUT41), .A2(n1343), .ZN(n1344) );
NAND2_X1 U1015 ( .A1(KEYINPUT37), .A2(n1347), .ZN(n1343) );
XOR2_X1 U1016 ( .A(n1348), .B(n1199), .Z(n1133) );
INV_X1 U1017 ( .A(G475), .ZN(n1199) );
OR2_X1 U1018 ( .A1(n1198), .A2(G902), .ZN(n1348) );
XNOR2_X1 U1019 ( .A(n1349), .B(n1350), .ZN(n1198) );
XNOR2_X1 U1020 ( .A(n1346), .B(n1351), .ZN(n1350) );
NOR2_X1 U1021 ( .A1(KEYINPUT31), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1022 ( .A(KEYINPUT7), .B(G113), .Z(n1352) );
XNOR2_X1 U1023 ( .A(n1353), .B(n1354), .ZN(n1349) );
NOR2_X1 U1024 ( .A1(G104), .A2(KEYINPUT8), .ZN(n1354) );
NOR2_X1 U1025 ( .A1(KEYINPUT56), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1026 ( .A(n1356), .B(n1357), .Z(n1355) );
XOR2_X1 U1027 ( .A(n1358), .B(n1359), .Z(n1357) );
AND2_X1 U1028 ( .A1(n1360), .A2(G214), .ZN(n1359) );
NAND2_X1 U1029 ( .A1(n1361), .A2(n1362), .ZN(n1358) );
NAND2_X1 U1030 ( .A1(G146), .A2(n1363), .ZN(n1362) );
XOR2_X1 U1031 ( .A(n1364), .B(KEYINPUT52), .Z(n1361) );
NAND2_X1 U1032 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
XNOR2_X1 U1033 ( .A(G131), .B(G143), .ZN(n1356) );
NAND2_X1 U1034 ( .A1(n1367), .A2(n1368), .ZN(n1320) );
OR2_X1 U1035 ( .A1(n1240), .A2(KEYINPUT61), .ZN(n1368) );
NAND3_X1 U1036 ( .A1(n1247), .A2(n1314), .A3(n1110), .ZN(n1240) );
NAND4_X1 U1037 ( .A1(n1110), .A2(n1247), .A3(n1248), .A4(KEYINPUT61), .ZN(n1367) );
INV_X1 U1038 ( .A(n1314), .ZN(n1248) );
NAND2_X1 U1039 ( .A1(n1093), .A2(n1369), .ZN(n1314) );
NAND4_X1 U1040 ( .A1(G953), .A2(G902), .A3(n1302), .A4(n1170), .ZN(n1369) );
INV_X1 U1041 ( .A(G898), .ZN(n1170) );
NAND3_X1 U1042 ( .A1(n1302), .A2(n1117), .A3(G952), .ZN(n1093) );
NAND2_X1 U1043 ( .A1(G237), .A2(G234), .ZN(n1302) );
XNOR2_X1 U1044 ( .A(n1121), .B(KEYINPUT22), .ZN(n1247) );
INV_X1 U1045 ( .A(n1252), .ZN(n1121) );
NOR2_X1 U1046 ( .A1(n1123), .A2(n1124), .ZN(n1252) );
INV_X1 U1047 ( .A(n1292), .ZN(n1124) );
NAND2_X1 U1048 ( .A1(G214), .A2(n1370), .ZN(n1292) );
XNOR2_X1 U1049 ( .A(n1371), .B(n1224), .ZN(n1123) );
NAND2_X1 U1050 ( .A1(G210), .A2(n1370), .ZN(n1224) );
NAND2_X1 U1051 ( .A1(n1372), .A2(n1325), .ZN(n1370) );
INV_X1 U1052 ( .A(G237), .ZN(n1372) );
NAND2_X1 U1053 ( .A1(n1222), .A2(n1325), .ZN(n1371) );
XNOR2_X1 U1054 ( .A(n1373), .B(n1374), .ZN(n1222) );
XOR2_X1 U1055 ( .A(n1375), .B(n1376), .Z(n1374) );
XOR2_X1 U1056 ( .A(G125), .B(n1377), .Z(n1376) );
NOR2_X1 U1057 ( .A1(KEYINPUT54), .A2(n1183), .ZN(n1377) );
XOR2_X1 U1058 ( .A(n1210), .B(n1178), .Z(n1183) );
AND2_X1 U1059 ( .A1(n1378), .A2(n1379), .ZN(n1178) );
NAND2_X1 U1060 ( .A1(KEYINPUT53), .A2(n1380), .ZN(n1379) );
OR3_X1 U1061 ( .A1(n1381), .A2(G107), .A3(KEYINPUT53), .ZN(n1378) );
NOR2_X1 U1062 ( .A1(G953), .A2(n1169), .ZN(n1375) );
INV_X1 U1063 ( .A(G224), .ZN(n1169) );
XOR2_X1 U1064 ( .A(n1382), .B(n1184), .Z(n1373) );
XNOR2_X1 U1065 ( .A(n1180), .B(n1383), .ZN(n1184) );
NAND2_X1 U1066 ( .A1(KEYINPUT26), .A2(n1346), .ZN(n1180) );
INV_X1 U1067 ( .A(G122), .ZN(n1346) );
XNOR2_X1 U1068 ( .A(n1181), .B(n1384), .ZN(n1382) );
NOR2_X1 U1069 ( .A1(n1095), .A2(n1130), .ZN(n1110) );
INV_X1 U1070 ( .A(n1094), .ZN(n1130) );
NAND2_X1 U1071 ( .A1(G221), .A2(n1385), .ZN(n1094) );
XOR2_X1 U1072 ( .A(n1141), .B(n1140), .Z(n1095) );
INV_X1 U1073 ( .A(G469), .ZN(n1140) );
AND2_X1 U1074 ( .A1(n1386), .A2(n1325), .ZN(n1141) );
XOR2_X1 U1075 ( .A(n1387), .B(n1388), .Z(n1386) );
XNOR2_X1 U1076 ( .A(n1220), .B(n1389), .ZN(n1388) );
NOR2_X1 U1077 ( .A1(KEYINPUT44), .A2(n1151), .ZN(n1389) );
XOR2_X1 U1078 ( .A(n1390), .B(n1391), .Z(n1151) );
NAND2_X1 U1079 ( .A1(n1392), .A2(n1393), .ZN(n1390) );
OR2_X1 U1080 ( .A1(n1394), .A2(G146), .ZN(n1393) );
XOR2_X1 U1081 ( .A(n1395), .B(KEYINPUT11), .Z(n1392) );
NAND2_X1 U1082 ( .A1(G146), .A2(n1394), .ZN(n1395) );
XOR2_X1 U1083 ( .A(G143), .B(KEYINPUT63), .Z(n1394) );
XNOR2_X1 U1084 ( .A(n1396), .B(n1397), .ZN(n1220) );
XNOR2_X1 U1085 ( .A(n1380), .B(n1398), .ZN(n1397) );
XOR2_X1 U1086 ( .A(G140), .B(n1399), .Z(n1398) );
AND2_X1 U1087 ( .A1(n1117), .A2(G227), .ZN(n1399) );
XNOR2_X1 U1088 ( .A(n1381), .B(n1347), .ZN(n1380) );
INV_X1 U1089 ( .A(G107), .ZN(n1347) );
INV_X1 U1090 ( .A(G104), .ZN(n1381) );
XNOR2_X1 U1091 ( .A(n1179), .B(n1400), .ZN(n1396) );
INV_X1 U1092 ( .A(n1156), .ZN(n1400) );
XNOR2_X1 U1093 ( .A(G101), .B(n1383), .ZN(n1179) );
XNOR2_X1 U1094 ( .A(KEYINPUT62), .B(KEYINPUT10), .ZN(n1387) );
INV_X1 U1095 ( .A(n1241), .ZN(n1107) );
NAND2_X1 U1096 ( .A1(n1312), .A2(n1132), .ZN(n1241) );
XOR2_X1 U1097 ( .A(n1401), .B(n1190), .Z(n1132) );
NAND2_X1 U1098 ( .A1(G217), .A2(n1385), .ZN(n1190) );
NAND2_X1 U1099 ( .A1(G234), .A2(n1325), .ZN(n1385) );
OR2_X1 U1100 ( .A1(n1187), .A2(G902), .ZN(n1401) );
XNOR2_X1 U1101 ( .A(n1402), .B(n1403), .ZN(n1187) );
XOR2_X1 U1102 ( .A(G137), .B(n1404), .Z(n1403) );
NOR2_X1 U1103 ( .A1(KEYINPUT1), .A2(n1405), .ZN(n1404) );
XOR2_X1 U1104 ( .A(n1406), .B(n1407), .Z(n1405) );
XNOR2_X1 U1105 ( .A(KEYINPUT47), .B(n1391), .ZN(n1407) );
INV_X1 U1106 ( .A(G128), .ZN(n1391) );
XNOR2_X1 U1107 ( .A(G119), .B(n1383), .ZN(n1406) );
XNOR2_X1 U1108 ( .A(n1321), .B(KEYINPUT36), .ZN(n1383) );
INV_X1 U1109 ( .A(G110), .ZN(n1321) );
XOR2_X1 U1110 ( .A(n1408), .B(n1409), .Z(n1402) );
NOR2_X1 U1111 ( .A1(n1333), .A2(n1410), .ZN(n1409) );
INV_X1 U1112 ( .A(G221), .ZN(n1410) );
NAND2_X1 U1113 ( .A1(G234), .A2(n1117), .ZN(n1333) );
INV_X1 U1114 ( .A(G953), .ZN(n1117) );
NAND3_X1 U1115 ( .A1(n1411), .A2(n1412), .A3(n1413), .ZN(n1408) );
OR2_X1 U1116 ( .A1(n1363), .A2(KEYINPUT39), .ZN(n1413) );
NAND3_X1 U1117 ( .A1(KEYINPUT39), .A2(n1414), .A3(n1366), .ZN(n1412) );
OR2_X1 U1118 ( .A1(n1366), .A2(n1414), .ZN(n1411) );
NOR2_X1 U1119 ( .A1(KEYINPUT34), .A2(n1365), .ZN(n1414) );
INV_X1 U1120 ( .A(n1363), .ZN(n1365) );
XOR2_X1 U1121 ( .A(n1152), .B(KEYINPUT14), .Z(n1363) );
XOR2_X1 U1122 ( .A(G125), .B(G140), .Z(n1152) );
XOR2_X1 U1123 ( .A(n1138), .B(n1137), .Z(n1312) );
INV_X1 U1124 ( .A(G472), .ZN(n1137) );
AND2_X1 U1125 ( .A1(n1415), .A2(n1325), .ZN(n1138) );
INV_X1 U1126 ( .A(G902), .ZN(n1325) );
XNOR2_X1 U1127 ( .A(n1416), .B(n1213), .ZN(n1415) );
XOR2_X1 U1128 ( .A(n1156), .B(n1384), .Z(n1213) );
XNOR2_X1 U1129 ( .A(n1417), .B(n1418), .ZN(n1384) );
XNOR2_X1 U1130 ( .A(KEYINPUT30), .B(n1366), .ZN(n1418) );
INV_X1 U1131 ( .A(G146), .ZN(n1366) );
XNOR2_X1 U1132 ( .A(G128), .B(G143), .ZN(n1417) );
XOR2_X1 U1133 ( .A(G131), .B(n1419), .Z(n1156) );
XNOR2_X1 U1134 ( .A(G137), .B(n1286), .ZN(n1419) );
INV_X1 U1135 ( .A(G134), .ZN(n1286) );
NAND3_X1 U1136 ( .A1(n1420), .A2(n1421), .A3(n1422), .ZN(n1416) );
NAND2_X1 U1137 ( .A1(n1207), .A2(n1181), .ZN(n1422) );
NOR2_X1 U1138 ( .A1(n1210), .A2(n1211), .ZN(n1207) );
NAND3_X1 U1139 ( .A1(n1175), .A2(n1211), .A3(G101), .ZN(n1421) );
INV_X1 U1140 ( .A(n1181), .ZN(n1175) );
NAND2_X1 U1141 ( .A1(n1423), .A2(n1210), .ZN(n1420) );
INV_X1 U1142 ( .A(G101), .ZN(n1210) );
XNOR2_X1 U1143 ( .A(n1211), .B(n1181), .ZN(n1423) );
XOR2_X1 U1144 ( .A(G113), .B(n1424), .Z(n1181) );
XNOR2_X1 U1145 ( .A(n1310), .B(G116), .ZN(n1424) );
INV_X1 U1146 ( .A(G119), .ZN(n1310) );
NAND2_X1 U1147 ( .A1(G210), .A2(n1360), .ZN(n1211) );
NOR2_X1 U1148 ( .A1(G953), .A2(G237), .ZN(n1360) );
endmodule


