//Key = 1000010011011000100001111001110100010001000001100010110010101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364;

XNOR2_X1 U746 ( .A(n1030), .B(n1031), .ZN(G9) );
NOR2_X1 U747 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U748 ( .A1(n1034), .A2(n1035), .ZN(G75) );
XOR2_X1 U749 ( .A(KEYINPUT14), .B(n1036), .Z(n1035) );
NOR3_X1 U750 ( .A1(n1037), .A2(G953), .A3(n1038), .ZN(n1036) );
INV_X1 U751 ( .A(n1039), .ZN(n1038) );
XNOR2_X1 U752 ( .A(KEYINPUT30), .B(n1040), .ZN(n1037) );
NOR3_X1 U753 ( .A1(n1041), .A2(n1040), .A3(n1042), .ZN(n1034) );
INV_X1 U754 ( .A(G952), .ZN(n1040) );
NAND3_X1 U755 ( .A1(n1039), .A2(n1043), .A3(n1044), .ZN(n1041) );
NAND2_X1 U756 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND3_X1 U758 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1048) );
NAND2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NAND2_X1 U760 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U761 ( .A1(n1056), .A2(n1033), .ZN(n1055) );
NAND2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1052) );
NAND2_X1 U763 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U764 ( .A1(n1057), .A2(n1061), .A3(n1054), .ZN(n1047) );
NAND3_X1 U765 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NAND2_X1 U766 ( .A1(n1049), .A2(n1065), .ZN(n1064) );
NAND2_X1 U767 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND3_X1 U768 ( .A1(G221), .A2(n1068), .A3(n1069), .ZN(n1067) );
NAND3_X1 U769 ( .A1(n1070), .A2(n1051), .A3(n1071), .ZN(n1062) );
INV_X1 U770 ( .A(n1072), .ZN(n1045) );
NAND4_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1039) );
NOR4_X1 U772 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
NOR2_X1 U773 ( .A1(G475), .A2(n1081), .ZN(n1079) );
INV_X1 U774 ( .A(n1082), .ZN(n1078) );
NOR2_X1 U775 ( .A1(n1083), .A2(n1084), .ZN(n1075) );
XOR2_X1 U776 ( .A(n1085), .B(n1086), .Z(n1084) );
NAND2_X1 U777 ( .A1(KEYINPUT23), .A2(G472), .ZN(n1086) );
XOR2_X1 U778 ( .A(n1087), .B(n1088), .Z(n1074) );
XOR2_X1 U779 ( .A(KEYINPUT15), .B(G478), .Z(n1088) );
XOR2_X1 U780 ( .A(n1089), .B(KEYINPUT20), .Z(n1073) );
XOR2_X1 U781 ( .A(n1090), .B(n1091), .Z(G72) );
XOR2_X1 U782 ( .A(n1092), .B(n1093), .Z(n1091) );
NAND2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U784 ( .A1(G953), .A2(n1096), .ZN(n1095) );
XOR2_X1 U785 ( .A(n1097), .B(n1098), .Z(n1094) );
XOR2_X1 U786 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U787 ( .A(KEYINPUT43), .B(n1101), .Z(n1100) );
NOR2_X1 U788 ( .A1(G131), .A2(KEYINPUT61), .ZN(n1099) );
XOR2_X1 U789 ( .A(n1102), .B(n1103), .Z(n1097) );
NAND2_X1 U790 ( .A1(n1104), .A2(n1043), .ZN(n1092) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1043), .ZN(n1090) );
NOR2_X1 U792 ( .A1(n1106), .A2(n1096), .ZN(n1105) );
NAND2_X1 U793 ( .A1(n1107), .A2(n1108), .ZN(G69) );
NAND2_X1 U794 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
OR2_X1 U795 ( .A1(n1043), .A2(G224), .ZN(n1110) );
NAND3_X1 U796 ( .A1(G953), .A2(n1111), .A3(n1112), .ZN(n1107) );
INV_X1 U797 ( .A(n1109), .ZN(n1112) );
XNOR2_X1 U798 ( .A(n1113), .B(n1114), .ZN(n1109) );
NOR2_X1 U799 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U800 ( .A(n1117), .B(n1118), .Z(n1116) );
XOR2_X1 U801 ( .A(KEYINPUT29), .B(G110), .Z(n1118) );
NOR2_X1 U802 ( .A1(G898), .A2(n1043), .ZN(n1115) );
NAND3_X1 U803 ( .A1(n1119), .A2(n1043), .A3(KEYINPUT9), .ZN(n1113) );
NAND2_X1 U804 ( .A1(n1120), .A2(n1121), .ZN(n1119) );
XOR2_X1 U805 ( .A(n1122), .B(KEYINPUT59), .Z(n1120) );
NAND2_X1 U806 ( .A1(G898), .A2(G224), .ZN(n1111) );
NOR2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(G66) );
XNOR2_X1 U808 ( .A(n1125), .B(n1126), .ZN(n1124) );
NAND2_X1 U809 ( .A1(KEYINPUT58), .A2(n1127), .ZN(n1125) );
NAND2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
XOR2_X1 U811 ( .A(KEYINPUT19), .B(G217), .Z(n1129) );
NOR2_X1 U812 ( .A1(n1123), .A2(n1130), .ZN(G63) );
NOR2_X1 U813 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U814 ( .A(n1133), .B(n1134), .Z(n1132) );
AND2_X1 U815 ( .A1(G478), .A2(n1128), .ZN(n1134) );
NOR2_X1 U816 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
XOR2_X1 U817 ( .A(KEYINPUT60), .B(n1137), .Z(n1136) );
INV_X1 U818 ( .A(KEYINPUT11), .ZN(n1135) );
NOR2_X1 U819 ( .A1(KEYINPUT11), .A2(n1138), .ZN(n1131) );
XNOR2_X1 U820 ( .A(n1137), .B(KEYINPUT60), .ZN(n1138) );
NOR3_X1 U821 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(G60) );
AND2_X1 U822 ( .A1(KEYINPUT5), .A2(n1123), .ZN(n1141) );
NOR3_X1 U823 ( .A1(KEYINPUT5), .A2(G953), .A3(G952), .ZN(n1140) );
XNOR2_X1 U824 ( .A(n1142), .B(n1143), .ZN(n1139) );
XOR2_X1 U825 ( .A(n1144), .B(KEYINPUT35), .Z(n1143) );
NAND3_X1 U826 ( .A1(G902), .A2(G475), .A3(n1145), .ZN(n1144) );
XOR2_X1 U827 ( .A(n1042), .B(KEYINPUT51), .Z(n1145) );
XNOR2_X1 U828 ( .A(n1146), .B(n1147), .ZN(G6) );
NOR2_X1 U829 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U830 ( .A1(n1123), .A2(n1150), .ZN(G57) );
XOR2_X1 U831 ( .A(n1151), .B(n1152), .Z(n1150) );
XOR2_X1 U832 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U833 ( .A1(KEYINPUT52), .A2(n1155), .ZN(n1153) );
XNOR2_X1 U834 ( .A(n1156), .B(n1157), .ZN(n1155) );
NAND2_X1 U835 ( .A1(KEYINPUT50), .A2(n1158), .ZN(n1156) );
XOR2_X1 U836 ( .A(KEYINPUT37), .B(n1159), .Z(n1151) );
AND2_X1 U837 ( .A1(G472), .A2(n1128), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1123), .A2(n1160), .ZN(G54) );
XOR2_X1 U839 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U840 ( .A(n1163), .B(n1158), .ZN(n1162) );
XOR2_X1 U841 ( .A(KEYINPUT41), .B(n1164), .Z(n1161) );
AND2_X1 U842 ( .A1(G469), .A2(n1128), .ZN(n1164) );
INV_X1 U843 ( .A(n1165), .ZN(n1128) );
NOR2_X1 U844 ( .A1(n1123), .A2(n1166), .ZN(G51) );
XOR2_X1 U845 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U846 ( .A(n1169), .B(n1157), .ZN(n1168) );
XNOR2_X1 U847 ( .A(n1170), .B(n1171), .ZN(n1167) );
NOR2_X1 U848 ( .A1(n1172), .A2(n1165), .ZN(n1171) );
NAND2_X1 U849 ( .A1(G902), .A2(n1042), .ZN(n1165) );
NAND3_X1 U850 ( .A1(n1121), .A2(n1122), .A3(n1173), .ZN(n1042) );
INV_X1 U851 ( .A(n1104), .ZN(n1173) );
NAND4_X1 U852 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1104) );
NOR4_X1 U853 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
NOR2_X1 U854 ( .A1(n1182), .A2(n1183), .ZN(n1176) );
OR3_X1 U855 ( .A1(n1184), .A2(n1033), .A3(n1080), .ZN(n1175) );
NAND2_X1 U856 ( .A1(n1185), .A2(n1186), .ZN(n1174) );
XOR2_X1 U857 ( .A(KEYINPUT3), .B(n1187), .Z(n1186) );
NOR4_X1 U858 ( .A1(n1056), .A2(n1059), .A3(n1083), .A4(n1188), .ZN(n1187) );
XNOR2_X1 U859 ( .A(KEYINPUT57), .B(n1189), .ZN(n1188) );
INV_X1 U860 ( .A(n1190), .ZN(n1059) );
NAND2_X1 U861 ( .A1(n1191), .A2(n1185), .ZN(n1122) );
XOR2_X1 U862 ( .A(n1149), .B(KEYINPUT24), .Z(n1191) );
NAND4_X1 U863 ( .A1(n1192), .A2(n1054), .A3(n1193), .A4(n1194), .ZN(n1149) );
AND4_X1 U864 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1121) );
NOR4_X1 U865 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NAND2_X1 U866 ( .A1(n1203), .A2(n1204), .ZN(n1197) );
XNOR2_X1 U867 ( .A(KEYINPUT34), .B(n1033), .ZN(n1204) );
INV_X1 U868 ( .A(n1032), .ZN(n1203) );
NAND2_X1 U869 ( .A1(n1054), .A2(n1205), .ZN(n1032) );
NAND3_X1 U870 ( .A1(n1205), .A2(n1057), .A3(n1190), .ZN(n1195) );
NOR2_X1 U871 ( .A1(n1043), .A2(G952), .ZN(n1123) );
XOR2_X1 U872 ( .A(G146), .B(n1182), .Z(G48) );
AND3_X1 U873 ( .A1(n1192), .A2(n1185), .A3(n1206), .ZN(n1182) );
XNOR2_X1 U874 ( .A(n1181), .B(n1207), .ZN(G45) );
XNOR2_X1 U875 ( .A(G143), .B(KEYINPUT17), .ZN(n1207) );
NOR4_X1 U876 ( .A1(n1184), .A2(n1148), .A3(n1208), .A4(n1209), .ZN(n1181) );
XOR2_X1 U877 ( .A(G140), .B(n1180), .Z(G42) );
NOR3_X1 U878 ( .A1(n1080), .A2(n1066), .A3(n1210), .ZN(n1180) );
NAND3_X1 U879 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(G39) );
OR2_X1 U880 ( .A1(n1214), .A2(KEYINPUT21), .ZN(n1213) );
NAND3_X1 U881 ( .A1(KEYINPUT21), .A2(n1214), .A3(n1183), .ZN(n1212) );
INV_X1 U882 ( .A(n1215), .ZN(n1183) );
NAND2_X1 U883 ( .A1(n1216), .A2(n1215), .ZN(n1211) );
NAND3_X1 U884 ( .A1(n1206), .A2(n1057), .A3(n1049), .ZN(n1215) );
INV_X1 U885 ( .A(n1080), .ZN(n1049) );
NAND2_X1 U886 ( .A1(n1217), .A2(KEYINPUT21), .ZN(n1216) );
XNOR2_X1 U887 ( .A(G137), .B(KEYINPUT7), .ZN(n1217) );
XOR2_X1 U888 ( .A(G134), .B(n1218), .Z(G36) );
NOR2_X1 U889 ( .A1(n1080), .A2(n1219), .ZN(n1218) );
XOR2_X1 U890 ( .A(KEYINPUT27), .B(n1220), .Z(n1219) );
NOR2_X1 U891 ( .A1(n1221), .A2(n1184), .ZN(n1220) );
XNOR2_X1 U892 ( .A(n1222), .B(KEYINPUT36), .ZN(n1221) );
XNOR2_X1 U893 ( .A(G131), .B(n1223), .ZN(G33) );
NAND2_X1 U894 ( .A1(KEYINPUT0), .A2(n1179), .ZN(n1223) );
NOR3_X1 U895 ( .A1(n1184), .A2(n1056), .A3(n1080), .ZN(n1179) );
NAND2_X1 U896 ( .A1(n1070), .A2(n1224), .ZN(n1080) );
NAND3_X1 U897 ( .A1(n1193), .A2(n1189), .A3(n1225), .ZN(n1184) );
XNOR2_X1 U898 ( .A(n1178), .B(n1226), .ZN(G30) );
NOR2_X1 U899 ( .A1(G128), .A2(KEYINPUT40), .ZN(n1226) );
AND3_X1 U900 ( .A1(n1222), .A2(n1185), .A3(n1206), .ZN(n1178) );
AND4_X1 U901 ( .A1(n1193), .A2(n1227), .A3(n1189), .A4(n1228), .ZN(n1206) );
XNOR2_X1 U902 ( .A(G101), .B(n1229), .ZN(G3) );
NAND2_X1 U903 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U904 ( .A1(KEYINPUT47), .A2(n1232), .ZN(n1231) );
OR2_X1 U905 ( .A1(KEYINPUT1), .A2(n1232), .ZN(n1230) );
INV_X1 U906 ( .A(n1196), .ZN(n1232) );
NAND3_X1 U907 ( .A1(n1205), .A2(n1057), .A3(n1225), .ZN(n1196) );
NOR3_X1 U908 ( .A1(n1148), .A2(n1233), .A3(n1066), .ZN(n1205) );
INV_X1 U909 ( .A(n1193), .ZN(n1066) );
XNOR2_X1 U910 ( .A(n1234), .B(n1235), .ZN(G27) );
NOR2_X1 U911 ( .A1(n1210), .A2(n1063), .ZN(n1235) );
NAND3_X1 U912 ( .A1(n1192), .A2(n1189), .A3(n1190), .ZN(n1210) );
NAND2_X1 U913 ( .A1(n1072), .A2(n1236), .ZN(n1189) );
NAND4_X1 U914 ( .A1(n1237), .A2(G953), .A3(G902), .A4(n1096), .ZN(n1236) );
INV_X1 U915 ( .A(G900), .ZN(n1096) );
XOR2_X1 U916 ( .A(n1238), .B(KEYINPUT42), .Z(n1237) );
NAND2_X1 U917 ( .A1(n1239), .A2(n1240), .ZN(G24) );
NAND2_X1 U918 ( .A1(n1201), .A2(n1241), .ZN(n1240) );
XOR2_X1 U919 ( .A(KEYINPUT39), .B(n1242), .Z(n1239) );
NOR2_X1 U920 ( .A1(n1201), .A2(n1241), .ZN(n1242) );
AND4_X1 U921 ( .A1(n1243), .A2(n1054), .A3(n1244), .A4(n1245), .ZN(n1201) );
NOR2_X1 U922 ( .A1(n1228), .A2(n1227), .ZN(n1054) );
XOR2_X1 U923 ( .A(n1246), .B(n1200), .Z(G21) );
AND4_X1 U924 ( .A1(n1243), .A2(n1057), .A3(n1227), .A4(n1228), .ZN(n1200) );
NAND2_X1 U925 ( .A1(KEYINPUT53), .A2(n1247), .ZN(n1246) );
NAND2_X1 U926 ( .A1(n1248), .A2(n1249), .ZN(G18) );
NAND2_X1 U927 ( .A1(G116), .A2(n1250), .ZN(n1249) );
XOR2_X1 U928 ( .A(n1251), .B(KEYINPUT49), .Z(n1248) );
NAND2_X1 U929 ( .A1(n1202), .A2(n1252), .ZN(n1251) );
INV_X1 U930 ( .A(n1250), .ZN(n1202) );
NAND3_X1 U931 ( .A1(n1225), .A2(n1222), .A3(n1243), .ZN(n1250) );
INV_X1 U932 ( .A(n1033), .ZN(n1222) );
NAND2_X1 U933 ( .A1(n1253), .A2(n1244), .ZN(n1033) );
XNOR2_X1 U934 ( .A(n1209), .B(KEYINPUT56), .ZN(n1253) );
XOR2_X1 U935 ( .A(G113), .B(n1199), .Z(G15) );
AND3_X1 U936 ( .A1(n1225), .A2(n1192), .A3(n1243), .ZN(n1199) );
NOR2_X1 U937 ( .A1(n1063), .A2(n1233), .ZN(n1243) );
INV_X1 U938 ( .A(n1194), .ZN(n1233) );
NAND2_X1 U939 ( .A1(n1051), .A2(n1185), .ZN(n1063) );
INV_X1 U940 ( .A(n1083), .ZN(n1051) );
NAND2_X1 U941 ( .A1(n1069), .A2(n1254), .ZN(n1083) );
NAND2_X1 U942 ( .A1(G221), .A2(n1068), .ZN(n1254) );
INV_X1 U943 ( .A(n1060), .ZN(n1225) );
NAND2_X1 U944 ( .A1(n1255), .A2(n1227), .ZN(n1060) );
XNOR2_X1 U945 ( .A(G110), .B(n1256), .ZN(G12) );
NAND4_X1 U946 ( .A1(n1190), .A2(n1193), .A3(n1257), .A4(n1258), .ZN(n1256) );
XNOR2_X1 U947 ( .A(KEYINPUT18), .B(n1148), .ZN(n1258) );
INV_X1 U948 ( .A(n1185), .ZN(n1148) );
NOR2_X1 U949 ( .A1(n1070), .A2(n1071), .ZN(n1185) );
INV_X1 U950 ( .A(n1224), .ZN(n1071) );
NAND2_X1 U951 ( .A1(G214), .A2(n1259), .ZN(n1224) );
XNOR2_X1 U952 ( .A(n1260), .B(n1172), .ZN(n1070) );
NAND2_X1 U953 ( .A1(G210), .A2(n1259), .ZN(n1172) );
NAND2_X1 U954 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
INV_X1 U955 ( .A(G237), .ZN(n1261) );
NAND2_X1 U956 ( .A1(n1263), .A2(n1262), .ZN(n1260) );
XOR2_X1 U957 ( .A(n1169), .B(n1264), .Z(n1263) );
XNOR2_X1 U958 ( .A(n1265), .B(n1266), .ZN(n1264) );
NAND2_X1 U959 ( .A1(KEYINPUT12), .A2(n1157), .ZN(n1266) );
NAND2_X1 U960 ( .A1(KEYINPUT8), .A2(n1170), .ZN(n1265) );
NAND2_X1 U961 ( .A1(G224), .A2(n1043), .ZN(n1170) );
XOR2_X1 U962 ( .A(n1117), .B(n1267), .Z(n1169) );
XOR2_X1 U963 ( .A(n1268), .B(n1269), .Z(n1117) );
XNOR2_X1 U964 ( .A(n1241), .B(G113), .ZN(n1269) );
XNOR2_X1 U965 ( .A(n1270), .B(n1271), .ZN(n1268) );
NAND3_X1 U966 ( .A1(n1272), .A2(n1273), .A3(n1274), .ZN(n1270) );
INV_X1 U967 ( .A(n1275), .ZN(n1274) );
NAND2_X1 U968 ( .A1(n1276), .A2(n1277), .ZN(n1273) );
INV_X1 U969 ( .A(KEYINPUT16), .ZN(n1277) );
XNOR2_X1 U970 ( .A(n1278), .B(n1279), .ZN(n1276) );
NOR2_X1 U971 ( .A1(G104), .A2(n1030), .ZN(n1279) );
NAND2_X1 U972 ( .A1(KEYINPUT16), .A2(n1280), .ZN(n1272) );
AND2_X1 U973 ( .A1(n1194), .A2(n1057), .ZN(n1257) );
NAND2_X1 U974 ( .A1(n1281), .A2(n1282), .ZN(n1057) );
OR2_X1 U975 ( .A1(n1056), .A2(KEYINPUT56), .ZN(n1282) );
INV_X1 U976 ( .A(n1192), .ZN(n1056) );
NOR2_X1 U977 ( .A1(n1244), .A2(n1209), .ZN(n1192) );
INV_X1 U978 ( .A(n1208), .ZN(n1244) );
NAND3_X1 U979 ( .A1(n1209), .A2(n1208), .A3(KEYINPUT56), .ZN(n1281) );
XNOR2_X1 U980 ( .A(n1087), .B(n1283), .ZN(n1208) );
NOR2_X1 U981 ( .A1(G478), .A2(KEYINPUT10), .ZN(n1283) );
NAND2_X1 U982 ( .A1(n1137), .A2(n1262), .ZN(n1087) );
XNOR2_X1 U983 ( .A(n1284), .B(n1285), .ZN(n1137) );
XOR2_X1 U984 ( .A(n1286), .B(n1287), .Z(n1285) );
NAND3_X1 U985 ( .A1(G217), .A2(n1043), .A3(G234), .ZN(n1287) );
NAND2_X1 U986 ( .A1(n1288), .A2(n1289), .ZN(n1286) );
NAND2_X1 U987 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XNOR2_X1 U988 ( .A(KEYINPUT31), .B(n1030), .ZN(n1291) );
XNOR2_X1 U989 ( .A(G116), .B(G122), .ZN(n1290) );
XOR2_X1 U990 ( .A(n1292), .B(KEYINPUT48), .Z(n1288) );
NAND2_X1 U991 ( .A1(n1293), .A2(n1294), .ZN(n1292) );
XNOR2_X1 U992 ( .A(n1241), .B(G116), .ZN(n1294) );
INV_X1 U993 ( .A(G122), .ZN(n1241) );
XNOR2_X1 U994 ( .A(KEYINPUT31), .B(G107), .ZN(n1293) );
XNOR2_X1 U995 ( .A(G128), .B(n1295), .ZN(n1284) );
XNOR2_X1 U996 ( .A(n1296), .B(G134), .ZN(n1295) );
INV_X1 U997 ( .A(n1245), .ZN(n1209) );
NAND2_X1 U998 ( .A1(n1297), .A2(n1089), .ZN(n1245) );
NAND2_X1 U999 ( .A1(G475), .A2(n1081), .ZN(n1089) );
OR2_X1 U1000 ( .A1(n1081), .A2(G475), .ZN(n1297) );
NAND2_X1 U1001 ( .A1(n1142), .A2(n1262), .ZN(n1081) );
XNOR2_X1 U1002 ( .A(n1298), .B(n1299), .ZN(n1142) );
XNOR2_X1 U1003 ( .A(n1146), .B(n1300), .ZN(n1299) );
XNOR2_X1 U1004 ( .A(KEYINPUT13), .B(n1301), .ZN(n1300) );
INV_X1 U1005 ( .A(G131), .ZN(n1301) );
XOR2_X1 U1006 ( .A(n1102), .B(n1302), .Z(n1298) );
XOR2_X1 U1007 ( .A(n1303), .B(n1304), .Z(n1302) );
AND2_X1 U1008 ( .A1(n1305), .A2(G214), .ZN(n1304) );
NOR2_X1 U1009 ( .A1(KEYINPUT4), .A2(n1306), .ZN(n1303) );
XOR2_X1 U1010 ( .A(G113), .B(n1307), .Z(n1306) );
NOR2_X1 U1011 ( .A1(G122), .A2(KEYINPUT26), .ZN(n1307) );
XNOR2_X1 U1012 ( .A(G125), .B(n1308), .ZN(n1102) );
NAND2_X1 U1013 ( .A1(n1072), .A2(n1309), .ZN(n1194) );
NAND4_X1 U1014 ( .A1(G953), .A2(G902), .A3(n1238), .A4(n1310), .ZN(n1309) );
INV_X1 U1015 ( .A(G898), .ZN(n1310) );
NAND3_X1 U1016 ( .A1(n1238), .A2(n1043), .A3(G952), .ZN(n1072) );
NAND2_X1 U1017 ( .A1(G237), .A2(G234), .ZN(n1238) );
NOR2_X1 U1018 ( .A1(n1069), .A2(n1311), .ZN(n1193) );
AND2_X1 U1019 ( .A1(G221), .A2(n1068), .ZN(n1311) );
XOR2_X1 U1020 ( .A(n1312), .B(G469), .Z(n1069) );
NAND2_X1 U1021 ( .A1(n1313), .A2(n1262), .ZN(n1312) );
XNOR2_X1 U1022 ( .A(n1314), .B(n1163), .ZN(n1313) );
XOR2_X1 U1023 ( .A(n1315), .B(n1316), .Z(n1163) );
XOR2_X1 U1024 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1025 ( .A(G110), .B(n1101), .Z(n1318) );
NOR2_X1 U1026 ( .A1(KEYINPUT32), .A2(n1319), .ZN(n1101) );
XOR2_X1 U1027 ( .A(KEYINPUT54), .B(G128), .Z(n1319) );
NOR2_X1 U1028 ( .A1(n1275), .A2(n1280), .ZN(n1317) );
NAND2_X1 U1029 ( .A1(n1320), .A2(n1321), .ZN(n1280) );
NAND3_X1 U1030 ( .A1(n1278), .A2(n1146), .A3(n1030), .ZN(n1321) );
INV_X1 U1031 ( .A(G107), .ZN(n1030) );
NAND2_X1 U1032 ( .A1(n1322), .A2(G107), .ZN(n1320) );
XNOR2_X1 U1033 ( .A(n1146), .B(G101), .ZN(n1322) );
NOR3_X1 U1034 ( .A1(n1146), .A2(G107), .A3(n1278), .ZN(n1275) );
INV_X1 U1035 ( .A(G104), .ZN(n1146) );
XNOR2_X1 U1036 ( .A(n1308), .B(n1323), .ZN(n1315) );
NOR2_X1 U1037 ( .A1(G953), .A2(n1106), .ZN(n1323) );
INV_X1 U1038 ( .A(G227), .ZN(n1106) );
XOR2_X1 U1039 ( .A(G143), .B(n1324), .Z(n1308) );
NAND2_X1 U1040 ( .A1(KEYINPUT45), .A2(n1158), .ZN(n1314) );
NOR2_X1 U1041 ( .A1(n1227), .A2(n1255), .ZN(n1190) );
INV_X1 U1042 ( .A(n1228), .ZN(n1255) );
NAND2_X1 U1043 ( .A1(n1325), .A2(n1082), .ZN(n1228) );
NAND3_X1 U1044 ( .A1(n1326), .A2(n1262), .A3(n1126), .ZN(n1082) );
XNOR2_X1 U1045 ( .A(n1077), .B(KEYINPUT6), .ZN(n1325) );
NOR2_X1 U1046 ( .A1(n1326), .A2(n1327), .ZN(n1077) );
AND2_X1 U1047 ( .A1(n1126), .A2(n1262), .ZN(n1327) );
XOR2_X1 U1048 ( .A(n1328), .B(n1329), .Z(n1126) );
XOR2_X1 U1049 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1050 ( .A(n1214), .B(G128), .ZN(n1331) );
INV_X1 U1051 ( .A(G137), .ZN(n1214) );
XOR2_X1 U1052 ( .A(KEYINPUT63), .B(KEYINPUT46), .Z(n1330) );
XOR2_X1 U1053 ( .A(n1332), .B(n1333), .Z(n1328) );
XOR2_X1 U1054 ( .A(n1334), .B(n1335), .Z(n1333) );
NOR2_X1 U1055 ( .A1(G119), .A2(KEYINPUT55), .ZN(n1335) );
AND3_X1 U1056 ( .A1(G221), .A2(n1043), .A3(G234), .ZN(n1334) );
INV_X1 U1057 ( .A(G953), .ZN(n1043) );
XNOR2_X1 U1058 ( .A(n1324), .B(n1267), .ZN(n1332) );
XNOR2_X1 U1059 ( .A(n1234), .B(G110), .ZN(n1267) );
INV_X1 U1060 ( .A(G125), .ZN(n1234) );
XNOR2_X1 U1061 ( .A(G140), .B(n1336), .ZN(n1324) );
NAND2_X1 U1062 ( .A1(n1337), .A2(n1068), .ZN(n1326) );
NAND2_X1 U1063 ( .A1(G234), .A2(n1262), .ZN(n1068) );
XOR2_X1 U1064 ( .A(KEYINPUT25), .B(G217), .Z(n1337) );
XNOR2_X1 U1065 ( .A(n1085), .B(G472), .ZN(n1227) );
NAND2_X1 U1066 ( .A1(n1338), .A2(n1262), .ZN(n1085) );
INV_X1 U1067 ( .A(G902), .ZN(n1262) );
XOR2_X1 U1068 ( .A(n1339), .B(n1154), .Z(n1338) );
XOR2_X1 U1069 ( .A(n1340), .B(n1341), .Z(n1154) );
XNOR2_X1 U1070 ( .A(G113), .B(n1278), .ZN(n1341) );
INV_X1 U1071 ( .A(G101), .ZN(n1278) );
XOR2_X1 U1072 ( .A(n1342), .B(n1343), .Z(n1340) );
NOR2_X1 U1073 ( .A1(KEYINPUT44), .A2(n1271), .ZN(n1343) );
XNOR2_X1 U1074 ( .A(n1247), .B(n1252), .ZN(n1271) );
INV_X1 U1075 ( .A(G116), .ZN(n1252) );
INV_X1 U1076 ( .A(G119), .ZN(n1247) );
NAND2_X1 U1077 ( .A1(G210), .A2(n1305), .ZN(n1342) );
NOR2_X1 U1078 ( .A1(G953), .A2(G237), .ZN(n1305) );
NAND2_X1 U1079 ( .A1(n1344), .A2(n1345), .ZN(n1339) );
NAND2_X1 U1080 ( .A1(n1346), .A2(n1158), .ZN(n1345) );
XOR2_X1 U1081 ( .A(KEYINPUT28), .B(n1347), .Z(n1344) );
NOR2_X1 U1082 ( .A1(n1158), .A2(n1346), .ZN(n1347) );
XNOR2_X1 U1083 ( .A(KEYINPUT22), .B(n1348), .ZN(n1346) );
INV_X1 U1084 ( .A(n1157), .ZN(n1348) );
XNOR2_X1 U1085 ( .A(n1349), .B(G128), .ZN(n1157) );
NAND3_X1 U1086 ( .A1(n1350), .A2(n1351), .A3(n1352), .ZN(n1349) );
NAND2_X1 U1087 ( .A1(n1336), .A2(n1353), .ZN(n1352) );
NAND3_X1 U1088 ( .A1(n1354), .A2(n1355), .A3(n1356), .ZN(n1353) );
NAND2_X1 U1089 ( .A1(KEYINPUT62), .A2(n1357), .ZN(n1356) );
NAND2_X1 U1090 ( .A1(KEYINPUT38), .A2(n1296), .ZN(n1355) );
NAND2_X1 U1091 ( .A1(n1358), .A2(n1359), .ZN(n1354) );
INV_X1 U1092 ( .A(KEYINPUT38), .ZN(n1359) );
NAND2_X1 U1093 ( .A1(n1296), .A2(n1360), .ZN(n1358) );
NAND2_X1 U1094 ( .A1(KEYINPUT33), .A2(n1361), .ZN(n1360) );
INV_X1 U1095 ( .A(n1362), .ZN(n1336) );
NAND4_X1 U1096 ( .A1(n1296), .A2(n1357), .A3(n1362), .A4(n1361), .ZN(n1351) );
INV_X1 U1097 ( .A(KEYINPUT62), .ZN(n1361) );
INV_X1 U1098 ( .A(KEYINPUT33), .ZN(n1357) );
NAND2_X1 U1099 ( .A1(KEYINPUT62), .A2(n1363), .ZN(n1350) );
NAND2_X1 U1100 ( .A1(n1296), .A2(n1364), .ZN(n1363) );
NAND2_X1 U1101 ( .A1(KEYINPUT33), .A2(n1362), .ZN(n1364) );
XOR2_X1 U1102 ( .A(G146), .B(KEYINPUT2), .Z(n1362) );
INV_X1 U1103 ( .A(G143), .ZN(n1296) );
XOR2_X1 U1104 ( .A(G131), .B(n1103), .Z(n1158) );
XOR2_X1 U1105 ( .A(G134), .B(G137), .Z(n1103) );
endmodule


