//Key = 1010011000010101110101001001110011101101110110000101000001110110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338;

NAND2_X1 U735 ( .A1(n1015), .A2(n1016), .ZN(G9) );
NAND2_X1 U736 ( .A1(G107), .A2(n1017), .ZN(n1016) );
NAND2_X1 U737 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
NAND2_X1 U738 ( .A1(KEYINPUT49), .A2(n1020), .ZN(n1019) );
OR2_X1 U739 ( .A1(n1021), .A2(KEYINPUT0), .ZN(n1018) );
NAND2_X1 U740 ( .A1(n1022), .A2(n1023), .ZN(n1015) );
NAND2_X1 U741 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NAND2_X1 U742 ( .A1(n1020), .A2(n1026), .ZN(n1025) );
INV_X1 U743 ( .A(KEYINPUT49), .ZN(n1026) );
XNOR2_X1 U744 ( .A(n1027), .B(KEYINPUT30), .ZN(n1020) );
NAND2_X1 U745 ( .A1(KEYINPUT0), .A2(n1027), .ZN(n1024) );
INV_X1 U746 ( .A(n1021), .ZN(n1027) );
NOR2_X1 U747 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR3_X1 U748 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1029) );
NAND3_X1 U749 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1030) );
NAND2_X1 U750 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND2_X1 U751 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NAND4_X1 U752 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1039) );
NOR2_X1 U753 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1046), .A2(n1047), .ZN(n1040) );
NAND2_X1 U755 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND3_X1 U756 ( .A1(n1048), .A2(n1050), .A3(n1051), .ZN(n1038) );
NAND2_X1 U757 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NAND4_X1 U758 ( .A1(n1054), .A2(n1042), .A3(n1055), .A4(n1056), .ZN(n1053) );
OR2_X1 U759 ( .A1(n1041), .A2(n1057), .ZN(n1056) );
NAND3_X1 U760 ( .A1(n1058), .A2(n1059), .A3(n1041), .ZN(n1055) );
NAND2_X1 U761 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U762 ( .A1(n1057), .A2(n1062), .ZN(n1052) );
NAND2_X1 U763 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NAND3_X1 U764 ( .A1(n1065), .A2(n1066), .A3(n1041), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1042), .A2(n1067), .ZN(n1066) );
NAND2_X1 U766 ( .A1(n1068), .A2(n1044), .ZN(n1065) );
INV_X1 U767 ( .A(n1069), .ZN(n1036) );
NOR3_X1 U768 ( .A1(n1070), .A2(G953), .A3(G952), .ZN(n1028) );
INV_X1 U769 ( .A(n1033), .ZN(n1070) );
NAND3_X1 U770 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1033) );
NOR4_X1 U771 ( .A1(n1074), .A2(n1060), .A3(n1075), .A4(n1076), .ZN(n1073) );
INV_X1 U772 ( .A(n1077), .ZN(n1060) );
NAND3_X1 U773 ( .A1(n1078), .A2(n1041), .A3(n1079), .ZN(n1074) );
NAND2_X1 U774 ( .A1(G469), .A2(n1080), .ZN(n1079) );
NAND2_X1 U775 ( .A1(G472), .A2(n1081), .ZN(n1078) );
NOR3_X1 U776 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1072) );
XOR2_X1 U777 ( .A(n1085), .B(KEYINPUT16), .Z(n1083) );
OR2_X1 U778 ( .A1(n1080), .A2(G469), .ZN(n1085) );
XNOR2_X1 U779 ( .A(n1086), .B(n1087), .ZN(n1082) );
NOR4_X1 U780 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1071) );
AND2_X1 U781 ( .A1(KEYINPUT40), .A2(n1092), .ZN(n1091) );
NOR2_X1 U782 ( .A1(KEYINPUT40), .A2(n1093), .ZN(n1090) );
NOR2_X1 U783 ( .A1(n1094), .A2(n1095), .ZN(n1089) );
NOR2_X1 U784 ( .A1(n1096), .A2(n1097), .ZN(n1088) );
NOR2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U786 ( .A1(KEYINPUT29), .A2(n1100), .ZN(n1099) );
AND2_X1 U787 ( .A1(n1095), .A2(KEYINPUT29), .ZN(n1098) );
OR2_X1 U788 ( .A1(KEYINPUT55), .A2(n1100), .ZN(n1095) );
XOR2_X1 U789 ( .A(n1101), .B(KEYINPUT54), .Z(n1100) );
XOR2_X1 U790 ( .A(n1102), .B(n1103), .Z(G72) );
XOR2_X1 U791 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U792 ( .A1(n1106), .A2(n1034), .ZN(n1105) );
XOR2_X1 U793 ( .A(n1107), .B(KEYINPUT19), .Z(n1106) );
NAND2_X1 U794 ( .A1(G900), .A2(G227), .ZN(n1107) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1104) );
NAND2_X1 U796 ( .A1(G953), .A2(n1110), .ZN(n1109) );
XOR2_X1 U797 ( .A(n1111), .B(n1112), .Z(n1108) );
NAND2_X1 U798 ( .A1(KEYINPUT43), .A2(n1113), .ZN(n1111) );
NAND2_X1 U799 ( .A1(n1034), .A2(n1031), .ZN(n1102) );
NAND2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(G69) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U802 ( .A1(G953), .A2(n1118), .ZN(n1117) );
NAND2_X1 U803 ( .A1(G898), .A2(G224), .ZN(n1118) );
NAND2_X1 U804 ( .A1(n1119), .A2(n1120), .ZN(n1114) );
NAND2_X1 U805 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NAND2_X1 U806 ( .A1(G953), .A2(n1123), .ZN(n1122) );
INV_X1 U807 ( .A(n1116), .ZN(n1119) );
XNOR2_X1 U808 ( .A(n1124), .B(n1125), .ZN(n1116) );
NOR2_X1 U809 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XNOR2_X1 U810 ( .A(KEYINPUT8), .B(n1034), .ZN(n1127) );
INV_X1 U811 ( .A(n1032), .ZN(n1126) );
NAND2_X1 U812 ( .A1(n1128), .A2(n1121), .ZN(n1124) );
INV_X1 U813 ( .A(n1129), .ZN(n1121) );
XOR2_X1 U814 ( .A(n1130), .B(n1131), .Z(n1128) );
XOR2_X1 U815 ( .A(n1132), .B(n1133), .Z(n1130) );
NAND2_X1 U816 ( .A1(KEYINPUT13), .A2(n1134), .ZN(n1132) );
NOR2_X1 U817 ( .A1(n1135), .A2(n1136), .ZN(G66) );
NOR3_X1 U818 ( .A1(n1101), .A2(n1137), .A3(n1138), .ZN(n1136) );
AND3_X1 U819 ( .A1(n1139), .A2(n1096), .A3(n1140), .ZN(n1138) );
INV_X1 U820 ( .A(n1094), .ZN(n1096) );
NOR2_X1 U821 ( .A1(n1141), .A2(n1139), .ZN(n1137) );
NOR2_X1 U822 ( .A1(n1142), .A2(n1094), .ZN(n1141) );
NOR2_X1 U823 ( .A1(n1031), .A2(n1032), .ZN(n1142) );
NOR2_X1 U824 ( .A1(n1135), .A2(n1143), .ZN(G63) );
XOR2_X1 U825 ( .A(n1144), .B(n1145), .Z(n1143) );
NAND2_X1 U826 ( .A1(n1140), .A2(G478), .ZN(n1145) );
NOR2_X1 U827 ( .A1(n1135), .A2(n1146), .ZN(G60) );
XOR2_X1 U828 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U829 ( .A(n1149), .B(KEYINPUT41), .Z(n1147) );
NAND2_X1 U830 ( .A1(n1140), .A2(G475), .ZN(n1149) );
XOR2_X1 U831 ( .A(n1150), .B(n1151), .Z(G6) );
NOR2_X1 U832 ( .A1(KEYINPUT38), .A2(n1152), .ZN(n1150) );
XNOR2_X1 U833 ( .A(KEYINPUT61), .B(n1153), .ZN(n1152) );
NOR3_X1 U834 ( .A1(n1135), .A2(n1154), .A3(n1155), .ZN(G57) );
NOR2_X1 U835 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
XNOR2_X1 U836 ( .A(n1158), .B(KEYINPUT22), .ZN(n1157) );
NOR2_X1 U837 ( .A1(G101), .A2(n1159), .ZN(n1154) );
XNOR2_X1 U838 ( .A(KEYINPUT14), .B(n1160), .ZN(n1159) );
INV_X1 U839 ( .A(n1158), .ZN(n1160) );
XNOR2_X1 U840 ( .A(n1161), .B(n1162), .ZN(n1158) );
XOR2_X1 U841 ( .A(n1163), .B(n1164), .Z(n1161) );
NAND2_X1 U842 ( .A1(n1140), .A2(G472), .ZN(n1163) );
NOR2_X1 U843 ( .A1(n1135), .A2(n1165), .ZN(G54) );
XOR2_X1 U844 ( .A(n1166), .B(n1167), .Z(n1165) );
NAND2_X1 U845 ( .A1(n1140), .A2(G469), .ZN(n1167) );
NAND2_X1 U846 ( .A1(n1168), .A2(n1169), .ZN(n1166) );
NAND2_X1 U847 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
XNOR2_X1 U848 ( .A(KEYINPUT3), .B(n1172), .ZN(n1170) );
XOR2_X1 U849 ( .A(n1173), .B(KEYINPUT56), .Z(n1168) );
NAND2_X1 U850 ( .A1(n1172), .A2(n1174), .ZN(n1173) );
XNOR2_X1 U851 ( .A(KEYINPUT26), .B(n1171), .ZN(n1174) );
NAND2_X1 U852 ( .A1(n1175), .A2(n1176), .ZN(n1171) );
NAND2_X1 U853 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XNOR2_X1 U854 ( .A(n1179), .B(KEYINPUT5), .ZN(n1177) );
XOR2_X1 U855 ( .A(n1180), .B(KEYINPUT53), .Z(n1175) );
NAND2_X1 U856 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U857 ( .A(KEYINPUT5), .B(n1183), .ZN(n1182) );
INV_X1 U858 ( .A(n1179), .ZN(n1183) );
XOR2_X1 U859 ( .A(n1184), .B(n1185), .Z(n1172) );
XNOR2_X1 U860 ( .A(n1186), .B(G110), .ZN(n1185) );
NOR2_X1 U861 ( .A1(n1187), .A2(n1188), .ZN(G51) );
XOR2_X1 U862 ( .A(KEYINPUT23), .B(n1135), .Z(n1188) );
NOR2_X1 U863 ( .A1(n1034), .A2(G952), .ZN(n1135) );
XOR2_X1 U864 ( .A(n1189), .B(n1190), .Z(n1187) );
XNOR2_X1 U865 ( .A(n1191), .B(n1192), .ZN(n1190) );
XNOR2_X1 U866 ( .A(n1193), .B(n1194), .ZN(n1189) );
NAND2_X1 U867 ( .A1(KEYINPUT44), .A2(n1195), .ZN(n1194) );
INV_X1 U868 ( .A(n1196), .ZN(n1195) );
NAND3_X1 U869 ( .A1(n1140), .A2(n1087), .A3(KEYINPUT15), .ZN(n1193) );
INV_X1 U870 ( .A(n1197), .ZN(n1087) );
AND2_X1 U871 ( .A1(G902), .A2(n1198), .ZN(n1140) );
OR2_X1 U872 ( .A1(n1032), .A2(n1031), .ZN(n1198) );
NAND4_X1 U873 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1031) );
NOR4_X1 U874 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1202) );
INV_X1 U875 ( .A(n1207), .ZN(n1206) );
NAND2_X1 U876 ( .A1(n1208), .A2(n1209), .ZN(n1201) );
NAND2_X1 U877 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
OR2_X1 U878 ( .A1(n1212), .A2(n1059), .ZN(n1211) );
NAND4_X1 U879 ( .A1(n1213), .A2(n1021), .A3(n1214), .A4(n1215), .ZN(n1032) );
NOR4_X1 U880 ( .A1(n1216), .A2(n1217), .A3(n1151), .A4(n1218), .ZN(n1215) );
NOR4_X1 U881 ( .A1(n1219), .A2(n1059), .A3(n1046), .A4(n1063), .ZN(n1218) );
INV_X1 U882 ( .A(n1220), .ZN(n1046) );
XOR2_X1 U883 ( .A(n1221), .B(KEYINPUT21), .Z(n1219) );
AND3_X1 U884 ( .A1(n1051), .A2(n1222), .A3(n1223), .ZN(n1151) );
AND2_X1 U885 ( .A1(n1224), .A2(n1225), .ZN(n1214) );
NAND3_X1 U886 ( .A1(n1051), .A2(n1222), .A3(n1208), .ZN(n1021) );
XOR2_X1 U887 ( .A(G146), .B(n1205), .Z(G48) );
NOR3_X1 U888 ( .A1(n1226), .A2(n1059), .A3(n1212), .ZN(n1205) );
XOR2_X1 U889 ( .A(G143), .B(n1227), .Z(G45) );
NOR2_X1 U890 ( .A1(KEYINPUT46), .A2(n1199), .ZN(n1227) );
NAND4_X1 U891 ( .A1(n1228), .A2(n1229), .A3(n1220), .A4(n1230), .ZN(n1199) );
NAND2_X1 U892 ( .A1(n1231), .A2(n1232), .ZN(G42) );
NAND2_X1 U893 ( .A1(G140), .A2(n1200), .ZN(n1232) );
XOR2_X1 U894 ( .A(n1233), .B(KEYINPUT48), .Z(n1231) );
OR2_X1 U895 ( .A1(n1200), .A2(G140), .ZN(n1233) );
NAND3_X1 U896 ( .A1(n1228), .A2(n1057), .A3(n1234), .ZN(n1200) );
NOR3_X1 U897 ( .A1(n1226), .A2(n1051), .A3(n1235), .ZN(n1234) );
XOR2_X1 U898 ( .A(G137), .B(n1204), .Z(G39) );
NOR3_X1 U899 ( .A1(n1045), .A2(n1044), .A3(n1212), .ZN(n1204) );
INV_X1 U900 ( .A(n1054), .ZN(n1044) );
XOR2_X1 U901 ( .A(G134), .B(n1236), .Z(G36) );
NOR3_X1 U902 ( .A1(n1210), .A2(KEYINPUT42), .A3(n1067), .ZN(n1236) );
XOR2_X1 U903 ( .A(G131), .B(n1203), .Z(G33) );
NOR2_X1 U904 ( .A1(n1210), .A2(n1226), .ZN(n1203) );
INV_X1 U905 ( .A(n1223), .ZN(n1226) );
NAND3_X1 U906 ( .A1(n1057), .A2(n1220), .A3(n1228), .ZN(n1210) );
INV_X1 U907 ( .A(n1045), .ZN(n1057) );
NAND2_X1 U908 ( .A1(n1061), .A2(n1077), .ZN(n1045) );
XOR2_X1 U909 ( .A(n1237), .B(KEYINPUT34), .Z(n1061) );
XNOR2_X1 U910 ( .A(n1238), .B(n1239), .ZN(G30) );
NOR3_X1 U911 ( .A1(n1212), .A2(n1240), .A3(n1067), .ZN(n1239) );
INV_X1 U912 ( .A(n1208), .ZN(n1067) );
XNOR2_X1 U913 ( .A(n1230), .B(KEYINPUT20), .ZN(n1240) );
NAND3_X1 U914 ( .A1(n1049), .A2(n1235), .A3(n1228), .ZN(n1212) );
AND3_X1 U915 ( .A1(n1241), .A2(n1041), .A3(n1068), .ZN(n1228) );
XNOR2_X1 U916 ( .A(n1217), .B(n1242), .ZN(G3) );
XNOR2_X1 U917 ( .A(KEYINPUT59), .B(n1156), .ZN(n1242) );
AND3_X1 U918 ( .A1(n1054), .A2(n1243), .A3(n1220), .ZN(n1217) );
XNOR2_X1 U919 ( .A(G125), .B(n1207), .ZN(G27) );
NAND4_X1 U920 ( .A1(n1049), .A2(n1241), .A3(n1230), .A4(n1244), .ZN(n1207) );
NOR2_X1 U921 ( .A1(n1235), .A2(n1063), .ZN(n1244) );
NAND2_X1 U922 ( .A1(n1069), .A2(n1245), .ZN(n1241) );
NAND4_X1 U923 ( .A1(G902), .A2(G953), .A3(n1246), .A4(n1110), .ZN(n1245) );
INV_X1 U924 ( .A(G900), .ZN(n1110) );
XOR2_X1 U925 ( .A(G122), .B(n1216), .Z(G24) );
AND4_X1 U926 ( .A1(n1229), .A2(n1247), .A3(n1051), .A4(n1048), .ZN(n1216) );
AND2_X1 U927 ( .A1(n1248), .A2(n1249), .ZN(n1229) );
XNOR2_X1 U928 ( .A(KEYINPUT52), .B(n1250), .ZN(n1248) );
XOR2_X1 U929 ( .A(n1225), .B(n1251), .Z(G21) );
NAND2_X1 U930 ( .A1(KEYINPUT32), .A2(G119), .ZN(n1251) );
NAND4_X1 U931 ( .A1(n1247), .A2(n1054), .A3(n1049), .A4(n1235), .ZN(n1225) );
XNOR2_X1 U932 ( .A(G116), .B(n1224), .ZN(G18) );
NAND3_X1 U933 ( .A1(n1247), .A2(n1208), .A3(n1220), .ZN(n1224) );
NOR2_X1 U934 ( .A1(n1084), .A2(n1252), .ZN(n1208) );
AND2_X1 U935 ( .A1(n1253), .A2(n1042), .ZN(n1247) );
XNOR2_X1 U936 ( .A(G113), .B(n1254), .ZN(G15) );
NAND4_X1 U937 ( .A1(n1255), .A2(n1220), .A3(n1230), .A4(n1221), .ZN(n1254) );
NOR2_X1 U938 ( .A1(n1049), .A2(n1048), .ZN(n1220) );
INV_X1 U939 ( .A(n1063), .ZN(n1255) );
NAND3_X1 U940 ( .A1(n1042), .A2(n1041), .A3(n1223), .ZN(n1063) );
NOR2_X1 U941 ( .A1(n1249), .A2(n1250), .ZN(n1223) );
INV_X1 U942 ( .A(n1084), .ZN(n1250) );
XNOR2_X1 U943 ( .A(G110), .B(n1213), .ZN(G12) );
NAND3_X1 U944 ( .A1(n1222), .A2(n1049), .A3(n1054), .ZN(n1213) );
NOR2_X1 U945 ( .A1(n1249), .A2(n1084), .ZN(n1054) );
XNOR2_X1 U946 ( .A(n1256), .B(G475), .ZN(n1084) );
OR2_X1 U947 ( .A1(n1148), .A2(G902), .ZN(n1256) );
XNOR2_X1 U948 ( .A(n1257), .B(n1258), .ZN(n1148) );
XOR2_X1 U949 ( .A(n1259), .B(n1260), .Z(n1258) );
XNOR2_X1 U950 ( .A(G113), .B(n1261), .ZN(n1260) );
NOR2_X1 U951 ( .A1(KEYINPUT47), .A2(n1262), .ZN(n1261) );
XOR2_X1 U952 ( .A(n1263), .B(n1264), .Z(n1262) );
AND3_X1 U953 ( .A1(G214), .A2(n1034), .A3(n1265), .ZN(n1264) );
XNOR2_X1 U954 ( .A(G131), .B(G143), .ZN(n1263) );
NAND2_X1 U955 ( .A1(KEYINPUT11), .A2(n1153), .ZN(n1259) );
XOR2_X1 U956 ( .A(n1113), .B(n1266), .Z(n1257) );
XOR2_X1 U957 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U958 ( .A(G125), .B(G140), .ZN(n1113) );
INV_X1 U959 ( .A(n1252), .ZN(n1249) );
NOR2_X1 U960 ( .A1(n1076), .A2(n1092), .ZN(n1252) );
AND2_X1 U961 ( .A1(n1269), .A2(n1093), .ZN(n1092) );
NOR2_X1 U962 ( .A1(n1093), .A2(n1269), .ZN(n1076) );
AND2_X1 U963 ( .A1(n1144), .A2(n1270), .ZN(n1269) );
NAND2_X1 U964 ( .A1(n1271), .A2(n1272), .ZN(n1144) );
NAND4_X1 U965 ( .A1(G234), .A2(G217), .A3(n1273), .A4(n1034), .ZN(n1272) );
NAND2_X1 U966 ( .A1(n1274), .A2(n1275), .ZN(n1271) );
NAND3_X1 U967 ( .A1(G217), .A2(n1034), .A3(G234), .ZN(n1275) );
XNOR2_X1 U968 ( .A(n1273), .B(KEYINPUT50), .ZN(n1274) );
XNOR2_X1 U969 ( .A(n1276), .B(n1277), .ZN(n1273) );
XOR2_X1 U970 ( .A(n1278), .B(n1279), .Z(n1277) );
XOR2_X1 U971 ( .A(G134), .B(G116), .Z(n1279) );
XOR2_X1 U972 ( .A(KEYINPUT63), .B(G143), .Z(n1278) );
XOR2_X1 U973 ( .A(n1280), .B(n1268), .Z(n1276) );
XNOR2_X1 U974 ( .A(n1281), .B(n1023), .ZN(n1280) );
NAND2_X1 U975 ( .A1(KEYINPUT36), .A2(n1238), .ZN(n1281) );
INV_X1 U976 ( .A(G478), .ZN(n1093) );
INV_X1 U977 ( .A(n1051), .ZN(n1049) );
XOR2_X1 U978 ( .A(n1101), .B(n1094), .Z(n1051) );
NAND2_X1 U979 ( .A1(G217), .A2(n1282), .ZN(n1094) );
NOR2_X1 U980 ( .A1(n1139), .A2(G902), .ZN(n1101) );
XOR2_X1 U981 ( .A(n1283), .B(n1284), .Z(n1139) );
XOR2_X1 U982 ( .A(n1285), .B(n1286), .Z(n1284) );
XNOR2_X1 U983 ( .A(n1238), .B(G119), .ZN(n1286) );
INV_X1 U984 ( .A(G128), .ZN(n1238) );
XOR2_X1 U985 ( .A(KEYINPUT45), .B(G137), .Z(n1285) );
XOR2_X1 U986 ( .A(n1287), .B(n1288), .Z(n1283) );
AND3_X1 U987 ( .A1(G221), .A2(n1034), .A3(G234), .ZN(n1288) );
XOR2_X1 U988 ( .A(n1289), .B(G110), .Z(n1287) );
NAND2_X1 U989 ( .A1(KEYINPUT58), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U990 ( .A(n1291), .B(n1267), .ZN(n1290) );
XOR2_X1 U991 ( .A(G146), .B(KEYINPUT12), .Z(n1267) );
NAND4_X1 U992 ( .A1(KEYINPUT62), .A2(n1292), .A3(n1293), .A4(n1294), .ZN(n1291) );
OR3_X1 U993 ( .A1(n1295), .A2(KEYINPUT25), .A3(G140), .ZN(n1294) );
NAND2_X1 U994 ( .A1(G140), .A2(n1295), .ZN(n1293) );
NAND2_X1 U995 ( .A1(KEYINPUT39), .A2(n1296), .ZN(n1295) );
NAND2_X1 U996 ( .A1(KEYINPUT25), .A2(G125), .ZN(n1292) );
AND2_X1 U997 ( .A1(n1243), .A2(n1048), .ZN(n1222) );
INV_X1 U998 ( .A(n1235), .ZN(n1048) );
NAND3_X1 U999 ( .A1(n1297), .A2(n1298), .A3(n1299), .ZN(n1235) );
INV_X1 U1000 ( .A(n1075), .ZN(n1299) );
NOR2_X1 U1001 ( .A1(n1081), .A2(G472), .ZN(n1075) );
OR2_X1 U1002 ( .A1(G472), .A2(KEYINPUT2), .ZN(n1298) );
NAND3_X1 U1003 ( .A1(G472), .A2(n1081), .A3(KEYINPUT2), .ZN(n1297) );
NAND2_X1 U1004 ( .A1(n1300), .A2(n1270), .ZN(n1081) );
XOR2_X1 U1005 ( .A(n1301), .B(n1302), .Z(n1300) );
XNOR2_X1 U1006 ( .A(G101), .B(n1303), .ZN(n1302) );
XNOR2_X1 U1007 ( .A(KEYINPUT7), .B(KEYINPUT33), .ZN(n1303) );
XNOR2_X1 U1008 ( .A(n1162), .B(n1164), .ZN(n1301) );
AND3_X1 U1009 ( .A1(n1265), .A2(n1034), .A3(G210), .ZN(n1164) );
XNOR2_X1 U1010 ( .A(n1304), .B(n1305), .ZN(n1162) );
XOR2_X1 U1011 ( .A(KEYINPUT60), .B(KEYINPUT18), .Z(n1305) );
XOR2_X1 U1012 ( .A(n1112), .B(n1133), .Z(n1304) );
XNOR2_X1 U1013 ( .A(n1191), .B(n1181), .ZN(n1112) );
INV_X1 U1014 ( .A(n1178), .ZN(n1181) );
AND2_X1 U1015 ( .A1(n1253), .A2(n1068), .ZN(n1243) );
INV_X1 U1016 ( .A(n1042), .ZN(n1068) );
XNOR2_X1 U1017 ( .A(n1080), .B(n1306), .ZN(n1042) );
XOR2_X1 U1018 ( .A(KEYINPUT17), .B(G469), .Z(n1306) );
NAND2_X1 U1019 ( .A1(n1307), .A2(n1270), .ZN(n1080) );
XOR2_X1 U1020 ( .A(n1308), .B(n1309), .Z(n1307) );
XNOR2_X1 U1021 ( .A(n1184), .B(n1178), .ZN(n1309) );
XOR2_X1 U1022 ( .A(G131), .B(n1310), .Z(n1178) );
XOR2_X1 U1023 ( .A(G137), .B(G134), .Z(n1310) );
NAND2_X1 U1024 ( .A1(G227), .A2(n1034), .ZN(n1184) );
XOR2_X1 U1025 ( .A(n1311), .B(n1312), .Z(n1308) );
NOR2_X1 U1026 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1027 ( .A(KEYINPUT9), .B(n1315), .Z(n1314) );
NOR2_X1 U1028 ( .A1(n1186), .A2(n1316), .ZN(n1315) );
AND2_X1 U1029 ( .A1(n1186), .A2(n1316), .ZN(n1313) );
XOR2_X1 U1030 ( .A(G110), .B(KEYINPUT4), .Z(n1316) );
INV_X1 U1031 ( .A(G140), .ZN(n1186) );
NAND2_X1 U1032 ( .A1(KEYINPUT37), .A2(n1179), .ZN(n1311) );
XNOR2_X1 U1033 ( .A(n1317), .B(n1318), .ZN(n1179) );
XNOR2_X1 U1034 ( .A(n1023), .B(G104), .ZN(n1318) );
INV_X1 U1035 ( .A(G107), .ZN(n1023) );
XNOR2_X1 U1036 ( .A(n1191), .B(n1156), .ZN(n1317) );
AND3_X1 U1037 ( .A1(n1041), .A2(n1221), .A3(n1230), .ZN(n1253) );
INV_X1 U1038 ( .A(n1059), .ZN(n1230) );
NAND2_X1 U1039 ( .A1(n1237), .A2(n1077), .ZN(n1059) );
NAND2_X1 U1040 ( .A1(G214), .A2(n1319), .ZN(n1077) );
XNOR2_X1 U1041 ( .A(n1320), .B(n1197), .ZN(n1237) );
NAND2_X1 U1042 ( .A1(G210), .A2(n1319), .ZN(n1197) );
NAND2_X1 U1043 ( .A1(n1265), .A2(n1270), .ZN(n1319) );
INV_X1 U1044 ( .A(G237), .ZN(n1265) );
NAND2_X1 U1045 ( .A1(n1321), .A2(n1086), .ZN(n1320) );
NAND3_X1 U1046 ( .A1(n1322), .A2(n1270), .A3(n1323), .ZN(n1086) );
XOR2_X1 U1047 ( .A(n1324), .B(KEYINPUT1), .Z(n1323) );
OR2_X1 U1048 ( .A1(n1325), .A2(n1196), .ZN(n1324) );
NAND2_X1 U1049 ( .A1(n1196), .A2(n1325), .ZN(n1322) );
XNOR2_X1 U1050 ( .A(n1326), .B(n1192), .ZN(n1325) );
XNOR2_X1 U1051 ( .A(n1296), .B(n1327), .ZN(n1192) );
NOR2_X1 U1052 ( .A1(G953), .A2(n1123), .ZN(n1327) );
INV_X1 U1053 ( .A(G224), .ZN(n1123) );
INV_X1 U1054 ( .A(G125), .ZN(n1296) );
NAND2_X1 U1055 ( .A1(KEYINPUT57), .A2(n1191), .ZN(n1326) );
XNOR2_X1 U1056 ( .A(G128), .B(n1328), .ZN(n1191) );
XOR2_X1 U1057 ( .A(G146), .B(G143), .Z(n1328) );
XNOR2_X1 U1058 ( .A(n1329), .B(n1131), .ZN(n1196) );
XOR2_X1 U1059 ( .A(G110), .B(n1268), .Z(n1131) );
XOR2_X1 U1060 ( .A(G122), .B(KEYINPUT31), .Z(n1268) );
XNOR2_X1 U1061 ( .A(n1134), .B(n1330), .ZN(n1329) );
NOR2_X1 U1062 ( .A1(KEYINPUT10), .A2(n1133), .ZN(n1330) );
XOR2_X1 U1063 ( .A(G113), .B(n1331), .Z(n1133) );
XOR2_X1 U1064 ( .A(G119), .B(G116), .Z(n1331) );
XOR2_X1 U1065 ( .A(n1332), .B(n1156), .Z(n1134) );
INV_X1 U1066 ( .A(G101), .ZN(n1156) );
NAND4_X1 U1067 ( .A1(KEYINPUT28), .A2(n1333), .A3(n1334), .A4(n1335), .ZN(n1332) );
NAND3_X1 U1068 ( .A1(KEYINPUT27), .A2(n1336), .A3(n1337), .ZN(n1335) );
OR2_X1 U1069 ( .A1(n1337), .A2(n1336), .ZN(n1334) );
AND2_X1 U1070 ( .A1(KEYINPUT6), .A2(n1153), .ZN(n1336) );
XOR2_X1 U1071 ( .A(G107), .B(KEYINPUT51), .Z(n1337) );
OR2_X1 U1072 ( .A1(n1153), .A2(KEYINPUT27), .ZN(n1333) );
INV_X1 U1073 ( .A(G104), .ZN(n1153) );
XOR2_X1 U1074 ( .A(KEYINPUT35), .B(KEYINPUT24), .Z(n1321) );
NAND2_X1 U1075 ( .A1(n1069), .A2(n1338), .ZN(n1221) );
NAND3_X1 U1076 ( .A1(n1129), .A2(n1246), .A3(G902), .ZN(n1338) );
NOR2_X1 U1077 ( .A1(n1034), .A2(G898), .ZN(n1129) );
NAND3_X1 U1078 ( .A1(n1246), .A2(n1034), .A3(G952), .ZN(n1069) );
INV_X1 U1079 ( .A(G953), .ZN(n1034) );
NAND2_X1 U1080 ( .A1(G237), .A2(G234), .ZN(n1246) );
NAND2_X1 U1081 ( .A1(G221), .A2(n1282), .ZN(n1041) );
NAND2_X1 U1082 ( .A1(G234), .A2(n1270), .ZN(n1282) );
INV_X1 U1083 ( .A(G902), .ZN(n1270) );
endmodule


