//Key = 1100101010011111010110001010111011110111100111011011110000000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352;

XNOR2_X1 U746 ( .A(G107), .B(n1029), .ZN(G9) );
NOR2_X1 U747 ( .A1(n1030), .A2(KEYINPUT61), .ZN(n1029) );
NOR2_X1 U748 ( .A1(n1031), .A2(n1032), .ZN(G75) );
XOR2_X1 U749 ( .A(KEYINPUT46), .B(n1033), .Z(n1032) );
NOR3_X1 U750 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NOR2_X1 U751 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U752 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR3_X1 U753 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1040) );
NOR3_X1 U754 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NOR2_X1 U755 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U756 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1045) );
NOR2_X1 U759 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U760 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NOR2_X1 U761 ( .A1(n1059), .A2(n1060), .ZN(n1042) );
NOR3_X1 U762 ( .A1(n1054), .A2(n1061), .A3(n1048), .ZN(n1060) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
INV_X1 U764 ( .A(n1064), .ZN(n1041) );
NOR4_X1 U765 ( .A1(n1065), .A2(n1048), .A3(n1044), .A4(n1054), .ZN(n1039) );
INV_X1 U766 ( .A(n1066), .ZN(n1054) );
INV_X1 U767 ( .A(n1067), .ZN(n1048) );
NOR2_X1 U768 ( .A1(n1068), .A2(n1069), .ZN(n1065) );
NOR2_X1 U769 ( .A1(G952), .A2(n1036), .ZN(n1031) );
NAND2_X1 U770 ( .A1(n1070), .A2(n1071), .ZN(n1036) );
NAND4_X1 U771 ( .A1(n1072), .A2(n1059), .A3(n1073), .A4(n1052), .ZN(n1071) );
XOR2_X1 U772 ( .A(KEYINPUT16), .B(n1074), .Z(n1073) );
NOR4_X1 U773 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
INV_X1 U774 ( .A(n1079), .ZN(n1077) );
NOR2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1076) );
XNOR2_X1 U776 ( .A(G478), .B(KEYINPUT55), .ZN(n1081) );
NAND3_X1 U777 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1075) );
NAND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
XNOR2_X1 U779 ( .A(n1087), .B(n1088), .ZN(n1072) );
XOR2_X1 U780 ( .A(n1089), .B(n1090), .Z(G72) );
XOR2_X1 U781 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U783 ( .A1(G953), .A2(n1095), .ZN(n1094) );
XOR2_X1 U784 ( .A(n1096), .B(n1097), .Z(n1093) );
XNOR2_X1 U785 ( .A(n1098), .B(n1099), .ZN(n1097) );
NAND2_X1 U786 ( .A1(KEYINPUT30), .A2(n1100), .ZN(n1098) );
XOR2_X1 U787 ( .A(n1101), .B(n1102), .Z(n1096) );
XNOR2_X1 U788 ( .A(n1103), .B(G125), .ZN(n1102) );
NOR2_X1 U789 ( .A1(KEYINPUT21), .A2(n1104), .ZN(n1101) );
NAND2_X1 U790 ( .A1(G953), .A2(n1105), .ZN(n1091) );
NAND2_X1 U791 ( .A1(n1106), .A2(G227), .ZN(n1105) );
XNOR2_X1 U792 ( .A(G900), .B(KEYINPUT32), .ZN(n1106) );
NOR2_X1 U793 ( .A1(n1107), .A2(G953), .ZN(n1089) );
NAND3_X1 U794 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(G69) );
OR2_X1 U795 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U796 ( .A1(n1113), .A2(n1114), .ZN(n1109) );
NAND2_X1 U797 ( .A1(KEYINPUT29), .A2(n1112), .ZN(n1114) );
INV_X1 U798 ( .A(n1115), .ZN(n1113) );
NAND2_X1 U799 ( .A1(n1116), .A2(n1115), .ZN(n1108) );
NAND2_X1 U800 ( .A1(G953), .A2(n1117), .ZN(n1115) );
NAND2_X1 U801 ( .A1(G898), .A2(G224), .ZN(n1117) );
NAND2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
OR2_X1 U803 ( .A1(n1111), .A2(KEYINPUT29), .ZN(n1119) );
NAND3_X1 U804 ( .A1(n1112), .A2(n1111), .A3(KEYINPUT29), .ZN(n1118) );
NAND2_X1 U805 ( .A1(n1070), .A2(n1120), .ZN(n1111) );
NAND2_X1 U806 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
AND2_X1 U807 ( .A1(n1123), .A2(n1124), .ZN(n1112) );
NAND2_X1 U808 ( .A1(G953), .A2(n1125), .ZN(n1124) );
XNOR2_X1 U809 ( .A(KEYINPUT14), .B(n1126), .ZN(n1125) );
XNOR2_X1 U810 ( .A(n1127), .B(n1128), .ZN(n1123) );
XNOR2_X1 U811 ( .A(n1129), .B(n1130), .ZN(n1128) );
NOR2_X1 U812 ( .A1(KEYINPUT10), .A2(n1131), .ZN(n1130) );
NAND2_X1 U813 ( .A1(KEYINPUT39), .A2(n1132), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1133), .A2(n1134), .ZN(G66) );
NOR3_X1 U815 ( .A1(n1085), .A2(n1135), .A3(n1136), .ZN(n1134) );
NOR3_X1 U816 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1136) );
INV_X1 U817 ( .A(n1140), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1141), .A2(n1140), .ZN(n1135) );
NOR2_X1 U819 ( .A1(n1142), .A2(n1138), .ZN(n1141) );
XOR2_X1 U820 ( .A(G217), .B(KEYINPUT12), .Z(n1138) );
NOR2_X1 U821 ( .A1(n1133), .A2(n1143), .ZN(G63) );
XNOR2_X1 U822 ( .A(n1144), .B(n1145), .ZN(n1143) );
NOR2_X1 U823 ( .A1(n1146), .A2(n1139), .ZN(n1145) );
NOR2_X1 U824 ( .A1(n1133), .A2(n1147), .ZN(G60) );
XNOR2_X1 U825 ( .A(n1148), .B(n1149), .ZN(n1147) );
AND2_X1 U826 ( .A1(G475), .A2(n1150), .ZN(n1149) );
XNOR2_X1 U827 ( .A(n1122), .B(n1151), .ZN(G6) );
NOR2_X1 U828 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U829 ( .A(KEYINPUT4), .B(KEYINPUT26), .Z(n1153) );
INV_X1 U830 ( .A(G104), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1133), .A2(n1154), .ZN(G57) );
XOR2_X1 U832 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U833 ( .A(n1157), .B(n1158), .ZN(n1156) );
AND2_X1 U834 ( .A1(G472), .A2(n1150), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1159), .B(KEYINPUT15), .Z(n1155) );
NAND2_X1 U836 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
NAND2_X1 U837 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U838 ( .A(KEYINPUT37), .B(n1164), .Z(n1160) );
NOR2_X1 U839 ( .A1(n1162), .A2(n1163), .ZN(n1164) );
XOR2_X1 U840 ( .A(n1165), .B(n1166), .Z(n1162) );
NOR2_X1 U841 ( .A1(n1133), .A2(n1167), .ZN(G54) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U844 ( .A(n1172), .B(n1173), .Z(n1170) );
NAND2_X1 U845 ( .A1(KEYINPUT43), .A2(n1100), .ZN(n1172) );
XOR2_X1 U846 ( .A(n1174), .B(n1175), .Z(n1168) );
NOR2_X1 U847 ( .A1(KEYINPUT25), .A2(n1176), .ZN(n1175) );
XOR2_X1 U848 ( .A(n1177), .B(KEYINPUT2), .Z(n1174) );
NAND2_X1 U849 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U850 ( .A1(n1180), .A2(G469), .A3(n1150), .ZN(n1179) );
INV_X1 U851 ( .A(KEYINPUT52), .ZN(n1180) );
NAND2_X1 U852 ( .A1(KEYINPUT6), .A2(n1181), .ZN(n1178) );
NAND2_X1 U853 ( .A1(n1150), .A2(G469), .ZN(n1181) );
NOR2_X1 U854 ( .A1(n1133), .A2(n1182), .ZN(G51) );
XOR2_X1 U855 ( .A(n1183), .B(n1184), .Z(n1182) );
XOR2_X1 U856 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U857 ( .A1(KEYINPUT63), .A2(n1187), .ZN(n1185) );
XOR2_X1 U858 ( .A(n1188), .B(n1189), .Z(n1183) );
NOR2_X1 U859 ( .A1(n1088), .A2(n1139), .ZN(n1189) );
INV_X1 U860 ( .A(n1150), .ZN(n1139) );
NOR2_X1 U861 ( .A1(n1190), .A2(n1142), .ZN(n1150) );
INV_X1 U862 ( .A(n1034), .ZN(n1142) );
NAND3_X1 U863 ( .A1(n1107), .A2(n1121), .A3(n1191), .ZN(n1034) );
XOR2_X1 U864 ( .A(n1122), .B(KEYINPUT42), .Z(n1191) );
NAND3_X1 U865 ( .A1(n1192), .A2(n1067), .A3(n1069), .ZN(n1122) );
AND4_X1 U866 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1121) );
NOR4_X1 U867 ( .A1(n1197), .A2(n1198), .A3(n1030), .A4(n1199), .ZN(n1196) );
AND3_X1 U868 ( .A1(n1068), .A2(n1067), .A3(n1192), .ZN(n1030) );
NAND2_X1 U869 ( .A1(n1050), .A2(n1200), .ZN(n1195) );
XOR2_X1 U870 ( .A(KEYINPUT18), .B(n1201), .Z(n1200) );
AND4_X1 U871 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1107) );
NOR4_X1 U872 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205) );
AND2_X1 U873 ( .A1(n1210), .A2(n1211), .ZN(n1204) );
NAND4_X1 U874 ( .A1(n1069), .A2(n1066), .A3(n1212), .A4(n1213), .ZN(n1202) );
XOR2_X1 U875 ( .A(n1214), .B(KEYINPUT27), .Z(n1188) );
NAND2_X1 U876 ( .A1(KEYINPUT1), .A2(n1215), .ZN(n1214) );
NOR2_X1 U877 ( .A1(n1070), .A2(G952), .ZN(n1133) );
XOR2_X1 U878 ( .A(n1216), .B(G146), .Z(G48) );
NAND2_X1 U879 ( .A1(KEYINPUT40), .A2(n1210), .ZN(n1216) );
NAND2_X1 U880 ( .A1(n1069), .A2(n1217), .ZN(n1210) );
XNOR2_X1 U881 ( .A(G143), .B(n1203), .ZN(G45) );
NAND4_X1 U882 ( .A1(n1218), .A2(n1050), .A3(n1219), .A4(n1220), .ZN(n1203) );
XNOR2_X1 U883 ( .A(G140), .B(n1221), .ZN(G42) );
NAND4_X1 U884 ( .A1(n1222), .A2(n1069), .A3(n1212), .A4(n1213), .ZN(n1221) );
XNOR2_X1 U885 ( .A(n1066), .B(KEYINPUT35), .ZN(n1222) );
XNOR2_X1 U886 ( .A(G137), .B(n1223), .ZN(G39) );
NAND2_X1 U887 ( .A1(KEYINPUT28), .A2(n1209), .ZN(n1223) );
AND4_X1 U888 ( .A1(n1064), .A2(n1066), .A3(n1212), .A4(n1224), .ZN(n1209) );
XOR2_X1 U889 ( .A(G134), .B(n1208), .Z(G36) );
AND3_X1 U890 ( .A1(n1218), .A2(n1068), .A3(n1066), .ZN(n1208) );
XOR2_X1 U891 ( .A(G131), .B(n1207), .Z(G33) );
AND3_X1 U892 ( .A1(n1066), .A2(n1218), .A3(n1069), .ZN(n1207) );
AND3_X1 U893 ( .A1(n1225), .A2(n1226), .A3(n1056), .ZN(n1218) );
NOR2_X1 U894 ( .A1(n1051), .A2(n1227), .ZN(n1066) );
INV_X1 U895 ( .A(n1052), .ZN(n1227) );
XNOR2_X1 U896 ( .A(G128), .B(n1228), .ZN(G30) );
NAND2_X1 U897 ( .A1(KEYINPUT11), .A2(n1206), .ZN(n1228) );
AND2_X1 U898 ( .A1(n1217), .A2(n1068), .ZN(n1206) );
AND3_X1 U899 ( .A1(n1050), .A2(n1224), .A3(n1212), .ZN(n1217) );
AND3_X1 U900 ( .A1(n1226), .A2(n1229), .A3(n1225), .ZN(n1212) );
XNOR2_X1 U901 ( .A(n1194), .B(n1230), .ZN(G3) );
NOR2_X1 U902 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
XOR2_X1 U903 ( .A(KEYINPUT34), .B(KEYINPUT24), .Z(n1232) );
NAND3_X1 U904 ( .A1(n1056), .A2(n1192), .A3(n1064), .ZN(n1194) );
XOR2_X1 U905 ( .A(n1211), .B(n1233), .Z(G27) );
XOR2_X1 U906 ( .A(KEYINPUT44), .B(G125), .Z(n1233) );
NAND4_X1 U907 ( .A1(n1059), .A2(n1050), .A3(n1069), .A4(n1234), .ZN(n1211) );
AND3_X1 U908 ( .A1(n1213), .A2(n1229), .A3(n1226), .ZN(n1234) );
NAND2_X1 U909 ( .A1(n1038), .A2(n1235), .ZN(n1226) );
NAND4_X1 U910 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1095), .ZN(n1235) );
INV_X1 U911 ( .A(G900), .ZN(n1095) );
XNOR2_X1 U912 ( .A(G122), .B(n1237), .ZN(G24) );
NOR2_X1 U913 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NOR2_X1 U914 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NAND4_X1 U915 ( .A1(n1050), .A2(n1219), .A3(n1067), .A4(n1242), .ZN(n1241) );
NOR3_X1 U916 ( .A1(n1243), .A2(n1244), .A3(n1059), .ZN(n1242) );
INV_X1 U917 ( .A(KEYINPUT22), .ZN(n1240) );
NOR2_X1 U918 ( .A1(KEYINPUT22), .A2(n1193), .ZN(n1238) );
NAND4_X1 U919 ( .A1(n1245), .A2(n1067), .A3(n1219), .A4(n1220), .ZN(n1193) );
NOR2_X1 U920 ( .A1(n1229), .A2(n1058), .ZN(n1067) );
INV_X1 U921 ( .A(n1213), .ZN(n1058) );
XNOR2_X1 U922 ( .A(G119), .B(n1246), .ZN(G21) );
NAND2_X1 U923 ( .A1(n1201), .A2(n1050), .ZN(n1246) );
AND3_X1 U924 ( .A1(n1064), .A2(n1059), .A3(n1247), .ZN(n1201) );
NOR3_X1 U925 ( .A1(n1084), .A2(n1057), .A3(n1243), .ZN(n1247) );
INV_X1 U926 ( .A(n1248), .ZN(n1243) );
NAND2_X1 U927 ( .A1(n1249), .A2(n1250), .ZN(G18) );
NAND2_X1 U928 ( .A1(n1198), .A2(n1251), .ZN(n1250) );
XOR2_X1 U929 ( .A(KEYINPUT19), .B(n1252), .Z(n1249) );
NOR2_X1 U930 ( .A1(n1198), .A2(n1251), .ZN(n1252) );
AND3_X1 U931 ( .A1(n1056), .A2(n1068), .A3(n1245), .ZN(n1198) );
NOR2_X1 U932 ( .A1(n1219), .A2(n1244), .ZN(n1068) );
INV_X1 U933 ( .A(n1220), .ZN(n1244) );
XOR2_X1 U934 ( .A(G113), .B(n1199), .Z(G15) );
AND3_X1 U935 ( .A1(n1069), .A2(n1056), .A3(n1245), .ZN(n1199) );
AND3_X1 U936 ( .A1(n1050), .A2(n1248), .A3(n1059), .ZN(n1245) );
INV_X1 U937 ( .A(n1044), .ZN(n1059) );
NAND2_X1 U938 ( .A1(n1062), .A2(n1063), .ZN(n1044) );
NOR2_X1 U939 ( .A1(n1229), .A2(n1084), .ZN(n1056) );
INV_X1 U940 ( .A(n1224), .ZN(n1084) );
NOR2_X1 U941 ( .A1(n1220), .A2(n1082), .ZN(n1069) );
INV_X1 U942 ( .A(n1219), .ZN(n1082) );
XOR2_X1 U943 ( .A(G110), .B(n1197), .Z(G12) );
AND4_X1 U944 ( .A1(n1064), .A2(n1192), .A3(n1213), .A4(n1229), .ZN(n1197) );
INV_X1 U945 ( .A(n1057), .ZN(n1229) );
NOR2_X1 U946 ( .A1(n1253), .A2(n1078), .ZN(n1057) );
NOR2_X1 U947 ( .A1(n1086), .A2(n1085), .ZN(n1078) );
AND2_X1 U948 ( .A1(n1254), .A2(n1086), .ZN(n1253) );
NAND2_X1 U949 ( .A1(G217), .A2(n1255), .ZN(n1086) );
XOR2_X1 U950 ( .A(KEYINPUT62), .B(n1085), .Z(n1254) );
NOR2_X1 U951 ( .A1(n1140), .A2(G902), .ZN(n1085) );
XNOR2_X1 U952 ( .A(n1256), .B(n1257), .ZN(n1140) );
XOR2_X1 U953 ( .A(n1258), .B(n1259), .Z(n1257) );
XOR2_X1 U954 ( .A(G137), .B(G125), .Z(n1259) );
XOR2_X1 U955 ( .A(KEYINPUT50), .B(KEYINPUT41), .Z(n1258) );
XOR2_X1 U956 ( .A(n1260), .B(n1261), .Z(n1256) );
XOR2_X1 U957 ( .A(n1262), .B(n1173), .Z(n1261) );
XNOR2_X1 U958 ( .A(G110), .B(n1103), .ZN(n1173) );
XOR2_X1 U959 ( .A(n1263), .B(G119), .Z(n1260) );
NAND3_X1 U960 ( .A1(n1264), .A2(n1070), .A3(G221), .ZN(n1263) );
XOR2_X1 U961 ( .A(KEYINPUT49), .B(G234), .Z(n1264) );
XOR2_X1 U962 ( .A(n1224), .B(KEYINPUT13), .Z(n1213) );
XNOR2_X1 U963 ( .A(n1265), .B(G472), .ZN(n1224) );
NAND2_X1 U964 ( .A1(n1266), .A2(n1190), .ZN(n1265) );
XOR2_X1 U965 ( .A(n1267), .B(n1268), .Z(n1266) );
XNOR2_X1 U966 ( .A(n1165), .B(n1269), .ZN(n1268) );
INV_X1 U967 ( .A(n1157), .ZN(n1269) );
XOR2_X1 U968 ( .A(n1270), .B(n1231), .Z(n1157) );
INV_X1 U969 ( .A(G101), .ZN(n1231) );
NAND2_X1 U970 ( .A1(n1271), .A2(G210), .ZN(n1270) );
XNOR2_X1 U971 ( .A(n1163), .B(n1272), .ZN(n1267) );
NOR2_X1 U972 ( .A1(KEYINPUT56), .A2(n1166), .ZN(n1272) );
XNOR2_X1 U973 ( .A(n1273), .B(n1274), .ZN(n1163) );
NOR2_X1 U974 ( .A1(KEYINPUT23), .A2(G116), .ZN(n1274) );
XNOR2_X1 U975 ( .A(G113), .B(G119), .ZN(n1273) );
AND3_X1 U976 ( .A1(n1225), .A2(n1248), .A3(n1050), .ZN(n1192) );
AND2_X1 U977 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U978 ( .A1(G214), .A2(n1275), .ZN(n1052) );
XNOR2_X1 U979 ( .A(n1276), .B(n1087), .ZN(n1051) );
NAND3_X1 U980 ( .A1(n1277), .A2(n1278), .A3(n1190), .ZN(n1087) );
NAND2_X1 U981 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
INV_X1 U982 ( .A(n1281), .ZN(n1279) );
NAND2_X1 U983 ( .A1(n1281), .A2(n1282), .ZN(n1277) );
NAND2_X1 U984 ( .A1(n1283), .A2(n1284), .ZN(n1282) );
NAND2_X1 U985 ( .A1(KEYINPUT5), .A2(n1285), .ZN(n1284) );
INV_X1 U986 ( .A(n1187), .ZN(n1285) );
OR2_X1 U987 ( .A1(n1280), .A2(KEYINPUT5), .ZN(n1283) );
NOR2_X1 U988 ( .A1(KEYINPUT59), .A2(n1187), .ZN(n1280) );
NAND2_X1 U989 ( .A1(n1286), .A2(n1287), .ZN(n1187) );
NAND2_X1 U990 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U991 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U992 ( .A1(KEYINPUT20), .A2(n1292), .ZN(n1291) );
INV_X1 U993 ( .A(KEYINPUT31), .ZN(n1290) );
NAND2_X1 U994 ( .A1(n1132), .A2(n1293), .ZN(n1286) );
NAND2_X1 U995 ( .A1(KEYINPUT20), .A2(n1294), .ZN(n1293) );
OR2_X1 U996 ( .A1(n1288), .A2(KEYINPUT31), .ZN(n1294) );
XNOR2_X1 U997 ( .A(n1131), .B(n1295), .ZN(n1288) );
INV_X1 U998 ( .A(n1127), .ZN(n1295) );
XOR2_X1 U999 ( .A(n1296), .B(G113), .Z(n1131) );
NAND2_X1 U1000 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
NAND2_X1 U1001 ( .A1(G119), .A2(n1299), .ZN(n1298) );
XOR2_X1 U1002 ( .A(KEYINPUT48), .B(n1300), .Z(n1297) );
NOR2_X1 U1003 ( .A1(G119), .A2(n1299), .ZN(n1300) );
XNOR2_X1 U1004 ( .A(KEYINPUT45), .B(n1251), .ZN(n1299) );
INV_X1 U1005 ( .A(n1292), .ZN(n1132) );
XOR2_X1 U1006 ( .A(n1301), .B(n1302), .Z(n1292) );
NAND2_X1 U1007 ( .A1(KEYINPUT33), .A2(G110), .ZN(n1301) );
XOR2_X1 U1008 ( .A(n1303), .B(n1215), .Z(n1281) );
XNOR2_X1 U1009 ( .A(G125), .B(KEYINPUT3), .ZN(n1215) );
XNOR2_X1 U1010 ( .A(n1186), .B(KEYINPUT36), .ZN(n1303) );
XNOR2_X1 U1011 ( .A(n1165), .B(n1304), .ZN(n1186) );
AND2_X1 U1012 ( .A1(n1070), .A2(G224), .ZN(n1304) );
XOR2_X1 U1013 ( .A(n1305), .B(n1306), .Z(n1165) );
XNOR2_X1 U1014 ( .A(G146), .B(n1307), .ZN(n1306) );
NAND2_X1 U1015 ( .A1(KEYINPUT47), .A2(n1308), .ZN(n1305) );
NAND2_X1 U1016 ( .A1(KEYINPUT17), .A2(n1088), .ZN(n1276) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1275), .ZN(n1088) );
NAND2_X1 U1018 ( .A1(n1309), .A2(n1190), .ZN(n1275) );
INV_X1 U1019 ( .A(G237), .ZN(n1309) );
NAND2_X1 U1020 ( .A1(n1310), .A2(n1038), .ZN(n1248) );
NAND3_X1 U1021 ( .A1(n1236), .A2(n1070), .A3(G952), .ZN(n1038) );
XOR2_X1 U1022 ( .A(n1311), .B(KEYINPUT60), .Z(n1310) );
NAND4_X1 U1023 ( .A1(G953), .A2(G902), .A3(n1236), .A4(n1126), .ZN(n1311) );
INV_X1 U1024 ( .A(G898), .ZN(n1126) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1236) );
NOR2_X1 U1026 ( .A1(n1062), .A2(n1312), .ZN(n1225) );
INV_X1 U1027 ( .A(n1063), .ZN(n1312) );
NAND2_X1 U1028 ( .A1(G221), .A2(n1255), .ZN(n1063) );
NAND2_X1 U1029 ( .A1(G234), .A2(n1190), .ZN(n1255) );
XOR2_X1 U1030 ( .A(n1313), .B(G469), .Z(n1062) );
NAND2_X1 U1031 ( .A1(n1314), .A2(n1190), .ZN(n1313) );
XOR2_X1 U1032 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1033 ( .A(n1317), .B(n1100), .ZN(n1316) );
XOR2_X1 U1034 ( .A(n1318), .B(n1262), .Z(n1100) );
XNOR2_X1 U1035 ( .A(n1308), .B(G146), .ZN(n1262) );
INV_X1 U1036 ( .A(G128), .ZN(n1308) );
NAND2_X1 U1037 ( .A1(KEYINPUT38), .A2(n1307), .ZN(n1318) );
XNOR2_X1 U1038 ( .A(n1171), .B(n1319), .ZN(n1317) );
NOR2_X1 U1039 ( .A1(G110), .A2(KEYINPUT57), .ZN(n1319) );
XOR2_X1 U1040 ( .A(n1127), .B(n1166), .Z(n1171) );
XNOR2_X1 U1041 ( .A(n1104), .B(n1099), .ZN(n1166) );
XOR2_X1 U1042 ( .A(G134), .B(G137), .Z(n1099) );
XOR2_X1 U1043 ( .A(G101), .B(n1320), .Z(n1127) );
XNOR2_X1 U1044 ( .A(n1321), .B(G104), .ZN(n1320) );
INV_X1 U1045 ( .A(G107), .ZN(n1321) );
XOR2_X1 U1046 ( .A(n1176), .B(n1322), .Z(n1315) );
XNOR2_X1 U1047 ( .A(KEYINPUT8), .B(n1103), .ZN(n1322) );
NAND2_X1 U1048 ( .A1(G227), .A2(n1070), .ZN(n1176) );
NOR2_X1 U1049 ( .A1(n1220), .A2(n1219), .ZN(n1064) );
XNOR2_X1 U1050 ( .A(n1323), .B(G475), .ZN(n1219) );
NAND2_X1 U1051 ( .A1(n1148), .A2(n1190), .ZN(n1323) );
XNOR2_X1 U1052 ( .A(n1324), .B(n1325), .ZN(n1148) );
XOR2_X1 U1053 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1054 ( .A(n1328), .B(n1329), .Z(n1327) );
NOR3_X1 U1055 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1329) );
NOR2_X1 U1056 ( .A1(n1333), .A2(n1103), .ZN(n1332) );
INV_X1 U1057 ( .A(G140), .ZN(n1103) );
NOR3_X1 U1058 ( .A1(G140), .A2(KEYINPUT58), .A3(n1334), .ZN(n1331) );
INV_X1 U1059 ( .A(n1333), .ZN(n1334) );
NOR2_X1 U1060 ( .A1(G125), .A2(KEYINPUT9), .ZN(n1333) );
AND2_X1 U1061 ( .A1(G125), .A2(KEYINPUT58), .ZN(n1330) );
NAND2_X1 U1062 ( .A1(n1335), .A2(KEYINPUT0), .ZN(n1328) );
XNOR2_X1 U1063 ( .A(n1336), .B(n1104), .ZN(n1335) );
XNOR2_X1 U1064 ( .A(G131), .B(KEYINPUT53), .ZN(n1104) );
XNOR2_X1 U1065 ( .A(n1337), .B(n1307), .ZN(n1336) );
NAND2_X1 U1066 ( .A1(n1271), .A2(G214), .ZN(n1337) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1271) );
NAND2_X1 U1068 ( .A1(KEYINPUT51), .A2(G113), .ZN(n1326) );
XOR2_X1 U1069 ( .A(n1338), .B(n1339), .Z(n1324) );
XOR2_X1 U1070 ( .A(KEYINPUT41), .B(G146), .Z(n1339) );
XNOR2_X1 U1071 ( .A(G104), .B(G122), .ZN(n1338) );
NAND2_X1 U1072 ( .A1(n1340), .A2(n1079), .ZN(n1220) );
NAND2_X1 U1073 ( .A1(n1080), .A2(n1146), .ZN(n1079) );
OR2_X1 U1074 ( .A1(n1146), .A2(n1080), .ZN(n1340) );
AND2_X1 U1075 ( .A1(n1190), .A2(n1144), .ZN(n1080) );
NAND2_X1 U1076 ( .A1(n1341), .A2(n1342), .ZN(n1144) );
NAND2_X1 U1077 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
XOR2_X1 U1078 ( .A(n1345), .B(KEYINPUT54), .Z(n1341) );
OR2_X1 U1079 ( .A1(n1344), .A2(n1343), .ZN(n1345) );
AND3_X1 U1080 ( .A1(G234), .A2(n1070), .A3(G217), .ZN(n1343) );
INV_X1 U1081 ( .A(G953), .ZN(n1070) );
XNOR2_X1 U1082 ( .A(n1346), .B(n1347), .ZN(n1344) );
XNOR2_X1 U1083 ( .A(G107), .B(n1348), .ZN(n1347) );
NAND2_X1 U1084 ( .A1(n1349), .A2(n1350), .ZN(n1348) );
NAND2_X1 U1085 ( .A1(G116), .A2(n1302), .ZN(n1350) );
INV_X1 U1086 ( .A(G122), .ZN(n1302) );
XOR2_X1 U1087 ( .A(n1351), .B(KEYINPUT7), .Z(n1349) );
NAND2_X1 U1088 ( .A1(G122), .A2(n1251), .ZN(n1351) );
INV_X1 U1089 ( .A(G116), .ZN(n1251) );
XNOR2_X1 U1090 ( .A(G128), .B(n1352), .ZN(n1346) );
XNOR2_X1 U1091 ( .A(n1307), .B(G134), .ZN(n1352) );
INV_X1 U1092 ( .A(G143), .ZN(n1307) );
INV_X1 U1093 ( .A(G902), .ZN(n1190) );
INV_X1 U1094 ( .A(G478), .ZN(n1146) );
endmodule


