//Key = 1000110011101010000101000000101010100110010110000100011010110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326;

XOR2_X1 U727 ( .A(G107), .B(n1002), .Z(G9) );
NOR2_X1 U728 ( .A1(n1003), .A2(n1004), .ZN(G75) );
NOR4_X1 U729 ( .A1(G953), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n1004) );
NOR2_X1 U730 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR2_X1 U731 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR3_X1 U732 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
NOR2_X1 U733 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U734 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR2_X1 U735 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NOR2_X1 U736 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NOR2_X1 U737 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NOR2_X1 U738 ( .A1(n1025), .A2(n1026), .ZN(n1023) );
NOR2_X1 U739 ( .A1(n1027), .A2(n1028), .ZN(n1019) );
NOR2_X1 U740 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NOR3_X1 U741 ( .A1(n1028), .A2(n1031), .A3(n1022), .ZN(n1015) );
NOR3_X1 U742 ( .A1(n1028), .A2(n1032), .A3(n1022), .ZN(n1010) );
INV_X1 U743 ( .A(n1033), .ZN(n1022) );
NOR2_X1 U744 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
NOR2_X1 U745 ( .A1(n1036), .A2(n1014), .ZN(n1035) );
NOR3_X1 U746 ( .A1(n1012), .A2(n1031), .A3(n1017), .ZN(n1034) );
NOR3_X1 U747 ( .A1(n1017), .A2(n1037), .A3(n1038), .ZN(n1031) );
NOR3_X1 U748 ( .A1(n1005), .A2(G953), .A3(G952), .ZN(n1003) );
AND4_X1 U749 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1005) );
NOR3_X1 U750 ( .A1(n1043), .A2(n1044), .A3(n1017), .ZN(n1042) );
INV_X1 U751 ( .A(n1045), .ZN(n1017) );
INV_X1 U752 ( .A(n1026), .ZN(n1043) );
NOR3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1041) );
NOR2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1047) );
XOR2_X1 U756 ( .A(n1053), .B(n1054), .Z(n1052) );
XOR2_X1 U757 ( .A(KEYINPUT50), .B(KEYINPUT5), .Z(n1054) );
INV_X1 U758 ( .A(n1055), .ZN(n1051) );
XOR2_X1 U759 ( .A(n1056), .B(n1057), .Z(n1046) );
NOR2_X1 U760 ( .A1(n1058), .A2(KEYINPUT48), .ZN(n1057) );
NOR3_X1 U761 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1040) );
XOR2_X1 U762 ( .A(n1062), .B(KEYINPUT37), .Z(n1061) );
XNOR2_X1 U763 ( .A(n1063), .B(KEYINPUT12), .ZN(n1060) );
NOR2_X1 U764 ( .A1(KEYINPUT44), .A2(n1064), .ZN(n1059) );
NOR3_X1 U765 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1039) );
NOR2_X1 U766 ( .A1(G478), .A2(n1068), .ZN(n1067) );
NOR2_X1 U767 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
XOR2_X1 U768 ( .A(KEYINPUT42), .B(n1071), .Z(n1070) );
NOR3_X1 U769 ( .A1(n1072), .A2(n1071), .A3(n1069), .ZN(n1066) );
INV_X1 U770 ( .A(KEYINPUT44), .ZN(n1069) );
XOR2_X1 U771 ( .A(KEYINPUT7), .B(n1073), .Z(n1065) );
XOR2_X1 U772 ( .A(n1074), .B(n1075), .Z(G72) );
NOR3_X1 U773 ( .A1(n1076), .A2(KEYINPUT22), .A3(n1077), .ZN(n1075) );
AND2_X1 U774 ( .A1(G227), .A2(G900), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
NAND3_X1 U776 ( .A1(n1080), .A2(n1081), .A3(n1082), .ZN(n1079) );
NAND2_X1 U777 ( .A1(G953), .A2(n1083), .ZN(n1081) );
XOR2_X1 U778 ( .A(KEYINPUT21), .B(n1084), .Z(n1080) );
NAND2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1078) );
INV_X1 U780 ( .A(n1082), .ZN(n1085) );
XOR2_X1 U781 ( .A(n1086), .B(n1087), .Z(n1082) );
XOR2_X1 U782 ( .A(n1088), .B(n1089), .Z(n1087) );
XOR2_X1 U783 ( .A(n1090), .B(n1091), .Z(n1086) );
NOR2_X1 U784 ( .A1(KEYINPUT25), .A2(n1092), .ZN(n1091) );
XOR2_X1 U785 ( .A(n1093), .B(KEYINPUT20), .Z(n1092) );
XOR2_X1 U786 ( .A(n1094), .B(G131), .Z(n1090) );
AND2_X1 U787 ( .A1(n1095), .A2(n1076), .ZN(n1084) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XOR2_X1 U789 ( .A(n1098), .B(n1099), .Z(G69) );
XOR2_X1 U790 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U791 ( .A1(G953), .A2(n1102), .ZN(n1101) );
NAND2_X1 U792 ( .A1(G898), .A2(G224), .ZN(n1102) );
NAND2_X1 U793 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
NAND2_X1 U794 ( .A1(G953), .A2(n1105), .ZN(n1104) );
XOR2_X1 U795 ( .A(n1106), .B(n1107), .Z(n1103) );
XOR2_X1 U796 ( .A(G113), .B(n1108), .Z(n1107) );
NOR2_X1 U797 ( .A1(KEYINPUT23), .A2(n1109), .ZN(n1108) );
INV_X1 U798 ( .A(n1110), .ZN(n1109) );
NOR2_X1 U799 ( .A1(n1111), .A2(G953), .ZN(n1098) );
NOR2_X1 U800 ( .A1(n1112), .A2(n1113), .ZN(G66) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U802 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NOR2_X1 U803 ( .A1(n1112), .A2(n1118), .ZN(G63) );
XOR2_X1 U804 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR2_X1 U805 ( .A1(KEYINPUT15), .A2(n1121), .ZN(n1120) );
XOR2_X1 U806 ( .A(n1122), .B(KEYINPUT57), .Z(n1121) );
NAND2_X1 U807 ( .A1(n1116), .A2(G478), .ZN(n1119) );
NOR2_X1 U808 ( .A1(n1112), .A2(n1123), .ZN(G60) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(n1123) );
NAND3_X1 U810 ( .A1(n1116), .A2(G475), .A3(KEYINPUT28), .ZN(n1124) );
XOR2_X1 U811 ( .A(n1126), .B(n1127), .Z(G6) );
NOR2_X1 U812 ( .A1(KEYINPUT18), .A2(n1128), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n1112), .A2(n1129), .ZN(G57) );
XOR2_X1 U814 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U815 ( .A(n1132), .B(G101), .Z(n1131) );
NAND2_X1 U816 ( .A1(n1116), .A2(G472), .ZN(n1132) );
NAND2_X1 U817 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
NAND2_X1 U818 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U819 ( .A(n1137), .B(KEYINPUT36), .Z(n1135) );
NAND2_X1 U820 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
INV_X1 U821 ( .A(n1136), .ZN(n1139) );
XOR2_X1 U822 ( .A(KEYINPUT46), .B(n1140), .Z(n1138) );
INV_X1 U823 ( .A(n1137), .ZN(n1140) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1137) );
NOR2_X1 U825 ( .A1(KEYINPUT3), .A2(n1143), .ZN(n1142) );
NOR2_X1 U826 ( .A1(n1112), .A2(n1144), .ZN(G54) );
XOR2_X1 U827 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U828 ( .A1(n1116), .A2(G469), .ZN(n1146) );
NAND2_X1 U829 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
NAND2_X1 U830 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XOR2_X1 U831 ( .A(n1088), .B(n1151), .Z(n1150) );
XNOR2_X1 U832 ( .A(n1152), .B(KEYINPUT24), .ZN(n1149) );
XOR2_X1 U833 ( .A(n1153), .B(KEYINPUT11), .Z(n1147) );
NAND2_X1 U834 ( .A1(n1154), .A2(n1152), .ZN(n1153) );
AND3_X1 U835 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1152) );
NAND3_X1 U836 ( .A1(n1158), .A2(n1159), .A3(n1160), .ZN(n1156) );
OR2_X1 U837 ( .A1(n1160), .A2(n1159), .ZN(n1155) );
INV_X1 U838 ( .A(KEYINPUT27), .ZN(n1160) );
XOR2_X1 U839 ( .A(n1161), .B(n1151), .Z(n1154) );
XNOR2_X1 U840 ( .A(n1162), .B(n1163), .ZN(n1151) );
NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n1164), .ZN(n1163) );
NAND2_X1 U842 ( .A1(KEYINPUT0), .A2(n1165), .ZN(n1162) );
NOR2_X1 U843 ( .A1(n1112), .A2(n1166), .ZN(G51) );
XOR2_X1 U844 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U845 ( .A(n1169), .B(n1170), .ZN(n1168) );
NAND2_X1 U846 ( .A1(n1116), .A2(n1171), .ZN(n1169) );
AND2_X1 U847 ( .A1(G902), .A2(n1007), .ZN(n1116) );
NAND3_X1 U848 ( .A1(n1111), .A2(n1096), .A3(n1172), .ZN(n1007) );
XOR2_X1 U849 ( .A(n1097), .B(KEYINPUT26), .Z(n1172) );
AND4_X1 U850 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1096) );
AND4_X1 U851 ( .A1(n1177), .A2(n1178), .A3(n1179), .A4(n1180), .ZN(n1176) );
AND2_X1 U852 ( .A1(n1181), .A2(n1182), .ZN(n1111) );
NOR4_X1 U853 ( .A1(n1183), .A2(n1126), .A3(n1184), .A4(n1002), .ZN(n1182) );
AND3_X1 U854 ( .A1(n1185), .A2(n1186), .A3(n1030), .ZN(n1002) );
NOR4_X1 U855 ( .A1(n1187), .A2(n1188), .A3(n1028), .A4(n1189), .ZN(n1184) );
AND3_X1 U856 ( .A1(n1185), .A2(n1186), .A3(n1029), .ZN(n1126) );
AND4_X1 U857 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1181) );
XOR2_X1 U858 ( .A(n1094), .B(n1194), .Z(n1167) );
NAND2_X1 U859 ( .A1(KEYINPUT38), .A2(n1195), .ZN(n1194) );
XOR2_X1 U860 ( .A(G113), .B(n1196), .Z(n1195) );
NOR2_X1 U861 ( .A1(n1197), .A2(G952), .ZN(n1112) );
XOR2_X1 U862 ( .A(G953), .B(KEYINPUT41), .Z(n1197) );
XNOR2_X1 U863 ( .A(G146), .B(n1175), .ZN(G48) );
NAND3_X1 U864 ( .A1(n1198), .A2(n1029), .A3(n1024), .ZN(n1175) );
XOR2_X1 U865 ( .A(n1173), .B(n1199), .Z(G45) );
XOR2_X1 U866 ( .A(n1200), .B(KEYINPUT16), .Z(n1199) );
NAND3_X1 U867 ( .A1(n1024), .A2(n1201), .A3(n1202), .ZN(n1173) );
NOR3_X1 U868 ( .A1(n1189), .A2(n1203), .A3(n1204), .ZN(n1202) );
INV_X1 U869 ( .A(n1037), .ZN(n1189) );
XNOR2_X1 U870 ( .A(G140), .B(n1174), .ZN(G42) );
NAND3_X1 U871 ( .A1(n1029), .A2(n1038), .A3(n1205), .ZN(n1174) );
XNOR2_X1 U872 ( .A(G137), .B(n1097), .ZN(G39) );
NAND2_X1 U873 ( .A1(n1205), .A2(n1206), .ZN(n1097) );
XOR2_X1 U874 ( .A(n1180), .B(n1207), .Z(G36) );
NOR2_X1 U875 ( .A1(G134), .A2(KEYINPUT63), .ZN(n1207) );
NAND3_X1 U876 ( .A1(n1037), .A2(n1030), .A3(n1205), .ZN(n1180) );
XOR2_X1 U877 ( .A(G131), .B(n1208), .Z(G33) );
NOR2_X1 U878 ( .A1(KEYINPUT2), .A2(n1179), .ZN(n1208) );
NAND3_X1 U879 ( .A1(n1037), .A2(n1029), .A3(n1205), .ZN(n1179) );
AND4_X1 U880 ( .A1(n1024), .A2(n1209), .A3(n1210), .A4(n1045), .ZN(n1205) );
INV_X1 U881 ( .A(n1012), .ZN(n1209) );
XOR2_X1 U882 ( .A(n1211), .B(KEYINPUT53), .Z(n1024) );
XNOR2_X1 U883 ( .A(G128), .B(n1178), .ZN(G30) );
NAND3_X1 U884 ( .A1(n1030), .A2(n1212), .A3(n1198), .ZN(n1178) );
AND3_X1 U885 ( .A1(n1073), .A2(n1063), .A3(n1201), .ZN(n1198) );
INV_X1 U886 ( .A(n1211), .ZN(n1212) );
NAND2_X1 U887 ( .A1(n1213), .A2(n1214), .ZN(G3) );
OR2_X1 U888 ( .A1(n1193), .A2(G101), .ZN(n1214) );
XOR2_X1 U889 ( .A(n1215), .B(KEYINPUT29), .Z(n1213) );
NAND2_X1 U890 ( .A1(G101), .A2(n1193), .ZN(n1215) );
NAND3_X1 U891 ( .A1(n1186), .A2(n1033), .A3(n1037), .ZN(n1193) );
XOR2_X1 U892 ( .A(n1094), .B(n1177), .Z(G27) );
NAND4_X1 U893 ( .A1(n1201), .A2(n1029), .A3(n1216), .A4(n1038), .ZN(n1177) );
AND2_X1 U894 ( .A1(n1217), .A2(n1210), .ZN(n1201) );
NAND2_X1 U895 ( .A1(n1009), .A2(n1218), .ZN(n1210) );
NAND4_X1 U896 ( .A1(G953), .A2(G902), .A3(n1219), .A4(n1083), .ZN(n1218) );
INV_X1 U897 ( .A(G900), .ZN(n1083) );
XOR2_X1 U898 ( .A(n1220), .B(G122), .Z(G24) );
NAND2_X1 U899 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND4_X1 U900 ( .A1(n1223), .A2(n1036), .A3(n1224), .A4(n1225), .ZN(n1222) );
INV_X1 U901 ( .A(KEYINPUT30), .ZN(n1225) );
NAND2_X1 U902 ( .A1(n1183), .A2(KEYINPUT30), .ZN(n1221) );
AND2_X1 U903 ( .A1(n1224), .A2(n1226), .ZN(n1183) );
NOR4_X1 U904 ( .A1(n1028), .A2(n1014), .A3(n1204), .A4(n1203), .ZN(n1224) );
XNOR2_X1 U905 ( .A(G119), .B(n1192), .ZN(G21) );
NAND3_X1 U906 ( .A1(n1216), .A2(n1226), .A3(n1206), .ZN(n1192) );
AND3_X1 U907 ( .A1(n1073), .A2(n1063), .A3(n1033), .ZN(n1206) );
XNOR2_X1 U908 ( .A(G116), .B(n1227), .ZN(G18) );
NAND4_X1 U909 ( .A1(n1228), .A2(n1037), .A3(n1229), .A4(n1216), .ZN(n1227) );
AND2_X1 U910 ( .A1(n1223), .A2(n1030), .ZN(n1229) );
XOR2_X1 U911 ( .A(n1036), .B(KEYINPUT43), .Z(n1228) );
XOR2_X1 U912 ( .A(n1230), .B(n1191), .Z(G15) );
NAND4_X1 U913 ( .A1(n1037), .A2(n1029), .A3(n1216), .A4(n1226), .ZN(n1191) );
INV_X1 U914 ( .A(n1187), .ZN(n1226) );
INV_X1 U915 ( .A(n1028), .ZN(n1216) );
NAND2_X1 U916 ( .A1(n1231), .A2(n1026), .ZN(n1028) );
AND2_X1 U917 ( .A1(n1232), .A2(n1233), .ZN(n1029) );
XNOR2_X1 U918 ( .A(KEYINPUT59), .B(n1204), .ZN(n1232) );
NOR2_X1 U919 ( .A1(n1063), .A2(n1234), .ZN(n1037) );
XOR2_X1 U920 ( .A(n1190), .B(n1235), .Z(G12) );
NAND2_X1 U921 ( .A1(KEYINPUT8), .A2(G110), .ZN(n1235) );
NAND3_X1 U922 ( .A1(n1033), .A2(n1038), .A3(n1186), .ZN(n1190) );
NOR2_X1 U923 ( .A1(n1187), .A2(n1211), .ZN(n1186) );
NAND2_X1 U924 ( .A1(n1025), .A2(n1026), .ZN(n1211) );
NAND2_X1 U925 ( .A1(G221), .A2(n1236), .ZN(n1026) );
INV_X1 U926 ( .A(n1231), .ZN(n1025) );
NOR2_X1 U927 ( .A1(n1237), .A2(n1044), .ZN(n1231) );
NOR2_X1 U928 ( .A1(n1055), .A2(n1053), .ZN(n1044) );
AND2_X1 U929 ( .A1(n1238), .A2(n1055), .ZN(n1237) );
NAND2_X1 U930 ( .A1(n1239), .A2(n1240), .ZN(n1055) );
XOR2_X1 U931 ( .A(n1241), .B(n1242), .Z(n1239) );
NAND2_X1 U932 ( .A1(KEYINPUT9), .A2(n1243), .ZN(n1242) );
XOR2_X1 U933 ( .A(n1244), .B(n1165), .Z(n1243) );
NOR2_X1 U934 ( .A1(KEYINPUT52), .A2(n1245), .ZN(n1244) );
XOR2_X1 U935 ( .A(n1164), .B(n1088), .Z(n1245) );
INV_X1 U936 ( .A(n1161), .ZN(n1088) );
XNOR2_X1 U937 ( .A(G128), .B(n1246), .ZN(n1161) );
NAND2_X1 U938 ( .A1(n1247), .A2(n1248), .ZN(n1164) );
NAND2_X1 U939 ( .A1(n1249), .A2(n1250), .ZN(n1248) );
INV_X1 U940 ( .A(KEYINPUT61), .ZN(n1250) );
NAND3_X1 U941 ( .A1(G101), .A2(n1251), .A3(KEYINPUT61), .ZN(n1247) );
NAND2_X1 U942 ( .A1(n1252), .A2(n1157), .ZN(n1241) );
OR2_X1 U943 ( .A1(n1159), .A2(n1158), .ZN(n1157) );
NAND2_X1 U944 ( .A1(n1158), .A2(n1159), .ZN(n1252) );
NAND2_X1 U945 ( .A1(G227), .A2(n1076), .ZN(n1159) );
XNOR2_X1 U946 ( .A(n1253), .B(n1089), .ZN(n1158) );
XNOR2_X1 U947 ( .A(n1053), .B(KEYINPUT49), .ZN(n1238) );
XOR2_X1 U948 ( .A(G469), .B(KEYINPUT13), .Z(n1053) );
NAND2_X1 U949 ( .A1(n1217), .A2(n1223), .ZN(n1187) );
NAND2_X1 U950 ( .A1(n1009), .A2(n1254), .ZN(n1223) );
NAND4_X1 U951 ( .A1(G953), .A2(G902), .A3(n1219), .A4(n1105), .ZN(n1254) );
INV_X1 U952 ( .A(G898), .ZN(n1105) );
NAND3_X1 U953 ( .A1(n1219), .A2(n1076), .A3(G952), .ZN(n1009) );
NAND2_X1 U954 ( .A1(G237), .A2(G234), .ZN(n1219) );
INV_X1 U955 ( .A(n1036), .ZN(n1217) );
NAND2_X1 U956 ( .A1(n1012), .A2(n1045), .ZN(n1036) );
NAND2_X1 U957 ( .A1(G214), .A2(n1255), .ZN(n1045) );
XOR2_X1 U958 ( .A(n1058), .B(n1171), .Z(n1012) );
INV_X1 U959 ( .A(n1056), .ZN(n1171) );
NAND2_X1 U960 ( .A1(G210), .A2(n1255), .ZN(n1056) );
NAND2_X1 U961 ( .A1(n1256), .A2(n1240), .ZN(n1255) );
INV_X1 U962 ( .A(G237), .ZN(n1256) );
AND2_X1 U963 ( .A1(n1257), .A2(n1240), .ZN(n1058) );
XOR2_X1 U964 ( .A(n1258), .B(n1259), .Z(n1257) );
XNOR2_X1 U965 ( .A(n1196), .B(n1170), .ZN(n1258) );
XNOR2_X1 U966 ( .A(n1260), .B(n1261), .ZN(n1170) );
NAND2_X1 U967 ( .A1(G224), .A2(n1076), .ZN(n1260) );
XNOR2_X1 U968 ( .A(n1262), .B(n1263), .ZN(n1196) );
INV_X1 U969 ( .A(n1106), .ZN(n1263) );
XNOR2_X1 U970 ( .A(n1249), .B(n1264), .ZN(n1106) );
XNOR2_X1 U971 ( .A(n1265), .B(n1251), .ZN(n1249) );
XOR2_X1 U972 ( .A(G104), .B(G107), .Z(n1251) );
NAND2_X1 U973 ( .A1(KEYINPUT10), .A2(n1110), .ZN(n1262) );
XOR2_X1 U974 ( .A(n1266), .B(n1267), .Z(n1110) );
XOR2_X1 U975 ( .A(KEYINPUT17), .B(G122), .Z(n1267) );
NAND2_X1 U976 ( .A1(KEYINPUT34), .A2(n1253), .ZN(n1266) );
INV_X1 U977 ( .A(G110), .ZN(n1253) );
NAND2_X1 U978 ( .A1(n1268), .A2(n1269), .ZN(n1038) );
OR2_X1 U979 ( .A1(n1014), .A2(KEYINPUT62), .ZN(n1269) );
INV_X1 U980 ( .A(n1185), .ZN(n1014) );
NOR2_X1 U981 ( .A1(n1063), .A2(n1073), .ZN(n1185) );
INV_X1 U982 ( .A(n1234), .ZN(n1073) );
NAND3_X1 U983 ( .A1(n1063), .A2(n1234), .A3(KEYINPUT62), .ZN(n1268) );
XOR2_X1 U984 ( .A(n1270), .B(G472), .Z(n1234) );
NAND2_X1 U985 ( .A1(n1271), .A2(n1272), .ZN(n1270) );
XOR2_X1 U986 ( .A(n1273), .B(n1274), .Z(n1272) );
INV_X1 U987 ( .A(n1141), .ZN(n1274) );
XNOR2_X1 U988 ( .A(n1165), .B(n1261), .ZN(n1141) );
XOR2_X1 U989 ( .A(n1246), .B(n1275), .Z(n1261) );
NOR2_X1 U990 ( .A1(G128), .A2(KEYINPUT1), .ZN(n1275) );
XOR2_X1 U991 ( .A(G143), .B(G146), .Z(n1246) );
XOR2_X1 U992 ( .A(G131), .B(n1276), .Z(n1165) );
INV_X1 U993 ( .A(n1093), .ZN(n1276) );
XNOR2_X1 U994 ( .A(G137), .B(G134), .ZN(n1093) );
XOR2_X1 U995 ( .A(n1277), .B(n1278), .Z(n1273) );
NOR2_X1 U996 ( .A1(KEYINPUT6), .A2(n1136), .ZN(n1278) );
XOR2_X1 U997 ( .A(n1279), .B(n1264), .Z(n1136) );
XOR2_X1 U998 ( .A(G116), .B(n1280), .Z(n1264) );
XOR2_X1 U999 ( .A(KEYINPUT51), .B(G119), .Z(n1280) );
NAND2_X1 U1000 ( .A1(KEYINPUT58), .A2(G113), .ZN(n1279) );
NAND2_X1 U1001 ( .A1(n1281), .A2(n1282), .ZN(n1277) );
NAND2_X1 U1002 ( .A1(n1143), .A2(n1265), .ZN(n1282) );
XOR2_X1 U1003 ( .A(n1283), .B(KEYINPUT55), .Z(n1281) );
OR2_X1 U1004 ( .A1(n1265), .A2(n1143), .ZN(n1283) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1284), .ZN(n1143) );
INV_X1 U1006 ( .A(G101), .ZN(n1265) );
XOR2_X1 U1007 ( .A(n1240), .B(KEYINPUT39), .Z(n1271) );
XNOR2_X1 U1008 ( .A(n1285), .B(n1117), .ZN(n1063) );
AND2_X1 U1009 ( .A1(G217), .A2(n1236), .ZN(n1117) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1240), .ZN(n1236) );
NAND2_X1 U1011 ( .A1(n1240), .A2(n1114), .ZN(n1285) );
NAND2_X1 U1012 ( .A1(n1286), .A2(n1287), .ZN(n1114) );
NAND2_X1 U1013 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XOR2_X1 U1014 ( .A(n1290), .B(KEYINPUT40), .Z(n1286) );
OR2_X1 U1015 ( .A1(n1289), .A2(n1288), .ZN(n1290) );
XNOR2_X1 U1016 ( .A(n1291), .B(n1292), .ZN(n1288) );
XOR2_X1 U1017 ( .A(KEYINPUT19), .B(G137), .Z(n1292) );
NAND2_X1 U1018 ( .A1(G221), .A2(n1293), .ZN(n1291) );
XNOR2_X1 U1019 ( .A(n1294), .B(n1295), .ZN(n1289) );
XOR2_X1 U1020 ( .A(G119), .B(n1296), .Z(n1295) );
XOR2_X1 U1021 ( .A(G146), .B(G128), .Z(n1296) );
XOR2_X1 U1022 ( .A(n1297), .B(G110), .Z(n1294) );
NAND2_X1 U1023 ( .A1(n1298), .A2(KEYINPUT54), .ZN(n1297) );
XOR2_X1 U1024 ( .A(n1299), .B(n1089), .Z(n1298) );
NAND2_X1 U1025 ( .A1(KEYINPUT32), .A2(n1094), .ZN(n1299) );
INV_X1 U1026 ( .A(G125), .ZN(n1094) );
NAND2_X1 U1027 ( .A1(n1300), .A2(n1301), .ZN(n1033) );
OR2_X1 U1028 ( .A1(n1188), .A2(KEYINPUT59), .ZN(n1301) );
INV_X1 U1029 ( .A(n1030), .ZN(n1188) );
NOR2_X1 U1030 ( .A1(n1233), .A2(n1204), .ZN(n1030) );
NAND3_X1 U1031 ( .A1(n1203), .A2(n1204), .A3(KEYINPUT59), .ZN(n1300) );
XOR2_X1 U1032 ( .A(n1071), .B(n1072), .Z(n1204) );
INV_X1 U1033 ( .A(G478), .ZN(n1072) );
INV_X1 U1034 ( .A(n1064), .ZN(n1071) );
NAND2_X1 U1035 ( .A1(n1302), .A2(n1240), .ZN(n1064) );
INV_X1 U1036 ( .A(n1122), .ZN(n1302) );
XOR2_X1 U1037 ( .A(n1303), .B(n1304), .Z(n1122) );
XOR2_X1 U1038 ( .A(G107), .B(n1305), .Z(n1304) );
XOR2_X1 U1039 ( .A(G122), .B(G116), .Z(n1305) );
XOR2_X1 U1040 ( .A(n1306), .B(n1307), .Z(n1303) );
NOR2_X1 U1041 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
XOR2_X1 U1042 ( .A(n1310), .B(KEYINPUT14), .Z(n1309) );
NAND2_X1 U1043 ( .A1(G134), .A2(n1311), .ZN(n1310) );
NOR2_X1 U1044 ( .A1(G134), .A2(n1311), .ZN(n1308) );
XOR2_X1 U1045 ( .A(G143), .B(G128), .Z(n1311) );
NAND2_X1 U1046 ( .A1(G217), .A2(n1293), .ZN(n1306) );
AND2_X1 U1047 ( .A1(G234), .A2(n1076), .ZN(n1293) );
INV_X1 U1048 ( .A(G953), .ZN(n1076) );
INV_X1 U1049 ( .A(n1233), .ZN(n1203) );
NAND2_X1 U1050 ( .A1(n1062), .A2(n1312), .ZN(n1233) );
NAND2_X1 U1051 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
XOR2_X1 U1052 ( .A(KEYINPUT60), .B(G475), .Z(n1313) );
NAND2_X1 U1053 ( .A1(n1049), .A2(n1050), .ZN(n1062) );
INV_X1 U1054 ( .A(G475), .ZN(n1050) );
INV_X1 U1055 ( .A(n1314), .ZN(n1049) );
NAND2_X1 U1056 ( .A1(n1125), .A2(n1240), .ZN(n1314) );
INV_X1 U1057 ( .A(G902), .ZN(n1240) );
XOR2_X1 U1058 ( .A(n1315), .B(n1316), .Z(n1125) );
XNOR2_X1 U1059 ( .A(n1259), .B(n1317), .ZN(n1316) );
XOR2_X1 U1060 ( .A(n1318), .B(n1089), .Z(n1317) );
XOR2_X1 U1061 ( .A(G140), .B(KEYINPUT35), .Z(n1089) );
NAND2_X1 U1062 ( .A1(KEYINPUT56), .A2(n1319), .ZN(n1318) );
XOR2_X1 U1063 ( .A(KEYINPUT4), .B(G122), .Z(n1319) );
XNOR2_X1 U1064 ( .A(n1230), .B(G125), .ZN(n1259) );
INV_X1 U1065 ( .A(G113), .ZN(n1230) );
XOR2_X1 U1066 ( .A(n1320), .B(n1321), .Z(n1315) );
NOR2_X1 U1067 ( .A1(KEYINPUT45), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1068 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1069 ( .A(KEYINPUT31), .B(G131), .Z(n1324) );
XOR2_X1 U1070 ( .A(n1325), .B(n1326), .Z(n1323) );
NOR2_X1 U1071 ( .A1(KEYINPUT47), .A2(n1200), .ZN(n1326) );
INV_X1 U1072 ( .A(G143), .ZN(n1200) );
NAND2_X1 U1073 ( .A1(G214), .A2(n1284), .ZN(n1325) );
NOR2_X1 U1074 ( .A1(G953), .A2(G237), .ZN(n1284) );
XOR2_X1 U1075 ( .A(n1128), .B(G146), .Z(n1320) );
INV_X1 U1076 ( .A(G104), .ZN(n1128) );
endmodule


