//Key = 1011110110110001000110001000000011101111101010110101100001000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286;

XOR2_X1 U709 ( .A(G107), .B(n973), .Z(G9) );
NOR3_X1 U710 ( .A1(n974), .A2(n975), .A3(n976), .ZN(n973) );
NOR2_X1 U711 ( .A1(n977), .A2(n978), .ZN(G75) );
NOR4_X1 U712 ( .A1(G953), .A2(n979), .A3(n980), .A4(n981), .ZN(n978) );
INV_X1 U713 ( .A(n982), .ZN(n981) );
NOR2_X1 U714 ( .A1(n983), .A2(n984), .ZN(n980) );
NOR2_X1 U715 ( .A1(n985), .A2(n986), .ZN(n983) );
NOR3_X1 U716 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
NOR2_X1 U717 ( .A1(n990), .A2(n991), .ZN(n988) );
AND2_X1 U718 ( .A1(n992), .A2(n993), .ZN(n991) );
NOR2_X1 U719 ( .A1(n994), .A2(n995), .ZN(n990) );
NOR2_X1 U720 ( .A1(n996), .A2(n997), .ZN(n994) );
AND2_X1 U721 ( .A1(n998), .A2(n992), .ZN(n997) );
NOR2_X1 U722 ( .A1(n999), .A2(n1000), .ZN(n996) );
NOR3_X1 U723 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n999) );
NOR3_X1 U724 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1003) );
INV_X1 U725 ( .A(KEYINPUT7), .ZN(n1004) );
NOR2_X1 U726 ( .A1(KEYINPUT7), .A2(n1007), .ZN(n1002) );
NOR4_X1 U727 ( .A1(n1008), .A2(n995), .A3(n1000), .A4(n1007), .ZN(n985) );
NOR2_X1 U728 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
NOR2_X1 U729 ( .A1(n1011), .A2(n989), .ZN(n1010) );
NOR2_X1 U730 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR2_X1 U731 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
XNOR2_X1 U732 ( .A(n1016), .B(KEYINPUT45), .ZN(n1014) );
NOR2_X1 U733 ( .A1(n1017), .A2(n987), .ZN(n1009) );
NOR3_X1 U734 ( .A1(n979), .A2(G953), .A3(G952), .ZN(n977) );
AND4_X1 U735 ( .A1(n1018), .A2(n1015), .A3(n1019), .A4(n1020), .ZN(n979) );
NOR4_X1 U736 ( .A1(n1021), .A2(n1022), .A3(n989), .A4(n1023), .ZN(n1020) );
XNOR2_X1 U737 ( .A(n1024), .B(n1025), .ZN(n1023) );
NOR2_X1 U738 ( .A1(n1026), .A2(n1027), .ZN(n1022) );
INV_X1 U739 ( .A(KEYINPUT31), .ZN(n1027) );
NOR2_X1 U740 ( .A1(n1005), .A2(n1006), .ZN(n1026) );
NOR2_X1 U741 ( .A1(KEYINPUT31), .A2(n992), .ZN(n1021) );
XOR2_X1 U742 ( .A(KEYINPUT38), .B(n1028), .Z(n1018) );
XOR2_X1 U743 ( .A(n1029), .B(n1030), .Z(G72) );
XOR2_X1 U744 ( .A(n1031), .B(n1032), .Z(n1030) );
NAND2_X1 U745 ( .A1(G953), .A2(n1033), .ZN(n1032) );
NAND2_X1 U746 ( .A1(G900), .A2(G227), .ZN(n1033) );
NAND2_X1 U747 ( .A1(n1034), .A2(n1035), .ZN(n1031) );
NAND2_X1 U748 ( .A1(G953), .A2(n1036), .ZN(n1035) );
XOR2_X1 U749 ( .A(n1037), .B(n1038), .Z(n1034) );
XOR2_X1 U750 ( .A(n1039), .B(n1040), .Z(n1038) );
XOR2_X1 U751 ( .A(n1041), .B(n1042), .Z(n1039) );
XOR2_X1 U752 ( .A(n1043), .B(n1044), .Z(n1037) );
NOR2_X1 U753 ( .A1(KEYINPUT23), .A2(G137), .ZN(n1044) );
XNOR2_X1 U754 ( .A(KEYINPUT26), .B(KEYINPUT21), .ZN(n1043) );
NOR2_X1 U755 ( .A1(n1045), .A2(G953), .ZN(n1029) );
NOR2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
XOR2_X1 U757 ( .A(n1048), .B(n1049), .Z(G69) );
XOR2_X1 U758 ( .A(n1050), .B(n1051), .Z(n1049) );
NAND2_X1 U759 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U760 ( .A1(G953), .A2(n1054), .ZN(n1053) );
XOR2_X1 U761 ( .A(n1055), .B(n1056), .Z(n1052) );
NAND2_X1 U762 ( .A1(KEYINPUT11), .A2(n1057), .ZN(n1055) );
NAND2_X1 U763 ( .A1(n1058), .A2(n1059), .ZN(n1050) );
NOR2_X1 U764 ( .A1(n1060), .A2(n1058), .ZN(n1048) );
AND2_X1 U765 ( .A1(G224), .A2(G898), .ZN(n1060) );
NOR2_X1 U766 ( .A1(n1061), .A2(n1062), .ZN(G66) );
NOR3_X1 U767 ( .A1(n1024), .A2(n1063), .A3(n1064), .ZN(n1062) );
NOR3_X1 U768 ( .A1(n1065), .A2(n1025), .A3(n1066), .ZN(n1064) );
INV_X1 U769 ( .A(n1067), .ZN(n1065) );
NOR2_X1 U770 ( .A1(n1068), .A2(n1067), .ZN(n1063) );
NOR2_X1 U771 ( .A1(n982), .A2(n1025), .ZN(n1068) );
NOR2_X1 U772 ( .A1(n1061), .A2(n1069), .ZN(G63) );
XOR2_X1 U773 ( .A(n1070), .B(n1071), .Z(n1069) );
NAND3_X1 U774 ( .A1(n1072), .A2(G478), .A3(KEYINPUT3), .ZN(n1071) );
NOR2_X1 U775 ( .A1(n1061), .A2(n1073), .ZN(G60) );
XOR2_X1 U776 ( .A(n1074), .B(n1075), .Z(n1073) );
NAND2_X1 U777 ( .A1(n1072), .A2(G475), .ZN(n1074) );
XNOR2_X1 U778 ( .A(G104), .B(n1076), .ZN(G6) );
NAND4_X1 U779 ( .A1(n1077), .A2(KEYINPUT39), .A3(n1078), .A4(n1079), .ZN(n1076) );
XNOR2_X1 U780 ( .A(n1013), .B(KEYINPUT4), .ZN(n1077) );
NOR2_X1 U781 ( .A1(n1061), .A2(n1080), .ZN(G57) );
XOR2_X1 U782 ( .A(n1081), .B(n1082), .Z(n1080) );
XOR2_X1 U783 ( .A(n1083), .B(n1084), .Z(n1082) );
XOR2_X1 U784 ( .A(n1085), .B(n1086), .Z(n1084) );
NOR2_X1 U785 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR3_X1 U786 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1088) );
NOR2_X1 U787 ( .A1(KEYINPUT16), .A2(n1092), .ZN(n1085) );
XNOR2_X1 U788 ( .A(n1093), .B(KEYINPUT20), .ZN(n1092) );
XOR2_X1 U789 ( .A(KEYINPUT28), .B(KEYINPUT18), .Z(n1083) );
XOR2_X1 U790 ( .A(n1094), .B(n1095), .Z(n1081) );
XOR2_X1 U791 ( .A(n1096), .B(n1097), .Z(n1094) );
NAND2_X1 U792 ( .A1(n1072), .A2(G472), .ZN(n1096) );
NOR2_X1 U793 ( .A1(n1098), .A2(n1099), .ZN(G54) );
XOR2_X1 U794 ( .A(n1100), .B(n1101), .Z(n1099) );
XNOR2_X1 U795 ( .A(n1102), .B(n1093), .ZN(n1101) );
XOR2_X1 U796 ( .A(n1103), .B(n1104), .Z(n1100) );
AND2_X1 U797 ( .A1(G469), .A2(n1072), .ZN(n1104) );
NAND3_X1 U798 ( .A1(KEYINPUT5), .A2(n1105), .A3(n1106), .ZN(n1103) );
XOR2_X1 U799 ( .A(n1107), .B(KEYINPUT53), .Z(n1106) );
NAND2_X1 U800 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
OR2_X1 U801 ( .A1(n1109), .A2(n1108), .ZN(n1105) );
XOR2_X1 U802 ( .A(n1110), .B(n1111), .Z(n1109) );
NAND2_X1 U803 ( .A1(KEYINPUT47), .A2(n1112), .ZN(n1110) );
NOR2_X1 U804 ( .A1(G952), .A2(n1113), .ZN(n1098) );
XNOR2_X1 U805 ( .A(KEYINPUT33), .B(n1058), .ZN(n1113) );
NOR2_X1 U806 ( .A1(n1061), .A2(n1114), .ZN(G51) );
NOR3_X1 U807 ( .A1(n1115), .A2(n1116), .A3(n1117), .ZN(n1114) );
AND2_X1 U808 ( .A1(n1118), .A2(KEYINPUT62), .ZN(n1117) );
NOR3_X1 U809 ( .A1(KEYINPUT62), .A2(n1119), .A3(n1118), .ZN(n1116) );
NOR4_X1 U810 ( .A1(KEYINPUT27), .A2(n1091), .A3(n1066), .A4(n1120), .ZN(n1119) );
INV_X1 U811 ( .A(KEYINPUT44), .ZN(n1120) );
NOR4_X1 U812 ( .A1(KEYINPUT27), .A2(n1121), .A3(n1091), .A4(n1066), .ZN(n1115) );
INV_X1 U813 ( .A(n1072), .ZN(n1066) );
NOR2_X1 U814 ( .A1(n1122), .A2(n982), .ZN(n1072) );
NOR3_X1 U815 ( .A1(n1047), .A2(n1059), .A3(n1123), .ZN(n982) );
XOR2_X1 U816 ( .A(n1046), .B(KEYINPUT56), .Z(n1123) );
NAND4_X1 U817 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1059) );
NOR4_X1 U818 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1127) );
NAND4_X1 U819 ( .A1(n1013), .A2(n1079), .A3(n1132), .A4(n1133), .ZN(n1126) );
NAND2_X1 U820 ( .A1(n1017), .A2(n1134), .ZN(n1133) );
INV_X1 U821 ( .A(KEYINPUT60), .ZN(n1134) );
NOR2_X1 U822 ( .A1(n1078), .A2(n1135), .ZN(n1017) );
NAND2_X1 U823 ( .A1(KEYINPUT60), .A2(n1135), .ZN(n1132) );
INV_X1 U824 ( .A(n975), .ZN(n1079) );
NAND4_X1 U825 ( .A1(n1001), .A2(n1136), .A3(n1019), .A4(n1137), .ZN(n975) );
NAND4_X1 U826 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1047) );
NOR4_X1 U827 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
INV_X1 U828 ( .A(n1146), .ZN(n1140) );
NOR2_X1 U829 ( .A1(n1147), .A2(KEYINPUT62), .ZN(n1121) );
AND2_X1 U830 ( .A1(n1118), .A2(KEYINPUT44), .ZN(n1147) );
XOR2_X1 U831 ( .A(n1148), .B(n1149), .Z(n1118) );
NOR2_X1 U832 ( .A1(KEYINPUT25), .A2(n1095), .ZN(n1149) );
NOR2_X1 U833 ( .A1(n1058), .A2(G952), .ZN(n1061) );
XNOR2_X1 U834 ( .A(G146), .B(n1138), .ZN(G48) );
NAND3_X1 U835 ( .A1(n1078), .A2(n1013), .A3(n1150), .ZN(n1138) );
XOR2_X1 U836 ( .A(n1151), .B(n1152), .Z(G45) );
XNOR2_X1 U837 ( .A(G143), .B(KEYINPUT6), .ZN(n1152) );
NAND2_X1 U838 ( .A1(KEYINPUT52), .A2(n1146), .ZN(n1151) );
NOR4_X1 U839 ( .A1(n1153), .A2(n974), .A3(n1154), .A4(n1155), .ZN(n1146) );
XNOR2_X1 U840 ( .A(G140), .B(n1139), .ZN(G42) );
NAND3_X1 U841 ( .A1(n1156), .A2(n1001), .A3(n1157), .ZN(n1139) );
XNOR2_X1 U842 ( .A(G137), .B(n1158), .ZN(G39) );
NAND2_X1 U843 ( .A1(KEYINPUT34), .A2(n1046), .ZN(n1158) );
AND3_X1 U844 ( .A1(n1150), .A2(n1159), .A3(n1157), .ZN(n1046) );
INV_X1 U845 ( .A(n987), .ZN(n1157) );
XOR2_X1 U846 ( .A(G134), .B(n1145), .Z(G36) );
NOR3_X1 U847 ( .A1(n987), .A2(n976), .A3(n1153), .ZN(n1145) );
XNOR2_X1 U848 ( .A(n1144), .B(n1160), .ZN(G33) );
XNOR2_X1 U849 ( .A(G131), .B(KEYINPUT48), .ZN(n1160) );
NOR3_X1 U850 ( .A1(n987), .A2(n1161), .A3(n1153), .ZN(n1144) );
NAND3_X1 U851 ( .A1(n1001), .A2(n1162), .A3(n993), .ZN(n1153) );
INV_X1 U852 ( .A(n1078), .ZN(n1161) );
NAND2_X1 U853 ( .A1(n1016), .A2(n1015), .ZN(n987) );
XNOR2_X1 U854 ( .A(n1163), .B(n1143), .ZN(G30) );
AND3_X1 U855 ( .A1(n1013), .A2(n1135), .A3(n1150), .ZN(n1143) );
AND4_X1 U856 ( .A1(n998), .A2(n1001), .A3(n995), .A4(n1162), .ZN(n1150) );
XNOR2_X1 U857 ( .A(n1090), .B(n1130), .ZN(G3) );
AND2_X1 U858 ( .A1(n1164), .A2(n993), .ZN(n1130) );
XOR2_X1 U859 ( .A(G125), .B(n1142), .Z(G27) );
AND3_X1 U860 ( .A1(n1156), .A2(n1013), .A3(n992), .ZN(n1142) );
AND4_X1 U861 ( .A1(n998), .A2(n1078), .A3(n1019), .A4(n1162), .ZN(n1156) );
NAND2_X1 U862 ( .A1(n984), .A2(n1165), .ZN(n1162) );
NAND2_X1 U863 ( .A1(n1166), .A2(n1036), .ZN(n1165) );
INV_X1 U864 ( .A(G900), .ZN(n1036) );
XOR2_X1 U865 ( .A(G122), .B(n1167), .Z(G24) );
NOR2_X1 U866 ( .A1(KEYINPUT41), .A2(n1124), .ZN(n1167) );
NAND3_X1 U867 ( .A1(n1168), .A2(n1136), .A3(n1169), .ZN(n1124) );
NOR3_X1 U868 ( .A1(n995), .A2(n1155), .A3(n1154), .ZN(n1169) );
NAND2_X1 U869 ( .A1(n1170), .A2(n1171), .ZN(G21) );
NAND2_X1 U870 ( .A1(G119), .A2(n1125), .ZN(n1171) );
XOR2_X1 U871 ( .A(n1172), .B(KEYINPUT14), .Z(n1170) );
OR2_X1 U872 ( .A1(n1125), .A2(G119), .ZN(n1172) );
NAND4_X1 U873 ( .A1(n998), .A2(n1168), .A3(n1159), .A4(n995), .ZN(n1125) );
XNOR2_X1 U874 ( .A(n1173), .B(n1131), .ZN(G18) );
AND3_X1 U875 ( .A1(n993), .A2(n1135), .A3(n1168), .ZN(n1131) );
INV_X1 U876 ( .A(n976), .ZN(n1135) );
NAND2_X1 U877 ( .A1(n1155), .A2(n1174), .ZN(n976) );
XOR2_X1 U878 ( .A(G113), .B(n1129), .Z(G15) );
AND3_X1 U879 ( .A1(n993), .A2(n1078), .A3(n1168), .ZN(n1129) );
AND3_X1 U880 ( .A1(n1013), .A2(n1137), .A3(n992), .ZN(n1168) );
INV_X1 U881 ( .A(n1007), .ZN(n992) );
NAND2_X1 U882 ( .A1(n1175), .A2(n1006), .ZN(n1007) );
INV_X1 U883 ( .A(n1005), .ZN(n1175) );
NOR2_X1 U884 ( .A1(n1174), .A2(n1155), .ZN(n1078) );
NOR2_X1 U885 ( .A1(n1000), .A2(n1019), .ZN(n993) );
XOR2_X1 U886 ( .A(G110), .B(n1128), .Z(G12) );
AND3_X1 U887 ( .A1(n998), .A2(n1019), .A3(n1164), .ZN(n1128) );
AND4_X1 U888 ( .A1(n1159), .A2(n1013), .A3(n1001), .A4(n1137), .ZN(n1164) );
NAND2_X1 U889 ( .A1(n984), .A2(n1176), .ZN(n1137) );
NAND2_X1 U890 ( .A1(n1166), .A2(n1054), .ZN(n1176) );
INV_X1 U891 ( .A(G898), .ZN(n1054) );
AND3_X1 U892 ( .A1(n1177), .A2(n1178), .A3(G953), .ZN(n1166) );
XNOR2_X1 U893 ( .A(KEYINPUT58), .B(n1122), .ZN(n1177) );
NAND3_X1 U894 ( .A1(n1178), .A2(n1058), .A3(n1179), .ZN(n984) );
XOR2_X1 U895 ( .A(KEYINPUT61), .B(G952), .Z(n1179) );
INV_X1 U896 ( .A(G953), .ZN(n1058) );
NAND2_X1 U897 ( .A1(G237), .A2(G234), .ZN(n1178) );
AND2_X1 U898 ( .A1(n1005), .A2(n1006), .ZN(n1001) );
NAND2_X1 U899 ( .A1(G221), .A2(n1180), .ZN(n1006) );
XNOR2_X1 U900 ( .A(n1181), .B(G469), .ZN(n1005) );
NAND2_X1 U901 ( .A1(n1182), .A2(n1122), .ZN(n1181) );
XOR2_X1 U902 ( .A(n1183), .B(n1184), .Z(n1182) );
XNOR2_X1 U903 ( .A(n1185), .B(n1112), .ZN(n1184) );
XOR2_X1 U904 ( .A(n1186), .B(n1187), .Z(n1183) );
NOR2_X1 U905 ( .A1(KEYINPUT9), .A2(n1111), .ZN(n1187) );
XNOR2_X1 U906 ( .A(G140), .B(KEYINPUT13), .ZN(n1111) );
XOR2_X1 U907 ( .A(n1188), .B(n1108), .Z(n1186) );
AND2_X1 U908 ( .A1(G227), .A2(n1189), .ZN(n1108) );
NAND2_X1 U909 ( .A1(KEYINPUT49), .A2(n1102), .ZN(n1188) );
XOR2_X1 U910 ( .A(n1190), .B(n1057), .Z(n1102) );
INV_X1 U911 ( .A(n1191), .ZN(n1057) );
XOR2_X1 U912 ( .A(n1041), .B(KEYINPUT32), .Z(n1190) );
NAND3_X1 U913 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1041) );
OR2_X1 U914 ( .A1(n1163), .A2(n1195), .ZN(n1194) );
NAND2_X1 U915 ( .A1(n1196), .A2(n1197), .ZN(n1193) );
INV_X1 U916 ( .A(KEYINPUT10), .ZN(n1197) );
NAND2_X1 U917 ( .A1(n1198), .A2(n1163), .ZN(n1196) );
XNOR2_X1 U918 ( .A(KEYINPUT46), .B(n1195), .ZN(n1198) );
NAND2_X1 U919 ( .A1(KEYINPUT10), .A2(n1199), .ZN(n1192) );
NAND2_X1 U920 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND3_X1 U921 ( .A1(KEYINPUT46), .A2(n1163), .A3(n1195), .ZN(n1201) );
OR2_X1 U922 ( .A1(n1195), .A2(KEYINPUT46), .ZN(n1200) );
INV_X1 U923 ( .A(n974), .ZN(n1013) );
NAND2_X1 U924 ( .A1(n1202), .A2(n1015), .ZN(n974) );
OR2_X1 U925 ( .A1(n1203), .A2(n1204), .ZN(n1015) );
INV_X1 U926 ( .A(n1016), .ZN(n1202) );
XOR2_X1 U927 ( .A(n1028), .B(KEYINPUT42), .Z(n1016) );
XNOR2_X1 U928 ( .A(n1205), .B(n1206), .ZN(n1028) );
NOR2_X1 U929 ( .A1(n1204), .A2(n1091), .ZN(n1206) );
INV_X1 U930 ( .A(G210), .ZN(n1091) );
NOR2_X1 U931 ( .A1(G902), .A2(G237), .ZN(n1204) );
NAND2_X1 U932 ( .A1(n1207), .A2(n1122), .ZN(n1205) );
XOR2_X1 U933 ( .A(n1148), .B(n1208), .Z(n1207) );
XNOR2_X1 U934 ( .A(n1095), .B(KEYINPUT8), .ZN(n1208) );
XOR2_X1 U935 ( .A(n1209), .B(n1210), .Z(n1148) );
XNOR2_X1 U936 ( .A(n1211), .B(n1056), .ZN(n1210) );
XOR2_X1 U937 ( .A(n1212), .B(n1213), .Z(n1056) );
XNOR2_X1 U938 ( .A(n1097), .B(G122), .ZN(n1212) );
NAND2_X1 U939 ( .A1(KEYINPUT51), .A2(n1191), .ZN(n1211) );
XOR2_X1 U940 ( .A(G101), .B(n1214), .Z(n1191) );
XOR2_X1 U941 ( .A(G107), .B(G104), .Z(n1214) );
XOR2_X1 U942 ( .A(n1215), .B(G125), .Z(n1209) );
NAND2_X1 U943 ( .A1(G224), .A2(n1189), .ZN(n1215) );
INV_X1 U944 ( .A(n989), .ZN(n1159) );
NAND2_X1 U945 ( .A1(n1154), .A2(n1155), .ZN(n989) );
XOR2_X1 U946 ( .A(n1216), .B(G475), .Z(n1155) );
NAND2_X1 U947 ( .A1(n1075), .A2(n1122), .ZN(n1216) );
XNOR2_X1 U948 ( .A(n1217), .B(n1218), .ZN(n1075) );
XOR2_X1 U949 ( .A(n1219), .B(n1220), .Z(n1218) );
XNOR2_X1 U950 ( .A(G104), .B(n1221), .ZN(n1220) );
NOR2_X1 U951 ( .A1(KEYINPUT50), .A2(n1222), .ZN(n1221) );
XOR2_X1 U952 ( .A(n1223), .B(G131), .Z(n1222) );
NAND2_X1 U953 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND2_X1 U954 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND2_X1 U955 ( .A1(n1228), .A2(G214), .ZN(n1227) );
XOR2_X1 U956 ( .A(KEYINPUT40), .B(n1229), .Z(n1224) );
NOR3_X1 U957 ( .A1(n1089), .A2(n1203), .A3(n1226), .ZN(n1229) );
INV_X1 U958 ( .A(G214), .ZN(n1203) );
NAND2_X1 U959 ( .A1(KEYINPUT2), .A2(n1230), .ZN(n1219) );
XNOR2_X1 U960 ( .A(G140), .B(n1231), .ZN(n1230) );
NAND2_X1 U961 ( .A1(KEYINPUT0), .A2(G125), .ZN(n1231) );
XNOR2_X1 U962 ( .A(G113), .B(n1232), .ZN(n1217) );
XOR2_X1 U963 ( .A(G146), .B(G122), .Z(n1232) );
INV_X1 U964 ( .A(n1174), .ZN(n1154) );
XNOR2_X1 U965 ( .A(n1233), .B(G478), .ZN(n1174) );
NAND2_X1 U966 ( .A1(n1122), .A2(n1070), .ZN(n1233) );
NAND2_X1 U967 ( .A1(n1234), .A2(n1235), .ZN(n1070) );
NAND2_X1 U968 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
XOR2_X1 U969 ( .A(n1238), .B(KEYINPUT1), .Z(n1234) );
OR2_X1 U970 ( .A1(n1237), .A2(n1236), .ZN(n1238) );
XOR2_X1 U971 ( .A(n1239), .B(n1240), .Z(n1236) );
XOR2_X1 U972 ( .A(G134), .B(G107), .Z(n1240) );
XOR2_X1 U973 ( .A(n1241), .B(n1242), .Z(n1239) );
NOR3_X1 U974 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1242) );
NOR2_X1 U975 ( .A1(KEYINPUT37), .A2(n1173), .ZN(n1245) );
NOR3_X1 U976 ( .A1(n1246), .A2(G122), .A3(n1247), .ZN(n1244) );
INV_X1 U977 ( .A(KEYINPUT37), .ZN(n1246) );
AND2_X1 U978 ( .A1(n1247), .A2(G122), .ZN(n1243) );
NAND2_X1 U979 ( .A1(KEYINPUT63), .A2(n1173), .ZN(n1247) );
NAND3_X1 U980 ( .A1(n1248), .A2(n1249), .A3(KEYINPUT19), .ZN(n1241) );
NAND2_X1 U981 ( .A1(n1250), .A2(n1226), .ZN(n1249) );
NAND2_X1 U982 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U983 ( .A1(KEYINPUT35), .A2(n1163), .ZN(n1252) );
OR2_X1 U984 ( .A1(n1253), .A2(KEYINPUT35), .ZN(n1251) );
NAND2_X1 U985 ( .A1(n1253), .A2(G143), .ZN(n1248) );
NOR2_X1 U986 ( .A1(G128), .A2(KEYINPUT30), .ZN(n1253) );
NAND3_X1 U987 ( .A1(G217), .A2(n1189), .A3(G234), .ZN(n1237) );
INV_X1 U988 ( .A(n995), .ZN(n1019) );
XNOR2_X1 U989 ( .A(n1254), .B(G472), .ZN(n995) );
NAND2_X1 U990 ( .A1(n1255), .A2(n1122), .ZN(n1254) );
XOR2_X1 U991 ( .A(n1256), .B(n1257), .Z(n1255) );
XNOR2_X1 U992 ( .A(n1097), .B(n1258), .ZN(n1257) );
NOR2_X1 U993 ( .A1(KEYINPUT59), .A2(n1259), .ZN(n1258) );
XNOR2_X1 U994 ( .A(n1095), .B(n1185), .ZN(n1259) );
INV_X1 U995 ( .A(n1093), .ZN(n1185) );
XNOR2_X1 U996 ( .A(n1260), .B(n1042), .ZN(n1093) );
XOR2_X1 U997 ( .A(G131), .B(G134), .Z(n1042) );
XNOR2_X1 U998 ( .A(G137), .B(KEYINPUT15), .ZN(n1260) );
XOR2_X1 U999 ( .A(G128), .B(n1261), .Z(n1095) );
NOR2_X1 U1000 ( .A1(KEYINPUT29), .A2(n1195), .ZN(n1261) );
XOR2_X1 U1001 ( .A(G146), .B(n1226), .Z(n1195) );
INV_X1 U1002 ( .A(G143), .ZN(n1226) );
XOR2_X1 U1003 ( .A(G113), .B(n1262), .Z(n1097) );
XNOR2_X1 U1004 ( .A(G119), .B(n1173), .ZN(n1262) );
INV_X1 U1005 ( .A(G116), .ZN(n1173) );
NAND2_X1 U1006 ( .A1(n1263), .A2(n1264), .ZN(n1256) );
NAND2_X1 U1007 ( .A1(n1087), .A2(n1265), .ZN(n1264) );
INV_X1 U1008 ( .A(n1266), .ZN(n1087) );
NAND2_X1 U1009 ( .A1(n1267), .A2(n1266), .ZN(n1263) );
NAND2_X1 U1010 ( .A1(n1090), .A2(n1268), .ZN(n1266) );
NAND2_X1 U1011 ( .A1(n1228), .A2(G210), .ZN(n1268) );
NAND2_X1 U1012 ( .A1(n1265), .A2(n1269), .ZN(n1267) );
NAND3_X1 U1013 ( .A1(G210), .A2(n1270), .A3(n1228), .ZN(n1269) );
INV_X1 U1014 ( .A(n1089), .ZN(n1228) );
NAND2_X1 U1015 ( .A1(n1189), .A2(n1271), .ZN(n1089) );
INV_X1 U1016 ( .A(G237), .ZN(n1271) );
XNOR2_X1 U1017 ( .A(KEYINPUT43), .B(n1090), .ZN(n1270) );
INV_X1 U1018 ( .A(G101), .ZN(n1090) );
INV_X1 U1019 ( .A(KEYINPUT17), .ZN(n1265) );
XNOR2_X1 U1020 ( .A(n1136), .B(KEYINPUT22), .ZN(n998) );
INV_X1 U1021 ( .A(n1000), .ZN(n1136) );
NAND2_X1 U1022 ( .A1(n1272), .A2(n1273), .ZN(n1000) );
NAND2_X1 U1023 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U1024 ( .A(n1276), .B(KEYINPUT12), .Z(n1272) );
OR2_X1 U1025 ( .A1(n1275), .A2(n1274), .ZN(n1276) );
XNOR2_X1 U1026 ( .A(n1025), .B(KEYINPUT55), .ZN(n1274) );
NAND2_X1 U1027 ( .A1(G217), .A2(n1180), .ZN(n1025) );
NAND2_X1 U1028 ( .A1(G234), .A2(n1122), .ZN(n1180) );
INV_X1 U1029 ( .A(G902), .ZN(n1122) );
INV_X1 U1030 ( .A(n1024), .ZN(n1275) );
NOR2_X1 U1031 ( .A1(n1067), .A2(G902), .ZN(n1024) );
XNOR2_X1 U1032 ( .A(n1277), .B(n1278), .ZN(n1067) );
XNOR2_X1 U1033 ( .A(n1040), .B(n1279), .ZN(n1278) );
XOR2_X1 U1034 ( .A(n1280), .B(n1281), .Z(n1279) );
AND3_X1 U1035 ( .A1(G221), .A2(n1189), .A3(G234), .ZN(n1281) );
XOR2_X1 U1036 ( .A(G953), .B(KEYINPUT36), .Z(n1189) );
NAND2_X1 U1037 ( .A1(n1282), .A2(n1283), .ZN(n1280) );
NAND2_X1 U1038 ( .A1(n1213), .A2(n1284), .ZN(n1283) );
XOR2_X1 U1039 ( .A(n1285), .B(KEYINPUT54), .Z(n1282) );
OR2_X1 U1040 ( .A1(n1284), .A2(n1213), .ZN(n1285) );
INV_X1 U1041 ( .A(n1112), .ZN(n1213) );
XOR2_X1 U1042 ( .A(G110), .B(KEYINPUT24), .Z(n1112) );
XNOR2_X1 U1043 ( .A(G119), .B(n1163), .ZN(n1284) );
INV_X1 U1044 ( .A(G128), .ZN(n1163) );
XOR2_X1 U1045 ( .A(G125), .B(G140), .Z(n1040) );
XNOR2_X1 U1046 ( .A(G137), .B(n1286), .ZN(n1277) );
XOR2_X1 U1047 ( .A(KEYINPUT57), .B(G146), .Z(n1286) );
endmodule


