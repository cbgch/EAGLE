//Key = 1110011101000000100101011011000101101100000100100110001101010011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
n1381, n1382;

XOR2_X1 U767 ( .A(G107), .B(n1051), .Z(G9) );
NOR2_X1 U768 ( .A1(n1052), .A2(n1053), .ZN(G75) );
NOR3_X1 U769 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
XOR2_X1 U770 ( .A(KEYINPUT29), .B(n1057), .Z(n1056) );
NOR2_X1 U771 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NOR2_X1 U772 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U773 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NOR2_X1 U774 ( .A1(n1064), .A2(n1065), .ZN(n1062) );
AND2_X1 U775 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR2_X1 U776 ( .A1(n1068), .A2(n1069), .ZN(n1064) );
NOR2_X1 U777 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
NOR2_X1 U778 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U779 ( .A1(n1074), .A2(n1075), .ZN(n1070) );
AND3_X1 U780 ( .A1(n1067), .A2(n1076), .A3(n1077), .ZN(n1060) );
NAND3_X1 U781 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1054) );
NAND2_X1 U782 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U783 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND3_X1 U784 ( .A1(n1085), .A2(n1067), .A3(n1086), .ZN(n1084) );
NOR3_X1 U785 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
XOR2_X1 U786 ( .A(n1063), .B(KEYINPUT14), .Z(n1089) );
NAND2_X1 U787 ( .A1(n1076), .A2(n1090), .ZN(n1083) );
NAND2_X1 U788 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U789 ( .A1(n1067), .A2(n1093), .ZN(n1092) );
NAND2_X1 U790 ( .A1(n1094), .A2(n1095), .ZN(n1091) );
NAND2_X1 U791 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
OR3_X1 U792 ( .A1(n1098), .A2(n1075), .A3(n1099), .ZN(n1097) );
NAND3_X1 U793 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1096) );
INV_X1 U794 ( .A(n1059), .ZN(n1081) );
NOR3_X1 U795 ( .A1(n1103), .A2(G953), .A3(G952), .ZN(n1052) );
INV_X1 U796 ( .A(n1078), .ZN(n1103) );
NAND4_X1 U797 ( .A1(n1104), .A2(n1076), .A3(n1105), .A4(n1106), .ZN(n1078) );
NOR3_X1 U798 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
NAND3_X1 U799 ( .A1(n1110), .A2(n1111), .A3(n1099), .ZN(n1107) );
NOR3_X1 U800 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1105) );
AND3_X1 U801 ( .A1(KEYINPUT23), .A2(n1115), .A3(G478), .ZN(n1114) );
NOR2_X1 U802 ( .A1(KEYINPUT23), .A2(G478), .ZN(n1113) );
XNOR2_X1 U803 ( .A(n1116), .B(n1117), .ZN(n1112) );
NOR2_X1 U804 ( .A1(KEYINPUT30), .A2(n1118), .ZN(n1117) );
INV_X1 U805 ( .A(G469), .ZN(n1118) );
XOR2_X1 U806 ( .A(n1119), .B(n1120), .Z(G72) );
XOR2_X1 U807 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1079), .ZN(n1122) );
AND2_X1 U809 ( .A1(G227), .A2(G900), .ZN(n1123) );
NAND2_X1 U810 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
NAND2_X1 U811 ( .A1(n1126), .A2(G953), .ZN(n1125) );
XOR2_X1 U812 ( .A(n1127), .B(n1128), .Z(n1124) );
NAND2_X1 U813 ( .A1(KEYINPUT33), .A2(n1129), .ZN(n1127) );
XOR2_X1 U814 ( .A(n1130), .B(n1131), .Z(n1129) );
XOR2_X1 U815 ( .A(KEYINPUT47), .B(G143), .Z(n1131) );
NAND2_X1 U816 ( .A1(n1079), .A2(n1132), .ZN(n1119) );
NAND3_X1 U817 ( .A1(n1133), .A2(n1134), .A3(n1135), .ZN(n1132) );
XOR2_X1 U818 ( .A(n1136), .B(KEYINPUT32), .Z(n1135) );
XNOR2_X1 U819 ( .A(KEYINPUT9), .B(n1137), .ZN(n1134) );
XOR2_X1 U820 ( .A(n1138), .B(n1139), .Z(G69) );
XOR2_X1 U821 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U822 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
NAND2_X1 U823 ( .A1(G953), .A2(n1144), .ZN(n1143) );
XOR2_X1 U824 ( .A(n1145), .B(n1146), .Z(n1142) );
NOR2_X1 U825 ( .A1(KEYINPUT51), .A2(n1147), .ZN(n1146) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
XOR2_X1 U827 ( .A(n1150), .B(KEYINPUT46), .Z(n1149) );
NAND2_X1 U828 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NOR2_X1 U829 ( .A1(n1151), .A2(n1152), .ZN(n1148) );
NAND2_X1 U830 ( .A1(n1153), .A2(n1079), .ZN(n1140) );
NOR2_X1 U831 ( .A1(n1154), .A2(n1079), .ZN(n1138) );
NOR2_X1 U832 ( .A1(n1155), .A2(n1144), .ZN(n1154) );
NOR3_X1 U833 ( .A1(n1156), .A2(n1157), .A3(n1158), .ZN(G66) );
NOR2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U835 ( .A(n1161), .B(KEYINPUT3), .Z(n1160) );
INV_X1 U836 ( .A(n1162), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1163), .A2(n1162), .ZN(n1157) );
NAND2_X1 U838 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
INV_X1 U839 ( .A(n1161), .ZN(n1163) );
NOR2_X1 U840 ( .A1(n1156), .A2(n1166), .ZN(G63) );
XOR2_X1 U841 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND3_X1 U842 ( .A1(n1164), .A2(G478), .A3(KEYINPUT6), .ZN(n1167) );
NOR2_X1 U843 ( .A1(n1156), .A2(n1169), .ZN(G60) );
XNOR2_X1 U844 ( .A(n1170), .B(n1171), .ZN(n1169) );
XNOR2_X1 U845 ( .A(n1172), .B(KEYINPUT31), .ZN(n1171) );
NAND2_X1 U846 ( .A1(KEYINPUT24), .A2(n1173), .ZN(n1172) );
NAND2_X1 U847 ( .A1(n1164), .A2(G475), .ZN(n1173) );
XOR2_X1 U848 ( .A(G104), .B(n1174), .Z(G6) );
NOR2_X1 U849 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
NOR2_X1 U850 ( .A1(KEYINPUT40), .A2(n1177), .ZN(n1176) );
INV_X1 U851 ( .A(n1178), .ZN(n1177) );
NOR2_X1 U852 ( .A1(KEYINPUT5), .A2(n1178), .ZN(n1175) );
NOR2_X1 U853 ( .A1(n1179), .A2(n1180), .ZN(G57) );
XOR2_X1 U854 ( .A(n1181), .B(n1182), .Z(n1180) );
XOR2_X1 U855 ( .A(n1183), .B(n1184), .Z(n1182) );
NAND2_X1 U856 ( .A1(n1164), .A2(G472), .ZN(n1184) );
NAND3_X1 U857 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1183) );
OR2_X1 U858 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NAND3_X1 U859 ( .A1(n1189), .A2(n1188), .A3(KEYINPUT34), .ZN(n1186) );
NOR2_X1 U860 ( .A1(KEYINPUT41), .A2(n1190), .ZN(n1189) );
NAND2_X1 U861 ( .A1(n1190), .A2(n1191), .ZN(n1185) );
INV_X1 U862 ( .A(KEYINPUT34), .ZN(n1191) );
XOR2_X1 U863 ( .A(n1192), .B(n1193), .Z(n1190) );
NAND2_X1 U864 ( .A1(KEYINPUT19), .A2(n1194), .ZN(n1192) );
XOR2_X1 U865 ( .A(G134), .B(n1195), .Z(n1194) );
NOR2_X1 U866 ( .A1(G952), .A2(n1196), .ZN(n1179) );
XOR2_X1 U867 ( .A(KEYINPUT59), .B(G953), .Z(n1196) );
NOR2_X1 U868 ( .A1(n1156), .A2(n1197), .ZN(G54) );
XOR2_X1 U869 ( .A(n1198), .B(n1199), .Z(n1197) );
NAND2_X1 U870 ( .A1(n1164), .A2(G469), .ZN(n1198) );
NOR2_X1 U871 ( .A1(n1156), .A2(n1200), .ZN(G51) );
XOR2_X1 U872 ( .A(n1201), .B(n1202), .Z(n1200) );
XOR2_X1 U873 ( .A(n1203), .B(n1204), .Z(n1202) );
NAND2_X1 U874 ( .A1(n1164), .A2(n1205), .ZN(n1203) );
AND2_X1 U875 ( .A1(G902), .A2(n1055), .ZN(n1164) );
NAND4_X1 U876 ( .A1(n1206), .A2(n1133), .A3(n1137), .A4(n1136), .ZN(n1055) );
AND4_X1 U877 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1133) );
NOR3_X1 U878 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1210) );
INV_X1 U879 ( .A(n1214), .ZN(n1213) );
NOR3_X1 U880 ( .A1(n1215), .A2(n1216), .A3(n1217), .ZN(n1211) );
XOR2_X1 U881 ( .A(KEYINPUT50), .B(n1076), .Z(n1215) );
INV_X1 U882 ( .A(n1153), .ZN(n1206) );
NAND4_X1 U883 ( .A1(n1218), .A2(n1178), .A3(n1219), .A4(n1220), .ZN(n1153) );
NOR4_X1 U884 ( .A1(n1051), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1220) );
AND2_X1 U885 ( .A1(n1093), .A2(n1224), .ZN(n1051) );
NAND2_X1 U886 ( .A1(n1225), .A2(n1226), .ZN(n1219) );
NAND2_X1 U887 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
NAND2_X1 U888 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
INV_X1 U889 ( .A(KEYINPUT13), .ZN(n1230) );
NAND2_X1 U890 ( .A1(n1102), .A2(n1231), .ZN(n1227) );
NAND2_X1 U891 ( .A1(n1232), .A2(n1233), .ZN(n1231) );
NAND2_X1 U892 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U893 ( .A1(n1077), .A2(n1236), .ZN(n1232) );
NAND2_X1 U894 ( .A1(n1077), .A2(n1224), .ZN(n1178) );
AND3_X1 U895 ( .A1(n1235), .A2(n1237), .A3(n1225), .ZN(n1224) );
INV_X1 U896 ( .A(n1075), .ZN(n1235) );
NAND3_X1 U897 ( .A1(n1066), .A2(n1238), .A3(KEYINPUT13), .ZN(n1218) );
NAND2_X1 U898 ( .A1(n1229), .A2(n1239), .ZN(n1238) );
XOR2_X1 U899 ( .A(n1240), .B(n1241), .Z(n1201) );
NAND2_X1 U900 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
NAND2_X1 U901 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
XOR2_X1 U902 ( .A(n1246), .B(KEYINPUT22), .Z(n1242) );
OR2_X1 U903 ( .A1(n1245), .A2(n1244), .ZN(n1246) );
NOR2_X1 U904 ( .A1(n1079), .A2(G952), .ZN(n1156) );
XNOR2_X1 U905 ( .A(G146), .B(n1137), .ZN(G48) );
NAND3_X1 U906 ( .A1(n1077), .A2(n1066), .A3(n1247), .ZN(n1137) );
XOR2_X1 U907 ( .A(n1248), .B(n1214), .Z(G45) );
NAND3_X1 U908 ( .A1(n1249), .A2(n1066), .A3(n1234), .ZN(n1214) );
XOR2_X1 U909 ( .A(G140), .B(n1212), .Z(G42) );
AND3_X1 U910 ( .A1(n1076), .A2(n1237), .A3(n1250), .ZN(n1212) );
XNOR2_X1 U911 ( .A(G137), .B(n1208), .ZN(G39) );
NAND3_X1 U912 ( .A1(n1247), .A2(n1076), .A3(n1094), .ZN(n1208) );
XOR2_X1 U913 ( .A(G134), .B(n1251), .Z(G36) );
NOR3_X1 U914 ( .A1(n1217), .A2(n1216), .A3(n1069), .ZN(n1251) );
INV_X1 U915 ( .A(n1093), .ZN(n1216) );
XNOR2_X1 U916 ( .A(G131), .B(n1136), .ZN(G33) );
NAND3_X1 U917 ( .A1(n1249), .A2(n1076), .A3(n1077), .ZN(n1136) );
INV_X1 U918 ( .A(n1069), .ZN(n1076) );
NAND2_X1 U919 ( .A1(n1085), .A2(n1252), .ZN(n1069) );
NAND2_X1 U920 ( .A1(G214), .A2(n1253), .ZN(n1252) );
INV_X1 U921 ( .A(n1217), .ZN(n1249) );
NAND3_X1 U922 ( .A1(n1237), .A2(n1254), .A3(n1236), .ZN(n1217) );
NAND3_X1 U923 ( .A1(n1255), .A2(n1256), .A3(n1257), .ZN(G30) );
OR2_X1 U924 ( .A1(n1209), .A2(G128), .ZN(n1257) );
NAND2_X1 U925 ( .A1(KEYINPUT58), .A2(n1258), .ZN(n1256) );
NAND2_X1 U926 ( .A1(G128), .A2(n1259), .ZN(n1258) );
XNOR2_X1 U927 ( .A(KEYINPUT1), .B(n1209), .ZN(n1259) );
NAND2_X1 U928 ( .A1(n1260), .A2(n1261), .ZN(n1255) );
INV_X1 U929 ( .A(KEYINPUT58), .ZN(n1261) );
NAND2_X1 U930 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
NAND3_X1 U931 ( .A1(KEYINPUT1), .A2(G128), .A3(n1209), .ZN(n1263) );
OR2_X1 U932 ( .A1(n1209), .A2(KEYINPUT1), .ZN(n1262) );
NAND3_X1 U933 ( .A1(n1093), .A2(n1066), .A3(n1247), .ZN(n1209) );
AND4_X1 U934 ( .A1(n1237), .A2(n1101), .A3(n1264), .A4(n1254), .ZN(n1247) );
XOR2_X1 U935 ( .A(n1265), .B(n1266), .Z(G3) );
XOR2_X1 U936 ( .A(KEYINPUT2), .B(G101), .Z(n1266) );
NAND3_X1 U937 ( .A1(n1229), .A2(n1066), .A3(n1267), .ZN(n1265) );
XOR2_X1 U938 ( .A(n1239), .B(KEYINPUT12), .Z(n1267) );
NOR3_X1 U939 ( .A1(n1072), .A2(n1074), .A3(n1063), .ZN(n1229) );
INV_X1 U940 ( .A(n1094), .ZN(n1063) );
XNOR2_X1 U941 ( .A(G125), .B(n1268), .ZN(G27) );
NAND2_X1 U942 ( .A1(KEYINPUT43), .A2(n1269), .ZN(n1268) );
INV_X1 U943 ( .A(n1207), .ZN(n1269) );
NAND3_X1 U944 ( .A1(n1102), .A2(n1066), .A3(n1250), .ZN(n1207) );
AND4_X1 U945 ( .A1(n1077), .A2(n1100), .A3(n1101), .A4(n1254), .ZN(n1250) );
NAND2_X1 U946 ( .A1(n1270), .A2(n1271), .ZN(n1254) );
NAND4_X1 U947 ( .A1(n1126), .A2(G953), .A3(G902), .A4(n1272), .ZN(n1271) );
XNOR2_X1 U948 ( .A(G900), .B(KEYINPUT61), .ZN(n1126) );
XOR2_X1 U949 ( .A(n1059), .B(KEYINPUT4), .Z(n1270) );
XNOR2_X1 U950 ( .A(G122), .B(n1273), .ZN(G24) );
NAND3_X1 U951 ( .A1(n1225), .A2(n1274), .A3(n1067), .ZN(n1273) );
NOR2_X1 U952 ( .A1(n1073), .A2(n1075), .ZN(n1067) );
NAND2_X1 U953 ( .A1(n1100), .A2(n1104), .ZN(n1075) );
XOR2_X1 U954 ( .A(KEYINPUT17), .B(n1234), .Z(n1274) );
AND2_X1 U955 ( .A1(n1109), .A2(n1275), .ZN(n1234) );
XOR2_X1 U956 ( .A(n1276), .B(n1223), .Z(G21) );
AND3_X1 U957 ( .A1(n1277), .A2(n1264), .A3(n1102), .ZN(n1223) );
XNOR2_X1 U958 ( .A(G119), .B(KEYINPUT21), .ZN(n1276) );
XNOR2_X1 U959 ( .A(n1222), .B(n1278), .ZN(G18) );
NOR2_X1 U960 ( .A1(G116), .A2(KEYINPUT38), .ZN(n1278) );
AND4_X1 U961 ( .A1(n1102), .A2(n1236), .A3(n1093), .A4(n1225), .ZN(n1222) );
NOR2_X1 U962 ( .A1(n1109), .A2(n1279), .ZN(n1093) );
XNOR2_X1 U963 ( .A(G113), .B(n1280), .ZN(G15) );
NAND4_X1 U964 ( .A1(n1077), .A2(n1236), .A3(n1225), .A4(n1281), .ZN(n1280) );
XOR2_X1 U965 ( .A(KEYINPUT60), .B(n1102), .Z(n1281) );
INV_X1 U966 ( .A(n1073), .ZN(n1102) );
NAND2_X1 U967 ( .A1(n1282), .A2(n1099), .ZN(n1073) );
INV_X1 U968 ( .A(n1072), .ZN(n1236) );
NAND2_X1 U969 ( .A1(n1104), .A2(n1264), .ZN(n1072) );
AND2_X1 U970 ( .A1(n1279), .A2(n1109), .ZN(n1077) );
INV_X1 U971 ( .A(n1275), .ZN(n1279) );
XOR2_X1 U972 ( .A(G110), .B(n1221), .Z(G12) );
AND3_X1 U973 ( .A1(n1237), .A2(n1100), .A3(n1277), .ZN(n1221) );
AND3_X1 U974 ( .A1(n1225), .A2(n1101), .A3(n1094), .ZN(n1277) );
NOR2_X1 U975 ( .A1(n1275), .A2(n1109), .ZN(n1094) );
XNOR2_X1 U976 ( .A(n1283), .B(G475), .ZN(n1109) );
NAND2_X1 U977 ( .A1(n1170), .A2(n1284), .ZN(n1283) );
XNOR2_X1 U978 ( .A(n1285), .B(n1286), .ZN(n1170) );
XOR2_X1 U979 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U980 ( .A(n1289), .B(G113), .Z(n1288) );
NAND2_X1 U981 ( .A1(KEYINPUT49), .A2(G146), .ZN(n1289) );
XNOR2_X1 U982 ( .A(G131), .B(KEYINPUT20), .ZN(n1287) );
XOR2_X1 U983 ( .A(n1290), .B(n1291), .Z(n1285) );
XNOR2_X1 U984 ( .A(n1292), .B(n1293), .ZN(n1291) );
NAND2_X1 U985 ( .A1(G214), .A2(n1294), .ZN(n1292) );
XNOR2_X1 U986 ( .A(n1128), .B(n1295), .ZN(n1290) );
NAND2_X1 U987 ( .A1(n1110), .A2(n1296), .ZN(n1275) );
NAND2_X1 U988 ( .A1(G478), .A2(n1115), .ZN(n1296) );
OR2_X1 U989 ( .A1(n1115), .A2(G478), .ZN(n1110) );
NAND2_X1 U990 ( .A1(n1168), .A2(n1284), .ZN(n1115) );
XOR2_X1 U991 ( .A(n1297), .B(n1298), .Z(n1168) );
XOR2_X1 U992 ( .A(G107), .B(n1299), .Z(n1298) );
XOR2_X1 U993 ( .A(G143), .B(G116), .Z(n1299) );
XOR2_X1 U994 ( .A(n1300), .B(n1295), .Z(n1297) );
XOR2_X1 U995 ( .A(n1301), .B(n1302), .Z(n1300) );
NAND2_X1 U996 ( .A1(G217), .A2(n1303), .ZN(n1301) );
INV_X1 U997 ( .A(n1104), .ZN(n1101) );
XOR2_X1 U998 ( .A(n1304), .B(n1165), .Z(n1104) );
AND2_X1 U999 ( .A1(G217), .A2(n1305), .ZN(n1165) );
NAND2_X1 U1000 ( .A1(n1161), .A2(n1284), .ZN(n1304) );
XOR2_X1 U1001 ( .A(n1306), .B(n1307), .Z(n1161) );
XOR2_X1 U1002 ( .A(n1308), .B(n1128), .Z(n1307) );
XOR2_X1 U1003 ( .A(G125), .B(n1309), .Z(n1128) );
XOR2_X1 U1004 ( .A(n1310), .B(n1311), .Z(n1306) );
AND2_X1 U1005 ( .A1(n1303), .A2(G221), .ZN(n1311) );
AND2_X1 U1006 ( .A1(G234), .A2(n1079), .ZN(n1303) );
XOR2_X1 U1007 ( .A(n1312), .B(G146), .Z(n1310) );
NAND3_X1 U1008 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1312) );
NAND2_X1 U1009 ( .A1(KEYINPUT45), .A2(n1316), .ZN(n1315) );
NAND3_X1 U1010 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(n1314) );
INV_X1 U1011 ( .A(KEYINPUT45), .ZN(n1318) );
OR2_X1 U1012 ( .A1(n1319), .A2(n1317), .ZN(n1313) );
NOR2_X1 U1013 ( .A1(KEYINPUT53), .A2(n1316), .ZN(n1317) );
XOR2_X1 U1014 ( .A(G128), .B(n1320), .Z(n1316) );
NOR2_X1 U1015 ( .A1(G119), .A2(KEYINPUT48), .ZN(n1320) );
AND2_X1 U1016 ( .A1(n1066), .A2(n1239), .ZN(n1225) );
NAND2_X1 U1017 ( .A1(n1059), .A2(n1321), .ZN(n1239) );
NAND4_X1 U1018 ( .A1(G953), .A2(G902), .A3(n1272), .A4(n1144), .ZN(n1321) );
INV_X1 U1019 ( .A(G898), .ZN(n1144) );
NAND3_X1 U1020 ( .A1(n1272), .A2(n1079), .A3(G952), .ZN(n1059) );
NAND2_X1 U1021 ( .A1(G237), .A2(G234), .ZN(n1272) );
NOR2_X1 U1022 ( .A1(n1085), .A2(n1322), .ZN(n1066) );
NOR2_X1 U1023 ( .A1(n1087), .A2(n1088), .ZN(n1322) );
INV_X1 U1024 ( .A(G214), .ZN(n1087) );
XOR2_X1 U1025 ( .A(n1323), .B(n1205), .Z(n1085) );
AND2_X1 U1026 ( .A1(G210), .A2(n1253), .ZN(n1205) );
INV_X1 U1027 ( .A(n1088), .ZN(n1253) );
NOR2_X1 U1028 ( .A1(n1324), .A2(G237), .ZN(n1088) );
XOR2_X1 U1029 ( .A(KEYINPUT28), .B(G902), .Z(n1324) );
NAND4_X1 U1030 ( .A1(n1325), .A2(n1284), .A3(n1326), .A4(n1327), .ZN(n1323) );
NAND2_X1 U1031 ( .A1(n1328), .A2(n1329), .ZN(n1327) );
INV_X1 U1032 ( .A(KEYINPUT27), .ZN(n1329) );
NAND2_X1 U1033 ( .A1(n1330), .A2(n1331), .ZN(n1328) );
INV_X1 U1034 ( .A(n1204), .ZN(n1331) );
XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n1332), .ZN(n1330) );
NAND2_X1 U1036 ( .A1(KEYINPUT27), .A2(n1333), .ZN(n1326) );
NAND2_X1 U1037 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
OR3_X1 U1038 ( .A1(n1332), .A2(n1204), .A3(KEYINPUT52), .ZN(n1335) );
NAND2_X1 U1039 ( .A1(KEYINPUT52), .A2(n1332), .ZN(n1334) );
NAND2_X1 U1040 ( .A1(n1204), .A2(n1332), .ZN(n1325) );
XNOR2_X1 U1041 ( .A(n1244), .B(n1336), .ZN(n1332) );
XOR2_X1 U1042 ( .A(n1241), .B(n1245), .Z(n1336) );
INV_X1 U1043 ( .A(n1193), .ZN(n1245) );
XOR2_X1 U1044 ( .A(n1337), .B(n1338), .Z(n1193) );
NOR2_X1 U1045 ( .A1(n1155), .A2(G953), .ZN(n1241) );
INV_X1 U1046 ( .A(G224), .ZN(n1155) );
XOR2_X1 U1047 ( .A(G125), .B(KEYINPUT39), .Z(n1244) );
XOR2_X1 U1048 ( .A(n1339), .B(n1340), .Z(n1204) );
INV_X1 U1049 ( .A(n1145), .ZN(n1340) );
XOR2_X1 U1050 ( .A(n1341), .B(n1342), .Z(n1145) );
XOR2_X1 U1051 ( .A(n1319), .B(n1295), .Z(n1342) );
XOR2_X1 U1052 ( .A(G122), .B(KEYINPUT7), .Z(n1295) );
XNOR2_X1 U1053 ( .A(KEYINPUT44), .B(KEYINPUT36), .ZN(n1341) );
XNOR2_X1 U1054 ( .A(n1152), .B(n1151), .ZN(n1339) );
AND2_X1 U1055 ( .A1(n1343), .A2(n1344), .ZN(n1151) );
NAND2_X1 U1056 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XNOR2_X1 U1057 ( .A(n1347), .B(KEYINPUT35), .ZN(n1346) );
XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(G113), .ZN(n1345) );
XOR2_X1 U1059 ( .A(n1348), .B(KEYINPUT8), .Z(n1343) );
NAND2_X1 U1060 ( .A1(n1349), .A2(n1347), .ZN(n1348) );
XOR2_X1 U1061 ( .A(G116), .B(n1350), .Z(n1347) );
NOR2_X1 U1062 ( .A1(G119), .A2(KEYINPUT25), .ZN(n1350) );
XOR2_X1 U1063 ( .A(KEYINPUT54), .B(G113), .Z(n1349) );
XNOR2_X1 U1064 ( .A(n1351), .B(G101), .ZN(n1152) );
NAND3_X1 U1065 ( .A1(n1352), .A2(n1353), .A3(n1354), .ZN(n1351) );
NAND2_X1 U1066 ( .A1(G107), .A2(n1355), .ZN(n1354) );
NAND2_X1 U1067 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
INV_X1 U1068 ( .A(n1358), .ZN(n1356) );
NAND3_X1 U1069 ( .A1(n1357), .A2(n1358), .A3(n1359), .ZN(n1353) );
XOR2_X1 U1070 ( .A(n1360), .B(G107), .Z(n1358) );
XNOR2_X1 U1071 ( .A(KEYINPUT18), .B(KEYINPUT11), .ZN(n1360) );
OR2_X1 U1072 ( .A1(n1359), .A2(n1357), .ZN(n1352) );
XOR2_X1 U1073 ( .A(G104), .B(KEYINPUT62), .Z(n1357) );
INV_X1 U1074 ( .A(KEYINPUT15), .ZN(n1359) );
INV_X1 U1075 ( .A(n1264), .ZN(n1100) );
NAND2_X1 U1076 ( .A1(n1361), .A2(n1111), .ZN(n1264) );
NAND3_X1 U1077 ( .A1(n1362), .A2(n1284), .A3(n1363), .ZN(n1111) );
INV_X1 U1078 ( .A(G472), .ZN(n1362) );
XNOR2_X1 U1079 ( .A(n1108), .B(KEYINPUT56), .ZN(n1361) );
AND2_X1 U1080 ( .A1(G472), .A2(n1364), .ZN(n1108) );
NAND2_X1 U1081 ( .A1(n1363), .A2(n1284), .ZN(n1364) );
XNOR2_X1 U1082 ( .A(n1365), .B(n1366), .ZN(n1363) );
XNOR2_X1 U1083 ( .A(n1181), .B(n1188), .ZN(n1366) );
XNOR2_X1 U1084 ( .A(G113), .B(n1367), .ZN(n1188) );
NOR2_X1 U1085 ( .A1(KEYINPUT10), .A2(n1368), .ZN(n1367) );
XOR2_X1 U1086 ( .A(G119), .B(G116), .Z(n1368) );
XNOR2_X1 U1087 ( .A(n1369), .B(G101), .ZN(n1181) );
NAND2_X1 U1088 ( .A1(G210), .A2(n1294), .ZN(n1369) );
NOR2_X1 U1089 ( .A1(G953), .A2(G237), .ZN(n1294) );
XOR2_X1 U1090 ( .A(n1370), .B(n1338), .Z(n1365) );
XNOR2_X1 U1091 ( .A(n1371), .B(KEYINPUT16), .ZN(n1338) );
NAND2_X1 U1092 ( .A1(n1372), .A2(KEYINPUT63), .ZN(n1371) );
XOR2_X1 U1093 ( .A(n1373), .B(G146), .Z(n1372) );
NAND2_X1 U1094 ( .A1(KEYINPUT37), .A2(n1248), .ZN(n1373) );
INV_X1 U1095 ( .A(G143), .ZN(n1248) );
XNOR2_X1 U1096 ( .A(n1374), .B(KEYINPUT55), .ZN(n1370) );
INV_X1 U1097 ( .A(n1074), .ZN(n1237) );
NAND2_X1 U1098 ( .A1(n1375), .A2(n1099), .ZN(n1074) );
NAND2_X1 U1099 ( .A1(G221), .A2(n1305), .ZN(n1099) );
NAND2_X1 U1100 ( .A1(n1376), .A2(G234), .ZN(n1305) );
XOR2_X1 U1101 ( .A(KEYINPUT28), .B(n1284), .Z(n1376) );
XOR2_X1 U1102 ( .A(KEYINPUT42), .B(n1098), .Z(n1375) );
INV_X1 U1103 ( .A(n1282), .ZN(n1098) );
XOR2_X1 U1104 ( .A(n1116), .B(G469), .Z(n1282) );
NAND2_X1 U1105 ( .A1(n1199), .A2(n1284), .ZN(n1116) );
INV_X1 U1106 ( .A(G902), .ZN(n1284) );
XOR2_X1 U1107 ( .A(n1377), .B(n1378), .Z(n1199) );
XOR2_X1 U1108 ( .A(n1379), .B(n1380), .Z(n1378) );
XOR2_X1 U1109 ( .A(n1381), .B(n1319), .Z(n1380) );
XOR2_X1 U1110 ( .A(G110), .B(KEYINPUT26), .Z(n1319) );
AND2_X1 U1111 ( .A1(n1079), .A2(G227), .ZN(n1381) );
INV_X1 U1112 ( .A(G953), .ZN(n1079) );
XOR2_X1 U1113 ( .A(G107), .B(G101), .Z(n1379) );
XOR2_X1 U1114 ( .A(n1382), .B(n1293), .Z(n1377) );
XOR2_X1 U1115 ( .A(G104), .B(G143), .Z(n1293) );
XNOR2_X1 U1116 ( .A(n1130), .B(n1309), .ZN(n1382) );
XOR2_X1 U1117 ( .A(G140), .B(KEYINPUT0), .Z(n1309) );
XOR2_X1 U1118 ( .A(G146), .B(n1374), .Z(n1130) );
XOR2_X1 U1119 ( .A(n1195), .B(n1302), .Z(n1374) );
XNOR2_X1 U1120 ( .A(G134), .B(n1337), .ZN(n1302) );
INV_X1 U1121 ( .A(G128), .ZN(n1337) );
XOR2_X1 U1122 ( .A(G131), .B(n1308), .Z(n1195) );
XOR2_X1 U1123 ( .A(G137), .B(KEYINPUT57), .Z(n1308) );
endmodule


