//Key = 1000100110011010101111000010110001111010110110001001101111001101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
n1467, n1468, n1469, n1470;

NAND3_X1 U797 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(G9) );
NAND2_X1 U798 ( .A1(G107), .A2(n1110), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U800 ( .A(KEYINPUT46), .ZN(n1112) );
XNOR2_X1 U801 ( .A(KEYINPUT24), .B(n1113), .ZN(n1111) );
OR3_X1 U802 ( .A1(n1113), .A2(G107), .A3(KEYINPUT46), .ZN(n1108) );
NAND2_X1 U803 ( .A1(KEYINPUT46), .A2(n1113), .ZN(n1107) );
NOR2_X1 U804 ( .A1(n1114), .A2(n1115), .ZN(G75) );
NOR3_X1 U805 ( .A1(n1116), .A2(G953), .A3(n1117), .ZN(n1115) );
XOR2_X1 U806 ( .A(KEYINPUT16), .B(n1118), .Z(n1116) );
NOR4_X1 U807 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
NOR2_X1 U808 ( .A1(n1123), .A2(n1124), .ZN(n1121) );
NOR2_X1 U809 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
AND2_X1 U810 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
NOR2_X1 U811 ( .A1(n1129), .A2(n1130), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(n1120) );
NOR2_X1 U815 ( .A1(n1137), .A2(n1138), .ZN(n1135) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1124), .ZN(n1138) );
NAND3_X1 U817 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1124) );
INV_X1 U818 ( .A(n1143), .ZN(n1142) );
NOR3_X1 U819 ( .A1(n1143), .A2(n1144), .A3(n1130), .ZN(n1137) );
NOR2_X1 U820 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
AND2_X1 U821 ( .A1(n1147), .A2(n1141), .ZN(n1146) );
AND2_X1 U822 ( .A1(n1140), .A2(n1148), .ZN(n1145) );
NOR4_X1 U823 ( .A1(n1149), .A2(n1143), .A3(n1150), .A4(n1151), .ZN(n1119) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XNOR2_X1 U825 ( .A(n1154), .B(KEYINPUT63), .ZN(n1153) );
NOR2_X1 U826 ( .A1(n1141), .A2(n1155), .ZN(n1150) );
OR3_X1 U827 ( .A1(n1156), .A2(n1136), .A3(n1130), .ZN(n1149) );
NOR3_X1 U828 ( .A1(n1117), .A2(G953), .A3(G952), .ZN(n1114) );
AND4_X1 U829 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1117) );
NOR4_X1 U830 ( .A1(n1161), .A2(n1152), .A3(n1162), .A4(n1163), .ZN(n1160) );
XNOR2_X1 U831 ( .A(n1164), .B(KEYINPUT18), .ZN(n1163) );
NOR2_X1 U832 ( .A1(n1165), .A2(n1166), .ZN(n1162) );
XOR2_X1 U833 ( .A(KEYINPUT52), .B(n1167), .Z(n1166) );
INV_X1 U834 ( .A(n1168), .ZN(n1165) );
NOR3_X1 U835 ( .A1(n1136), .A2(n1169), .A3(n1170), .ZN(n1159) );
NOR2_X1 U836 ( .A1(G475), .A2(n1171), .ZN(n1170) );
XNOR2_X1 U837 ( .A(n1172), .B(n1173), .ZN(n1171) );
XNOR2_X1 U838 ( .A(KEYINPUT27), .B(KEYINPUT19), .ZN(n1173) );
NOR2_X1 U839 ( .A1(n1172), .A2(n1174), .ZN(n1169) );
XOR2_X1 U840 ( .A(n1175), .B(n1176), .Z(n1158) );
XNOR2_X1 U841 ( .A(n1177), .B(KEYINPUT48), .ZN(n1176) );
INV_X1 U842 ( .A(n1178), .ZN(n1177) );
NAND2_X1 U843 ( .A1(KEYINPUT54), .A2(n1179), .ZN(n1175) );
XOR2_X1 U844 ( .A(n1180), .B(n1181), .Z(G72) );
NOR2_X1 U845 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NOR2_X1 U846 ( .A1(n1184), .A2(n1185), .ZN(n1182) );
NAND2_X1 U847 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
NAND2_X1 U848 ( .A1(n1188), .A2(n1183), .ZN(n1187) );
XNOR2_X1 U849 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND3_X1 U850 ( .A1(G900), .A2(n1190), .A3(G953), .ZN(n1186) );
XNOR2_X1 U851 ( .A(n1191), .B(n1192), .ZN(n1190) );
XNOR2_X1 U852 ( .A(n1193), .B(n1194), .ZN(n1192) );
NOR2_X1 U853 ( .A1(n1195), .A2(n1196), .ZN(n1194) );
XOR2_X1 U854 ( .A(n1197), .B(KEYINPUT29), .Z(n1196) );
NAND2_X1 U855 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
XNOR2_X1 U856 ( .A(KEYINPUT37), .B(n1200), .ZN(n1198) );
XOR2_X1 U857 ( .A(n1201), .B(n1202), .Z(n1191) );
NAND3_X1 U858 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1201) );
NAND2_X1 U859 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND2_X1 U860 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
XNOR2_X1 U861 ( .A(KEYINPUT31), .B(n1210), .ZN(n1208) );
NAND3_X1 U862 ( .A1(G125), .A2(n1211), .A3(n1209), .ZN(n1204) );
INV_X1 U863 ( .A(KEYINPUT49), .ZN(n1209) );
NAND2_X1 U864 ( .A1(KEYINPUT49), .A2(n1210), .ZN(n1203) );
NAND2_X1 U865 ( .A1(n1212), .A2(n1213), .ZN(G69) );
NAND2_X1 U866 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U867 ( .A(KEYINPUT7), .B(n1216), .Z(n1212) );
NOR2_X1 U868 ( .A1(n1214), .A2(n1217), .ZN(n1216) );
NOR2_X1 U869 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
INV_X1 U870 ( .A(n1215), .ZN(n1219) );
NAND3_X1 U871 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1215) );
NAND2_X1 U872 ( .A1(G953), .A2(n1223), .ZN(n1221) );
NAND2_X1 U873 ( .A1(n1224), .A2(n1183), .ZN(n1220) );
NOR3_X1 U874 ( .A1(n1222), .A2(G953), .A3(n1225), .ZN(n1218) );
XNOR2_X1 U875 ( .A(n1226), .B(n1227), .ZN(n1222) );
NAND2_X1 U876 ( .A1(n1228), .A2(n1229), .ZN(n1226) );
NAND2_X1 U877 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
XOR2_X1 U878 ( .A(KEYINPUT14), .B(n1232), .Z(n1228) );
NOR2_X1 U879 ( .A1(n1231), .A2(n1230), .ZN(n1232) );
AND2_X1 U880 ( .A1(G953), .A2(n1233), .ZN(n1214) );
NAND2_X1 U881 ( .A1(G898), .A2(G224), .ZN(n1233) );
NOR2_X1 U882 ( .A1(n1234), .A2(n1235), .ZN(G66) );
XOR2_X1 U883 ( .A(KEYINPUT59), .B(n1236), .Z(n1235) );
NOR3_X1 U884 ( .A1(n1167), .A2(n1237), .A3(n1238), .ZN(n1234) );
NOR3_X1 U885 ( .A1(n1239), .A2(n1168), .A3(n1240), .ZN(n1238) );
INV_X1 U886 ( .A(n1241), .ZN(n1239) );
NOR2_X1 U887 ( .A1(n1242), .A2(n1241), .ZN(n1237) );
NOR2_X1 U888 ( .A1(n1243), .A2(n1168), .ZN(n1242) );
NOR2_X1 U889 ( .A1(n1236), .A2(n1244), .ZN(G63) );
NOR2_X1 U890 ( .A1(n1245), .A2(n1246), .ZN(n1244) );
XOR2_X1 U891 ( .A(n1247), .B(n1248), .Z(n1246) );
NOR2_X1 U892 ( .A1(n1249), .A2(n1240), .ZN(n1248) );
INV_X1 U893 ( .A(G478), .ZN(n1249) );
NOR2_X1 U894 ( .A1(n1250), .A2(KEYINPUT6), .ZN(n1247) );
AND2_X1 U895 ( .A1(n1250), .A2(KEYINPUT6), .ZN(n1245) );
NOR2_X1 U896 ( .A1(n1236), .A2(n1251), .ZN(G60) );
NOR3_X1 U897 ( .A1(n1172), .A2(n1252), .A3(n1253), .ZN(n1251) );
NOR2_X1 U898 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NOR2_X1 U899 ( .A1(n1243), .A2(n1174), .ZN(n1254) );
INV_X1 U900 ( .A(n1122), .ZN(n1243) );
NOR3_X1 U901 ( .A1(n1256), .A2(n1174), .A3(n1240), .ZN(n1252) );
INV_X1 U902 ( .A(G475), .ZN(n1174) );
INV_X1 U903 ( .A(n1255), .ZN(n1256) );
XNOR2_X1 U904 ( .A(G104), .B(n1257), .ZN(G6) );
NOR2_X1 U905 ( .A1(n1236), .A2(n1258), .ZN(G57) );
XOR2_X1 U906 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U907 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U908 ( .A(n1263), .B(n1264), .Z(n1259) );
NOR2_X1 U909 ( .A1(n1265), .A2(n1240), .ZN(n1264) );
NAND2_X1 U910 ( .A1(n1266), .A2(n1267), .ZN(n1263) );
XOR2_X1 U911 ( .A(n1268), .B(KEYINPUT39), .Z(n1266) );
NOR2_X1 U912 ( .A1(n1236), .A2(n1269), .ZN(G54) );
XOR2_X1 U913 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U914 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U915 ( .A(KEYINPUT57), .B(n1274), .Z(n1270) );
NOR2_X1 U916 ( .A1(n1275), .A2(n1240), .ZN(n1274) );
NOR2_X1 U917 ( .A1(n1236), .A2(n1276), .ZN(G51) );
XOR2_X1 U918 ( .A(n1277), .B(n1278), .Z(n1276) );
XNOR2_X1 U919 ( .A(n1279), .B(n1280), .ZN(n1278) );
NAND3_X1 U920 ( .A1(n1281), .A2(n1282), .A3(n1283), .ZN(n1279) );
NAND2_X1 U921 ( .A1(n1284), .A2(n1210), .ZN(n1283) );
NAND2_X1 U922 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
XNOR2_X1 U923 ( .A(KEYINPUT3), .B(n1287), .ZN(n1285) );
NAND3_X1 U924 ( .A1(n1287), .A2(n1288), .A3(n1289), .ZN(n1282) );
INV_X1 U925 ( .A(KEYINPUT60), .ZN(n1289) );
NAND2_X1 U926 ( .A1(KEYINPUT3), .A2(n1290), .ZN(n1288) );
NAND3_X1 U927 ( .A1(n1291), .A2(n1292), .A3(KEYINPUT60), .ZN(n1281) );
NAND2_X1 U928 ( .A1(n1293), .A2(n1290), .ZN(n1292) );
NAND2_X1 U929 ( .A1(G125), .A2(n1286), .ZN(n1290) );
INV_X1 U930 ( .A(KEYINPUT45), .ZN(n1286) );
INV_X1 U931 ( .A(KEYINPUT3), .ZN(n1293) );
XOR2_X1 U932 ( .A(n1294), .B(n1295), .Z(n1277) );
NOR2_X1 U933 ( .A1(n1240), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U934 ( .A(KEYINPUT44), .B(n1178), .ZN(n1296) );
NAND2_X1 U935 ( .A1(G902), .A2(n1122), .ZN(n1240) );
NAND3_X1 U936 ( .A1(n1297), .A2(n1298), .A3(n1189), .ZN(n1122) );
AND2_X1 U937 ( .A1(n1299), .A2(n1300), .ZN(n1189) );
AND4_X1 U938 ( .A1(n1301), .A2(n1302), .A3(n1303), .A4(n1304), .ZN(n1300) );
NOR4_X1 U939 ( .A1(n1305), .A2(n1306), .A3(n1307), .A4(n1308), .ZN(n1299) );
NOR2_X1 U940 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
INV_X1 U941 ( .A(n1311), .ZN(n1306) );
INV_X1 U942 ( .A(n1312), .ZN(n1305) );
NAND2_X1 U943 ( .A1(KEYINPUT62), .A2(n1313), .ZN(n1298) );
OR2_X1 U944 ( .A1(n1225), .A2(KEYINPUT62), .ZN(n1297) );
INV_X1 U945 ( .A(n1224), .ZN(n1225) );
NAND2_X1 U946 ( .A1(n1314), .A2(n1315), .ZN(n1224) );
AND4_X1 U947 ( .A1(n1113), .A2(n1313), .A3(n1316), .A4(n1317), .ZN(n1315) );
NAND3_X1 U948 ( .A1(n1141), .A2(n1318), .A3(n1127), .ZN(n1113) );
NOR4_X1 U949 ( .A1(n1319), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1314) );
NOR2_X1 U950 ( .A1(KEYINPUT1), .A2(n1257), .ZN(n1322) );
NAND3_X1 U951 ( .A1(n1141), .A2(n1318), .A3(n1323), .ZN(n1257) );
NOR4_X1 U952 ( .A1(n1324), .A2(n1325), .A3(n1326), .A4(n1327), .ZN(n1321) );
NOR2_X1 U953 ( .A1(n1328), .A2(n1329), .ZN(n1325) );
NOR2_X1 U954 ( .A1(n1330), .A2(n1331), .ZN(n1324) );
AND3_X1 U955 ( .A1(KEYINPUT1), .A2(n1141), .A3(n1323), .ZN(n1330) );
NOR3_X1 U956 ( .A1(n1332), .A2(n1309), .A3(n1333), .ZN(n1320) );
INV_X1 U957 ( .A(n1334), .ZN(n1333) );
XNOR2_X1 U958 ( .A(KEYINPUT26), .B(n1130), .ZN(n1332) );
NAND2_X1 U959 ( .A1(KEYINPUT51), .A2(n1335), .ZN(n1294) );
NOR2_X1 U960 ( .A1(n1183), .A2(G952), .ZN(n1236) );
XNOR2_X1 U961 ( .A(n1336), .B(n1337), .ZN(G48) );
NOR2_X1 U962 ( .A1(n1338), .A2(n1310), .ZN(n1337) );
NAND3_X1 U963 ( .A1(n1339), .A2(n1147), .A3(n1323), .ZN(n1310) );
XNOR2_X1 U964 ( .A(n1340), .B(KEYINPUT47), .ZN(n1338) );
XOR2_X1 U965 ( .A(n1341), .B(G143), .Z(G45) );
NAND2_X1 U966 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
NAND2_X1 U967 ( .A1(n1307), .A2(n1344), .ZN(n1343) );
INV_X1 U968 ( .A(KEYINPUT53), .ZN(n1344) );
NOR2_X1 U969 ( .A1(n1345), .A2(n1327), .ZN(n1307) );
NAND3_X1 U970 ( .A1(n1147), .A2(n1345), .A3(KEYINPUT53), .ZN(n1342) );
NAND4_X1 U971 ( .A1(n1148), .A2(n1339), .A3(n1346), .A4(n1347), .ZN(n1345) );
XNOR2_X1 U972 ( .A(G140), .B(n1303), .ZN(G42) );
NAND3_X1 U973 ( .A1(n1348), .A2(n1323), .A3(n1154), .ZN(n1303) );
XNOR2_X1 U974 ( .A(G137), .B(n1302), .ZN(G39) );
NAND3_X1 U975 ( .A1(n1340), .A2(n1348), .A3(n1349), .ZN(n1302) );
XNOR2_X1 U976 ( .A(G134), .B(n1311), .ZN(G36) );
NAND3_X1 U977 ( .A1(n1148), .A2(n1127), .A3(n1348), .ZN(n1311) );
XNOR2_X1 U978 ( .A(G131), .B(n1301), .ZN(G33) );
NAND3_X1 U979 ( .A1(n1323), .A2(n1148), .A3(n1348), .ZN(n1301) );
AND2_X1 U980 ( .A1(n1140), .A2(n1339), .ZN(n1348) );
AND2_X1 U981 ( .A1(n1132), .A2(n1350), .ZN(n1339) );
NOR2_X1 U982 ( .A1(n1156), .A2(n1152), .ZN(n1140) );
INV_X1 U983 ( .A(n1155), .ZN(n1152) );
XNOR2_X1 U984 ( .A(G128), .B(n1312), .ZN(G30) );
NAND4_X1 U985 ( .A1(n1351), .A2(n1340), .A3(n1127), .A4(n1352), .ZN(n1312) );
XNOR2_X1 U986 ( .A(G101), .B(n1353), .ZN(G3) );
NAND4_X1 U987 ( .A1(n1352), .A2(n1331), .A3(n1354), .A4(n1329), .ZN(n1353) );
NOR2_X1 U988 ( .A1(n1355), .A2(n1130), .ZN(n1329) );
INV_X1 U989 ( .A(n1349), .ZN(n1130) );
XNOR2_X1 U990 ( .A(KEYINPUT9), .B(n1327), .ZN(n1354) );
XNOR2_X1 U991 ( .A(G125), .B(n1304), .ZN(G27) );
NAND4_X1 U992 ( .A1(n1351), .A2(n1154), .A3(n1323), .A4(n1128), .ZN(n1304) );
AND2_X1 U993 ( .A1(n1147), .A2(n1350), .ZN(n1351) );
NAND2_X1 U994 ( .A1(n1356), .A2(n1143), .ZN(n1350) );
NAND3_X1 U995 ( .A1(n1357), .A2(n1185), .A3(n1358), .ZN(n1356) );
XNOR2_X1 U996 ( .A(G953), .B(KEYINPUT0), .ZN(n1358) );
INV_X1 U997 ( .A(G900), .ZN(n1185) );
INV_X1 U998 ( .A(n1327), .ZN(n1147) );
NAND2_X1 U999 ( .A1(n1359), .A2(n1360), .ZN(G24) );
NAND2_X1 U1000 ( .A1(G122), .A2(n1361), .ZN(n1360) );
XOR2_X1 U1001 ( .A(n1362), .B(KEYINPUT22), .Z(n1359) );
NAND2_X1 U1002 ( .A1(n1319), .A2(n1363), .ZN(n1362) );
INV_X1 U1003 ( .A(n1361), .ZN(n1319) );
NAND4_X1 U1004 ( .A1(n1334), .A2(n1141), .A3(n1346), .A4(n1347), .ZN(n1361) );
NOR2_X1 U1005 ( .A1(n1364), .A2(n1164), .ZN(n1141) );
XOR2_X1 U1006 ( .A(n1365), .B(n1366), .Z(G21) );
XNOR2_X1 U1007 ( .A(G119), .B(KEYINPUT42), .ZN(n1366) );
NAND3_X1 U1008 ( .A1(n1349), .A2(n1340), .A3(n1334), .ZN(n1365) );
INV_X1 U1009 ( .A(n1309), .ZN(n1340) );
NAND2_X1 U1010 ( .A1(n1164), .A2(n1364), .ZN(n1309) );
INV_X1 U1011 ( .A(n1367), .ZN(n1364) );
XNOR2_X1 U1012 ( .A(G116), .B(n1317), .ZN(G18) );
NAND3_X1 U1013 ( .A1(n1148), .A2(n1127), .A3(n1334), .ZN(n1317) );
NOR2_X1 U1014 ( .A1(n1347), .A2(n1157), .ZN(n1127) );
XNOR2_X1 U1015 ( .A(G113), .B(n1313), .ZN(G15) );
NAND3_X1 U1016 ( .A1(n1323), .A2(n1148), .A3(n1334), .ZN(n1313) );
NOR3_X1 U1017 ( .A1(n1327), .A2(n1328), .A3(n1136), .ZN(n1334) );
INV_X1 U1018 ( .A(n1128), .ZN(n1136) );
NOR2_X1 U1019 ( .A1(n1133), .A2(n1368), .ZN(n1128) );
INV_X1 U1020 ( .A(n1134), .ZN(n1368) );
INV_X1 U1021 ( .A(n1355), .ZN(n1148) );
NAND2_X1 U1022 ( .A1(n1367), .A2(n1164), .ZN(n1355) );
INV_X1 U1023 ( .A(n1139), .ZN(n1323) );
NAND2_X1 U1024 ( .A1(n1157), .A2(n1347), .ZN(n1139) );
INV_X1 U1025 ( .A(n1346), .ZN(n1157) );
XNOR2_X1 U1026 ( .A(G110), .B(n1316), .ZN(G12) );
NAND3_X1 U1027 ( .A1(n1349), .A2(n1318), .A3(n1154), .ZN(n1316) );
NOR2_X1 U1028 ( .A1(n1164), .A2(n1367), .ZN(n1154) );
NOR2_X1 U1029 ( .A1(n1369), .A2(n1161), .ZN(n1367) );
NOR2_X1 U1030 ( .A1(n1168), .A2(n1167), .ZN(n1161) );
AND2_X1 U1031 ( .A1(n1167), .A2(n1168), .ZN(n1369) );
NAND2_X1 U1032 ( .A1(G217), .A2(n1370), .ZN(n1168) );
NOR2_X1 U1033 ( .A1(n1241), .A2(G902), .ZN(n1167) );
XNOR2_X1 U1034 ( .A(n1371), .B(n1372), .ZN(n1241) );
XOR2_X1 U1035 ( .A(n1373), .B(n1374), .Z(n1372) );
XOR2_X1 U1036 ( .A(n1375), .B(n1376), .Z(n1374) );
XNOR2_X1 U1037 ( .A(n1211), .B(n1377), .ZN(n1376) );
XOR2_X1 U1038 ( .A(G119), .B(n1378), .Z(n1377) );
AND3_X1 U1039 ( .A1(G221), .A2(n1183), .A3(G234), .ZN(n1378) );
INV_X1 U1040 ( .A(n1206), .ZN(n1211) );
XNOR2_X1 U1041 ( .A(G128), .B(n1379), .ZN(n1375) );
XNOR2_X1 U1042 ( .A(KEYINPUT58), .B(n1336), .ZN(n1379) );
NAND2_X1 U1043 ( .A1(KEYINPUT8), .A2(n1380), .ZN(n1373) );
XNOR2_X1 U1044 ( .A(KEYINPUT21), .B(n1210), .ZN(n1380) );
XNOR2_X1 U1045 ( .A(n1381), .B(n1382), .ZN(n1371) );
NAND2_X1 U1046 ( .A1(KEYINPUT36), .A2(n1383), .ZN(n1382) );
NAND2_X1 U1047 ( .A1(KEYINPUT38), .A2(n1199), .ZN(n1381) );
XOR2_X1 U1048 ( .A(n1384), .B(n1265), .Z(n1164) );
INV_X1 U1049 ( .A(G472), .ZN(n1265) );
NAND2_X1 U1050 ( .A1(n1385), .A2(n1386), .ZN(n1384) );
XOR2_X1 U1051 ( .A(n1387), .B(n1388), .Z(n1385) );
XNOR2_X1 U1052 ( .A(n1389), .B(n1262), .ZN(n1388) );
XOR2_X1 U1053 ( .A(G113), .B(n1390), .Z(n1262) );
NAND2_X1 U1054 ( .A1(n1267), .A2(n1268), .ZN(n1389) );
NAND2_X1 U1055 ( .A1(n1391), .A2(n1392), .ZN(n1268) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1393), .ZN(n1392) );
NAND3_X1 U1057 ( .A1(G210), .A2(n1393), .A3(G101), .ZN(n1267) );
NAND2_X1 U1058 ( .A1(n1394), .A2(n1395), .ZN(n1387) );
NAND2_X1 U1059 ( .A1(n1261), .A2(n1396), .ZN(n1395) );
INV_X1 U1060 ( .A(KEYINPUT13), .ZN(n1396) );
XNOR2_X1 U1061 ( .A(n1273), .B(n1397), .ZN(n1261) );
XNOR2_X1 U1062 ( .A(n1398), .B(n1202), .ZN(n1273) );
XOR2_X1 U1063 ( .A(n1399), .B(n1400), .Z(n1202) );
NAND3_X1 U1064 ( .A1(n1401), .A2(n1291), .A3(KEYINPUT13), .ZN(n1394) );
NOR3_X1 U1065 ( .A1(n1326), .A2(n1328), .A3(n1327), .ZN(n1318) );
NAND2_X1 U1066 ( .A1(n1156), .A2(n1155), .ZN(n1327) );
NAND2_X1 U1067 ( .A1(G214), .A2(n1402), .ZN(n1155) );
XNOR2_X1 U1068 ( .A(n1179), .B(n1178), .ZN(n1156) );
NAND2_X1 U1069 ( .A1(G210), .A2(n1402), .ZN(n1178) );
NAND2_X1 U1070 ( .A1(n1403), .A2(n1386), .ZN(n1402) );
INV_X1 U1071 ( .A(G237), .ZN(n1403) );
AND2_X1 U1072 ( .A1(n1404), .A2(n1386), .ZN(n1179) );
XNOR2_X1 U1073 ( .A(n1405), .B(n1406), .ZN(n1404) );
XOR2_X1 U1074 ( .A(n1407), .B(n1335), .Z(n1406) );
NAND2_X1 U1075 ( .A1(G224), .A2(n1183), .ZN(n1335) );
NAND3_X1 U1076 ( .A1(n1408), .A2(n1409), .A3(n1410), .ZN(n1407) );
NAND2_X1 U1077 ( .A1(n1287), .A2(n1411), .ZN(n1410) );
NAND2_X1 U1078 ( .A1(KEYINPUT34), .A2(n1412), .ZN(n1411) );
XNOR2_X1 U1079 ( .A(KEYINPUT40), .B(n1210), .ZN(n1412) );
NAND3_X1 U1080 ( .A1(KEYINPUT34), .A2(n1291), .A3(n1210), .ZN(n1409) );
INV_X1 U1081 ( .A(n1287), .ZN(n1291) );
XOR2_X1 U1082 ( .A(n1397), .B(n1400), .Z(n1287) );
AND2_X1 U1083 ( .A1(KEYINPUT20), .A2(n1193), .ZN(n1397) );
OR2_X1 U1084 ( .A1(n1210), .A2(KEYINPUT34), .ZN(n1408) );
INV_X1 U1085 ( .A(G125), .ZN(n1210) );
INV_X1 U1086 ( .A(n1280), .ZN(n1405) );
XOR2_X1 U1087 ( .A(n1231), .B(n1413), .Z(n1280) );
XNOR2_X1 U1088 ( .A(n1227), .B(n1414), .ZN(n1413) );
NAND2_X1 U1089 ( .A1(KEYINPUT33), .A2(n1230), .ZN(n1414) );
XNOR2_X1 U1090 ( .A(n1415), .B(n1416), .ZN(n1230) );
XNOR2_X1 U1091 ( .A(G107), .B(n1417), .ZN(n1416) );
NAND2_X1 U1092 ( .A1(n1418), .A2(n1391), .ZN(n1415) );
XNOR2_X1 U1093 ( .A(KEYINPUT25), .B(KEYINPUT10), .ZN(n1418) );
AND2_X1 U1094 ( .A1(n1419), .A2(n1420), .ZN(n1227) );
NAND2_X1 U1095 ( .A1(G122), .A2(n1383), .ZN(n1420) );
XOR2_X1 U1096 ( .A(n1421), .B(KEYINPUT17), .Z(n1419) );
NAND2_X1 U1097 ( .A1(n1422), .A2(n1363), .ZN(n1421) );
XNOR2_X1 U1098 ( .A(G110), .B(KEYINPUT41), .ZN(n1422) );
XNOR2_X1 U1099 ( .A(n1423), .B(n1390), .ZN(n1231) );
XOR2_X1 U1100 ( .A(G116), .B(G119), .Z(n1390) );
NAND2_X1 U1101 ( .A1(KEYINPUT61), .A2(n1424), .ZN(n1423) );
INV_X1 U1102 ( .A(G113), .ZN(n1424) );
INV_X1 U1103 ( .A(n1331), .ZN(n1328) );
NAND2_X1 U1104 ( .A1(n1425), .A2(n1143), .ZN(n1331) );
NAND3_X1 U1105 ( .A1(n1426), .A2(n1183), .A3(G952), .ZN(n1143) );
NAND3_X1 U1106 ( .A1(n1357), .A2(n1223), .A3(G953), .ZN(n1425) );
INV_X1 U1107 ( .A(G898), .ZN(n1223) );
AND2_X1 U1108 ( .A1(G902), .A2(n1426), .ZN(n1357) );
NAND2_X1 U1109 ( .A1(G237), .A2(G234), .ZN(n1426) );
INV_X1 U1110 ( .A(n1352), .ZN(n1326) );
XOR2_X1 U1111 ( .A(n1132), .B(KEYINPUT15), .Z(n1352) );
AND2_X1 U1112 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U1113 ( .A1(G221), .A2(n1370), .ZN(n1134) );
NAND2_X1 U1114 ( .A1(G234), .A2(n1386), .ZN(n1370) );
XOR2_X1 U1115 ( .A(n1427), .B(n1275), .Z(n1133) );
INV_X1 U1116 ( .A(G469), .ZN(n1275) );
NAND2_X1 U1117 ( .A1(n1428), .A2(n1386), .ZN(n1427) );
INV_X1 U1118 ( .A(G902), .ZN(n1386) );
XOR2_X1 U1119 ( .A(n1400), .B(n1429), .Z(n1428) );
XNOR2_X1 U1120 ( .A(n1430), .B(n1272), .ZN(n1429) );
XNOR2_X1 U1121 ( .A(n1431), .B(n1432), .ZN(n1272) );
XOR2_X1 U1122 ( .A(n1433), .B(n1434), .Z(n1432) );
XNOR2_X1 U1123 ( .A(n1383), .B(G104), .ZN(n1434) );
INV_X1 U1124 ( .A(G110), .ZN(n1383) );
XOR2_X1 U1125 ( .A(KEYINPUT50), .B(KEYINPUT2), .Z(n1433) );
XOR2_X1 U1126 ( .A(n1435), .B(n1436), .Z(n1431) );
XNOR2_X1 U1127 ( .A(n1391), .B(n1437), .ZN(n1436) );
NOR2_X1 U1128 ( .A1(n1184), .A2(n1438), .ZN(n1437) );
XNOR2_X1 U1129 ( .A(KEYINPUT23), .B(n1183), .ZN(n1438) );
INV_X1 U1130 ( .A(G227), .ZN(n1184) );
INV_X1 U1131 ( .A(G101), .ZN(n1391) );
XNOR2_X1 U1132 ( .A(n1439), .B(n1206), .ZN(n1435) );
NAND2_X1 U1133 ( .A1(KEYINPUT4), .A2(n1401), .ZN(n1430) );
XNOR2_X1 U1134 ( .A(n1398), .B(n1399), .ZN(n1401) );
NAND2_X1 U1135 ( .A1(n1440), .A2(n1441), .ZN(n1398) );
INV_X1 U1136 ( .A(n1195), .ZN(n1441) );
NOR2_X1 U1137 ( .A1(n1199), .A2(G134), .ZN(n1195) );
INV_X1 U1138 ( .A(G137), .ZN(n1199) );
XOR2_X1 U1139 ( .A(KEYINPUT55), .B(n1442), .Z(n1440) );
NOR2_X1 U1140 ( .A1(G137), .A2(n1200), .ZN(n1442) );
XOR2_X1 U1141 ( .A(G143), .B(G146), .Z(n1400) );
NOR2_X1 U1142 ( .A1(n1346), .A2(n1347), .ZN(n1349) );
XOR2_X1 U1143 ( .A(n1443), .B(n1444), .Z(n1347) );
INV_X1 U1144 ( .A(n1172), .ZN(n1444) );
NOR2_X1 U1145 ( .A1(n1255), .A2(G902), .ZN(n1172) );
XNOR2_X1 U1146 ( .A(n1445), .B(n1446), .ZN(n1255) );
XOR2_X1 U1147 ( .A(n1447), .B(n1448), .Z(n1446) );
NAND2_X1 U1148 ( .A1(n1449), .A2(n1450), .ZN(n1448) );
NAND2_X1 U1149 ( .A1(n1451), .A2(n1417), .ZN(n1450) );
XOR2_X1 U1150 ( .A(KEYINPUT56), .B(n1452), .Z(n1449) );
NOR2_X1 U1151 ( .A1(n1451), .A2(n1417), .ZN(n1452) );
INV_X1 U1152 ( .A(G104), .ZN(n1417) );
XNOR2_X1 U1153 ( .A(G113), .B(G122), .ZN(n1451) );
NAND2_X1 U1154 ( .A1(n1453), .A2(KEYINPUT28), .ZN(n1447) );
XOR2_X1 U1155 ( .A(n1454), .B(G143), .Z(n1453) );
NAND2_X1 U1156 ( .A1(G214), .A2(n1393), .ZN(n1454) );
NOR2_X1 U1157 ( .A1(G953), .A2(G237), .ZN(n1393) );
XOR2_X1 U1158 ( .A(n1455), .B(n1399), .Z(n1445) );
XOR2_X1 U1159 ( .A(G131), .B(KEYINPUT11), .Z(n1399) );
NAND2_X1 U1160 ( .A1(n1456), .A2(n1457), .ZN(n1455) );
NAND2_X1 U1161 ( .A1(n1458), .A2(n1336), .ZN(n1457) );
INV_X1 U1162 ( .A(G146), .ZN(n1336) );
XOR2_X1 U1163 ( .A(n1459), .B(KEYINPUT35), .Z(n1458) );
NAND2_X1 U1164 ( .A1(G146), .A2(n1460), .ZN(n1456) );
XOR2_X1 U1165 ( .A(n1459), .B(KEYINPUT5), .Z(n1460) );
XNOR2_X1 U1166 ( .A(G125), .B(n1206), .ZN(n1459) );
XOR2_X1 U1167 ( .A(G140), .B(KEYINPUT32), .Z(n1206) );
NAND2_X1 U1168 ( .A1(KEYINPUT12), .A2(G475), .ZN(n1443) );
XOR2_X1 U1169 ( .A(G478), .B(n1461), .Z(n1346) );
NOR2_X1 U1170 ( .A1(n1250), .A2(G902), .ZN(n1461) );
AND2_X1 U1171 ( .A1(n1462), .A2(n1463), .ZN(n1250) );
NAND2_X1 U1172 ( .A1(n1464), .A2(n1465), .ZN(n1463) );
XOR2_X1 U1173 ( .A(KEYINPUT43), .B(n1466), .Z(n1462) );
NOR2_X1 U1174 ( .A1(n1464), .A2(n1465), .ZN(n1466) );
XOR2_X1 U1175 ( .A(n1467), .B(n1468), .Z(n1465) );
XOR2_X1 U1176 ( .A(n1469), .B(n1439), .Z(n1468) );
XNOR2_X1 U1177 ( .A(G107), .B(n1193), .ZN(n1439) );
INV_X1 U1178 ( .A(G128), .ZN(n1193) );
NOR2_X1 U1179 ( .A1(KEYINPUT30), .A2(n1363), .ZN(n1469) );
INV_X1 U1180 ( .A(G122), .ZN(n1363) );
XNOR2_X1 U1181 ( .A(G116), .B(n1470), .ZN(n1467) );
XNOR2_X1 U1182 ( .A(G143), .B(n1200), .ZN(n1470) );
INV_X1 U1183 ( .A(G134), .ZN(n1200) );
AND3_X1 U1184 ( .A1(G217), .A2(n1183), .A3(G234), .ZN(n1464) );
INV_X1 U1185 ( .A(G953), .ZN(n1183) );
endmodule


