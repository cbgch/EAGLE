//Key = 1010011110110100010100101011110001000111100000101010100101010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;

XOR2_X1 U720 ( .A(G107), .B(n992), .Z(G9) );
NOR2_X1 U721 ( .A1(n993), .A2(n994), .ZN(G75) );
NOR3_X1 U722 ( .A1(n995), .A2(n996), .A3(n997), .ZN(n994) );
NOR2_X1 U723 ( .A1(n998), .A2(n999), .ZN(n996) );
NOR2_X1 U724 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR2_X1 U725 ( .A1(KEYINPUT50), .A2(n1002), .ZN(n1001) );
NOR4_X1 U726 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n1002) );
NOR2_X1 U727 ( .A1(n1007), .A2(n1006), .ZN(n1000) );
NOR2_X1 U728 ( .A1(n1008), .A2(n1009), .ZN(n1007) );
AND2_X1 U729 ( .A1(n1010), .A2(n1011), .ZN(n1009) );
NOR2_X1 U730 ( .A1(n1012), .A2(n1003), .ZN(n1008) );
NOR2_X1 U731 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
AND2_X1 U732 ( .A1(n1011), .A2(n1015), .ZN(n1014) );
AND3_X1 U733 ( .A1(KEYINPUT50), .A2(n1016), .A3(n1017), .ZN(n1013) );
NAND3_X1 U734 ( .A1(n1018), .A2(n1019), .A3(n1020), .ZN(n995) );
NAND3_X1 U735 ( .A1(n1017), .A2(n1021), .A3(n1022), .ZN(n1020) );
INV_X1 U736 ( .A(n1006), .ZN(n1022) );
NAND2_X1 U737 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
NAND3_X1 U738 ( .A1(n1025), .A2(n1026), .A3(n1011), .ZN(n1024) );
NAND2_X1 U739 ( .A1(n1027), .A2(n1028), .ZN(n1023) );
NAND2_X1 U740 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
NAND4_X1 U741 ( .A1(KEYINPUT33), .A2(n1031), .A3(n1032), .A4(n1025), .ZN(n1030) );
NAND2_X1 U742 ( .A1(n1011), .A2(n1033), .ZN(n1029) );
NAND3_X1 U743 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
OR2_X1 U744 ( .A1(n999), .A2(KEYINPUT33), .ZN(n1036) );
NAND3_X1 U745 ( .A1(G214), .A2(n1037), .A3(n1038), .ZN(n1034) );
NOR3_X1 U746 ( .A1(n1039), .A2(G953), .A3(G952), .ZN(n993) );
INV_X1 U747 ( .A(n1018), .ZN(n1039) );
NAND4_X1 U748 ( .A1(n1040), .A2(n1041), .A3(n1042), .A4(n1043), .ZN(n1018) );
NOR4_X1 U749 ( .A1(n1044), .A2(n1045), .A3(n999), .A4(n1046), .ZN(n1043) );
NOR2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U751 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
AND2_X1 U752 ( .A1(n1051), .A2(KEYINPUT6), .ZN(n1050) );
NOR2_X1 U753 ( .A1(KEYINPUT6), .A2(n1052), .ZN(n1049) );
INV_X1 U754 ( .A(G478), .ZN(n1047) );
NOR2_X1 U755 ( .A1(G478), .A2(n1051), .ZN(n1044) );
NAND2_X1 U756 ( .A1(KEYINPUT39), .A2(n1053), .ZN(n1051) );
XNOR2_X1 U757 ( .A(KEYINPUT0), .B(n1054), .ZN(n1041) );
XOR2_X1 U758 ( .A(KEYINPUT27), .B(n1055), .Z(n1040) );
XOR2_X1 U759 ( .A(n1056), .B(n1057), .Z(G72) );
XOR2_X1 U760 ( .A(n1058), .B(n1059), .Z(n1057) );
NOR2_X1 U761 ( .A1(n1060), .A2(G953), .ZN(n1059) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1062), .ZN(n1058) );
XOR2_X1 U763 ( .A(n1063), .B(n1064), .Z(n1062) );
XNOR2_X1 U764 ( .A(n1065), .B(n1066), .ZN(n1064) );
INV_X1 U765 ( .A(n1067), .ZN(n1066) );
XOR2_X1 U766 ( .A(n1068), .B(n1069), .Z(n1063) );
XNOR2_X1 U767 ( .A(G131), .B(KEYINPUT36), .ZN(n1069) );
NAND3_X1 U768 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1068) );
NAND2_X1 U769 ( .A1(KEYINPUT23), .A2(G134), .ZN(n1072) );
NAND3_X1 U770 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1071) );
INV_X1 U771 ( .A(KEYINPUT23), .ZN(n1074) );
OR2_X1 U772 ( .A1(n1075), .A2(n1073), .ZN(n1070) );
NOR2_X1 U773 ( .A1(G134), .A2(KEYINPUT25), .ZN(n1073) );
XNOR2_X1 U774 ( .A(G137), .B(KEYINPUT44), .ZN(n1075) );
XOR2_X1 U775 ( .A(KEYINPUT21), .B(n1076), .Z(n1061) );
NOR2_X1 U776 ( .A1(n1077), .A2(n1019), .ZN(n1056) );
AND2_X1 U777 ( .A1(G227), .A2(G900), .ZN(n1077) );
XOR2_X1 U778 ( .A(n1078), .B(n1079), .Z(G69) );
NOR2_X1 U779 ( .A1(n1080), .A2(n1019), .ZN(n1079) );
AND2_X1 U780 ( .A1(G224), .A2(G898), .ZN(n1080) );
NAND2_X1 U781 ( .A1(n1081), .A2(n1082), .ZN(n1078) );
NAND3_X1 U782 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
NAND2_X1 U783 ( .A1(G953), .A2(n1086), .ZN(n1084) );
XOR2_X1 U784 ( .A(KEYINPUT55), .B(n1087), .Z(n1081) );
NOR3_X1 U785 ( .A1(n1083), .A2(G953), .A3(n1085), .ZN(n1087) );
XOR2_X1 U786 ( .A(n1088), .B(KEYINPUT53), .Z(n1083) );
NOR2_X1 U787 ( .A1(n1089), .A2(n1090), .ZN(G66) );
XOR2_X1 U788 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND3_X1 U789 ( .A1(n1093), .A2(n997), .A3(n1094), .ZN(n1091) );
XNOR2_X1 U790 ( .A(KEYINPUT62), .B(n1095), .ZN(n1093) );
NOR2_X1 U791 ( .A1(n1089), .A2(n1096), .ZN(G63) );
NOR3_X1 U792 ( .A1(n1053), .A2(n1097), .A3(n1098), .ZN(n1096) );
NOR3_X1 U793 ( .A1(n1099), .A2(n1100), .A3(n1095), .ZN(n1098) );
AND2_X1 U794 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NAND2_X1 U795 ( .A1(G478), .A2(n997), .ZN(n1099) );
INV_X1 U796 ( .A(n1052), .ZN(n1053) );
NOR2_X1 U797 ( .A1(n1101), .A2(n1102), .ZN(G60) );
XOR2_X1 U798 ( .A(n1103), .B(n1104), .Z(n1102) );
NAND3_X1 U799 ( .A1(G475), .A2(n997), .A3(n1105), .ZN(n1103) );
XNOR2_X1 U800 ( .A(G902), .B(KEYINPUT17), .ZN(n1105) );
XNOR2_X1 U801 ( .A(n1089), .B(KEYINPUT7), .ZN(n1101) );
XNOR2_X1 U802 ( .A(G104), .B(n1106), .ZN(G6) );
NAND4_X1 U803 ( .A1(n1107), .A2(n1017), .A3(n1108), .A4(n1109), .ZN(n1106) );
OR2_X1 U804 ( .A1(n1110), .A2(KEYINPUT60), .ZN(n1109) );
NAND2_X1 U805 ( .A1(KEYINPUT60), .A2(n1111), .ZN(n1108) );
NAND3_X1 U806 ( .A1(n1004), .A2(n1112), .A3(n1113), .ZN(n1111) );
NOR2_X1 U807 ( .A1(n1089), .A2(n1114), .ZN(G57) );
XOR2_X1 U808 ( .A(n1115), .B(n1116), .Z(n1114) );
XNOR2_X1 U809 ( .A(n1117), .B(n1118), .ZN(n1116) );
XNOR2_X1 U810 ( .A(n1119), .B(n1120), .ZN(n1115) );
XOR2_X1 U811 ( .A(KEYINPUT34), .B(n1121), .Z(n1120) );
NOR3_X1 U812 ( .A1(n1095), .A2(n1122), .A3(n1123), .ZN(n1121) );
XOR2_X1 U813 ( .A(n997), .B(KEYINPUT63), .Z(n1122) );
NOR2_X1 U814 ( .A1(n1089), .A2(n1124), .ZN(G54) );
XOR2_X1 U815 ( .A(n1125), .B(n1126), .Z(n1124) );
XNOR2_X1 U816 ( .A(n1067), .B(n1127), .ZN(n1126) );
XOR2_X1 U817 ( .A(n1128), .B(n1129), .Z(n1127) );
XNOR2_X1 U818 ( .A(n1130), .B(n1131), .ZN(n1125) );
XOR2_X1 U819 ( .A(n1132), .B(KEYINPUT18), .Z(n1131) );
NAND3_X1 U820 ( .A1(G902), .A2(n997), .A3(G469), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1089), .A2(n1133), .ZN(G51) );
XOR2_X1 U822 ( .A(n1088), .B(n1134), .Z(n1133) );
XOR2_X1 U823 ( .A(n1135), .B(n1136), .Z(n1134) );
NAND3_X1 U824 ( .A1(G902), .A2(n997), .A3(n1137), .ZN(n1136) );
NAND2_X1 U825 ( .A1(n1085), .A2(n1060), .ZN(n997) );
AND4_X1 U826 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1060) );
NOR4_X1 U827 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
AND2_X1 U828 ( .A1(n1146), .A2(n1147), .ZN(n1140) );
NAND2_X1 U829 ( .A1(n1148), .A2(n1025), .ZN(n1138) );
INV_X1 U830 ( .A(n999), .ZN(n1025) );
XOR2_X1 U831 ( .A(n1149), .B(KEYINPUT59), .Z(n1148) );
AND4_X1 U832 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1153), .ZN(n1085) );
NOR4_X1 U833 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n992), .ZN(n1153) );
NOR3_X1 U834 ( .A1(n1157), .A2(n1158), .A3(n1005), .ZN(n992) );
NOR2_X1 U835 ( .A1(n1159), .A2(n1160), .ZN(n1152) );
NOR3_X1 U836 ( .A1(n1161), .A2(n1011), .A3(n1162), .ZN(n1160) );
INV_X1 U837 ( .A(n1046), .ZN(n1011) );
AND2_X1 U838 ( .A1(n1161), .A2(n1163), .ZN(n1159) );
INV_X1 U839 ( .A(KEYINPUT15), .ZN(n1161) );
NAND3_X1 U840 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1151) );
XNOR2_X1 U841 ( .A(n1003), .B(KEYINPUT35), .ZN(n1164) );
NAND2_X1 U842 ( .A1(n1110), .A2(n1010), .ZN(n1150) );
NAND2_X1 U843 ( .A1(n1167), .A2(n1168), .ZN(n1010) );
NAND2_X1 U844 ( .A1(n1107), .A2(n1017), .ZN(n1168) );
NAND2_X1 U845 ( .A1(n1169), .A2(n1027), .ZN(n1167) );
NAND2_X1 U846 ( .A1(KEYINPUT28), .A2(n1170), .ZN(n1135) );
NAND2_X1 U847 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND2_X1 U848 ( .A1(n1173), .A2(n1174), .ZN(n1172) );
XOR2_X1 U849 ( .A(KEYINPUT46), .B(n1175), .Z(n1171) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1173), .ZN(n1175) );
XNOR2_X1 U851 ( .A(n1176), .B(n1177), .ZN(n1173) );
NOR2_X1 U852 ( .A1(n1019), .A2(G952), .ZN(n1089) );
XNOR2_X1 U853 ( .A(n1139), .B(n1178), .ZN(G48) );
NOR2_X1 U854 ( .A1(KEYINPUT51), .A2(n1179), .ZN(n1178) );
NAND3_X1 U855 ( .A1(n1166), .A2(n1107), .A3(n1180), .ZN(n1139) );
XNOR2_X1 U856 ( .A(G143), .B(n1147), .ZN(G45) );
NAND4_X1 U857 ( .A1(n1181), .A2(n1180), .A3(n1015), .A4(n1182), .ZN(n1147) );
XNOR2_X1 U858 ( .A(n1183), .B(KEYINPUT29), .ZN(n1181) );
XOR2_X1 U859 ( .A(G140), .B(n1184), .Z(G42) );
NOR2_X1 U860 ( .A1(n999), .A2(n1149), .ZN(n1184) );
NAND4_X1 U861 ( .A1(n1169), .A2(n1107), .A3(n1016), .A4(n1185), .ZN(n1149) );
XNOR2_X1 U862 ( .A(G137), .B(n1186), .ZN(G39) );
NOR2_X1 U863 ( .A1(n1145), .A2(KEYINPUT9), .ZN(n1186) );
AND3_X1 U864 ( .A1(n1166), .A2(n1027), .A3(n1187), .ZN(n1145) );
XNOR2_X1 U865 ( .A(n1144), .B(n1188), .ZN(G36) );
XNOR2_X1 U866 ( .A(G134), .B(KEYINPUT43), .ZN(n1188) );
AND3_X1 U867 ( .A1(n1015), .A2(n1026), .A3(n1187), .ZN(n1144) );
XNOR2_X1 U868 ( .A(G131), .B(n1189), .ZN(G33) );
NOR2_X1 U869 ( .A1(n1143), .A2(KEYINPUT54), .ZN(n1189) );
AND3_X1 U870 ( .A1(n1107), .A2(n1015), .A3(n1187), .ZN(n1143) );
NOR3_X1 U871 ( .A1(n1004), .A2(n1190), .A3(n999), .ZN(n1187) );
NAND2_X1 U872 ( .A1(n1038), .A2(n1191), .ZN(n999) );
NAND2_X1 U873 ( .A1(G214), .A2(n1037), .ZN(n1191) );
NAND2_X1 U874 ( .A1(n1192), .A2(n1193), .ZN(G30) );
NAND2_X1 U875 ( .A1(G128), .A2(n1146), .ZN(n1193) );
XOR2_X1 U876 ( .A(KEYINPUT5), .B(n1194), .Z(n1192) );
NOR2_X1 U877 ( .A1(G128), .A2(n1146), .ZN(n1194) );
NAND3_X1 U878 ( .A1(n1166), .A2(n1026), .A3(n1180), .ZN(n1146) );
NOR3_X1 U879 ( .A1(n1035), .A2(n1190), .A3(n1004), .ZN(n1180) );
INV_X1 U880 ( .A(n1016), .ZN(n1004) );
XNOR2_X1 U881 ( .A(G101), .B(n1195), .ZN(G3) );
NOR2_X1 U882 ( .A1(n1156), .A2(KEYINPUT20), .ZN(n1195) );
AND3_X1 U883 ( .A1(n1110), .A2(n1027), .A3(n1015), .ZN(n1156) );
INV_X1 U884 ( .A(n1157), .ZN(n1110) );
NAND3_X1 U885 ( .A1(n1113), .A2(n1112), .A3(n1016), .ZN(n1157) );
XNOR2_X1 U886 ( .A(G125), .B(n1196), .ZN(G27) );
NAND2_X1 U887 ( .A1(KEYINPUT37), .A2(n1142), .ZN(n1196) );
AND3_X1 U888 ( .A1(n1169), .A2(n1107), .A3(n1197), .ZN(n1142) );
NOR3_X1 U889 ( .A1(n1046), .A2(n1190), .A3(n1035), .ZN(n1197) );
INV_X1 U890 ( .A(n1185), .ZN(n1190) );
NAND2_X1 U891 ( .A1(n1006), .A2(n1198), .ZN(n1185) );
NAND3_X1 U892 ( .A1(G902), .A2(n1199), .A3(n1076), .ZN(n1198) );
NOR2_X1 U893 ( .A1(n1019), .A2(G900), .ZN(n1076) );
XOR2_X1 U894 ( .A(G122), .B(n1155), .Z(G24) );
AND4_X1 U895 ( .A1(n1165), .A2(n1017), .A3(n1200), .A4(n1201), .ZN(n1155) );
OR2_X1 U896 ( .A1(n1026), .A2(KEYINPUT29), .ZN(n1201) );
NAND2_X1 U897 ( .A1(KEYINPUT29), .A2(n1202), .ZN(n1200) );
NAND2_X1 U898 ( .A1(n1183), .A2(n1182), .ZN(n1202) );
INV_X1 U899 ( .A(n1005), .ZN(n1017) );
NAND2_X1 U900 ( .A1(n1203), .A2(n1042), .ZN(n1005) );
XOR2_X1 U901 ( .A(G119), .B(n1204), .Z(G21) );
AND3_X1 U902 ( .A1(n1166), .A2(n1027), .A3(n1165), .ZN(n1204) );
NOR2_X1 U903 ( .A1(n1042), .A2(n1203), .ZN(n1166) );
INV_X1 U904 ( .A(n1205), .ZN(n1203) );
XNOR2_X1 U905 ( .A(G116), .B(n1206), .ZN(G18) );
NOR2_X1 U906 ( .A1(n1154), .A2(KEYINPUT47), .ZN(n1206) );
AND3_X1 U907 ( .A1(n1165), .A2(n1026), .A3(n1015), .ZN(n1154) );
INV_X1 U908 ( .A(n1158), .ZN(n1026) );
NAND2_X1 U909 ( .A1(n1054), .A2(n1182), .ZN(n1158) );
NOR3_X1 U910 ( .A1(n1035), .A2(n1207), .A3(n1046), .ZN(n1165) );
XOR2_X1 U911 ( .A(n1208), .B(n1163), .Z(G15) );
NOR2_X1 U912 ( .A1(n1162), .A2(n1046), .ZN(n1163) );
NAND2_X1 U913 ( .A1(n1032), .A2(n1209), .ZN(n1046) );
NAND4_X1 U914 ( .A1(n1107), .A2(n1015), .A3(n1113), .A4(n1112), .ZN(n1162) );
AND2_X1 U915 ( .A1(n1042), .A2(n1205), .ZN(n1015) );
XNOR2_X1 U916 ( .A(G113), .B(KEYINPUT57), .ZN(n1208) );
XNOR2_X1 U917 ( .A(G110), .B(n1210), .ZN(G12) );
NAND4_X1 U918 ( .A1(n1211), .A2(n1169), .A3(n1212), .A4(n1016), .ZN(n1210) );
NOR2_X1 U919 ( .A1(n1032), .A2(n1031), .ZN(n1016) );
INV_X1 U920 ( .A(n1209), .ZN(n1031) );
NAND2_X1 U921 ( .A1(G221), .A2(n1213), .ZN(n1209) );
XOR2_X1 U922 ( .A(n1214), .B(G469), .Z(n1032) );
NAND2_X1 U923 ( .A1(n1215), .A2(n1095), .ZN(n1214) );
XOR2_X1 U924 ( .A(n1128), .B(n1216), .Z(n1215) );
XNOR2_X1 U925 ( .A(n1217), .B(n1218), .ZN(n1216) );
NAND3_X1 U926 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1217) );
NAND2_X1 U927 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
INV_X1 U928 ( .A(KEYINPUT48), .ZN(n1223) );
NAND3_X1 U929 ( .A1(KEYINPUT48), .A2(n1224), .A3(n1067), .ZN(n1220) );
OR2_X1 U930 ( .A1(n1067), .A2(n1224), .ZN(n1219) );
NOR2_X1 U931 ( .A1(n1225), .A2(n1222), .ZN(n1224) );
XOR2_X1 U932 ( .A(G101), .B(n1129), .Z(n1222) );
INV_X1 U933 ( .A(KEYINPUT40), .ZN(n1225) );
XOR2_X1 U934 ( .A(G128), .B(n1226), .Z(n1067) );
NOR2_X1 U935 ( .A1(KEYINPUT45), .A2(n1227), .ZN(n1226) );
XNOR2_X1 U936 ( .A(G146), .B(G143), .ZN(n1227) );
XNOR2_X1 U937 ( .A(n1228), .B(n1229), .ZN(n1128) );
INV_X1 U938 ( .A(n1117), .ZN(n1229) );
XNOR2_X1 U939 ( .A(G140), .B(n1230), .ZN(n1228) );
AND2_X1 U940 ( .A1(n1019), .A2(G227), .ZN(n1230) );
NOR2_X1 U941 ( .A1(n1207), .A2(n1003), .ZN(n1212) );
INV_X1 U942 ( .A(n1027), .ZN(n1003) );
NAND2_X1 U943 ( .A1(n1231), .A2(n1232), .ZN(n1027) );
OR3_X1 U944 ( .A1(n1183), .A2(n1182), .A3(KEYINPUT31), .ZN(n1232) );
NAND2_X1 U945 ( .A1(KEYINPUT31), .A2(n1107), .ZN(n1231) );
NOR2_X1 U946 ( .A1(n1182), .A2(n1054), .ZN(n1107) );
INV_X1 U947 ( .A(n1183), .ZN(n1054) );
XNOR2_X1 U948 ( .A(n1233), .B(G475), .ZN(n1183) );
NAND2_X1 U949 ( .A1(n1104), .A2(n1095), .ZN(n1233) );
XOR2_X1 U950 ( .A(n1234), .B(n1235), .Z(n1104) );
XOR2_X1 U951 ( .A(G104), .B(n1236), .Z(n1235) );
NOR3_X1 U952 ( .A1(KEYINPUT56), .A2(n1237), .A3(n1238), .ZN(n1236) );
NOR2_X1 U953 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
XOR2_X1 U954 ( .A(n1241), .B(KEYINPUT3), .Z(n1240) );
NOR2_X1 U955 ( .A1(G143), .A2(n1242), .ZN(n1237) );
XOR2_X1 U956 ( .A(n1241), .B(KEYINPUT13), .Z(n1242) );
XOR2_X1 U957 ( .A(n1243), .B(n1244), .Z(n1241) );
XNOR2_X1 U958 ( .A(n1245), .B(n1246), .ZN(n1244) );
AND3_X1 U959 ( .A1(G214), .A2(n1019), .A3(n1247), .ZN(n1246) );
INV_X1 U960 ( .A(G131), .ZN(n1245) );
NAND2_X1 U961 ( .A1(n1248), .A2(KEYINPUT2), .ZN(n1243) );
XNOR2_X1 U962 ( .A(G146), .B(n1065), .ZN(n1248) );
NAND3_X1 U963 ( .A1(n1249), .A2(n1250), .A3(KEYINPUT10), .ZN(n1234) );
NAND2_X1 U964 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
XNOR2_X1 U965 ( .A(G113), .B(n1253), .ZN(n1251) );
OR3_X1 U966 ( .A1(n1254), .A2(n1253), .A3(n1252), .ZN(n1249) );
INV_X1 U967 ( .A(KEYINPUT12), .ZN(n1252) );
XOR2_X1 U968 ( .A(G122), .B(KEYINPUT30), .Z(n1253) );
XNOR2_X1 U969 ( .A(n1052), .B(G478), .ZN(n1182) );
NAND2_X1 U970 ( .A1(n1100), .A2(n1095), .ZN(n1052) );
XOR2_X1 U971 ( .A(n1255), .B(n1256), .Z(n1100) );
XOR2_X1 U972 ( .A(n1257), .B(n1258), .Z(n1256) );
NAND2_X1 U973 ( .A1(n1259), .A2(G217), .ZN(n1258) );
NAND2_X1 U974 ( .A1(n1260), .A2(KEYINPUT61), .ZN(n1257) );
XOR2_X1 U975 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U976 ( .A(KEYINPUT24), .B(G107), .Z(n1262) );
XNOR2_X1 U977 ( .A(G128), .B(n1263), .ZN(n1255) );
XNOR2_X1 U978 ( .A(n1239), .B(G134), .ZN(n1263) );
INV_X1 U979 ( .A(G143), .ZN(n1239) );
INV_X1 U980 ( .A(n1112), .ZN(n1207) );
NAND2_X1 U981 ( .A1(n1006), .A2(n1264), .ZN(n1112) );
NAND4_X1 U982 ( .A1(G953), .A2(G902), .A3(n1199), .A4(n1086), .ZN(n1264) );
INV_X1 U983 ( .A(G898), .ZN(n1086) );
NAND3_X1 U984 ( .A1(n1199), .A2(n1019), .A3(G952), .ZN(n1006) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1199) );
NOR2_X1 U986 ( .A1(n1205), .A2(n1042), .ZN(n1169) );
XOR2_X1 U987 ( .A(n1265), .B(n1094), .Z(n1042) );
AND2_X1 U988 ( .A1(G217), .A2(n1213), .ZN(n1094) );
NAND2_X1 U989 ( .A1(G234), .A2(n1266), .ZN(n1213) );
NAND2_X1 U990 ( .A1(n1092), .A2(n1095), .ZN(n1265) );
XOR2_X1 U991 ( .A(n1267), .B(n1268), .Z(n1092) );
XOR2_X1 U992 ( .A(n1269), .B(n1270), .Z(n1268) );
XOR2_X1 U993 ( .A(n1271), .B(G119), .Z(n1270) );
NAND2_X1 U994 ( .A1(G221), .A2(n1259), .ZN(n1271) );
AND2_X1 U995 ( .A1(G234), .A2(n1019), .ZN(n1259) );
XNOR2_X1 U996 ( .A(G137), .B(KEYINPUT32), .ZN(n1269) );
XOR2_X1 U997 ( .A(n1272), .B(n1273), .Z(n1267) );
XOR2_X1 U998 ( .A(n1274), .B(n1065), .Z(n1272) );
XNOR2_X1 U999 ( .A(G140), .B(n1176), .ZN(n1065) );
INV_X1 U1000 ( .A(G125), .ZN(n1176) );
NAND2_X1 U1001 ( .A1(KEYINPUT8), .A2(n1218), .ZN(n1274) );
XOR2_X1 U1002 ( .A(n1055), .B(KEYINPUT49), .Z(n1205) );
XOR2_X1 U1003 ( .A(n1275), .B(n1123), .Z(n1055) );
INV_X1 U1004 ( .A(G472), .ZN(n1123) );
NAND2_X1 U1005 ( .A1(n1276), .A2(n1095), .ZN(n1275) );
XNOR2_X1 U1006 ( .A(n1277), .B(n1118), .ZN(n1276) );
XOR2_X1 U1007 ( .A(n1278), .B(n1279), .Z(n1118) );
XNOR2_X1 U1008 ( .A(n1254), .B(G101), .ZN(n1279) );
INV_X1 U1009 ( .A(G113), .ZN(n1254) );
XOR2_X1 U1010 ( .A(n1280), .B(n1281), .Z(n1278) );
NOR2_X1 U1011 ( .A1(KEYINPUT14), .A2(n1282), .ZN(n1281) );
XNOR2_X1 U1012 ( .A(n1283), .B(n1284), .ZN(n1282) );
NOR2_X1 U1013 ( .A1(G119), .A2(KEYINPUT41), .ZN(n1284) );
NAND3_X1 U1014 ( .A1(n1247), .A2(n1019), .A3(G210), .ZN(n1280) );
NOR2_X1 U1015 ( .A1(n1285), .A2(n1286), .ZN(n1277) );
XOR2_X1 U1016 ( .A(n1287), .B(KEYINPUT19), .Z(n1286) );
NAND2_X1 U1017 ( .A1(n1288), .A2(n1177), .ZN(n1287) );
NOR2_X1 U1018 ( .A1(n1288), .A2(n1177), .ZN(n1285) );
XNOR2_X1 U1019 ( .A(KEYINPUT58), .B(n1117), .ZN(n1288) );
XNOR2_X1 U1020 ( .A(n1289), .B(n1290), .ZN(n1117) );
XOR2_X1 U1021 ( .A(KEYINPUT22), .B(G137), .Z(n1290) );
XNOR2_X1 U1022 ( .A(G131), .B(G134), .ZN(n1289) );
XOR2_X1 U1023 ( .A(n1113), .B(KEYINPUT4), .Z(n1211) );
XOR2_X1 U1024 ( .A(n1035), .B(KEYINPUT52), .Z(n1113) );
OR2_X1 U1025 ( .A1(n1038), .A2(n1291), .ZN(n1035) );
AND2_X1 U1026 ( .A1(G214), .A2(n1037), .ZN(n1291) );
XOR2_X1 U1027 ( .A(n1292), .B(n1137), .Z(n1038) );
AND2_X1 U1028 ( .A1(G210), .A2(n1037), .ZN(n1137) );
NAND2_X1 U1029 ( .A1(n1266), .A2(n1247), .ZN(n1037) );
INV_X1 U1030 ( .A(G237), .ZN(n1247) );
XNOR2_X1 U1031 ( .A(G902), .B(KEYINPUT1), .ZN(n1266) );
NAND2_X1 U1032 ( .A1(n1293), .A2(n1095), .ZN(n1292) );
INV_X1 U1033 ( .A(G902), .ZN(n1095) );
XOR2_X1 U1034 ( .A(n1294), .B(n1295), .Z(n1293) );
XNOR2_X1 U1035 ( .A(G125), .B(n1174), .ZN(n1295) );
NAND2_X1 U1036 ( .A1(G224), .A2(n1019), .ZN(n1174) );
INV_X1 U1037 ( .A(G953), .ZN(n1019) );
XNOR2_X1 U1038 ( .A(n1088), .B(n1296), .ZN(n1294) );
NOR2_X1 U1039 ( .A1(KEYINPUT42), .A2(n1119), .ZN(n1296) );
INV_X1 U1040 ( .A(n1177), .ZN(n1119) );
XOR2_X1 U1041 ( .A(G143), .B(n1273), .Z(n1177) );
XNOR2_X1 U1042 ( .A(G128), .B(n1179), .ZN(n1273) );
INV_X1 U1043 ( .A(G146), .ZN(n1179) );
XNOR2_X1 U1044 ( .A(n1297), .B(n1298), .ZN(n1088) );
XOR2_X1 U1045 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U1046 ( .A(G119), .B(KEYINPUT26), .ZN(n1300) );
NAND2_X1 U1047 ( .A1(KEYINPUT38), .A2(G113), .ZN(n1299) );
XOR2_X1 U1048 ( .A(n1301), .B(n1130), .Z(n1297) );
XNOR2_X1 U1049 ( .A(G101), .B(n1218), .ZN(n1130) );
INV_X1 U1050 ( .A(G110), .ZN(n1218) );
XOR2_X1 U1051 ( .A(n1261), .B(n1302), .Z(n1301) );
NOR2_X1 U1052 ( .A1(KEYINPUT16), .A2(n1129), .ZN(n1302) );
XOR2_X1 U1053 ( .A(G104), .B(G107), .Z(n1129) );
XNOR2_X1 U1054 ( .A(G122), .B(n1283), .ZN(n1261) );
XOR2_X1 U1055 ( .A(G116), .B(KEYINPUT11), .Z(n1283) );
endmodule


