//Key = 0110110110011101111001101110100111011100011000000101010010111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;

XNOR2_X1 U748 ( .A(G107), .B(n1030), .ZN(G9) );
NOR2_X1 U749 ( .A1(n1031), .A2(KEYINPUT52), .ZN(n1030) );
NOR2_X1 U750 ( .A1(n1032), .A2(n1033), .ZN(G75) );
NOR3_X1 U751 ( .A1(n1034), .A2(G953), .A3(n1035), .ZN(n1033) );
XOR2_X1 U752 ( .A(n1036), .B(KEYINPUT30), .Z(n1034) );
NAND3_X1 U753 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NAND2_X1 U754 ( .A1(n1040), .A2(n1041), .ZN(n1038) );
NAND2_X1 U755 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U756 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U757 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U758 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
OR2_X1 U759 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1047) );
NAND2_X1 U761 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U762 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
INV_X1 U763 ( .A(n1059), .ZN(n1055) );
NAND3_X1 U764 ( .A1(n1049), .A2(n1060), .A3(n1053), .ZN(n1042) );
NAND3_X1 U765 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND2_X1 U766 ( .A1(n1064), .A2(n1046), .ZN(n1063) );
NAND2_X1 U767 ( .A1(n1065), .A2(n1066), .ZN(n1062) );
XNOR2_X1 U768 ( .A(n1046), .B(KEYINPUT36), .ZN(n1065) );
NAND2_X1 U769 ( .A1(n1044), .A2(n1067), .ZN(n1061) );
NAND3_X1 U770 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
OR3_X1 U771 ( .A1(n1071), .A2(n1072), .A3(KEYINPUT54), .ZN(n1069) );
NAND2_X1 U772 ( .A1(KEYINPUT54), .A2(n1046), .ZN(n1068) );
INV_X1 U773 ( .A(n1073), .ZN(n1040) );
NOR3_X1 U774 ( .A1(n1035), .A2(G953), .A3(G952), .ZN(n1032) );
AND4_X1 U775 ( .A1(n1074), .A2(n1049), .A3(n1075), .A4(n1076), .ZN(n1035) );
NOR4_X1 U776 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
XNOR2_X1 U777 ( .A(n1072), .B(KEYINPUT13), .ZN(n1079) );
NOR2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1078) );
XOR2_X1 U779 ( .A(KEYINPUT7), .B(G475), .Z(n1082) );
INV_X1 U780 ( .A(n1083), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1084), .B(KEYINPUT29), .Z(n1075) );
XNOR2_X1 U782 ( .A(n1085), .B(G478), .ZN(n1074) );
XOR2_X1 U783 ( .A(n1086), .B(n1087), .Z(G72) );
NOR2_X1 U784 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U785 ( .A(n1090), .B(KEYINPUT25), .Z(n1089) );
NAND3_X1 U786 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1090) );
NOR2_X1 U787 ( .A1(n1094), .A2(n1091), .ZN(n1088) );
NAND2_X1 U788 ( .A1(n1095), .A2(n1096), .ZN(n1091) );
NAND2_X1 U789 ( .A1(G953), .A2(n1097), .ZN(n1096) );
XOR2_X1 U790 ( .A(n1098), .B(n1099), .Z(n1095) );
XOR2_X1 U791 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND4_X1 U792 ( .A1(n1102), .A2(n1103), .A3(n1104), .A4(n1105), .ZN(n1101) );
NAND3_X1 U793 ( .A1(G134), .A2(n1106), .A3(n1107), .ZN(n1105) );
NAND3_X1 U794 ( .A1(n1108), .A2(n1109), .A3(G131), .ZN(n1104) );
NAND2_X1 U795 ( .A1(KEYINPUT12), .A2(n1110), .ZN(n1108) );
OR2_X1 U796 ( .A1(n1111), .A2(n1106), .ZN(n1102) );
INV_X1 U797 ( .A(KEYINPUT12), .ZN(n1106) );
NAND3_X1 U798 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1100) );
NAND2_X1 U799 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NAND2_X1 U800 ( .A1(n1117), .A2(n1118), .ZN(n1113) );
INV_X1 U801 ( .A(KEYINPUT49), .ZN(n1118) );
NAND2_X1 U802 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
XNOR2_X1 U803 ( .A(KEYINPUT11), .B(G125), .ZN(n1119) );
NAND2_X1 U804 ( .A1(KEYINPUT49), .A2(n1121), .ZN(n1112) );
NAND2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
OR2_X1 U806 ( .A1(G125), .A2(KEYINPUT11), .ZN(n1123) );
NAND3_X1 U807 ( .A1(G125), .A2(n1120), .A3(KEYINPUT11), .ZN(n1122) );
INV_X1 U808 ( .A(n1115), .ZN(n1120) );
AND2_X1 U809 ( .A1(n1092), .A2(n1093), .ZN(n1094) );
XOR2_X1 U810 ( .A(n1039), .B(KEYINPUT60), .Z(n1093) );
NAND3_X1 U811 ( .A1(G953), .A2(n1124), .A3(KEYINPUT28), .ZN(n1086) );
XOR2_X1 U812 ( .A(KEYINPUT5), .B(n1125), .Z(n1124) );
NOR2_X1 U813 ( .A1(n1126), .A2(n1097), .ZN(n1125) );
XOR2_X1 U814 ( .A(n1127), .B(n1128), .Z(G69) );
NOR2_X1 U815 ( .A1(n1129), .A2(n1092), .ZN(n1128) );
NOR2_X1 U816 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U817 ( .A1(n1132), .A2(n1133), .ZN(n1127) );
NAND2_X1 U818 ( .A1(n1134), .A2(n1092), .ZN(n1133) );
XNOR2_X1 U819 ( .A(n1037), .B(n1135), .ZN(n1134) );
NAND3_X1 U820 ( .A1(G898), .A2(n1135), .A3(G953), .ZN(n1132) );
NOR2_X1 U821 ( .A1(n1136), .A2(n1137), .ZN(G66) );
XOR2_X1 U822 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U823 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NOR2_X1 U824 ( .A1(n1136), .A2(n1142), .ZN(G63) );
XOR2_X1 U825 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U826 ( .A1(n1145), .A2(KEYINPUT20), .ZN(n1144) );
NAND3_X1 U827 ( .A1(n1146), .A2(n1147), .A3(G478), .ZN(n1143) );
XNOR2_X1 U828 ( .A(KEYINPUT6), .B(n1148), .ZN(n1146) );
NOR2_X1 U829 ( .A1(n1136), .A2(n1149), .ZN(G60) );
XOR2_X1 U830 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U831 ( .A1(n1140), .A2(G475), .ZN(n1150) );
XNOR2_X1 U832 ( .A(n1152), .B(n1153), .ZN(G6) );
NOR2_X1 U833 ( .A1(n1070), .A2(n1154), .ZN(n1153) );
NOR2_X1 U834 ( .A1(n1136), .A2(n1155), .ZN(G57) );
XOR2_X1 U835 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U836 ( .A(n1158), .B(n1159), .Z(n1157) );
XNOR2_X1 U837 ( .A(n1160), .B(n1161), .ZN(n1156) );
XNOR2_X1 U838 ( .A(KEYINPUT57), .B(n1162), .ZN(n1161) );
NOR3_X1 U839 ( .A1(n1163), .A2(KEYINPUT39), .A3(n1164), .ZN(n1162) );
NOR2_X1 U840 ( .A1(n1136), .A2(n1165), .ZN(G54) );
XOR2_X1 U841 ( .A(n1166), .B(n1167), .Z(n1165) );
XOR2_X1 U842 ( .A(n1168), .B(n1169), .Z(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
NAND2_X1 U844 ( .A1(KEYINPUT2), .A2(n1172), .ZN(n1170) );
XNOR2_X1 U845 ( .A(n1173), .B(G110), .ZN(n1168) );
XOR2_X1 U846 ( .A(n1174), .B(n1098), .Z(n1166) );
XOR2_X1 U847 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U848 ( .A1(n1140), .A2(G469), .ZN(n1175) );
NOR2_X1 U849 ( .A1(n1136), .A2(n1177), .ZN(G51) );
XNOR2_X1 U850 ( .A(n1178), .B(n1179), .ZN(n1177) );
XOR2_X1 U851 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U852 ( .A1(n1140), .A2(n1182), .ZN(n1180) );
INV_X1 U853 ( .A(n1163), .ZN(n1140) );
NAND2_X1 U854 ( .A1(G902), .A2(n1147), .ZN(n1163) );
NAND2_X1 U855 ( .A1(n1039), .A2(n1037), .ZN(n1147) );
AND4_X1 U856 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1037) );
NOR4_X1 U857 ( .A1(n1187), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1186) );
NOR2_X1 U858 ( .A1(n1031), .A2(n1191), .ZN(n1185) );
INV_X1 U859 ( .A(n1192), .ZN(n1191) );
AND3_X1 U860 ( .A1(n1044), .A2(n1193), .A3(n1052), .ZN(n1031) );
NAND2_X1 U861 ( .A1(n1194), .A2(n1195), .ZN(n1183) );
XNOR2_X1 U862 ( .A(KEYINPUT3), .B(n1154), .ZN(n1195) );
NAND4_X1 U863 ( .A1(n1051), .A2(n1044), .A3(n1059), .A4(n1196), .ZN(n1154) );
AND2_X1 U864 ( .A1(n1197), .A2(n1198), .ZN(n1039) );
NOR4_X1 U865 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1198) );
NOR4_X1 U866 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1197) );
NOR3_X1 U867 ( .A1(n1207), .A2(n1208), .A3(n1209), .ZN(n1206) );
XNOR2_X1 U868 ( .A(n1052), .B(KEYINPUT27), .ZN(n1208) );
XOR2_X1 U869 ( .A(KEYINPUT8), .B(n1046), .Z(n1207) );
NOR2_X1 U870 ( .A1(n1092), .A2(G952), .ZN(n1136) );
XOR2_X1 U871 ( .A(n1202), .B(n1210), .Z(G48) );
XOR2_X1 U872 ( .A(KEYINPUT38), .B(G146), .Z(n1210) );
AND3_X1 U873 ( .A1(n1211), .A2(n1194), .A3(n1051), .ZN(n1202) );
XOR2_X1 U874 ( .A(G143), .B(n1201), .Z(G45) );
NOR3_X1 U875 ( .A1(n1212), .A2(n1070), .A3(n1209), .ZN(n1201) );
XOR2_X1 U876 ( .A(n1213), .B(G140), .Z(G42) );
NAND2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND3_X1 U878 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1215) );
INV_X1 U879 ( .A(KEYINPUT15), .ZN(n1218) );
NAND2_X1 U880 ( .A1(n1203), .A2(KEYINPUT15), .ZN(n1214) );
AND2_X1 U881 ( .A1(n1066), .A2(n1216), .ZN(n1203) );
XNOR2_X1 U882 ( .A(n1110), .B(n1205), .ZN(G39) );
AND3_X1 U883 ( .A1(n1046), .A2(n1211), .A3(n1053), .ZN(n1205) );
XNOR2_X1 U884 ( .A(G134), .B(n1219), .ZN(G36) );
NAND3_X1 U885 ( .A1(n1046), .A2(n1052), .A3(n1220), .ZN(n1219) );
INV_X1 U886 ( .A(n1209), .ZN(n1220) );
NAND3_X1 U887 ( .A1(n1059), .A2(n1221), .A3(n1064), .ZN(n1209) );
XOR2_X1 U888 ( .A(n1200), .B(n1222), .Z(G33) );
XNOR2_X1 U889 ( .A(KEYINPUT19), .B(n1107), .ZN(n1222) );
AND2_X1 U890 ( .A1(n1064), .A2(n1216), .ZN(n1200) );
AND4_X1 U891 ( .A1(n1046), .A2(n1051), .A3(n1059), .A4(n1221), .ZN(n1216) );
NOR2_X1 U892 ( .A1(n1072), .A2(n1077), .ZN(n1046) );
INV_X1 U893 ( .A(n1071), .ZN(n1077) );
XOR2_X1 U894 ( .A(n1199), .B(n1223), .Z(G30) );
NOR2_X1 U895 ( .A1(KEYINPUT43), .A2(n1224), .ZN(n1223) );
AND3_X1 U896 ( .A1(n1052), .A2(n1194), .A3(n1211), .ZN(n1199) );
AND4_X1 U897 ( .A1(n1059), .A2(n1225), .A3(n1226), .A4(n1221), .ZN(n1211) );
XNOR2_X1 U898 ( .A(G101), .B(n1227), .ZN(G3) );
NAND2_X1 U899 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
NAND2_X1 U900 ( .A1(KEYINPUT46), .A2(n1190), .ZN(n1229) );
OR2_X1 U901 ( .A1(KEYINPUT47), .A2(n1190), .ZN(n1228) );
AND3_X1 U902 ( .A1(n1064), .A2(n1193), .A3(n1053), .ZN(n1190) );
XNOR2_X1 U903 ( .A(n1204), .B(n1230), .ZN(G27) );
XNOR2_X1 U904 ( .A(KEYINPUT53), .B(n1116), .ZN(n1230) );
AND4_X1 U905 ( .A1(n1066), .A2(n1051), .A3(n1231), .A4(n1049), .ZN(n1204) );
AND2_X1 U906 ( .A1(n1221), .A2(n1194), .ZN(n1231) );
NAND2_X1 U907 ( .A1(n1073), .A2(n1232), .ZN(n1221) );
NAND4_X1 U908 ( .A1(G953), .A2(G902), .A3(n1233), .A4(n1097), .ZN(n1232) );
INV_X1 U909 ( .A(G900), .ZN(n1097) );
XOR2_X1 U910 ( .A(n1234), .B(G122), .Z(G24) );
NAND2_X1 U911 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND4_X1 U912 ( .A1(n1044), .A2(n1212), .A3(n1237), .A4(n1238), .ZN(n1236) );
INV_X1 U913 ( .A(KEYINPUT56), .ZN(n1238) );
NAND2_X1 U914 ( .A1(n1189), .A2(KEYINPUT56), .ZN(n1235) );
NOR3_X1 U915 ( .A1(n1212), .A2(n1080), .A3(n1239), .ZN(n1189) );
INV_X1 U916 ( .A(n1044), .ZN(n1080) );
NOR2_X1 U917 ( .A1(n1226), .A2(n1225), .ZN(n1044) );
NAND2_X1 U918 ( .A1(n1240), .A2(n1241), .ZN(n1212) );
XNOR2_X1 U919 ( .A(G119), .B(n1184), .ZN(G21) );
NAND4_X1 U920 ( .A1(n1237), .A2(n1053), .A3(n1225), .A4(n1226), .ZN(n1184) );
XNOR2_X1 U921 ( .A(n1188), .B(n1242), .ZN(G18) );
NAND2_X1 U922 ( .A1(G116), .A2(n1243), .ZN(n1242) );
XOR2_X1 U923 ( .A(KEYINPUT50), .B(KEYINPUT22), .Z(n1243) );
AND3_X1 U924 ( .A1(n1064), .A2(n1052), .A3(n1237), .ZN(n1188) );
NOR2_X1 U925 ( .A1(n1241), .A2(n1244), .ZN(n1052) );
XNOR2_X1 U926 ( .A(G113), .B(n1192), .ZN(G15) );
NAND3_X1 U927 ( .A1(n1064), .A2(n1051), .A3(n1237), .ZN(n1192) );
INV_X1 U928 ( .A(n1239), .ZN(n1237) );
NAND3_X1 U929 ( .A1(n1194), .A2(n1196), .A3(n1049), .ZN(n1239) );
NOR2_X1 U930 ( .A1(n1245), .A2(n1057), .ZN(n1049) );
AND2_X1 U931 ( .A1(n1244), .A2(n1241), .ZN(n1051) );
NOR2_X1 U932 ( .A1(n1225), .A2(n1246), .ZN(n1064) );
XOR2_X1 U933 ( .A(n1247), .B(n1187), .Z(G12) );
AND3_X1 U934 ( .A1(n1066), .A2(n1193), .A3(n1053), .ZN(n1187) );
NOR2_X1 U935 ( .A1(n1241), .A2(n1240), .ZN(n1053) );
INV_X1 U936 ( .A(n1244), .ZN(n1240) );
XNOR2_X1 U937 ( .A(n1248), .B(n1085), .ZN(n1244) );
NOR2_X1 U938 ( .A1(n1145), .A2(G902), .ZN(n1085) );
AND2_X1 U939 ( .A1(n1249), .A2(n1250), .ZN(n1145) );
NAND3_X1 U940 ( .A1(n1251), .A2(n1252), .A3(G217), .ZN(n1250) );
XOR2_X1 U941 ( .A(KEYINPUT35), .B(n1253), .Z(n1252) );
NAND2_X1 U942 ( .A1(n1253), .A2(n1254), .ZN(n1249) );
NAND2_X1 U943 ( .A1(G217), .A2(n1251), .ZN(n1254) );
XNOR2_X1 U944 ( .A(n1255), .B(n1256), .ZN(n1253) );
XOR2_X1 U945 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U946 ( .A(G107), .B(G143), .ZN(n1258) );
NAND2_X1 U947 ( .A1(KEYINPUT21), .A2(n1224), .ZN(n1257) );
XNOR2_X1 U948 ( .A(n1259), .B(n1260), .ZN(n1255) );
NAND2_X1 U949 ( .A1(KEYINPUT51), .A2(n1109), .ZN(n1260) );
NAND2_X1 U950 ( .A1(KEYINPUT17), .A2(n1261), .ZN(n1259) );
NAND2_X1 U951 ( .A1(KEYINPUT32), .A2(n1262), .ZN(n1248) );
INV_X1 U952 ( .A(G478), .ZN(n1262) );
NAND2_X1 U953 ( .A1(n1084), .A2(n1263), .ZN(n1241) );
NAND2_X1 U954 ( .A1(G475), .A2(n1083), .ZN(n1263) );
OR2_X1 U955 ( .A1(n1083), .A2(G475), .ZN(n1084) );
NAND2_X1 U956 ( .A1(n1151), .A2(n1148), .ZN(n1083) );
AND3_X1 U957 ( .A1(n1264), .A2(n1265), .A3(n1266), .ZN(n1151) );
OR2_X1 U958 ( .A1(n1267), .A2(KEYINPUT4), .ZN(n1266) );
OR3_X1 U959 ( .A1(n1268), .A2(n1269), .A3(n1270), .ZN(n1265) );
INV_X1 U960 ( .A(KEYINPUT4), .ZN(n1268) );
NAND2_X1 U961 ( .A1(n1270), .A2(n1269), .ZN(n1264) );
NAND2_X1 U962 ( .A1(KEYINPUT42), .A2(n1267), .ZN(n1269) );
NAND2_X1 U963 ( .A1(n1271), .A2(n1272), .ZN(n1267) );
NAND2_X1 U964 ( .A1(n1273), .A2(n1152), .ZN(n1272) );
XOR2_X1 U965 ( .A(KEYINPUT26), .B(n1274), .Z(n1271) );
NOR2_X1 U966 ( .A1(n1273), .A2(n1152), .ZN(n1274) );
AND2_X1 U967 ( .A1(n1275), .A2(n1276), .ZN(n1273) );
NAND2_X1 U968 ( .A1(G122), .A2(n1277), .ZN(n1276) );
XOR2_X1 U969 ( .A(n1278), .B(KEYINPUT55), .Z(n1275) );
OR2_X1 U970 ( .A1(n1277), .A2(G122), .ZN(n1278) );
XNOR2_X1 U971 ( .A(n1279), .B(n1280), .ZN(n1270) );
XNOR2_X1 U972 ( .A(G131), .B(n1281), .ZN(n1280) );
NAND2_X1 U973 ( .A1(KEYINPUT18), .A2(G146), .ZN(n1281) );
XOR2_X1 U974 ( .A(n1282), .B(n1283), .Z(n1279) );
NAND2_X1 U975 ( .A1(n1284), .A2(n1285), .ZN(n1282) );
NAND4_X1 U976 ( .A1(G214), .A2(G143), .A3(n1286), .A4(n1092), .ZN(n1285) );
NAND2_X1 U977 ( .A1(n1287), .A2(n1288), .ZN(n1284) );
NAND3_X1 U978 ( .A1(n1286), .A2(n1092), .A3(G214), .ZN(n1288) );
XNOR2_X1 U979 ( .A(G143), .B(KEYINPUT45), .ZN(n1287) );
AND3_X1 U980 ( .A1(n1194), .A2(n1196), .A3(n1059), .ZN(n1193) );
NOR2_X1 U981 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
AND2_X1 U982 ( .A1(G221), .A2(n1289), .ZN(n1057) );
INV_X1 U983 ( .A(n1245), .ZN(n1058) );
XNOR2_X1 U984 ( .A(n1290), .B(G469), .ZN(n1245) );
NAND2_X1 U985 ( .A1(n1291), .A2(n1148), .ZN(n1290) );
XOR2_X1 U986 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U987 ( .A(n1171), .B(n1294), .ZN(n1293) );
XNOR2_X1 U988 ( .A(n1295), .B(n1296), .ZN(n1294) );
NAND2_X1 U989 ( .A1(KEYINPUT58), .A2(n1297), .ZN(n1296) );
NAND2_X1 U990 ( .A1(KEYINPUT59), .A2(n1173), .ZN(n1295) );
NOR2_X1 U991 ( .A1(n1126), .A2(G953), .ZN(n1171) );
INV_X1 U992 ( .A(G227), .ZN(n1126) );
XNOR2_X1 U993 ( .A(n1172), .B(n1298), .ZN(n1292) );
XNOR2_X1 U994 ( .A(n1299), .B(n1176), .ZN(n1298) );
XNOR2_X1 U995 ( .A(n1300), .B(n1301), .ZN(n1176) );
NAND2_X1 U996 ( .A1(KEYINPUT1), .A2(n1302), .ZN(n1300) );
NAND2_X1 U997 ( .A1(KEYINPUT63), .A2(n1098), .ZN(n1299) );
XNOR2_X1 U998 ( .A(n1303), .B(n1304), .ZN(n1098) );
XNOR2_X1 U999 ( .A(G146), .B(n1224), .ZN(n1304) );
NAND2_X1 U1000 ( .A1(KEYINPUT16), .A2(n1305), .ZN(n1303) );
XOR2_X1 U1001 ( .A(n1115), .B(KEYINPUT44), .Z(n1172) );
NAND2_X1 U1002 ( .A1(n1073), .A2(n1306), .ZN(n1196) );
NAND4_X1 U1003 ( .A1(G953), .A2(G902), .A3(n1233), .A4(n1131), .ZN(n1306) );
INV_X1 U1004 ( .A(G898), .ZN(n1131) );
NAND3_X1 U1005 ( .A1(n1233), .A2(n1092), .A3(G952), .ZN(n1073) );
NAND2_X1 U1006 ( .A1(G237), .A2(G234), .ZN(n1233) );
INV_X1 U1007 ( .A(n1070), .ZN(n1194) );
NAND2_X1 U1008 ( .A1(n1307), .A2(n1071), .ZN(n1070) );
NAND2_X1 U1009 ( .A1(G214), .A2(n1308), .ZN(n1071) );
XNOR2_X1 U1010 ( .A(KEYINPUT34), .B(n1309), .ZN(n1307) );
INV_X1 U1011 ( .A(n1072), .ZN(n1309) );
XNOR2_X1 U1012 ( .A(n1310), .B(n1182), .ZN(n1072) );
AND2_X1 U1013 ( .A1(G210), .A2(n1308), .ZN(n1182) );
NAND2_X1 U1014 ( .A1(n1286), .A2(n1148), .ZN(n1308) );
NAND2_X1 U1015 ( .A1(n1311), .A2(n1148), .ZN(n1310) );
XOR2_X1 U1016 ( .A(n1312), .B(n1181), .Z(n1311) );
XNOR2_X1 U1017 ( .A(n1160), .B(n1313), .ZN(n1181) );
XNOR2_X1 U1018 ( .A(n1116), .B(n1314), .ZN(n1313) );
NOR2_X1 U1019 ( .A1(G953), .A2(n1130), .ZN(n1314) );
INV_X1 U1020 ( .A(G224), .ZN(n1130) );
NAND2_X1 U1021 ( .A1(KEYINPUT41), .A2(n1178), .ZN(n1312) );
INV_X1 U1022 ( .A(n1135), .ZN(n1178) );
XNOR2_X1 U1023 ( .A(n1315), .B(n1316), .ZN(n1135) );
XOR2_X1 U1024 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1025 ( .A(n1302), .B(n1261), .Z(n1318) );
XOR2_X1 U1026 ( .A(G116), .B(G122), .Z(n1261) );
XNOR2_X1 U1027 ( .A(n1319), .B(KEYINPUT9), .ZN(n1302) );
INV_X1 U1028 ( .A(G101), .ZN(n1319) );
XOR2_X1 U1029 ( .A(n1320), .B(n1301), .Z(n1317) );
XNOR2_X1 U1030 ( .A(G107), .B(n1152), .ZN(n1301) );
INV_X1 U1031 ( .A(G104), .ZN(n1152) );
NOR2_X1 U1032 ( .A1(KEYINPUT14), .A2(n1297), .ZN(n1320) );
XOR2_X1 U1033 ( .A(n1321), .B(n1322), .Z(n1315) );
XNOR2_X1 U1034 ( .A(n1323), .B(G113), .ZN(n1322) );
XNOR2_X1 U1035 ( .A(KEYINPUT31), .B(KEYINPUT0), .ZN(n1321) );
INV_X1 U1036 ( .A(n1217), .ZN(n1066) );
NAND2_X1 U1037 ( .A1(n1246), .A2(n1225), .ZN(n1217) );
XNOR2_X1 U1038 ( .A(n1324), .B(n1141), .ZN(n1225) );
AND2_X1 U1039 ( .A1(G217), .A2(n1289), .ZN(n1141) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1148), .ZN(n1289) );
NAND2_X1 U1041 ( .A1(n1139), .A2(n1148), .ZN(n1324) );
XNOR2_X1 U1042 ( .A(n1325), .B(n1326), .ZN(n1139) );
XOR2_X1 U1043 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1044 ( .A(n1297), .B(n1329), .ZN(n1328) );
NOR2_X1 U1045 ( .A1(KEYINPUT10), .A2(n1330), .ZN(n1329) );
XOR2_X1 U1046 ( .A(n1331), .B(G146), .Z(n1330) );
NAND2_X1 U1047 ( .A1(KEYINPUT33), .A2(n1283), .ZN(n1331) );
XNOR2_X1 U1048 ( .A(n1116), .B(n1115), .ZN(n1283) );
XOR2_X1 U1049 ( .A(G140), .B(KEYINPUT48), .Z(n1115) );
INV_X1 U1050 ( .A(G125), .ZN(n1116) );
AND2_X1 U1051 ( .A1(n1251), .A2(G221), .ZN(n1327) );
AND2_X1 U1052 ( .A1(G234), .A2(n1092), .ZN(n1251) );
XNOR2_X1 U1053 ( .A(G119), .B(n1332), .ZN(n1325) );
XNOR2_X1 U1054 ( .A(n1110), .B(G128), .ZN(n1332) );
INV_X1 U1055 ( .A(n1226), .ZN(n1246) );
XOR2_X1 U1056 ( .A(n1333), .B(n1164), .Z(n1226) );
INV_X1 U1057 ( .A(G472), .ZN(n1164) );
NAND2_X1 U1058 ( .A1(n1334), .A2(n1148), .ZN(n1333) );
INV_X1 U1059 ( .A(G902), .ZN(n1148) );
XNOR2_X1 U1060 ( .A(n1159), .B(n1335), .ZN(n1334) );
XNOR2_X1 U1061 ( .A(n1158), .B(n1336), .ZN(n1335) );
NOR2_X1 U1062 ( .A1(KEYINPUT23), .A2(n1160), .ZN(n1336) );
XOR2_X1 U1063 ( .A(n1337), .B(n1305), .Z(n1160) );
XNOR2_X1 U1064 ( .A(G143), .B(KEYINPUT62), .ZN(n1305) );
XOR2_X1 U1065 ( .A(n1338), .B(G146), .Z(n1337) );
NAND2_X1 U1066 ( .A1(KEYINPUT24), .A2(n1224), .ZN(n1338) );
INV_X1 U1067 ( .A(G128), .ZN(n1224) );
XNOR2_X1 U1068 ( .A(n1339), .B(n1340), .ZN(n1158) );
NOR2_X1 U1069 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1070 ( .A(KEYINPUT61), .B(n1343), .Z(n1342) );
NOR2_X1 U1071 ( .A1(G116), .A2(n1323), .ZN(n1343) );
AND2_X1 U1072 ( .A1(n1323), .A2(G116), .ZN(n1341) );
INV_X1 U1073 ( .A(G119), .ZN(n1323) );
XNOR2_X1 U1074 ( .A(n1173), .B(n1344), .ZN(n1339) );
NOR2_X1 U1075 ( .A1(KEYINPUT40), .A2(n1277), .ZN(n1344) );
INV_X1 U1076 ( .A(G113), .ZN(n1277) );
AND3_X1 U1077 ( .A1(n1103), .A2(n1111), .A3(n1345), .ZN(n1173) );
NAND3_X1 U1078 ( .A1(G131), .A2(n1109), .A3(G137), .ZN(n1345) );
INV_X1 U1079 ( .A(G134), .ZN(n1109) );
NAND2_X1 U1080 ( .A1(n1346), .A2(n1110), .ZN(n1111) );
INV_X1 U1081 ( .A(G137), .ZN(n1110) );
XNOR2_X1 U1082 ( .A(G131), .B(G134), .ZN(n1346) );
NAND3_X1 U1083 ( .A1(G134), .A2(n1107), .A3(G137), .ZN(n1103) );
INV_X1 U1084 ( .A(G131), .ZN(n1107) );
XOR2_X1 U1085 ( .A(G101), .B(n1347), .Z(n1159) );
AND3_X1 U1086 ( .A1(G210), .A2(n1092), .A3(n1286), .ZN(n1347) );
INV_X1 U1087 ( .A(G237), .ZN(n1286) );
INV_X1 U1088 ( .A(G953), .ZN(n1092) );
NAND2_X1 U1089 ( .A1(KEYINPUT37), .A2(n1297), .ZN(n1247) );
INV_X1 U1090 ( .A(G110), .ZN(n1297) );
endmodule


