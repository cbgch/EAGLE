//Key = 0101001011011101001111000110011110100101000010110101110011011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;

XNOR2_X1 U788 ( .A(G107), .B(n1083), .ZN(G9) );
NOR2_X1 U789 ( .A1(n1084), .A2(n1085), .ZN(G75) );
XOR2_X1 U790 ( .A(KEYINPUT16), .B(n1086), .Z(n1085) );
AND3_X1 U791 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1086) );
NOR4_X1 U792 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1089), .ZN(n1084) );
INV_X1 U793 ( .A(G952), .ZN(n1089) );
NOR2_X1 U794 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NOR3_X1 U795 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1093) );
NOR4_X1 U796 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
NOR2_X1 U797 ( .A1(n1102), .A2(n1103), .ZN(n1098) );
NOR2_X1 U798 ( .A1(n1104), .A2(n1105), .ZN(n1096) );
NOR2_X1 U799 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
NOR2_X1 U800 ( .A1(n1108), .A2(n1100), .ZN(n1107) );
NOR2_X1 U801 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U802 ( .A1(KEYINPUT22), .A2(n1111), .ZN(n1109) );
NOR2_X1 U803 ( .A1(n1112), .A2(n1099), .ZN(n1106) );
INV_X1 U804 ( .A(n1113), .ZN(n1099) );
NOR2_X1 U805 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NOR2_X1 U806 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
XNOR2_X1 U807 ( .A(n1118), .B(KEYINPUT46), .ZN(n1116) );
NOR2_X1 U808 ( .A1(n1119), .A2(n1120), .ZN(n1095) );
INV_X1 U809 ( .A(KEYINPUT22), .ZN(n1120) );
NOR3_X1 U810 ( .A1(n1105), .A2(n1100), .A3(n1111), .ZN(n1119) );
INV_X1 U811 ( .A(n1121), .ZN(n1105) );
NAND4_X1 U812 ( .A1(n1122), .A2(n1087), .A3(n1123), .A4(n1088), .ZN(n1090) );
NAND4_X1 U813 ( .A1(n1124), .A2(n1125), .A3(n1121), .A4(n1113), .ZN(n1123) );
XOR2_X1 U814 ( .A(n1126), .B(KEYINPUT21), .Z(n1125) );
NAND2_X1 U815 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U816 ( .A(n1129), .B(KEYINPUT49), .ZN(n1124) );
NAND2_X1 U817 ( .A1(n1130), .A2(n1131), .ZN(n1087) );
NOR4_X1 U818 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1131) );
XNOR2_X1 U819 ( .A(G469), .B(n1136), .ZN(n1135) );
NOR2_X1 U820 ( .A1(n1137), .A2(KEYINPUT45), .ZN(n1136) );
NOR2_X1 U821 ( .A1(n1138), .A2(n1139), .ZN(n1134) );
INV_X1 U822 ( .A(n1140), .ZN(n1132) );
NOR4_X1 U823 ( .A1(n1141), .A2(n1142), .A3(n1094), .A4(n1143), .ZN(n1130) );
XOR2_X1 U824 ( .A(n1144), .B(n1145), .Z(n1143) );
XNOR2_X1 U825 ( .A(KEYINPUT36), .B(n1146), .ZN(n1145) );
NOR3_X1 U826 ( .A1(n1147), .A2(KEYINPUT58), .A3(G902), .ZN(n1144) );
NAND4_X1 U827 ( .A1(n1121), .A2(n1129), .A3(n1113), .A4(n1148), .ZN(n1122) );
NOR2_X1 U828 ( .A1(n1101), .A2(n1149), .ZN(n1121) );
XOR2_X1 U829 ( .A(n1150), .B(n1151), .Z(G72) );
NOR2_X1 U830 ( .A1(n1152), .A2(n1088), .ZN(n1151) );
AND2_X1 U831 ( .A1(G227), .A2(G900), .ZN(n1152) );
NAND2_X1 U832 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
NAND2_X1 U833 ( .A1(n1155), .A2(n1088), .ZN(n1154) );
XOR2_X1 U834 ( .A(n1156), .B(n1157), .Z(n1155) );
OR3_X1 U835 ( .A1(n1158), .A2(n1157), .A3(n1088), .ZN(n1153) );
XNOR2_X1 U836 ( .A(n1159), .B(n1160), .ZN(n1157) );
XOR2_X1 U837 ( .A(G131), .B(n1161), .Z(n1160) );
XOR2_X1 U838 ( .A(KEYINPUT4), .B(G137), .Z(n1161) );
XOR2_X1 U839 ( .A(n1162), .B(n1163), .Z(n1159) );
XNOR2_X1 U840 ( .A(n1164), .B(n1165), .ZN(n1163) );
NOR2_X1 U841 ( .A1(KEYINPUT14), .A2(n1166), .ZN(n1165) );
XNOR2_X1 U842 ( .A(G134), .B(KEYINPUT9), .ZN(n1166) );
NAND2_X1 U843 ( .A1(KEYINPUT59), .A2(n1167), .ZN(n1164) );
INV_X1 U844 ( .A(n1168), .ZN(n1167) );
XOR2_X1 U845 ( .A(n1169), .B(n1170), .Z(G69) );
NOR2_X1 U846 ( .A1(n1171), .A2(n1088), .ZN(n1170) );
NOR2_X1 U847 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND2_X1 U848 ( .A1(n1174), .A2(n1175), .ZN(n1169) );
NAND3_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1175) );
NAND2_X1 U850 ( .A1(G953), .A2(n1173), .ZN(n1177) );
NAND2_X1 U851 ( .A1(n1179), .A2(n1088), .ZN(n1176) );
XOR2_X1 U852 ( .A(KEYINPUT15), .B(n1180), .Z(n1174) );
NOR3_X1 U853 ( .A1(n1178), .A2(G953), .A3(n1181), .ZN(n1180) );
INV_X1 U854 ( .A(n1179), .ZN(n1181) );
NAND3_X1 U855 ( .A1(n1182), .A2(n1183), .A3(n1184), .ZN(n1179) );
XOR2_X1 U856 ( .A(n1185), .B(KEYINPUT5), .Z(n1184) );
XNOR2_X1 U857 ( .A(KEYINPUT8), .B(n1186), .ZN(n1183) );
XNOR2_X1 U858 ( .A(n1187), .B(n1188), .ZN(n1178) );
XOR2_X1 U859 ( .A(KEYINPUT43), .B(n1189), .Z(n1188) );
NOR2_X1 U860 ( .A1(KEYINPUT41), .A2(n1190), .ZN(n1189) );
XNOR2_X1 U861 ( .A(n1191), .B(n1192), .ZN(n1187) );
NOR2_X1 U862 ( .A1(n1193), .A2(n1194), .ZN(G66) );
XOR2_X1 U863 ( .A(n1195), .B(n1196), .Z(n1194) );
NOR2_X1 U864 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
NOR2_X1 U865 ( .A1(n1193), .A2(n1199), .ZN(G63) );
XOR2_X1 U866 ( .A(n1200), .B(n1147), .Z(n1199) );
NOR2_X1 U867 ( .A1(n1146), .A2(n1198), .ZN(n1200) );
NOR2_X1 U868 ( .A1(n1193), .A2(n1201), .ZN(G60) );
XOR2_X1 U869 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U870 ( .A1(n1204), .A2(n1198), .ZN(n1202) );
XNOR2_X1 U871 ( .A(G104), .B(n1186), .ZN(G6) );
NOR2_X1 U872 ( .A1(n1193), .A2(n1205), .ZN(G57) );
XOR2_X1 U873 ( .A(n1206), .B(n1207), .Z(n1205) );
NOR2_X1 U874 ( .A1(KEYINPUT33), .A2(n1208), .ZN(n1207) );
XNOR2_X1 U875 ( .A(n1209), .B(n1210), .ZN(n1208) );
XOR2_X1 U876 ( .A(n1211), .B(n1212), .Z(n1210) );
NOR2_X1 U877 ( .A1(n1139), .A2(n1198), .ZN(n1212) );
NOR2_X1 U878 ( .A1(KEYINPUT23), .A2(n1213), .ZN(n1211) );
NOR3_X1 U879 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1206) );
NOR2_X1 U880 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
AND3_X1 U881 ( .A1(n1217), .A2(n1218), .A3(KEYINPUT51), .ZN(n1215) );
AND2_X1 U882 ( .A1(KEYINPUT53), .A2(n1219), .ZN(n1218) );
INV_X1 U883 ( .A(n1220), .ZN(n1217) );
NOR2_X1 U884 ( .A1(KEYINPUT51), .A2(n1219), .ZN(n1214) );
NOR2_X1 U885 ( .A1(n1193), .A2(n1221), .ZN(G54) );
XOR2_X1 U886 ( .A(n1222), .B(n1223), .Z(n1221) );
XOR2_X1 U887 ( .A(n1224), .B(n1225), .Z(n1222) );
NOR2_X1 U888 ( .A1(n1226), .A2(n1198), .ZN(n1225) );
NAND2_X1 U889 ( .A1(KEYINPUT12), .A2(n1227), .ZN(n1224) );
NOR2_X1 U890 ( .A1(n1193), .A2(n1228), .ZN(G51) );
XNOR2_X1 U891 ( .A(n1229), .B(n1230), .ZN(n1228) );
XNOR2_X1 U892 ( .A(n1231), .B(n1232), .ZN(n1230) );
NOR2_X1 U893 ( .A1(n1198), .A2(n1233), .ZN(n1231) );
XOR2_X1 U894 ( .A(KEYINPUT20), .B(n1234), .Z(n1233) );
NAND2_X1 U895 ( .A1(G902), .A2(n1091), .ZN(n1198) );
NAND4_X1 U896 ( .A1(n1156), .A2(n1182), .A3(n1186), .A4(n1185), .ZN(n1091) );
NAND3_X1 U897 ( .A1(n1235), .A2(n1113), .A3(n1103), .ZN(n1186) );
AND4_X1 U898 ( .A1(n1236), .A2(n1083), .A3(n1237), .A4(n1238), .ZN(n1182) );
NOR3_X1 U899 ( .A1(n1239), .A2(n1240), .A3(n1241), .ZN(n1238) );
NOR3_X1 U900 ( .A1(n1242), .A2(n1111), .A3(n1243), .ZN(n1241) );
XNOR2_X1 U901 ( .A(KEYINPUT13), .B(n1244), .ZN(n1242) );
NOR4_X1 U902 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1149), .ZN(n1240) );
INV_X1 U903 ( .A(n1248), .ZN(n1149) );
NOR2_X1 U904 ( .A1(n1249), .A2(n1250), .ZN(n1246) );
INV_X1 U905 ( .A(KEYINPUT38), .ZN(n1250) );
NOR3_X1 U906 ( .A1(n1251), .A2(n1252), .A3(n1148), .ZN(n1249) );
NOR2_X1 U907 ( .A1(KEYINPUT38), .A2(n1235), .ZN(n1245) );
NOR2_X1 U908 ( .A1(n1253), .A2(n1254), .ZN(n1239) );
INV_X1 U909 ( .A(n1255), .ZN(n1237) );
NAND3_X1 U910 ( .A1(n1102), .A2(n1113), .A3(n1235), .ZN(n1083) );
AND4_X1 U911 ( .A1(n1256), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1156) );
NOR4_X1 U912 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1259) );
NOR2_X1 U913 ( .A1(n1264), .A2(n1094), .ZN(n1263) );
NOR3_X1 U914 ( .A1(n1265), .A2(n1266), .A3(n1267), .ZN(n1264) );
NOR4_X1 U915 ( .A1(n1268), .A2(n1269), .A3(n1251), .A4(n1270), .ZN(n1261) );
AND2_X1 U916 ( .A1(n1268), .A2(n1271), .ZN(n1260) );
INV_X1 U917 ( .A(KEYINPUT27), .ZN(n1268) );
NOR2_X1 U918 ( .A1(n1088), .A2(G952), .ZN(n1193) );
XNOR2_X1 U919 ( .A(G146), .B(n1257), .ZN(G48) );
NAND3_X1 U920 ( .A1(n1103), .A2(n1148), .A3(n1272), .ZN(n1257) );
XOR2_X1 U921 ( .A(G143), .B(n1271), .Z(G45) );
NOR2_X1 U922 ( .A1(n1269), .A2(n1273), .ZN(n1271) );
NAND4_X1 U923 ( .A1(n1274), .A2(n1148), .A3(n1275), .A4(n1142), .ZN(n1269) );
NAND2_X1 U924 ( .A1(n1276), .A2(n1277), .ZN(G42) );
NAND3_X1 U925 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
XOR2_X1 U926 ( .A(n1281), .B(KEYINPUT7), .Z(n1276) );
NAND2_X1 U927 ( .A1(G140), .A2(n1282), .ZN(n1281) );
NAND2_X1 U928 ( .A1(n1280), .A2(n1278), .ZN(n1282) );
NAND2_X1 U929 ( .A1(n1283), .A2(n1284), .ZN(n1278) );
NAND2_X1 U930 ( .A1(n1267), .A2(n1285), .ZN(n1284) );
NOR3_X1 U931 ( .A1(n1286), .A2(n1273), .A3(n1247), .ZN(n1267) );
OR4_X1 U932 ( .A1(n1273), .A2(n1103), .A3(n1247), .A4(n1285), .ZN(n1283) );
INV_X1 U933 ( .A(KEYINPUT62), .ZN(n1285) );
XNOR2_X1 U934 ( .A(G137), .B(n1287), .ZN(G39) );
NAND2_X1 U935 ( .A1(n1288), .A2(n1265), .ZN(n1287) );
AND2_X1 U936 ( .A1(n1248), .A2(n1272), .ZN(n1265) );
XNOR2_X1 U937 ( .A(n1280), .B(KEYINPUT52), .ZN(n1288) );
XNOR2_X1 U938 ( .A(n1289), .B(n1290), .ZN(G36) );
NOR2_X1 U939 ( .A1(KEYINPUT42), .A2(n1291), .ZN(n1290) );
INV_X1 U940 ( .A(n1262), .ZN(n1291) );
NOR4_X1 U941 ( .A1(n1111), .A2(n1094), .A3(n1273), .A4(n1244), .ZN(n1262) );
XNOR2_X1 U942 ( .A(G131), .B(n1292), .ZN(G33) );
NAND2_X1 U943 ( .A1(n1280), .A2(n1293), .ZN(n1292) );
XOR2_X1 U944 ( .A(KEYINPUT0), .B(n1266), .Z(n1293) );
NOR3_X1 U945 ( .A1(n1286), .A2(n1273), .A3(n1111), .ZN(n1266) );
INV_X1 U946 ( .A(n1094), .ZN(n1280) );
NAND2_X1 U947 ( .A1(n1128), .A2(n1294), .ZN(n1094) );
NAND2_X1 U948 ( .A1(n1295), .A2(n1296), .ZN(G30) );
NAND2_X1 U949 ( .A1(G128), .A2(n1258), .ZN(n1296) );
XOR2_X1 U950 ( .A(n1297), .B(KEYINPUT63), .Z(n1295) );
OR2_X1 U951 ( .A1(n1258), .A2(G128), .ZN(n1297) );
NAND3_X1 U952 ( .A1(n1102), .A2(n1148), .A3(n1272), .ZN(n1258) );
NOR3_X1 U953 ( .A1(n1298), .A2(n1299), .A3(n1273), .ZN(n1272) );
NAND2_X1 U954 ( .A1(n1115), .A2(n1270), .ZN(n1273) );
INV_X1 U955 ( .A(n1251), .ZN(n1115) );
XNOR2_X1 U956 ( .A(n1219), .B(n1255), .ZN(G3) );
NOR2_X1 U957 ( .A1(n1300), .A2(n1111), .ZN(n1255) );
INV_X1 U958 ( .A(n1274), .ZN(n1111) );
XNOR2_X1 U959 ( .A(G125), .B(n1256), .ZN(G27) );
NAND3_X1 U960 ( .A1(n1110), .A2(n1129), .A3(n1301), .ZN(n1256) );
AND3_X1 U961 ( .A1(n1103), .A2(n1270), .A3(n1148), .ZN(n1301) );
NAND2_X1 U962 ( .A1(n1101), .A2(n1302), .ZN(n1270) );
NAND4_X1 U963 ( .A1(G953), .A2(G902), .A3(n1303), .A4(n1158), .ZN(n1302) );
INV_X1 U964 ( .A(G900), .ZN(n1158) );
XNOR2_X1 U965 ( .A(G122), .B(n1236), .ZN(G24) );
NAND4_X1 U966 ( .A1(n1304), .A2(n1113), .A3(n1275), .A4(n1142), .ZN(n1236) );
NOR2_X1 U967 ( .A1(n1305), .A2(n1141), .ZN(n1113) );
XNOR2_X1 U968 ( .A(n1306), .B(n1307), .ZN(G21) );
NOR2_X1 U969 ( .A1(n1308), .A2(n1253), .ZN(n1307) );
XOR2_X1 U970 ( .A(n1254), .B(KEYINPUT2), .Z(n1308) );
NAND3_X1 U971 ( .A1(n1248), .A2(n1129), .A3(n1309), .ZN(n1254) );
NOR3_X1 U972 ( .A1(n1298), .A2(n1252), .A3(n1299), .ZN(n1309) );
XNOR2_X1 U973 ( .A(n1310), .B(n1311), .ZN(G18) );
NOR3_X1 U974 ( .A1(n1243), .A2(n1312), .A3(n1244), .ZN(n1311) );
INV_X1 U975 ( .A(n1102), .ZN(n1244) );
NOR2_X1 U976 ( .A1(n1142), .A2(n1313), .ZN(n1102) );
XNOR2_X1 U977 ( .A(n1274), .B(KEYINPUT40), .ZN(n1312) );
INV_X1 U978 ( .A(n1304), .ZN(n1243) );
XNOR2_X1 U979 ( .A(G113), .B(n1185), .ZN(G15) );
NAND3_X1 U980 ( .A1(n1274), .A2(n1103), .A3(n1304), .ZN(n1185) );
NOR3_X1 U981 ( .A1(n1253), .A2(n1252), .A3(n1100), .ZN(n1304) );
INV_X1 U982 ( .A(n1129), .ZN(n1100) );
NOR2_X1 U983 ( .A1(n1118), .A2(n1133), .ZN(n1129) );
INV_X1 U984 ( .A(n1117), .ZN(n1133) );
INV_X1 U985 ( .A(n1286), .ZN(n1103) );
NAND2_X1 U986 ( .A1(n1313), .A2(n1314), .ZN(n1286) );
XOR2_X1 U987 ( .A(KEYINPUT35), .B(n1142), .Z(n1314) );
INV_X1 U988 ( .A(n1275), .ZN(n1313) );
NOR2_X1 U989 ( .A1(n1141), .A2(n1299), .ZN(n1274) );
INV_X1 U990 ( .A(n1305), .ZN(n1299) );
XOR2_X1 U991 ( .A(G110), .B(n1315), .Z(G12) );
NOR2_X1 U992 ( .A1(n1247), .A2(n1300), .ZN(n1315) );
NAND2_X1 U993 ( .A1(n1248), .A2(n1235), .ZN(n1300) );
NOR3_X1 U994 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1235) );
INV_X1 U995 ( .A(n1148), .ZN(n1253) );
NOR2_X1 U996 ( .A1(n1128), .A2(n1127), .ZN(n1148) );
INV_X1 U997 ( .A(n1294), .ZN(n1127) );
NAND2_X1 U998 ( .A1(G214), .A2(n1316), .ZN(n1294) );
XOR2_X1 U999 ( .A(n1317), .B(n1234), .Z(n1128) );
AND2_X1 U1000 ( .A1(G210), .A2(n1316), .ZN(n1234) );
NAND2_X1 U1001 ( .A1(n1318), .A2(n1319), .ZN(n1316) );
NAND3_X1 U1002 ( .A1(n1320), .A2(n1321), .A3(n1319), .ZN(n1317) );
NAND2_X1 U1003 ( .A1(n1322), .A2(n1232), .ZN(n1321) );
NAND2_X1 U1004 ( .A1(n1323), .A2(n1324), .ZN(n1322) );
NAND2_X1 U1005 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
INV_X1 U1006 ( .A(KEYINPUT24), .ZN(n1326) );
NAND2_X1 U1007 ( .A1(KEYINPUT24), .A2(n1229), .ZN(n1323) );
OR2_X1 U1008 ( .A1(n1232), .A2(n1325), .ZN(n1320) );
NAND2_X1 U1009 ( .A1(KEYINPUT25), .A2(n1229), .ZN(n1325) );
XNOR2_X1 U1010 ( .A(n1327), .B(n1328), .ZN(n1229) );
XNOR2_X1 U1011 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR2_X1 U1012 ( .A1(G953), .A2(n1172), .ZN(n1330) );
INV_X1 U1013 ( .A(G224), .ZN(n1172) );
INV_X1 U1014 ( .A(G125), .ZN(n1329) );
XOR2_X1 U1015 ( .A(n1331), .B(n1192), .Z(n1232) );
XNOR2_X1 U1016 ( .A(n1332), .B(n1333), .ZN(n1192) );
NOR2_X1 U1017 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1018 ( .A(KEYINPUT50), .B(n1336), .Z(n1335) );
NOR2_X1 U1019 ( .A1(G119), .A2(n1337), .ZN(n1336) );
AND2_X1 U1020 ( .A1(n1337), .A2(G119), .ZN(n1334) );
XOR2_X1 U1021 ( .A(G116), .B(KEYINPUT34), .Z(n1337) );
XOR2_X1 U1022 ( .A(n1338), .B(n1191), .Z(n1331) );
XNOR2_X1 U1023 ( .A(G110), .B(n1339), .ZN(n1191) );
NAND2_X1 U1024 ( .A1(KEYINPUT26), .A2(n1340), .ZN(n1338) );
INV_X1 U1025 ( .A(n1190), .ZN(n1340) );
XNOR2_X1 U1026 ( .A(n1341), .B(n1342), .ZN(n1190) );
NOR3_X1 U1027 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1342) );
AND2_X1 U1028 ( .A1(n1346), .A2(G107), .ZN(n1345) );
NOR3_X1 U1029 ( .A1(G107), .A2(KEYINPUT54), .A3(n1346), .ZN(n1344) );
NAND2_X1 U1030 ( .A1(KEYINPUT30), .A2(n1347), .ZN(n1346) );
AND2_X1 U1031 ( .A1(G104), .A2(KEYINPUT54), .ZN(n1343) );
NAND2_X1 U1032 ( .A1(KEYINPUT60), .A2(n1219), .ZN(n1341) );
AND2_X1 U1033 ( .A1(n1348), .A2(n1101), .ZN(n1252) );
NAND3_X1 U1034 ( .A1(n1303), .A2(n1088), .A3(G952), .ZN(n1101) );
NAND4_X1 U1035 ( .A1(G953), .A2(G902), .A3(n1303), .A4(n1173), .ZN(n1348) );
INV_X1 U1036 ( .A(G898), .ZN(n1173) );
NAND2_X1 U1037 ( .A1(G237), .A2(G234), .ZN(n1303) );
NAND2_X1 U1038 ( .A1(n1118), .A2(n1117), .ZN(n1251) );
NAND2_X1 U1039 ( .A1(G221), .A2(n1349), .ZN(n1117) );
XOR2_X1 U1040 ( .A(KEYINPUT47), .B(n1350), .Z(n1349) );
AND2_X1 U1041 ( .A1(n1319), .A2(G234), .ZN(n1350) );
XNOR2_X1 U1042 ( .A(n1137), .B(n1226), .ZN(n1118) );
INV_X1 U1043 ( .A(G469), .ZN(n1226) );
AND2_X1 U1044 ( .A1(n1351), .A2(n1319), .ZN(n1137) );
XOR2_X1 U1045 ( .A(n1223), .B(n1227), .Z(n1351) );
XNOR2_X1 U1046 ( .A(n1352), .B(n1353), .ZN(n1223) );
XOR2_X1 U1047 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1048 ( .A(G107), .B(n1219), .ZN(n1355) );
INV_X1 U1049 ( .A(G101), .ZN(n1219) );
XNOR2_X1 U1050 ( .A(n1279), .B(G110), .ZN(n1354) );
XOR2_X1 U1051 ( .A(n1162), .B(n1356), .Z(n1352) );
XOR2_X1 U1052 ( .A(n1357), .B(n1358), .Z(n1356) );
NAND2_X1 U1053 ( .A1(KEYINPUT1), .A2(G104), .ZN(n1358) );
NAND2_X1 U1054 ( .A1(n1359), .A2(n1088), .ZN(n1357) );
XOR2_X1 U1055 ( .A(KEYINPUT17), .B(G227), .Z(n1359) );
XOR2_X1 U1056 ( .A(n1360), .B(n1361), .Z(n1162) );
NAND2_X1 U1057 ( .A1(n1362), .A2(n1363), .ZN(n1360) );
NAND2_X1 U1058 ( .A1(G143), .A2(n1364), .ZN(n1363) );
XOR2_X1 U1059 ( .A(KEYINPUT3), .B(n1365), .Z(n1362) );
NOR2_X1 U1060 ( .A1(G143), .A2(n1364), .ZN(n1365) );
NOR2_X1 U1061 ( .A1(n1275), .A2(n1142), .ZN(n1248) );
XOR2_X1 U1062 ( .A(n1366), .B(n1204), .Z(n1142) );
INV_X1 U1063 ( .A(G475), .ZN(n1204) );
OR2_X1 U1064 ( .A1(n1203), .A2(G902), .ZN(n1366) );
XNOR2_X1 U1065 ( .A(n1367), .B(n1368), .ZN(n1203) );
XOR2_X1 U1066 ( .A(n1369), .B(n1370), .Z(n1368) );
AND3_X1 U1067 ( .A1(G214), .A2(n1088), .A3(n1318), .ZN(n1369) );
XOR2_X1 U1068 ( .A(n1371), .B(n1372), .Z(n1367) );
XOR2_X1 U1069 ( .A(G143), .B(G131), .Z(n1372) );
NAND3_X1 U1070 ( .A1(n1373), .A2(n1374), .A3(n1375), .ZN(n1371) );
OR2_X1 U1071 ( .A1(n1376), .A2(KEYINPUT37), .ZN(n1375) );
NAND3_X1 U1072 ( .A1(KEYINPUT37), .A2(n1377), .A3(n1347), .ZN(n1374) );
INV_X1 U1073 ( .A(G104), .ZN(n1347) );
INV_X1 U1074 ( .A(n1378), .ZN(n1377) );
NAND2_X1 U1075 ( .A1(G104), .A2(n1378), .ZN(n1373) );
NAND2_X1 U1076 ( .A1(KEYINPUT56), .A2(n1376), .ZN(n1378) );
XNOR2_X1 U1077 ( .A(G113), .B(n1339), .ZN(n1376) );
XOR2_X1 U1078 ( .A(n1379), .B(n1146), .Z(n1275) );
INV_X1 U1079 ( .A(G478), .ZN(n1146) );
OR2_X1 U1080 ( .A1(n1147), .A2(G902), .ZN(n1379) );
XNOR2_X1 U1081 ( .A(n1380), .B(n1381), .ZN(n1147) );
NOR2_X1 U1082 ( .A1(n1382), .A2(n1383), .ZN(n1381) );
INV_X1 U1083 ( .A(G217), .ZN(n1383) );
NAND2_X1 U1084 ( .A1(n1384), .A2(KEYINPUT39), .ZN(n1380) );
XOR2_X1 U1085 ( .A(n1385), .B(n1386), .Z(n1384) );
XNOR2_X1 U1086 ( .A(n1289), .B(n1387), .ZN(n1386) );
XOR2_X1 U1087 ( .A(KEYINPUT18), .B(G143), .Z(n1387) );
INV_X1 U1088 ( .A(G134), .ZN(n1289) );
XNOR2_X1 U1089 ( .A(n1361), .B(n1388), .ZN(n1385) );
XOR2_X1 U1090 ( .A(G107), .B(n1389), .Z(n1388) );
NOR4_X1 U1091 ( .A1(n1390), .A2(n1391), .A3(KEYINPUT61), .A4(n1392), .ZN(n1389) );
NOR2_X1 U1092 ( .A1(KEYINPUT31), .A2(n1310), .ZN(n1392) );
NOR2_X1 U1093 ( .A1(n1393), .A2(n1339), .ZN(n1391) );
AND2_X1 U1094 ( .A1(n1310), .A2(KEYINPUT57), .ZN(n1393) );
AND4_X1 U1095 ( .A1(n1339), .A2(KEYINPUT31), .A3(n1310), .A4(KEYINPUT57), .ZN(n1390) );
INV_X1 U1096 ( .A(G122), .ZN(n1339) );
INV_X1 U1097 ( .A(n1110), .ZN(n1247) );
NOR2_X1 U1098 ( .A1(n1305), .A2(n1298), .ZN(n1110) );
INV_X1 U1099 ( .A(n1141), .ZN(n1298) );
XOR2_X1 U1100 ( .A(n1394), .B(n1197), .Z(n1141) );
NAND2_X1 U1101 ( .A1(G217), .A2(n1395), .ZN(n1197) );
NAND2_X1 U1102 ( .A1(G234), .A2(n1319), .ZN(n1395) );
OR2_X1 U1103 ( .A1(n1196), .A2(G902), .ZN(n1394) );
XNOR2_X1 U1104 ( .A(n1396), .B(n1397), .ZN(n1196) );
XOR2_X1 U1105 ( .A(n1398), .B(n1370), .Z(n1397) );
XNOR2_X1 U1106 ( .A(n1364), .B(n1168), .ZN(n1370) );
XNOR2_X1 U1107 ( .A(G125), .B(n1279), .ZN(n1168) );
INV_X1 U1108 ( .A(G140), .ZN(n1279) );
NOR2_X1 U1109 ( .A1(n1399), .A2(n1382), .ZN(n1398) );
NAND2_X1 U1110 ( .A1(G234), .A2(n1088), .ZN(n1382) );
INV_X1 U1111 ( .A(G221), .ZN(n1399) );
XOR2_X1 U1112 ( .A(n1400), .B(n1401), .Z(n1396) );
XOR2_X1 U1113 ( .A(G137), .B(G110), .Z(n1401) );
NAND2_X1 U1114 ( .A1(n1402), .A2(n1403), .ZN(n1400) );
NAND2_X1 U1115 ( .A1(G119), .A2(n1361), .ZN(n1403) );
XOR2_X1 U1116 ( .A(KEYINPUT11), .B(n1404), .Z(n1402) );
NOR2_X1 U1117 ( .A1(G119), .A2(n1361), .ZN(n1404) );
NAND3_X1 U1118 ( .A1(n1405), .A2(n1406), .A3(n1140), .ZN(n1305) );
NAND2_X1 U1119 ( .A1(n1138), .A2(n1139), .ZN(n1140) );
NAND2_X1 U1120 ( .A1(KEYINPUT28), .A2(n1139), .ZN(n1406) );
OR3_X1 U1121 ( .A1(n1138), .A2(KEYINPUT28), .A3(n1139), .ZN(n1405) );
INV_X1 U1122 ( .A(G472), .ZN(n1139) );
AND2_X1 U1123 ( .A1(n1407), .A2(n1319), .ZN(n1138) );
INV_X1 U1124 ( .A(G902), .ZN(n1319) );
XOR2_X1 U1125 ( .A(n1408), .B(n1409), .Z(n1407) );
XNOR2_X1 U1126 ( .A(G101), .B(n1220), .ZN(n1409) );
NAND3_X1 U1127 ( .A1(n1318), .A2(n1088), .A3(n1410), .ZN(n1220) );
XOR2_X1 U1128 ( .A(KEYINPUT48), .B(G210), .Z(n1410) );
INV_X1 U1129 ( .A(G953), .ZN(n1088) );
INV_X1 U1130 ( .A(G237), .ZN(n1318) );
XNOR2_X1 U1131 ( .A(n1411), .B(n1412), .ZN(n1408) );
INV_X1 U1132 ( .A(n1209), .ZN(n1412) );
XNOR2_X1 U1133 ( .A(n1413), .B(n1414), .ZN(n1209) );
XNOR2_X1 U1134 ( .A(KEYINPUT29), .B(n1310), .ZN(n1414) );
INV_X1 U1135 ( .A(G116), .ZN(n1310) );
XNOR2_X1 U1136 ( .A(n1415), .B(n1332), .ZN(n1413) );
INV_X1 U1137 ( .A(G113), .ZN(n1332) );
NAND2_X1 U1138 ( .A1(KEYINPUT44), .A2(n1306), .ZN(n1415) );
INV_X1 U1139 ( .A(G119), .ZN(n1306) );
NAND3_X1 U1140 ( .A1(n1416), .A2(n1417), .A3(KEYINPUT19), .ZN(n1411) );
OR2_X1 U1141 ( .A1(n1213), .A2(KEYINPUT10), .ZN(n1417) );
XNOR2_X1 U1142 ( .A(n1327), .B(n1227), .ZN(n1213) );
NAND3_X1 U1143 ( .A1(n1227), .A2(n1327), .A3(KEYINPUT10), .ZN(n1416) );
XOR2_X1 U1144 ( .A(n1418), .B(n1361), .Z(n1327) );
XOR2_X1 U1145 ( .A(G128), .B(KEYINPUT6), .Z(n1361) );
XNOR2_X1 U1146 ( .A(n1419), .B(n1364), .ZN(n1418) );
INV_X1 U1147 ( .A(G146), .ZN(n1364) );
NAND2_X1 U1148 ( .A1(KEYINPUT32), .A2(G143), .ZN(n1419) );
XOR2_X1 U1149 ( .A(n1420), .B(n1421), .Z(n1227) );
NOR2_X1 U1150 ( .A1(KEYINPUT55), .A2(G131), .ZN(n1421) );
XNOR2_X1 U1151 ( .A(G134), .B(G137), .ZN(n1420) );
endmodule


