//Key = 1000101110110110100000001000011110100101001000100000010000000110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372;

XNOR2_X1 U766 ( .A(G107), .B(n1050), .ZN(G9) );
NAND3_X1 U767 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n1050) );
XNOR2_X1 U768 ( .A(n1054), .B(KEYINPUT33), .ZN(n1053) );
NOR2_X1 U769 ( .A1(n1055), .A2(n1056), .ZN(G75) );
NOR4_X1 U770 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR2_X1 U771 ( .A1(n1061), .A2(n1062), .ZN(n1059) );
NOR3_X1 U772 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NOR2_X1 U773 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U774 ( .A(KEYINPUT2), .ZN(n1067) );
NOR2_X1 U775 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NOR4_X1 U776 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1064) );
NOR2_X1 U777 ( .A1(n1074), .A2(n1075), .ZN(n1070) );
NOR2_X1 U778 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NOR2_X1 U779 ( .A1(n1078), .A2(n1069), .ZN(n1063) );
INV_X1 U780 ( .A(n1079), .ZN(n1069) );
NOR4_X1 U781 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1078) );
NOR2_X1 U782 ( .A1(n1071), .A2(n1084), .ZN(n1083) );
NOR2_X1 U783 ( .A1(KEYINPUT2), .A2(n1068), .ZN(n1082) );
INV_X1 U784 ( .A(n1052), .ZN(n1068) );
NOR2_X1 U785 ( .A1(n1085), .A2(n1071), .ZN(n1052) );
INV_X1 U786 ( .A(n1086), .ZN(n1071) );
NOR3_X1 U787 ( .A1(n1087), .A2(KEYINPUT42), .A3(n1088), .ZN(n1081) );
NOR2_X1 U788 ( .A1(n1089), .A2(n1072), .ZN(n1080) );
NOR2_X1 U789 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XNOR2_X1 U790 ( .A(n1092), .B(KEYINPUT0), .ZN(n1091) );
AND2_X1 U791 ( .A1(n1093), .A2(KEYINPUT42), .ZN(n1090) );
XNOR2_X1 U792 ( .A(KEYINPUT53), .B(n1094), .ZN(n1058) );
NAND3_X1 U793 ( .A1(n1095), .A2(n1096), .A3(n1097), .ZN(n1057) );
NAND4_X1 U794 ( .A1(n1079), .A2(n1087), .A3(n1086), .A4(n1098), .ZN(n1097) );
NAND2_X1 U795 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NAND2_X1 U796 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U797 ( .A1(n1073), .A2(n1103), .ZN(n1079) );
NOR3_X1 U798 ( .A1(n1104), .A2(G953), .A3(G952), .ZN(n1055) );
INV_X1 U799 ( .A(n1095), .ZN(n1104) );
NAND4_X1 U800 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1095) );
NOR4_X1 U801 ( .A1(n1109), .A2(n1110), .A3(n1062), .A4(n1111), .ZN(n1108) );
XNOR2_X1 U802 ( .A(KEYINPUT36), .B(n1112), .ZN(n1111) );
XNOR2_X1 U803 ( .A(n1113), .B(KEYINPUT39), .ZN(n1109) );
NOR3_X1 U804 ( .A1(n1114), .A2(n1115), .A3(n1116), .ZN(n1107) );
NOR2_X1 U805 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
INV_X1 U806 ( .A(G475), .ZN(n1118) );
NOR2_X1 U807 ( .A1(G902), .A2(n1119), .ZN(n1117) );
NAND2_X1 U808 ( .A1(G478), .A2(n1120), .ZN(n1106) );
NAND3_X1 U809 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
NAND2_X1 U810 ( .A1(n1124), .A2(n1122), .ZN(n1105) );
INV_X1 U811 ( .A(KEYINPUT27), .ZN(n1122) );
XOR2_X1 U812 ( .A(n1125), .B(n1126), .Z(G72) );
NOR2_X1 U813 ( .A1(n1127), .A2(n1096), .ZN(n1126) );
NOR2_X1 U814 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U815 ( .A1(n1130), .A2(n1131), .ZN(n1125) );
NAND2_X1 U816 ( .A1(n1132), .A2(n1096), .ZN(n1131) );
XNOR2_X1 U817 ( .A(n1133), .B(n1134), .ZN(n1132) );
NAND3_X1 U818 ( .A1(n1134), .A2(G900), .A3(G953), .ZN(n1130) );
AND2_X1 U819 ( .A1(n1135), .A2(KEYINPUT46), .ZN(n1134) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
XNOR2_X1 U821 ( .A(n1138), .B(n1139), .ZN(n1137) );
NOR2_X1 U822 ( .A1(KEYINPUT45), .A2(n1140), .ZN(n1139) );
XOR2_X1 U823 ( .A(KEYINPUT22), .B(n1141), .Z(n1140) );
NAND2_X1 U824 ( .A1(n1142), .A2(KEYINPUT34), .ZN(n1138) );
XNOR2_X1 U825 ( .A(n1143), .B(KEYINPUT13), .ZN(n1142) );
XOR2_X1 U826 ( .A(n1144), .B(n1145), .Z(G69) );
XOR2_X1 U827 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND3_X1 U828 ( .A1(n1094), .A2(n1096), .A3(KEYINPUT6), .ZN(n1147) );
NAND2_X1 U829 ( .A1(n1148), .A2(n1149), .ZN(n1146) );
NAND2_X1 U830 ( .A1(G953), .A2(n1150), .ZN(n1149) );
XNOR2_X1 U831 ( .A(n1151), .B(n1152), .ZN(n1148) );
NAND2_X1 U832 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
INV_X1 U833 ( .A(n1155), .ZN(n1154) );
NAND2_X1 U834 ( .A1(n1156), .A2(n1157), .ZN(n1153) );
XNOR2_X1 U835 ( .A(n1158), .B(KEYINPUT24), .ZN(n1156) );
NOR2_X1 U836 ( .A1(n1159), .A2(n1096), .ZN(n1144) );
NOR2_X1 U837 ( .A1(n1160), .A2(n1150), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1161), .A2(n1162), .ZN(G66) );
XOR2_X1 U839 ( .A(n1163), .B(n1164), .Z(n1162) );
NAND2_X1 U840 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
NOR2_X1 U841 ( .A1(n1161), .A2(n1167), .ZN(G63) );
XNOR2_X1 U842 ( .A(n1168), .B(n1169), .ZN(n1167) );
NAND4_X1 U843 ( .A1(KEYINPUT8), .A2(G478), .A3(n1170), .A4(n1171), .ZN(n1168) );
XNOR2_X1 U844 ( .A(KEYINPUT23), .B(n1121), .ZN(n1170) );
NOR2_X1 U845 ( .A1(n1161), .A2(n1172), .ZN(G60) );
XNOR2_X1 U846 ( .A(n1173), .B(n1119), .ZN(n1172) );
NAND2_X1 U847 ( .A1(n1165), .A2(G475), .ZN(n1173) );
XNOR2_X1 U848 ( .A(G104), .B(n1174), .ZN(G6) );
NAND4_X1 U849 ( .A1(n1175), .A2(n1051), .A3(n1086), .A4(n1176), .ZN(n1174) );
NOR2_X1 U850 ( .A1(n1161), .A2(n1177), .ZN(G57) );
XOR2_X1 U851 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U852 ( .A(n1180), .B(n1181), .ZN(n1179) );
XOR2_X1 U853 ( .A(n1182), .B(n1183), .Z(n1180) );
NOR2_X1 U854 ( .A1(KEYINPUT56), .A2(n1184), .ZN(n1183) );
NAND2_X1 U855 ( .A1(n1165), .A2(G472), .ZN(n1182) );
XOR2_X1 U856 ( .A(n1185), .B(n1186), .Z(n1178) );
NOR2_X1 U857 ( .A1(KEYINPUT40), .A2(n1187), .ZN(n1186) );
XNOR2_X1 U858 ( .A(n1188), .B(G101), .ZN(n1185) );
NOR2_X1 U859 ( .A1(n1161), .A2(n1189), .ZN(G54) );
XOR2_X1 U860 ( .A(n1190), .B(n1191), .Z(n1189) );
XNOR2_X1 U861 ( .A(n1192), .B(n1193), .ZN(n1191) );
XOR2_X1 U862 ( .A(n1194), .B(n1195), .Z(n1190) );
NAND2_X1 U863 ( .A1(n1165), .A2(G469), .ZN(n1194) );
NOR2_X1 U864 ( .A1(n1196), .A2(n1197), .ZN(G51) );
XOR2_X1 U865 ( .A(KEYINPUT21), .B(n1161), .Z(n1197) );
NOR2_X1 U866 ( .A1(n1096), .A2(G952), .ZN(n1161) );
XOR2_X1 U867 ( .A(n1198), .B(n1199), .Z(n1196) );
XNOR2_X1 U868 ( .A(KEYINPUT58), .B(n1200), .ZN(n1199) );
XOR2_X1 U869 ( .A(n1201), .B(n1202), .Z(n1198) );
NOR2_X1 U870 ( .A1(n1203), .A2(n1204), .ZN(n1202) );
AND2_X1 U871 ( .A1(KEYINPUT43), .A2(n1205), .ZN(n1204) );
NOR2_X1 U872 ( .A1(KEYINPUT44), .A2(n1205), .ZN(n1203) );
XOR2_X1 U873 ( .A(n1206), .B(n1207), .Z(n1205) );
NAND2_X1 U874 ( .A1(KEYINPUT37), .A2(n1208), .ZN(n1206) );
INV_X1 U875 ( .A(n1187), .ZN(n1208) );
NAND2_X1 U876 ( .A1(n1165), .A2(n1209), .ZN(n1201) );
AND2_X1 U877 ( .A1(G902), .A2(n1171), .ZN(n1165) );
NAND2_X1 U878 ( .A1(n1133), .A2(n1210), .ZN(n1171) );
INV_X1 U879 ( .A(n1094), .ZN(n1210) );
NAND4_X1 U880 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1094) );
NOR4_X1 U881 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1214) );
NAND3_X1 U882 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1213) );
OR2_X1 U883 ( .A1(n1222), .A2(KEYINPUT57), .ZN(n1220) );
NAND2_X1 U884 ( .A1(KEYINPUT57), .A2(n1223), .ZN(n1219) );
NAND3_X1 U885 ( .A1(n1176), .A2(n1099), .A3(n1224), .ZN(n1223) );
NAND4_X1 U886 ( .A1(n1051), .A2(n1086), .A3(n1225), .A4(n1226), .ZN(n1211) );
NAND2_X1 U887 ( .A1(n1054), .A2(n1227), .ZN(n1226) );
NAND2_X1 U888 ( .A1(KEYINPUT59), .A2(n1175), .ZN(n1227) );
NAND3_X1 U889 ( .A1(n1228), .A2(n1085), .A3(n1176), .ZN(n1225) );
OR2_X1 U890 ( .A1(n1084), .A2(KEYINPUT59), .ZN(n1228) );
INV_X1 U891 ( .A(n1060), .ZN(n1133) );
NAND4_X1 U892 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1060) );
NOR4_X1 U893 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1232) );
NAND2_X1 U894 ( .A1(n1092), .A2(n1237), .ZN(n1231) );
NAND2_X1 U895 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NAND2_X1 U896 ( .A1(n1240), .A2(n1175), .ZN(n1238) );
NAND2_X1 U897 ( .A1(n1241), .A2(n1242), .ZN(n1229) );
XNOR2_X1 U898 ( .A(KEYINPUT26), .B(n1243), .ZN(n1242) );
XNOR2_X1 U899 ( .A(G146), .B(n1230), .ZN(G48) );
NAND2_X1 U900 ( .A1(n1244), .A2(n1175), .ZN(n1230) );
XOR2_X1 U901 ( .A(n1245), .B(n1246), .Z(G45) );
NOR2_X1 U902 ( .A1(G143), .A2(KEYINPUT60), .ZN(n1246) );
NAND2_X1 U903 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
XNOR2_X1 U904 ( .A(KEYINPUT9), .B(n1249), .ZN(n1248) );
INV_X1 U905 ( .A(n1239), .ZN(n1247) );
NAND4_X1 U906 ( .A1(n1250), .A2(n1051), .A3(n1251), .A4(n1252), .ZN(n1239) );
XOR2_X1 U907 ( .A(G140), .B(n1236), .Z(G42) );
AND2_X1 U908 ( .A1(n1240), .A2(n1253), .ZN(n1236) );
XNOR2_X1 U909 ( .A(G137), .B(n1254), .ZN(G39) );
NAND2_X1 U910 ( .A1(KEYINPUT11), .A2(n1235), .ZN(n1254) );
AND2_X1 U911 ( .A1(n1240), .A2(n1221), .ZN(n1235) );
XOR2_X1 U912 ( .A(G134), .B(n1255), .Z(G36) );
NOR2_X1 U913 ( .A1(n1062), .A2(n1243), .ZN(n1255) );
NAND4_X1 U914 ( .A1(n1092), .A2(n1256), .A3(n1075), .A4(n1251), .ZN(n1243) );
XNOR2_X1 U915 ( .A(G131), .B(n1257), .ZN(G33) );
NAND3_X1 U916 ( .A1(n1092), .A2(n1240), .A3(n1258), .ZN(n1257) );
XNOR2_X1 U917 ( .A(n1175), .B(KEYINPUT10), .ZN(n1258) );
INV_X1 U918 ( .A(n1084), .ZN(n1175) );
AND3_X1 U919 ( .A1(n1075), .A2(n1251), .A3(n1241), .ZN(n1240) );
INV_X1 U920 ( .A(n1062), .ZN(n1241) );
NAND2_X1 U921 ( .A1(n1102), .A2(n1259), .ZN(n1062) );
XOR2_X1 U922 ( .A(G128), .B(n1234), .Z(G30) );
AND2_X1 U923 ( .A1(n1244), .A2(n1256), .ZN(n1234) );
INV_X1 U924 ( .A(n1085), .ZN(n1256) );
AND4_X1 U925 ( .A1(n1051), .A2(n1260), .A3(n1113), .A4(n1251), .ZN(n1244) );
XNOR2_X1 U926 ( .A(n1261), .B(n1216), .ZN(G3) );
AND2_X1 U927 ( .A1(n1262), .A2(n1092), .ZN(n1216) );
XNOR2_X1 U928 ( .A(n1233), .B(n1263), .ZN(G27) );
XNOR2_X1 U929 ( .A(G125), .B(KEYINPUT49), .ZN(n1263) );
AND4_X1 U930 ( .A1(n1224), .A2(n1253), .A3(n1264), .A4(n1251), .ZN(n1233) );
NAND2_X1 U931 ( .A1(n1073), .A2(n1265), .ZN(n1251) );
NAND4_X1 U932 ( .A1(G953), .A2(G902), .A3(n1266), .A4(n1129), .ZN(n1265) );
INV_X1 U933 ( .A(G900), .ZN(n1129) );
NOR2_X1 U934 ( .A1(n1088), .A2(n1084), .ZN(n1253) );
INV_X1 U935 ( .A(n1093), .ZN(n1088) );
INV_X1 U936 ( .A(n1103), .ZN(n1224) );
XNOR2_X1 U937 ( .A(G122), .B(n1212), .ZN(G24) );
NAND4_X1 U938 ( .A1(n1250), .A2(n1222), .A3(n1086), .A4(n1252), .ZN(n1212) );
NOR2_X1 U939 ( .A1(n1113), .A2(n1260), .ZN(n1086) );
XOR2_X1 U940 ( .A(n1267), .B(n1268), .Z(G21) );
XOR2_X1 U941 ( .A(KEYINPUT35), .B(G119), .Z(n1268) );
AND2_X1 U942 ( .A1(n1221), .A2(n1222), .ZN(n1267) );
NOR3_X1 U943 ( .A1(n1269), .A2(n1270), .A3(n1072), .ZN(n1221) );
XNOR2_X1 U944 ( .A(n1271), .B(n1218), .ZN(G18) );
NOR3_X1 U945 ( .A1(n1249), .A2(n1085), .A3(n1272), .ZN(n1218) );
NAND2_X1 U946 ( .A1(n1273), .A2(n1252), .ZN(n1085) );
INV_X1 U947 ( .A(n1274), .ZN(n1252) );
XNOR2_X1 U948 ( .A(n1275), .B(n1217), .ZN(G15) );
NOR3_X1 U949 ( .A1(n1249), .A2(n1084), .A3(n1272), .ZN(n1217) );
INV_X1 U950 ( .A(n1222), .ZN(n1272) );
NOR3_X1 U951 ( .A1(n1099), .A2(n1054), .A3(n1103), .ZN(n1222) );
NAND2_X1 U952 ( .A1(n1112), .A2(n1276), .ZN(n1103) );
INV_X1 U953 ( .A(n1077), .ZN(n1112) );
INV_X1 U954 ( .A(n1176), .ZN(n1054) );
INV_X1 U955 ( .A(n1264), .ZN(n1099) );
NAND2_X1 U956 ( .A1(n1274), .A2(n1250), .ZN(n1084) );
XNOR2_X1 U957 ( .A(n1273), .B(KEYINPUT52), .ZN(n1250) );
INV_X1 U958 ( .A(n1092), .ZN(n1249) );
NOR2_X1 U959 ( .A1(n1260), .A2(n1270), .ZN(n1092) );
INV_X1 U960 ( .A(n1113), .ZN(n1270) );
XOR2_X1 U961 ( .A(G110), .B(n1215), .Z(G12) );
AND2_X1 U962 ( .A1(n1262), .A2(n1093), .ZN(n1215) );
NOR2_X1 U963 ( .A1(n1113), .A2(n1269), .ZN(n1093) );
INV_X1 U964 ( .A(n1260), .ZN(n1269) );
XOR2_X1 U965 ( .A(n1110), .B(KEYINPUT47), .Z(n1260) );
XNOR2_X1 U966 ( .A(n1277), .B(n1166), .ZN(n1110) );
AND2_X1 U967 ( .A1(G217), .A2(n1278), .ZN(n1166) );
NAND2_X1 U968 ( .A1(n1121), .A2(n1163), .ZN(n1277) );
NAND2_X1 U969 ( .A1(n1279), .A2(n1280), .ZN(n1163) );
NAND2_X1 U970 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U971 ( .A(n1283), .B(KEYINPUT54), .Z(n1279) );
OR2_X1 U972 ( .A1(n1282), .A2(n1281), .ZN(n1283) );
XOR2_X1 U973 ( .A(n1284), .B(G137), .Z(n1281) );
NAND3_X1 U974 ( .A1(G234), .A2(n1096), .A3(G221), .ZN(n1284) );
XNOR2_X1 U975 ( .A(n1285), .B(n1286), .ZN(n1282) );
XNOR2_X1 U976 ( .A(G110), .B(n1287), .ZN(n1286) );
NAND2_X1 U977 ( .A1(KEYINPUT14), .A2(n1288), .ZN(n1287) );
XOR2_X1 U978 ( .A(G146), .B(n1141), .Z(n1288) );
XNOR2_X1 U979 ( .A(G119), .B(G128), .ZN(n1285) );
XNOR2_X1 U980 ( .A(n1289), .B(G472), .ZN(n1113) );
NAND2_X1 U981 ( .A1(n1290), .A2(n1121), .ZN(n1289) );
XOR2_X1 U982 ( .A(n1291), .B(n1292), .Z(n1290) );
XNOR2_X1 U983 ( .A(KEYINPUT48), .B(n1261), .ZN(n1292) );
XNOR2_X1 U984 ( .A(n1293), .B(n1184), .ZN(n1291) );
NAND2_X1 U985 ( .A1(n1294), .A2(n1295), .ZN(n1184) );
XOR2_X1 U986 ( .A(KEYINPUT15), .B(G210), .Z(n1295) );
NAND2_X1 U987 ( .A1(n1296), .A2(KEYINPUT61), .ZN(n1293) );
XNOR2_X1 U988 ( .A(n1187), .B(n1297), .ZN(n1296) );
XNOR2_X1 U989 ( .A(n1298), .B(n1299), .ZN(n1297) );
NOR2_X1 U990 ( .A1(n1188), .A2(KEYINPUT19), .ZN(n1299) );
AND2_X1 U991 ( .A1(n1300), .A2(n1301), .ZN(n1188) );
XOR2_X1 U992 ( .A(n1302), .B(KEYINPUT25), .Z(n1300) );
NAND2_X1 U993 ( .A1(n1303), .A2(n1275), .ZN(n1302) );
INV_X1 U994 ( .A(G113), .ZN(n1275) );
XOR2_X1 U995 ( .A(KEYINPUT16), .B(n1304), .Z(n1303) );
NAND2_X1 U996 ( .A1(KEYINPUT30), .A2(n1181), .ZN(n1298) );
AND3_X1 U997 ( .A1(n1051), .A2(n1176), .A3(n1087), .ZN(n1262) );
INV_X1 U998 ( .A(n1072), .ZN(n1087) );
NAND2_X1 U999 ( .A1(n1274), .A2(n1273), .ZN(n1072) );
NOR2_X1 U1000 ( .A1(n1305), .A2(n1115), .ZN(n1273) );
NOR3_X1 U1001 ( .A1(G475), .A2(G902), .A3(n1119), .ZN(n1115) );
AND2_X1 U1002 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U1003 ( .A1(n1308), .A2(n1121), .ZN(n1307) );
INV_X1 U1004 ( .A(n1119), .ZN(n1308) );
XNOR2_X1 U1005 ( .A(n1309), .B(n1310), .ZN(n1119) );
XNOR2_X1 U1006 ( .A(n1311), .B(n1312), .ZN(n1310) );
NAND2_X1 U1007 ( .A1(KEYINPUT29), .A2(n1141), .ZN(n1311) );
XOR2_X1 U1008 ( .A(G140), .B(G125), .Z(n1141) );
XOR2_X1 U1009 ( .A(n1313), .B(n1314), .Z(n1309) );
NOR2_X1 U1010 ( .A1(n1315), .A2(n1316), .ZN(n1314) );
XOR2_X1 U1011 ( .A(KEYINPUT28), .B(n1317), .Z(n1316) );
NOR2_X1 U1012 ( .A1(G104), .A2(n1318), .ZN(n1317) );
AND2_X1 U1013 ( .A1(n1318), .A2(G104), .ZN(n1315) );
XNOR2_X1 U1014 ( .A(G113), .B(n1319), .ZN(n1318) );
XOR2_X1 U1015 ( .A(n1320), .B(n1321), .Z(n1313) );
NOR2_X1 U1016 ( .A1(G131), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1017 ( .A(KEYINPUT51), .B(KEYINPUT38), .Z(n1322) );
NAND2_X1 U1018 ( .A1(n1294), .A2(G214), .ZN(n1320) );
NOR2_X1 U1019 ( .A1(G953), .A2(G237), .ZN(n1294) );
XNOR2_X1 U1020 ( .A(G475), .B(KEYINPUT31), .ZN(n1306) );
NOR2_X1 U1021 ( .A1(n1323), .A2(n1124), .ZN(n1274) );
NOR3_X1 U1022 ( .A1(G478), .A2(G902), .A3(n1169), .ZN(n1124) );
INV_X1 U1023 ( .A(n1123), .ZN(n1169) );
AND2_X1 U1024 ( .A1(G478), .A2(n1324), .ZN(n1323) );
NAND2_X1 U1025 ( .A1(n1123), .A2(n1121), .ZN(n1324) );
XOR2_X1 U1026 ( .A(n1325), .B(n1326), .Z(n1123) );
XOR2_X1 U1027 ( .A(n1327), .B(n1328), .Z(n1326) );
NOR2_X1 U1028 ( .A1(G143), .A2(KEYINPUT41), .ZN(n1328) );
AND3_X1 U1029 ( .A1(G217), .A2(n1096), .A3(G234), .ZN(n1327) );
XOR2_X1 U1030 ( .A(n1329), .B(n1330), .Z(n1325) );
NOR2_X1 U1031 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1032 ( .A(KEYINPUT63), .B(n1333), .Z(n1332) );
NOR2_X1 U1033 ( .A1(G107), .A2(n1334), .ZN(n1333) );
AND2_X1 U1034 ( .A1(n1334), .A2(G107), .ZN(n1331) );
NAND2_X1 U1035 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
NAND2_X1 U1036 ( .A1(G116), .A2(n1319), .ZN(n1336) );
INV_X1 U1037 ( .A(G122), .ZN(n1319) );
XOR2_X1 U1038 ( .A(n1337), .B(KEYINPUT3), .Z(n1335) );
NAND2_X1 U1039 ( .A1(G122), .A2(n1271), .ZN(n1337) );
XNOR2_X1 U1040 ( .A(G134), .B(G128), .ZN(n1329) );
NAND2_X1 U1041 ( .A1(n1073), .A2(n1338), .ZN(n1176) );
NAND4_X1 U1042 ( .A1(G953), .A2(G902), .A3(n1266), .A4(n1150), .ZN(n1338) );
INV_X1 U1043 ( .A(G898), .ZN(n1150) );
NAND3_X1 U1044 ( .A1(n1266), .A2(n1096), .A3(G952), .ZN(n1073) );
INV_X1 U1045 ( .A(G953), .ZN(n1096) );
NAND2_X1 U1046 ( .A1(G237), .A2(n1339), .ZN(n1266) );
AND2_X1 U1047 ( .A1(n1264), .A2(n1075), .ZN(n1051) );
AND2_X1 U1048 ( .A1(n1276), .A2(n1077), .ZN(n1075) );
XNOR2_X1 U1049 ( .A(n1340), .B(n1341), .ZN(n1077) );
XOR2_X1 U1050 ( .A(KEYINPUT50), .B(G469), .Z(n1341) );
NAND2_X1 U1051 ( .A1(n1342), .A2(n1121), .ZN(n1340) );
XOR2_X1 U1052 ( .A(n1343), .B(n1195), .Z(n1342) );
XNOR2_X1 U1053 ( .A(n1344), .B(n1345), .ZN(n1195) );
XOR2_X1 U1054 ( .A(G140), .B(G110), .Z(n1345) );
XOR2_X1 U1055 ( .A(n1181), .B(n1346), .Z(n1344) );
NOR2_X1 U1056 ( .A1(G953), .A2(n1128), .ZN(n1346) );
INV_X1 U1057 ( .A(G227), .ZN(n1128) );
XOR2_X1 U1058 ( .A(n1136), .B(KEYINPUT20), .Z(n1181) );
XNOR2_X1 U1059 ( .A(G131), .B(n1347), .ZN(n1136) );
XOR2_X1 U1060 ( .A(G137), .B(G134), .Z(n1347) );
NAND4_X1 U1061 ( .A1(KEYINPUT32), .A2(n1348), .A3(n1349), .A4(n1350), .ZN(n1343) );
NAND3_X1 U1062 ( .A1(KEYINPUT62), .A2(n1351), .A3(n1193), .ZN(n1350) );
OR2_X1 U1063 ( .A1(n1193), .A2(n1351), .ZN(n1349) );
NOR2_X1 U1064 ( .A1(KEYINPUT5), .A2(n1143), .ZN(n1351) );
XNOR2_X1 U1065 ( .A(n1352), .B(n1353), .ZN(n1193) );
NAND2_X1 U1066 ( .A1(KEYINPUT4), .A2(n1261), .ZN(n1352) );
INV_X1 U1067 ( .A(G101), .ZN(n1261) );
OR2_X1 U1068 ( .A1(n1192), .A2(KEYINPUT62), .ZN(n1348) );
INV_X1 U1069 ( .A(n1143), .ZN(n1192) );
XNOR2_X1 U1070 ( .A(n1354), .B(n1355), .ZN(n1143) );
NOR2_X1 U1071 ( .A1(G146), .A2(KEYINPUT55), .ZN(n1355) );
XNOR2_X1 U1072 ( .A(G128), .B(G143), .ZN(n1354) );
XNOR2_X1 U1073 ( .A(n1116), .B(KEYINPUT1), .ZN(n1276) );
INV_X1 U1074 ( .A(n1076), .ZN(n1116) );
NAND2_X1 U1075 ( .A1(G221), .A2(n1278), .ZN(n1076) );
NAND2_X1 U1076 ( .A1(n1339), .A2(n1121), .ZN(n1278) );
XNOR2_X1 U1077 ( .A(G234), .B(KEYINPUT7), .ZN(n1339) );
NOR2_X1 U1078 ( .A1(n1102), .A2(n1101), .ZN(n1264) );
INV_X1 U1079 ( .A(n1259), .ZN(n1101) );
NAND2_X1 U1080 ( .A1(G214), .A2(n1356), .ZN(n1259) );
XOR2_X1 U1081 ( .A(n1357), .B(n1209), .Z(n1102) );
AND2_X1 U1082 ( .A1(G210), .A2(n1356), .ZN(n1209) );
NAND2_X1 U1083 ( .A1(n1358), .A2(n1121), .ZN(n1356) );
INV_X1 U1084 ( .A(G237), .ZN(n1358) );
NAND2_X1 U1085 ( .A1(n1359), .A2(n1121), .ZN(n1357) );
INV_X1 U1086 ( .A(G902), .ZN(n1121) );
XOR2_X1 U1087 ( .A(n1207), .B(n1360), .Z(n1359) );
XNOR2_X1 U1088 ( .A(n1200), .B(n1187), .ZN(n1360) );
XOR2_X1 U1089 ( .A(n1361), .B(n1362), .Z(n1187) );
INV_X1 U1090 ( .A(n1312), .ZN(n1362) );
XOR2_X1 U1091 ( .A(G143), .B(G146), .Z(n1312) );
XNOR2_X1 U1092 ( .A(G128), .B(KEYINPUT18), .ZN(n1361) );
NAND3_X1 U1093 ( .A1(n1363), .A2(n1364), .A3(n1365), .ZN(n1200) );
NAND2_X1 U1094 ( .A1(n1155), .A2(n1152), .ZN(n1365) );
NOR2_X1 U1095 ( .A1(n1158), .A2(n1157), .ZN(n1155) );
NAND3_X1 U1096 ( .A1(n1157), .A2(n1366), .A3(n1367), .ZN(n1364) );
INV_X1 U1097 ( .A(n1158), .ZN(n1367) );
INV_X1 U1098 ( .A(n1152), .ZN(n1366) );
NAND2_X1 U1099 ( .A1(n1158), .A2(n1368), .ZN(n1363) );
XNOR2_X1 U1100 ( .A(n1157), .B(n1152), .ZN(n1368) );
XOR2_X1 U1101 ( .A(G110), .B(n1369), .Z(n1152) );
NOR2_X1 U1102 ( .A1(G122), .A2(KEYINPUT12), .ZN(n1369) );
AND2_X1 U1103 ( .A1(n1370), .A2(n1371), .ZN(n1157) );
OR2_X1 U1104 ( .A1(n1304), .A2(G113), .ZN(n1371) );
XOR2_X1 U1105 ( .A(n1301), .B(KEYINPUT17), .Z(n1370) );
NAND2_X1 U1106 ( .A1(G113), .A2(n1304), .ZN(n1301) );
XNOR2_X1 U1107 ( .A(G119), .B(n1271), .ZN(n1304) );
INV_X1 U1108 ( .A(G116), .ZN(n1271) );
XOR2_X1 U1109 ( .A(G101), .B(n1353), .Z(n1158) );
XOR2_X1 U1110 ( .A(G104), .B(G107), .Z(n1353) );
XOR2_X1 U1111 ( .A(G125), .B(n1372), .Z(n1207) );
NOR2_X1 U1112 ( .A1(n1160), .A2(G953), .ZN(n1372) );
INV_X1 U1113 ( .A(G224), .ZN(n1160) );
endmodule


