//Key = 1000111110101101011001010111011000011001011101111000110000111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353;

XOR2_X1 U743 ( .A(G107), .B(n1025), .Z(G9) );
NOR3_X1 U744 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1025) );
XOR2_X1 U745 ( .A(KEYINPUT15), .B(n1029), .Z(n1026) );
NOR2_X1 U746 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U747 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
NOR2_X1 U748 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U749 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR2_X1 U750 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR2_X1 U751 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
NOR2_X1 U752 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR3_X1 U753 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1044) );
NOR2_X1 U754 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U755 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR2_X1 U756 ( .A1(n1053), .A2(n1054), .ZN(n1046) );
AND3_X1 U757 ( .A1(n1055), .A2(n1056), .A3(n1029), .ZN(n1042) );
NOR4_X1 U758 ( .A1(n1057), .A2(n1050), .A3(n1053), .A4(n1045), .ZN(n1038) );
NAND4_X1 U759 ( .A1(n1058), .A2(n1059), .A3(n1060), .A4(n1061), .ZN(n1032) );
NAND4_X1 U760 ( .A1(n1062), .A2(n1063), .A3(n1029), .A4(n1064), .ZN(n1059) );
NOR3_X1 U761 ( .A1(n1065), .A2(n1045), .A3(n1037), .ZN(n1064) );
XOR2_X1 U762 ( .A(KEYINPUT60), .B(n1066), .Z(n1065) );
XOR2_X1 U763 ( .A(KEYINPUT16), .B(n1055), .Z(n1062) );
NAND3_X1 U764 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1058) );
XOR2_X1 U765 ( .A(n1070), .B(KEYINPUT62), .Z(n1069) );
NAND4_X1 U766 ( .A1(n1071), .A2(n1072), .A3(n1055), .A4(n1029), .ZN(n1070) );
XOR2_X1 U767 ( .A(n1037), .B(KEYINPUT18), .Z(n1071) );
AND3_X1 U768 ( .A1(n1060), .A2(n1061), .A3(n1073), .ZN(n1030) );
NAND4_X1 U769 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1060) );
NOR4_X1 U770 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
XOR2_X1 U771 ( .A(KEYINPUT9), .B(n1082), .Z(n1081) );
XNOR2_X1 U772 ( .A(n1083), .B(n1084), .ZN(n1080) );
NOR3_X1 U773 ( .A1(n1085), .A2(n1068), .A3(n1066), .ZN(n1076) );
NOR2_X1 U774 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NOR2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR2_X1 U776 ( .A1(KEYINPUT59), .A2(n1090), .ZN(n1088) );
NAND3_X1 U777 ( .A1(n1091), .A2(n1092), .A3(KEYINPUT59), .ZN(n1075) );
NAND2_X1 U778 ( .A1(n1093), .A2(n1090), .ZN(n1092) );
INV_X1 U779 ( .A(KEYINPUT36), .ZN(n1090) );
NAND2_X1 U780 ( .A1(KEYINPUT36), .A2(n1094), .ZN(n1091) );
NAND2_X1 U781 ( .A1(n1086), .A2(n1093), .ZN(n1094) );
XOR2_X1 U782 ( .A(n1095), .B(n1096), .Z(G72) );
XOR2_X1 U783 ( .A(n1097), .B(n1098), .Z(n1096) );
NAND2_X1 U784 ( .A1(G953), .A2(n1099), .ZN(n1098) );
NAND2_X1 U785 ( .A1(G900), .A2(G227), .ZN(n1099) );
NAND4_X1 U786 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1097) );
NAND2_X1 U787 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
INV_X1 U788 ( .A(KEYINPUT58), .ZN(n1105) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1104) );
XNOR2_X1 U790 ( .A(KEYINPUT21), .B(n1108), .ZN(n1107) );
NAND2_X1 U791 ( .A1(KEYINPUT58), .A2(n1109), .ZN(n1102) );
NAND2_X1 U792 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND3_X1 U793 ( .A1(KEYINPUT21), .A2(n1106), .A3(n1108), .ZN(n1111) );
OR2_X1 U794 ( .A1(n1108), .A2(KEYINPUT21), .ZN(n1110) );
OR2_X1 U795 ( .A1(n1108), .A2(n1106), .ZN(n1101) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(n1106) );
XNOR2_X1 U797 ( .A(KEYINPUT53), .B(KEYINPUT13), .ZN(n1112) );
XNOR2_X1 U798 ( .A(n1114), .B(n1115), .ZN(n1108) );
NAND2_X1 U799 ( .A1(n1116), .A2(KEYINPUT63), .ZN(n1114) );
XOR2_X1 U800 ( .A(n1117), .B(n1118), .Z(n1116) );
XNOR2_X1 U801 ( .A(KEYINPUT6), .B(n1119), .ZN(n1117) );
NOR2_X1 U802 ( .A1(G134), .A2(KEYINPUT2), .ZN(n1119) );
XOR2_X1 U803 ( .A(KEYINPUT35), .B(n1120), .Z(n1100) );
NOR2_X1 U804 ( .A1(G900), .A2(n1061), .ZN(n1120) );
AND2_X1 U805 ( .A1(n1035), .A2(n1061), .ZN(n1095) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(G69) );
XOR2_X1 U807 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U808 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U809 ( .A(n1127), .B(n1128), .Z(n1126) );
XOR2_X1 U810 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U811 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
OR2_X1 U812 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
XOR2_X1 U813 ( .A(n1135), .B(KEYINPUT40), .Z(n1131) );
NAND2_X1 U814 ( .A1(n1134), .A2(n1133), .ZN(n1135) );
XNOR2_X1 U815 ( .A(n1136), .B(KEYINPUT14), .ZN(n1133) );
XOR2_X1 U816 ( .A(n1137), .B(G122), .Z(n1127) );
XNOR2_X1 U817 ( .A(KEYINPUT47), .B(KEYINPUT25), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1061), .A2(n1138), .ZN(n1125) );
XOR2_X1 U819 ( .A(KEYINPUT19), .B(G898), .Z(n1138) );
NAND3_X1 U820 ( .A1(n1033), .A2(n1061), .A3(KEYINPUT42), .ZN(n1123) );
NAND2_X1 U821 ( .A1(G953), .A2(n1139), .ZN(n1121) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1139) );
NOR2_X1 U823 ( .A1(n1140), .A2(n1141), .ZN(G66) );
NOR3_X1 U824 ( .A1(n1083), .A2(n1142), .A3(n1143), .ZN(n1141) );
NOR3_X1 U825 ( .A1(n1144), .A2(n1084), .A3(n1145), .ZN(n1143) );
INV_X1 U826 ( .A(n1146), .ZN(n1144) );
NOR2_X1 U827 ( .A1(n1147), .A2(n1146), .ZN(n1142) );
NOR2_X1 U828 ( .A1(n1148), .A2(n1084), .ZN(n1147) );
NOR2_X1 U829 ( .A1(n1035), .A2(n1033), .ZN(n1148) );
NOR2_X1 U830 ( .A1(n1140), .A2(n1149), .ZN(G63) );
XOR2_X1 U831 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U832 ( .A1(n1152), .A2(G478), .ZN(n1150) );
NOR2_X1 U833 ( .A1(n1140), .A2(n1153), .ZN(G60) );
XOR2_X1 U834 ( .A(n1154), .B(n1155), .Z(n1153) );
NAND2_X1 U835 ( .A1(n1152), .A2(G475), .ZN(n1154) );
XOR2_X1 U836 ( .A(G104), .B(n1156), .Z(G6) );
NOR2_X1 U837 ( .A1(n1140), .A2(n1157), .ZN(G57) );
XOR2_X1 U838 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U839 ( .A(n1160), .B(n1161), .Z(n1159) );
AND2_X1 U840 ( .A1(G472), .A2(n1152), .ZN(n1161) );
NOR2_X1 U841 ( .A1(KEYINPUT1), .A2(n1162), .ZN(n1160) );
XOR2_X1 U842 ( .A(n1163), .B(G101), .Z(n1162) );
NAND2_X1 U843 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U844 ( .A1(KEYINPUT51), .A2(n1166), .ZN(n1165) );
NAND2_X1 U845 ( .A1(KEYINPUT61), .A2(n1167), .ZN(n1164) );
INV_X1 U846 ( .A(n1166), .ZN(n1167) );
NOR3_X1 U847 ( .A1(n1168), .A2(n1169), .A3(n1170), .ZN(G54) );
NOR3_X1 U848 ( .A1(n1171), .A2(n1061), .A3(n1073), .ZN(n1170) );
INV_X1 U849 ( .A(G952), .ZN(n1073) );
AND2_X1 U850 ( .A1(n1171), .A2(n1140), .ZN(n1169) );
INV_X1 U851 ( .A(KEYINPUT32), .ZN(n1171) );
XOR2_X1 U852 ( .A(n1172), .B(n1173), .Z(n1168) );
XOR2_X1 U853 ( .A(n1174), .B(n1175), .Z(n1173) );
NAND2_X1 U854 ( .A1(n1152), .A2(G469), .ZN(n1174) );
INV_X1 U855 ( .A(n1145), .ZN(n1152) );
XOR2_X1 U856 ( .A(n1176), .B(n1177), .Z(n1172) );
NAND2_X1 U857 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
OR2_X1 U858 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U859 ( .A(n1182), .B(KEYINPUT20), .Z(n1178) );
NAND2_X1 U860 ( .A1(n1180), .A2(n1181), .ZN(n1182) );
XNOR2_X1 U861 ( .A(n1183), .B(G140), .ZN(n1180) );
NAND2_X1 U862 ( .A1(KEYINPUT8), .A2(n1130), .ZN(n1183) );
NOR2_X1 U863 ( .A1(n1140), .A2(n1184), .ZN(G51) );
XOR2_X1 U864 ( .A(n1185), .B(n1186), .Z(n1184) );
NOR2_X1 U865 ( .A1(n1093), .A2(n1145), .ZN(n1186) );
NAND2_X1 U866 ( .A1(G902), .A2(n1187), .ZN(n1145) );
OR2_X1 U867 ( .A1(n1033), .A2(n1035), .ZN(n1187) );
NAND4_X1 U868 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1035) );
NOR4_X1 U869 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
AND2_X1 U870 ( .A1(n1196), .A2(n1197), .ZN(n1190) );
NAND4_X1 U871 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1033) );
NOR4_X1 U872 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1156), .ZN(n1201) );
NOR3_X1 U873 ( .A1(n1028), .A2(n1050), .A3(n1205), .ZN(n1156) );
INV_X1 U874 ( .A(n1029), .ZN(n1050) );
INV_X1 U875 ( .A(n1206), .ZN(n1204) );
NAND2_X1 U876 ( .A1(n1207), .A2(n1208), .ZN(n1200) );
NAND2_X1 U877 ( .A1(n1209), .A2(n1205), .ZN(n1208) );
XOR2_X1 U878 ( .A(n1027), .B(KEYINPUT49), .Z(n1209) );
NAND4_X1 U879 ( .A1(n1210), .A2(n1055), .A3(n1211), .A4(n1212), .ZN(n1199) );
OR2_X1 U880 ( .A1(n1213), .A2(KEYINPUT54), .ZN(n1212) );
NAND2_X1 U881 ( .A1(KEYINPUT54), .A2(n1214), .ZN(n1211) );
NAND2_X1 U882 ( .A1(n1215), .A2(n1057), .ZN(n1214) );
INV_X1 U883 ( .A(n1216), .ZN(n1057) );
NAND3_X1 U884 ( .A1(n1051), .A2(n1029), .A3(n1213), .ZN(n1198) );
NOR2_X1 U885 ( .A1(KEYINPUT24), .A2(n1217), .ZN(n1185) );
XOR2_X1 U886 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U887 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U888 ( .A(n1222), .B(n1223), .Z(n1218) );
NOR2_X1 U889 ( .A1(n1061), .A2(G952), .ZN(n1140) );
XOR2_X1 U890 ( .A(n1188), .B(n1224), .Z(G48) );
NAND2_X1 U891 ( .A1(KEYINPUT29), .A2(G146), .ZN(n1224) );
NAND3_X1 U892 ( .A1(n1052), .A2(n1056), .A3(n1225), .ZN(n1188) );
XOR2_X1 U893 ( .A(n1226), .B(n1189), .Z(G45) );
NAND4_X1 U894 ( .A1(n1227), .A2(n1228), .A3(n1056), .A4(n1079), .ZN(n1189) );
XOR2_X1 U895 ( .A(n1229), .B(n1196), .Z(G42) );
NAND3_X1 U896 ( .A1(n1230), .A2(n1216), .A3(n1231), .ZN(n1196) );
XOR2_X1 U897 ( .A(G137), .B(n1195), .Z(G39) );
AND3_X1 U898 ( .A1(n1231), .A2(n1055), .A3(n1225), .ZN(n1195) );
XOR2_X1 U899 ( .A(n1232), .B(n1233), .Z(G36) );
NAND2_X1 U900 ( .A1(KEYINPUT52), .A2(n1194), .ZN(n1233) );
AND3_X1 U901 ( .A1(n1228), .A2(n1051), .A3(n1231), .ZN(n1194) );
XOR2_X1 U902 ( .A(G131), .B(n1193), .Z(G33) );
AND3_X1 U903 ( .A1(n1228), .A2(n1052), .A3(n1231), .ZN(n1193) );
INV_X1 U904 ( .A(n1045), .ZN(n1231) );
NAND2_X1 U905 ( .A1(n1067), .A2(n1234), .ZN(n1045) );
AND2_X1 U906 ( .A1(n1235), .A2(n1236), .ZN(n1228) );
NAND2_X1 U907 ( .A1(n1237), .A2(n1238), .ZN(G30) );
NAND2_X1 U908 ( .A1(G128), .A2(n1197), .ZN(n1238) );
XOR2_X1 U909 ( .A(n1239), .B(KEYINPUT33), .Z(n1237) );
OR2_X1 U910 ( .A1(n1197), .A2(G128), .ZN(n1239) );
NAND3_X1 U911 ( .A1(n1051), .A2(n1056), .A3(n1225), .ZN(n1197) );
AND2_X1 U912 ( .A1(n1235), .A2(n1240), .ZN(n1225) );
AND3_X1 U913 ( .A1(n1078), .A2(n1241), .A3(n1216), .ZN(n1235) );
XOR2_X1 U914 ( .A(G101), .B(n1202), .Z(G3) );
AND2_X1 U915 ( .A1(n1047), .A2(n1213), .ZN(n1202) );
INV_X1 U916 ( .A(n1028), .ZN(n1213) );
AND3_X1 U917 ( .A1(n1236), .A2(n1078), .A3(n1055), .ZN(n1047) );
XOR2_X1 U918 ( .A(G125), .B(n1192), .Z(G27) );
AND3_X1 U919 ( .A1(n1072), .A2(n1056), .A3(n1230), .ZN(n1192) );
AND3_X1 U920 ( .A1(n1052), .A2(n1241), .A3(n1210), .ZN(n1230) );
INV_X1 U921 ( .A(n1054), .ZN(n1210) );
NAND2_X1 U922 ( .A1(n1037), .A2(n1242), .ZN(n1241) );
NAND4_X1 U923 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1244), .ZN(n1242) );
INV_X1 U924 ( .A(G900), .ZN(n1244) );
XOR2_X1 U925 ( .A(n1245), .B(n1206), .Z(G24) );
NAND4_X1 U926 ( .A1(n1215), .A2(n1079), .A3(n1029), .A4(n1246), .ZN(n1206) );
AND2_X1 U927 ( .A1(n1072), .A2(n1227), .ZN(n1246) );
NOR2_X1 U928 ( .A1(n1240), .A2(n1078), .ZN(n1029) );
XOR2_X1 U929 ( .A(G119), .B(n1203), .Z(G21) );
AND3_X1 U930 ( .A1(n1055), .A2(n1240), .A3(n1247), .ZN(n1203) );
INV_X1 U931 ( .A(n1053), .ZN(n1055) );
XNOR2_X1 U932 ( .A(G116), .B(n1248), .ZN(G18) );
NAND2_X1 U933 ( .A1(n1207), .A2(n1051), .ZN(n1248) );
INV_X1 U934 ( .A(n1027), .ZN(n1051) );
NAND2_X1 U935 ( .A1(n1079), .A2(n1249), .ZN(n1027) );
INV_X1 U936 ( .A(n1250), .ZN(n1079) );
XNOR2_X1 U937 ( .A(G113), .B(n1251), .ZN(G15) );
NAND2_X1 U938 ( .A1(n1207), .A2(n1052), .ZN(n1251) );
INV_X1 U939 ( .A(n1205), .ZN(n1052) );
NAND2_X1 U940 ( .A1(n1227), .A2(n1250), .ZN(n1205) );
XOR2_X1 U941 ( .A(n1252), .B(KEYINPUT4), .Z(n1227) );
AND2_X1 U942 ( .A1(n1247), .A2(n1236), .ZN(n1207) );
INV_X1 U943 ( .A(n1240), .ZN(n1236) );
AND3_X1 U944 ( .A1(n1215), .A2(n1078), .A3(n1072), .ZN(n1247) );
INV_X1 U945 ( .A(n1041), .ZN(n1072) );
NAND2_X1 U946 ( .A1(n1063), .A2(n1253), .ZN(n1041) );
XOR2_X1 U947 ( .A(G110), .B(n1254), .Z(G12) );
NOR3_X1 U948 ( .A1(n1054), .A2(n1028), .A3(n1053), .ZN(n1254) );
NAND2_X1 U949 ( .A1(n1250), .A2(n1249), .ZN(n1053) );
XOR2_X1 U950 ( .A(n1082), .B(KEYINPUT41), .Z(n1249) );
INV_X1 U951 ( .A(n1252), .ZN(n1082) );
XOR2_X1 U952 ( .A(n1255), .B(G475), .Z(n1252) );
NAND2_X1 U953 ( .A1(n1155), .A2(n1256), .ZN(n1255) );
XOR2_X1 U954 ( .A(n1257), .B(n1258), .Z(n1155) );
XOR2_X1 U955 ( .A(n1259), .B(n1260), .Z(n1258) );
XOR2_X1 U956 ( .A(n1261), .B(n1221), .Z(n1260) );
XOR2_X1 U957 ( .A(G122), .B(G125), .Z(n1221) );
NAND2_X1 U958 ( .A1(KEYINPUT39), .A2(n1262), .ZN(n1261) );
XOR2_X1 U959 ( .A(KEYINPUT28), .B(G140), .Z(n1262) );
XOR2_X1 U960 ( .A(n1263), .B(n1264), .Z(n1259) );
AND3_X1 U961 ( .A1(G214), .A2(n1061), .A3(n1265), .ZN(n1264) );
NAND2_X1 U962 ( .A1(KEYINPUT48), .A2(n1226), .ZN(n1263) );
INV_X1 U963 ( .A(G143), .ZN(n1226) );
XOR2_X1 U964 ( .A(n1266), .B(n1267), .Z(n1257) );
XOR2_X1 U965 ( .A(G146), .B(G131), .Z(n1267) );
XNOR2_X1 U966 ( .A(G104), .B(G113), .ZN(n1266) );
XOR2_X1 U967 ( .A(n1268), .B(G478), .Z(n1250) );
NAND2_X1 U968 ( .A1(n1269), .A2(n1151), .ZN(n1268) );
XOR2_X1 U969 ( .A(n1270), .B(n1271), .Z(n1151) );
XOR2_X1 U970 ( .A(n1272), .B(n1273), .Z(n1271) );
NAND2_X1 U971 ( .A1(KEYINPUT0), .A2(n1245), .ZN(n1273) );
INV_X1 U972 ( .A(G122), .ZN(n1245) );
NAND3_X1 U973 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1272) );
NAND2_X1 U974 ( .A1(G134), .A2(n1277), .ZN(n1276) );
NAND2_X1 U975 ( .A1(KEYINPUT30), .A2(n1278), .ZN(n1277) );
XOR2_X1 U976 ( .A(KEYINPUT56), .B(n1279), .Z(n1278) );
NAND3_X1 U977 ( .A1(KEYINPUT30), .A2(n1232), .A3(n1279), .ZN(n1275) );
OR2_X1 U978 ( .A1(n1279), .A2(KEYINPUT30), .ZN(n1274) );
XOR2_X1 U979 ( .A(n1280), .B(KEYINPUT23), .Z(n1279) );
XOR2_X1 U980 ( .A(n1281), .B(n1282), .Z(n1270) );
AND3_X1 U981 ( .A1(G217), .A2(n1061), .A3(G234), .ZN(n1282) );
XNOR2_X1 U982 ( .A(G107), .B(G116), .ZN(n1281) );
XOR2_X1 U983 ( .A(n1256), .B(KEYINPUT11), .Z(n1269) );
NAND2_X1 U984 ( .A1(n1215), .A2(n1216), .ZN(n1028) );
NOR2_X1 U985 ( .A1(n1063), .A2(n1066), .ZN(n1216) );
INV_X1 U986 ( .A(n1253), .ZN(n1066) );
NAND2_X1 U987 ( .A1(G221), .A2(n1283), .ZN(n1253) );
XNOR2_X1 U988 ( .A(n1074), .B(KEYINPUT17), .ZN(n1063) );
XOR2_X1 U989 ( .A(n1284), .B(G469), .Z(n1074) );
NAND2_X1 U990 ( .A1(n1285), .A2(n1256), .ZN(n1284) );
XOR2_X1 U991 ( .A(n1286), .B(n1287), .Z(n1285) );
NOR2_X1 U992 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
XOR2_X1 U993 ( .A(KEYINPUT37), .B(n1290), .Z(n1289) );
AND2_X1 U994 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
NOR2_X1 U995 ( .A1(n1292), .A2(n1291), .ZN(n1288) );
XNOR2_X1 U996 ( .A(n1293), .B(n1294), .ZN(n1291) );
XOR2_X1 U997 ( .A(n1229), .B(KEYINPUT34), .Z(n1293) );
INV_X1 U998 ( .A(G140), .ZN(n1229) );
INV_X1 U999 ( .A(n1181), .ZN(n1292) );
NAND2_X1 U1000 ( .A1(G227), .A2(n1061), .ZN(n1181) );
NAND2_X1 U1001 ( .A1(n1295), .A2(n1296), .ZN(n1286) );
NAND2_X1 U1002 ( .A1(n1175), .A2(n1297), .ZN(n1296) );
NAND2_X1 U1003 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
XOR2_X1 U1004 ( .A(n1300), .B(n1301), .Z(n1298) );
NAND2_X1 U1005 ( .A1(n1302), .A2(n1303), .ZN(n1295) );
NAND2_X1 U1006 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U1007 ( .A1(n1306), .A2(n1300), .ZN(n1305) );
OR2_X1 U1008 ( .A1(n1176), .A2(n1300), .ZN(n1304) );
INV_X1 U1009 ( .A(KEYINPUT12), .ZN(n1300) );
NAND2_X1 U1010 ( .A1(n1299), .A2(n1301), .ZN(n1176) );
INV_X1 U1011 ( .A(n1306), .ZN(n1301) );
NOR2_X1 U1012 ( .A1(n1307), .A2(n1115), .ZN(n1306) );
NAND2_X1 U1013 ( .A1(n1115), .A2(n1307), .ZN(n1299) );
XOR2_X1 U1014 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1015 ( .A(n1310), .B(KEYINPUT5), .Z(n1308) );
INV_X1 U1016 ( .A(G101), .ZN(n1310) );
XNOR2_X1 U1017 ( .A(G146), .B(n1280), .ZN(n1115) );
XOR2_X1 U1018 ( .A(G128), .B(G143), .Z(n1280) );
INV_X1 U1019 ( .A(n1175), .ZN(n1302) );
AND2_X1 U1020 ( .A1(n1056), .A2(n1311), .ZN(n1215) );
NAND2_X1 U1021 ( .A1(n1037), .A2(n1312), .ZN(n1311) );
NAND4_X1 U1022 ( .A1(G953), .A2(G902), .A3(n1243), .A4(n1313), .ZN(n1312) );
INV_X1 U1023 ( .A(G898), .ZN(n1313) );
NAND3_X1 U1024 ( .A1(n1243), .A2(n1061), .A3(G952), .ZN(n1037) );
NAND2_X1 U1025 ( .A1(G237), .A2(G234), .ZN(n1243) );
NOR2_X1 U1026 ( .A1(n1067), .A2(n1068), .ZN(n1056) );
INV_X1 U1027 ( .A(n1234), .ZN(n1068) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1314), .ZN(n1234) );
XNOR2_X1 U1029 ( .A(n1086), .B(n1089), .ZN(n1067) );
INV_X1 U1030 ( .A(n1093), .ZN(n1089) );
NAND2_X1 U1031 ( .A1(G210), .A2(n1314), .ZN(n1093) );
NAND2_X1 U1032 ( .A1(n1256), .A2(n1265), .ZN(n1314) );
AND2_X1 U1033 ( .A1(n1315), .A2(n1256), .ZN(n1086) );
XOR2_X1 U1034 ( .A(n1316), .B(n1317), .Z(n1315) );
XNOR2_X1 U1035 ( .A(n1222), .B(n1318), .ZN(n1317) );
XOR2_X1 U1036 ( .A(G122), .B(n1319), .Z(n1318) );
NOR2_X1 U1037 ( .A1(KEYINPUT55), .A2(n1320), .ZN(n1319) );
XOR2_X1 U1038 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1039 ( .A(KEYINPUT3), .B(G125), .Z(n1322) );
NAND2_X1 U1040 ( .A1(G224), .A2(n1061), .ZN(n1222) );
XNOR2_X1 U1041 ( .A(n1220), .B(n1134), .ZN(n1316) );
XOR2_X1 U1042 ( .A(n1136), .B(n1294), .Z(n1220) );
XOR2_X1 U1043 ( .A(n1323), .B(KEYINPUT43), .Z(n1136) );
NAND2_X1 U1044 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
NAND2_X1 U1045 ( .A1(n1309), .A2(n1326), .ZN(n1325) );
XOR2_X1 U1046 ( .A(KEYINPUT7), .B(n1327), .Z(n1324) );
NOR2_X1 U1047 ( .A1(n1309), .A2(n1326), .ZN(n1327) );
XOR2_X1 U1048 ( .A(KEYINPUT27), .B(G101), .Z(n1326) );
XNOR2_X1 U1049 ( .A(G104), .B(G107), .ZN(n1309) );
NAND2_X1 U1050 ( .A1(n1328), .A2(n1240), .ZN(n1054) );
NAND2_X1 U1051 ( .A1(n1329), .A2(n1330), .ZN(n1240) );
NAND2_X1 U1052 ( .A1(n1083), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1053 ( .A(n1332), .B(KEYINPUT38), .Z(n1329) );
OR2_X1 U1054 ( .A1(n1331), .A2(n1083), .ZN(n1332) );
NOR2_X1 U1055 ( .A1(n1146), .A2(G902), .ZN(n1083) );
XOR2_X1 U1056 ( .A(n1333), .B(n1334), .Z(n1146) );
XOR2_X1 U1057 ( .A(n1335), .B(n1113), .Z(n1334) );
XOR2_X1 U1058 ( .A(G125), .B(G140), .Z(n1113) );
AND3_X1 U1059 ( .A1(n1336), .A2(G234), .A3(G221), .ZN(n1335) );
XOR2_X1 U1060 ( .A(KEYINPUT31), .B(n1061), .Z(n1336) );
XOR2_X1 U1061 ( .A(n1337), .B(n1338), .Z(n1333) );
NOR2_X1 U1062 ( .A1(KEYINPUT57), .A2(n1339), .ZN(n1338) );
XOR2_X1 U1063 ( .A(n1294), .B(n1340), .Z(n1339) );
XOR2_X1 U1064 ( .A(G128), .B(G119), .Z(n1340) );
INV_X1 U1065 ( .A(n1130), .ZN(n1294) );
XNOR2_X1 U1066 ( .A(G110), .B(KEYINPUT45), .ZN(n1130) );
XNOR2_X1 U1067 ( .A(G137), .B(G146), .ZN(n1337) );
XNOR2_X1 U1068 ( .A(n1084), .B(KEYINPUT26), .ZN(n1331) );
NAND2_X1 U1069 ( .A1(G217), .A2(n1283), .ZN(n1084) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1256), .ZN(n1283) );
XOR2_X1 U1071 ( .A(KEYINPUT10), .B(n1078), .Z(n1328) );
XNOR2_X1 U1072 ( .A(n1341), .B(n1342), .ZN(n1078) );
XOR2_X1 U1073 ( .A(KEYINPUT44), .B(G472), .Z(n1342) );
NAND2_X1 U1074 ( .A1(n1343), .A2(n1256), .ZN(n1341) );
INV_X1 U1075 ( .A(G902), .ZN(n1256) );
XOR2_X1 U1076 ( .A(n1344), .B(n1345), .Z(n1343) );
NOR2_X1 U1077 ( .A1(KEYINPUT50), .A2(n1346), .ZN(n1345) );
XOR2_X1 U1078 ( .A(n1166), .B(G101), .Z(n1346) );
NAND3_X1 U1079 ( .A1(n1265), .A2(n1061), .A3(G210), .ZN(n1166) );
INV_X1 U1080 ( .A(G953), .ZN(n1061) );
INV_X1 U1081 ( .A(G237), .ZN(n1265) );
NAND2_X1 U1082 ( .A1(n1347), .A2(n1348), .ZN(n1344) );
NAND2_X1 U1083 ( .A1(n1158), .A2(n1349), .ZN(n1348) );
INV_X1 U1084 ( .A(KEYINPUT22), .ZN(n1349) );
XNOR2_X1 U1085 ( .A(n1223), .B(n1175), .ZN(n1158) );
XNOR2_X1 U1086 ( .A(n1134), .B(n1321), .ZN(n1223) );
NAND3_X1 U1087 ( .A1(n1350), .A2(n1134), .A3(KEYINPUT22), .ZN(n1347) );
XNOR2_X1 U1088 ( .A(G113), .B(n1351), .ZN(n1134) );
XOR2_X1 U1089 ( .A(G119), .B(G116), .Z(n1351) );
XOR2_X1 U1090 ( .A(n1175), .B(n1321), .Z(n1350) );
XNOR2_X1 U1091 ( .A(n1352), .B(G128), .ZN(n1321) );
NAND2_X1 U1092 ( .A1(KEYINPUT46), .A2(n1353), .ZN(n1352) );
XOR2_X1 U1093 ( .A(G146), .B(G143), .Z(n1353) );
XOR2_X1 U1094 ( .A(n1232), .B(n1118), .Z(n1175) );
XOR2_X1 U1095 ( .A(G131), .B(G137), .Z(n1118) );
INV_X1 U1096 ( .A(G134), .ZN(n1232) );
endmodule


