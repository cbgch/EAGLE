//Key = 0001111100100100110110101010111010000101110100011111011100101100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;

XNOR2_X1 U713 ( .A(G107), .B(n984), .ZN(G9) );
NOR2_X1 U714 ( .A1(n985), .A2(n986), .ZN(G75) );
NOR4_X1 U715 ( .A1(n987), .A2(n988), .A3(n989), .A4(n990), .ZN(n986) );
NOR4_X1 U716 ( .A1(n991), .A2(n992), .A3(n993), .A4(n994), .ZN(n989) );
NOR4_X1 U717 ( .A1(n995), .A2(n996), .A3(n997), .A4(n998), .ZN(n992) );
NOR2_X1 U718 ( .A1(n999), .A2(n1000), .ZN(n998) );
INV_X1 U719 ( .A(KEYINPUT26), .ZN(n1000) );
NOR2_X1 U720 ( .A1(KEYINPUT14), .A2(n1001), .ZN(n997) );
NAND2_X1 U721 ( .A1(n1002), .A2(n1003), .ZN(n996) );
NAND2_X1 U722 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NOR3_X1 U723 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n991) );
NOR2_X1 U724 ( .A1(KEYINPUT26), .A2(n999), .ZN(n1008) );
NAND3_X1 U725 ( .A1(n1004), .A2(n1009), .A3(n1010), .ZN(n999) );
NOR2_X1 U726 ( .A1(n1001), .A2(n1011), .ZN(n1007) );
INV_X1 U727 ( .A(KEYINPUT14), .ZN(n1011) );
NAND3_X1 U728 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1001) );
NAND3_X1 U729 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n987) );
NAND4_X1 U730 ( .A1(n1006), .A2(n1014), .A3(n1004), .A4(n1018), .ZN(n1017) );
NAND2_X1 U731 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND2_X1 U732 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
OR2_X1 U733 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U734 ( .A1(n1025), .A2(n1026), .ZN(n1019) );
NAND2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND2_X1 U736 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
INV_X1 U737 ( .A(n995), .ZN(n1006) );
NOR3_X1 U738 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n985) );
INV_X1 U739 ( .A(n1015), .ZN(n1031) );
NAND4_X1 U740 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1015) );
NOR4_X1 U741 ( .A1(n1010), .A2(n1029), .A3(n1036), .A4(n1037), .ZN(n1035) );
XOR2_X1 U742 ( .A(n1038), .B(n1039), .Z(n1036) );
XOR2_X1 U743 ( .A(KEYINPUT1), .B(n1040), .Z(n1039) );
NOR2_X1 U744 ( .A1(KEYINPUT46), .A2(G469), .ZN(n1040) );
NOR2_X1 U745 ( .A1(n1013), .A2(n1041), .ZN(n1034) );
XOR2_X1 U746 ( .A(n1042), .B(KEYINPUT6), .Z(n1033) );
NAND2_X1 U747 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND2_X1 U748 ( .A1(G472), .A2(n1045), .ZN(n1044) );
XOR2_X1 U749 ( .A(n1046), .B(KEYINPUT18), .Z(n1043) );
OR2_X1 U750 ( .A1(n1045), .A2(G472), .ZN(n1046) );
XOR2_X1 U751 ( .A(n1047), .B(G475), .Z(n1032) );
XOR2_X1 U752 ( .A(n1048), .B(n1049), .Z(G72) );
NOR2_X1 U753 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
XNOR2_X1 U755 ( .A(G227), .B(KEYINPUT42), .ZN(n1052) );
NAND3_X1 U756 ( .A1(n1054), .A2(n1055), .A3(KEYINPUT41), .ZN(n1048) );
NAND2_X1 U757 ( .A1(n1056), .A2(n1016), .ZN(n1055) );
XOR2_X1 U758 ( .A(n990), .B(n1057), .Z(n1056) );
NAND3_X1 U759 ( .A1(G900), .A2(n1057), .A3(G953), .ZN(n1054) );
XOR2_X1 U760 ( .A(n1058), .B(n1059), .Z(n1057) );
XOR2_X1 U761 ( .A(n1060), .B(n1061), .Z(n1059) );
NOR2_X1 U762 ( .A1(KEYINPUT25), .A2(n1062), .ZN(n1061) );
XOR2_X1 U763 ( .A(n1063), .B(n1064), .Z(n1058) );
NAND2_X1 U764 ( .A1(KEYINPUT50), .A2(n1065), .ZN(n1063) );
XOR2_X1 U765 ( .A(n1066), .B(n1067), .Z(G69) );
XOR2_X1 U766 ( .A(n1068), .B(n1069), .Z(n1067) );
NOR2_X1 U767 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U768 ( .A(n1016), .B(KEYINPUT20), .Z(n1071) );
INV_X1 U769 ( .A(n988), .ZN(n1070) );
NAND3_X1 U770 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1068) );
XOR2_X1 U771 ( .A(n1075), .B(KEYINPUT62), .Z(n1074) );
NAND2_X1 U772 ( .A1(G953), .A2(n1076), .ZN(n1075) );
XOR2_X1 U773 ( .A(KEYINPUT53), .B(n1077), .Z(n1072) );
NOR2_X1 U774 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1080), .A2(n1081), .ZN(n1066) );
NAND2_X1 U776 ( .A1(G898), .A2(G224), .ZN(n1081) );
INV_X1 U777 ( .A(n1051), .ZN(n1080) );
XOR2_X1 U778 ( .A(n1016), .B(KEYINPUT27), .Z(n1051) );
NOR2_X1 U779 ( .A1(n1082), .A2(n1083), .ZN(G66) );
XOR2_X1 U780 ( .A(n1084), .B(n1085), .Z(n1083) );
XOR2_X1 U781 ( .A(KEYINPUT9), .B(KEYINPUT39), .Z(n1085) );
XOR2_X1 U782 ( .A(n1086), .B(n1087), .Z(n1084) );
NAND2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
NOR2_X1 U784 ( .A1(n1082), .A2(n1090), .ZN(G63) );
XOR2_X1 U785 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U786 ( .A1(n1088), .A2(G478), .ZN(n1092) );
NOR2_X1 U787 ( .A1(n1082), .A2(n1093), .ZN(G60) );
XOR2_X1 U788 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U789 ( .A1(KEYINPUT43), .A2(n1096), .ZN(n1095) );
NAND2_X1 U790 ( .A1(n1088), .A2(G475), .ZN(n1094) );
XOR2_X1 U791 ( .A(G104), .B(n1097), .Z(G6) );
NOR2_X1 U792 ( .A1(n1082), .A2(n1098), .ZN(G57) );
XOR2_X1 U793 ( .A(n1099), .B(n1100), .Z(n1098) );
XOR2_X1 U794 ( .A(n1101), .B(n1102), .Z(n1100) );
XOR2_X1 U795 ( .A(n1103), .B(n1104), .Z(n1101) );
NOR2_X1 U796 ( .A1(KEYINPUT8), .A2(n1105), .ZN(n1104) );
NAND2_X1 U797 ( .A1(n1088), .A2(G472), .ZN(n1103) );
XNOR2_X1 U798 ( .A(n1106), .B(n1107), .ZN(n1099) );
XOR2_X1 U799 ( .A(KEYINPUT11), .B(G101), .Z(n1107) );
NOR2_X1 U800 ( .A1(n1082), .A2(n1108), .ZN(G54) );
XOR2_X1 U801 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U802 ( .A1(n1088), .A2(G469), .ZN(n1110) );
NAND2_X1 U803 ( .A1(n1111), .A2(KEYINPUT13), .ZN(n1109) );
XOR2_X1 U804 ( .A(n1112), .B(n1113), .Z(n1111) );
XNOR2_X1 U805 ( .A(n1114), .B(n1115), .ZN(n1113) );
XOR2_X1 U806 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND2_X1 U807 ( .A1(KEYINPUT16), .A2(n1118), .ZN(n1116) );
XOR2_X1 U808 ( .A(n1119), .B(n1120), .Z(n1112) );
XOR2_X1 U809 ( .A(KEYINPUT37), .B(G140), .Z(n1120) );
XOR2_X1 U810 ( .A(n1121), .B(n1122), .Z(n1119) );
NOR2_X1 U811 ( .A1(KEYINPUT12), .A2(n1123), .ZN(n1122) );
XOR2_X1 U812 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U813 ( .A1(n1082), .A2(n1126), .ZN(G51) );
NOR2_X1 U814 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U815 ( .A(KEYINPUT36), .B(n1129), .Z(n1128) );
NOR2_X1 U816 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
AND2_X1 U817 ( .A1(n1131), .A2(n1130), .ZN(n1127) );
XOR2_X1 U818 ( .A(n1132), .B(n1133), .Z(n1130) );
NOR2_X1 U819 ( .A1(n1134), .A2(KEYINPUT38), .ZN(n1133) );
NOR2_X1 U820 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XOR2_X1 U821 ( .A(n1137), .B(KEYINPUT24), .Z(n1136) );
XNOR2_X1 U822 ( .A(n1138), .B(n1139), .ZN(n1132) );
NAND2_X1 U823 ( .A1(n1088), .A2(n1140), .ZN(n1131) );
AND2_X1 U824 ( .A1(G902), .A2(n1141), .ZN(n1088) );
NAND2_X1 U825 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
INV_X1 U826 ( .A(n990), .ZN(n1143) );
NAND4_X1 U827 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n990) );
AND3_X1 U828 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NAND2_X1 U829 ( .A1(n1151), .A2(n1152), .ZN(n1146) );
NAND2_X1 U830 ( .A1(n1153), .A2(n1154), .ZN(n1144) );
NAND3_X1 U831 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1154) );
NAND2_X1 U832 ( .A1(n1021), .A2(n1025), .ZN(n1157) );
NAND2_X1 U833 ( .A1(n1158), .A2(n1024), .ZN(n1156) );
XOR2_X1 U834 ( .A(n1027), .B(KEYINPUT32), .Z(n1158) );
NAND2_X1 U835 ( .A1(n1023), .A2(n1159), .ZN(n1155) );
XOR2_X1 U836 ( .A(KEYINPUT63), .B(n1152), .Z(n1159) );
XOR2_X1 U837 ( .A(n988), .B(KEYINPUT4), .Z(n1142) );
NAND2_X1 U838 ( .A1(n1160), .A2(n1161), .ZN(n988) );
AND4_X1 U839 ( .A1(n1162), .A2(n984), .A3(n1163), .A4(n1164), .ZN(n1161) );
NAND3_X1 U840 ( .A1(n1024), .A2(n1004), .A3(n1165), .ZN(n984) );
NOR4_X1 U841 ( .A1(n1166), .A2(n1097), .A3(n1167), .A4(n1168), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1027), .A2(n1169), .ZN(n1168) );
NOR4_X1 U843 ( .A1(n1170), .A2(n1002), .A3(n1171), .A4(n1172), .ZN(n1167) );
XOR2_X1 U844 ( .A(KEYINPUT58), .B(n1173), .Z(n1172) );
AND3_X1 U845 ( .A1(n1165), .A2(n1004), .A3(n1023), .ZN(n1097) );
NOR2_X1 U846 ( .A1(n1016), .A2(G952), .ZN(n1082) );
XNOR2_X1 U847 ( .A(G146), .B(n1174), .ZN(G48) );
NAND2_X1 U848 ( .A1(n1175), .A2(n1023), .ZN(n1174) );
XOR2_X1 U849 ( .A(G143), .B(n1176), .Z(G45) );
NOR2_X1 U850 ( .A1(n1027), .A2(n1177), .ZN(n1176) );
XOR2_X1 U851 ( .A(KEYINPUT51), .B(n1151), .Z(n1177) );
AND4_X1 U852 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1041), .ZN(n1151) );
INV_X1 U853 ( .A(n1181), .ZN(n1041) );
XNOR2_X1 U854 ( .A(G140), .B(n1145), .ZN(G42) );
NAND2_X1 U855 ( .A1(n1182), .A2(n1183), .ZN(n1145) );
XOR2_X1 U856 ( .A(n1184), .B(n1185), .Z(G39) );
NAND3_X1 U857 ( .A1(n1021), .A2(n1025), .A3(n1153), .ZN(n1185) );
XNOR2_X1 U858 ( .A(G134), .B(n1148), .ZN(G36) );
NAND3_X1 U859 ( .A1(n1180), .A2(n1024), .A3(n1182), .ZN(n1148) );
XNOR2_X1 U860 ( .A(G131), .B(n1150), .ZN(G33) );
NAND3_X1 U861 ( .A1(n1023), .A2(n1180), .A3(n1182), .ZN(n1150) );
AND2_X1 U862 ( .A1(n1021), .A2(n1179), .ZN(n1182) );
INV_X1 U863 ( .A(n994), .ZN(n1021) );
NAND2_X1 U864 ( .A1(n1030), .A2(n1186), .ZN(n994) );
XOR2_X1 U865 ( .A(n1124), .B(n1187), .Z(G30) );
NAND2_X1 U866 ( .A1(n1175), .A2(n1024), .ZN(n1187) );
AND2_X1 U867 ( .A1(n1153), .A2(n1152), .ZN(n1175) );
AND3_X1 U868 ( .A1(n1188), .A2(n1013), .A3(n1179), .ZN(n1153) );
AND2_X1 U869 ( .A1(n1005), .A2(n1189), .ZN(n1179) );
XOR2_X1 U870 ( .A(G101), .B(n1166), .Z(G3) );
AND3_X1 U871 ( .A1(n1025), .A2(n1165), .A3(n1180), .ZN(n1166) );
XNOR2_X1 U872 ( .A(G125), .B(n1149), .ZN(G27) );
NAND4_X1 U873 ( .A1(n1183), .A2(n1014), .A3(n1152), .A4(n1189), .ZN(n1149) );
NAND2_X1 U874 ( .A1(n995), .A2(n1190), .ZN(n1189) );
NAND2_X1 U875 ( .A1(n1191), .A2(n1053), .ZN(n1190) );
INV_X1 U876 ( .A(G900), .ZN(n1053) );
AND3_X1 U877 ( .A1(n1012), .A2(n1013), .A3(n1023), .ZN(n1183) );
XOR2_X1 U878 ( .A(G122), .B(n1192), .Z(G24) );
NOR2_X1 U879 ( .A1(n1027), .A2(n1193), .ZN(n1192) );
XNOR2_X1 U880 ( .A(KEYINPUT5), .B(n1169), .ZN(n1193) );
NAND4_X1 U881 ( .A1(n1178), .A2(n1014), .A3(n1194), .A4(n1004), .ZN(n1169) );
NOR2_X1 U882 ( .A1(n1013), .A2(n1188), .ZN(n1004) );
NOR2_X1 U883 ( .A1(n1170), .A2(n1181), .ZN(n1194) );
XOR2_X1 U884 ( .A(n1162), .B(n1195), .Z(G21) );
XOR2_X1 U885 ( .A(KEYINPUT55), .B(G119), .Z(n1195) );
NAND4_X1 U886 ( .A1(n1188), .A2(n1014), .A3(n1025), .A4(n1196), .ZN(n1162) );
AND3_X1 U887 ( .A1(n1152), .A2(n1197), .A3(n1013), .ZN(n1196) );
XOR2_X1 U888 ( .A(n1198), .B(n1164), .Z(G18) );
NAND4_X1 U889 ( .A1(n1199), .A2(n1024), .A3(n1152), .A4(n1197), .ZN(n1164) );
INV_X1 U890 ( .A(n1027), .ZN(n1152) );
XNOR2_X1 U891 ( .A(n1173), .B(KEYINPUT23), .ZN(n1027) );
NOR2_X1 U892 ( .A1(n1178), .A2(n1181), .ZN(n1024) );
XNOR2_X1 U893 ( .A(G113), .B(n1200), .ZN(G15) );
NAND4_X1 U894 ( .A1(n1023), .A2(n1199), .A3(n1173), .A4(n1201), .ZN(n1200) );
XOR2_X1 U895 ( .A(KEYINPUT28), .B(n1170), .Z(n1201) );
INV_X1 U896 ( .A(n1197), .ZN(n1170) );
INV_X1 U897 ( .A(n1002), .ZN(n1199) );
NAND2_X1 U898 ( .A1(n1180), .A2(n1014), .ZN(n1002) );
AND2_X1 U899 ( .A1(n1009), .A2(n1202), .ZN(n1014) );
NOR2_X1 U900 ( .A1(n1012), .A2(n1013), .ZN(n1180) );
INV_X1 U901 ( .A(n1171), .ZN(n1023) );
NAND2_X1 U902 ( .A1(n1178), .A2(n1181), .ZN(n1171) );
XOR2_X1 U903 ( .A(n1118), .B(n1163), .Z(G12) );
NAND4_X1 U904 ( .A1(n1025), .A2(n1165), .A3(n1012), .A4(n1013), .ZN(n1163) );
XNOR2_X1 U905 ( .A(n1203), .B(n1089), .ZN(n1013) );
AND2_X1 U906 ( .A1(G217), .A2(n1204), .ZN(n1089) );
OR2_X1 U907 ( .A1(n1087), .A2(G902), .ZN(n1203) );
XNOR2_X1 U908 ( .A(n1205), .B(n1206), .ZN(n1087) );
XOR2_X1 U909 ( .A(n1184), .B(n1207), .Z(n1206) );
NAND2_X1 U910 ( .A1(n1208), .A2(n1209), .ZN(n1207) );
NAND2_X1 U911 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
XOR2_X1 U912 ( .A(n1212), .B(KEYINPUT59), .Z(n1208) );
OR2_X1 U913 ( .A1(n1211), .A2(n1210), .ZN(n1212) );
XNOR2_X1 U914 ( .A(n1213), .B(n1065), .ZN(n1210) );
XNOR2_X1 U915 ( .A(G140), .B(G125), .ZN(n1065) );
XNOR2_X1 U916 ( .A(G146), .B(KEYINPUT60), .ZN(n1213) );
XNOR2_X1 U917 ( .A(n1214), .B(n1215), .ZN(n1211) );
NOR2_X1 U918 ( .A1(KEYINPUT21), .A2(G110), .ZN(n1215) );
XOR2_X1 U919 ( .A(G119), .B(n1124), .Z(n1214) );
INV_X1 U920 ( .A(G137), .ZN(n1184) );
NAND3_X1 U921 ( .A1(G221), .A2(G234), .A3(n1216), .ZN(n1205) );
INV_X1 U922 ( .A(n1188), .ZN(n1012) );
XNOR2_X1 U923 ( .A(G472), .B(n1217), .ZN(n1188) );
NOR2_X1 U924 ( .A1(n1218), .A2(KEYINPUT44), .ZN(n1217) );
INV_X1 U925 ( .A(n1045), .ZN(n1218) );
NAND2_X1 U926 ( .A1(n1219), .A2(n1220), .ZN(n1045) );
XOR2_X1 U927 ( .A(n1221), .B(n1222), .Z(n1219) );
XOR2_X1 U928 ( .A(n1102), .B(n1105), .Z(n1222) );
XNOR2_X1 U929 ( .A(n1223), .B(n1224), .ZN(n1102) );
XNOR2_X1 U930 ( .A(KEYINPUT34), .B(n1225), .ZN(n1221) );
NOR2_X1 U931 ( .A1(KEYINPUT31), .A2(n1226), .ZN(n1225) );
XNOR2_X1 U932 ( .A(G101), .B(n1227), .ZN(n1226) );
NAND2_X1 U933 ( .A1(KEYINPUT19), .A2(n1106), .ZN(n1227) );
AND3_X1 U934 ( .A1(n1216), .A2(n1228), .A3(G210), .ZN(n1106) );
AND3_X1 U935 ( .A1(n1173), .A2(n1197), .A3(n1005), .ZN(n1165) );
NOR2_X1 U936 ( .A1(n1009), .A2(n1010), .ZN(n1005) );
INV_X1 U937 ( .A(n1202), .ZN(n1010) );
NAND2_X1 U938 ( .A1(G221), .A2(n1204), .ZN(n1202) );
NAND2_X1 U939 ( .A1(G234), .A2(n1220), .ZN(n1204) );
XNOR2_X1 U940 ( .A(n1038), .B(n1229), .ZN(n1009) );
XOR2_X1 U941 ( .A(KEYINPUT10), .B(G469), .Z(n1229) );
NAND2_X1 U942 ( .A1(n1230), .A2(n1220), .ZN(n1038) );
XOR2_X1 U943 ( .A(n1231), .B(n1232), .Z(n1230) );
XNOR2_X1 U944 ( .A(n1233), .B(KEYINPUT3), .ZN(n1232) );
NAND2_X1 U945 ( .A1(KEYINPUT22), .A2(n1234), .ZN(n1233) );
XOR2_X1 U946 ( .A(n1117), .B(n1235), .Z(n1234) );
XOR2_X1 U947 ( .A(G140), .B(G110), .Z(n1235) );
AND2_X1 U948 ( .A1(G227), .A2(n1216), .ZN(n1117) );
XOR2_X1 U949 ( .A(n1223), .B(n1125), .Z(n1231) );
XNOR2_X1 U950 ( .A(n1236), .B(n1237), .ZN(n1125) );
XOR2_X1 U951 ( .A(G101), .B(n1060), .Z(n1237) );
NOR2_X1 U952 ( .A1(KEYINPUT56), .A2(n1224), .ZN(n1060) );
XOR2_X1 U953 ( .A(n1064), .B(n1121), .Z(n1223) );
NAND2_X1 U954 ( .A1(KEYINPUT30), .A2(n1062), .ZN(n1121) );
XOR2_X1 U955 ( .A(G134), .B(KEYINPUT47), .Z(n1062) );
XOR2_X1 U956 ( .A(G128), .B(n1114), .Z(n1064) );
XOR2_X1 U957 ( .A(G131), .B(G137), .Z(n1114) );
NAND2_X1 U958 ( .A1(n995), .A2(n1238), .ZN(n1197) );
NAND2_X1 U959 ( .A1(n1191), .A2(n1076), .ZN(n1238) );
INV_X1 U960 ( .A(G898), .ZN(n1076) );
AND3_X1 U961 ( .A1(G953), .A2(n1239), .A3(n1240), .ZN(n1191) );
XOR2_X1 U962 ( .A(n1220), .B(KEYINPUT61), .Z(n1240) );
NAND3_X1 U963 ( .A1(n1239), .A2(n1016), .A3(G952), .ZN(n995) );
NAND2_X1 U964 ( .A1(G237), .A2(G234), .ZN(n1239) );
NOR2_X1 U965 ( .A1(n1030), .A2(n1029), .ZN(n1173) );
INV_X1 U966 ( .A(n1186), .ZN(n1029) );
NAND2_X1 U967 ( .A1(G214), .A2(n1241), .ZN(n1186) );
XOR2_X1 U968 ( .A(n1037), .B(KEYINPUT54), .Z(n1030) );
XNOR2_X1 U969 ( .A(n1242), .B(n1140), .ZN(n1037) );
AND2_X1 U970 ( .A1(G210), .A2(n1241), .ZN(n1140) );
NAND2_X1 U971 ( .A1(n1243), .A2(n1228), .ZN(n1241) );
XOR2_X1 U972 ( .A(n1220), .B(KEYINPUT52), .Z(n1243) );
NAND2_X1 U973 ( .A1(n1244), .A2(n1220), .ZN(n1242) );
XOR2_X1 U974 ( .A(n1139), .B(n1245), .Z(n1244) );
XOR2_X1 U975 ( .A(n1138), .B(n1246), .Z(n1245) );
NOR2_X1 U976 ( .A1(n1135), .A2(n1247), .ZN(n1246) );
XOR2_X1 U977 ( .A(n1137), .B(KEYINPUT7), .Z(n1247) );
NAND2_X1 U978 ( .A1(G125), .A2(n1248), .ZN(n1137) );
NOR2_X1 U979 ( .A1(G125), .A2(n1248), .ZN(n1135) );
XOR2_X1 U980 ( .A(n1124), .B(n1224), .Z(n1248) );
NAND2_X1 U981 ( .A1(n1073), .A2(n1249), .ZN(n1138) );
OR2_X1 U982 ( .A1(n1079), .A2(n1078), .ZN(n1249) );
NAND2_X1 U983 ( .A1(n1078), .A2(n1079), .ZN(n1073) );
XNOR2_X1 U984 ( .A(n1250), .B(n1251), .ZN(n1079) );
XOR2_X1 U985 ( .A(KEYINPUT57), .B(G110), .Z(n1251) );
NAND2_X1 U986 ( .A1(KEYINPUT49), .A2(n1252), .ZN(n1250) );
XNOR2_X1 U987 ( .A(n1253), .B(n1105), .ZN(n1078) );
XNOR2_X1 U988 ( .A(G113), .B(n1254), .ZN(n1105) );
XOR2_X1 U989 ( .A(G119), .B(G116), .Z(n1254) );
XOR2_X1 U990 ( .A(n1255), .B(G101), .Z(n1253) );
NAND2_X1 U991 ( .A1(KEYINPUT40), .A2(n1236), .ZN(n1255) );
XOR2_X1 U992 ( .A(G104), .B(n1256), .Z(n1236) );
NAND2_X1 U993 ( .A1(G224), .A2(n1216), .ZN(n1139) );
INV_X1 U994 ( .A(n993), .ZN(n1025) );
NAND2_X1 U995 ( .A1(n1181), .A2(n1257), .ZN(n993) );
INV_X1 U996 ( .A(n1178), .ZN(n1257) );
XOR2_X1 U997 ( .A(n1047), .B(n1258), .Z(n1178) );
NOR2_X1 U998 ( .A1(G475), .A2(KEYINPUT45), .ZN(n1258) );
OR2_X1 U999 ( .A1(n1096), .A2(G902), .ZN(n1047) );
XOR2_X1 U1000 ( .A(n1259), .B(n1260), .Z(n1096) );
XOR2_X1 U1001 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U1002 ( .A(n1263), .B(n1264), .Z(n1262) );
XNOR2_X1 U1003 ( .A(G104), .B(n1265), .ZN(n1264) );
NOR2_X1 U1004 ( .A1(KEYINPUT2), .A2(G125), .ZN(n1265) );
XOR2_X1 U1005 ( .A(G113), .B(n1252), .Z(n1263) );
INV_X1 U1006 ( .A(G122), .ZN(n1252) );
XOR2_X1 U1007 ( .A(n1266), .B(n1267), .Z(n1261) );
XOR2_X1 U1008 ( .A(G140), .B(G131), .Z(n1267) );
XOR2_X1 U1009 ( .A(KEYINPUT60), .B(KEYINPUT33), .Z(n1266) );
XNOR2_X1 U1010 ( .A(n1224), .B(n1268), .ZN(n1259) );
AND3_X1 U1011 ( .A1(G214), .A2(n1228), .A3(n1216), .ZN(n1268) );
INV_X1 U1012 ( .A(G237), .ZN(n1228) );
XOR2_X1 U1013 ( .A(G146), .B(G143), .Z(n1224) );
XNOR2_X1 U1014 ( .A(G478), .B(n1269), .ZN(n1181) );
AND2_X1 U1015 ( .A1(n1091), .A2(n1220), .ZN(n1269) );
INV_X1 U1016 ( .A(G902), .ZN(n1220) );
NAND2_X1 U1017 ( .A1(n1270), .A2(n1271), .ZN(n1091) );
NAND2_X1 U1018 ( .A1(n1272), .A2(n1273), .ZN(n1271) );
XOR2_X1 U1019 ( .A(KEYINPUT48), .B(n1274), .Z(n1270) );
NOR2_X1 U1020 ( .A1(n1272), .A2(n1273), .ZN(n1274) );
NAND3_X1 U1021 ( .A1(n1216), .A2(G234), .A3(G217), .ZN(n1273) );
XOR2_X1 U1022 ( .A(n1016), .B(KEYINPUT15), .Z(n1216) );
INV_X1 U1023 ( .A(G953), .ZN(n1016) );
XOR2_X1 U1024 ( .A(n1275), .B(n1276), .Z(n1272) );
XOR2_X1 U1025 ( .A(n1277), .B(n1278), .Z(n1276) );
NAND2_X1 U1026 ( .A1(KEYINPUT29), .A2(n1256), .ZN(n1278) );
XNOR2_X1 U1027 ( .A(G107), .B(KEYINPUT35), .ZN(n1256) );
NAND3_X1 U1028 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1277) );
NAND2_X1 U1029 ( .A1(G143), .A2(n1282), .ZN(n1281) );
OR3_X1 U1030 ( .A1(n1282), .A2(G143), .A3(KEYINPUT0), .ZN(n1280) );
NAND2_X1 U1031 ( .A1(KEYINPUT17), .A2(n1124), .ZN(n1282) );
INV_X1 U1032 ( .A(G128), .ZN(n1124) );
NAND2_X1 U1033 ( .A1(G128), .A2(KEYINPUT0), .ZN(n1279) );
XOR2_X1 U1034 ( .A(n1198), .B(n1283), .Z(n1275) );
XOR2_X1 U1035 ( .A(G134), .B(G122), .Z(n1283) );
INV_X1 U1036 ( .A(G116), .ZN(n1198) );
INV_X1 U1037 ( .A(G110), .ZN(n1118) );
endmodule


