//Key = 1110000111100001100110011101011110011101001000000011111101100111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423;

XNOR2_X1 U790 ( .A(G107), .B(n1094), .ZN(G9) );
NAND2_X1 U791 ( .A1(KEYINPUT19), .A2(n1095), .ZN(n1094) );
NOR2_X1 U792 ( .A1(n1096), .A2(n1097), .ZN(G75) );
NOR4_X1 U793 ( .A1(G953), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1097) );
NOR2_X1 U794 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U795 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NOR3_X1 U796 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1104) );
NOR2_X1 U797 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NOR2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(n1110) );
NOR2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NOR2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1112) );
NOR2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NOR4_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1115), .A4(n1122), .ZN(n1108) );
NOR3_X1 U804 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1121) );
NOR2_X1 U805 ( .A1(n1126), .A2(n1127), .ZN(n1120) );
NOR3_X1 U806 ( .A1(n1111), .A2(n1116), .A3(n1128), .ZN(n1103) );
NOR2_X1 U807 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NOR2_X1 U808 ( .A1(n1131), .A2(n1115), .ZN(n1129) );
NOR2_X1 U809 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NOR2_X1 U810 ( .A1(n1105), .A2(n1134), .ZN(n1133) );
NOR2_X1 U811 ( .A1(KEYINPUT47), .A2(n1135), .ZN(n1132) );
AND2_X1 U812 ( .A1(n1130), .A2(n1136), .ZN(n1116) );
NAND3_X1 U813 ( .A1(n1137), .A2(n1138), .A3(KEYINPUT47), .ZN(n1136) );
NOR3_X1 U814 ( .A1(n1098), .A2(G953), .A3(G952), .ZN(n1096) );
AND4_X1 U815 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1098) );
NOR3_X1 U816 ( .A1(n1143), .A2(n1106), .A3(n1144), .ZN(n1142) );
NOR2_X1 U817 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XNOR2_X1 U818 ( .A(G469), .B(KEYINPUT28), .ZN(n1146) );
AND2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
NAND3_X1 U820 ( .A1(n1149), .A2(n1150), .A3(n1127), .ZN(n1143) );
NOR3_X1 U821 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1141) );
XNOR2_X1 U822 ( .A(n1154), .B(n1155), .ZN(n1153) );
XNOR2_X1 U823 ( .A(KEYINPUT50), .B(n1156), .ZN(n1155) );
XNOR2_X1 U824 ( .A(n1157), .B(KEYINPUT25), .ZN(n1152) );
XOR2_X1 U825 ( .A(n1158), .B(n1159), .Z(n1151) );
NOR2_X1 U826 ( .A1(KEYINPUT33), .A2(n1160), .ZN(n1159) );
XNOR2_X1 U827 ( .A(G472), .B(KEYINPUT39), .ZN(n1158) );
XOR2_X1 U828 ( .A(n1161), .B(KEYINPUT14), .Z(n1139) );
XOR2_X1 U829 ( .A(n1162), .B(n1163), .Z(G72) );
NOR3_X1 U830 ( .A1(n1164), .A2(KEYINPUT11), .A3(n1165), .ZN(n1163) );
AND2_X1 U831 ( .A1(G227), .A2(G900), .ZN(n1165) );
NAND2_X1 U832 ( .A1(n1166), .A2(n1167), .ZN(n1162) );
NAND2_X1 U833 ( .A1(n1168), .A2(n1164), .ZN(n1167) );
XOR2_X1 U834 ( .A(n1169), .B(n1170), .Z(n1168) );
NAND3_X1 U835 ( .A1(n1170), .A2(G900), .A3(G953), .ZN(n1166) );
NOR3_X1 U836 ( .A1(KEYINPUT56), .A2(n1171), .A3(n1172), .ZN(n1170) );
XOR2_X1 U837 ( .A(n1173), .B(KEYINPUT24), .Z(n1172) );
NAND2_X1 U838 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U839 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
XOR2_X1 U840 ( .A(n1176), .B(n1177), .Z(n1175) );
NAND2_X1 U841 ( .A1(n1178), .A2(KEYINPUT63), .ZN(n1176) );
XNOR2_X1 U842 ( .A(G137), .B(n1179), .ZN(n1178) );
XOR2_X1 U843 ( .A(n1180), .B(n1181), .Z(G69) );
XOR2_X1 U844 ( .A(n1182), .B(n1183), .Z(n1181) );
NAND2_X1 U845 ( .A1(G953), .A2(n1184), .ZN(n1183) );
NAND2_X1 U846 ( .A1(G898), .A2(G224), .ZN(n1184) );
NAND2_X1 U847 ( .A1(n1185), .A2(n1186), .ZN(n1182) );
NAND2_X1 U848 ( .A1(G953), .A2(n1187), .ZN(n1186) );
XNOR2_X1 U849 ( .A(n1188), .B(n1189), .ZN(n1185) );
NAND2_X1 U850 ( .A1(KEYINPUT20), .A2(n1190), .ZN(n1188) );
AND2_X1 U851 ( .A1(n1191), .A2(n1164), .ZN(n1180) );
NOR3_X1 U852 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(G66) );
AND2_X1 U853 ( .A1(KEYINPUT27), .A2(n1195), .ZN(n1194) );
NOR3_X1 U854 ( .A1(KEYINPUT27), .A2(n1196), .A3(n1164), .ZN(n1193) );
INV_X1 U855 ( .A(G952), .ZN(n1196) );
XOR2_X1 U856 ( .A(n1197), .B(n1198), .Z(n1192) );
NOR2_X1 U857 ( .A1(n1199), .A2(n1200), .ZN(n1197) );
NOR2_X1 U858 ( .A1(n1195), .A2(n1201), .ZN(G63) );
XOR2_X1 U859 ( .A(n1202), .B(n1203), .Z(n1201) );
NOR2_X1 U860 ( .A1(n1204), .A2(n1200), .ZN(n1202) );
NOR2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(G60) );
XNOR2_X1 U862 ( .A(n1195), .B(KEYINPUT42), .ZN(n1206) );
NOR3_X1 U863 ( .A1(n1154), .A2(n1207), .A3(n1208), .ZN(n1205) );
NOR3_X1 U864 ( .A1(n1209), .A2(n1156), .A3(n1200), .ZN(n1208) );
INV_X1 U865 ( .A(n1210), .ZN(n1209) );
NOR2_X1 U866 ( .A1(n1211), .A2(n1210), .ZN(n1207) );
NOR2_X1 U867 ( .A1(n1212), .A2(n1156), .ZN(n1211) );
XNOR2_X1 U868 ( .A(G104), .B(n1213), .ZN(G6) );
NOR2_X1 U869 ( .A1(n1195), .A2(n1214), .ZN(G57) );
XOR2_X1 U870 ( .A(n1215), .B(n1216), .Z(n1214) );
NAND2_X1 U871 ( .A1(KEYINPUT0), .A2(n1217), .ZN(n1215) );
XOR2_X1 U872 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U873 ( .A(n1220), .B(n1221), .Z(n1218) );
NOR2_X1 U874 ( .A1(n1222), .A2(n1200), .ZN(n1221) );
NAND2_X1 U875 ( .A1(KEYINPUT2), .A2(n1223), .ZN(n1220) );
NOR3_X1 U876 ( .A1(n1195), .A2(n1224), .A3(n1225), .ZN(G54) );
NOR4_X1 U877 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1200), .ZN(n1225) );
INV_X1 U878 ( .A(n1229), .ZN(n1226) );
NOR2_X1 U879 ( .A1(n1229), .A2(n1230), .ZN(n1224) );
NOR3_X1 U880 ( .A1(n1200), .A2(n1231), .A3(n1228), .ZN(n1230) );
AND2_X1 U881 ( .A1(n1227), .A2(n1232), .ZN(n1231) );
INV_X1 U882 ( .A(KEYINPUT7), .ZN(n1227) );
NAND2_X1 U883 ( .A1(G902), .A2(n1100), .ZN(n1200) );
INV_X1 U884 ( .A(n1212), .ZN(n1100) );
NOR2_X1 U885 ( .A1(KEYINPUT34), .A2(n1232), .ZN(n1229) );
NAND2_X1 U886 ( .A1(n1233), .A2(n1234), .ZN(n1232) );
OR2_X1 U887 ( .A1(n1148), .A2(KEYINPUT18), .ZN(n1234) );
NAND2_X1 U888 ( .A1(KEYINPUT18), .A2(n1235), .ZN(n1233) );
NAND2_X1 U889 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
OR2_X1 U890 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
NOR2_X1 U891 ( .A1(n1195), .A2(n1240), .ZN(G51) );
XOR2_X1 U892 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U893 ( .A1(KEYINPUT49), .A2(n1243), .ZN(n1242) );
XOR2_X1 U894 ( .A(n1244), .B(n1245), .Z(n1243) );
XNOR2_X1 U895 ( .A(n1246), .B(n1247), .ZN(n1245) );
NAND2_X1 U896 ( .A1(KEYINPUT30), .A2(n1248), .ZN(n1247) );
NAND2_X1 U897 ( .A1(KEYINPUT9), .A2(n1249), .ZN(n1246) );
XNOR2_X1 U898 ( .A(G125), .B(n1250), .ZN(n1244) );
NOR3_X1 U899 ( .A1(n1251), .A2(KEYINPUT48), .A3(G953), .ZN(n1250) );
INV_X1 U900 ( .A(G224), .ZN(n1251) );
NAND3_X1 U901 ( .A1(G902), .A2(G210), .A3(n1252), .ZN(n1241) );
XNOR2_X1 U902 ( .A(n1212), .B(KEYINPUT22), .ZN(n1252) );
NOR2_X1 U903 ( .A1(n1191), .A2(n1169), .ZN(n1212) );
NAND4_X1 U904 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1169) );
NOR4_X1 U905 ( .A1(n1257), .A2(n1258), .A3(n1259), .A4(n1260), .ZN(n1256) );
NOR3_X1 U906 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1255) );
NOR2_X1 U907 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
AND3_X1 U908 ( .A1(n1264), .A2(n1266), .A3(KEYINPUT12), .ZN(n1262) );
NOR2_X1 U909 ( .A1(KEYINPUT12), .A2(n1267), .ZN(n1261) );
NAND4_X1 U910 ( .A1(n1213), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1191) );
NOR4_X1 U911 ( .A1(n1271), .A2(n1272), .A3(n1095), .A4(n1273), .ZN(n1270) );
NOR2_X1 U912 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
NOR2_X1 U913 ( .A1(n1276), .A2(n1277), .ZN(n1274) );
NOR2_X1 U914 ( .A1(n1111), .A2(n1278), .ZN(n1277) );
NOR2_X1 U915 ( .A1(n1279), .A2(n1280), .ZN(n1276) );
XNOR2_X1 U916 ( .A(n1125), .B(KEYINPUT40), .ZN(n1279) );
AND3_X1 U917 ( .A1(n1281), .A2(n1126), .A3(n1118), .ZN(n1095) );
AND3_X1 U918 ( .A1(KEYINPUT5), .A2(n1282), .A3(n1283), .ZN(n1272) );
NOR2_X1 U919 ( .A1(KEYINPUT5), .A2(n1284), .ZN(n1271) );
NOR2_X1 U920 ( .A1(n1285), .A2(n1286), .ZN(n1269) );
NAND3_X1 U921 ( .A1(n1281), .A2(n1126), .A3(n1119), .ZN(n1213) );
INV_X1 U922 ( .A(n1111), .ZN(n1126) );
NOR2_X1 U923 ( .A1(n1164), .A2(G952), .ZN(n1195) );
NAND2_X1 U924 ( .A1(n1287), .A2(n1288), .ZN(G48) );
NAND2_X1 U925 ( .A1(n1289), .A2(n1260), .ZN(n1288) );
XOR2_X1 U926 ( .A(KEYINPUT31), .B(n1290), .Z(n1287) );
NOR2_X1 U927 ( .A1(n1260), .A2(n1289), .ZN(n1290) );
XNOR2_X1 U928 ( .A(KEYINPUT13), .B(G146), .ZN(n1289) );
AND3_X1 U929 ( .A1(n1119), .A2(n1138), .A3(n1291), .ZN(n1260) );
XNOR2_X1 U930 ( .A(G143), .B(n1267), .ZN(G45) );
NAND2_X1 U931 ( .A1(n1266), .A2(n1292), .ZN(n1267) );
NOR4_X1 U932 ( .A1(n1278), .A2(n1282), .A3(n1135), .A4(n1114), .ZN(n1266) );
NAND2_X1 U933 ( .A1(n1293), .A2(n1294), .ZN(G42) );
OR2_X1 U934 ( .A1(n1253), .A2(G140), .ZN(n1294) );
XOR2_X1 U935 ( .A(n1295), .B(KEYINPUT41), .Z(n1293) );
NAND2_X1 U936 ( .A1(G140), .A2(n1253), .ZN(n1295) );
NAND3_X1 U937 ( .A1(n1119), .A2(n1124), .A3(n1296), .ZN(n1253) );
XNOR2_X1 U938 ( .A(G137), .B(n1254), .ZN(G39) );
NAND4_X1 U939 ( .A1(n1296), .A2(n1137), .A3(n1297), .A4(n1298), .ZN(n1254) );
XOR2_X1 U940 ( .A(n1299), .B(n1259), .Z(G36) );
AND3_X1 U941 ( .A1(n1125), .A2(n1118), .A3(n1296), .ZN(n1259) );
XNOR2_X1 U942 ( .A(G134), .B(KEYINPUT37), .ZN(n1299) );
XOR2_X1 U943 ( .A(G131), .B(n1258), .Z(G33) );
AND3_X1 U944 ( .A1(n1119), .A2(n1125), .A3(n1296), .ZN(n1258) );
NOR3_X1 U945 ( .A1(n1135), .A2(n1264), .A3(n1130), .ZN(n1296) );
OR2_X1 U946 ( .A1(n1122), .A2(n1123), .ZN(n1130) );
INV_X1 U947 ( .A(n1127), .ZN(n1123) );
NAND2_X1 U948 ( .A1(n1300), .A2(n1301), .ZN(G30) );
NAND2_X1 U949 ( .A1(n1257), .A2(n1302), .ZN(n1301) );
XOR2_X1 U950 ( .A(n1303), .B(KEYINPUT17), .Z(n1300) );
OR2_X1 U951 ( .A1(n1302), .A2(n1257), .ZN(n1303) );
AND3_X1 U952 ( .A1(n1118), .A2(n1304), .A3(n1291), .ZN(n1257) );
NOR4_X1 U953 ( .A1(n1114), .A2(n1305), .A3(n1140), .A4(n1264), .ZN(n1291) );
INV_X1 U954 ( .A(n1292), .ZN(n1264) );
XOR2_X1 U955 ( .A(G128), .B(KEYINPUT53), .Z(n1302) );
XOR2_X1 U956 ( .A(n1284), .B(n1306), .Z(G3) );
NOR2_X1 U957 ( .A1(G101), .A2(KEYINPUT59), .ZN(n1306) );
NAND2_X1 U958 ( .A1(n1125), .A2(n1283), .ZN(n1284) );
INV_X1 U959 ( .A(n1282), .ZN(n1125) );
XOR2_X1 U960 ( .A(G125), .B(n1307), .Z(G27) );
NOR2_X1 U961 ( .A1(n1265), .A2(n1308), .ZN(n1307) );
XNOR2_X1 U962 ( .A(KEYINPUT46), .B(n1292), .ZN(n1308) );
NAND2_X1 U963 ( .A1(n1102), .A2(n1309), .ZN(n1292) );
NAND4_X1 U964 ( .A1(G953), .A2(G902), .A3(n1310), .A4(n1311), .ZN(n1309) );
INV_X1 U965 ( .A(G900), .ZN(n1311) );
NAND4_X1 U966 ( .A1(n1119), .A2(n1312), .A3(n1313), .A4(n1124), .ZN(n1265) );
NOR2_X1 U967 ( .A1(n1106), .A2(n1114), .ZN(n1313) );
INV_X1 U968 ( .A(n1314), .ZN(n1119) );
XOR2_X1 U969 ( .A(G122), .B(n1315), .Z(G24) );
NOR3_X1 U970 ( .A1(n1316), .A2(n1111), .A3(n1275), .ZN(n1315) );
NAND2_X1 U971 ( .A1(n1305), .A2(n1317), .ZN(n1111) );
XNOR2_X1 U972 ( .A(KEYINPUT32), .B(n1278), .ZN(n1316) );
NAND2_X1 U973 ( .A1(n1157), .A2(n1318), .ZN(n1278) );
XNOR2_X1 U974 ( .A(n1268), .B(n1319), .ZN(G21) );
XNOR2_X1 U975 ( .A(KEYINPUT44), .B(n1320), .ZN(n1319) );
OR4_X1 U976 ( .A1(n1275), .A2(n1115), .A3(n1305), .A4(n1140), .ZN(n1268) );
INV_X1 U977 ( .A(n1297), .ZN(n1305) );
INV_X1 U978 ( .A(n1137), .ZN(n1115) );
XOR2_X1 U979 ( .A(G116), .B(n1321), .Z(G18) );
NOR3_X1 U980 ( .A1(n1282), .A2(n1280), .A3(n1275), .ZN(n1321) );
INV_X1 U981 ( .A(n1118), .ZN(n1280) );
NOR2_X1 U982 ( .A1(n1318), .A2(n1322), .ZN(n1118) );
XOR2_X1 U983 ( .A(G113), .B(n1286), .Z(G15) );
NOR3_X1 U984 ( .A1(n1282), .A2(n1275), .A3(n1314), .ZN(n1286) );
NAND2_X1 U985 ( .A1(n1322), .A2(n1318), .ZN(n1314) );
INV_X1 U986 ( .A(n1157), .ZN(n1322) );
NAND3_X1 U987 ( .A1(n1323), .A2(n1134), .A3(n1312), .ZN(n1275) );
NAND2_X1 U988 ( .A1(n1297), .A2(n1317), .ZN(n1282) );
XNOR2_X1 U989 ( .A(n1140), .B(KEYINPUT16), .ZN(n1317) );
XOR2_X1 U990 ( .A(G110), .B(n1285), .Z(G12) );
AND2_X1 U991 ( .A1(n1124), .A2(n1283), .ZN(n1285) );
AND2_X1 U992 ( .A1(n1137), .A2(n1281), .ZN(n1283) );
AND2_X1 U993 ( .A1(n1323), .A2(n1304), .ZN(n1281) );
XNOR2_X1 U994 ( .A(n1135), .B(KEYINPUT45), .ZN(n1304) );
INV_X1 U995 ( .A(n1138), .ZN(n1135) );
NOR2_X1 U996 ( .A1(n1312), .A2(n1106), .ZN(n1138) );
INV_X1 U997 ( .A(n1134), .ZN(n1106) );
NAND2_X1 U998 ( .A1(G221), .A2(n1324), .ZN(n1134) );
INV_X1 U999 ( .A(n1105), .ZN(n1312) );
NAND2_X1 U1000 ( .A1(n1149), .A2(n1325), .ZN(n1105) );
NAND2_X1 U1001 ( .A1(G469), .A2(n1326), .ZN(n1325) );
NAND2_X1 U1002 ( .A1(n1147), .A2(n1148), .ZN(n1326) );
NAND3_X1 U1003 ( .A1(n1228), .A2(n1147), .A3(n1148), .ZN(n1149) );
NAND3_X1 U1004 ( .A1(n1327), .A2(n1328), .A3(n1236), .ZN(n1148) );
NAND2_X1 U1005 ( .A1(n1239), .A2(n1238), .ZN(n1236) );
NOR2_X1 U1006 ( .A1(n1329), .A2(n1330), .ZN(n1239) );
NAND2_X1 U1007 ( .A1(n1331), .A2(n1329), .ZN(n1328) );
XNOR2_X1 U1008 ( .A(n1238), .B(n1330), .ZN(n1331) );
NAND3_X1 U1009 ( .A1(n1330), .A2(n1332), .A3(n1333), .ZN(n1327) );
INV_X1 U1010 ( .A(n1238), .ZN(n1332) );
XNOR2_X1 U1011 ( .A(n1334), .B(n1335), .ZN(n1238) );
XOR2_X1 U1012 ( .A(G140), .B(G110), .Z(n1335) );
NAND2_X1 U1013 ( .A1(G227), .A2(n1336), .ZN(n1334) );
XNOR2_X1 U1014 ( .A(KEYINPUT10), .B(n1164), .ZN(n1336) );
XOR2_X1 U1015 ( .A(n1337), .B(n1338), .Z(n1330) );
XNOR2_X1 U1016 ( .A(n1177), .B(n1339), .ZN(n1337) );
XOR2_X1 U1017 ( .A(n1340), .B(n1341), .Z(n1177) );
NAND2_X1 U1018 ( .A1(KEYINPUT58), .A2(n1342), .ZN(n1340) );
INV_X1 U1019 ( .A(G469), .ZN(n1228) );
NOR2_X1 U1020 ( .A1(n1114), .A2(n1343), .ZN(n1323) );
AND2_X1 U1021 ( .A1(n1344), .A2(n1102), .ZN(n1343) );
NAND3_X1 U1022 ( .A1(n1310), .A2(n1164), .A3(G952), .ZN(n1102) );
NAND4_X1 U1023 ( .A1(G953), .A2(G902), .A3(n1187), .A4(n1310), .ZN(n1344) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1310) );
XOR2_X1 U1025 ( .A(KEYINPUT61), .B(G898), .Z(n1187) );
NAND2_X1 U1026 ( .A1(n1127), .A2(n1122), .ZN(n1114) );
NAND2_X1 U1027 ( .A1(n1161), .A2(n1150), .ZN(n1122) );
NAND2_X1 U1028 ( .A1(G210), .A2(n1345), .ZN(n1150) );
NAND2_X1 U1029 ( .A1(n1147), .A2(n1346), .ZN(n1345) );
NAND2_X1 U1030 ( .A1(G237), .A2(n1347), .ZN(n1346) );
NAND3_X1 U1031 ( .A1(n1348), .A2(n1147), .A3(n1349), .ZN(n1161) );
INV_X1 U1032 ( .A(n1347), .ZN(n1349) );
XNOR2_X1 U1033 ( .A(n1350), .B(n1351), .ZN(n1347) );
XNOR2_X1 U1034 ( .A(n1352), .B(n1248), .ZN(n1351) );
XOR2_X1 U1035 ( .A(n1190), .B(n1353), .Z(n1248) );
NOR2_X1 U1036 ( .A1(KEYINPUT6), .A2(n1189), .ZN(n1353) );
XNOR2_X1 U1037 ( .A(n1354), .B(n1355), .ZN(n1189) );
NOR2_X1 U1038 ( .A1(n1356), .A2(n1357), .ZN(n1355) );
XOR2_X1 U1039 ( .A(n1358), .B(KEYINPUT23), .Z(n1357) );
NAND2_X1 U1040 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
NOR2_X1 U1041 ( .A1(n1359), .A2(n1360), .ZN(n1356) );
NAND3_X1 U1042 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1360) );
OR2_X1 U1043 ( .A1(n1364), .A2(KEYINPUT62), .ZN(n1363) );
NAND3_X1 U1044 ( .A1(KEYINPUT62), .A2(n1364), .A3(G119), .ZN(n1362) );
NAND2_X1 U1045 ( .A1(n1365), .A2(n1320), .ZN(n1361) );
NAND2_X1 U1046 ( .A1(n1366), .A2(KEYINPUT62), .ZN(n1365) );
XNOR2_X1 U1047 ( .A(n1364), .B(KEYINPUT36), .ZN(n1366) );
NAND2_X1 U1048 ( .A1(n1367), .A2(n1368), .ZN(n1354) );
NAND2_X1 U1049 ( .A1(n1369), .A2(n1339), .ZN(n1368) );
XOR2_X1 U1050 ( .A(KEYINPUT15), .B(n1338), .Z(n1369) );
NAND2_X1 U1051 ( .A1(n1338), .A2(G107), .ZN(n1367) );
XOR2_X1 U1052 ( .A(G101), .B(G104), .Z(n1338) );
XOR2_X1 U1053 ( .A(G110), .B(n1370), .Z(n1190) );
NAND2_X1 U1054 ( .A1(G224), .A2(n1164), .ZN(n1352) );
XNOR2_X1 U1055 ( .A(G125), .B(n1371), .ZN(n1350) );
NOR2_X1 U1056 ( .A1(KEYINPUT38), .A2(n1372), .ZN(n1371) );
NAND2_X1 U1057 ( .A1(G210), .A2(G237), .ZN(n1348) );
NAND2_X1 U1058 ( .A1(G214), .A2(n1373), .ZN(n1127) );
OR2_X1 U1059 ( .A1(G237), .A2(G902), .ZN(n1373) );
NOR2_X1 U1060 ( .A1(n1157), .A2(n1318), .ZN(n1137) );
NAND2_X1 U1061 ( .A1(n1374), .A2(n1375), .ZN(n1318) );
NAND2_X1 U1062 ( .A1(n1154), .A2(n1156), .ZN(n1375) );
INV_X1 U1063 ( .A(G475), .ZN(n1156) );
XOR2_X1 U1064 ( .A(n1376), .B(KEYINPUT43), .Z(n1374) );
NAND2_X1 U1065 ( .A1(G475), .A2(n1377), .ZN(n1376) );
INV_X1 U1066 ( .A(n1154), .ZN(n1377) );
NOR2_X1 U1067 ( .A1(n1210), .A2(G902), .ZN(n1154) );
XNOR2_X1 U1068 ( .A(n1378), .B(n1379), .ZN(n1210) );
XOR2_X1 U1069 ( .A(n1370), .B(n1380), .Z(n1379) );
XNOR2_X1 U1070 ( .A(n1174), .B(n1359), .ZN(n1380) );
XOR2_X1 U1071 ( .A(n1381), .B(n1382), .Z(n1378) );
XNOR2_X1 U1072 ( .A(G104), .B(n1383), .ZN(n1382) );
NAND2_X1 U1073 ( .A1(KEYINPUT52), .A2(n1384), .ZN(n1383) );
XOR2_X1 U1074 ( .A(n1385), .B(n1386), .Z(n1384) );
XNOR2_X1 U1075 ( .A(G143), .B(n1387), .ZN(n1386) );
NAND2_X1 U1076 ( .A1(G214), .A2(n1388), .ZN(n1387) );
NOR2_X1 U1077 ( .A1(G131), .A2(KEYINPUT60), .ZN(n1385) );
NAND2_X1 U1078 ( .A1(KEYINPUT8), .A2(n1389), .ZN(n1381) );
XOR2_X1 U1079 ( .A(n1390), .B(n1204), .Z(n1157) );
INV_X1 U1080 ( .A(G478), .ZN(n1204) );
NAND2_X1 U1081 ( .A1(n1391), .A2(n1147), .ZN(n1390) );
XNOR2_X1 U1082 ( .A(n1203), .B(KEYINPUT3), .ZN(n1391) );
XNOR2_X1 U1083 ( .A(n1392), .B(n1393), .ZN(n1203) );
XOR2_X1 U1084 ( .A(n1394), .B(n1395), .Z(n1393) );
XOR2_X1 U1085 ( .A(G128), .B(G116), .Z(n1395) );
XNOR2_X1 U1086 ( .A(n1396), .B(G134), .ZN(n1394) );
INV_X1 U1087 ( .A(G143), .ZN(n1396) );
XOR2_X1 U1088 ( .A(n1397), .B(n1370), .Z(n1392) );
XOR2_X1 U1089 ( .A(G122), .B(KEYINPUT57), .Z(n1370) );
XNOR2_X1 U1090 ( .A(n1398), .B(n1339), .ZN(n1397) );
INV_X1 U1091 ( .A(G107), .ZN(n1339) );
NAND2_X1 U1092 ( .A1(G217), .A2(n1399), .ZN(n1398) );
NOR2_X1 U1093 ( .A1(n1297), .A2(n1140), .ZN(n1124) );
INV_X1 U1094 ( .A(n1298), .ZN(n1140) );
XOR2_X1 U1095 ( .A(n1400), .B(n1199), .Z(n1298) );
NAND2_X1 U1096 ( .A1(G217), .A2(n1324), .ZN(n1199) );
NAND2_X1 U1097 ( .A1(G234), .A2(n1147), .ZN(n1324) );
OR2_X1 U1098 ( .A1(n1198), .A2(G902), .ZN(n1400) );
XNOR2_X1 U1099 ( .A(n1401), .B(n1402), .ZN(n1198) );
XNOR2_X1 U1100 ( .A(G137), .B(n1403), .ZN(n1402) );
NAND2_X1 U1101 ( .A1(n1404), .A2(n1405), .ZN(n1403) );
NAND2_X1 U1102 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
XOR2_X1 U1103 ( .A(n1408), .B(KEYINPUT4), .Z(n1404) );
OR2_X1 U1104 ( .A1(n1407), .A2(n1406), .ZN(n1408) );
XNOR2_X1 U1105 ( .A(G110), .B(n1409), .ZN(n1406) );
XNOR2_X1 U1106 ( .A(G128), .B(n1320), .ZN(n1409) );
INV_X1 U1107 ( .A(G119), .ZN(n1320) );
XNOR2_X1 U1108 ( .A(G146), .B(n1174), .ZN(n1407) );
XNOR2_X1 U1109 ( .A(G125), .B(G140), .ZN(n1174) );
NAND2_X1 U1110 ( .A1(G221), .A2(n1399), .ZN(n1401) );
AND2_X1 U1111 ( .A1(G234), .A2(n1164), .ZN(n1399) );
INV_X1 U1112 ( .A(G953), .ZN(n1164) );
XOR2_X1 U1113 ( .A(n1160), .B(n1222), .Z(n1297) );
INV_X1 U1114 ( .A(G472), .ZN(n1222) );
NAND2_X1 U1115 ( .A1(n1410), .A2(n1147), .ZN(n1160) );
INV_X1 U1116 ( .A(G902), .ZN(n1147) );
XNOR2_X1 U1117 ( .A(n1223), .B(n1411), .ZN(n1410) );
XNOR2_X1 U1118 ( .A(n1412), .B(n1216), .ZN(n1411) );
XNOR2_X1 U1119 ( .A(n1413), .B(G101), .ZN(n1216) );
NAND2_X1 U1120 ( .A1(G210), .A2(n1388), .ZN(n1413) );
NOR2_X1 U1121 ( .A1(G953), .A2(G237), .ZN(n1388) );
NAND3_X1 U1122 ( .A1(n1414), .A2(n1415), .A3(KEYINPUT55), .ZN(n1412) );
NAND3_X1 U1123 ( .A1(n1329), .A2(n1372), .A3(n1416), .ZN(n1415) );
OR2_X1 U1124 ( .A1(n1219), .A2(n1416), .ZN(n1414) );
INV_X1 U1125 ( .A(KEYINPUT51), .ZN(n1416) );
XNOR2_X1 U1126 ( .A(n1329), .B(n1372), .ZN(n1219) );
INV_X1 U1127 ( .A(n1249), .ZN(n1372) );
XOR2_X1 U1128 ( .A(n1342), .B(n1341), .Z(n1249) );
XNOR2_X1 U1129 ( .A(G128), .B(n1389), .ZN(n1341) );
INV_X1 U1130 ( .A(G146), .ZN(n1389) );
XOR2_X1 U1131 ( .A(G143), .B(KEYINPUT1), .Z(n1342) );
INV_X1 U1132 ( .A(n1333), .ZN(n1329) );
NAND2_X1 U1133 ( .A1(n1417), .A2(n1418), .ZN(n1333) );
NAND2_X1 U1134 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
INV_X1 U1135 ( .A(G137), .ZN(n1420) );
XOR2_X1 U1136 ( .A(KEYINPUT35), .B(n1179), .Z(n1419) );
NAND2_X1 U1137 ( .A1(n1179), .A2(G137), .ZN(n1417) );
XOR2_X1 U1138 ( .A(G131), .B(G134), .Z(n1179) );
XOR2_X1 U1139 ( .A(n1421), .B(n1422), .Z(n1223) );
XOR2_X1 U1140 ( .A(n1359), .B(n1364), .Z(n1422) );
XOR2_X1 U1141 ( .A(G116), .B(KEYINPUT54), .Z(n1364) );
XOR2_X1 U1142 ( .A(G113), .B(KEYINPUT21), .Z(n1359) );
XNOR2_X1 U1143 ( .A(KEYINPUT29), .B(n1423), .ZN(n1421) );
NOR2_X1 U1144 ( .A1(G119), .A2(KEYINPUT26), .ZN(n1423) );
endmodule


