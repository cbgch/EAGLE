//Key = 0110010100001000111000101011111101011011110101010100001001000000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350;

XNOR2_X1 U731 ( .A(G107), .B(n1029), .ZN(G9) );
NAND4_X1 U732 ( .A1(n1030), .A2(n1031), .A3(n1032), .A4(n1033), .ZN(n1029) );
XNOR2_X1 U733 ( .A(n1034), .B(KEYINPUT45), .ZN(n1030) );
NOR2_X1 U734 ( .A1(n1035), .A2(n1036), .ZN(G75) );
XOR2_X1 U735 ( .A(KEYINPUT9), .B(n1037), .Z(n1036) );
AND3_X1 U736 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NOR4_X1 U737 ( .A1(n1041), .A2(n1042), .A3(n1039), .A4(n1043), .ZN(n1035) );
INV_X1 U738 ( .A(G952), .ZN(n1039) );
NAND4_X1 U739 ( .A1(n1038), .A2(n1044), .A3(n1045), .A4(n1040), .ZN(n1041) );
NAND4_X1 U740 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1040) );
NOR4_X1 U741 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1049) );
XOR2_X1 U742 ( .A(n1054), .B(n1055), .Z(n1051) );
NOR2_X1 U743 ( .A1(n1056), .A2(KEYINPUT32), .ZN(n1055) );
INV_X1 U744 ( .A(n1057), .ZN(n1056) );
NOR2_X1 U745 ( .A1(n1058), .A2(n1059), .ZN(n1048) );
AND3_X1 U746 ( .A1(n1060), .A2(n1061), .A3(KEYINPUT49), .ZN(n1059) );
NOR2_X1 U747 ( .A1(n1062), .A2(n1060), .ZN(n1058) );
NOR2_X1 U748 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
NOR2_X1 U749 ( .A1(KEYINPUT49), .A2(n1065), .ZN(n1063) );
INV_X1 U750 ( .A(n1061), .ZN(n1065) );
XNOR2_X1 U751 ( .A(n1064), .B(KEYINPUT44), .ZN(n1061) );
XNOR2_X1 U752 ( .A(n1066), .B(G475), .ZN(n1046) );
NAND3_X1 U753 ( .A1(n1047), .A2(n1067), .A3(n1068), .ZN(n1045) );
NAND2_X1 U754 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
NAND2_X1 U755 ( .A1(n1032), .A2(n1071), .ZN(n1070) );
NAND2_X1 U756 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND2_X1 U757 ( .A1(n1074), .A2(n1033), .ZN(n1073) );
XNOR2_X1 U758 ( .A(n1075), .B(KEYINPUT1), .ZN(n1074) );
NAND2_X1 U759 ( .A1(n1075), .A2(n1076), .ZN(n1072) );
NAND2_X1 U760 ( .A1(n1077), .A2(n1078), .ZN(n1069) );
NAND2_X1 U761 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U762 ( .A1(n1032), .A2(n1081), .ZN(n1080) );
NAND2_X1 U763 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U764 ( .A1(n1050), .A2(n1084), .ZN(n1083) );
NAND2_X1 U765 ( .A1(n1075), .A2(n1085), .ZN(n1079) );
NAND2_X1 U766 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U767 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XNOR2_X1 U768 ( .A(n1090), .B(KEYINPUT34), .ZN(n1086) );
NAND2_X1 U769 ( .A1(n1075), .A2(n1091), .ZN(n1044) );
NAND2_X1 U770 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND2_X1 U771 ( .A1(n1094), .A2(n1034), .ZN(n1093) );
XOR2_X1 U772 ( .A(n1095), .B(KEYINPUT62), .Z(n1092) );
NAND3_X1 U773 ( .A1(n1096), .A2(n1094), .A3(n1097), .ZN(n1095) );
AND3_X1 U774 ( .A1(n1077), .A2(n1032), .A3(n1068), .ZN(n1094) );
INV_X1 U775 ( .A(n1098), .ZN(n1068) );
XOR2_X1 U776 ( .A(n1099), .B(n1100), .Z(G72) );
NOR2_X1 U777 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
NOR2_X1 U778 ( .A1(n1103), .A2(n1104), .ZN(n1101) );
NAND2_X1 U779 ( .A1(n1105), .A2(n1106), .ZN(n1099) );
NAND3_X1 U780 ( .A1(n1107), .A2(n1108), .A3(n1043), .ZN(n1106) );
NAND2_X1 U781 ( .A1(G953), .A2(n1109), .ZN(n1108) );
NAND2_X1 U782 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U783 ( .A1(G900), .A2(n1112), .ZN(n1110) );
NAND2_X1 U784 ( .A1(n1113), .A2(n1114), .ZN(n1107) );
OR2_X1 U785 ( .A1(n1111), .A2(n1112), .ZN(n1113) );
INV_X1 U786 ( .A(KEYINPUT24), .ZN(n1111) );
NAND2_X1 U787 ( .A1(n1112), .A2(n1115), .ZN(n1105) );
NAND2_X1 U788 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U789 ( .A1(G900), .A2(n1118), .ZN(n1117) );
NAND2_X1 U790 ( .A1(n1043), .A2(n1119), .ZN(n1118) );
NAND2_X1 U791 ( .A1(KEYINPUT24), .A2(G953), .ZN(n1119) );
NAND2_X1 U792 ( .A1(n1120), .A2(n1114), .ZN(n1116) );
NAND2_X1 U793 ( .A1(KEYINPUT24), .A2(n1043), .ZN(n1120) );
XOR2_X1 U794 ( .A(n1121), .B(n1122), .Z(n1112) );
XOR2_X1 U795 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U796 ( .A(n1125), .B(n1126), .Z(n1121) );
NAND2_X1 U797 ( .A1(n1127), .A2(n1128), .ZN(n1125) );
XOR2_X1 U798 ( .A(KEYINPUT36), .B(n1129), .Z(n1127) );
XOR2_X1 U799 ( .A(n1130), .B(n1131), .Z(G69) );
NOR2_X1 U800 ( .A1(n1132), .A2(n1102), .ZN(n1131) );
XNOR2_X1 U801 ( .A(G953), .B(KEYINPUT46), .ZN(n1102) );
NOR2_X1 U802 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U803 ( .A1(n1135), .A2(n1136), .ZN(n1130) );
NAND2_X1 U804 ( .A1(n1137), .A2(n1114), .ZN(n1136) );
XOR2_X1 U805 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U806 ( .A(n1042), .B(KEYINPUT6), .Z(n1138) );
NAND3_X1 U807 ( .A1(n1139), .A2(G898), .A3(G953), .ZN(n1135) );
NOR2_X1 U808 ( .A1(KEYINPUT59), .A2(n1140), .ZN(n1139) );
NOR2_X1 U809 ( .A1(n1141), .A2(n1142), .ZN(G66) );
XOR2_X1 U810 ( .A(KEYINPUT51), .B(n1143), .Z(n1142) );
XNOR2_X1 U811 ( .A(n1144), .B(n1145), .ZN(n1141) );
NOR2_X1 U812 ( .A1(n1064), .A2(n1146), .ZN(n1145) );
NOR2_X1 U813 ( .A1(n1143), .A2(n1147), .ZN(G63) );
XOR2_X1 U814 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U815 ( .A1(n1150), .A2(n1146), .ZN(n1148) );
INV_X1 U816 ( .A(G478), .ZN(n1150) );
NOR2_X1 U817 ( .A1(n1143), .A2(n1151), .ZN(G60) );
NOR3_X1 U818 ( .A1(n1152), .A2(n1153), .A3(n1154), .ZN(n1151) );
AND2_X1 U819 ( .A1(n1155), .A2(KEYINPUT3), .ZN(n1154) );
NOR2_X1 U820 ( .A1(KEYINPUT3), .A2(n1156), .ZN(n1153) );
NOR2_X1 U821 ( .A1(n1157), .A2(n1066), .ZN(n1156) );
NOR2_X1 U822 ( .A1(n1158), .A2(n1155), .ZN(n1157) );
NOR2_X1 U823 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
NOR2_X1 U824 ( .A1(n1043), .A2(n1042), .ZN(n1159) );
NOR3_X1 U825 ( .A1(n1146), .A2(n1161), .A3(n1160), .ZN(n1152) );
INV_X1 U826 ( .A(G475), .ZN(n1160) );
NOR2_X1 U827 ( .A1(KEYINPUT3), .A2(n1155), .ZN(n1161) );
XNOR2_X1 U828 ( .A(G104), .B(n1162), .ZN(G6) );
NOR2_X1 U829 ( .A1(n1143), .A2(n1163), .ZN(G57) );
XOR2_X1 U830 ( .A(n1164), .B(n1165), .Z(n1163) );
XNOR2_X1 U831 ( .A(KEYINPUT43), .B(n1166), .ZN(n1165) );
NOR2_X1 U832 ( .A1(n1167), .A2(KEYINPUT52), .ZN(n1166) );
NOR2_X1 U833 ( .A1(n1168), .A2(n1146), .ZN(n1167) );
NOR2_X1 U834 ( .A1(n1143), .A2(n1169), .ZN(G54) );
XOR2_X1 U835 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U836 ( .A(n1172), .B(n1173), .ZN(n1171) );
XOR2_X1 U837 ( .A(n1174), .B(n1175), .Z(n1170) );
NOR2_X1 U838 ( .A1(KEYINPUT58), .A2(n1176), .ZN(n1175) );
NOR2_X1 U839 ( .A1(n1177), .A2(n1146), .ZN(n1176) );
XNOR2_X1 U840 ( .A(KEYINPUT61), .B(KEYINPUT2), .ZN(n1174) );
NOR2_X1 U841 ( .A1(n1143), .A2(n1178), .ZN(G51) );
XOR2_X1 U842 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U843 ( .A(n1181), .B(n1182), .Z(n1180) );
NOR2_X1 U844 ( .A1(n1057), .A2(n1146), .ZN(n1182) );
NAND2_X1 U845 ( .A1(G902), .A2(n1183), .ZN(n1146) );
OR2_X1 U846 ( .A1(n1042), .A2(n1043), .ZN(n1183) );
NAND4_X1 U847 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1043) );
NOR4_X1 U848 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NOR2_X1 U849 ( .A1(n1082), .A2(n1192), .ZN(n1191) );
NOR2_X1 U850 ( .A1(n1193), .A2(n1194), .ZN(n1190) );
INV_X1 U851 ( .A(KEYINPUT40), .ZN(n1194) );
AND3_X1 U852 ( .A1(KEYINPUT31), .A2(n1033), .A3(n1195), .ZN(n1189) );
NOR3_X1 U853 ( .A1(n1196), .A2(n1034), .A3(n1197), .ZN(n1188) );
NOR2_X1 U854 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
NOR4_X1 U855 ( .A1(KEYINPUT31), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1199) );
NOR4_X1 U856 ( .A1(KEYINPUT40), .A2(n1082), .A3(n1203), .A4(n1204), .ZN(n1198) );
AND3_X1 U857 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1186) );
NAND4_X1 U858 ( .A1(n1208), .A2(n1162), .A3(n1209), .A4(n1210), .ZN(n1042) );
NOR4_X1 U859 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
NOR3_X1 U860 ( .A1(n1204), .A2(n1215), .A3(n1216), .ZN(n1214) );
NOR4_X1 U861 ( .A1(n1217), .A2(n1200), .A3(n1218), .A4(n1219), .ZN(n1213) );
XOR2_X1 U862 ( .A(KEYINPUT28), .B(n1032), .Z(n1219) );
NOR2_X1 U863 ( .A1(n1220), .A2(n1221), .ZN(n1209) );
NAND4_X1 U864 ( .A1(n1076), .A2(n1031), .A3(n1032), .A4(n1034), .ZN(n1162) );
INV_X1 U865 ( .A(n1218), .ZN(n1031) );
NOR2_X1 U866 ( .A1(KEYINPUT42), .A2(n1222), .ZN(n1181) );
XNOR2_X1 U867 ( .A(n1223), .B(n1224), .ZN(n1222) );
XOR2_X1 U868 ( .A(KEYINPUT33), .B(n1225), .Z(n1224) );
NOR2_X1 U869 ( .A1(n1114), .A2(G952), .ZN(n1143) );
XNOR2_X1 U870 ( .A(G146), .B(n1193), .ZN(G48) );
NAND3_X1 U871 ( .A1(n1076), .A2(n1226), .A3(n1227), .ZN(n1193) );
XNOR2_X1 U872 ( .A(n1228), .B(n1229), .ZN(G45) );
NOR2_X1 U873 ( .A1(n1230), .A2(n1082), .ZN(n1229) );
XOR2_X1 U874 ( .A(n1192), .B(KEYINPUT55), .Z(n1230) );
NAND2_X1 U875 ( .A1(n1231), .A2(n1232), .ZN(n1192) );
XNOR2_X1 U876 ( .A(G140), .B(n1184), .ZN(G42) );
NAND3_X1 U877 ( .A1(n1075), .A2(n1034), .A3(n1233), .ZN(n1184) );
XNOR2_X1 U878 ( .A(G137), .B(n1185), .ZN(G39) );
NAND3_X1 U879 ( .A1(n1075), .A2(n1077), .A3(n1227), .ZN(n1185) );
XNOR2_X1 U880 ( .A(G134), .B(n1234), .ZN(G36) );
NAND2_X1 U881 ( .A1(n1195), .A2(n1033), .ZN(n1234) );
XOR2_X1 U882 ( .A(n1206), .B(n1235), .Z(G33) );
XOR2_X1 U883 ( .A(KEYINPUT38), .B(G131), .Z(n1235) );
NAND2_X1 U884 ( .A1(n1195), .A2(n1076), .ZN(n1206) );
AND2_X1 U885 ( .A1(n1075), .A2(n1231), .ZN(n1195) );
NOR3_X1 U886 ( .A1(n1217), .A2(n1197), .A3(n1201), .ZN(n1231) );
INV_X1 U887 ( .A(n1202), .ZN(n1075) );
NAND2_X1 U888 ( .A1(n1084), .A2(n1236), .ZN(n1202) );
NAND2_X1 U889 ( .A1(n1237), .A2(n1238), .ZN(G30) );
NAND2_X1 U890 ( .A1(n1239), .A2(n1205), .ZN(n1238) );
XNOR2_X1 U891 ( .A(G128), .B(KEYINPUT7), .ZN(n1239) );
XOR2_X1 U892 ( .A(KEYINPUT18), .B(n1240), .Z(n1237) );
NOR2_X1 U893 ( .A1(n1241), .A2(n1205), .ZN(n1240) );
NAND3_X1 U894 ( .A1(n1033), .A2(n1226), .A3(n1227), .ZN(n1205) );
NOR3_X1 U895 ( .A1(n1217), .A2(n1197), .A3(n1204), .ZN(n1227) );
INV_X1 U896 ( .A(n1242), .ZN(n1197) );
XNOR2_X1 U897 ( .A(G128), .B(KEYINPUT54), .ZN(n1241) );
XNOR2_X1 U898 ( .A(n1243), .B(n1212), .ZN(G3) );
AND2_X1 U899 ( .A1(n1090), .A2(n1244), .ZN(n1212) );
XNOR2_X1 U900 ( .A(G125), .B(n1207), .ZN(G27) );
NAND3_X1 U901 ( .A1(n1047), .A2(n1226), .A3(n1233), .ZN(n1207) );
AND4_X1 U902 ( .A1(n1088), .A2(n1076), .A3(n1089), .A4(n1242), .ZN(n1233) );
NAND2_X1 U903 ( .A1(n1098), .A2(n1245), .ZN(n1242) );
NAND4_X1 U904 ( .A1(G953), .A2(G902), .A3(n1246), .A4(n1104), .ZN(n1245) );
INV_X1 U905 ( .A(G900), .ZN(n1104) );
INV_X1 U906 ( .A(n1247), .ZN(n1047) );
XOR2_X1 U907 ( .A(G122), .B(n1211), .Z(G24) );
AND3_X1 U908 ( .A1(n1248), .A2(n1032), .A3(n1232), .ZN(n1211) );
AND2_X1 U909 ( .A1(n1249), .A2(n1052), .ZN(n1232) );
XNOR2_X1 U910 ( .A(n1250), .B(KEYINPUT56), .ZN(n1249) );
NOR2_X1 U911 ( .A1(n1053), .A2(n1089), .ZN(n1032) );
XOR2_X1 U912 ( .A(n1251), .B(n1252), .Z(G21) );
NOR2_X1 U913 ( .A1(G119), .A2(KEYINPUT48), .ZN(n1252) );
NAND4_X1 U914 ( .A1(n1253), .A2(n1254), .A3(n1077), .A4(n1255), .ZN(n1251) );
NOR2_X1 U915 ( .A1(n1247), .A2(n1204), .ZN(n1255) );
NAND2_X1 U916 ( .A1(n1089), .A2(n1053), .ZN(n1204) );
XNOR2_X1 U917 ( .A(KEYINPUT25), .B(n1082), .ZN(n1253) );
INV_X1 U918 ( .A(n1226), .ZN(n1082) );
XOR2_X1 U919 ( .A(n1221), .B(n1256), .Z(G18) );
NOR2_X1 U920 ( .A1(KEYINPUT23), .A2(n1257), .ZN(n1256) );
NOR3_X1 U921 ( .A1(n1216), .A2(n1200), .A3(n1201), .ZN(n1221) );
INV_X1 U922 ( .A(n1033), .ZN(n1200) );
NOR2_X1 U923 ( .A1(n1258), .A2(n1259), .ZN(n1033) );
INV_X1 U924 ( .A(n1052), .ZN(n1258) );
XOR2_X1 U925 ( .A(G113), .B(n1220), .Z(G15) );
NOR3_X1 U926 ( .A1(n1216), .A2(n1203), .A3(n1201), .ZN(n1220) );
INV_X1 U927 ( .A(n1090), .ZN(n1201) );
NOR2_X1 U928 ( .A1(n1089), .A2(n1088), .ZN(n1090) );
INV_X1 U929 ( .A(n1076), .ZN(n1203) );
NOR2_X1 U930 ( .A1(n1250), .A2(n1052), .ZN(n1076) );
INV_X1 U931 ( .A(n1248), .ZN(n1216) );
NOR2_X1 U932 ( .A1(n1247), .A2(n1218), .ZN(n1248) );
NAND2_X1 U933 ( .A1(n1096), .A2(n1260), .ZN(n1247) );
XNOR2_X1 U934 ( .A(G110), .B(n1208), .ZN(G12) );
NAND3_X1 U935 ( .A1(n1088), .A2(n1089), .A3(n1244), .ZN(n1208) );
NOR3_X1 U936 ( .A1(n1218), .A2(n1217), .A3(n1215), .ZN(n1244) );
INV_X1 U937 ( .A(n1077), .ZN(n1215) );
NOR2_X1 U938 ( .A1(n1052), .A2(n1259), .ZN(n1077) );
INV_X1 U939 ( .A(n1250), .ZN(n1259) );
XOR2_X1 U940 ( .A(n1066), .B(n1261), .Z(n1250) );
NOR2_X1 U941 ( .A1(G475), .A2(KEYINPUT15), .ZN(n1261) );
NOR2_X1 U942 ( .A1(n1155), .A2(G902), .ZN(n1066) );
XOR2_X1 U943 ( .A(n1262), .B(n1263), .Z(n1155) );
XNOR2_X1 U944 ( .A(n1264), .B(n1265), .ZN(n1263) );
XNOR2_X1 U945 ( .A(n1123), .B(n1266), .ZN(n1265) );
NOR2_X1 U946 ( .A1(KEYINPUT4), .A2(n1124), .ZN(n1266) );
XNOR2_X1 U947 ( .A(n1267), .B(G125), .ZN(n1124) );
INV_X1 U948 ( .A(G140), .ZN(n1267) );
XOR2_X1 U949 ( .A(n1268), .B(n1269), .Z(n1262) );
XNOR2_X1 U950 ( .A(n1270), .B(G143), .ZN(n1269) );
XOR2_X1 U951 ( .A(n1271), .B(G104), .Z(n1268) );
NAND2_X1 U952 ( .A1(n1272), .A2(G214), .ZN(n1271) );
XOR2_X1 U953 ( .A(G478), .B(n1273), .Z(n1052) );
NOR2_X1 U954 ( .A1(G902), .A2(n1149), .ZN(n1273) );
XNOR2_X1 U955 ( .A(n1274), .B(n1275), .ZN(n1149) );
XOR2_X1 U956 ( .A(n1276), .B(n1277), .Z(n1275) );
NOR3_X1 U957 ( .A1(n1278), .A2(KEYINPUT0), .A3(n1279), .ZN(n1276) );
INV_X1 U958 ( .A(G217), .ZN(n1278) );
XOR2_X1 U959 ( .A(n1280), .B(n1281), .Z(n1274) );
NOR2_X1 U960 ( .A1(KEYINPUT63), .A2(n1282), .ZN(n1281) );
XOR2_X1 U961 ( .A(G134), .B(n1283), .Z(n1282) );
XNOR2_X1 U962 ( .A(G107), .B(G116), .ZN(n1280) );
INV_X1 U963 ( .A(n1034), .ZN(n1217) );
NOR2_X1 U964 ( .A1(n1096), .A2(n1097), .ZN(n1034) );
INV_X1 U965 ( .A(n1260), .ZN(n1097) );
NAND2_X1 U966 ( .A1(G221), .A2(n1284), .ZN(n1260) );
XNOR2_X1 U967 ( .A(n1285), .B(n1177), .ZN(n1096) );
INV_X1 U968 ( .A(G469), .ZN(n1177) );
NAND2_X1 U969 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
XOR2_X1 U970 ( .A(n1288), .B(n1172), .Z(n1286) );
XNOR2_X1 U971 ( .A(n1289), .B(n1290), .ZN(n1172) );
XNOR2_X1 U972 ( .A(n1243), .B(n1291), .ZN(n1290) );
XOR2_X1 U973 ( .A(G107), .B(G104), .Z(n1291) );
XOR2_X1 U974 ( .A(n1292), .B(n1293), .Z(n1289) );
XOR2_X1 U975 ( .A(n1126), .B(n1294), .Z(n1293) );
NOR2_X1 U976 ( .A1(G953), .A2(n1103), .ZN(n1294) );
INV_X1 U977 ( .A(G227), .ZN(n1103) );
AND2_X1 U978 ( .A1(n1295), .A2(n1296), .ZN(n1126) );
NAND2_X1 U979 ( .A1(n1297), .A2(G128), .ZN(n1296) );
XOR2_X1 U980 ( .A(KEYINPUT26), .B(n1298), .Z(n1295) );
NOR2_X1 U981 ( .A1(G128), .A2(n1299), .ZN(n1298) );
XOR2_X1 U982 ( .A(n1297), .B(KEYINPUT11), .Z(n1299) );
XNOR2_X1 U983 ( .A(n1300), .B(n1270), .ZN(n1297) );
NAND2_X1 U984 ( .A1(KEYINPUT41), .A2(n1228), .ZN(n1300) );
NOR2_X1 U985 ( .A1(KEYINPUT13), .A2(n1173), .ZN(n1288) );
NAND2_X1 U986 ( .A1(n1226), .A2(n1254), .ZN(n1218) );
NAND2_X1 U987 ( .A1(n1301), .A2(n1098), .ZN(n1254) );
NAND3_X1 U988 ( .A1(n1038), .A2(n1246), .A3(G952), .ZN(n1098) );
XOR2_X1 U989 ( .A(n1114), .B(KEYINPUT37), .Z(n1038) );
NAND4_X1 U990 ( .A1(G953), .A2(G902), .A3(n1246), .A4(n1134), .ZN(n1301) );
INV_X1 U991 ( .A(G898), .ZN(n1134) );
NAND2_X1 U992 ( .A1(G237), .A2(n1302), .ZN(n1246) );
XOR2_X1 U993 ( .A(KEYINPUT21), .B(G234), .Z(n1302) );
NOR2_X1 U994 ( .A1(n1084), .A2(n1050), .ZN(n1226) );
INV_X1 U995 ( .A(n1236), .ZN(n1050) );
NAND2_X1 U996 ( .A1(G214), .A2(n1303), .ZN(n1236) );
XOR2_X1 U997 ( .A(n1304), .B(n1057), .Z(n1084) );
NAND2_X1 U998 ( .A1(G210), .A2(n1303), .ZN(n1057) );
NAND2_X1 U999 ( .A1(n1305), .A2(n1287), .ZN(n1303) );
XOR2_X1 U1000 ( .A(KEYINPUT39), .B(G237), .Z(n1305) );
XOR2_X1 U1001 ( .A(n1054), .B(KEYINPUT30), .Z(n1304) );
NAND2_X1 U1002 ( .A1(n1306), .A2(n1287), .ZN(n1054) );
XOR2_X1 U1003 ( .A(n1307), .B(n1308), .Z(n1306) );
XOR2_X1 U1004 ( .A(n1309), .B(n1179), .Z(n1308) );
XNOR2_X1 U1005 ( .A(n1140), .B(KEYINPUT22), .ZN(n1179) );
XNOR2_X1 U1006 ( .A(n1310), .B(n1311), .ZN(n1140) );
XOR2_X1 U1007 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1008 ( .A(G110), .B(G104), .Z(n1313) );
XNOR2_X1 U1009 ( .A(KEYINPUT29), .B(n1257), .ZN(n1312) );
INV_X1 U1010 ( .A(G116), .ZN(n1257) );
XOR2_X1 U1011 ( .A(n1314), .B(n1315), .Z(n1310) );
XNOR2_X1 U1012 ( .A(G101), .B(n1316), .ZN(n1315) );
NAND2_X1 U1013 ( .A1(KEYINPUT47), .A2(G107), .ZN(n1316) );
XNOR2_X1 U1014 ( .A(n1317), .B(n1318), .ZN(n1314) );
INV_X1 U1015 ( .A(n1264), .ZN(n1318) );
XOR2_X1 U1016 ( .A(G113), .B(n1277), .Z(n1264) );
XOR2_X1 U1017 ( .A(G122), .B(KEYINPUT20), .Z(n1277) );
NAND2_X1 U1018 ( .A1(KEYINPUT27), .A2(n1319), .ZN(n1317) );
NAND2_X1 U1019 ( .A1(KEYINPUT57), .A2(n1223), .ZN(n1309) );
XNOR2_X1 U1020 ( .A(n1320), .B(n1321), .ZN(n1223) );
XNOR2_X1 U1021 ( .A(G125), .B(KEYINPUT8), .ZN(n1320) );
XNOR2_X1 U1022 ( .A(n1225), .B(KEYINPUT19), .ZN(n1307) );
NOR2_X1 U1023 ( .A1(n1133), .A2(G953), .ZN(n1225) );
INV_X1 U1024 ( .A(G224), .ZN(n1133) );
XOR2_X1 U1025 ( .A(n1060), .B(n1064), .Z(n1089) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1284), .ZN(n1064) );
NAND2_X1 U1027 ( .A1(G234), .A2(n1287), .ZN(n1284) );
NAND2_X1 U1028 ( .A1(n1144), .A2(n1287), .ZN(n1060) );
NAND2_X1 U1029 ( .A1(n1322), .A2(n1323), .ZN(n1144) );
NAND2_X1 U1030 ( .A1(n1324), .A2(n1325), .ZN(n1323) );
XOR2_X1 U1031 ( .A(n1326), .B(KEYINPUT50), .Z(n1322) );
OR2_X1 U1032 ( .A1(n1325), .A2(n1324), .ZN(n1326) );
XOR2_X1 U1033 ( .A(n1327), .B(n1328), .Z(n1324) );
XNOR2_X1 U1034 ( .A(n1329), .B(n1173), .ZN(n1328) );
XNOR2_X1 U1035 ( .A(G110), .B(G140), .ZN(n1173) );
NOR2_X1 U1036 ( .A1(G128), .A2(KEYINPUT14), .ZN(n1329) );
XOR2_X1 U1037 ( .A(n1330), .B(n1331), .Z(n1327) );
XNOR2_X1 U1038 ( .A(n1332), .B(G119), .ZN(n1331) );
INV_X1 U1039 ( .A(G125), .ZN(n1332) );
NAND2_X1 U1040 ( .A1(KEYINPUT17), .A2(n1270), .ZN(n1330) );
XOR2_X1 U1041 ( .A(n1333), .B(n1334), .Z(n1325) );
NAND2_X1 U1042 ( .A1(G221), .A2(n1335), .ZN(n1333) );
INV_X1 U1043 ( .A(n1279), .ZN(n1335) );
NAND2_X1 U1044 ( .A1(G234), .A2(n1114), .ZN(n1279) );
INV_X1 U1045 ( .A(G953), .ZN(n1114) );
INV_X1 U1046 ( .A(n1053), .ZN(n1088) );
XOR2_X1 U1047 ( .A(n1336), .B(n1168), .Z(n1053) );
INV_X1 U1048 ( .A(G472), .ZN(n1168) );
NAND2_X1 U1049 ( .A1(n1337), .A2(n1287), .ZN(n1336) );
INV_X1 U1050 ( .A(G902), .ZN(n1287) );
XOR2_X1 U1051 ( .A(n1164), .B(n1338), .Z(n1337) );
XOR2_X1 U1052 ( .A(KEYINPUT5), .B(KEYINPUT16), .Z(n1338) );
XOR2_X1 U1053 ( .A(n1339), .B(n1340), .Z(n1164) );
XOR2_X1 U1054 ( .A(n1321), .B(n1341), .Z(n1340) );
XOR2_X1 U1055 ( .A(n1342), .B(n1292), .Z(n1341) );
XNOR2_X1 U1056 ( .A(n1123), .B(n1343), .ZN(n1292) );
NOR3_X1 U1057 ( .A1(n1129), .A2(KEYINPUT10), .A3(n1344), .ZN(n1343) );
INV_X1 U1058 ( .A(n1128), .ZN(n1344) );
NAND2_X1 U1059 ( .A1(G134), .A2(n1334), .ZN(n1128) );
NOR2_X1 U1060 ( .A1(n1334), .A2(G134), .ZN(n1129) );
XNOR2_X1 U1061 ( .A(G137), .B(KEYINPUT60), .ZN(n1334) );
XOR2_X1 U1062 ( .A(G131), .B(KEYINPUT12), .Z(n1123) );
NAND2_X1 U1063 ( .A1(n1272), .A2(G210), .ZN(n1342) );
NOR2_X1 U1064 ( .A1(G953), .A2(G237), .ZN(n1272) );
XOR2_X1 U1065 ( .A(n1283), .B(n1345), .Z(n1321) );
NOR2_X1 U1066 ( .A1(KEYINPUT53), .A2(n1270), .ZN(n1345) );
INV_X1 U1067 ( .A(G146), .ZN(n1270) );
XNOR2_X1 U1068 ( .A(n1228), .B(G128), .ZN(n1283) );
INV_X1 U1069 ( .A(G143), .ZN(n1228) );
XOR2_X1 U1070 ( .A(n1346), .B(n1347), .Z(n1339) );
XNOR2_X1 U1071 ( .A(G113), .B(n1243), .ZN(n1347) );
INV_X1 U1072 ( .A(G101), .ZN(n1243) );
NAND2_X1 U1073 ( .A1(n1348), .A2(n1349), .ZN(n1346) );
NAND2_X1 U1074 ( .A1(G116), .A2(n1319), .ZN(n1349) );
XOR2_X1 U1075 ( .A(KEYINPUT35), .B(n1350), .Z(n1348) );
NOR2_X1 U1076 ( .A1(G116), .A2(n1319), .ZN(n1350) );
INV_X1 U1077 ( .A(G119), .ZN(n1319) );
endmodule


