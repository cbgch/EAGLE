//Key = 0110100101000000101111110110011011010011000110111011001010011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355;

XOR2_X1 U741 ( .A(n1033), .B(n1034), .Z(G9) );
XNOR2_X1 U742 ( .A(KEYINPUT6), .B(n1035), .ZN(n1034) );
NOR2_X1 U743 ( .A1(n1036), .A2(n1037), .ZN(G75) );
NOR3_X1 U744 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
INV_X1 U745 ( .A(G952), .ZN(n1039) );
NAND3_X1 U746 ( .A1(n1041), .A2(n1042), .A3(n1043), .ZN(n1038) );
NAND2_X1 U747 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U748 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND4_X1 U749 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
NAND2_X1 U750 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND3_X1 U751 ( .A1(n1054), .A2(n1055), .A3(KEYINPUT9), .ZN(n1053) );
INV_X1 U752 ( .A(n1056), .ZN(n1052) );
NAND2_X1 U753 ( .A1(n1057), .A2(n1058), .ZN(n1046) );
NAND3_X1 U754 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
NAND3_X1 U755 ( .A1(n1050), .A2(n1062), .A3(n1048), .ZN(n1061) );
NAND3_X1 U756 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1062) );
NAND2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
INV_X1 U758 ( .A(n1068), .ZN(n1064) );
NAND2_X1 U759 ( .A1(n1049), .A2(n1069), .ZN(n1063) );
INV_X1 U760 ( .A(KEYINPUT9), .ZN(n1069) );
NAND2_X1 U761 ( .A1(n1049), .A2(n1070), .ZN(n1060) );
NAND3_X1 U762 ( .A1(n1071), .A2(n1072), .A3(n1073), .ZN(n1070) );
NAND2_X1 U763 ( .A1(KEYINPUT21), .A2(n1074), .ZN(n1073) );
NAND3_X1 U764 ( .A1(n1075), .A2(n1050), .A3(n1076), .ZN(n1072) );
NAND2_X1 U765 ( .A1(n1048), .A2(n1077), .ZN(n1071) );
NAND2_X1 U766 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
OR3_X1 U767 ( .A1(n1080), .A2(KEYINPUT21), .A3(n1049), .ZN(n1059) );
INV_X1 U768 ( .A(n1081), .ZN(n1044) );
NOR3_X1 U769 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1036) );
NOR2_X1 U770 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U771 ( .A(KEYINPUT19), .ZN(n1086) );
NOR2_X1 U772 ( .A1(G953), .A2(G952), .ZN(n1085) );
NOR2_X1 U773 ( .A1(KEYINPUT19), .A2(n1087), .ZN(n1083) );
INV_X1 U774 ( .A(n1041), .ZN(n1082) );
NAND4_X1 U775 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1041) );
NOR4_X1 U776 ( .A1(n1076), .A2(n1054), .A3(n1092), .A4(n1093), .ZN(n1091) );
NOR2_X1 U777 ( .A1(n1094), .A2(n1095), .ZN(n1090) );
XOR2_X1 U778 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U779 ( .A1(KEYINPUT56), .A2(G472), .ZN(n1097) );
XNOR2_X1 U780 ( .A(n1098), .B(n1099), .ZN(n1089) );
XOR2_X1 U781 ( .A(n1100), .B(n1101), .Z(n1088) );
XOR2_X1 U782 ( .A(n1102), .B(n1103), .Z(G72) );
XOR2_X1 U783 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR3_X1 U784 ( .A1(n1106), .A2(KEYINPUT53), .A3(G953), .ZN(n1105) );
NOR3_X1 U785 ( .A1(n1107), .A2(n1108), .A3(n1109), .ZN(n1106) );
NAND2_X1 U786 ( .A1(n1110), .A2(n1111), .ZN(n1104) );
NAND2_X1 U787 ( .A1(G900), .A2(G227), .ZN(n1111) );
XNOR2_X1 U788 ( .A(G953), .B(KEYINPUT51), .ZN(n1110) );
NAND2_X1 U789 ( .A1(n1112), .A2(n1113), .ZN(n1102) );
NAND2_X1 U790 ( .A1(G953), .A2(n1114), .ZN(n1113) );
XOR2_X1 U791 ( .A(n1115), .B(n1116), .Z(n1112) );
XNOR2_X1 U792 ( .A(n1117), .B(n1118), .ZN(n1116) );
XNOR2_X1 U793 ( .A(KEYINPUT37), .B(n1119), .ZN(n1118) );
INV_X1 U794 ( .A(G140), .ZN(n1119) );
XOR2_X1 U795 ( .A(n1120), .B(n1121), .Z(n1115) );
NOR2_X1 U796 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U797 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XNOR2_X1 U798 ( .A(G134), .B(KEYINPUT39), .ZN(n1125) );
NOR2_X1 U799 ( .A1(G137), .A2(n1126), .ZN(n1122) );
XNOR2_X1 U800 ( .A(G134), .B(KEYINPUT40), .ZN(n1126) );
XNOR2_X1 U801 ( .A(n1127), .B(n1128), .ZN(n1120) );
NAND2_X1 U802 ( .A1(KEYINPUT50), .A2(n1129), .ZN(n1127) );
NAND2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(G69) );
NAND2_X1 U804 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
OR2_X1 U805 ( .A1(n1042), .A2(G224), .ZN(n1133) );
NAND3_X1 U806 ( .A1(G953), .A2(n1134), .A3(n1135), .ZN(n1130) );
INV_X1 U807 ( .A(n1132), .ZN(n1135) );
XNOR2_X1 U808 ( .A(n1136), .B(n1137), .ZN(n1132) );
NOR3_X1 U809 ( .A1(n1138), .A2(KEYINPUT24), .A3(n1139), .ZN(n1137) );
XOR2_X1 U810 ( .A(n1140), .B(n1141), .Z(n1138) );
NAND2_X1 U811 ( .A1(n1142), .A2(KEYINPUT47), .ZN(n1141) );
XNOR2_X1 U812 ( .A(G110), .B(G122), .ZN(n1142) );
NAND3_X1 U813 ( .A1(n1143), .A2(n1144), .A3(n1145), .ZN(n1140) );
OR2_X1 U814 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
NAND3_X1 U815 ( .A1(n1147), .A2(n1146), .A3(KEYINPUT4), .ZN(n1144) );
NOR2_X1 U816 ( .A1(KEYINPUT14), .A2(n1148), .ZN(n1147) );
NAND2_X1 U817 ( .A1(n1148), .A2(n1149), .ZN(n1143) );
INV_X1 U818 ( .A(KEYINPUT4), .ZN(n1149) );
XNOR2_X1 U819 ( .A(n1150), .B(G107), .ZN(n1148) );
NAND2_X1 U820 ( .A1(n1151), .A2(n1042), .ZN(n1136) );
XOR2_X1 U821 ( .A(KEYINPUT44), .B(n1152), .Z(n1151) );
NAND2_X1 U822 ( .A1(G898), .A2(G224), .ZN(n1134) );
NOR2_X1 U823 ( .A1(n1153), .A2(n1154), .ZN(G66) );
XNOR2_X1 U824 ( .A(n1087), .B(KEYINPUT16), .ZN(n1154) );
XOR2_X1 U825 ( .A(n1155), .B(n1156), .Z(n1153) );
XOR2_X1 U826 ( .A(KEYINPUT63), .B(n1157), .Z(n1156) );
NOR2_X1 U827 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
NOR2_X1 U828 ( .A1(n1087), .A2(n1160), .ZN(G63) );
XNOR2_X1 U829 ( .A(n1161), .B(n1162), .ZN(n1160) );
NOR2_X1 U830 ( .A1(n1163), .A2(n1159), .ZN(n1161) );
NOR2_X1 U831 ( .A1(n1087), .A2(n1164), .ZN(G60) );
XOR2_X1 U832 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND3_X1 U833 ( .A1(G475), .A2(n1040), .A3(n1167), .ZN(n1165) );
XNOR2_X1 U834 ( .A(G902), .B(KEYINPUT59), .ZN(n1167) );
XOR2_X1 U835 ( .A(n1168), .B(G104), .Z(G6) );
NAND2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NAND2_X1 U837 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
INV_X1 U838 ( .A(KEYINPUT12), .ZN(n1172) );
NAND3_X1 U839 ( .A1(n1173), .A2(n1079), .A3(KEYINPUT12), .ZN(n1169) );
NOR2_X1 U840 ( .A1(n1087), .A2(n1174), .ZN(G57) );
XOR2_X1 U841 ( .A(n1175), .B(n1176), .Z(n1174) );
XNOR2_X1 U842 ( .A(n1177), .B(n1178), .ZN(n1176) );
XOR2_X1 U843 ( .A(n1179), .B(n1180), .Z(n1175) );
NOR2_X1 U844 ( .A1(n1181), .A2(n1159), .ZN(n1180) );
NAND2_X1 U845 ( .A1(KEYINPUT33), .A2(n1182), .ZN(n1179) );
NOR2_X1 U846 ( .A1(n1087), .A2(n1183), .ZN(G54) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U848 ( .A(KEYINPUT11), .B(n1186), .Z(n1185) );
NOR2_X1 U849 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U850 ( .A(n1189), .B(n1190), .Z(n1188) );
INV_X1 U851 ( .A(n1191), .ZN(n1187) );
NOR2_X1 U852 ( .A1(n1192), .A2(n1191), .ZN(n1184) );
NAND3_X1 U853 ( .A1(n1193), .A2(n1194), .A3(G469), .ZN(n1191) );
NAND2_X1 U854 ( .A1(KEYINPUT30), .A2(n1159), .ZN(n1194) );
NAND2_X1 U855 ( .A1(n1195), .A2(n1196), .ZN(n1193) );
INV_X1 U856 ( .A(KEYINPUT30), .ZN(n1196) );
OR2_X1 U857 ( .A1(n1040), .A2(n1197), .ZN(n1195) );
XNOR2_X1 U858 ( .A(n1190), .B(n1189), .ZN(n1192) );
NOR2_X1 U859 ( .A1(KEYINPUT34), .A2(n1198), .ZN(n1189) );
XOR2_X1 U860 ( .A(n1199), .B(n1200), .Z(n1198) );
NOR2_X1 U861 ( .A1(KEYINPUT62), .A2(n1201), .ZN(n1200) );
NOR2_X1 U862 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
XOR2_X1 U863 ( .A(n1204), .B(KEYINPUT35), .Z(n1203) );
NAND2_X1 U864 ( .A1(n1128), .A2(n1205), .ZN(n1204) );
NOR2_X1 U865 ( .A1(n1128), .A2(n1205), .ZN(n1202) );
NOR2_X1 U866 ( .A1(n1087), .A2(n1206), .ZN(G51) );
NOR2_X1 U867 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U868 ( .A(n1209), .B(KEYINPUT48), .Z(n1208) );
NAND2_X1 U869 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NOR2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(n1207) );
AND2_X1 U871 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND2_X1 U872 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
NAND2_X1 U873 ( .A1(n1216), .A2(n1217), .ZN(n1215) );
NAND3_X1 U874 ( .A1(n1216), .A2(n1217), .A3(n1218), .ZN(n1212) );
XOR2_X1 U875 ( .A(n1219), .B(KEYINPUT15), .Z(n1216) );
NOR2_X1 U876 ( .A1(n1159), .A2(n1101), .ZN(n1210) );
NAND2_X1 U877 ( .A1(G902), .A2(n1040), .ZN(n1159) );
NAND3_X1 U878 ( .A1(n1152), .A2(n1220), .A3(n1221), .ZN(n1040) );
XOR2_X1 U879 ( .A(n1222), .B(KEYINPUT20), .Z(n1221) );
NAND2_X1 U880 ( .A1(n1223), .A2(n1224), .ZN(n1222) );
INV_X1 U881 ( .A(n1109), .ZN(n1224) );
NAND3_X1 U882 ( .A1(n1225), .A2(n1226), .A3(n1227), .ZN(n1109) );
NAND2_X1 U883 ( .A1(n1228), .A2(n1057), .ZN(n1227) );
NAND3_X1 U884 ( .A1(n1229), .A2(n1056), .A3(n1230), .ZN(n1225) );
XNOR2_X1 U885 ( .A(n1108), .B(KEYINPUT17), .ZN(n1223) );
INV_X1 U886 ( .A(n1107), .ZN(n1220) );
NAND3_X1 U887 ( .A1(n1231), .A2(n1232), .A3(n1233), .ZN(n1107) );
NAND2_X1 U888 ( .A1(n1234), .A2(n1235), .ZN(n1233) );
NAND2_X1 U889 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
NAND2_X1 U890 ( .A1(n1238), .A2(n1057), .ZN(n1237) );
NAND2_X1 U891 ( .A1(n1230), .A2(n1056), .ZN(n1236) );
AND2_X1 U892 ( .A1(n1239), .A2(n1240), .ZN(n1152) );
AND4_X1 U893 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1240) );
NOR4_X1 U894 ( .A1(n1245), .A2(n1246), .A3(n1033), .A4(n1171), .ZN(n1239) );
AND2_X1 U895 ( .A1(n1229), .A2(n1173), .ZN(n1171) );
AND2_X1 U896 ( .A1(n1234), .A2(n1173), .ZN(n1033) );
AND4_X1 U897 ( .A1(n1056), .A2(n1247), .A3(n1049), .A4(n1248), .ZN(n1173) );
NOR2_X1 U898 ( .A1(n1042), .A2(G952), .ZN(n1087) );
XOR2_X1 U899 ( .A(G146), .B(n1249), .Z(G48) );
NOR3_X1 U900 ( .A1(n1250), .A2(n1251), .A3(n1079), .ZN(n1249) );
XNOR2_X1 U901 ( .A(n1056), .B(KEYINPUT5), .ZN(n1251) );
XNOR2_X1 U902 ( .A(G143), .B(n1252), .ZN(G45) );
NOR2_X1 U903 ( .A1(n1108), .A2(KEYINPUT8), .ZN(n1252) );
AND4_X1 U904 ( .A1(n1253), .A2(n1238), .A3(n1056), .A4(n1094), .ZN(n1108) );
XNOR2_X1 U905 ( .A(G140), .B(n1254), .ZN(G42) );
NAND2_X1 U906 ( .A1(n1057), .A2(n1255), .ZN(n1254) );
XOR2_X1 U907 ( .A(KEYINPUT58), .B(n1228), .Z(n1255) );
AND2_X1 U908 ( .A1(n1256), .A2(n1247), .ZN(n1228) );
XNOR2_X1 U909 ( .A(G137), .B(n1226), .ZN(G39) );
NAND3_X1 U910 ( .A1(n1057), .A2(n1050), .A3(n1230), .ZN(n1226) );
INV_X1 U911 ( .A(n1250), .ZN(n1230) );
XNOR2_X1 U912 ( .A(G134), .B(n1257), .ZN(G36) );
NAND3_X1 U913 ( .A1(n1234), .A2(n1258), .A3(n1238), .ZN(n1257) );
XOR2_X1 U914 ( .A(KEYINPUT10), .B(n1057), .Z(n1258) );
XNOR2_X1 U915 ( .A(G131), .B(n1231), .ZN(G33) );
NAND3_X1 U916 ( .A1(n1057), .A2(n1229), .A3(n1238), .ZN(n1231) );
AND3_X1 U917 ( .A1(n1247), .A2(n1259), .A3(n1068), .ZN(n1238) );
AND2_X1 U918 ( .A1(n1055), .A2(n1260), .ZN(n1057) );
XNOR2_X1 U919 ( .A(G128), .B(n1261), .ZN(G30) );
NAND2_X1 U920 ( .A1(n1056), .A2(n1262), .ZN(n1261) );
XOR2_X1 U921 ( .A(KEYINPUT0), .B(n1263), .Z(n1262) );
NOR2_X1 U922 ( .A1(n1078), .A2(n1250), .ZN(n1263) );
NAND4_X1 U923 ( .A1(n1066), .A2(n1247), .A3(n1264), .A4(n1259), .ZN(n1250) );
INV_X1 U924 ( .A(n1234), .ZN(n1078) );
XOR2_X1 U925 ( .A(G101), .B(n1246), .Z(G3) );
AND2_X1 U926 ( .A1(n1068), .A2(n1265), .ZN(n1246) );
XNOR2_X1 U927 ( .A(G125), .B(n1232), .ZN(G27) );
NAND3_X1 U928 ( .A1(n1048), .A2(n1056), .A3(n1256), .ZN(n1232) );
AND4_X1 U929 ( .A1(n1066), .A2(n1229), .A3(n1067), .A4(n1259), .ZN(n1256) );
NAND2_X1 U930 ( .A1(n1081), .A2(n1266), .ZN(n1259) );
NAND4_X1 U931 ( .A1(G953), .A2(G902), .A3(n1267), .A4(n1114), .ZN(n1266) );
INV_X1 U932 ( .A(G900), .ZN(n1114) );
XOR2_X1 U933 ( .A(G122), .B(n1245), .Z(G24) );
AND4_X1 U934 ( .A1(n1253), .A2(n1268), .A3(n1049), .A4(n1094), .ZN(n1245) );
NOR2_X1 U935 ( .A1(n1264), .A2(n1066), .ZN(n1049) );
XOR2_X1 U936 ( .A(n1244), .B(n1269), .Z(G21) );
NAND2_X1 U937 ( .A1(KEYINPUT23), .A2(G119), .ZN(n1269) );
NAND4_X1 U938 ( .A1(n1066), .A2(n1268), .A3(n1050), .A4(n1264), .ZN(n1244) );
XNOR2_X1 U939 ( .A(G116), .B(n1243), .ZN(G18) );
NAND3_X1 U940 ( .A1(n1068), .A2(n1234), .A3(n1268), .ZN(n1243) );
XNOR2_X1 U941 ( .A(G113), .B(n1242), .ZN(G15) );
NAND3_X1 U942 ( .A1(n1068), .A2(n1229), .A3(n1268), .ZN(n1242) );
AND3_X1 U943 ( .A1(n1056), .A2(n1248), .A3(n1048), .ZN(n1268) );
NOR2_X1 U944 ( .A1(n1270), .A2(n1076), .ZN(n1048) );
INV_X1 U945 ( .A(n1079), .ZN(n1229) );
NAND2_X1 U946 ( .A1(n1253), .A2(n1271), .ZN(n1079) );
XNOR2_X1 U947 ( .A(n1093), .B(KEYINPUT2), .ZN(n1253) );
NOR2_X1 U948 ( .A1(n1066), .A2(n1067), .ZN(n1068) );
XNOR2_X1 U949 ( .A(G110), .B(n1241), .ZN(G12) );
NAND3_X1 U950 ( .A1(n1067), .A2(n1066), .A3(n1265), .ZN(n1241) );
AND3_X1 U951 ( .A1(n1056), .A2(n1248), .A3(n1074), .ZN(n1265) );
INV_X1 U952 ( .A(n1080), .ZN(n1074) );
NAND2_X1 U953 ( .A1(n1247), .A2(n1050), .ZN(n1080) );
NAND2_X1 U954 ( .A1(n1272), .A2(n1273), .ZN(n1050) );
OR3_X1 U955 ( .A1(n1093), .A2(n1094), .A3(KEYINPUT42), .ZN(n1273) );
NAND2_X1 U956 ( .A1(KEYINPUT42), .A2(n1234), .ZN(n1272) );
NOR2_X1 U957 ( .A1(n1093), .A2(n1271), .ZN(n1234) );
INV_X1 U958 ( .A(n1094), .ZN(n1271) );
XOR2_X1 U959 ( .A(n1274), .B(n1163), .Z(n1094) );
INV_X1 U960 ( .A(G478), .ZN(n1163) );
NAND2_X1 U961 ( .A1(n1162), .A2(n1275), .ZN(n1274) );
XOR2_X1 U962 ( .A(n1276), .B(n1277), .Z(n1162) );
XOR2_X1 U963 ( .A(n1278), .B(n1279), .Z(n1277) );
NOR4_X1 U964 ( .A1(KEYINPUT27), .A2(G953), .A3(n1280), .A4(n1281), .ZN(n1278) );
INV_X1 U965 ( .A(G217), .ZN(n1280) );
XNOR2_X1 U966 ( .A(G116), .B(n1282), .ZN(n1276) );
NOR2_X1 U967 ( .A1(KEYINPUT28), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U968 ( .A(n1284), .B(n1285), .ZN(n1283) );
XOR2_X1 U969 ( .A(KEYINPUT57), .B(G134), .Z(n1285) );
XNOR2_X1 U970 ( .A(n1286), .B(G475), .ZN(n1093) );
NAND2_X1 U971 ( .A1(n1166), .A2(n1275), .ZN(n1286) );
XNOR2_X1 U972 ( .A(n1287), .B(n1288), .ZN(n1166) );
XNOR2_X1 U973 ( .A(G140), .B(n1289), .ZN(n1288) );
NAND2_X1 U974 ( .A1(n1290), .A2(KEYINPUT18), .ZN(n1289) );
XOR2_X1 U975 ( .A(n1291), .B(n1292), .Z(n1290) );
NAND2_X1 U976 ( .A1(KEYINPUT43), .A2(n1293), .ZN(n1291) );
XOR2_X1 U977 ( .A(G122), .B(G113), .Z(n1293) );
XOR2_X1 U978 ( .A(n1294), .B(n1295), .Z(n1287) );
NAND2_X1 U979 ( .A1(KEYINPUT32), .A2(n1296), .ZN(n1294) );
XNOR2_X1 U980 ( .A(n1117), .B(n1297), .ZN(n1296) );
NOR2_X1 U981 ( .A1(KEYINPUT13), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U982 ( .A(G143), .B(n1299), .ZN(n1298) );
NAND3_X1 U983 ( .A1(n1300), .A2(n1042), .A3(G214), .ZN(n1299) );
NOR2_X1 U984 ( .A1(n1076), .A2(n1075), .ZN(n1247) );
INV_X1 U985 ( .A(n1270), .ZN(n1075) );
NAND3_X1 U986 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1270) );
OR2_X1 U987 ( .A1(n1098), .A2(KEYINPUT46), .ZN(n1303) );
NAND3_X1 U988 ( .A1(KEYINPUT46), .A2(n1098), .A3(G469), .ZN(n1302) );
NAND2_X1 U989 ( .A1(n1304), .A2(n1099), .ZN(n1301) );
INV_X1 U990 ( .A(G469), .ZN(n1099) );
NAND2_X1 U991 ( .A1(KEYINPUT46), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U992 ( .A(KEYINPUT29), .B(n1098), .ZN(n1305) );
NAND2_X1 U993 ( .A1(n1306), .A2(n1275), .ZN(n1098) );
XOR2_X1 U994 ( .A(n1307), .B(n1308), .Z(n1306) );
XNOR2_X1 U995 ( .A(n1190), .B(n1205), .ZN(n1308) );
XNOR2_X1 U996 ( .A(n1309), .B(G101), .ZN(n1205) );
NAND2_X1 U997 ( .A1(n1310), .A2(KEYINPUT1), .ZN(n1309) );
XNOR2_X1 U998 ( .A(G107), .B(n1292), .ZN(n1310) );
XNOR2_X1 U999 ( .A(n1311), .B(n1312), .ZN(n1190) );
NAND2_X1 U1000 ( .A1(G227), .A2(n1042), .ZN(n1311) );
XOR2_X1 U1001 ( .A(n1182), .B(KEYINPUT25), .Z(n1307) );
AND2_X1 U1002 ( .A1(G221), .A2(n1313), .ZN(n1076) );
NAND2_X1 U1003 ( .A1(n1081), .A2(n1314), .ZN(n1248) );
NAND3_X1 U1004 ( .A1(G902), .A2(n1267), .A3(n1139), .ZN(n1314) );
NOR2_X1 U1005 ( .A1(n1042), .A2(G898), .ZN(n1139) );
NAND3_X1 U1006 ( .A1(n1267), .A2(n1042), .A3(G952), .ZN(n1081) );
NAND2_X1 U1007 ( .A1(G237), .A2(n1315), .ZN(n1267) );
NOR2_X1 U1008 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
INV_X1 U1009 ( .A(n1260), .ZN(n1054) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1316), .ZN(n1260) );
XNOR2_X1 U1011 ( .A(n1101), .B(n1317), .ZN(n1055) );
NOR2_X1 U1012 ( .A1(n1100), .A2(KEYINPUT45), .ZN(n1317) );
AND2_X1 U1013 ( .A1(n1318), .A2(n1275), .ZN(n1100) );
XNOR2_X1 U1014 ( .A(n1319), .B(n1214), .ZN(n1318) );
INV_X1 U1015 ( .A(n1218), .ZN(n1214) );
XNOR2_X1 U1016 ( .A(n1320), .B(n1321), .ZN(n1218) );
XNOR2_X1 U1017 ( .A(n1322), .B(n1279), .ZN(n1321) );
XNOR2_X1 U1018 ( .A(n1035), .B(G122), .ZN(n1279) );
INV_X1 U1019 ( .A(G107), .ZN(n1035) );
INV_X1 U1020 ( .A(n1150), .ZN(n1322) );
XOR2_X1 U1021 ( .A(G101), .B(n1292), .Z(n1150) );
XOR2_X1 U1022 ( .A(G104), .B(KEYINPUT31), .Z(n1292) );
XOR2_X1 U1023 ( .A(n1323), .B(n1324), .Z(n1320) );
NOR2_X1 U1024 ( .A1(KEYINPUT61), .A2(n1325), .ZN(n1324) );
XNOR2_X1 U1025 ( .A(KEYINPUT3), .B(n1146), .ZN(n1325) );
NAND2_X1 U1026 ( .A1(n1326), .A2(n1327), .ZN(n1146) );
NAND2_X1 U1027 ( .A1(n1328), .A2(G119), .ZN(n1327) );
NAND2_X1 U1028 ( .A1(n1329), .A2(n1330), .ZN(n1326) );
INV_X1 U1029 ( .A(G119), .ZN(n1330) );
XNOR2_X1 U1030 ( .A(n1328), .B(KEYINPUT49), .ZN(n1329) );
XNOR2_X1 U1031 ( .A(G110), .B(KEYINPUT54), .ZN(n1323) );
NOR2_X1 U1032 ( .A1(n1331), .A2(KEYINPUT52), .ZN(n1319) );
AND2_X1 U1033 ( .A1(n1219), .A2(n1217), .ZN(n1331) );
NAND3_X1 U1034 ( .A1(G224), .A2(n1042), .A3(n1332), .ZN(n1217) );
XOR2_X1 U1035 ( .A(n1284), .B(n1295), .Z(n1332) );
NAND2_X1 U1036 ( .A1(n1333), .A2(n1334), .ZN(n1219) );
NAND2_X1 U1037 ( .A1(G224), .A2(n1042), .ZN(n1334) );
XNOR2_X1 U1038 ( .A(n1295), .B(n1284), .ZN(n1333) );
NAND2_X1 U1039 ( .A1(G210), .A2(n1316), .ZN(n1101) );
NAND2_X1 U1040 ( .A1(n1335), .A2(n1197), .ZN(n1316) );
INV_X1 U1041 ( .A(G237), .ZN(n1335) );
XNOR2_X1 U1042 ( .A(n1092), .B(KEYINPUT26), .ZN(n1066) );
XOR2_X1 U1043 ( .A(n1336), .B(n1158), .Z(n1092) );
NAND2_X1 U1044 ( .A1(G217), .A2(n1313), .ZN(n1158) );
NAND2_X1 U1045 ( .A1(n1315), .A2(n1197), .ZN(n1313) );
XOR2_X1 U1046 ( .A(G234), .B(KEYINPUT55), .Z(n1315) );
NAND2_X1 U1047 ( .A1(n1155), .A2(n1275), .ZN(n1336) );
XOR2_X1 U1048 ( .A(n1337), .B(n1338), .Z(n1155) );
XOR2_X1 U1049 ( .A(n1295), .B(n1312), .Z(n1338) );
XNOR2_X1 U1050 ( .A(n1339), .B(G140), .ZN(n1312) );
INV_X1 U1051 ( .A(G110), .ZN(n1339) );
XNOR2_X1 U1052 ( .A(n1129), .B(G146), .ZN(n1295) );
INV_X1 U1053 ( .A(G125), .ZN(n1129) );
XOR2_X1 U1054 ( .A(n1340), .B(n1341), .Z(n1337) );
NOR3_X1 U1055 ( .A1(n1342), .A2(G953), .A3(n1281), .ZN(n1341) );
XOR2_X1 U1056 ( .A(G234), .B(KEYINPUT38), .Z(n1281) );
INV_X1 U1057 ( .A(G221), .ZN(n1342) );
XNOR2_X1 U1058 ( .A(n1343), .B(n1124), .ZN(n1340) );
INV_X1 U1059 ( .A(G137), .ZN(n1124) );
NAND2_X1 U1060 ( .A1(n1344), .A2(KEYINPUT60), .ZN(n1343) );
XNOR2_X1 U1061 ( .A(G128), .B(G119), .ZN(n1344) );
INV_X1 U1062 ( .A(n1264), .ZN(n1067) );
XOR2_X1 U1063 ( .A(n1096), .B(n1181), .Z(n1264) );
INV_X1 U1064 ( .A(G472), .ZN(n1181) );
NAND2_X1 U1065 ( .A1(n1345), .A2(n1346), .ZN(n1096) );
XNOR2_X1 U1066 ( .A(n1178), .B(n1347), .ZN(n1346) );
XNOR2_X1 U1067 ( .A(n1182), .B(n1348), .ZN(n1347) );
INV_X1 U1068 ( .A(n1177), .ZN(n1348) );
XNOR2_X1 U1069 ( .A(n1349), .B(G101), .ZN(n1177) );
NAND3_X1 U1070 ( .A1(n1300), .A2(n1042), .A3(G210), .ZN(n1349) );
INV_X1 U1071 ( .A(G953), .ZN(n1042) );
XNOR2_X1 U1072 ( .A(G237), .B(KEYINPUT36), .ZN(n1300) );
XNOR2_X1 U1073 ( .A(n1199), .B(n1128), .ZN(n1182) );
XOR2_X1 U1074 ( .A(G146), .B(n1284), .Z(n1128) );
XOR2_X1 U1075 ( .A(G128), .B(n1350), .Z(n1284) );
INV_X1 U1076 ( .A(G143), .ZN(n1350) );
NAND2_X1 U1077 ( .A1(n1351), .A2(n1352), .ZN(n1199) );
NAND2_X1 U1078 ( .A1(n1353), .A2(n1117), .ZN(n1352) );
XOR2_X1 U1079 ( .A(KEYINPUT22), .B(n1354), .Z(n1351) );
NOR2_X1 U1080 ( .A1(n1353), .A2(n1117), .ZN(n1354) );
INV_X1 U1081 ( .A(G131), .ZN(n1117) );
XNOR2_X1 U1082 ( .A(G134), .B(G137), .ZN(n1353) );
XOR2_X1 U1083 ( .A(G119), .B(n1328), .Z(n1178) );
XNOR2_X1 U1084 ( .A(G113), .B(n1355), .ZN(n1328) );
INV_X1 U1085 ( .A(G116), .ZN(n1355) );
XOR2_X1 U1086 ( .A(KEYINPUT41), .B(n1275), .Z(n1345) );
XNOR2_X1 U1087 ( .A(n1197), .B(KEYINPUT7), .ZN(n1275) );
INV_X1 U1088 ( .A(G902), .ZN(n1197) );
endmodule


