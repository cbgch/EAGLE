//Key = 1111000011101001100101011101011010111001110010001000101000011110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
n1396, n1397, n1398, n1399;

NAND2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(G9) );
NAND2_X1 U770 ( .A1(G107), .A2(n1068), .ZN(n1067) );
XOR2_X1 U771 ( .A(n1069), .B(KEYINPUT55), .Z(n1066) );
OR2_X1 U772 ( .A1(n1068), .A2(G107), .ZN(n1069) );
NOR2_X1 U773 ( .A1(n1070), .A2(n1071), .ZN(G75) );
NOR4_X1 U774 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1071) );
NOR3_X1 U775 ( .A1(n1076), .A2(n1077), .A3(n1078), .ZN(n1074) );
NOR3_X1 U776 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
AND3_X1 U777 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1081) );
OR2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U779 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR2_X1 U780 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
NOR2_X1 U781 ( .A1(n1091), .A2(n1092), .ZN(n1085) );
NOR2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NOR2_X1 U783 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
AND3_X1 U784 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1080) );
XNOR2_X1 U785 ( .A(n1083), .B(KEYINPUT41), .ZN(n1098) );
XOR2_X1 U786 ( .A(n1100), .B(KEYINPUT48), .Z(n1079) );
NAND3_X1 U787 ( .A1(n1101), .A2(n1083), .A3(n1097), .ZN(n1100) );
NAND3_X1 U788 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1072) );
NAND4_X1 U789 ( .A1(n1097), .A2(n1082), .A3(n1105), .A4(n1083), .ZN(n1104) );
NAND2_X1 U790 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
NAND2_X1 U791 ( .A1(n1077), .A2(n1108), .ZN(n1107) );
NOR3_X1 U792 ( .A1(n1109), .A2(G953), .A3(G952), .ZN(n1070) );
INV_X1 U793 ( .A(n1102), .ZN(n1109) );
NAND4_X1 U794 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1102) );
NOR4_X1 U795 ( .A1(n1114), .A2(n1077), .A3(n1115), .A4(n1116), .ZN(n1113) );
NOR2_X1 U796 ( .A1(KEYINPUT2), .A2(n1117), .ZN(n1116) );
XOR2_X1 U797 ( .A(n1118), .B(KEYINPUT52), .Z(n1115) );
INV_X1 U798 ( .A(n1119), .ZN(n1077) );
NOR3_X1 U799 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1112) );
NOR2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1122) );
NOR2_X1 U801 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
XOR2_X1 U802 ( .A(n1117), .B(KEYINPUT59), .Z(n1125) );
NOR3_X1 U803 ( .A1(n1127), .A2(n1128), .A3(n1126), .ZN(n1121) );
INV_X1 U804 ( .A(KEYINPUT2), .ZN(n1126) );
INV_X1 U805 ( .A(n1117), .ZN(n1128) );
XOR2_X1 U806 ( .A(n1129), .B(n1130), .Z(n1120) );
XOR2_X1 U807 ( .A(n1131), .B(KEYINPUT53), .Z(n1130) );
XNOR2_X1 U808 ( .A(n1132), .B(n1133), .ZN(n1110) );
XOR2_X1 U809 ( .A(KEYINPUT49), .B(G478), .Z(n1133) );
XOR2_X1 U810 ( .A(n1134), .B(n1135), .Z(G72) );
NOR2_X1 U811 ( .A1(n1136), .A2(n1103), .ZN(n1135) );
AND2_X1 U812 ( .A1(G227), .A2(G900), .ZN(n1136) );
NOR3_X1 U813 ( .A1(KEYINPUT13), .A2(n1137), .A3(n1138), .ZN(n1134) );
NOR2_X1 U814 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U816 ( .A1(G900), .A2(n1103), .ZN(n1141) );
INV_X1 U817 ( .A(n1143), .ZN(n1139) );
NOR2_X1 U818 ( .A1(n1142), .A2(n1143), .ZN(n1137) );
XOR2_X1 U819 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U820 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U821 ( .A(n1148), .B(n1149), .Z(n1144) );
NAND2_X1 U822 ( .A1(KEYINPUT61), .A2(n1150), .ZN(n1148) );
NOR2_X1 U823 ( .A1(G953), .A2(n1151), .ZN(n1142) );
NAND2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(G69) );
NAND3_X1 U825 ( .A1(n1154), .A2(n1155), .A3(n1156), .ZN(n1153) );
OR2_X1 U826 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
NAND2_X1 U827 ( .A1(n1159), .A2(n1158), .ZN(n1154) );
XOR2_X1 U828 ( .A(KEYINPUT29), .B(n1160), .Z(n1152) );
NOR3_X1 U829 ( .A1(n1156), .A2(n1158), .A3(n1157), .ZN(n1160) );
XNOR2_X1 U830 ( .A(n1159), .B(KEYINPUT34), .ZN(n1157) );
NOR2_X1 U831 ( .A1(G953), .A2(n1161), .ZN(n1159) );
AND3_X1 U832 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1158) );
NAND2_X1 U833 ( .A1(G953), .A2(n1165), .ZN(n1164) );
NAND2_X1 U834 ( .A1(KEYINPUT57), .A2(n1166), .ZN(n1163) );
NAND2_X1 U835 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
NAND2_X1 U836 ( .A1(n1169), .A2(n1170), .ZN(n1162) );
INV_X1 U837 ( .A(KEYINPUT57), .ZN(n1170) );
NAND2_X1 U838 ( .A1(G953), .A2(n1171), .ZN(n1156) );
NAND2_X1 U839 ( .A1(G898), .A2(G224), .ZN(n1171) );
NOR2_X1 U840 ( .A1(n1172), .A2(n1173), .ZN(G66) );
XOR2_X1 U841 ( .A(n1174), .B(n1175), .Z(n1173) );
NOR2_X1 U842 ( .A1(n1176), .A2(n1177), .ZN(n1174) );
NOR2_X1 U843 ( .A1(n1172), .A2(n1178), .ZN(G63) );
NOR3_X1 U844 ( .A1(n1132), .A2(n1179), .A3(n1180), .ZN(n1178) );
NOR3_X1 U845 ( .A1(n1181), .A2(n1182), .A3(n1177), .ZN(n1180) );
INV_X1 U846 ( .A(n1183), .ZN(n1181) );
NOR2_X1 U847 ( .A1(n1184), .A2(n1183), .ZN(n1179) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1182), .ZN(n1184) );
NOR2_X1 U849 ( .A1(n1075), .A2(n1073), .ZN(n1185) );
NOR2_X1 U850 ( .A1(n1172), .A2(n1186), .ZN(G60) );
XOR2_X1 U851 ( .A(n1187), .B(n1188), .Z(n1186) );
XNOR2_X1 U852 ( .A(KEYINPUT4), .B(n1189), .ZN(n1188) );
NOR2_X1 U853 ( .A1(n1190), .A2(n1177), .ZN(n1187) );
INV_X1 U854 ( .A(G475), .ZN(n1190) );
XNOR2_X1 U855 ( .A(G104), .B(n1191), .ZN(G6) );
NOR2_X1 U856 ( .A1(n1172), .A2(n1192), .ZN(G57) );
XOR2_X1 U857 ( .A(n1193), .B(n1194), .Z(n1192) );
XOR2_X1 U858 ( .A(n1195), .B(n1196), .Z(n1194) );
XOR2_X1 U859 ( .A(n1197), .B(n1198), .Z(n1195) );
NOR3_X1 U860 ( .A1(n1177), .A2(KEYINPUT43), .A3(n1199), .ZN(n1198) );
INV_X1 U861 ( .A(G472), .ZN(n1199) );
XOR2_X1 U862 ( .A(n1200), .B(n1201), .Z(n1193) );
XNOR2_X1 U863 ( .A(G101), .B(n1202), .ZN(n1201) );
NAND2_X1 U864 ( .A1(n1203), .A2(n1204), .ZN(n1200) );
NAND2_X1 U865 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U866 ( .A(KEYINPUT3), .B(n1207), .Z(n1203) );
NOR2_X1 U867 ( .A1(n1205), .A2(n1206), .ZN(n1207) );
NOR3_X1 U868 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(G54) );
NOR2_X1 U869 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
XOR2_X1 U870 ( .A(KEYINPUT11), .B(n1213), .Z(n1211) );
NOR2_X1 U871 ( .A1(n1214), .A2(n1215), .ZN(n1209) );
XNOR2_X1 U872 ( .A(n1213), .B(KEYINPUT14), .ZN(n1215) );
XNOR2_X1 U873 ( .A(n1216), .B(n1217), .ZN(n1213) );
XOR2_X1 U874 ( .A(n1218), .B(n1219), .Z(n1217) );
NOR2_X1 U875 ( .A1(n1131), .A2(n1177), .ZN(n1219) );
INV_X1 U876 ( .A(G469), .ZN(n1131) );
NOR2_X1 U877 ( .A1(KEYINPUT6), .A2(n1220), .ZN(n1218) );
INV_X1 U878 ( .A(n1212), .ZN(n1214) );
XOR2_X1 U879 ( .A(n1221), .B(n1222), .Z(n1212) );
XOR2_X1 U880 ( .A(KEYINPUT24), .B(KEYINPUT0), .Z(n1222) );
XOR2_X1 U881 ( .A(n1223), .B(n1224), .Z(n1221) );
XNOR2_X1 U882 ( .A(n1172), .B(KEYINPUT19), .ZN(n1208) );
NOR2_X1 U883 ( .A1(n1172), .A2(n1225), .ZN(G51) );
XOR2_X1 U884 ( .A(n1226), .B(n1227), .Z(n1225) );
XNOR2_X1 U885 ( .A(n1206), .B(n1228), .ZN(n1227) );
XOR2_X1 U886 ( .A(n1229), .B(n1230), .Z(n1226) );
NOR2_X1 U887 ( .A1(n1117), .A2(n1177), .ZN(n1229) );
NAND2_X1 U888 ( .A1(G902), .A2(n1231), .ZN(n1177) );
NAND2_X1 U889 ( .A1(n1161), .A2(n1151), .ZN(n1231) );
INV_X1 U890 ( .A(n1075), .ZN(n1151) );
NAND4_X1 U891 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1075) );
NOR4_X1 U892 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235) );
NOR2_X1 U893 ( .A1(n1240), .A2(n1241), .ZN(n1234) );
NOR3_X1 U894 ( .A1(n1242), .A2(n1243), .A3(n1244), .ZN(n1241) );
XOR2_X1 U895 ( .A(KEYINPUT15), .B(n1101), .Z(n1242) );
NAND2_X1 U896 ( .A1(n1245), .A2(n1246), .ZN(n1233) );
NAND2_X1 U897 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND4_X1 U898 ( .A1(n1249), .A2(n1250), .A3(n1251), .A4(n1252), .ZN(n1248) );
INV_X1 U899 ( .A(KEYINPUT9), .ZN(n1252) );
XNOR2_X1 U900 ( .A(n1253), .B(KEYINPUT26), .ZN(n1247) );
NAND2_X1 U901 ( .A1(KEYINPUT9), .A2(n1254), .ZN(n1232) );
INV_X1 U902 ( .A(n1073), .ZN(n1161) );
NAND4_X1 U903 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1073) );
AND4_X1 U904 ( .A1(n1259), .A2(n1191), .A3(n1068), .A4(n1260), .ZN(n1258) );
NAND3_X1 U905 ( .A1(n1111), .A2(n1099), .A3(n1261), .ZN(n1068) );
NAND3_X1 U906 ( .A1(n1261), .A2(n1111), .A3(n1101), .ZN(n1191) );
NOR2_X1 U907 ( .A1(n1262), .A2(n1263), .ZN(n1257) );
NOR2_X1 U908 ( .A1(n1264), .A2(n1243), .ZN(n1263) );
NOR2_X1 U909 ( .A1(n1265), .A2(n1106), .ZN(n1262) );
XOR2_X1 U910 ( .A(n1266), .B(KEYINPUT18), .Z(n1265) );
NAND3_X1 U911 ( .A1(n1090), .A2(n1099), .A3(n1267), .ZN(n1255) );
NOR2_X1 U912 ( .A1(n1103), .A2(G952), .ZN(n1172) );
XOR2_X1 U913 ( .A(n1268), .B(n1269), .Z(G48) );
NAND2_X1 U914 ( .A1(n1253), .A2(n1245), .ZN(n1269) );
AND2_X1 U915 ( .A1(n1270), .A2(n1101), .ZN(n1253) );
NAND3_X1 U916 ( .A1(n1271), .A2(n1272), .A3(n1273), .ZN(G45) );
OR2_X1 U917 ( .A1(n1274), .A2(n1254), .ZN(n1273) );
NAND2_X1 U918 ( .A1(n1275), .A2(n1276), .ZN(n1272) );
INV_X1 U919 ( .A(KEYINPUT25), .ZN(n1276) );
NAND2_X1 U920 ( .A1(n1277), .A2(n1254), .ZN(n1275) );
XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n1274), .ZN(n1277) );
NAND2_X1 U922 ( .A1(KEYINPUT25), .A2(n1278), .ZN(n1271) );
NAND2_X1 U923 ( .A1(n1279), .A2(n1280), .ZN(n1278) );
OR2_X1 U924 ( .A1(n1274), .A2(KEYINPUT39), .ZN(n1280) );
NAND3_X1 U925 ( .A1(n1254), .A2(n1274), .A3(KEYINPUT39), .ZN(n1279) );
XOR2_X1 U926 ( .A(G143), .B(KEYINPUT10), .Z(n1274) );
AND4_X1 U927 ( .A1(n1250), .A2(n1090), .A3(n1249), .A4(n1245), .ZN(n1254) );
AND3_X1 U928 ( .A1(n1094), .A2(n1281), .A3(n1282), .ZN(n1250) );
XOR2_X1 U929 ( .A(G140), .B(n1283), .Z(G42) );
NOR3_X1 U930 ( .A1(n1244), .A2(n1284), .A3(n1243), .ZN(n1283) );
XOR2_X1 U931 ( .A(G137), .B(n1240), .Z(G39) );
AND4_X1 U932 ( .A1(n1270), .A2(n1082), .A3(n1108), .A4(n1119), .ZN(n1240) );
XOR2_X1 U933 ( .A(G134), .B(n1239), .Z(G36) );
NOR3_X1 U934 ( .A1(n1251), .A2(n1285), .A3(n1244), .ZN(n1239) );
INV_X1 U935 ( .A(n1099), .ZN(n1285) );
XOR2_X1 U936 ( .A(G131), .B(n1238), .Z(G33) );
NOR3_X1 U937 ( .A1(n1284), .A2(n1251), .A3(n1244), .ZN(n1238) );
NAND4_X1 U938 ( .A1(n1282), .A2(n1094), .A3(n1108), .A4(n1119), .ZN(n1244) );
INV_X1 U939 ( .A(n1076), .ZN(n1108) );
XOR2_X1 U940 ( .A(G128), .B(n1237), .Z(G30) );
AND3_X1 U941 ( .A1(n1099), .A2(n1245), .A3(n1270), .ZN(n1237) );
AND4_X1 U942 ( .A1(n1282), .A2(n1094), .A3(n1286), .A4(n1287), .ZN(n1270) );
XNOR2_X1 U943 ( .A(G101), .B(n1259), .ZN(G3) );
OR2_X1 U944 ( .A1(n1251), .A2(n1264), .ZN(n1259) );
INV_X1 U945 ( .A(n1090), .ZN(n1251) );
XOR2_X1 U946 ( .A(G125), .B(n1236), .Z(G27) );
AND4_X1 U947 ( .A1(n1282), .A2(n1089), .A3(n1288), .A4(n1289), .ZN(n1236) );
NOR2_X1 U948 ( .A1(n1106), .A2(n1284), .ZN(n1288) );
INV_X1 U949 ( .A(n1243), .ZN(n1089) );
AND2_X1 U950 ( .A1(n1083), .A2(n1290), .ZN(n1282) );
NAND2_X1 U951 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
OR3_X1 U952 ( .A1(n1293), .A2(G900), .A3(n1103), .ZN(n1291) );
XOR2_X1 U953 ( .A(G122), .B(n1294), .Z(G24) );
NOR2_X1 U954 ( .A1(n1106), .A2(n1266), .ZN(n1294) );
NAND4_X1 U955 ( .A1(n1249), .A2(n1097), .A3(n1295), .A4(n1281), .ZN(n1266) );
NOR2_X1 U956 ( .A1(n1088), .A2(n1092), .ZN(n1097) );
INV_X1 U957 ( .A(n1111), .ZN(n1092) );
NOR2_X1 U958 ( .A1(n1287), .A2(n1286), .ZN(n1111) );
INV_X1 U959 ( .A(n1289), .ZN(n1088) );
XOR2_X1 U960 ( .A(n1256), .B(n1296), .Z(G21) );
NAND2_X1 U961 ( .A1(KEYINPUT36), .A2(G119), .ZN(n1296) );
NAND4_X1 U962 ( .A1(n1267), .A2(n1082), .A3(n1286), .A4(n1287), .ZN(n1256) );
INV_X1 U963 ( .A(n1297), .ZN(n1286) );
XOR2_X1 U964 ( .A(n1298), .B(n1299), .Z(G18) );
NAND4_X1 U965 ( .A1(KEYINPUT60), .A2(n1267), .A3(n1090), .A4(n1099), .ZN(n1299) );
NOR2_X1 U966 ( .A1(n1300), .A2(n1281), .ZN(n1099) );
XOR2_X1 U967 ( .A(n1260), .B(n1301), .Z(G15) );
NAND2_X1 U968 ( .A1(KEYINPUT16), .A2(G113), .ZN(n1301) );
NAND3_X1 U969 ( .A1(n1101), .A2(n1090), .A3(n1267), .ZN(n1260) );
AND3_X1 U970 ( .A1(n1295), .A2(n1245), .A3(n1289), .ZN(n1267) );
NOR2_X1 U971 ( .A1(n1302), .A2(n1095), .ZN(n1289) );
NOR2_X1 U972 ( .A1(n1287), .A2(n1297), .ZN(n1090) );
INV_X1 U973 ( .A(n1284), .ZN(n1101) );
NAND2_X1 U974 ( .A1(n1281), .A2(n1300), .ZN(n1284) );
INV_X1 U975 ( .A(n1249), .ZN(n1300) );
XOR2_X1 U976 ( .A(G110), .B(n1303), .Z(G12) );
NOR3_X1 U977 ( .A1(n1243), .A2(KEYINPUT51), .A3(n1264), .ZN(n1303) );
NAND2_X1 U978 ( .A1(n1082), .A2(n1261), .ZN(n1264) );
AND3_X1 U979 ( .A1(n1295), .A2(n1245), .A3(n1094), .ZN(n1261) );
NOR2_X1 U980 ( .A1(n1304), .A2(n1302), .ZN(n1094) );
XNOR2_X1 U981 ( .A(n1114), .B(KEYINPUT44), .ZN(n1302) );
INV_X1 U982 ( .A(n1096), .ZN(n1114) );
NAND2_X1 U983 ( .A1(G221), .A2(n1305), .ZN(n1096) );
INV_X1 U984 ( .A(n1095), .ZN(n1304) );
XOR2_X1 U985 ( .A(n1306), .B(G469), .Z(n1095) );
NAND2_X1 U986 ( .A1(KEYINPUT54), .A2(n1129), .ZN(n1306) );
NAND2_X1 U987 ( .A1(n1293), .A2(n1307), .ZN(n1129) );
NAND2_X1 U988 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
OR2_X1 U989 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U990 ( .A(n1312), .B(KEYINPUT28), .Z(n1308) );
NAND2_X1 U991 ( .A1(n1311), .A2(n1310), .ZN(n1312) );
XNOR2_X1 U992 ( .A(n1220), .B(n1313), .ZN(n1310) );
INV_X1 U993 ( .A(n1216), .ZN(n1313) );
XOR2_X1 U994 ( .A(n1205), .B(n1147), .Z(n1216) );
XNOR2_X1 U995 ( .A(n1206), .B(KEYINPUT47), .ZN(n1147) );
XOR2_X1 U996 ( .A(n1314), .B(n1315), .Z(n1220) );
XOR2_X1 U997 ( .A(KEYINPUT35), .B(G107), .Z(n1315) );
XNOR2_X1 U998 ( .A(G101), .B(G104), .ZN(n1314) );
XOR2_X1 U999 ( .A(n1316), .B(n1223), .Z(n1311) );
NAND2_X1 U1000 ( .A1(G227), .A2(n1103), .ZN(n1223) );
NAND2_X1 U1001 ( .A1(KEYINPUT12), .A2(n1224), .ZN(n1316) );
XOR2_X1 U1002 ( .A(G140), .B(G110), .Z(n1224) );
INV_X1 U1003 ( .A(n1106), .ZN(n1245) );
NAND2_X1 U1004 ( .A1(n1317), .A2(n1119), .ZN(n1106) );
NAND2_X1 U1005 ( .A1(G214), .A2(n1318), .ZN(n1119) );
XOR2_X1 U1006 ( .A(n1076), .B(KEYINPUT17), .Z(n1317) );
XOR2_X1 U1007 ( .A(n1117), .B(n1319), .Z(n1076) );
NOR2_X1 U1008 ( .A1(n1123), .A2(KEYINPUT42), .ZN(n1319) );
INV_X1 U1009 ( .A(n1127), .ZN(n1123) );
NAND2_X1 U1010 ( .A1(n1320), .A2(n1293), .ZN(n1127) );
XOR2_X1 U1011 ( .A(n1228), .B(n1321), .Z(n1320) );
XOR2_X1 U1012 ( .A(n1322), .B(n1323), .Z(n1321) );
NAND2_X1 U1013 ( .A1(KEYINPUT32), .A2(n1206), .ZN(n1322) );
XNOR2_X1 U1014 ( .A(n1324), .B(n1169), .ZN(n1228) );
XNOR2_X1 U1015 ( .A(n1168), .B(n1167), .ZN(n1169) );
XOR2_X1 U1016 ( .A(n1325), .B(n1326), .Z(n1167) );
NOR2_X1 U1017 ( .A1(KEYINPUT56), .A2(G110), .ZN(n1326) );
XOR2_X1 U1018 ( .A(n1327), .B(KEYINPUT50), .Z(n1325) );
INV_X1 U1019 ( .A(G122), .ZN(n1327) );
XNOR2_X1 U1020 ( .A(n1328), .B(n1329), .ZN(n1168) );
XOR2_X1 U1021 ( .A(KEYINPUT40), .B(n1330), .Z(n1329) );
NOR2_X1 U1022 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
XOR2_X1 U1023 ( .A(n1333), .B(KEYINPUT30), .Z(n1332) );
NAND2_X1 U1024 ( .A1(G104), .A2(n1334), .ZN(n1333) );
NOR2_X1 U1025 ( .A1(G104), .A2(n1334), .ZN(n1331) );
XOR2_X1 U1026 ( .A(n1335), .B(n1336), .Z(n1328) );
NOR2_X1 U1027 ( .A1(G116), .A2(KEYINPUT58), .ZN(n1336) );
NAND2_X1 U1028 ( .A1(G224), .A2(n1103), .ZN(n1324) );
NAND2_X1 U1029 ( .A1(G210), .A2(n1318), .ZN(n1117) );
NAND2_X1 U1030 ( .A1(n1337), .A2(n1293), .ZN(n1318) );
INV_X1 U1031 ( .A(G237), .ZN(n1337) );
AND2_X1 U1032 ( .A1(n1338), .A2(n1083), .ZN(n1295) );
NAND2_X1 U1033 ( .A1(G237), .A2(G234), .ZN(n1083) );
NAND2_X1 U1034 ( .A1(n1292), .A2(n1339), .ZN(n1338) );
NAND3_X1 U1035 ( .A1(G902), .A2(n1165), .A3(G953), .ZN(n1339) );
INV_X1 U1036 ( .A(G898), .ZN(n1165) );
NAND2_X1 U1037 ( .A1(n1340), .A2(n1103), .ZN(n1292) );
XOR2_X1 U1038 ( .A(KEYINPUT22), .B(G952), .Z(n1340) );
NOR2_X1 U1039 ( .A1(n1281), .A2(n1249), .ZN(n1082) );
XOR2_X1 U1040 ( .A(n1182), .B(n1341), .Z(n1249) );
NOR2_X1 U1041 ( .A1(n1132), .A2(KEYINPUT33), .ZN(n1341) );
NOR2_X1 U1042 ( .A1(n1183), .A2(G902), .ZN(n1132) );
XOR2_X1 U1043 ( .A(n1342), .B(n1343), .Z(n1183) );
XOR2_X1 U1044 ( .A(G116), .B(n1344), .Z(n1343) );
XOR2_X1 U1045 ( .A(G134), .B(G122), .Z(n1344) );
XOR2_X1 U1046 ( .A(n1345), .B(n1346), .Z(n1342) );
NOR2_X1 U1047 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
INV_X1 U1048 ( .A(G217), .ZN(n1347) );
XOR2_X1 U1049 ( .A(n1334), .B(n1349), .Z(n1345) );
NOR2_X1 U1050 ( .A1(KEYINPUT31), .A2(n1350), .ZN(n1349) );
INV_X1 U1051 ( .A(G107), .ZN(n1334) );
INV_X1 U1052 ( .A(G478), .ZN(n1182) );
XNOR2_X1 U1053 ( .A(n1118), .B(KEYINPUT37), .ZN(n1281) );
XOR2_X1 U1054 ( .A(n1351), .B(G475), .Z(n1118) );
NAND2_X1 U1055 ( .A1(n1293), .A2(n1189), .ZN(n1351) );
NAND2_X1 U1056 ( .A1(n1352), .A2(n1353), .ZN(n1189) );
NAND2_X1 U1057 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
XOR2_X1 U1058 ( .A(n1356), .B(KEYINPUT20), .Z(n1352) );
OR2_X1 U1059 ( .A1(n1355), .A2(n1354), .ZN(n1356) );
XNOR2_X1 U1060 ( .A(n1357), .B(n1358), .ZN(n1354) );
XOR2_X1 U1061 ( .A(KEYINPUT45), .B(G122), .Z(n1358) );
XNOR2_X1 U1062 ( .A(G113), .B(G104), .ZN(n1357) );
XNOR2_X1 U1063 ( .A(n1359), .B(n1360), .ZN(n1355) );
XOR2_X1 U1064 ( .A(n1361), .B(n1362), .Z(n1360) );
NAND2_X1 U1065 ( .A1(n1363), .A2(G214), .ZN(n1362) );
NAND3_X1 U1066 ( .A1(n1364), .A2(n1365), .A3(n1366), .ZN(n1361) );
NAND2_X1 U1067 ( .A1(KEYINPUT38), .A2(n1149), .ZN(n1366) );
NAND3_X1 U1068 ( .A1(n1367), .A2(n1368), .A3(n1268), .ZN(n1365) );
INV_X1 U1069 ( .A(KEYINPUT38), .ZN(n1368) );
OR2_X1 U1070 ( .A1(n1268), .A2(n1367), .ZN(n1364) );
NOR2_X1 U1071 ( .A1(n1369), .A2(n1149), .ZN(n1367) );
INV_X1 U1072 ( .A(KEYINPUT23), .ZN(n1369) );
XOR2_X1 U1073 ( .A(n1370), .B(G143), .Z(n1359) );
INV_X1 U1074 ( .A(G131), .ZN(n1370) );
NAND2_X1 U1075 ( .A1(n1297), .A2(n1287), .ZN(n1243) );
XOR2_X1 U1076 ( .A(n1371), .B(n1176), .Z(n1287) );
NAND2_X1 U1077 ( .A1(G217), .A2(n1305), .ZN(n1176) );
NAND2_X1 U1078 ( .A1(G234), .A2(n1293), .ZN(n1305) );
OR2_X1 U1079 ( .A1(n1175), .A2(G902), .ZN(n1371) );
XNOR2_X1 U1080 ( .A(n1372), .B(n1373), .ZN(n1175) );
XOR2_X1 U1081 ( .A(G110), .B(n1374), .Z(n1373) );
XOR2_X1 U1082 ( .A(G128), .B(G119), .Z(n1374) );
XNOR2_X1 U1083 ( .A(n1375), .B(n1376), .ZN(n1372) );
NOR2_X1 U1084 ( .A1(KEYINPUT46), .A2(n1377), .ZN(n1376) );
XOR2_X1 U1085 ( .A(n1149), .B(n1268), .Z(n1377) );
XOR2_X1 U1086 ( .A(G140), .B(n1230), .Z(n1149) );
INV_X1 U1087 ( .A(n1323), .ZN(n1230) );
XNOR2_X1 U1088 ( .A(G125), .B(KEYINPUT21), .ZN(n1323) );
NOR2_X1 U1089 ( .A1(KEYINPUT7), .A2(n1378), .ZN(n1375) );
XOR2_X1 U1090 ( .A(n1379), .B(KEYINPUT5), .Z(n1378) );
NAND3_X1 U1091 ( .A1(n1380), .A2(n1381), .A3(n1382), .ZN(n1379) );
OR2_X1 U1092 ( .A1(n1383), .A2(G137), .ZN(n1382) );
NAND2_X1 U1093 ( .A1(n1384), .A2(n1385), .ZN(n1381) );
INV_X1 U1094 ( .A(KEYINPUT1), .ZN(n1385) );
NAND2_X1 U1095 ( .A1(n1386), .A2(G137), .ZN(n1384) );
XNOR2_X1 U1096 ( .A(n1383), .B(KEYINPUT62), .ZN(n1386) );
NAND2_X1 U1097 ( .A1(KEYINPUT1), .A2(n1387), .ZN(n1380) );
NAND2_X1 U1098 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
OR2_X1 U1099 ( .A1(n1383), .A2(KEYINPUT62), .ZN(n1389) );
NAND3_X1 U1100 ( .A1(n1383), .A2(G137), .A3(KEYINPUT62), .ZN(n1388) );
NOR2_X1 U1101 ( .A1(n1348), .A2(n1390), .ZN(n1383) );
INV_X1 U1102 ( .A(G221), .ZN(n1390) );
NAND2_X1 U1103 ( .A1(G234), .A2(n1103), .ZN(n1348) );
INV_X1 U1104 ( .A(G953), .ZN(n1103) );
XOR2_X1 U1105 ( .A(n1391), .B(G472), .Z(n1297) );
NAND2_X1 U1106 ( .A1(n1392), .A2(n1293), .ZN(n1391) );
INV_X1 U1107 ( .A(G902), .ZN(n1293) );
XOR2_X1 U1108 ( .A(n1393), .B(n1394), .Z(n1392) );
XOR2_X1 U1109 ( .A(n1395), .B(n1396), .Z(n1394) );
INV_X1 U1110 ( .A(n1335), .ZN(n1396) );
XNOR2_X1 U1111 ( .A(G101), .B(n1196), .ZN(n1335) );
XOR2_X1 U1112 ( .A(G113), .B(G119), .Z(n1196) );
XOR2_X1 U1113 ( .A(n1205), .B(n1397), .Z(n1395) );
INV_X1 U1114 ( .A(n1197), .ZN(n1397) );
XOR2_X1 U1115 ( .A(n1298), .B(KEYINPUT27), .Z(n1197) );
INV_X1 U1116 ( .A(G116), .ZN(n1298) );
XOR2_X1 U1117 ( .A(n1150), .B(n1146), .Z(n1205) );
XOR2_X1 U1118 ( .A(G131), .B(G137), .Z(n1146) );
INV_X1 U1119 ( .A(G134), .ZN(n1150) );
XNOR2_X1 U1120 ( .A(n1398), .B(n1206), .ZN(n1393) );
XNOR2_X1 U1121 ( .A(n1399), .B(n1350), .ZN(n1206) );
XNOR2_X1 U1122 ( .A(G128), .B(G143), .ZN(n1350) );
XOR2_X1 U1123 ( .A(n1268), .B(KEYINPUT63), .Z(n1399) );
INV_X1 U1124 ( .A(G146), .ZN(n1268) );
XOR2_X1 U1125 ( .A(n1202), .B(KEYINPUT8), .Z(n1398) );
NAND2_X1 U1126 ( .A1(n1363), .A2(G210), .ZN(n1202) );
NOR2_X1 U1127 ( .A1(G953), .A2(G237), .ZN(n1363) );
endmodule


