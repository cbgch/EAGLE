//Key = 0111001101001000101011010101111010111110011101100010101011100010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303;

XNOR2_X1 U716 ( .A(G107), .B(n994), .ZN(G9) );
NOR2_X1 U717 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR4_X1 U718 ( .A1(n997), .A2(n998), .A3(G953), .A4(n999), .ZN(n996) );
NOR3_X1 U719 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n998) );
NOR2_X1 U720 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR2_X1 U721 ( .A1(KEYINPUT47), .A2(n1005), .ZN(n1003) );
NAND4_X1 U722 ( .A1(n1006), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n997) );
NAND3_X1 U723 ( .A1(KEYINPUT47), .A2(n1010), .A3(n1011), .ZN(n1009) );
NAND3_X1 U724 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
OR2_X1 U725 ( .A1(n1011), .A2(KEYINPUT47), .ZN(n1008) );
NAND2_X1 U726 ( .A1(n1015), .A2(n1016), .ZN(n1011) );
NAND2_X1 U727 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND3_X1 U728 ( .A1(n1012), .A2(n1019), .A3(n1020), .ZN(n1018) );
NAND2_X1 U729 ( .A1(n1021), .A2(n1022), .ZN(n1019) );
NAND2_X1 U730 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND2_X1 U731 ( .A1(n1014), .A2(n1025), .ZN(n1017) );
NAND2_X1 U732 ( .A1(n1015), .A2(n1026), .ZN(n1007) );
NAND2_X1 U733 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND4_X1 U734 ( .A1(n1029), .A2(n1020), .A3(n1030), .A4(n1031), .ZN(n1028) );
NAND2_X1 U735 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U736 ( .A1(n1012), .A2(n1034), .ZN(n1032) );
NAND2_X1 U737 ( .A1(n1035), .A2(n1036), .ZN(n1030) );
NAND2_X1 U738 ( .A1(n1023), .A2(n1037), .ZN(n1036) );
XOR2_X1 U739 ( .A(KEYINPUT13), .B(n1012), .Z(n1037) );
NAND3_X1 U740 ( .A1(n1014), .A2(n1038), .A3(n1039), .ZN(n1027) );
INV_X1 U741 ( .A(n1000), .ZN(n1014) );
NAND4_X1 U742 ( .A1(n1020), .A2(n1023), .A3(n1029), .A4(n1033), .ZN(n1000) );
INV_X1 U743 ( .A(n1040), .ZN(n1020) );
INV_X1 U744 ( .A(n1041), .ZN(n1006) );
NOR3_X1 U745 ( .A1(n999), .A2(G953), .A3(G952), .ZN(n995) );
AND4_X1 U746 ( .A1(n1033), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n999) );
NOR2_X1 U747 ( .A1(n1045), .A2(n1046), .ZN(n1044) );
XOR2_X1 U748 ( .A(n1047), .B(KEYINPUT53), .Z(n1045) );
NAND4_X1 U749 ( .A1(n1048), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1047) );
XOR2_X1 U750 ( .A(n1052), .B(n1053), .Z(n1051) );
XOR2_X1 U751 ( .A(n1054), .B(KEYINPUT31), .Z(n1053) );
NAND2_X1 U752 ( .A1(KEYINPUT58), .A2(n1055), .ZN(n1052) );
XOR2_X1 U753 ( .A(KEYINPUT45), .B(n1056), .Z(n1050) );
XOR2_X1 U754 ( .A(n1057), .B(KEYINPUT35), .Z(n1048) );
XOR2_X1 U755 ( .A(n1058), .B(n1059), .Z(n1043) );
NAND2_X1 U756 ( .A1(KEYINPUT46), .A2(n1060), .ZN(n1059) );
XOR2_X1 U757 ( .A(n1061), .B(n1062), .Z(G72) );
XOR2_X1 U758 ( .A(n1063), .B(n1064), .Z(n1062) );
NOR2_X1 U759 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
XOR2_X1 U760 ( .A(n1067), .B(n1068), .Z(n1066) );
XOR2_X1 U761 ( .A(n1069), .B(n1070), .Z(n1068) );
XOR2_X1 U762 ( .A(n1071), .B(n1072), .Z(n1067) );
XNOR2_X1 U763 ( .A(KEYINPUT10), .B(n1073), .ZN(n1072) );
NOR2_X1 U764 ( .A1(G900), .A2(n1074), .ZN(n1065) );
NAND2_X1 U765 ( .A1(n1074), .A2(n1075), .ZN(n1063) );
NAND2_X1 U766 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
XOR2_X1 U767 ( .A(n1078), .B(KEYINPUT11), .Z(n1076) );
NAND2_X1 U768 ( .A1(G953), .A2(n1079), .ZN(n1061) );
NAND2_X1 U769 ( .A1(G900), .A2(G227), .ZN(n1079) );
XOR2_X1 U770 ( .A(n1080), .B(n1081), .Z(G69) );
XOR2_X1 U771 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U772 ( .A1(n1084), .A2(n1074), .ZN(n1083) );
NOR2_X1 U773 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
XOR2_X1 U774 ( .A(KEYINPUT36), .B(G224), .Z(n1086) );
NAND2_X1 U775 ( .A1(n1087), .A2(n1088), .ZN(n1082) );
XOR2_X1 U776 ( .A(KEYINPUT54), .B(n1089), .Z(n1088) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(n1087) );
NAND3_X1 U778 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1090) );
NAND2_X1 U779 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NAND2_X1 U780 ( .A1(KEYINPUT14), .A2(n1097), .ZN(n1093) );
NAND2_X1 U781 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
XOR2_X1 U782 ( .A(KEYINPUT56), .B(n1096), .Z(n1099) );
NAND2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1092) );
INV_X1 U784 ( .A(KEYINPUT14), .ZN(n1101) );
NAND2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND3_X1 U786 ( .A1(KEYINPUT56), .A2(n1098), .A3(n1104), .ZN(n1103) );
OR2_X1 U787 ( .A1(n1104), .A2(KEYINPUT56), .ZN(n1102) );
NAND2_X1 U788 ( .A1(n1074), .A2(n1105), .ZN(n1080) );
NAND2_X1 U789 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XNOR2_X1 U790 ( .A(KEYINPUT3), .B(n1108), .ZN(n1107) );
NOR2_X1 U791 ( .A1(n1109), .A2(n1110), .ZN(G66) );
XOR2_X1 U792 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR3_X1 U793 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1111) );
XNOR2_X1 U794 ( .A(G217), .B(KEYINPUT8), .ZN(n1115) );
NOR2_X1 U795 ( .A1(n1109), .A2(n1116), .ZN(G63) );
XNOR2_X1 U796 ( .A(n1117), .B(n1118), .ZN(n1116) );
NOR2_X1 U797 ( .A1(n1055), .A2(n1113), .ZN(n1118) );
INV_X1 U798 ( .A(G478), .ZN(n1055) );
NOR2_X1 U799 ( .A1(n1109), .A2(n1119), .ZN(G60) );
XOR2_X1 U800 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U801 ( .A1(n1122), .A2(n1113), .ZN(n1120) );
INV_X1 U802 ( .A(G475), .ZN(n1122) );
XNOR2_X1 U803 ( .A(G104), .B(n1123), .ZN(G6) );
NAND2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
NOR2_X1 U805 ( .A1(n1126), .A2(n1127), .ZN(G57) );
XNOR2_X1 U806 ( .A(n1109), .B(KEYINPUT41), .ZN(n1127) );
XOR2_X1 U807 ( .A(n1128), .B(n1129), .Z(n1126) );
XOR2_X1 U808 ( .A(n1130), .B(n1131), .Z(n1129) );
XNOR2_X1 U809 ( .A(KEYINPUT24), .B(n1132), .ZN(n1131) );
NOR2_X1 U810 ( .A1(n1133), .A2(n1113), .ZN(n1130) );
INV_X1 U811 ( .A(G472), .ZN(n1133) );
XOR2_X1 U812 ( .A(n1134), .B(n1135), .Z(n1128) );
XOR2_X1 U813 ( .A(n1136), .B(n1137), .Z(n1134) );
NOR2_X1 U814 ( .A1(KEYINPUT49), .A2(n1138), .ZN(n1137) );
NOR2_X1 U815 ( .A1(n1109), .A2(n1139), .ZN(G54) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1139) );
XOR2_X1 U817 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U818 ( .A1(n1058), .A2(n1113), .ZN(n1142) );
INV_X1 U819 ( .A(G469), .ZN(n1058) );
XNOR2_X1 U820 ( .A(n1144), .B(n1145), .ZN(n1140) );
NOR2_X1 U821 ( .A1(KEYINPUT5), .A2(n1146), .ZN(n1145) );
XNOR2_X1 U822 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U823 ( .A(G140), .B(G110), .Z(n1148) );
NAND2_X1 U824 ( .A1(KEYINPUT32), .A2(n1149), .ZN(n1144) );
NOR2_X1 U825 ( .A1(n1109), .A2(n1150), .ZN(G51) );
XOR2_X1 U826 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U827 ( .A(n1153), .B(n1154), .ZN(n1152) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1151) );
NOR2_X1 U829 ( .A1(n1157), .A2(n1113), .ZN(n1156) );
NAND2_X1 U830 ( .A1(n1158), .A2(n1041), .ZN(n1113) );
NAND4_X1 U831 ( .A1(n1077), .A2(n1106), .A3(n1078), .A4(n1108), .ZN(n1041) );
AND4_X1 U832 ( .A1(n1159), .A2(n1160), .A3(n1161), .A4(n1162), .ZN(n1106) );
AND4_X1 U833 ( .A1(n994), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1162) );
NAND2_X1 U834 ( .A1(n1034), .A2(n1125), .ZN(n994) );
AND2_X1 U835 ( .A1(n1166), .A2(n1015), .ZN(n1125) );
NAND3_X1 U836 ( .A1(n1013), .A2(n1166), .A3(n1023), .ZN(n1161) );
NAND4_X1 U837 ( .A1(n1124), .A2(n1015), .A3(n1167), .A4(n1024), .ZN(n1159) );
NOR2_X1 U838 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
XOR2_X1 U839 ( .A(n1170), .B(KEYINPUT18), .Z(n1169) );
AND4_X1 U840 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1077) );
NOR4_X1 U841 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
INV_X1 U842 ( .A(n1179), .ZN(n1176) );
NAND4_X1 U843 ( .A1(n1180), .A2(n1004), .A3(n1025), .A4(n1181), .ZN(n1173) );
XOR2_X1 U844 ( .A(n1182), .B(KEYINPUT25), .Z(n1158) );
NOR2_X1 U845 ( .A1(n1074), .A2(G952), .ZN(n1109) );
XNOR2_X1 U846 ( .A(G146), .B(n1171), .ZN(G48) );
NAND3_X1 U847 ( .A1(n1183), .A2(n1025), .A3(n1124), .ZN(n1171) );
XOR2_X1 U848 ( .A(n1172), .B(n1184), .Z(G45) );
XNOR2_X1 U849 ( .A(G143), .B(KEYINPUT60), .ZN(n1184) );
NAND4_X1 U850 ( .A1(n1024), .A2(n1025), .A3(n1013), .A4(n1185), .ZN(n1172) );
AND3_X1 U851 ( .A1(n1186), .A2(n1181), .A3(n1187), .ZN(n1185) );
NAND2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(G42) );
OR2_X1 U853 ( .A1(n1190), .A2(G140), .ZN(n1189) );
NAND2_X1 U854 ( .A1(n1191), .A2(G140), .ZN(n1188) );
NAND2_X1 U855 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NAND2_X1 U856 ( .A1(n1178), .A2(n1194), .ZN(n1193) );
INV_X1 U857 ( .A(KEYINPUT1), .ZN(n1194) );
NAND2_X1 U858 ( .A1(KEYINPUT1), .A2(n1190), .ZN(n1192) );
NAND2_X1 U859 ( .A1(KEYINPUT57), .A2(n1178), .ZN(n1190) );
AND3_X1 U860 ( .A1(n1124), .A2(n1195), .A3(n1004), .ZN(n1178) );
XOR2_X1 U861 ( .A(G137), .B(n1177), .Z(G39) );
AND3_X1 U862 ( .A1(n1183), .A2(n1012), .A3(n1023), .ZN(n1177) );
XNOR2_X1 U863 ( .A(G134), .B(n1078), .ZN(G36) );
NAND3_X1 U864 ( .A1(n1013), .A2(n1034), .A3(n1195), .ZN(n1078) );
NAND3_X1 U865 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(G33) );
NAND2_X1 U866 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
INV_X1 U867 ( .A(G131), .ZN(n1200) );
NAND2_X1 U868 ( .A1(n1201), .A2(KEYINPUT38), .ZN(n1199) );
XOR2_X1 U869 ( .A(n1179), .B(KEYINPUT33), .Z(n1201) );
NAND3_X1 U870 ( .A1(KEYINPUT38), .A2(G131), .A3(n1179), .ZN(n1197) );
OR2_X1 U871 ( .A1(n1179), .A2(KEYINPUT38), .ZN(n1196) );
NAND3_X1 U872 ( .A1(n1195), .A2(n1013), .A3(n1124), .ZN(n1179) );
AND3_X1 U873 ( .A1(n1024), .A2(n1181), .A3(n1012), .ZN(n1195) );
INV_X1 U874 ( .A(n1002), .ZN(n1012) );
NAND2_X1 U875 ( .A1(n1038), .A2(n1042), .ZN(n1002) );
XOR2_X1 U876 ( .A(n1202), .B(n1203), .Z(G30) );
NAND2_X1 U877 ( .A1(KEYINPUT20), .A2(n1175), .ZN(n1203) );
AND3_X1 U878 ( .A1(n1034), .A2(n1025), .A3(n1183), .ZN(n1175) );
AND4_X1 U879 ( .A1(n1057), .A2(n1024), .A3(n1056), .A4(n1181), .ZN(n1183) );
XOR2_X1 U880 ( .A(G101), .B(n1204), .Z(G3) );
NOR4_X1 U881 ( .A1(KEYINPUT40), .A2(n1205), .A3(n1005), .A4(n1206), .ZN(n1204) );
XOR2_X1 U882 ( .A(G125), .B(n1207), .Z(G27) );
NOR4_X1 U883 ( .A1(n1208), .A2(n1209), .A3(n1021), .A4(n1210), .ZN(n1207) );
XNOR2_X1 U884 ( .A(KEYINPUT0), .B(n1181), .ZN(n1210) );
NAND2_X1 U885 ( .A1(n1040), .A2(n1211), .ZN(n1181) );
NAND4_X1 U886 ( .A1(G902), .A2(G953), .A3(n1212), .A4(n1213), .ZN(n1211) );
INV_X1 U887 ( .A(G900), .ZN(n1213) );
INV_X1 U888 ( .A(n1004), .ZN(n1209) );
XOR2_X1 U889 ( .A(n1214), .B(KEYINPUT22), .Z(n1208) );
XNOR2_X1 U890 ( .A(G122), .B(n1160), .ZN(G24) );
NAND4_X1 U891 ( .A1(n1215), .A2(n1015), .A3(n1186), .A4(n1187), .ZN(n1160) );
NOR2_X1 U892 ( .A1(n1056), .A2(n1057), .ZN(n1015) );
XOR2_X1 U893 ( .A(n1216), .B(G119), .Z(G21) );
NAND2_X1 U894 ( .A1(KEYINPUT7), .A2(n1165), .ZN(n1216) );
NAND4_X1 U895 ( .A1(n1023), .A2(n1215), .A3(n1057), .A4(n1056), .ZN(n1165) );
INV_X1 U896 ( .A(n1217), .ZN(n1056) );
XNOR2_X1 U897 ( .A(n1218), .B(n1108), .ZN(G18) );
NAND3_X1 U898 ( .A1(n1013), .A2(n1034), .A3(n1215), .ZN(n1108) );
NOR4_X1 U899 ( .A1(n1219), .A2(n1214), .A3(n1035), .A4(n1168), .ZN(n1215) );
INV_X1 U900 ( .A(n1220), .ZN(n1168) );
INV_X1 U901 ( .A(n1029), .ZN(n1219) );
AND2_X1 U902 ( .A1(n1049), .A2(n1186), .ZN(n1034) );
NAND2_X1 U903 ( .A1(KEYINPUT62), .A2(n1221), .ZN(n1218) );
INV_X1 U904 ( .A(G116), .ZN(n1221) );
XNOR2_X1 U905 ( .A(G113), .B(n1164), .ZN(G15) );
NAND4_X1 U906 ( .A1(n1180), .A2(n1013), .A3(n1170), .A4(n1220), .ZN(n1164) );
INV_X1 U907 ( .A(n1005), .ZN(n1013) );
NAND2_X1 U908 ( .A1(n1057), .A2(n1217), .ZN(n1005) );
INV_X1 U909 ( .A(n1021), .ZN(n1180) );
NAND3_X1 U910 ( .A1(n1029), .A2(n1033), .A3(n1124), .ZN(n1021) );
AND2_X1 U911 ( .A1(n1222), .A2(n1187), .ZN(n1124) );
XNOR2_X1 U912 ( .A(n1163), .B(n1223), .ZN(G12) );
XOR2_X1 U913 ( .A(KEYINPUT61), .B(G110), .Z(n1223) );
NAND3_X1 U914 ( .A1(n1023), .A2(n1166), .A3(n1004), .ZN(n1163) );
NOR2_X1 U915 ( .A1(n1057), .A2(n1217), .ZN(n1004) );
XOR2_X1 U916 ( .A(n1224), .B(n1225), .Z(n1217) );
NOR2_X1 U917 ( .A1(n1114), .A2(n1226), .ZN(n1225) );
XOR2_X1 U918 ( .A(KEYINPUT52), .B(G217), .Z(n1226) );
INV_X1 U919 ( .A(n1227), .ZN(n1114) );
OR2_X1 U920 ( .A1(n1112), .A2(G902), .ZN(n1224) );
XNOR2_X1 U921 ( .A(n1228), .B(n1229), .ZN(n1112) );
XOR2_X1 U922 ( .A(n1070), .B(n1230), .Z(n1229) );
XOR2_X1 U923 ( .A(n1231), .B(n1232), .Z(n1230) );
NAND2_X1 U924 ( .A1(n1233), .A2(KEYINPUT23), .ZN(n1232) );
XOR2_X1 U925 ( .A(n1234), .B(G137), .Z(n1233) );
NAND2_X1 U926 ( .A1(G221), .A2(n1235), .ZN(n1234) );
XOR2_X1 U927 ( .A(G125), .B(G140), .Z(n1070) );
XOR2_X1 U928 ( .A(n1236), .B(n1237), .Z(n1228) );
XOR2_X1 U929 ( .A(G146), .B(G128), .Z(n1237) );
INV_X1 U930 ( .A(G119), .ZN(n1236) );
XOR2_X1 U931 ( .A(n1238), .B(n1239), .Z(n1057) );
XOR2_X1 U932 ( .A(KEYINPUT43), .B(G472), .Z(n1239) );
NAND2_X1 U933 ( .A1(n1240), .A2(n1182), .ZN(n1238) );
XOR2_X1 U934 ( .A(n1241), .B(n1136), .Z(n1240) );
XOR2_X1 U935 ( .A(n1242), .B(G101), .Z(n1136) );
NAND3_X1 U936 ( .A1(G210), .A2(n1074), .A3(n1243), .ZN(n1242) );
XOR2_X1 U937 ( .A(n1244), .B(KEYINPUT48), .Z(n1243) );
NAND2_X1 U938 ( .A1(n1245), .A2(KEYINPUT6), .ZN(n1241) );
XOR2_X1 U939 ( .A(n1246), .B(n1138), .Z(n1245) );
XOR2_X1 U940 ( .A(n1135), .B(n1132), .Z(n1246) );
XNOR2_X1 U941 ( .A(n1104), .B(KEYINPUT29), .ZN(n1135) );
INV_X1 U942 ( .A(n1205), .ZN(n1166) );
NAND3_X1 U943 ( .A1(n1170), .A2(n1220), .A3(n1024), .ZN(n1205) );
NOR2_X1 U944 ( .A1(n1029), .A2(n1035), .ZN(n1024) );
INV_X1 U945 ( .A(n1033), .ZN(n1035) );
NAND2_X1 U946 ( .A1(G221), .A2(n1227), .ZN(n1033) );
NAND2_X1 U947 ( .A1(G234), .A2(n1182), .ZN(n1227) );
XOR2_X1 U948 ( .A(n1060), .B(n1247), .Z(n1029) );
XOR2_X1 U949 ( .A(KEYINPUT17), .B(G469), .Z(n1247) );
NAND2_X1 U950 ( .A1(n1248), .A2(n1182), .ZN(n1060) );
XNOR2_X1 U951 ( .A(n1143), .B(n1249), .ZN(n1248) );
XOR2_X1 U952 ( .A(n1250), .B(n1149), .Z(n1249) );
INV_X1 U953 ( .A(n1069), .ZN(n1149) );
XOR2_X1 U954 ( .A(n1251), .B(n1252), .Z(n1069) );
NAND2_X1 U955 ( .A1(KEYINPUT42), .A2(G128), .ZN(n1251) );
NOR2_X1 U956 ( .A1(KEYINPUT44), .A2(n1253), .ZN(n1250) );
NOR2_X1 U957 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
XOR2_X1 U958 ( .A(n1256), .B(KEYINPUT27), .Z(n1255) );
NAND2_X1 U959 ( .A1(n1147), .A2(n1257), .ZN(n1256) );
NOR2_X1 U960 ( .A1(n1147), .A2(n1257), .ZN(n1254) );
XOR2_X1 U961 ( .A(n1258), .B(n1231), .Z(n1257) );
INV_X1 U962 ( .A(G110), .ZN(n1231) );
NAND2_X1 U963 ( .A1(KEYINPUT34), .A2(n1259), .ZN(n1258) );
AND2_X1 U964 ( .A1(G227), .A2(n1074), .ZN(n1147) );
XNOR2_X1 U965 ( .A(n1132), .B(n1260), .ZN(n1143) );
XOR2_X1 U966 ( .A(G101), .B(n1261), .Z(n1260) );
NOR2_X1 U967 ( .A1(KEYINPUT39), .A2(n1262), .ZN(n1261) );
XNOR2_X1 U968 ( .A(n1263), .B(KEYINPUT30), .ZN(n1262) );
NAND2_X1 U969 ( .A1(n1264), .A2(n1265), .ZN(n1132) );
NAND2_X1 U970 ( .A1(n1071), .A2(n1073), .ZN(n1265) );
XOR2_X1 U971 ( .A(KEYINPUT9), .B(n1266), .Z(n1264) );
NOR2_X1 U972 ( .A1(n1071), .A2(n1073), .ZN(n1266) );
XNOR2_X1 U973 ( .A(G131), .B(KEYINPUT4), .ZN(n1073) );
XNOR2_X1 U974 ( .A(G134), .B(G137), .ZN(n1071) );
NAND2_X1 U975 ( .A1(n1040), .A2(n1267), .ZN(n1220) );
NAND3_X1 U976 ( .A1(n1089), .A2(n1212), .A3(G902), .ZN(n1267) );
AND2_X1 U977 ( .A1(n1268), .A2(G953), .ZN(n1089) );
XOR2_X1 U978 ( .A(n1085), .B(KEYINPUT19), .Z(n1268) );
INV_X1 U979 ( .A(G898), .ZN(n1085) );
NAND3_X1 U980 ( .A1(n1212), .A2(n1074), .A3(G952), .ZN(n1040) );
NAND2_X1 U981 ( .A1(G237), .A2(G234), .ZN(n1212) );
XOR2_X1 U982 ( .A(n1214), .B(KEYINPUT12), .Z(n1170) );
INV_X1 U983 ( .A(n1025), .ZN(n1214) );
NOR2_X1 U984 ( .A1(n1038), .A2(n1039), .ZN(n1025) );
INV_X1 U985 ( .A(n1042), .ZN(n1039) );
NAND2_X1 U986 ( .A1(G214), .A2(n1269), .ZN(n1042) );
XOR2_X1 U987 ( .A(n1046), .B(KEYINPUT37), .Z(n1038) );
XOR2_X1 U988 ( .A(n1270), .B(n1157), .Z(n1046) );
NAND2_X1 U989 ( .A1(G210), .A2(n1269), .ZN(n1157) );
NAND2_X1 U990 ( .A1(n1244), .A2(n1182), .ZN(n1269) );
NAND2_X1 U991 ( .A1(n1271), .A2(n1182), .ZN(n1270) );
XOR2_X1 U992 ( .A(n1272), .B(n1273), .Z(n1271) );
XOR2_X1 U993 ( .A(n1274), .B(n1155), .Z(n1273) );
AND2_X1 U994 ( .A1(G224), .A2(n1074), .ZN(n1155) );
NOR2_X1 U995 ( .A1(KEYINPUT26), .A2(n1153), .ZN(n1274) );
XOR2_X1 U996 ( .A(n1275), .B(n1098), .Z(n1153) );
INV_X1 U997 ( .A(n1095), .ZN(n1098) );
XOR2_X1 U998 ( .A(G101), .B(n1263), .Z(n1095) );
XOR2_X1 U999 ( .A(G104), .B(G107), .Z(n1263) );
XNOR2_X1 U1000 ( .A(n1091), .B(n1276), .ZN(n1275) );
NOR2_X1 U1001 ( .A1(KEYINPUT59), .A2(n1096), .ZN(n1276) );
INV_X1 U1002 ( .A(n1104), .ZN(n1096) );
XNOR2_X1 U1003 ( .A(G113), .B(n1277), .ZN(n1104) );
XOR2_X1 U1004 ( .A(G119), .B(G116), .Z(n1277) );
XNOR2_X1 U1005 ( .A(n1278), .B(G110), .ZN(n1091) );
NAND2_X1 U1006 ( .A1(KEYINPUT28), .A2(G122), .ZN(n1278) );
NOR2_X1 U1007 ( .A1(KEYINPUT15), .A2(n1154), .ZN(n1272) );
XNOR2_X1 U1008 ( .A(G125), .B(n1138), .ZN(n1154) );
XNOR2_X1 U1009 ( .A(n1279), .B(n1252), .ZN(n1138) );
XOR2_X1 U1010 ( .A(G143), .B(G146), .Z(n1252) );
XOR2_X1 U1011 ( .A(n1202), .B(KEYINPUT55), .Z(n1279) );
INV_X1 U1012 ( .A(G128), .ZN(n1202) );
INV_X1 U1013 ( .A(n1206), .ZN(n1023) );
NAND2_X1 U1014 ( .A1(n1280), .A2(n1222), .ZN(n1206) );
XNOR2_X1 U1015 ( .A(n1186), .B(KEYINPUT51), .ZN(n1222) );
XOR2_X1 U1016 ( .A(n1281), .B(G478), .Z(n1186) );
NAND2_X1 U1017 ( .A1(KEYINPUT21), .A2(n1054), .ZN(n1281) );
NAND2_X1 U1018 ( .A1(n1117), .A2(n1182), .ZN(n1054) );
INV_X1 U1019 ( .A(G902), .ZN(n1182) );
XNOR2_X1 U1020 ( .A(n1282), .B(n1283), .ZN(n1117) );
XOR2_X1 U1021 ( .A(n1284), .B(n1285), .Z(n1283) );
XOR2_X1 U1022 ( .A(G128), .B(G122), .Z(n1285) );
XOR2_X1 U1023 ( .A(G143), .B(G134), .Z(n1284) );
XOR2_X1 U1024 ( .A(n1286), .B(n1287), .Z(n1282) );
XOR2_X1 U1025 ( .A(G116), .B(G107), .Z(n1287) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1235), .ZN(n1286) );
AND2_X1 U1027 ( .A1(G234), .A2(n1074), .ZN(n1235) );
XOR2_X1 U1028 ( .A(KEYINPUT50), .B(n1187), .Z(n1280) );
INV_X1 U1029 ( .A(n1049), .ZN(n1187) );
XOR2_X1 U1030 ( .A(n1288), .B(G475), .Z(n1049) );
OR2_X1 U1031 ( .A1(n1121), .A2(G902), .ZN(n1288) );
XNOR2_X1 U1032 ( .A(n1289), .B(n1290), .ZN(n1121) );
XNOR2_X1 U1033 ( .A(G104), .B(n1291), .ZN(n1290) );
NAND3_X1 U1034 ( .A1(n1292), .A2(n1293), .A3(n1294), .ZN(n1291) );
OR2_X1 U1035 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND3_X1 U1036 ( .A1(n1296), .A2(n1295), .A3(KEYINPUT2), .ZN(n1293) );
XNOR2_X1 U1037 ( .A(n1297), .B(n1298), .ZN(n1295) );
XOR2_X1 U1038 ( .A(G143), .B(G131), .Z(n1298) );
NAND3_X1 U1039 ( .A1(n1244), .A2(n1074), .A3(G214), .ZN(n1297) );
INV_X1 U1040 ( .A(G953), .ZN(n1074) );
INV_X1 U1041 ( .A(G237), .ZN(n1244) );
AND2_X1 U1042 ( .A1(KEYINPUT16), .A2(n1299), .ZN(n1296) );
OR2_X1 U1043 ( .A1(n1299), .A2(KEYINPUT2), .ZN(n1292) );
XNOR2_X1 U1044 ( .A(n1300), .B(G146), .ZN(n1299) );
NAND2_X1 U1045 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1046 ( .A1(G125), .A2(n1259), .ZN(n1302) );
XOR2_X1 U1047 ( .A(n1303), .B(KEYINPUT63), .Z(n1301) );
OR2_X1 U1048 ( .A1(n1259), .A2(G125), .ZN(n1303) );
INV_X1 U1049 ( .A(G140), .ZN(n1259) );
XNOR2_X1 U1050 ( .A(G113), .B(G122), .ZN(n1289) );
endmodule


