//Key = 0000011110111011100101001011000001111110100101011001101000011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295;

XOR2_X1 U710 ( .A(n986), .B(n987), .Z(G9) );
NAND4_X1 U711 ( .A1(n988), .A2(n989), .A3(n990), .A4(n991), .ZN(n987) );
NOR2_X1 U712 ( .A1(KEYINPUT31), .A2(n992), .ZN(n990) );
NAND3_X1 U713 ( .A1(n993), .A2(n994), .A3(n995), .ZN(G75) );
NAND2_X1 U714 ( .A1(G952), .A2(n996), .ZN(n995) );
NAND3_X1 U715 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n996) );
XOR2_X1 U716 ( .A(n1000), .B(KEYINPUT23), .Z(n999) );
NAND4_X1 U717 ( .A1(n989), .A2(n1001), .A3(n1002), .A4(n1003), .ZN(n1000) );
NOR2_X1 U718 ( .A1(n1004), .A2(n1005), .ZN(n1003) );
NAND2_X1 U719 ( .A1(n1001), .A2(n1006), .ZN(n998) );
NAND2_X1 U720 ( .A1(n1007), .A2(n1008), .ZN(n1006) );
NAND3_X1 U721 ( .A1(n989), .A2(n1009), .A3(n1010), .ZN(n1008) );
NAND3_X1 U722 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1009) );
NAND2_X1 U723 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NAND3_X1 U724 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1012) );
XOR2_X1 U725 ( .A(n1004), .B(KEYINPUT19), .Z(n1018) );
XOR2_X1 U726 ( .A(n1019), .B(KEYINPUT10), .Z(n1016) );
NAND2_X1 U727 ( .A1(n1002), .A2(n1020), .ZN(n1011) );
NAND2_X1 U728 ( .A1(n1021), .A2(n1022), .ZN(n1020) );
NAND2_X1 U729 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NAND3_X1 U730 ( .A1(n1002), .A2(n1025), .A3(n1014), .ZN(n1007) );
NAND2_X1 U731 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NAND2_X1 U732 ( .A1(n1028), .A2(n1010), .ZN(n1027) );
INV_X1 U733 ( .A(n1029), .ZN(n1026) );
XNOR2_X1 U734 ( .A(n1030), .B(KEYINPUT54), .ZN(n1001) );
NAND4_X1 U735 ( .A1(n1031), .A2(n1032), .A3(n1033), .A4(n1034), .ZN(n993) );
NOR4_X1 U736 ( .A1(n1023), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1034) );
XOR2_X1 U737 ( .A(n1038), .B(n1039), .Z(n1037) );
NOR2_X1 U738 ( .A1(n1040), .A2(KEYINPUT63), .ZN(n1039) );
XNOR2_X1 U739 ( .A(n1041), .B(n1042), .ZN(n1036) );
NAND2_X1 U740 ( .A1(KEYINPUT36), .A2(n1043), .ZN(n1041) );
INV_X1 U741 ( .A(G472), .ZN(n1043) );
NOR2_X1 U742 ( .A1(n1044), .A2(n1045), .ZN(n1033) );
XOR2_X1 U743 ( .A(n1046), .B(n1047), .Z(n1045) );
NAND2_X1 U744 ( .A1(KEYINPUT7), .A2(G475), .ZN(n1047) );
XOR2_X1 U745 ( .A(n1048), .B(n1049), .Z(n1032) );
XOR2_X1 U746 ( .A(n1050), .B(KEYINPUT24), .Z(n1049) );
XOR2_X1 U747 ( .A(n1051), .B(n1052), .Z(G72) );
NOR2_X1 U748 ( .A1(n1053), .A2(n994), .ZN(n1052) );
NOR2_X1 U749 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NAND2_X1 U750 ( .A1(n1056), .A2(n1057), .ZN(n1051) );
NAND2_X1 U751 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
XOR2_X1 U752 ( .A(n1060), .B(n1061), .Z(n1056) );
NOR2_X1 U753 ( .A1(n1058), .A2(n1059), .ZN(n1061) );
INV_X1 U754 ( .A(KEYINPUT62), .ZN(n1059) );
NAND2_X1 U755 ( .A1(n1062), .A2(n1063), .ZN(n1058) );
NAND2_X1 U756 ( .A1(G953), .A2(n1064), .ZN(n1063) );
XOR2_X1 U757 ( .A(KEYINPUT33), .B(G900), .Z(n1064) );
XOR2_X1 U758 ( .A(n1065), .B(n1066), .Z(n1062) );
XOR2_X1 U759 ( .A(n1067), .B(n1068), .Z(n1066) );
NAND2_X1 U760 ( .A1(n1069), .A2(KEYINPUT16), .ZN(n1067) );
XOR2_X1 U761 ( .A(n1070), .B(n1071), .Z(n1069) );
XOR2_X1 U762 ( .A(KEYINPUT43), .B(G140), .Z(n1071) );
NAND2_X1 U763 ( .A1(KEYINPUT15), .A2(n1072), .ZN(n1070) );
XOR2_X1 U764 ( .A(KEYINPUT5), .B(G125), .Z(n1072) );
XOR2_X1 U765 ( .A(KEYINPUT59), .B(n1073), .Z(n1065) );
NOR2_X1 U766 ( .A1(KEYINPUT53), .A2(n1074), .ZN(n1073) );
XOR2_X1 U767 ( .A(n1075), .B(G131), .Z(n1074) );
NAND2_X1 U768 ( .A1(KEYINPUT11), .A2(n1076), .ZN(n1075) );
XOR2_X1 U769 ( .A(G134), .B(n1077), .Z(n1076) );
NOR2_X1 U770 ( .A1(G137), .A2(KEYINPUT9), .ZN(n1077) );
NAND2_X1 U771 ( .A1(n994), .A2(n1078), .ZN(n1060) );
XOR2_X1 U772 ( .A(n1079), .B(n1080), .Z(G69) );
NOR2_X1 U773 ( .A1(n1081), .A2(n994), .ZN(n1080) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
NAND3_X1 U776 ( .A1(n1086), .A2(n1087), .A3(n1088), .ZN(n1085) );
NAND2_X1 U777 ( .A1(G953), .A2(n1083), .ZN(n1087) );
INV_X1 U778 ( .A(G898), .ZN(n1083) );
OR2_X1 U779 ( .A1(n1086), .A2(n1088), .ZN(n1084) );
NAND2_X1 U780 ( .A1(n994), .A2(n1089), .ZN(n1088) );
NAND4_X1 U781 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n1094), .ZN(n1090) );
XNOR2_X1 U783 ( .A(n1095), .B(n1096), .ZN(n1086) );
XOR2_X1 U784 ( .A(KEYINPUT14), .B(n1097), .Z(n1096) );
NOR2_X1 U785 ( .A1(n1098), .A2(n1099), .ZN(G66) );
XOR2_X1 U786 ( .A(n1100), .B(n1101), .Z(n1099) );
NAND2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NOR2_X1 U788 ( .A1(n1098), .A2(n1104), .ZN(G63) );
XOR2_X1 U789 ( .A(n1105), .B(n1106), .Z(n1104) );
NAND2_X1 U790 ( .A1(n1102), .A2(G478), .ZN(n1105) );
NOR2_X1 U791 ( .A1(n1098), .A2(n1107), .ZN(G60) );
XOR2_X1 U792 ( .A(n1108), .B(n1109), .Z(n1107) );
NAND2_X1 U793 ( .A1(n1102), .A2(G475), .ZN(n1108) );
XNOR2_X1 U794 ( .A(G104), .B(n1110), .ZN(G6) );
NOR2_X1 U795 ( .A1(n1098), .A2(n1111), .ZN(G57) );
XOR2_X1 U796 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U797 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND2_X1 U798 ( .A1(n1102), .A2(G472), .ZN(n1115) );
NAND2_X1 U799 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
XOR2_X1 U800 ( .A(KEYINPUT45), .B(KEYINPUT0), .Z(n1117) );
XOR2_X1 U801 ( .A(n1118), .B(KEYINPUT55), .Z(n1116) );
XOR2_X1 U802 ( .A(n1119), .B(n1120), .Z(n1112) );
NOR2_X1 U803 ( .A1(n1098), .A2(n1121), .ZN(G54) );
XOR2_X1 U804 ( .A(n1122), .B(n1123), .Z(n1121) );
XOR2_X1 U805 ( .A(KEYINPUT3), .B(n1124), .Z(n1123) );
NOR2_X1 U806 ( .A1(KEYINPUT58), .A2(n1125), .ZN(n1124) );
XOR2_X1 U807 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U808 ( .A1(n1128), .A2(KEYINPUT27), .ZN(n1126) );
XNOR2_X1 U809 ( .A(n1129), .B(KEYINPUT4), .ZN(n1128) );
NAND2_X1 U810 ( .A1(n1102), .A2(G469), .ZN(n1122) );
NOR2_X1 U811 ( .A1(n1098), .A2(n1130), .ZN(G51) );
XOR2_X1 U812 ( .A(n1131), .B(n1132), .Z(n1130) );
NAND2_X1 U813 ( .A1(n1102), .A2(n1133), .ZN(n1131) );
INV_X1 U814 ( .A(n1048), .ZN(n1133) );
NOR2_X1 U815 ( .A1(n1134), .A2(n997), .ZN(n1102) );
AND4_X1 U816 ( .A1(n1092), .A2(n1093), .A3(n1091), .A4(n1135), .ZN(n997) );
NOR2_X1 U817 ( .A1(n1094), .A2(n1078), .ZN(n1135) );
NAND4_X1 U818 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1078) );
NOR4_X1 U819 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
NOR2_X1 U820 ( .A1(n1005), .A2(n1144), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1021), .A2(n1145), .ZN(n1142) );
INV_X1 U822 ( .A(n1146), .ZN(n1140) );
AND2_X1 U823 ( .A1(n1147), .A2(n1148), .ZN(n1138) );
NAND3_X1 U824 ( .A1(n1110), .A2(n1149), .A3(n1150), .ZN(n1094) );
NAND3_X1 U825 ( .A1(n1151), .A2(n1029), .A3(n991), .ZN(n1150) );
NAND2_X1 U826 ( .A1(n1152), .A2(n1153), .ZN(n1029) );
NAND3_X1 U827 ( .A1(n1154), .A2(n1155), .A3(n1010), .ZN(n1153) );
NAND2_X1 U828 ( .A1(n988), .A2(n989), .ZN(n1152) );
NAND4_X1 U829 ( .A1(n1156), .A2(n989), .A3(n1151), .A4(n991), .ZN(n1110) );
NAND2_X1 U830 ( .A1(n1157), .A2(n1158), .ZN(n1091) );
NAND2_X1 U831 ( .A1(n1159), .A2(n1005), .ZN(n1158) );
XNOR2_X1 U832 ( .A(n988), .B(KEYINPUT17), .ZN(n1159) );
NOR2_X1 U833 ( .A1(n994), .A2(G952), .ZN(n1098) );
XOR2_X1 U834 ( .A(G146), .B(n1141), .Z(G48) );
AND3_X1 U835 ( .A1(n1015), .A2(n1160), .A3(n1161), .ZN(n1141) );
XNOR2_X1 U836 ( .A(G143), .B(n1147), .ZN(G45) );
NAND4_X1 U837 ( .A1(n1162), .A2(n1044), .A3(n1163), .A4(n1164), .ZN(n1147) );
AND3_X1 U838 ( .A1(n1165), .A2(n1015), .A3(n1028), .ZN(n1164) );
XNOR2_X1 U839 ( .A(G140), .B(n1136), .ZN(G42) );
NAND3_X1 U840 ( .A1(n1154), .A2(n1166), .A3(n1156), .ZN(n1136) );
XNOR2_X1 U841 ( .A(G137), .B(n1137), .ZN(G39) );
NAND3_X1 U842 ( .A1(n1010), .A2(n1160), .A3(n1166), .ZN(n1137) );
AND4_X1 U843 ( .A1(n1165), .A2(n1014), .A3(n1015), .A4(n1155), .ZN(n1166) );
NAND2_X1 U844 ( .A1(n1167), .A2(n1168), .ZN(G36) );
OR2_X1 U845 ( .A1(n1148), .A2(G134), .ZN(n1168) );
XOR2_X1 U846 ( .A(n1169), .B(KEYINPUT20), .Z(n1167) );
NAND2_X1 U847 ( .A1(G134), .A2(n1148), .ZN(n1169) );
NAND2_X1 U848 ( .A1(n1170), .A2(n988), .ZN(n1148) );
INV_X1 U849 ( .A(n1144), .ZN(n1170) );
XOR2_X1 U850 ( .A(G131), .B(n1171), .Z(G33) );
NOR2_X1 U851 ( .A1(n1144), .A2(n1172), .ZN(n1171) );
XOR2_X1 U852 ( .A(KEYINPUT60), .B(n1156), .Z(n1172) );
INV_X1 U853 ( .A(n1005), .ZN(n1156) );
NAND4_X1 U854 ( .A1(n1165), .A2(n1014), .A3(n1028), .A4(n1015), .ZN(n1144) );
INV_X1 U855 ( .A(n1004), .ZN(n1014) );
NAND2_X1 U856 ( .A1(n1024), .A2(n1173), .ZN(n1004) );
XNOR2_X1 U857 ( .A(G128), .B(n1174), .ZN(G30) );
NAND2_X1 U858 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
INV_X1 U859 ( .A(n1145), .ZN(n1176) );
NAND4_X1 U860 ( .A1(n1165), .A2(n988), .A3(n1177), .A4(n1151), .ZN(n1145) );
NOR2_X1 U861 ( .A1(n1154), .A2(n1031), .ZN(n1177) );
INV_X1 U862 ( .A(n1178), .ZN(n1165) );
XOR2_X1 U863 ( .A(n1021), .B(KEYINPUT38), .Z(n1175) );
XNOR2_X1 U864 ( .A(G101), .B(n1149), .ZN(G3) );
NAND3_X1 U865 ( .A1(n1151), .A2(n1179), .A3(n1028), .ZN(n1149) );
NAND2_X1 U866 ( .A1(n1180), .A2(n1181), .ZN(G27) );
NAND2_X1 U867 ( .A1(n1182), .A2(n1146), .ZN(n1181) );
XOR2_X1 U868 ( .A(n1183), .B(KEYINPUT22), .Z(n1180) );
OR2_X1 U869 ( .A1(n1146), .A2(n1182), .ZN(n1183) );
XNOR2_X1 U870 ( .A(n1184), .B(KEYINPUT39), .ZN(n1182) );
NAND3_X1 U871 ( .A1(n1154), .A2(n1002), .A3(n1161), .ZN(n1146) );
NOR4_X1 U872 ( .A1(n1005), .A2(n1178), .A3(n1021), .A4(n1031), .ZN(n1161) );
INV_X1 U873 ( .A(n1163), .ZN(n1021) );
NAND2_X1 U874 ( .A1(n1185), .A2(n1186), .ZN(n1178) );
NAND2_X1 U875 ( .A1(n1187), .A2(G953), .ZN(n1186) );
XOR2_X1 U876 ( .A(n1055), .B(KEYINPUT33), .Z(n1187) );
INV_X1 U877 ( .A(G900), .ZN(n1055) );
XOR2_X1 U878 ( .A(n1188), .B(n1092), .Z(G24) );
NAND4_X1 U879 ( .A1(n1002), .A2(n989), .A3(n1189), .A4(n991), .ZN(n1092) );
AND2_X1 U880 ( .A1(n1044), .A2(n1162), .ZN(n1189) );
NOR2_X1 U881 ( .A1(n1160), .A2(n1155), .ZN(n989) );
XNOR2_X1 U882 ( .A(n1190), .B(n1093), .ZN(G21) );
NAND4_X1 U883 ( .A1(n1179), .A2(n1002), .A3(n1155), .A4(n1160), .ZN(n1093) );
NAND2_X1 U884 ( .A1(KEYINPUT47), .A2(n1191), .ZN(n1190) );
NAND2_X1 U885 ( .A1(n1192), .A2(n1193), .ZN(G18) );
NAND2_X1 U886 ( .A1(G116), .A2(n1194), .ZN(n1193) );
XOR2_X1 U887 ( .A(KEYINPUT35), .B(n1195), .Z(n1192) );
NOR2_X1 U888 ( .A1(G116), .A2(n1194), .ZN(n1195) );
NAND2_X1 U889 ( .A1(n1157), .A2(n988), .ZN(n1194) );
NOR2_X1 U890 ( .A1(n1162), .A2(n1196), .ZN(n988) );
INV_X1 U891 ( .A(n1197), .ZN(n1157) );
XOR2_X1 U892 ( .A(G113), .B(n1198), .Z(G15) );
NOR2_X1 U893 ( .A1(n1197), .A2(n1005), .ZN(n1198) );
NAND2_X1 U894 ( .A1(n1196), .A2(n1162), .ZN(n1005) );
NAND3_X1 U895 ( .A1(n1002), .A2(n991), .A3(n1028), .ZN(n1197) );
NOR2_X1 U896 ( .A1(n1155), .A2(n1154), .ZN(n1028) );
INV_X1 U897 ( .A(n1031), .ZN(n1155) );
AND2_X1 U898 ( .A1(n1017), .A2(n1019), .ZN(n1002) );
XNOR2_X1 U899 ( .A(G110), .B(n1199), .ZN(G12) );
NAND3_X1 U900 ( .A1(KEYINPUT51), .A2(n1179), .A3(n1200), .ZN(n1199) );
NOR3_X1 U901 ( .A1(n992), .A2(n1031), .A3(n1160), .ZN(n1200) );
INV_X1 U902 ( .A(n1154), .ZN(n1160) );
XOR2_X1 U903 ( .A(n1042), .B(G472), .Z(n1154) );
NAND2_X1 U904 ( .A1(n1201), .A2(n1134), .ZN(n1042) );
XOR2_X1 U905 ( .A(n1118), .B(n1202), .Z(n1201) );
XNOR2_X1 U906 ( .A(KEYINPUT49), .B(n1203), .ZN(n1202) );
NOR2_X1 U907 ( .A1(KEYINPUT25), .A2(n1204), .ZN(n1203) );
XOR2_X1 U908 ( .A(n1205), .B(n1120), .Z(n1204) );
XNOR2_X1 U909 ( .A(n1206), .B(G113), .ZN(n1120) );
NAND2_X1 U910 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U911 ( .A1(G119), .A2(n1209), .ZN(n1208) );
INV_X1 U912 ( .A(G116), .ZN(n1209) );
XOR2_X1 U913 ( .A(n1210), .B(KEYINPUT42), .Z(n1207) );
NAND2_X1 U914 ( .A1(G116), .A2(n1191), .ZN(n1210) );
NAND2_X1 U915 ( .A1(KEYINPUT48), .A2(n1119), .ZN(n1205) );
XNOR2_X1 U916 ( .A(n1211), .B(n1212), .ZN(n1118) );
NAND2_X1 U917 ( .A1(G210), .A2(n1213), .ZN(n1211) );
XOR2_X1 U918 ( .A(n1214), .B(n1103), .Z(n1031) );
AND2_X1 U919 ( .A1(G217), .A2(n1215), .ZN(n1103) );
NAND2_X1 U920 ( .A1(n1101), .A2(n1134), .ZN(n1214) );
XNOR2_X1 U921 ( .A(n1216), .B(n1217), .ZN(n1101) );
XOR2_X1 U922 ( .A(n1218), .B(n1219), .Z(n1217) );
XNOR2_X1 U923 ( .A(n1129), .B(n1220), .ZN(n1219) );
AND4_X1 U924 ( .A1(n1221), .A2(n994), .A3(n1222), .A4(G221), .ZN(n1220) );
INV_X1 U925 ( .A(KEYINPUT13), .ZN(n1221) );
XOR2_X1 U926 ( .A(n1191), .B(n1223), .Z(n1216) );
XOR2_X1 U927 ( .A(G137), .B(G128), .Z(n1223) );
INV_X1 U928 ( .A(n1151), .ZN(n992) );
XNOR2_X1 U929 ( .A(n1015), .B(KEYINPUT8), .ZN(n1151) );
NOR2_X1 U930 ( .A1(n1017), .A2(n1035), .ZN(n1015) );
INV_X1 U931 ( .A(n1019), .ZN(n1035) );
NAND2_X1 U932 ( .A1(G221), .A2(n1215), .ZN(n1019) );
NAND2_X1 U933 ( .A1(G234), .A2(n1134), .ZN(n1215) );
XNOR2_X1 U934 ( .A(n1224), .B(n1040), .ZN(n1017) );
AND2_X1 U935 ( .A1(n1225), .A2(n1134), .ZN(n1040) );
XNOR2_X1 U936 ( .A(n1127), .B(n1129), .ZN(n1225) );
XOR2_X1 U937 ( .A(G110), .B(G140), .Z(n1129) );
XNOR2_X1 U938 ( .A(n1226), .B(n1227), .ZN(n1127) );
XOR2_X1 U939 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U940 ( .A(KEYINPUT59), .B(n1230), .Z(n1229) );
NOR2_X1 U941 ( .A1(KEYINPUT50), .A2(n1231), .ZN(n1230) );
NOR2_X1 U942 ( .A1(G953), .A2(n1054), .ZN(n1228) );
INV_X1 U943 ( .A(G227), .ZN(n1054) );
XNOR2_X1 U944 ( .A(n1119), .B(n1212), .ZN(n1226) );
XOR2_X1 U945 ( .A(n1232), .B(n1233), .Z(n1119) );
XNOR2_X1 U946 ( .A(G137), .B(n1234), .ZN(n1233) );
XNOR2_X1 U947 ( .A(KEYINPUT52), .B(KEYINPUT32), .ZN(n1234) );
XOR2_X1 U948 ( .A(n1235), .B(n1236), .Z(n1232) );
INV_X1 U949 ( .A(n1068), .ZN(n1236) );
XOR2_X1 U950 ( .A(n1237), .B(n1238), .Z(n1235) );
NOR2_X1 U951 ( .A1(G131), .A2(KEYINPUT29), .ZN(n1238) );
INV_X1 U952 ( .A(G134), .ZN(n1237) );
NAND2_X1 U953 ( .A1(KEYINPUT21), .A2(n1038), .ZN(n1224) );
INV_X1 U954 ( .A(G469), .ZN(n1038) );
AND2_X1 U955 ( .A1(n1010), .A2(n991), .ZN(n1179) );
AND3_X1 U956 ( .A1(n1185), .A2(n1239), .A3(n1163), .ZN(n991) );
NOR2_X1 U957 ( .A1(n1024), .A2(n1023), .ZN(n1163) );
INV_X1 U958 ( .A(n1173), .ZN(n1023) );
NAND2_X1 U959 ( .A1(G214), .A2(n1240), .ZN(n1173) );
XOR2_X1 U960 ( .A(n1241), .B(n1050), .Z(n1024) );
NAND2_X1 U961 ( .A1(n1242), .A2(n1134), .ZN(n1050) );
XOR2_X1 U962 ( .A(KEYINPUT2), .B(n1132), .Z(n1242) );
XNOR2_X1 U963 ( .A(n1243), .B(n1244), .ZN(n1132) );
XOR2_X1 U964 ( .A(n1245), .B(n1068), .Z(n1244) );
XOR2_X1 U965 ( .A(n1246), .B(n1247), .Z(n1068) );
XNOR2_X1 U966 ( .A(G146), .B(KEYINPUT46), .ZN(n1246) );
NAND3_X1 U967 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1245) );
NAND2_X1 U968 ( .A1(n1095), .A2(n1251), .ZN(n1250) );
NAND2_X1 U969 ( .A1(KEYINPUT34), .A2(n1252), .ZN(n1251) );
XOR2_X1 U970 ( .A(KEYINPUT1), .B(n1097), .Z(n1252) );
INV_X1 U971 ( .A(n1253), .ZN(n1095) );
NAND3_X1 U972 ( .A1(KEYINPUT44), .A2(n1254), .A3(n1255), .ZN(n1249) );
INV_X1 U973 ( .A(n1097), .ZN(n1255) );
NAND2_X1 U974 ( .A1(KEYINPUT1), .A2(n1256), .ZN(n1254) );
NAND3_X1 U975 ( .A1(n1257), .A2(n1258), .A3(n1097), .ZN(n1248) );
XOR2_X1 U976 ( .A(G110), .B(G122), .Z(n1097) );
INV_X1 U977 ( .A(KEYINPUT44), .ZN(n1258) );
NAND2_X1 U978 ( .A1(n1259), .A2(n1256), .ZN(n1257) );
NAND2_X1 U979 ( .A1(n1253), .A2(KEYINPUT34), .ZN(n1256) );
XOR2_X1 U980 ( .A(n1260), .B(n1261), .Z(n1253) );
XOR2_X1 U981 ( .A(G113), .B(n1262), .Z(n1261) );
NOR2_X1 U982 ( .A1(n1263), .A2(n1264), .ZN(n1262) );
XOR2_X1 U983 ( .A(n1265), .B(KEYINPUT37), .Z(n1264) );
NAND2_X1 U984 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
XOR2_X1 U985 ( .A(KEYINPUT6), .B(G119), .Z(n1266) );
NOR2_X1 U986 ( .A1(n1191), .A2(n1267), .ZN(n1263) );
XOR2_X1 U987 ( .A(KEYINPUT41), .B(G116), .Z(n1267) );
INV_X1 U988 ( .A(G119), .ZN(n1191) );
XNOR2_X1 U989 ( .A(n1212), .B(n1231), .ZN(n1260) );
XNOR2_X1 U990 ( .A(G104), .B(G107), .ZN(n1231) );
XNOR2_X1 U991 ( .A(G101), .B(KEYINPUT30), .ZN(n1212) );
INV_X1 U992 ( .A(KEYINPUT1), .ZN(n1259) );
XOR2_X1 U993 ( .A(n1184), .B(n1268), .Z(n1243) );
NOR2_X1 U994 ( .A1(G953), .A2(n1082), .ZN(n1268) );
INV_X1 U995 ( .A(G224), .ZN(n1082) );
NAND2_X1 U996 ( .A1(KEYINPUT12), .A2(n1048), .ZN(n1241) );
NAND2_X1 U997 ( .A1(G210), .A2(n1240), .ZN(n1048) );
NAND2_X1 U998 ( .A1(n1269), .A2(n1134), .ZN(n1240) );
INV_X1 U999 ( .A(G237), .ZN(n1269) );
NAND2_X1 U1000 ( .A1(G898), .A2(G953), .ZN(n1239) );
AND3_X1 U1001 ( .A1(n1270), .A2(n1271), .A3(n1030), .ZN(n1185) );
NAND2_X1 U1002 ( .A1(G237), .A2(G234), .ZN(n1030) );
OR2_X1 U1003 ( .A1(G952), .A2(G953), .ZN(n1271) );
NAND2_X1 U1004 ( .A1(G953), .A2(n1134), .ZN(n1270) );
NOR2_X1 U1005 ( .A1(n1044), .A2(n1162), .ZN(n1010) );
XNOR2_X1 U1006 ( .A(n1046), .B(G475), .ZN(n1162) );
NAND2_X1 U1007 ( .A1(n1109), .A2(n1134), .ZN(n1046) );
XOR2_X1 U1008 ( .A(n1272), .B(n1273), .Z(n1109) );
XOR2_X1 U1009 ( .A(G113), .B(n1274), .Z(n1273) );
XOR2_X1 U1010 ( .A(KEYINPUT57), .B(G122), .Z(n1274) );
XOR2_X1 U1011 ( .A(n1275), .B(G104), .Z(n1272) );
NAND2_X1 U1012 ( .A1(n1276), .A2(KEYINPUT40), .ZN(n1275) );
XOR2_X1 U1013 ( .A(n1218), .B(n1277), .Z(n1276) );
XOR2_X1 U1014 ( .A(G140), .B(n1278), .Z(n1277) );
NOR2_X1 U1015 ( .A1(KEYINPUT18), .A2(n1279), .ZN(n1278) );
XOR2_X1 U1016 ( .A(n1280), .B(n1281), .Z(n1279) );
XOR2_X1 U1017 ( .A(G143), .B(G131), .Z(n1281) );
NAND2_X1 U1018 ( .A1(G214), .A2(n1213), .ZN(n1280) );
NOR2_X1 U1019 ( .A1(G953), .A2(G237), .ZN(n1213) );
XOR2_X1 U1020 ( .A(G146), .B(n1184), .Z(n1218) );
INV_X1 U1021 ( .A(G125), .ZN(n1184) );
INV_X1 U1022 ( .A(n1196), .ZN(n1044) );
XOR2_X1 U1023 ( .A(n1282), .B(G478), .Z(n1196) );
NAND2_X1 U1024 ( .A1(n1106), .A2(n1134), .ZN(n1282) );
INV_X1 U1025 ( .A(G902), .ZN(n1134) );
XOR2_X1 U1026 ( .A(n1283), .B(n1284), .Z(n1106) );
XNOR2_X1 U1027 ( .A(n1285), .B(n1247), .ZN(n1284) );
XOR2_X1 U1028 ( .A(G128), .B(G143), .Z(n1247) );
NAND2_X1 U1029 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
NAND2_X1 U1030 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U1031 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
NAND2_X1 U1032 ( .A1(KEYINPUT26), .A2(G107), .ZN(n1291) );
INV_X1 U1033 ( .A(n1292), .ZN(n1288) );
NAND2_X1 U1034 ( .A1(n1293), .A2(n986), .ZN(n1286) );
INV_X1 U1035 ( .A(G107), .ZN(n986) );
NAND2_X1 U1036 ( .A1(KEYINPUT26), .A2(n1294), .ZN(n1293) );
NAND2_X1 U1037 ( .A1(n1292), .A2(n1290), .ZN(n1294) );
INV_X1 U1038 ( .A(KEYINPUT56), .ZN(n1290) );
XNOR2_X1 U1039 ( .A(n1188), .B(G116), .ZN(n1292) );
INV_X1 U1040 ( .A(G122), .ZN(n1188) );
XOR2_X1 U1041 ( .A(n1295), .B(G134), .Z(n1283) );
NAND3_X1 U1042 ( .A1(n1222), .A2(n994), .A3(G217), .ZN(n1295) );
INV_X1 U1043 ( .A(G953), .ZN(n994) );
XOR2_X1 U1044 ( .A(G234), .B(KEYINPUT28), .Z(n1222) );
endmodule


