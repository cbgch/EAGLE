//Key = 0110100001101001110100110100001101011100010001101000011011101001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
n1388, n1389;

NAND3_X1 U760 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(G9) );
OR2_X1 U761 ( .A1(n1051), .A2(KEYINPUT45), .ZN(n1050) );
NAND3_X1 U762 ( .A1(KEYINPUT45), .A2(n1051), .A3(G107), .ZN(n1049) );
NAND2_X1 U763 ( .A1(n1052), .A2(n1053), .ZN(n1048) );
INV_X1 U764 ( .A(G107), .ZN(n1053) );
NAND2_X1 U765 ( .A1(n1054), .A2(KEYINPUT45), .ZN(n1052) );
XOR2_X1 U766 ( .A(n1051), .B(KEYINPUT20), .Z(n1054) );
NOR2_X1 U767 ( .A1(n1055), .A2(n1056), .ZN(G75) );
NOR4_X1 U768 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR2_X1 U769 ( .A1(KEYINPUT10), .A2(n1061), .ZN(n1059) );
AND3_X1 U770 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NAND4_X1 U771 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1057) );
NAND2_X1 U772 ( .A1(n1069), .A2(n1070), .ZN(n1066) );
NAND2_X1 U773 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NAND3_X1 U774 ( .A1(n1064), .A2(n1073), .A3(n1074), .ZN(n1072) );
NAND2_X1 U775 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NAND2_X1 U776 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
OR2_X1 U777 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U778 ( .A1(n1081), .A2(n1082), .ZN(n1075) );
NAND2_X1 U779 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NAND2_X1 U780 ( .A1(KEYINPUT10), .A2(n1063), .ZN(n1084) );
NAND2_X1 U781 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND3_X1 U782 ( .A1(n1077), .A2(n1087), .A3(n1081), .ZN(n1071) );
NAND3_X1 U783 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
NAND2_X1 U784 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XNOR2_X1 U785 ( .A(n1074), .B(KEYINPUT46), .ZN(n1091) );
OR3_X1 U786 ( .A1(n1093), .A2(KEYINPUT39), .A3(n1094), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1064), .A2(n1095), .ZN(n1088) );
NAND2_X1 U788 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
NAND2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
INV_X1 U790 ( .A(n1100), .ZN(n1069) );
NAND2_X1 U791 ( .A1(KEYINPUT39), .A2(n1101), .ZN(n1065) );
NAND2_X1 U792 ( .A1(n1062), .A2(n1102), .ZN(n1101) );
NOR3_X1 U793 ( .A1(n1093), .A2(n1103), .A3(n1100), .ZN(n1062) );
INV_X1 U794 ( .A(n1081), .ZN(n1103) );
NOR3_X1 U795 ( .A1(n1104), .A2(G953), .A3(G952), .ZN(n1055) );
INV_X1 U796 ( .A(n1067), .ZN(n1104) );
NAND4_X1 U797 ( .A1(n1105), .A2(n1106), .A3(n1107), .A4(n1108), .ZN(n1067) );
NOR4_X1 U798 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1108) );
XNOR2_X1 U799 ( .A(n1113), .B(n1114), .ZN(n1112) );
NAND2_X1 U800 ( .A1(n1115), .A2(KEYINPUT4), .ZN(n1113) );
XOR2_X1 U801 ( .A(G475), .B(n1116), .Z(n1111) );
NOR2_X1 U802 ( .A1(G902), .A2(n1117), .ZN(n1116) );
NOR3_X1 U803 ( .A1(n1118), .A2(n1119), .A3(n1098), .ZN(n1107) );
INV_X1 U804 ( .A(n1120), .ZN(n1119) );
NOR2_X1 U805 ( .A1(KEYINPUT4), .A2(n1115), .ZN(n1118) );
XNOR2_X1 U806 ( .A(KEYINPUT12), .B(G472), .ZN(n1115) );
OR2_X1 U807 ( .A1(n1121), .A2(n1122), .ZN(n1106) );
XOR2_X1 U808 ( .A(KEYINPUT37), .B(n1123), .Z(n1105) );
XOR2_X1 U809 ( .A(n1124), .B(n1125), .Z(G72) );
NOR2_X1 U810 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
XOR2_X1 U811 ( .A(n1128), .B(KEYINPUT17), .Z(n1127) );
NAND3_X1 U812 ( .A1(n1060), .A2(n1068), .A3(n1129), .ZN(n1128) );
XNOR2_X1 U813 ( .A(KEYINPUT16), .B(n1130), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1131), .A2(n1130), .ZN(n1126) );
NAND3_X1 U815 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1130) );
XOR2_X1 U816 ( .A(n1135), .B(KEYINPUT38), .Z(n1134) );
NAND2_X1 U817 ( .A1(n1136), .A2(n1137), .ZN(n1135) );
OR2_X1 U818 ( .A1(n1137), .A2(n1136), .ZN(n1133) );
XNOR2_X1 U819 ( .A(n1138), .B(n1139), .ZN(n1137) );
XOR2_X1 U820 ( .A(G134), .B(n1140), .Z(n1139) );
NOR2_X1 U821 ( .A1(KEYINPUT29), .A2(n1141), .ZN(n1140) );
XNOR2_X1 U822 ( .A(n1142), .B(n1143), .ZN(n1138) );
NOR2_X1 U823 ( .A1(G131), .A2(KEYINPUT49), .ZN(n1143) );
NOR2_X1 U824 ( .A1(G137), .A2(KEYINPUT14), .ZN(n1142) );
NAND2_X1 U825 ( .A1(G953), .A2(n1144), .ZN(n1132) );
AND2_X1 U826 ( .A1(n1068), .A2(n1060), .ZN(n1131) );
NAND2_X1 U827 ( .A1(G953), .A2(n1145), .ZN(n1124) );
NAND2_X1 U828 ( .A1(G900), .A2(G227), .ZN(n1145) );
XOR2_X1 U829 ( .A(n1146), .B(n1147), .Z(G69) );
XOR2_X1 U830 ( .A(n1148), .B(n1149), .Z(n1147) );
NOR2_X1 U831 ( .A1(n1150), .A2(n1068), .ZN(n1149) );
NOR2_X1 U832 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND2_X1 U833 ( .A1(n1153), .A2(n1154), .ZN(n1148) );
NAND2_X1 U834 ( .A1(G953), .A2(n1152), .ZN(n1154) );
XNOR2_X1 U835 ( .A(n1155), .B(n1156), .ZN(n1153) );
NAND2_X1 U836 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
NAND2_X1 U837 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
XOR2_X1 U838 ( .A(KEYINPUT53), .B(n1161), .Z(n1157) );
NOR2_X1 U839 ( .A1(n1159), .A2(n1160), .ZN(n1161) );
NAND2_X1 U840 ( .A1(n1068), .A2(n1058), .ZN(n1146) );
NOR2_X1 U841 ( .A1(n1162), .A2(n1163), .ZN(G66) );
XOR2_X1 U842 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U843 ( .A1(n1166), .A2(G217), .ZN(n1164) );
NOR2_X1 U844 ( .A1(n1162), .A2(n1167), .ZN(G63) );
XOR2_X1 U845 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U846 ( .A1(n1166), .A2(G478), .ZN(n1168) );
NOR2_X1 U847 ( .A1(n1162), .A2(n1170), .ZN(G60) );
XNOR2_X1 U848 ( .A(n1171), .B(n1117), .ZN(n1170) );
NAND2_X1 U849 ( .A1(n1166), .A2(G475), .ZN(n1171) );
XNOR2_X1 U850 ( .A(n1172), .B(n1173), .ZN(G6) );
NOR2_X1 U851 ( .A1(KEYINPUT0), .A2(n1174), .ZN(n1173) );
INV_X1 U852 ( .A(G104), .ZN(n1174) );
NOR2_X1 U853 ( .A1(n1162), .A2(n1175), .ZN(G57) );
XOR2_X1 U854 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U855 ( .A(n1178), .B(n1179), .Z(n1176) );
NOR2_X1 U856 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
XOR2_X1 U857 ( .A(n1182), .B(KEYINPUT36), .Z(n1181) );
INV_X1 U858 ( .A(n1183), .ZN(n1180) );
NAND2_X1 U859 ( .A1(n1166), .A2(G472), .ZN(n1178) );
NOR2_X1 U860 ( .A1(n1162), .A2(n1184), .ZN(G54) );
XOR2_X1 U861 ( .A(n1185), .B(n1186), .Z(n1184) );
XNOR2_X1 U862 ( .A(n1187), .B(n1188), .ZN(n1186) );
NAND4_X1 U863 ( .A1(KEYINPUT15), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187) );
NAND3_X1 U864 ( .A1(KEYINPUT57), .A2(n1192), .A3(n1193), .ZN(n1191) );
INV_X1 U865 ( .A(n1194), .ZN(n1192) );
NAND2_X1 U866 ( .A1(n1195), .A2(n1194), .ZN(n1190) );
NAND2_X1 U867 ( .A1(KEYINPUT63), .A2(n1196), .ZN(n1194) );
OR2_X1 U868 ( .A1(n1196), .A2(KEYINPUT57), .ZN(n1189) );
XOR2_X1 U869 ( .A(n1197), .B(n1198), .Z(n1196) );
XOR2_X1 U870 ( .A(n1141), .B(KEYINPUT31), .Z(n1197) );
XOR2_X1 U871 ( .A(n1199), .B(n1200), .Z(n1185) );
NOR3_X1 U872 ( .A1(n1201), .A2(KEYINPUT27), .A3(n1202), .ZN(n1200) );
NOR2_X1 U873 ( .A1(n1162), .A2(n1203), .ZN(G51) );
XOR2_X1 U874 ( .A(n1204), .B(n1205), .Z(n1203) );
XOR2_X1 U875 ( .A(n1206), .B(n1207), .Z(n1205) );
NAND2_X1 U876 ( .A1(n1166), .A2(n1122), .ZN(n1207) );
INV_X1 U877 ( .A(n1201), .ZN(n1166) );
NAND2_X1 U878 ( .A1(G902), .A2(n1208), .ZN(n1201) );
OR2_X1 U879 ( .A1(n1058), .A2(n1060), .ZN(n1208) );
NAND4_X1 U880 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1060) );
NOR4_X1 U881 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n1212) );
INV_X1 U882 ( .A(n1217), .ZN(n1216) );
NAND2_X1 U883 ( .A1(n1074), .A2(n1218), .ZN(n1211) );
NAND2_X1 U884 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND3_X1 U885 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1220) );
OR2_X1 U886 ( .A1(n1224), .A2(KEYINPUT50), .ZN(n1222) );
NAND2_X1 U887 ( .A1(KEYINPUT50), .A2(n1225), .ZN(n1221) );
NAND3_X1 U888 ( .A1(n1063), .A2(n1100), .A3(n1226), .ZN(n1225) );
XNOR2_X1 U889 ( .A(KEYINPUT60), .B(n1227), .ZN(n1219) );
NAND4_X1 U890 ( .A1(n1172), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1058) );
AND4_X1 U891 ( .A1(n1051), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1230) );
NAND3_X1 U892 ( .A1(n1064), .A2(n1234), .A3(n1080), .ZN(n1051) );
NAND3_X1 U893 ( .A1(n1234), .A2(n1235), .A3(n1081), .ZN(n1229) );
NAND2_X1 U894 ( .A1(n1094), .A2(n1236), .ZN(n1235) );
NAND3_X1 U895 ( .A1(n1064), .A2(n1234), .A3(n1079), .ZN(n1172) );
NAND2_X1 U896 ( .A1(n1237), .A2(KEYINPUT22), .ZN(n1206) );
XOR2_X1 U897 ( .A(n1238), .B(n1239), .Z(n1237) );
NAND2_X1 U898 ( .A1(n1240), .A2(n1241), .ZN(n1238) );
NAND2_X1 U899 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
XOR2_X1 U900 ( .A(KEYINPUT48), .B(n1244), .Z(n1240) );
NOR2_X1 U901 ( .A1(n1243), .A2(n1242), .ZN(n1244) );
NOR2_X1 U902 ( .A1(n1068), .A2(G952), .ZN(n1162) );
XNOR2_X1 U903 ( .A(G146), .B(n1209), .ZN(G48) );
NAND2_X1 U904 ( .A1(n1245), .A2(n1079), .ZN(n1209) );
NAND2_X1 U905 ( .A1(n1246), .A2(n1247), .ZN(G45) );
NAND2_X1 U906 ( .A1(G143), .A2(n1210), .ZN(n1247) );
XOR2_X1 U907 ( .A(n1248), .B(KEYINPUT59), .Z(n1246) );
OR2_X1 U908 ( .A1(n1210), .A2(G143), .ZN(n1248) );
NAND3_X1 U909 ( .A1(n1224), .A2(n1092), .A3(n1249), .ZN(n1210) );
NOR3_X1 U910 ( .A1(n1250), .A2(n1096), .A3(n1251), .ZN(n1249) );
INV_X1 U911 ( .A(n1252), .ZN(n1096) );
XOR2_X1 U912 ( .A(G140), .B(n1253), .Z(G42) );
NOR2_X1 U913 ( .A1(n1093), .A2(n1227), .ZN(n1253) );
NAND3_X1 U914 ( .A1(n1224), .A2(n1079), .A3(n1254), .ZN(n1227) );
NAND2_X1 U915 ( .A1(n1255), .A2(n1256), .ZN(G39) );
NAND2_X1 U916 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U917 ( .A1(G137), .A2(n1259), .ZN(n1258) );
NAND2_X1 U918 ( .A1(KEYINPUT62), .A2(KEYINPUT35), .ZN(n1259) );
INV_X1 U919 ( .A(n1260), .ZN(n1257) );
NAND3_X1 U920 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1255) );
INV_X1 U921 ( .A(KEYINPUT62), .ZN(n1263) );
NAND2_X1 U922 ( .A1(G137), .A2(n1264), .ZN(n1262) );
INV_X1 U923 ( .A(KEYINPUT35), .ZN(n1264) );
NAND2_X1 U924 ( .A1(KEYINPUT35), .A2(n1265), .ZN(n1261) );
NAND2_X1 U925 ( .A1(G137), .A2(n1260), .ZN(n1265) );
NAND2_X1 U926 ( .A1(n1074), .A2(n1266), .ZN(n1260) );
XOR2_X1 U927 ( .A(KEYINPUT5), .B(n1267), .Z(n1266) );
NOR2_X1 U928 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND2_X1 U929 ( .A1(n1270), .A2(n1271), .ZN(G36) );
NAND2_X1 U930 ( .A1(G134), .A2(n1272), .ZN(n1271) );
NAND2_X1 U931 ( .A1(n1215), .A2(n1273), .ZN(n1272) );
NAND2_X1 U932 ( .A1(KEYINPUT7), .A2(n1274), .ZN(n1273) );
NAND3_X1 U933 ( .A1(n1275), .A2(n1276), .A3(n1277), .ZN(n1270) );
INV_X1 U934 ( .A(KEYINPUT7), .ZN(n1277) );
NAND2_X1 U935 ( .A1(n1278), .A2(n1274), .ZN(n1276) );
INV_X1 U936 ( .A(KEYINPUT3), .ZN(n1274) );
NAND2_X1 U937 ( .A1(n1215), .A2(n1279), .ZN(n1275) );
OR2_X1 U938 ( .A1(G134), .A2(KEYINPUT3), .ZN(n1279) );
INV_X1 U939 ( .A(n1278), .ZN(n1215) );
NAND2_X1 U940 ( .A1(n1280), .A2(n1080), .ZN(n1278) );
XOR2_X1 U941 ( .A(G131), .B(n1214), .Z(G33) );
AND2_X1 U942 ( .A1(n1280), .A2(n1079), .ZN(n1214) );
NOR3_X1 U943 ( .A1(n1269), .A2(n1236), .A3(n1093), .ZN(n1280) );
INV_X1 U944 ( .A(n1074), .ZN(n1093) );
NOR2_X1 U945 ( .A1(n1281), .A2(n1098), .ZN(n1074) );
XNOR2_X1 U946 ( .A(n1282), .B(n1213), .ZN(G30) );
AND2_X1 U947 ( .A1(n1245), .A2(n1080), .ZN(n1213) );
AND4_X1 U948 ( .A1(n1283), .A2(n1224), .A3(n1252), .A4(n1109), .ZN(n1245) );
INV_X1 U949 ( .A(n1269), .ZN(n1224) );
NAND2_X1 U950 ( .A1(n1063), .A2(n1284), .ZN(n1269) );
XNOR2_X1 U951 ( .A(G101), .B(n1285), .ZN(G3) );
NAND3_X1 U952 ( .A1(n1092), .A2(n1234), .A3(n1286), .ZN(n1285) );
XNOR2_X1 U953 ( .A(n1081), .B(KEYINPUT58), .ZN(n1286) );
XNOR2_X1 U954 ( .A(G125), .B(n1217), .ZN(G27) );
NAND4_X1 U955 ( .A1(n1102), .A2(n1079), .A3(n1252), .A4(n1284), .ZN(n1217) );
NAND2_X1 U956 ( .A1(n1226), .A2(n1100), .ZN(n1284) );
XOR2_X1 U957 ( .A(n1287), .B(KEYINPUT11), .Z(n1226) );
NAND4_X1 U958 ( .A1(G953), .A2(n1288), .A3(n1289), .A4(n1144), .ZN(n1287) );
INV_X1 U959 ( .A(G900), .ZN(n1144) );
XNOR2_X1 U960 ( .A(KEYINPUT28), .B(n1290), .ZN(n1288) );
NOR2_X1 U961 ( .A1(n1094), .A2(n1110), .ZN(n1102) );
XNOR2_X1 U962 ( .A(G122), .B(n1228), .ZN(G24) );
NAND4_X1 U963 ( .A1(n1291), .A2(n1292), .A3(n1293), .A4(n1064), .ZN(n1228) );
NOR2_X1 U964 ( .A1(n1109), .A2(n1283), .ZN(n1064) );
XNOR2_X1 U965 ( .A(G119), .B(n1233), .ZN(G21) );
NAND2_X1 U966 ( .A1(n1223), .A2(n1292), .ZN(n1233) );
INV_X1 U967 ( .A(n1268), .ZN(n1223) );
NAND3_X1 U968 ( .A1(n1283), .A2(n1109), .A3(n1081), .ZN(n1268) );
NAND2_X1 U969 ( .A1(n1294), .A2(n1295), .ZN(G18) );
NAND2_X1 U970 ( .A1(G116), .A2(n1232), .ZN(n1295) );
XOR2_X1 U971 ( .A(n1296), .B(KEYINPUT61), .Z(n1294) );
OR2_X1 U972 ( .A1(n1232), .A2(G116), .ZN(n1296) );
NAND3_X1 U973 ( .A1(n1092), .A2(n1080), .A3(n1292), .ZN(n1232) );
NOR2_X1 U974 ( .A1(n1251), .A2(n1291), .ZN(n1080) );
XNOR2_X1 U975 ( .A(G113), .B(n1231), .ZN(G15) );
NAND3_X1 U976 ( .A1(n1079), .A2(n1092), .A3(n1292), .ZN(n1231) );
AND3_X1 U977 ( .A1(n1252), .A2(n1297), .A3(n1077), .ZN(n1292) );
INV_X1 U978 ( .A(n1110), .ZN(n1077) );
NAND2_X1 U979 ( .A1(n1086), .A2(n1298), .ZN(n1110) );
INV_X1 U980 ( .A(n1236), .ZN(n1092) );
NAND2_X1 U981 ( .A1(n1283), .A2(n1299), .ZN(n1236) );
NOR2_X1 U982 ( .A1(n1250), .A2(n1293), .ZN(n1079) );
XOR2_X1 U983 ( .A(n1300), .B(n1301), .Z(G12) );
NAND2_X1 U984 ( .A1(KEYINPUT23), .A2(G110), .ZN(n1301) );
NAND3_X1 U985 ( .A1(n1234), .A2(n1302), .A3(n1081), .ZN(n1300) );
NOR2_X1 U986 ( .A1(n1293), .A2(n1291), .ZN(n1081) );
INV_X1 U987 ( .A(n1250), .ZN(n1291) );
XNOR2_X1 U988 ( .A(n1303), .B(G475), .ZN(n1250) );
NAND2_X1 U989 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
NAND2_X1 U990 ( .A1(n1306), .A2(n1290), .ZN(n1305) );
INV_X1 U991 ( .A(n1117), .ZN(n1306) );
XNOR2_X1 U992 ( .A(n1307), .B(n1308), .ZN(n1117) );
XOR2_X1 U993 ( .A(n1136), .B(n1309), .Z(n1308) );
XNOR2_X1 U994 ( .A(n1310), .B(n1311), .ZN(n1309) );
XOR2_X1 U995 ( .A(n1312), .B(n1313), .Z(n1307) );
NOR2_X1 U996 ( .A1(KEYINPUT13), .A2(n1314), .ZN(n1313) );
XOR2_X1 U997 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U998 ( .A(n1317), .B(G131), .ZN(n1316) );
NAND4_X1 U999 ( .A1(KEYINPUT54), .A2(G214), .A3(n1318), .A4(n1068), .ZN(n1315) );
XNOR2_X1 U1000 ( .A(G113), .B(G122), .ZN(n1312) );
XNOR2_X1 U1001 ( .A(KEYINPUT52), .B(KEYINPUT47), .ZN(n1304) );
INV_X1 U1002 ( .A(n1251), .ZN(n1293) );
XOR2_X1 U1003 ( .A(n1123), .B(KEYINPUT30), .Z(n1251) );
XNOR2_X1 U1004 ( .A(n1319), .B(G478), .ZN(n1123) );
NAND2_X1 U1005 ( .A1(n1169), .A2(n1290), .ZN(n1319) );
XOR2_X1 U1006 ( .A(n1320), .B(n1321), .Z(n1169) );
NOR2_X1 U1007 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
XOR2_X1 U1008 ( .A(KEYINPUT24), .B(n1324), .Z(n1323) );
NOR2_X1 U1009 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
AND2_X1 U1010 ( .A1(n1326), .A2(n1325), .ZN(n1322) );
XNOR2_X1 U1011 ( .A(n1327), .B(n1328), .ZN(n1325) );
XNOR2_X1 U1012 ( .A(KEYINPUT25), .B(n1329), .ZN(n1328) );
INV_X1 U1013 ( .A(G122), .ZN(n1329) );
XNOR2_X1 U1014 ( .A(G107), .B(G116), .ZN(n1327) );
XOR2_X1 U1015 ( .A(G128), .B(n1330), .Z(n1326) );
XNOR2_X1 U1016 ( .A(n1317), .B(G134), .ZN(n1330) );
NAND2_X1 U1017 ( .A1(G217), .A2(n1331), .ZN(n1320) );
XNOR2_X1 U1018 ( .A(KEYINPUT40), .B(n1094), .ZN(n1302) );
INV_X1 U1019 ( .A(n1254), .ZN(n1094) );
NOR2_X1 U1020 ( .A1(n1283), .A2(n1299), .ZN(n1254) );
INV_X1 U1021 ( .A(n1109), .ZN(n1299) );
NAND3_X1 U1022 ( .A1(n1332), .A2(n1333), .A3(n1334), .ZN(n1109) );
NAND2_X1 U1023 ( .A1(G902), .A2(G217), .ZN(n1334) );
NAND3_X1 U1024 ( .A1(n1165), .A2(n1290), .A3(n1335), .ZN(n1333) );
OR2_X1 U1025 ( .A1(n1165), .A2(n1335), .ZN(n1332) );
NAND2_X1 U1026 ( .A1(G217), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1027 ( .A(n1337), .B(n1338), .Z(n1165) );
XNOR2_X1 U1028 ( .A(n1339), .B(n1136), .ZN(n1338) );
XOR2_X1 U1029 ( .A(G140), .B(n1243), .Z(n1136) );
XOR2_X1 U1030 ( .A(n1340), .B(n1341), .Z(n1337) );
XNOR2_X1 U1031 ( .A(G119), .B(n1342), .ZN(n1341) );
NAND2_X1 U1032 ( .A1(KEYINPUT1), .A2(n1343), .ZN(n1342) );
XNOR2_X1 U1033 ( .A(G137), .B(n1344), .ZN(n1343) );
NAND2_X1 U1034 ( .A1(G221), .A2(n1331), .ZN(n1344) );
NOR2_X1 U1035 ( .A1(n1336), .A2(G953), .ZN(n1331) );
INV_X1 U1036 ( .A(G234), .ZN(n1336) );
NAND2_X1 U1037 ( .A1(KEYINPUT2), .A2(n1345), .ZN(n1340) );
XOR2_X1 U1038 ( .A(G472), .B(n1346), .Z(n1283) );
NOR2_X1 U1039 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
NOR2_X1 U1040 ( .A1(KEYINPUT34), .A2(n1114), .ZN(n1348) );
AND2_X1 U1041 ( .A1(KEYINPUT51), .A2(n1114), .ZN(n1347) );
AND2_X1 U1042 ( .A1(n1349), .A2(n1290), .ZN(n1114) );
XNOR2_X1 U1043 ( .A(n1350), .B(n1177), .ZN(n1349) );
XOR2_X1 U1044 ( .A(G101), .B(n1351), .Z(n1177) );
AND3_X1 U1045 ( .A1(G210), .A2(n1068), .A3(n1318), .ZN(n1351) );
INV_X1 U1046 ( .A(G237), .ZN(n1318) );
NAND2_X1 U1047 ( .A1(n1182), .A2(n1183), .ZN(n1350) );
NAND2_X1 U1048 ( .A1(n1352), .A2(n1353), .ZN(n1183) );
OR2_X1 U1049 ( .A1(n1353), .A2(n1352), .ZN(n1182) );
XOR2_X1 U1050 ( .A(G113), .B(n1354), .Z(n1352) );
XOR2_X1 U1051 ( .A(n1193), .B(n1242), .Z(n1353) );
AND3_X1 U1052 ( .A1(n1252), .A2(n1297), .A3(n1063), .ZN(n1234) );
NOR2_X1 U1053 ( .A1(n1086), .A2(n1085), .ZN(n1063) );
INV_X1 U1054 ( .A(n1298), .ZN(n1085) );
NAND2_X1 U1055 ( .A1(G221), .A2(n1355), .ZN(n1298) );
NAND2_X1 U1056 ( .A1(G234), .A2(n1290), .ZN(n1355) );
XNOR2_X1 U1057 ( .A(n1356), .B(n1202), .ZN(n1086) );
INV_X1 U1058 ( .A(G469), .ZN(n1202) );
NAND2_X1 U1059 ( .A1(n1357), .A2(n1290), .ZN(n1356) );
XOR2_X1 U1060 ( .A(n1358), .B(n1359), .Z(n1357) );
XNOR2_X1 U1061 ( .A(n1360), .B(n1195), .ZN(n1359) );
INV_X1 U1062 ( .A(n1193), .ZN(n1195) );
XOR2_X1 U1063 ( .A(G131), .B(n1361), .Z(n1193) );
XOR2_X1 U1064 ( .A(G137), .B(G134), .Z(n1361) );
XOR2_X1 U1065 ( .A(n1362), .B(n1198), .Z(n1360) );
XNOR2_X1 U1066 ( .A(n1363), .B(G101), .ZN(n1198) );
NAND2_X1 U1067 ( .A1(KEYINPUT41), .A2(n1188), .ZN(n1362) );
XOR2_X1 U1068 ( .A(G140), .B(n1345), .Z(n1188) );
XOR2_X1 U1069 ( .A(n1364), .B(n1365), .Z(n1358) );
NOR2_X1 U1070 ( .A1(KEYINPUT55), .A2(n1141), .ZN(n1365) );
NAND2_X1 U1071 ( .A1(n1366), .A2(n1367), .ZN(n1141) );
OR2_X1 U1072 ( .A1(n1368), .A2(G128), .ZN(n1367) );
XOR2_X1 U1073 ( .A(n1369), .B(KEYINPUT21), .Z(n1366) );
NAND2_X1 U1074 ( .A1(G128), .A2(n1368), .ZN(n1369) );
NAND2_X1 U1075 ( .A1(n1370), .A2(n1371), .ZN(n1368) );
OR2_X1 U1076 ( .A1(n1311), .A2(n1317), .ZN(n1371) );
XOR2_X1 U1077 ( .A(n1372), .B(KEYINPUT8), .Z(n1370) );
NAND2_X1 U1078 ( .A1(n1311), .A2(n1317), .ZN(n1372) );
XOR2_X1 U1079 ( .A(n1199), .B(KEYINPUT32), .Z(n1364) );
NAND2_X1 U1080 ( .A1(G227), .A2(n1068), .ZN(n1199) );
NAND2_X1 U1081 ( .A1(n1100), .A2(n1373), .ZN(n1297) );
NAND4_X1 U1082 ( .A1(G953), .A2(G902), .A3(n1289), .A4(n1152), .ZN(n1373) );
INV_X1 U1083 ( .A(G898), .ZN(n1152) );
NAND3_X1 U1084 ( .A1(n1289), .A2(n1068), .A3(G952), .ZN(n1100) );
INV_X1 U1085 ( .A(G953), .ZN(n1068) );
NAND2_X1 U1086 ( .A1(G237), .A2(G234), .ZN(n1289) );
NOR2_X1 U1087 ( .A1(n1099), .A2(n1098), .ZN(n1252) );
AND2_X1 U1088 ( .A1(G214), .A2(n1374), .ZN(n1098) );
INV_X1 U1089 ( .A(n1281), .ZN(n1099) );
NAND3_X1 U1090 ( .A1(n1375), .A2(n1376), .A3(n1120), .ZN(n1281) );
NAND2_X1 U1091 ( .A1(n1122), .A2(n1121), .ZN(n1120) );
NAND2_X1 U1092 ( .A1(KEYINPUT6), .A2(n1121), .ZN(n1376) );
OR3_X1 U1093 ( .A1(n1122), .A2(KEYINPUT6), .A3(n1121), .ZN(n1375) );
NAND2_X1 U1094 ( .A1(n1377), .A2(n1290), .ZN(n1121) );
XOR2_X1 U1095 ( .A(n1204), .B(n1378), .Z(n1377) );
NOR2_X1 U1096 ( .A1(KEYINPUT44), .A2(n1379), .ZN(n1378) );
XOR2_X1 U1097 ( .A(n1380), .B(n1381), .Z(n1379) );
XOR2_X1 U1098 ( .A(n1239), .B(n1242), .Z(n1381) );
XNOR2_X1 U1099 ( .A(n1317), .B(n1339), .ZN(n1242) );
XNOR2_X1 U1100 ( .A(n1282), .B(n1311), .ZN(n1339) );
XOR2_X1 U1101 ( .A(G146), .B(KEYINPUT26), .Z(n1311) );
INV_X1 U1102 ( .A(G128), .ZN(n1282) );
INV_X1 U1103 ( .A(G143), .ZN(n1317) );
NOR2_X1 U1104 ( .A1(n1151), .A2(G953), .ZN(n1239) );
INV_X1 U1105 ( .A(G224), .ZN(n1151) );
XNOR2_X1 U1106 ( .A(KEYINPUT18), .B(n1243), .ZN(n1380) );
INV_X1 U1107 ( .A(G125), .ZN(n1243) );
XNOR2_X1 U1108 ( .A(n1382), .B(n1383), .ZN(n1204) );
INV_X1 U1109 ( .A(n1156), .ZN(n1383) );
XOR2_X1 U1110 ( .A(G122), .B(n1345), .Z(n1156) );
XOR2_X1 U1111 ( .A(G110), .B(KEYINPUT19), .Z(n1345) );
XNOR2_X1 U1112 ( .A(n1384), .B(n1159), .ZN(n1382) );
XOR2_X1 U1113 ( .A(n1363), .B(n1385), .Z(n1159) );
NOR2_X1 U1114 ( .A1(G101), .A2(KEYINPUT43), .ZN(n1385) );
XNOR2_X1 U1115 ( .A(G107), .B(n1310), .ZN(n1363) );
XOR2_X1 U1116 ( .A(G104), .B(KEYINPUT9), .Z(n1310) );
NAND2_X1 U1117 ( .A1(KEYINPUT33), .A2(n1160), .ZN(n1384) );
XNOR2_X1 U1118 ( .A(n1386), .B(n1387), .ZN(n1160) );
INV_X1 U1119 ( .A(G113), .ZN(n1387) );
NAND2_X1 U1120 ( .A1(KEYINPUT56), .A2(n1354), .ZN(n1386) );
XNOR2_X1 U1121 ( .A(n1388), .B(G116), .ZN(n1354) );
INV_X1 U1122 ( .A(G119), .ZN(n1388) );
AND2_X1 U1123 ( .A1(G210), .A2(n1374), .ZN(n1122) );
NAND2_X1 U1124 ( .A1(n1389), .A2(n1290), .ZN(n1374) );
INV_X1 U1125 ( .A(G902), .ZN(n1290) );
XNOR2_X1 U1126 ( .A(G237), .B(KEYINPUT42), .ZN(n1389) );
endmodule


