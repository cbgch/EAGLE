//Key = 1101111111110101011110000011010011001000110011000111011100111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272;

XNOR2_X1 U704 ( .A(G107), .B(n964), .ZN(G9) );
NAND4_X1 U705 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(n964) );
XOR2_X1 U706 ( .A(KEYINPUT16), .B(n969), .Z(n968) );
NOR2_X1 U707 ( .A1(n970), .A2(n971), .ZN(G75) );
NOR4_X1 U708 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(n971) );
NOR2_X1 U709 ( .A1(n976), .A2(n977), .ZN(n975) );
NOR2_X1 U710 ( .A1(n978), .A2(n979), .ZN(n974) );
NOR4_X1 U711 ( .A1(n980), .A2(n981), .A3(n982), .A4(n983), .ZN(n978) );
NAND3_X1 U712 ( .A1(n984), .A2(n985), .A3(n986), .ZN(n972) );
NAND3_X1 U713 ( .A1(n987), .A2(n988), .A3(n989), .ZN(n986) );
NAND2_X1 U714 ( .A1(n990), .A2(n991), .ZN(n988) );
INV_X1 U715 ( .A(n980), .ZN(n991) );
NAND2_X1 U716 ( .A1(n992), .A2(n993), .ZN(n990) );
NAND2_X1 U717 ( .A1(n994), .A2(n995), .ZN(n993) );
NAND3_X1 U718 ( .A1(n996), .A2(n997), .A3(n966), .ZN(n995) );
NAND2_X1 U719 ( .A1(n998), .A2(n999), .ZN(n994) );
NAND2_X1 U720 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NAND2_X1 U721 ( .A1(n966), .A2(n1002), .ZN(n1001) );
NAND2_X1 U722 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
NAND2_X1 U723 ( .A1(n1005), .A2(n1006), .ZN(n1004) );
XNOR2_X1 U724 ( .A(n1007), .B(n1008), .ZN(n1006) );
NAND2_X1 U725 ( .A1(n1009), .A2(n979), .ZN(n1003) );
INV_X1 U726 ( .A(KEYINPUT30), .ZN(n979) );
NAND2_X1 U727 ( .A1(n996), .A2(n1010), .ZN(n1000) );
OR2_X1 U728 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NAND2_X1 U729 ( .A1(n980), .A2(n1013), .ZN(n987) );
XOR2_X1 U730 ( .A(n977), .B(KEYINPUT23), .Z(n1013) );
OR2_X1 U731 ( .A1(n982), .A2(n1014), .ZN(n977) );
NAND3_X1 U732 ( .A1(n998), .A2(n966), .A3(n992), .ZN(n982) );
INV_X1 U733 ( .A(n1015), .ZN(n992) );
NOR3_X1 U734 ( .A1(n1016), .A2(G953), .A3(G952), .ZN(n970) );
INV_X1 U735 ( .A(n984), .ZN(n1016) );
NAND4_X1 U736 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n984) );
NOR3_X1 U737 ( .A1(n1021), .A2(n980), .A3(n1022), .ZN(n1020) );
XOR2_X1 U738 ( .A(n1023), .B(KEYINPUT54), .Z(n1022) );
NAND3_X1 U739 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1021) );
NOR3_X1 U740 ( .A1(n983), .A2(n1027), .A3(n1028), .ZN(n1019) );
NOR2_X1 U741 ( .A1(n1029), .A2(n1030), .ZN(n1028) );
XOR2_X1 U742 ( .A(KEYINPUT29), .B(n1031), .Z(n1030) );
NOR2_X1 U743 ( .A1(G469), .A2(n1032), .ZN(n1027) );
XNOR2_X1 U744 ( .A(n1031), .B(KEYINPUT7), .ZN(n1032) );
XNOR2_X1 U745 ( .A(n1033), .B(KEYINPUT13), .ZN(n1031) );
XNOR2_X1 U746 ( .A(KEYINPUT61), .B(n1034), .ZN(n1018) );
XOR2_X1 U747 ( .A(n1035), .B(n1036), .Z(G72) );
XOR2_X1 U748 ( .A(n1037), .B(n1038), .Z(n1036) );
NOR2_X1 U749 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
XNOR2_X1 U750 ( .A(KEYINPUT40), .B(n985), .ZN(n1040) );
NOR2_X1 U751 ( .A1(n1041), .A2(n1042), .ZN(n1039) );
NAND2_X1 U752 ( .A1(n1043), .A2(n1044), .ZN(n1037) );
NAND2_X1 U753 ( .A1(n1045), .A2(n1042), .ZN(n1044) );
XOR2_X1 U754 ( .A(n1046), .B(n1047), .Z(n1043) );
XNOR2_X1 U755 ( .A(n1048), .B(n1049), .ZN(n1047) );
XOR2_X1 U756 ( .A(n1050), .B(n1051), .Z(n1046) );
NAND2_X1 U757 ( .A1(n985), .A2(n1052), .ZN(n1035) );
XOR2_X1 U758 ( .A(n1053), .B(n1054), .Z(G69) );
XOR2_X1 U759 ( .A(n1055), .B(n1056), .Z(n1054) );
NOR2_X1 U760 ( .A1(n1057), .A2(G953), .ZN(n1056) );
NOR3_X1 U761 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1057) );
INV_X1 U762 ( .A(n1061), .ZN(n1059) );
NOR2_X1 U763 ( .A1(n1062), .A2(n1063), .ZN(n1055) );
XOR2_X1 U764 ( .A(n1064), .B(KEYINPUT28), .Z(n1063) );
NAND2_X1 U765 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U767 ( .A(n1069), .B(KEYINPUT37), .Z(n1065) );
OR2_X1 U768 ( .A1(n1068), .A2(n1067), .ZN(n1069) );
INV_X1 U769 ( .A(n1070), .ZN(n1067) );
AND2_X1 U770 ( .A1(n1071), .A2(n1045), .ZN(n1062) );
NOR2_X1 U771 ( .A1(n1072), .A2(n985), .ZN(n1053) );
NOR2_X1 U772 ( .A1(n1073), .A2(n1071), .ZN(n1072) );
NOR2_X1 U773 ( .A1(n1074), .A2(n1075), .ZN(G66) );
XNOR2_X1 U774 ( .A(n1076), .B(n1077), .ZN(n1075) );
NOR2_X1 U775 ( .A1(n1078), .A2(n1079), .ZN(n1076) );
NOR2_X1 U776 ( .A1(n1074), .A2(n1080), .ZN(G63) );
XNOR2_X1 U777 ( .A(n1081), .B(n1082), .ZN(n1080) );
XOR2_X1 U778 ( .A(KEYINPUT47), .B(n1083), .Z(n1082) );
NOR2_X1 U779 ( .A1(n1084), .A2(n1079), .ZN(n1083) );
NOR2_X1 U780 ( .A1(n1074), .A2(n1085), .ZN(G60) );
XNOR2_X1 U781 ( .A(n1086), .B(n1087), .ZN(n1085) );
NOR2_X1 U782 ( .A1(n1088), .A2(n1079), .ZN(n1087) );
XOR2_X1 U783 ( .A(G104), .B(n1089), .Z(G6) );
NOR4_X1 U784 ( .A1(KEYINPUT31), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1089) );
NOR2_X1 U785 ( .A1(n1074), .A2(n1093), .ZN(G57) );
XOR2_X1 U786 ( .A(n1094), .B(n1095), .Z(n1093) );
XOR2_X1 U787 ( .A(n1096), .B(n1097), .Z(n1095) );
XNOR2_X1 U788 ( .A(n1098), .B(n1099), .ZN(n1097) );
NOR2_X1 U789 ( .A1(KEYINPUT35), .A2(n1100), .ZN(n1099) );
XOR2_X1 U790 ( .A(KEYINPUT62), .B(KEYINPUT58), .Z(n1096) );
XOR2_X1 U791 ( .A(n1101), .B(n1102), .Z(n1094) );
XNOR2_X1 U792 ( .A(n1103), .B(n1104), .ZN(n1101) );
NOR2_X1 U793 ( .A1(n1079), .A2(n1105), .ZN(n1104) );
XOR2_X1 U794 ( .A(KEYINPUT50), .B(G472), .Z(n1105) );
NOR2_X1 U795 ( .A1(n1074), .A2(n1106), .ZN(G54) );
XOR2_X1 U796 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U797 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XOR2_X1 U799 ( .A(KEYINPUT2), .B(n1113), .Z(n1112) );
NOR2_X1 U800 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
XOR2_X1 U801 ( .A(n1116), .B(KEYINPUT18), .Z(n1115) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1117), .ZN(n1111) );
XOR2_X1 U803 ( .A(n1118), .B(n1119), .Z(n1116) );
NOR2_X1 U804 ( .A1(KEYINPUT43), .A2(n1120), .ZN(n1109) );
XOR2_X1 U805 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U806 ( .A(n1123), .B(n1124), .ZN(n1122) );
INV_X1 U807 ( .A(G110), .ZN(n1123) );
NAND2_X1 U808 ( .A1(KEYINPUT1), .A2(n1048), .ZN(n1121) );
NAND2_X1 U809 ( .A1(KEYINPUT9), .A2(n1125), .ZN(n1107) );
OR2_X1 U810 ( .A1(n1079), .A2(n1029), .ZN(n1125) );
NOR2_X1 U811 ( .A1(n1074), .A2(n1126), .ZN(G51) );
XNOR2_X1 U812 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U813 ( .A1(n1129), .A2(n1079), .ZN(n1128) );
NAND2_X1 U814 ( .A1(G902), .A2(n973), .ZN(n1079) );
NAND4_X1 U815 ( .A1(n1130), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n973) );
XNOR2_X1 U816 ( .A(KEYINPUT56), .B(n1060), .ZN(n1133) );
NAND4_X1 U817 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1060) );
NAND4_X1 U818 ( .A1(n1138), .A2(n1011), .A3(n965), .A4(n1139), .ZN(n1134) );
XNOR2_X1 U819 ( .A(KEYINPUT52), .B(n976), .ZN(n1139) );
INV_X1 U820 ( .A(n1140), .ZN(n976) );
XNOR2_X1 U821 ( .A(KEYINPUT63), .B(n1061), .ZN(n1132) );
INV_X1 U822 ( .A(n1058), .ZN(n1131) );
NAND2_X1 U823 ( .A1(n1141), .A2(n1142), .ZN(n1058) );
NAND3_X1 U824 ( .A1(n966), .A2(n997), .A3(n1143), .ZN(n1142) );
NAND2_X1 U825 ( .A1(n1091), .A2(n1144), .ZN(n997) );
INV_X1 U826 ( .A(n1052), .ZN(n1130) );
NAND4_X1 U827 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1052) );
NOR4_X1 U828 ( .A1(n1149), .A2(n1150), .A3(n1151), .A4(n1152), .ZN(n1148) );
INV_X1 U829 ( .A(n1153), .ZN(n1149) );
AND2_X1 U830 ( .A1(n1154), .A2(n1155), .ZN(n1147) );
NOR2_X1 U831 ( .A1(n985), .A2(G952), .ZN(n1074) );
XNOR2_X1 U832 ( .A(G146), .B(n1155), .ZN(G48) );
NAND4_X1 U833 ( .A1(n1156), .A2(n1157), .A3(n1009), .A4(n1158), .ZN(n1155) );
XNOR2_X1 U834 ( .A(G143), .B(n1154), .ZN(G45) );
NAND4_X1 U835 ( .A1(n1159), .A2(n1011), .A3(n1009), .A4(n1158), .ZN(n1154) );
NAND2_X1 U836 ( .A1(n1160), .A2(n1161), .ZN(G42) );
NAND2_X1 U837 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XNOR2_X1 U838 ( .A(G140), .B(KEYINPUT19), .ZN(n1163) );
XOR2_X1 U839 ( .A(n1145), .B(KEYINPUT39), .Z(n1162) );
NAND2_X1 U840 ( .A1(n1164), .A2(n1048), .ZN(n1160) );
XOR2_X1 U841 ( .A(n1145), .B(KEYINPUT17), .Z(n1164) );
NAND3_X1 U842 ( .A1(n1012), .A2(n1157), .A3(n1165), .ZN(n1145) );
XNOR2_X1 U843 ( .A(G137), .B(n1146), .ZN(G39) );
NAND4_X1 U844 ( .A1(n1166), .A2(n998), .A3(n1165), .A4(n1167), .ZN(n1146) );
XOR2_X1 U845 ( .A(G134), .B(n1151), .Z(G36) );
AND3_X1 U846 ( .A1(n1011), .A2(n965), .A3(n1165), .ZN(n1151) );
XOR2_X1 U847 ( .A(G131), .B(n1150), .Z(G33) );
AND3_X1 U848 ( .A1(n1011), .A2(n1157), .A3(n1165), .ZN(n1150) );
NOR4_X1 U849 ( .A1(n983), .A2(n981), .A3(n1168), .A4(n980), .ZN(n1165) );
INV_X1 U850 ( .A(n1009), .ZN(n981) );
XOR2_X1 U851 ( .A(n969), .B(KEYINPUT46), .Z(n1009) );
XOR2_X1 U852 ( .A(G128), .B(n1152), .Z(G30) );
AND4_X1 U853 ( .A1(n1156), .A2(n965), .A3(n969), .A4(n1158), .ZN(n1152) );
XNOR2_X1 U854 ( .A(G101), .B(n1141), .ZN(G3) );
NAND3_X1 U855 ( .A1(n998), .A2(n1011), .A3(n1143), .ZN(n1141) );
XNOR2_X1 U856 ( .A(G125), .B(n1153), .ZN(G27) );
NAND4_X1 U857 ( .A1(n1012), .A2(n1157), .A3(n1169), .A4(n1140), .ZN(n1153) );
NOR2_X1 U858 ( .A1(n1168), .A2(n1014), .ZN(n1169) );
INV_X1 U859 ( .A(n996), .ZN(n1014) );
INV_X1 U860 ( .A(n1158), .ZN(n1168) );
NAND2_X1 U861 ( .A1(n1015), .A2(n1170), .ZN(n1158) );
NAND2_X1 U862 ( .A1(n1171), .A2(n1042), .ZN(n1170) );
INV_X1 U863 ( .A(G900), .ZN(n1042) );
XNOR2_X1 U864 ( .A(G122), .B(n1135), .ZN(G24) );
NAND3_X1 U865 ( .A1(n1159), .A2(n966), .A3(n1138), .ZN(n1135) );
INV_X1 U866 ( .A(n1090), .ZN(n966) );
NAND2_X1 U867 ( .A1(n1023), .A2(n1034), .ZN(n1090) );
INV_X1 U868 ( .A(n1167), .ZN(n1034) );
AND3_X1 U869 ( .A1(n1140), .A2(n1172), .A3(n1173), .ZN(n1159) );
XNOR2_X1 U870 ( .A(G119), .B(n1136), .ZN(G21) );
NAND3_X1 U871 ( .A1(n998), .A2(n1156), .A3(n1138), .ZN(n1136) );
AND3_X1 U872 ( .A1(n1140), .A2(n1167), .A3(n1166), .ZN(n1156) );
XOR2_X1 U873 ( .A(n1174), .B(KEYINPUT60), .Z(n1166) );
XNOR2_X1 U874 ( .A(G116), .B(n1175), .ZN(G18) );
NAND4_X1 U875 ( .A1(n1138), .A2(n1011), .A3(n965), .A4(n1140), .ZN(n1175) );
XOR2_X1 U876 ( .A(n1176), .B(KEYINPUT42), .Z(n1140) );
INV_X1 U877 ( .A(n1144), .ZN(n965) );
NAND2_X1 U878 ( .A1(n1177), .A2(n1172), .ZN(n1144) );
XOR2_X1 U879 ( .A(n1173), .B(KEYINPUT5), .Z(n1177) );
XNOR2_X1 U880 ( .A(G113), .B(n1137), .ZN(G15) );
NAND4_X1 U881 ( .A1(n1138), .A2(n1011), .A3(n1157), .A4(n1176), .ZN(n1137) );
INV_X1 U882 ( .A(n1091), .ZN(n1157) );
NAND2_X1 U883 ( .A1(n1178), .A2(n1173), .ZN(n1091) );
INV_X1 U884 ( .A(n1172), .ZN(n1178) );
AND2_X1 U885 ( .A1(n1023), .A2(n1167), .ZN(n1011) );
AND2_X1 U886 ( .A1(n996), .A2(n1179), .ZN(n1138) );
NAND2_X1 U887 ( .A1(n1180), .A2(n1181), .ZN(n996) );
NAND3_X1 U888 ( .A1(n1008), .A2(n1026), .A3(n1007), .ZN(n1181) );
INV_X1 U889 ( .A(KEYINPUT12), .ZN(n1007) );
NAND2_X1 U890 ( .A1(KEYINPUT12), .A2(n969), .ZN(n1180) );
XNOR2_X1 U891 ( .A(G110), .B(n1061), .ZN(G12) );
NAND3_X1 U892 ( .A1(n998), .A2(n1012), .A3(n1143), .ZN(n1061) );
INV_X1 U893 ( .A(n1092), .ZN(n1143) );
NAND2_X1 U894 ( .A1(n967), .A2(n969), .ZN(n1092) );
NOR2_X1 U895 ( .A1(n1008), .A2(n1005), .ZN(n969) );
INV_X1 U896 ( .A(n1026), .ZN(n1005) );
NAND2_X1 U897 ( .A1(G221), .A2(n1182), .ZN(n1026) );
XOR2_X1 U898 ( .A(n1183), .B(n1029), .Z(n1008) );
INV_X1 U899 ( .A(G469), .ZN(n1029) );
NAND2_X1 U900 ( .A1(KEYINPUT36), .A2(n1033), .ZN(n1183) );
NAND2_X1 U901 ( .A1(n1184), .A2(n1185), .ZN(n1033) );
XOR2_X1 U902 ( .A(n1186), .B(n1187), .Z(n1184) );
XNOR2_X1 U903 ( .A(n1114), .B(n1119), .ZN(n1187) );
XNOR2_X1 U904 ( .A(n1188), .B(n1189), .ZN(n1186) );
XOR2_X1 U905 ( .A(n1124), .B(n1190), .Z(n1189) );
NOR2_X1 U906 ( .A1(KEYINPUT38), .A2(n1118), .ZN(n1190) );
XNOR2_X1 U907 ( .A(n1049), .B(G128), .ZN(n1118) );
AND2_X1 U908 ( .A1(n1191), .A2(n1192), .ZN(n1049) );
NAND2_X1 U909 ( .A1(G146), .A2(n1193), .ZN(n1192) );
XOR2_X1 U910 ( .A(KEYINPUT11), .B(n1194), .Z(n1191) );
NOR2_X1 U911 ( .A1(n1195), .A2(n1193), .ZN(n1194) );
XNOR2_X1 U912 ( .A(G146), .B(KEYINPUT41), .ZN(n1195) );
NOR2_X1 U913 ( .A1(n1041), .A2(G953), .ZN(n1124) );
INV_X1 U914 ( .A(G227), .ZN(n1041) );
AND2_X1 U915 ( .A1(n1176), .A2(n1179), .ZN(n967) );
NAND2_X1 U916 ( .A1(n1015), .A2(n1196), .ZN(n1179) );
NAND2_X1 U917 ( .A1(n1171), .A2(n1071), .ZN(n1196) );
INV_X1 U918 ( .A(G898), .ZN(n1071) );
AND3_X1 U919 ( .A1(n1045), .A2(n1197), .A3(n1198), .ZN(n1171) );
XNOR2_X1 U920 ( .A(G902), .B(KEYINPUT6), .ZN(n1198) );
XOR2_X1 U921 ( .A(G953), .B(KEYINPUT25), .Z(n1045) );
NAND3_X1 U922 ( .A1(n1197), .A2(n985), .A3(G952), .ZN(n1015) );
NAND2_X1 U923 ( .A1(G237), .A2(G234), .ZN(n1197) );
NOR2_X1 U924 ( .A1(n989), .A2(n980), .ZN(n1176) );
NOR2_X1 U925 ( .A1(n1199), .A2(n1200), .ZN(n980) );
INV_X1 U926 ( .A(G214), .ZN(n1199) );
INV_X1 U927 ( .A(n983), .ZN(n989) );
XNOR2_X1 U928 ( .A(n1201), .B(n1202), .ZN(n983) );
NOR2_X1 U929 ( .A1(n1200), .A2(n1203), .ZN(n1202) );
XNOR2_X1 U930 ( .A(KEYINPUT45), .B(n1129), .ZN(n1203) );
INV_X1 U931 ( .A(G210), .ZN(n1129) );
NOR2_X1 U932 ( .A1(G902), .A2(G237), .ZN(n1200) );
NAND2_X1 U933 ( .A1(n1204), .A2(n1127), .ZN(n1201) );
XNOR2_X1 U934 ( .A(n1205), .B(n1206), .ZN(n1127) );
XNOR2_X1 U935 ( .A(n1207), .B(n1068), .ZN(n1206) );
XOR2_X1 U936 ( .A(n1119), .B(n1208), .Z(n1068) );
NOR2_X1 U937 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
XOR2_X1 U938 ( .A(KEYINPUT48), .B(n1211), .Z(n1210) );
NOR2_X1 U939 ( .A1(G113), .A2(n1212), .ZN(n1211) );
AND2_X1 U940 ( .A1(n1212), .A2(G113), .ZN(n1209) );
XOR2_X1 U941 ( .A(G116), .B(G119), .Z(n1212) );
XOR2_X1 U942 ( .A(G101), .B(n1213), .Z(n1119) );
XNOR2_X1 U943 ( .A(n1214), .B(G104), .ZN(n1213) );
INV_X1 U944 ( .A(G107), .ZN(n1214) );
INV_X1 U945 ( .A(n1103), .ZN(n1207) );
XOR2_X1 U946 ( .A(n1215), .B(n1216), .Z(n1205) );
XNOR2_X1 U947 ( .A(n1217), .B(n1218), .ZN(n1216) );
NOR2_X1 U948 ( .A1(G953), .A2(n1073), .ZN(n1218) );
INV_X1 U949 ( .A(G224), .ZN(n1073) );
INV_X1 U950 ( .A(G125), .ZN(n1217) );
NAND2_X1 U951 ( .A1(KEYINPUT33), .A2(n1070), .ZN(n1215) );
XNOR2_X1 U952 ( .A(G110), .B(n1219), .ZN(n1070) );
XNOR2_X1 U953 ( .A(KEYINPUT0), .B(n1185), .ZN(n1204) );
NOR2_X1 U954 ( .A1(n1167), .A2(n1174), .ZN(n1012) );
XOR2_X1 U955 ( .A(n1023), .B(KEYINPUT57), .Z(n1174) );
XNOR2_X1 U956 ( .A(n1220), .B(n1078), .ZN(n1023) );
NAND2_X1 U957 ( .A1(G217), .A2(n1182), .ZN(n1078) );
NAND2_X1 U958 ( .A1(G234), .A2(n1185), .ZN(n1182) );
NAND2_X1 U959 ( .A1(n1077), .A2(n1221), .ZN(n1220) );
XNOR2_X1 U960 ( .A(KEYINPUT27), .B(n1185), .ZN(n1221) );
XOR2_X1 U961 ( .A(n1222), .B(n1223), .Z(n1077) );
XOR2_X1 U962 ( .A(n1050), .B(n1224), .Z(n1223) );
XOR2_X1 U963 ( .A(n1225), .B(n1188), .Z(n1224) );
XOR2_X1 U964 ( .A(G110), .B(G140), .Z(n1188) );
NAND2_X1 U965 ( .A1(KEYINPUT10), .A2(n1226), .ZN(n1225) );
INV_X1 U966 ( .A(G137), .ZN(n1226) );
XNOR2_X1 U967 ( .A(G125), .B(G128), .ZN(n1050) );
XOR2_X1 U968 ( .A(n1227), .B(n1228), .Z(n1222) );
XOR2_X1 U969 ( .A(KEYINPUT14), .B(G146), .Z(n1228) );
XOR2_X1 U970 ( .A(n1229), .B(G119), .Z(n1227) );
NAND2_X1 U971 ( .A1(G221), .A2(n1230), .ZN(n1229) );
XNOR2_X1 U972 ( .A(n1231), .B(G472), .ZN(n1167) );
NAND2_X1 U973 ( .A1(n1232), .A2(n1185), .ZN(n1231) );
XOR2_X1 U974 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U975 ( .A(n1100), .B(n1235), .Z(n1234) );
NAND2_X1 U976 ( .A1(n1236), .A2(KEYINPUT26), .ZN(n1235) );
XNOR2_X1 U977 ( .A(n1102), .B(n1237), .ZN(n1236) );
XNOR2_X1 U978 ( .A(n1238), .B(KEYINPUT22), .ZN(n1237) );
NAND2_X1 U979 ( .A1(KEYINPUT8), .A2(n1103), .ZN(n1238) );
XNOR2_X1 U980 ( .A(n1239), .B(n1240), .ZN(n1103) );
XOR2_X1 U981 ( .A(KEYINPUT24), .B(G146), .Z(n1240) );
XNOR2_X1 U982 ( .A(G128), .B(G143), .ZN(n1239) );
XNOR2_X1 U983 ( .A(n1241), .B(n1242), .ZN(n1102) );
XNOR2_X1 U984 ( .A(n1243), .B(n1244), .ZN(n1242) );
XOR2_X1 U985 ( .A(KEYINPUT15), .B(G119), .Z(n1244) );
XNOR2_X1 U986 ( .A(n1245), .B(n1114), .ZN(n1241) );
INV_X1 U987 ( .A(n1117), .ZN(n1114) );
XOR2_X1 U988 ( .A(n1051), .B(KEYINPUT55), .Z(n1117) );
XNOR2_X1 U989 ( .A(n1246), .B(n1247), .ZN(n1051) );
XNOR2_X1 U990 ( .A(G131), .B(G137), .ZN(n1246) );
NAND2_X1 U991 ( .A1(KEYINPUT32), .A2(G116), .ZN(n1245) );
NAND2_X1 U992 ( .A1(G210), .A2(n1248), .ZN(n1100) );
NAND2_X1 U993 ( .A1(KEYINPUT4), .A2(n1098), .ZN(n1233) );
INV_X1 U994 ( .A(G101), .ZN(n1098) );
NOR2_X1 U995 ( .A1(n1172), .A2(n1173), .ZN(n998) );
XOR2_X1 U996 ( .A(n1017), .B(KEYINPUT59), .Z(n1173) );
XNOR2_X1 U997 ( .A(n1249), .B(n1088), .ZN(n1017) );
INV_X1 U998 ( .A(G475), .ZN(n1088) );
NAND2_X1 U999 ( .A1(n1086), .A2(n1185), .ZN(n1249) );
XNOR2_X1 U1000 ( .A(n1250), .B(n1251), .ZN(n1086) );
XOR2_X1 U1001 ( .A(n1252), .B(n1253), .Z(n1251) );
XNOR2_X1 U1002 ( .A(n1219), .B(G104), .ZN(n1253) );
XNOR2_X1 U1003 ( .A(n1193), .B(G131), .ZN(n1252) );
XOR2_X1 U1004 ( .A(n1254), .B(n1255), .Z(n1250) );
XOR2_X1 U1005 ( .A(n1256), .B(n1257), .Z(n1255) );
NAND2_X1 U1006 ( .A1(G214), .A2(n1248), .ZN(n1257) );
NOR2_X1 U1007 ( .A1(G953), .A2(G237), .ZN(n1248) );
NAND2_X1 U1008 ( .A1(KEYINPUT51), .A2(n1258), .ZN(n1256) );
XOR2_X1 U1009 ( .A(n1259), .B(n1260), .Z(n1258) );
XNOR2_X1 U1010 ( .A(G125), .B(G146), .ZN(n1260) );
NAND2_X1 U1011 ( .A1(KEYINPUT3), .A2(n1048), .ZN(n1259) );
INV_X1 U1012 ( .A(G140), .ZN(n1048) );
NAND2_X1 U1013 ( .A1(KEYINPUT20), .A2(n1243), .ZN(n1254) );
INV_X1 U1014 ( .A(G113), .ZN(n1243) );
NAND2_X1 U1015 ( .A1(n1261), .A2(n1024), .ZN(n1172) );
NAND3_X1 U1016 ( .A1(n1084), .A2(n1185), .A3(n1081), .ZN(n1024) );
INV_X1 U1017 ( .A(G478), .ZN(n1084) );
XNOR2_X1 U1018 ( .A(KEYINPUT53), .B(n1025), .ZN(n1261) );
NAND2_X1 U1019 ( .A1(G478), .A2(n1262), .ZN(n1025) );
NAND2_X1 U1020 ( .A1(n1081), .A2(n1185), .ZN(n1262) );
INV_X1 U1021 ( .A(G902), .ZN(n1185) );
XNOR2_X1 U1022 ( .A(n1263), .B(n1264), .ZN(n1081) );
XOR2_X1 U1023 ( .A(n1265), .B(n1266), .Z(n1264) );
XNOR2_X1 U1024 ( .A(G107), .B(G128), .ZN(n1266) );
NAND3_X1 U1025 ( .A1(KEYINPUT44), .A2(n1267), .A3(n1268), .ZN(n1265) );
XOR2_X1 U1026 ( .A(n1269), .B(KEYINPUT34), .Z(n1268) );
NAND2_X1 U1027 ( .A1(G116), .A2(n1219), .ZN(n1269) );
OR2_X1 U1028 ( .A1(n1219), .A2(G116), .ZN(n1267) );
INV_X1 U1029 ( .A(G122), .ZN(n1219) );
XOR2_X1 U1030 ( .A(n1270), .B(n1247), .Z(n1263) );
XOR2_X1 U1031 ( .A(G134), .B(KEYINPUT49), .Z(n1247) );
XOR2_X1 U1032 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U1033 ( .A1(KEYINPUT21), .A2(n1193), .ZN(n1272) );
INV_X1 U1034 ( .A(G143), .ZN(n1193) );
NAND2_X1 U1035 ( .A1(G217), .A2(n1230), .ZN(n1271) );
AND2_X1 U1036 ( .A1(G234), .A2(n985), .ZN(n1230) );
INV_X1 U1037 ( .A(G953), .ZN(n985) );
endmodule


