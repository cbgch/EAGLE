//Key = 0101000111011011110010011001001011010111011101101010010111000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;

XNOR2_X1 U742 ( .A(G107), .B(n1009), .ZN(G9) );
NOR2_X1 U743 ( .A1(n1010), .A2(n1011), .ZN(G75) );
NOR4_X1 U744 ( .A1(n1012), .A2(n1013), .A3(n1014), .A4(n1015), .ZN(n1011) );
NAND4_X1 U745 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1012) );
NAND3_X1 U746 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1017) );
NAND2_X1 U747 ( .A1(n1023), .A2(n1024), .ZN(n1020) );
NAND4_X1 U748 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
INV_X1 U749 ( .A(KEYINPUT17), .ZN(n1028) );
NAND2_X1 U750 ( .A1(n1029), .A2(n1030), .ZN(n1023) );
NAND2_X1 U751 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
OR2_X1 U752 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
NAND2_X1 U753 ( .A1(n1035), .A2(n1036), .ZN(n1031) );
NAND2_X1 U754 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U755 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U756 ( .A1(n1025), .A2(n1041), .ZN(n1016) );
NAND2_X1 U757 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U758 ( .A1(n1027), .A2(n1021), .A3(n1035), .ZN(n1043) );
NAND3_X1 U759 ( .A1(n1044), .A2(n1045), .A3(n1035), .ZN(n1027) );
NAND2_X1 U760 ( .A1(n1029), .A2(n1046), .ZN(n1045) );
OR2_X1 U761 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NAND2_X1 U762 ( .A1(n1022), .A2(n1049), .ZN(n1044) );
NAND2_X1 U763 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U764 ( .A1(KEYINPUT17), .A2(n1026), .ZN(n1051) );
XOR2_X1 U765 ( .A(n1052), .B(KEYINPUT40), .Z(n1042) );
NAND4_X1 U766 ( .A1(n1029), .A2(n1021), .A3(n1053), .A4(n1054), .ZN(n1052) );
NOR2_X1 U767 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR3_X1 U768 ( .A1(n1057), .A2(G953), .A3(n1058), .ZN(n1010) );
INV_X1 U769 ( .A(n1018), .ZN(n1058) );
NAND4_X1 U770 ( .A1(n1039), .A2(n1035), .A3(n1059), .A4(n1060), .ZN(n1018) );
NOR4_X1 U771 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1060) );
XNOR2_X1 U772 ( .A(n1065), .B(n1066), .ZN(n1062) );
NOR2_X1 U773 ( .A1(n1067), .A2(KEYINPUT63), .ZN(n1066) );
XOR2_X1 U774 ( .A(n1068), .B(n1069), .Z(n1061) );
XOR2_X1 U775 ( .A(KEYINPUT44), .B(G475), .Z(n1069) );
NAND2_X1 U776 ( .A1(KEYINPUT27), .A2(n1070), .ZN(n1068) );
XNOR2_X1 U777 ( .A(n1040), .B(KEYINPUT34), .ZN(n1059) );
XNOR2_X1 U778 ( .A(KEYINPUT0), .B(n1014), .ZN(n1057) );
INV_X1 U779 ( .A(G952), .ZN(n1014) );
XOR2_X1 U780 ( .A(n1071), .B(n1072), .Z(G72) );
NOR2_X1 U781 ( .A1(n1073), .A2(n1019), .ZN(n1072) );
AND2_X1 U782 ( .A1(G227), .A2(G900), .ZN(n1073) );
NAND2_X1 U783 ( .A1(n1074), .A2(n1075), .ZN(n1071) );
NAND2_X1 U784 ( .A1(n1076), .A2(n1019), .ZN(n1075) );
XOR2_X1 U785 ( .A(n1077), .B(n1015), .Z(n1076) );
NAND3_X1 U786 ( .A1(n1077), .A2(G900), .A3(G953), .ZN(n1074) );
NOR2_X1 U787 ( .A1(KEYINPUT22), .A2(n1078), .ZN(n1077) );
XOR2_X1 U788 ( .A(n1079), .B(n1080), .Z(n1078) );
XNOR2_X1 U789 ( .A(n1081), .B(n1082), .ZN(n1080) );
XOR2_X1 U790 ( .A(n1083), .B(n1084), .Z(n1079) );
XNOR2_X1 U791 ( .A(G137), .B(n1085), .ZN(n1084) );
NAND2_X1 U792 ( .A1(KEYINPUT38), .A2(n1086), .ZN(n1085) );
NAND2_X1 U793 ( .A1(KEYINPUT15), .A2(n1087), .ZN(n1083) );
XOR2_X1 U794 ( .A(n1088), .B(n1089), .Z(G69) );
XOR2_X1 U795 ( .A(n1090), .B(n1091), .Z(n1089) );
NAND3_X1 U796 ( .A1(n1013), .A2(n1019), .A3(KEYINPUT11), .ZN(n1091) );
NAND2_X1 U797 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
XOR2_X1 U798 ( .A(KEYINPUT24), .B(n1094), .Z(n1093) );
NOR2_X1 U799 ( .A1(n1095), .A2(n1019), .ZN(n1088) );
AND2_X1 U800 ( .A1(G224), .A2(G898), .ZN(n1095) );
NOR2_X1 U801 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XOR2_X1 U802 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U803 ( .A1(KEYINPUT53), .A2(n1100), .ZN(n1099) );
NAND2_X1 U804 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
XOR2_X1 U805 ( .A(n1103), .B(G217), .Z(n1101) );
XNOR2_X1 U806 ( .A(KEYINPUT9), .B(KEYINPUT19), .ZN(n1103) );
NOR2_X1 U807 ( .A1(n1096), .A2(n1104), .ZN(G63) );
XNOR2_X1 U808 ( .A(n1105), .B(n1106), .ZN(n1104) );
AND2_X1 U809 ( .A1(G478), .A2(n1102), .ZN(n1105) );
NOR2_X1 U810 ( .A1(n1096), .A2(n1107), .ZN(G60) );
XNOR2_X1 U811 ( .A(n1108), .B(n1109), .ZN(n1107) );
AND2_X1 U812 ( .A1(G475), .A2(n1102), .ZN(n1108) );
XNOR2_X1 U813 ( .A(G104), .B(n1110), .ZN(G6) );
NOR2_X1 U814 ( .A1(n1096), .A2(n1111), .ZN(G57) );
NOR2_X1 U815 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U816 ( .A(KEYINPUT18), .B(n1114), .Z(n1113) );
NOR2_X1 U817 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
XOR2_X1 U818 ( .A(KEYINPUT4), .B(n1117), .Z(n1116) );
AND2_X1 U819 ( .A1(n1115), .A2(n1117), .ZN(n1112) );
XNOR2_X1 U820 ( .A(n1118), .B(n1119), .ZN(n1117) );
NOR2_X1 U821 ( .A1(KEYINPUT5), .A2(n1120), .ZN(n1119) );
XOR2_X1 U822 ( .A(n1121), .B(n1122), .Z(n1120) );
XNOR2_X1 U823 ( .A(KEYINPUT6), .B(n1123), .ZN(n1121) );
NOR2_X1 U824 ( .A1(KEYINPUT36), .A2(n1124), .ZN(n1123) );
NAND2_X1 U825 ( .A1(n1102), .A2(G472), .ZN(n1118) );
NAND3_X1 U826 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1115) );
NAND2_X1 U827 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
OR3_X1 U828 ( .A1(n1129), .A2(n1130), .A3(G101), .ZN(n1126) );
INV_X1 U829 ( .A(KEYINPUT41), .ZN(n1129) );
NAND2_X1 U830 ( .A1(G101), .A2(n1130), .ZN(n1125) );
NAND2_X1 U831 ( .A1(KEYINPUT23), .A2(n1131), .ZN(n1130) );
NOR2_X1 U832 ( .A1(n1096), .A2(n1132), .ZN(G54) );
XOR2_X1 U833 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U834 ( .A(n1135), .B(n1136), .Z(n1134) );
XOR2_X1 U835 ( .A(n1137), .B(n1138), .Z(n1136) );
NAND2_X1 U836 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U837 ( .A1(n1141), .A2(n1082), .ZN(n1140) );
XOR2_X1 U838 ( .A(KEYINPUT12), .B(n1142), .Z(n1139) );
NOR2_X1 U839 ( .A1(n1082), .A2(n1141), .ZN(n1142) );
INV_X1 U840 ( .A(n1143), .ZN(n1141) );
INV_X1 U841 ( .A(n1144), .ZN(n1082) );
AND2_X1 U842 ( .A1(G469), .A2(n1102), .ZN(n1135) );
INV_X1 U843 ( .A(n1145), .ZN(n1102) );
XNOR2_X1 U844 ( .A(n1146), .B(n1147), .ZN(n1133) );
NAND2_X1 U845 ( .A1(n1148), .A2(KEYINPUT14), .ZN(n1146) );
XOR2_X1 U846 ( .A(n1149), .B(G110), .Z(n1148) );
NAND2_X1 U847 ( .A1(KEYINPUT16), .A2(n1150), .ZN(n1149) );
NOR2_X1 U848 ( .A1(n1096), .A2(n1151), .ZN(G51) );
XNOR2_X1 U849 ( .A(n1152), .B(n1153), .ZN(n1151) );
XNOR2_X1 U850 ( .A(n1154), .B(n1155), .ZN(n1153) );
NOR3_X1 U851 ( .A1(n1145), .A2(KEYINPUT21), .A3(n1156), .ZN(n1155) );
NAND2_X1 U852 ( .A1(G902), .A2(n1157), .ZN(n1145) );
OR2_X1 U853 ( .A1(n1013), .A2(n1015), .ZN(n1157) );
NAND2_X1 U854 ( .A1(n1158), .A2(n1159), .ZN(n1015) );
NOR4_X1 U855 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1159) );
INV_X1 U856 ( .A(n1164), .ZN(n1163) );
INV_X1 U857 ( .A(n1165), .ZN(n1160) );
NOR4_X1 U858 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1158) );
NOR2_X1 U859 ( .A1(n1033), .A2(n1170), .ZN(n1169) );
NOR2_X1 U860 ( .A1(n1171), .A2(n1172), .ZN(n1168) );
INV_X1 U861 ( .A(n1173), .ZN(n1167) );
NAND4_X1 U862 ( .A1(n1174), .A2(n1110), .A3(n1175), .A4(n1176), .ZN(n1013) );
AND4_X1 U863 ( .A1(n1009), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1176) );
NAND3_X1 U864 ( .A1(n1048), .A2(n1029), .A3(n1180), .ZN(n1009) );
NAND2_X1 U865 ( .A1(n1022), .A2(n1181), .ZN(n1175) );
NAND2_X1 U866 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U867 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U868 ( .A1(n1186), .A2(n1180), .ZN(n1182) );
NAND3_X1 U869 ( .A1(n1180), .A2(n1029), .A3(n1047), .ZN(n1110) );
NAND4_X1 U870 ( .A1(n1187), .A2(n1184), .A3(n1029), .A4(n1064), .ZN(n1174) );
INV_X1 U871 ( .A(n1188), .ZN(n1187) );
NAND2_X1 U872 ( .A1(KEYINPUT39), .A2(n1189), .ZN(n1154) );
XNOR2_X1 U873 ( .A(n1190), .B(n1191), .ZN(n1189) );
NOR2_X1 U874 ( .A1(n1019), .A2(G952), .ZN(n1096) );
XNOR2_X1 U875 ( .A(G146), .B(n1173), .ZN(G48) );
NAND4_X1 U876 ( .A1(n1192), .A2(n1047), .A3(n1185), .A4(n1193), .ZN(n1173) );
XOR2_X1 U877 ( .A(G143), .B(n1166), .Z(G45) );
AND3_X1 U878 ( .A1(n1192), .A2(n1186), .A3(n1194), .ZN(n1166) );
NOR3_X1 U879 ( .A1(n1188), .A2(n1195), .A3(n1037), .ZN(n1194) );
XNOR2_X1 U880 ( .A(n1150), .B(n1162), .ZN(G42) );
AND2_X1 U881 ( .A1(n1196), .A2(n1026), .ZN(n1162) );
XNOR2_X1 U882 ( .A(n1197), .B(n1198), .ZN(G39) );
NOR2_X1 U883 ( .A1(n1199), .A2(n1033), .ZN(n1198) );
INV_X1 U884 ( .A(n1025), .ZN(n1033) );
XOR2_X1 U885 ( .A(n1170), .B(KEYINPUT26), .Z(n1199) );
NAND3_X1 U886 ( .A1(n1022), .A2(n1185), .A3(n1192), .ZN(n1170) );
XNOR2_X1 U887 ( .A(G134), .B(n1164), .ZN(G36) );
NAND4_X1 U888 ( .A1(n1025), .A2(n1192), .A3(n1186), .A4(n1048), .ZN(n1164) );
XNOR2_X1 U889 ( .A(n1086), .B(n1161), .ZN(G33) );
AND2_X1 U890 ( .A1(n1196), .A2(n1186), .ZN(n1161) );
AND3_X1 U891 ( .A1(n1192), .A2(n1047), .A3(n1025), .ZN(n1196) );
NOR2_X1 U892 ( .A1(n1200), .A2(n1040), .ZN(n1025) );
XNOR2_X1 U893 ( .A(G128), .B(n1165), .ZN(G30) );
NAND4_X1 U894 ( .A1(n1192), .A2(n1185), .A3(n1048), .A4(n1193), .ZN(n1165) );
NOR2_X1 U895 ( .A1(n1034), .A2(n1171), .ZN(n1192) );
XOR2_X1 U896 ( .A(G101), .B(n1201), .Z(G3) );
NOR2_X1 U897 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NOR2_X1 U898 ( .A1(KEYINPUT51), .A2(n1204), .ZN(n1203) );
INV_X1 U899 ( .A(n1205), .ZN(n1204) );
NOR2_X1 U900 ( .A1(KEYINPUT55), .A2(n1205), .ZN(n1202) );
NAND3_X1 U901 ( .A1(n1186), .A2(n1022), .A3(n1206), .ZN(n1205) );
NOR3_X1 U902 ( .A1(n1034), .A2(n1207), .A3(n1208), .ZN(n1206) );
XNOR2_X1 U903 ( .A(n1193), .B(KEYINPUT47), .ZN(n1208) );
XNOR2_X1 U904 ( .A(n1209), .B(n1210), .ZN(G27) );
NOR2_X1 U905 ( .A1(n1211), .A2(n1172), .ZN(n1210) );
NAND4_X1 U906 ( .A1(n1047), .A2(n1035), .A3(n1193), .A4(n1026), .ZN(n1172) );
INV_X1 U907 ( .A(n1212), .ZN(n1035) );
XNOR2_X1 U908 ( .A(n1171), .B(KEYINPUT32), .ZN(n1211) );
AND2_X1 U909 ( .A1(n1213), .A2(n1214), .ZN(n1171) );
NAND4_X1 U910 ( .A1(G953), .A2(G902), .A3(n1021), .A4(n1215), .ZN(n1213) );
INV_X1 U911 ( .A(G900), .ZN(n1215) );
XNOR2_X1 U912 ( .A(G122), .B(n1216), .ZN(G24) );
NAND4_X1 U913 ( .A1(n1064), .A2(n1217), .A3(n1029), .A4(n1218), .ZN(n1216) );
NOR3_X1 U914 ( .A1(n1219), .A2(n1212), .A3(n1188), .ZN(n1218) );
XNOR2_X1 U915 ( .A(KEYINPUT56), .B(n1037), .ZN(n1219) );
AND2_X1 U916 ( .A1(n1220), .A2(n1221), .ZN(n1029) );
XNOR2_X1 U917 ( .A(n1063), .B(KEYINPUT13), .ZN(n1220) );
XNOR2_X1 U918 ( .A(G119), .B(n1222), .ZN(G21) );
NAND3_X1 U919 ( .A1(n1184), .A2(n1185), .A3(n1223), .ZN(n1222) );
XNOR2_X1 U920 ( .A(n1022), .B(KEYINPUT30), .ZN(n1223) );
XOR2_X1 U921 ( .A(n1179), .B(n1224), .Z(G18) );
XNOR2_X1 U922 ( .A(G116), .B(KEYINPUT31), .ZN(n1224) );
NAND3_X1 U923 ( .A1(n1186), .A2(n1048), .A3(n1184), .ZN(n1179) );
AND2_X1 U924 ( .A1(n1225), .A2(n1064), .ZN(n1048) );
XOR2_X1 U925 ( .A(n1178), .B(n1226), .Z(G15) );
XOR2_X1 U926 ( .A(KEYINPUT8), .B(G113), .Z(n1226) );
NAND3_X1 U927 ( .A1(n1184), .A2(n1186), .A3(n1047), .ZN(n1178) );
NOR2_X1 U928 ( .A1(n1188), .A2(n1064), .ZN(n1047) );
XNOR2_X1 U929 ( .A(n1225), .B(KEYINPUT37), .ZN(n1188) );
INV_X1 U930 ( .A(n1050), .ZN(n1186) );
NAND2_X1 U931 ( .A1(n1063), .A2(n1221), .ZN(n1050) );
NOR3_X1 U932 ( .A1(n1037), .A2(n1207), .A3(n1212), .ZN(n1184) );
NAND2_X1 U933 ( .A1(n1053), .A2(n1056), .ZN(n1212) );
XOR2_X1 U934 ( .A(G110), .B(n1227), .Z(G12) );
NOR2_X1 U935 ( .A1(KEYINPUT49), .A2(n1177), .ZN(n1227) );
NAND3_X1 U936 ( .A1(n1180), .A2(n1026), .A3(n1022), .ZN(n1177) );
INV_X1 U937 ( .A(n1055), .ZN(n1022) );
NAND2_X1 U938 ( .A1(n1195), .A2(n1225), .ZN(n1055) );
XOR2_X1 U939 ( .A(n1070), .B(n1228), .Z(n1225) );
XOR2_X1 U940 ( .A(KEYINPUT28), .B(G475), .Z(n1228) );
NAND2_X1 U941 ( .A1(n1109), .A2(n1229), .ZN(n1070) );
XOR2_X1 U942 ( .A(n1230), .B(n1231), .Z(n1109) );
XOR2_X1 U943 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U944 ( .A(n1234), .B(n1086), .ZN(n1233) );
NAND2_X1 U945 ( .A1(KEYINPUT7), .A2(n1235), .ZN(n1234) );
NAND2_X1 U946 ( .A1(n1236), .A2(G214), .ZN(n1232) );
XOR2_X1 U947 ( .A(n1237), .B(n1238), .Z(n1230) );
XOR2_X1 U948 ( .A(n1239), .B(n1081), .Z(n1237) );
INV_X1 U949 ( .A(n1064), .ZN(n1195) );
XNOR2_X1 U950 ( .A(n1240), .B(G478), .ZN(n1064) );
NAND2_X1 U951 ( .A1(n1106), .A2(n1229), .ZN(n1240) );
XOR2_X1 U952 ( .A(n1241), .B(n1242), .Z(n1106) );
XOR2_X1 U953 ( .A(n1243), .B(n1244), .Z(n1242) );
XNOR2_X1 U954 ( .A(n1245), .B(n1246), .ZN(n1244) );
NOR2_X1 U955 ( .A1(KEYINPUT60), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U956 ( .A(G116), .B(G122), .ZN(n1247) );
NAND2_X1 U957 ( .A1(KEYINPUT46), .A2(n1248), .ZN(n1245) );
XNOR2_X1 U958 ( .A(n1249), .B(n1250), .ZN(n1248) );
AND2_X1 U959 ( .A1(n1251), .A2(G217), .ZN(n1243) );
XNOR2_X1 U960 ( .A(G107), .B(n1252), .ZN(n1241) );
XNOR2_X1 U961 ( .A(KEYINPUT43), .B(n1087), .ZN(n1252) );
NAND2_X1 U962 ( .A1(n1253), .A2(n1254), .ZN(n1026) );
OR3_X1 U963 ( .A1(n1221), .A2(n1063), .A3(KEYINPUT13), .ZN(n1254) );
NAND2_X1 U964 ( .A1(KEYINPUT13), .A2(n1185), .ZN(n1253) );
NOR2_X1 U965 ( .A1(n1221), .A2(n1255), .ZN(n1185) );
INV_X1 U966 ( .A(n1063), .ZN(n1255) );
XNOR2_X1 U967 ( .A(n1256), .B(G472), .ZN(n1063) );
NAND2_X1 U968 ( .A1(n1257), .A2(n1229), .ZN(n1256) );
XOR2_X1 U969 ( .A(n1258), .B(n1259), .Z(n1257) );
XNOR2_X1 U970 ( .A(n1122), .B(n1124), .ZN(n1259) );
XOR2_X1 U971 ( .A(n1260), .B(n1261), .Z(n1124) );
XOR2_X1 U972 ( .A(KEYINPUT33), .B(G119), .Z(n1261) );
XNOR2_X1 U973 ( .A(G113), .B(G116), .ZN(n1260) );
XNOR2_X1 U974 ( .A(n1147), .B(n1262), .ZN(n1122) );
XNOR2_X1 U975 ( .A(n1131), .B(G101), .ZN(n1258) );
INV_X1 U976 ( .A(n1128), .ZN(n1131) );
NAND2_X1 U977 ( .A1(n1236), .A2(G210), .ZN(n1128) );
NOR2_X1 U978 ( .A1(G953), .A2(G237), .ZN(n1236) );
NAND3_X1 U979 ( .A1(n1263), .A2(n1264), .A3(n1265), .ZN(n1221) );
NAND2_X1 U980 ( .A1(KEYINPUT10), .A2(n1065), .ZN(n1265) );
NAND3_X1 U981 ( .A1(n1266), .A2(n1267), .A3(n1268), .ZN(n1264) );
INV_X1 U982 ( .A(KEYINPUT10), .ZN(n1267) );
OR2_X1 U983 ( .A1(n1268), .A2(n1266), .ZN(n1263) );
NOR2_X1 U984 ( .A1(n1065), .A2(KEYINPUT52), .ZN(n1266) );
AND2_X1 U985 ( .A1(G217), .A2(n1269), .ZN(n1065) );
XNOR2_X1 U986 ( .A(n1067), .B(KEYINPUT62), .ZN(n1268) );
NOR2_X1 U987 ( .A1(n1100), .A2(n1270), .ZN(n1067) );
XOR2_X1 U988 ( .A(n1271), .B(n1272), .Z(n1100) );
XOR2_X1 U989 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U990 ( .A(n1249), .B(G119), .ZN(n1274) );
INV_X1 U991 ( .A(G128), .ZN(n1249) );
XNOR2_X1 U992 ( .A(n1275), .B(G137), .ZN(n1273) );
INV_X1 U993 ( .A(G146), .ZN(n1275) );
XOR2_X1 U994 ( .A(n1276), .B(n1277), .Z(n1271) );
NOR3_X1 U995 ( .A1(KEYINPUT25), .A2(n1278), .A3(n1279), .ZN(n1277) );
NOR3_X1 U996 ( .A1(KEYINPUT57), .A2(G140), .A3(n1209), .ZN(n1279) );
AND2_X1 U997 ( .A1(n1081), .A2(KEYINPUT57), .ZN(n1278) );
XOR2_X1 U998 ( .A(n1209), .B(G140), .Z(n1081) );
INV_X1 U999 ( .A(G125), .ZN(n1209) );
XOR2_X1 U1000 ( .A(n1280), .B(G110), .Z(n1276) );
NAND2_X1 U1001 ( .A1(n1251), .A2(G221), .ZN(n1280) );
AND2_X1 U1002 ( .A1(G234), .A2(n1019), .ZN(n1251) );
NOR3_X1 U1003 ( .A1(n1034), .A2(n1207), .A3(n1037), .ZN(n1180) );
INV_X1 U1004 ( .A(n1193), .ZN(n1037) );
NOR2_X1 U1005 ( .A1(n1039), .A2(n1040), .ZN(n1193) );
NOR2_X1 U1006 ( .A1(n1281), .A2(n1282), .ZN(n1040) );
INV_X1 U1007 ( .A(G214), .ZN(n1281) );
INV_X1 U1008 ( .A(n1200), .ZN(n1039) );
XNOR2_X1 U1009 ( .A(n1283), .B(n1284), .ZN(n1200) );
NOR2_X1 U1010 ( .A1(n1282), .A2(n1156), .ZN(n1284) );
INV_X1 U1011 ( .A(G210), .ZN(n1156) );
NOR2_X1 U1012 ( .A1(G902), .A2(G237), .ZN(n1282) );
NAND2_X1 U1013 ( .A1(n1285), .A2(n1229), .ZN(n1283) );
XNOR2_X1 U1014 ( .A(n1286), .B(n1092), .ZN(n1285) );
INV_X1 U1015 ( .A(n1152), .ZN(n1092) );
XNOR2_X1 U1016 ( .A(n1287), .B(n1288), .ZN(n1152) );
XOR2_X1 U1017 ( .A(G110), .B(n1289), .Z(n1288) );
XNOR2_X1 U1018 ( .A(KEYINPUT35), .B(n1235), .ZN(n1289) );
INV_X1 U1019 ( .A(G122), .ZN(n1235) );
XOR2_X1 U1020 ( .A(n1290), .B(n1291), .Z(n1287) );
XOR2_X1 U1021 ( .A(n1292), .B(n1238), .Z(n1290) );
XOR2_X1 U1022 ( .A(G104), .B(G113), .Z(n1238) );
NAND2_X1 U1023 ( .A1(n1293), .A2(KEYINPUT45), .ZN(n1292) );
XNOR2_X1 U1024 ( .A(n1294), .B(n1295), .ZN(n1293) );
INV_X1 U1025 ( .A(G116), .ZN(n1295) );
NAND2_X1 U1026 ( .A1(KEYINPUT3), .A2(G119), .ZN(n1294) );
NAND2_X1 U1027 ( .A1(n1296), .A2(n1297), .ZN(n1286) );
NAND2_X1 U1028 ( .A1(n1262), .A2(n1298), .ZN(n1297) );
NAND2_X1 U1029 ( .A1(n1299), .A2(n1190), .ZN(n1296) );
INV_X1 U1030 ( .A(n1262), .ZN(n1190) );
XOR2_X1 U1031 ( .A(n1144), .B(KEYINPUT59), .Z(n1262) );
XNOR2_X1 U1032 ( .A(KEYINPUT2), .B(n1298), .ZN(n1299) );
INV_X1 U1033 ( .A(n1191), .ZN(n1298) );
XOR2_X1 U1034 ( .A(G125), .B(n1300), .Z(n1191) );
AND2_X1 U1035 ( .A1(n1019), .A2(G224), .ZN(n1300) );
INV_X1 U1036 ( .A(n1217), .ZN(n1207) );
NAND2_X1 U1037 ( .A1(n1214), .A2(n1301), .ZN(n1217) );
NAND3_X1 U1038 ( .A1(G902), .A2(n1021), .A3(n1094), .ZN(n1301) );
NOR2_X1 U1039 ( .A1(n1019), .A2(G898), .ZN(n1094) );
NAND3_X1 U1040 ( .A1(n1302), .A2(n1019), .A3(G952), .ZN(n1214) );
XNOR2_X1 U1041 ( .A(KEYINPUT50), .B(n1021), .ZN(n1302) );
NAND2_X1 U1042 ( .A1(G237), .A2(G234), .ZN(n1021) );
NAND2_X1 U1043 ( .A1(n1303), .A2(n1056), .ZN(n1034) );
NAND2_X1 U1044 ( .A1(G221), .A2(n1269), .ZN(n1056) );
NAND2_X1 U1045 ( .A1(G234), .A2(n1304), .ZN(n1269) );
INV_X1 U1046 ( .A(n1053), .ZN(n1303) );
XOR2_X1 U1047 ( .A(n1305), .B(G469), .Z(n1053) );
NAND4_X1 U1048 ( .A1(n1229), .A2(n1306), .A3(n1307), .A4(n1308), .ZN(n1305) );
NAND4_X1 U1049 ( .A1(n1309), .A2(n1310), .A3(KEYINPUT48), .A4(n1311), .ZN(n1308) );
XNOR2_X1 U1050 ( .A(n1312), .B(n1147), .ZN(n1309) );
INV_X1 U1051 ( .A(n1313), .ZN(n1147) );
OR2_X1 U1052 ( .A1(n1311), .A2(n1310), .ZN(n1307) );
INV_X1 U1053 ( .A(KEYINPUT58), .ZN(n1311) );
NAND2_X1 U1054 ( .A1(n1314), .A2(n1315), .ZN(n1306) );
NAND2_X1 U1055 ( .A1(KEYINPUT48), .A2(n1310), .ZN(n1315) );
XOR2_X1 U1056 ( .A(n1316), .B(n1137), .Z(n1310) );
NAND2_X1 U1057 ( .A1(G227), .A2(n1019), .ZN(n1137) );
INV_X1 U1058 ( .A(G953), .ZN(n1019) );
NAND2_X1 U1059 ( .A1(n1317), .A2(n1318), .ZN(n1316) );
NAND2_X1 U1060 ( .A1(G110), .A2(n1150), .ZN(n1318) );
XOR2_X1 U1061 ( .A(KEYINPUT1), .B(n1319), .Z(n1317) );
NOR2_X1 U1062 ( .A1(G110), .A2(n1150), .ZN(n1319) );
INV_X1 U1063 ( .A(G140), .ZN(n1150) );
XNOR2_X1 U1064 ( .A(n1312), .B(n1313), .ZN(n1314) );
XOR2_X1 U1065 ( .A(n1320), .B(n1086), .Z(n1313) );
INV_X1 U1066 ( .A(G131), .ZN(n1086) );
NAND2_X1 U1067 ( .A1(KEYINPUT20), .A2(n1321), .ZN(n1320) );
XNOR2_X1 U1068 ( .A(n1197), .B(n1322), .ZN(n1321) );
NOR2_X1 U1069 ( .A1(KEYINPUT54), .A2(n1087), .ZN(n1322) );
INV_X1 U1070 ( .A(G134), .ZN(n1087) );
INV_X1 U1071 ( .A(G137), .ZN(n1197) );
NAND2_X1 U1072 ( .A1(n1323), .A2(n1324), .ZN(n1312) );
NAND2_X1 U1073 ( .A1(n1143), .A2(n1144), .ZN(n1324) );
XOR2_X1 U1074 ( .A(KEYINPUT42), .B(n1325), .Z(n1323) );
NOR2_X1 U1075 ( .A1(n1144), .A2(n1143), .ZN(n1325) );
XOR2_X1 U1076 ( .A(G104), .B(n1291), .Z(n1143) );
XNOR2_X1 U1077 ( .A(n1326), .B(G101), .ZN(n1291) );
INV_X1 U1078 ( .A(G107), .ZN(n1326) );
XOR2_X1 U1079 ( .A(G128), .B(n1239), .Z(n1144) );
XOR2_X1 U1080 ( .A(G146), .B(n1250), .Z(n1239) );
XOR2_X1 U1081 ( .A(G143), .B(KEYINPUT29), .Z(n1250) );
INV_X1 U1082 ( .A(n1270), .ZN(n1229) );
XOR2_X1 U1083 ( .A(n1304), .B(KEYINPUT61), .Z(n1270) );
INV_X1 U1084 ( .A(G902), .ZN(n1304) );
endmodule


