//Key = 1011011100010001011001110000100000000001101000001011001011111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
n1331, n1332;

XNOR2_X1 U736 ( .A(G107), .B(n1011), .ZN(G9) );
NAND2_X1 U737 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
XOR2_X1 U738 ( .A(KEYINPUT10), .B(n1014), .Z(n1013) );
NAND4_X1 U739 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(G75) );
NAND3_X1 U740 ( .A1(KEYINPUT45), .A2(n1019), .A3(n1020), .ZN(n1018) );
INV_X1 U741 ( .A(G952), .ZN(n1019) );
OR2_X1 U742 ( .A1(n1020), .A2(KEYINPUT45), .ZN(n1017) );
NAND2_X1 U743 ( .A1(G952), .A2(n1021), .ZN(n1015) );
NAND3_X1 U744 ( .A1(n1022), .A2(n1020), .A3(n1023), .ZN(n1021) );
XOR2_X1 U745 ( .A(n1024), .B(KEYINPUT4), .Z(n1023) );
NAND2_X1 U746 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U747 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
NAND3_X1 U748 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
NOR3_X1 U749 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NOR3_X1 U750 ( .A1(n1035), .A2(n1036), .A3(n1014), .ZN(n1034) );
NOR2_X1 U751 ( .A1(n1037), .A2(n1038), .ZN(n1033) );
NAND2_X1 U752 ( .A1(n1039), .A2(n1040), .ZN(n1030) );
NAND4_X1 U753 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1027) );
NOR2_X1 U754 ( .A1(n1045), .A2(n1035), .ZN(n1044) );
INV_X1 U755 ( .A(n1038), .ZN(n1035) );
OR2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1043) );
NAND2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1042) );
NAND2_X1 U758 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NAND3_X1 U759 ( .A1(n1029), .A2(n1052), .A3(n1053), .ZN(n1051) );
NAND2_X1 U760 ( .A1(n1054), .A2(n1032), .ZN(n1041) );
NAND2_X1 U761 ( .A1(n1047), .A2(n1046), .ZN(n1032) );
INV_X1 U762 ( .A(n1055), .ZN(n1025) );
NAND4_X1 U763 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1020) );
NOR4_X1 U764 ( .A1(n1060), .A2(n1039), .A3(n1061), .A4(n1062), .ZN(n1059) );
XOR2_X1 U765 ( .A(n1063), .B(KEYINPUT17), .Z(n1062) );
XOR2_X1 U766 ( .A(n1064), .B(n1065), .Z(n1061) );
NOR2_X1 U767 ( .A1(G472), .A2(KEYINPUT16), .ZN(n1065) );
INV_X1 U768 ( .A(n1052), .ZN(n1060) );
NOR2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(n1058) );
XOR2_X1 U770 ( .A(n1068), .B(KEYINPUT28), .Z(n1066) );
XNOR2_X1 U771 ( .A(n1069), .B(n1070), .ZN(n1056) );
XOR2_X1 U772 ( .A(n1071), .B(n1072), .Z(G72) );
NOR2_X1 U773 ( .A1(n1073), .A2(n1016), .ZN(n1072) );
AND2_X1 U774 ( .A1(G227), .A2(G900), .ZN(n1073) );
NOR2_X1 U775 ( .A1(KEYINPUT55), .A2(n1074), .ZN(n1071) );
XOR2_X1 U776 ( .A(n1075), .B(n1076), .Z(n1074) );
NOR2_X1 U777 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U778 ( .A(n1079), .B(n1080), .Z(n1078) );
XNOR2_X1 U779 ( .A(n1081), .B(n1082), .ZN(n1080) );
NAND2_X1 U780 ( .A1(KEYINPUT2), .A2(n1083), .ZN(n1081) );
XOR2_X1 U781 ( .A(n1084), .B(n1085), .Z(n1083) );
XOR2_X1 U782 ( .A(G134), .B(G131), .Z(n1085) );
NOR2_X1 U783 ( .A1(G137), .A2(KEYINPUT29), .ZN(n1084) );
XOR2_X1 U784 ( .A(KEYINPUT13), .B(n1086), .Z(n1079) );
NOR2_X1 U785 ( .A1(KEYINPUT14), .A2(n1087), .ZN(n1086) );
XOR2_X1 U786 ( .A(G140), .B(G125), .Z(n1087) );
NOR2_X1 U787 ( .A1(G900), .A2(n1016), .ZN(n1077) );
NAND2_X1 U788 ( .A1(n1088), .A2(n1016), .ZN(n1075) );
XOR2_X1 U789 ( .A(KEYINPUT18), .B(n1089), .Z(n1088) );
NOR3_X1 U790 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1089) );
XNOR2_X1 U791 ( .A(KEYINPUT7), .B(n1093), .ZN(n1090) );
XOR2_X1 U792 ( .A(n1094), .B(n1095), .Z(G69) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1016), .ZN(n1095) );
AND2_X1 U794 ( .A1(G224), .A2(G898), .ZN(n1096) );
NAND2_X1 U795 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
NAND2_X1 U796 ( .A1(n1099), .A2(n1016), .ZN(n1098) );
XOR2_X1 U797 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR3_X1 U798 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1100) );
OR3_X1 U799 ( .A1(n1105), .A2(n1101), .A3(n1016), .ZN(n1097) );
XNOR2_X1 U800 ( .A(n1106), .B(n1107), .ZN(n1101) );
NOR2_X1 U801 ( .A1(n1108), .A2(n1109), .ZN(G66) );
XOR2_X1 U802 ( .A(n1110), .B(n1111), .Z(n1109) );
NOR2_X1 U803 ( .A1(n1112), .A2(KEYINPUT9), .ZN(n1111) );
NAND3_X1 U804 ( .A1(G217), .A2(n1113), .A3(n1114), .ZN(n1110) );
NOR2_X1 U805 ( .A1(n1108), .A2(n1115), .ZN(G63) );
XOR2_X1 U806 ( .A(n1116), .B(n1117), .Z(n1115) );
AND2_X1 U807 ( .A1(G478), .A2(n1114), .ZN(n1116) );
NOR2_X1 U808 ( .A1(n1108), .A2(n1118), .ZN(G60) );
XNOR2_X1 U809 ( .A(n1119), .B(n1120), .ZN(n1118) );
AND2_X1 U810 ( .A1(G475), .A2(n1114), .ZN(n1120) );
XNOR2_X1 U811 ( .A(n1103), .B(n1121), .ZN(G6) );
NOR2_X1 U812 ( .A1(G104), .A2(KEYINPUT26), .ZN(n1121) );
NOR2_X1 U813 ( .A1(n1108), .A2(n1122), .ZN(G57) );
XOR2_X1 U814 ( .A(n1123), .B(n1124), .Z(n1122) );
XNOR2_X1 U815 ( .A(G101), .B(n1125), .ZN(n1124) );
XNOR2_X1 U816 ( .A(KEYINPUT62), .B(KEYINPUT46), .ZN(n1125) );
XOR2_X1 U817 ( .A(n1126), .B(n1127), .Z(n1123) );
NOR2_X1 U818 ( .A1(KEYINPUT19), .A2(n1128), .ZN(n1127) );
XOR2_X1 U819 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U820 ( .A(n1131), .B(n1132), .Z(n1129) );
AND2_X1 U821 ( .A1(G472), .A2(n1114), .ZN(n1132) );
NAND2_X1 U822 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
XOR2_X1 U823 ( .A(KEYINPUT63), .B(KEYINPUT1), .Z(n1134) );
XNOR2_X1 U824 ( .A(G113), .B(n1135), .ZN(n1133) );
NOR2_X1 U825 ( .A1(n1108), .A2(n1136), .ZN(G54) );
XOR2_X1 U826 ( .A(n1137), .B(n1138), .Z(n1136) );
XNOR2_X1 U827 ( .A(n1139), .B(n1140), .ZN(n1138) );
NOR3_X1 U828 ( .A1(n1141), .A2(KEYINPUT31), .A3(n1142), .ZN(n1140) );
INV_X1 U829 ( .A(G469), .ZN(n1142) );
NOR2_X1 U830 ( .A1(KEYINPUT53), .A2(n1143), .ZN(n1139) );
XNOR2_X1 U831 ( .A(n1144), .B(n1145), .ZN(n1143) );
XOR2_X1 U832 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND2_X1 U833 ( .A1(n1148), .A2(KEYINPUT56), .ZN(n1146) );
XNOR2_X1 U834 ( .A(n1082), .B(KEYINPUT58), .ZN(n1148) );
NOR3_X1 U835 ( .A1(n1108), .A2(n1149), .A3(n1150), .ZN(G51) );
NOR2_X1 U836 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U837 ( .A(n1153), .B(n1154), .Z(n1151) );
NOR2_X1 U838 ( .A1(KEYINPUT49), .A2(n1155), .ZN(n1153) );
INV_X1 U839 ( .A(n1156), .ZN(n1155) );
NOR2_X1 U840 ( .A1(n1157), .A2(n1158), .ZN(n1149) );
XOR2_X1 U841 ( .A(n1159), .B(n1154), .Z(n1158) );
XOR2_X1 U842 ( .A(n1160), .B(n1161), .Z(n1154) );
NOR2_X1 U843 ( .A1(n1070), .A2(n1141), .ZN(n1161) );
INV_X1 U844 ( .A(n1114), .ZN(n1141) );
NOR2_X1 U845 ( .A1(n1162), .A2(n1022), .ZN(n1114) );
NOR4_X1 U846 ( .A1(n1102), .A2(n1163), .A3(n1092), .A4(n1164), .ZN(n1022) );
OR2_X1 U847 ( .A1(n1093), .A2(n1165), .ZN(n1164) );
XOR2_X1 U848 ( .A(KEYINPUT52), .B(n1091), .Z(n1165) );
NAND4_X1 U849 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1093) );
NAND2_X1 U850 ( .A1(n1170), .A2(n1036), .ZN(n1166) );
NAND3_X1 U851 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1092) );
NAND2_X1 U852 ( .A1(n1174), .A2(n1170), .ZN(n1173) );
INV_X1 U853 ( .A(n1175), .ZN(n1170) );
XOR2_X1 U854 ( .A(n1176), .B(KEYINPUT60), .Z(n1174) );
XNOR2_X1 U855 ( .A(KEYINPUT43), .B(n1177), .ZN(n1163) );
NOR2_X1 U856 ( .A1(n1178), .A2(n1104), .ZN(n1177) );
NAND3_X1 U857 ( .A1(n1179), .A2(n1180), .A3(n1181), .ZN(n1104) );
NAND2_X1 U858 ( .A1(n1012), .A2(n1014), .ZN(n1181) );
XNOR2_X1 U859 ( .A(n1103), .B(KEYINPUT21), .ZN(n1178) );
AND2_X1 U860 ( .A1(n1036), .A2(n1012), .ZN(n1103) );
AND3_X1 U861 ( .A1(n1047), .A2(n1182), .A3(n1183), .ZN(n1012) );
NAND4_X1 U862 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1102) );
XOR2_X1 U863 ( .A(KEYINPUT27), .B(n1188), .Z(n1162) );
NOR2_X1 U864 ( .A1(KEYINPUT49), .A2(n1156), .ZN(n1159) );
XNOR2_X1 U865 ( .A(n1189), .B(n1190), .ZN(n1156) );
NAND2_X1 U866 ( .A1(KEYINPUT5), .A2(G125), .ZN(n1189) );
NOR2_X1 U867 ( .A1(n1016), .A2(G952), .ZN(n1108) );
XOR2_X1 U868 ( .A(G146), .B(n1191), .Z(G48) );
NOR2_X1 U869 ( .A1(n1192), .A2(n1175), .ZN(n1191) );
XOR2_X1 U870 ( .A(n1193), .B(n1167), .Z(G45) );
NAND4_X1 U871 ( .A1(n1194), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1167) );
AND2_X1 U872 ( .A1(n1183), .A2(n1198), .ZN(n1197) );
XNOR2_X1 U873 ( .A(n1199), .B(n1168), .ZN(G42) );
NAND2_X1 U874 ( .A1(n1200), .A2(n1201), .ZN(n1168) );
XOR2_X1 U875 ( .A(n1202), .B(KEYINPUT22), .Z(n1199) );
XNOR2_X1 U876 ( .A(G137), .B(n1169), .ZN(G39) );
NAND2_X1 U877 ( .A1(n1201), .A2(n1203), .ZN(n1169) );
XOR2_X1 U878 ( .A(G134), .B(n1091), .Z(G36) );
AND3_X1 U879 ( .A1(n1201), .A2(n1014), .A3(n1198), .ZN(n1091) );
XNOR2_X1 U880 ( .A(n1171), .B(n1204), .ZN(G33) );
NOR2_X1 U881 ( .A1(KEYINPUT36), .A2(n1205), .ZN(n1204) );
INV_X1 U882 ( .A(G131), .ZN(n1205) );
NAND3_X1 U883 ( .A1(n1036), .A2(n1201), .A3(n1198), .ZN(n1171) );
AND4_X1 U884 ( .A1(n1046), .A2(n1040), .A3(n1206), .A4(n1029), .ZN(n1201) );
NOR2_X1 U885 ( .A1(n1039), .A2(n1207), .ZN(n1206) );
XOR2_X1 U886 ( .A(G128), .B(n1208), .Z(G30) );
NOR2_X1 U887 ( .A1(n1176), .A2(n1175), .ZN(n1208) );
NAND4_X1 U888 ( .A1(n1183), .A2(n1209), .A3(n1195), .A4(n1067), .ZN(n1175) );
XNOR2_X1 U889 ( .A(G101), .B(n1179), .ZN(G3) );
NAND2_X1 U890 ( .A1(n1210), .A2(n1198), .ZN(n1179) );
XNOR2_X1 U891 ( .A(G125), .B(n1172), .ZN(G27) );
NAND3_X1 U892 ( .A1(n1038), .A2(n1200), .A3(n1211), .ZN(n1172) );
NOR3_X1 U893 ( .A1(n1029), .A2(n1207), .A3(n1212), .ZN(n1211) );
INV_X1 U894 ( .A(n1195), .ZN(n1207) );
NAND2_X1 U895 ( .A1(n1055), .A2(n1213), .ZN(n1195) );
NAND4_X1 U896 ( .A1(G953), .A2(G902), .A3(n1214), .A4(n1215), .ZN(n1213) );
INV_X1 U897 ( .A(G900), .ZN(n1215) );
NOR3_X1 U898 ( .A1(n1209), .A2(n1053), .A3(n1192), .ZN(n1200) );
XNOR2_X1 U899 ( .A(G122), .B(n1184), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1216), .A2(n1047), .A3(n1196), .A4(n1194), .ZN(n1184) );
NOR2_X1 U901 ( .A1(n1067), .A2(n1209), .ZN(n1047) );
XNOR2_X1 U902 ( .A(n1185), .B(n1217), .ZN(G21) );
NOR2_X1 U903 ( .A1(KEYINPUT30), .A2(n1218), .ZN(n1217) );
NAND2_X1 U904 ( .A1(n1216), .A2(n1203), .ZN(n1185) );
NOR3_X1 U905 ( .A1(n1050), .A2(n1053), .A3(n1045), .ZN(n1203) );
NAND2_X1 U906 ( .A1(n1219), .A2(n1220), .ZN(G18) );
NAND2_X1 U907 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
INV_X1 U908 ( .A(G116), .ZN(n1222) );
XNOR2_X1 U909 ( .A(KEYINPUT47), .B(n1186), .ZN(n1221) );
NAND2_X1 U910 ( .A1(n1223), .A2(G116), .ZN(n1219) );
XNOR2_X1 U911 ( .A(KEYINPUT15), .B(n1186), .ZN(n1223) );
NAND3_X1 U912 ( .A1(n1198), .A2(n1014), .A3(n1216), .ZN(n1186) );
INV_X1 U913 ( .A(n1176), .ZN(n1014) );
NAND2_X1 U914 ( .A1(n1057), .A2(n1196), .ZN(n1176) );
INV_X1 U915 ( .A(n1063), .ZN(n1196) );
XNOR2_X1 U916 ( .A(G113), .B(n1187), .ZN(G15) );
NAND3_X1 U917 ( .A1(n1198), .A2(n1036), .A3(n1216), .ZN(n1187) );
AND4_X1 U918 ( .A1(n1054), .A2(n1038), .A3(n1046), .A4(n1182), .ZN(n1216) );
INV_X1 U919 ( .A(n1212), .ZN(n1046) );
NOR2_X1 U920 ( .A1(n1040), .A2(n1039), .ZN(n1038) );
INV_X1 U921 ( .A(n1068), .ZN(n1040) );
INV_X1 U922 ( .A(n1192), .ZN(n1036) );
NAND2_X1 U923 ( .A1(n1063), .A2(n1194), .ZN(n1192) );
INV_X1 U924 ( .A(n1057), .ZN(n1194) );
INV_X1 U925 ( .A(n1049), .ZN(n1198) );
NAND2_X1 U926 ( .A1(n1053), .A2(n1209), .ZN(n1049) );
INV_X1 U927 ( .A(n1050), .ZN(n1209) );
INV_X1 U928 ( .A(n1067), .ZN(n1053) );
XOR2_X1 U929 ( .A(n1224), .B(n1180), .Z(G12) );
NAND3_X1 U930 ( .A1(n1050), .A2(n1067), .A3(n1210), .ZN(n1180) );
AND3_X1 U931 ( .A1(n1183), .A2(n1182), .A3(n1037), .ZN(n1210) );
INV_X1 U932 ( .A(n1045), .ZN(n1037) );
NAND2_X1 U933 ( .A1(n1063), .A2(n1057), .ZN(n1045) );
XOR2_X1 U934 ( .A(n1225), .B(n1226), .Z(n1057) );
XOR2_X1 U935 ( .A(KEYINPUT33), .B(G475), .Z(n1226) );
NAND2_X1 U936 ( .A1(n1119), .A2(n1188), .ZN(n1225) );
XNOR2_X1 U937 ( .A(n1227), .B(n1228), .ZN(n1119) );
XOR2_X1 U938 ( .A(G122), .B(G113), .Z(n1228) );
XNOR2_X1 U939 ( .A(n1229), .B(n1230), .ZN(n1227) );
NOR2_X1 U940 ( .A1(G104), .A2(KEYINPUT44), .ZN(n1230) );
NOR2_X1 U941 ( .A1(KEYINPUT38), .A2(n1231), .ZN(n1229) );
XOR2_X1 U942 ( .A(n1232), .B(n1233), .Z(n1231) );
XOR2_X1 U943 ( .A(n1234), .B(n1235), .Z(n1233) );
NOR2_X1 U944 ( .A1(G131), .A2(KEYINPUT35), .ZN(n1235) );
NAND2_X1 U945 ( .A1(n1236), .A2(n1237), .ZN(n1234) );
XOR2_X1 U946 ( .A(n1238), .B(KEYINPUT32), .Z(n1236) );
XOR2_X1 U947 ( .A(n1239), .B(n1240), .Z(n1232) );
NAND2_X1 U948 ( .A1(n1241), .A2(G214), .ZN(n1239) );
XOR2_X1 U949 ( .A(n1242), .B(G478), .Z(n1063) );
OR2_X1 U950 ( .A1(n1117), .A2(G902), .ZN(n1242) );
XNOR2_X1 U951 ( .A(n1243), .B(n1244), .ZN(n1117) );
XOR2_X1 U952 ( .A(G116), .B(n1245), .Z(n1244) );
XOR2_X1 U953 ( .A(G134), .B(G122), .Z(n1245) );
XOR2_X1 U954 ( .A(n1246), .B(n1247), .Z(n1243) );
NOR2_X1 U955 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
XOR2_X1 U956 ( .A(n1250), .B(G107), .Z(n1246) );
NAND2_X1 U957 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U958 ( .A1(G143), .A2(n1253), .ZN(n1252) );
XOR2_X1 U959 ( .A(KEYINPUT48), .B(n1254), .Z(n1251) );
NOR2_X1 U960 ( .A1(G143), .A2(n1253), .ZN(n1254) );
NAND2_X1 U961 ( .A1(n1055), .A2(n1255), .ZN(n1182) );
NAND4_X1 U962 ( .A1(G953), .A2(G902), .A3(n1214), .A4(n1105), .ZN(n1255) );
INV_X1 U963 ( .A(G898), .ZN(n1105) );
NAND3_X1 U964 ( .A1(n1214), .A2(n1016), .A3(G952), .ZN(n1055) );
NAND2_X1 U965 ( .A1(G237), .A2(G234), .ZN(n1214) );
NOR4_X1 U966 ( .A1(n1029), .A2(n1212), .A3(n1068), .A4(n1039), .ZN(n1183) );
AND2_X1 U967 ( .A1(G221), .A2(n1113), .ZN(n1039) );
NAND2_X1 U968 ( .A1(G234), .A2(n1188), .ZN(n1113) );
XOR2_X1 U969 ( .A(n1256), .B(n1257), .Z(n1068) );
XOR2_X1 U970 ( .A(KEYINPUT8), .B(G469), .Z(n1257) );
NAND2_X1 U971 ( .A1(n1258), .A2(n1188), .ZN(n1256) );
XOR2_X1 U972 ( .A(n1259), .B(n1260), .Z(n1258) );
INV_X1 U973 ( .A(n1137), .ZN(n1260) );
XOR2_X1 U974 ( .A(n1261), .B(n1262), .Z(n1137) );
XOR2_X1 U975 ( .A(G140), .B(G110), .Z(n1262) );
NAND2_X1 U976 ( .A1(G227), .A2(n1016), .ZN(n1261) );
XOR2_X1 U977 ( .A(n1263), .B(n1264), .Z(n1259) );
INV_X1 U978 ( .A(n1147), .ZN(n1264) );
NAND2_X1 U979 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
NAND2_X1 U980 ( .A1(n1144), .A2(n1082), .ZN(n1266) );
XOR2_X1 U981 ( .A(KEYINPUT59), .B(n1267), .Z(n1265) );
NOR2_X1 U982 ( .A1(n1144), .A2(n1082), .ZN(n1267) );
XNOR2_X1 U983 ( .A(n1253), .B(n1240), .ZN(n1082) );
XOR2_X1 U984 ( .A(G146), .B(G143), .Z(n1240) );
NAND2_X1 U985 ( .A1(n1268), .A2(n1269), .ZN(n1144) );
NAND2_X1 U986 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
INV_X1 U987 ( .A(KEYINPUT34), .ZN(n1271) );
XOR2_X1 U988 ( .A(G101), .B(n1272), .Z(n1270) );
NAND3_X1 U989 ( .A1(G101), .A2(n1272), .A3(KEYINPUT34), .ZN(n1268) );
XOR2_X1 U990 ( .A(n1052), .B(KEYINPUT23), .Z(n1212) );
NAND2_X1 U991 ( .A1(G214), .A2(n1273), .ZN(n1052) );
INV_X1 U992 ( .A(n1054), .ZN(n1029) );
XNOR2_X1 U993 ( .A(n1274), .B(n1069), .ZN(n1054) );
NAND2_X1 U994 ( .A1(n1275), .A2(n1188), .ZN(n1069) );
XOR2_X1 U995 ( .A(n1276), .B(n1277), .Z(n1275) );
XOR2_X1 U996 ( .A(n1157), .B(n1278), .Z(n1277) );
XOR2_X1 U997 ( .A(KEYINPUT6), .B(G125), .Z(n1278) );
INV_X1 U998 ( .A(n1152), .ZN(n1157) );
NAND2_X1 U999 ( .A1(G224), .A2(n1016), .ZN(n1152) );
XOR2_X1 U1000 ( .A(n1190), .B(n1160), .Z(n1276) );
XNOR2_X1 U1001 ( .A(n1279), .B(n1280), .ZN(n1160) );
XOR2_X1 U1002 ( .A(KEYINPUT50), .B(n1107), .Z(n1280) );
AND2_X1 U1003 ( .A1(n1281), .A2(n1282), .ZN(n1107) );
OR2_X1 U1004 ( .A1(n1224), .A2(G122), .ZN(n1282) );
XOR2_X1 U1005 ( .A(n1283), .B(KEYINPUT25), .Z(n1281) );
NAND2_X1 U1006 ( .A1(G122), .A2(n1224), .ZN(n1283) );
NAND2_X1 U1007 ( .A1(KEYINPUT54), .A2(n1106), .ZN(n1279) );
XOR2_X1 U1008 ( .A(n1284), .B(n1285), .Z(n1106) );
XOR2_X1 U1009 ( .A(G119), .B(n1286), .Z(n1285) );
NOR2_X1 U1010 ( .A1(G116), .A2(KEYINPUT37), .ZN(n1286) );
XNOR2_X1 U1011 ( .A(n1272), .B(n1287), .ZN(n1284) );
XOR2_X1 U1012 ( .A(G104), .B(n1288), .Z(n1272) );
XOR2_X1 U1013 ( .A(KEYINPUT20), .B(G107), .Z(n1288) );
NAND2_X1 U1014 ( .A1(KEYINPUT40), .A2(n1070), .ZN(n1274) );
NAND2_X1 U1015 ( .A1(G210), .A2(n1273), .ZN(n1070) );
NAND2_X1 U1016 ( .A1(n1289), .A2(n1188), .ZN(n1273) );
XOR2_X1 U1017 ( .A(KEYINPUT0), .B(G237), .Z(n1289) );
NAND3_X1 U1018 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1067) );
NAND2_X1 U1019 ( .A1(n1112), .A2(n1293), .ZN(n1292) );
OR3_X1 U1020 ( .A1(n1293), .A2(n1112), .A3(G902), .ZN(n1291) );
AND2_X1 U1021 ( .A1(n1294), .A2(n1295), .ZN(n1112) );
NAND2_X1 U1022 ( .A1(n1296), .A2(n1297), .ZN(n1295) );
XOR2_X1 U1023 ( .A(KEYINPUT42), .B(n1298), .Z(n1294) );
NOR2_X1 U1024 ( .A1(n1296), .A2(n1297), .ZN(n1298) );
XOR2_X1 U1025 ( .A(n1299), .B(n1300), .Z(n1297) );
XOR2_X1 U1026 ( .A(n1224), .B(n1301), .Z(n1300) );
NAND3_X1 U1027 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1301) );
NAND2_X1 U1028 ( .A1(G146), .A2(n1305), .ZN(n1304) );
NAND2_X1 U1029 ( .A1(KEYINPUT24), .A2(n1306), .ZN(n1303) );
NAND2_X1 U1030 ( .A1(n1307), .A2(n1308), .ZN(n1306) );
XOR2_X1 U1031 ( .A(KEYINPUT3), .B(G146), .Z(n1308) );
NAND2_X1 U1032 ( .A1(n1309), .A2(n1310), .ZN(n1302) );
INV_X1 U1033 ( .A(KEYINPUT24), .ZN(n1310) );
NAND2_X1 U1034 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
NAND3_X1 U1035 ( .A1(KEYINPUT3), .A2(n1307), .A3(n1313), .ZN(n1312) );
INV_X1 U1036 ( .A(n1305), .ZN(n1307) );
NAND2_X1 U1037 ( .A1(n1237), .A2(n1238), .ZN(n1305) );
NAND2_X1 U1038 ( .A1(n1314), .A2(G125), .ZN(n1238) );
OR2_X1 U1039 ( .A1(n1314), .A2(G125), .ZN(n1237) );
XOR2_X1 U1040 ( .A(n1202), .B(KEYINPUT41), .Z(n1314) );
INV_X1 U1041 ( .A(G140), .ZN(n1202) );
OR2_X1 U1042 ( .A1(n1313), .A2(KEYINPUT3), .ZN(n1311) );
INV_X1 U1043 ( .A(G146), .ZN(n1313) );
XOR2_X1 U1044 ( .A(n1218), .B(G128), .Z(n1299) );
AND2_X1 U1045 ( .A1(n1315), .A2(n1316), .ZN(n1296) );
NAND3_X1 U1046 ( .A1(G137), .A2(G221), .A3(n1317), .ZN(n1316) );
NAND2_X1 U1047 ( .A1(n1318), .A2(n1319), .ZN(n1315) );
NAND2_X1 U1048 ( .A1(n1317), .A2(G221), .ZN(n1319) );
INV_X1 U1049 ( .A(n1249), .ZN(n1317) );
NAND2_X1 U1050 ( .A1(G234), .A2(n1016), .ZN(n1249) );
INV_X1 U1051 ( .A(G953), .ZN(n1016) );
XOR2_X1 U1052 ( .A(KEYINPUT61), .B(G137), .Z(n1318) );
NOR2_X1 U1053 ( .A1(n1248), .A2(G234), .ZN(n1293) );
INV_X1 U1054 ( .A(G217), .ZN(n1248) );
NAND2_X1 U1055 ( .A1(G217), .A2(G902), .ZN(n1290) );
XOR2_X1 U1056 ( .A(n1064), .B(G472), .Z(n1050) );
NAND2_X1 U1057 ( .A1(n1320), .A2(n1188), .ZN(n1064) );
INV_X1 U1058 ( .A(G902), .ZN(n1188) );
XOR2_X1 U1059 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1060 ( .A(n1130), .B(n1135), .ZN(n1322) );
XOR2_X1 U1061 ( .A(G116), .B(n1323), .Z(n1135) );
NOR2_X1 U1062 ( .A1(KEYINPUT12), .A2(n1324), .ZN(n1323) );
XOR2_X1 U1063 ( .A(n1218), .B(KEYINPUT51), .Z(n1324) );
INV_X1 U1064 ( .A(G119), .ZN(n1218) );
XOR2_X1 U1065 ( .A(n1147), .B(n1190), .Z(n1130) );
XOR2_X1 U1066 ( .A(n1325), .B(n1326), .Z(n1190) );
NOR2_X1 U1067 ( .A1(n1327), .A2(n1328), .ZN(n1326) );
XOR2_X1 U1068 ( .A(n1329), .B(KEYINPUT39), .Z(n1328) );
NAND2_X1 U1069 ( .A1(G146), .A2(n1193), .ZN(n1329) );
NOR2_X1 U1070 ( .A1(G146), .A2(n1193), .ZN(n1327) );
INV_X1 U1071 ( .A(G143), .ZN(n1193) );
NAND2_X1 U1072 ( .A1(KEYINPUT11), .A2(n1253), .ZN(n1325) );
INV_X1 U1073 ( .A(G128), .ZN(n1253) );
XOR2_X1 U1074 ( .A(n1330), .B(n1331), .Z(n1147) );
XOR2_X1 U1075 ( .A(G137), .B(G131), .Z(n1331) );
NAND2_X1 U1076 ( .A1(KEYINPUT57), .A2(n1332), .ZN(n1330) );
INV_X1 U1077 ( .A(G134), .ZN(n1332) );
XOR2_X1 U1078 ( .A(n1126), .B(n1287), .Z(n1321) );
XOR2_X1 U1079 ( .A(G101), .B(G113), .Z(n1287) );
NAND2_X1 U1080 ( .A1(n1241), .A2(G210), .ZN(n1126) );
NOR2_X1 U1081 ( .A1(G953), .A2(G237), .ZN(n1241) );
INV_X1 U1082 ( .A(G110), .ZN(n1224) );
endmodule


