//Key = 0101111110010110010001101001011010000101110001000111011000100110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313;

XNOR2_X1 U721 ( .A(G107), .B(n998), .ZN(G9) );
NOR2_X1 U722 ( .A1(n999), .A2(n1000), .ZN(G75) );
NOR4_X1 U723 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n1000) );
NOR2_X1 U724 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
NAND4_X1 U725 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1001) );
NAND3_X1 U726 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n1008) );
NAND2_X1 U727 ( .A1(n1014), .A2(n1015), .ZN(n1012) );
NAND3_X1 U728 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n1015) );
OR2_X1 U729 ( .A1(n1019), .A2(n1020), .ZN(n1017) );
NAND2_X1 U730 ( .A1(n1021), .A2(n1022), .ZN(n1014) );
NAND3_X1 U731 ( .A1(n1023), .A2(n1024), .A3(n1025), .ZN(n1022) );
NAND2_X1 U732 ( .A1(n1016), .A2(n1026), .ZN(n1025) );
NAND3_X1 U733 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1024) );
XNOR2_X1 U734 ( .A(n1016), .B(KEYINPUT21), .ZN(n1029) );
NAND2_X1 U735 ( .A1(n1018), .A2(n1030), .ZN(n1023) );
OR2_X1 U736 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND3_X1 U737 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1007) );
XOR2_X1 U738 ( .A(n1006), .B(KEYINPUT39), .Z(n1035) );
NAND4_X1 U739 ( .A1(n1013), .A2(n1018), .A3(n1016), .A4(n1021), .ZN(n1006) );
INV_X1 U740 ( .A(n1036), .ZN(n1013) );
NOR3_X1 U741 ( .A1(n1037), .A2(G953), .A3(n1038), .ZN(n999) );
INV_X1 U742 ( .A(n1009), .ZN(n1038) );
NAND4_X1 U743 ( .A1(n1039), .A2(n1040), .A3(n1041), .A4(n1042), .ZN(n1009) );
NOR4_X1 U744 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
AND3_X1 U745 ( .A1(KEYINPUT4), .A2(n1047), .A3(n1048), .ZN(n1046) );
NOR2_X1 U746 ( .A1(KEYINPUT4), .A2(n1048), .ZN(n1045) );
XNOR2_X1 U747 ( .A(KEYINPUT12), .B(n1033), .ZN(n1044) );
NAND3_X1 U748 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1043) );
XNOR2_X1 U749 ( .A(G472), .B(n1052), .ZN(n1051) );
NAND2_X1 U750 ( .A1(KEYINPUT22), .A2(n1053), .ZN(n1052) );
NAND2_X1 U751 ( .A1(n1054), .A2(n1055), .ZN(n1050) );
XOR2_X1 U752 ( .A(KEYINPUT11), .B(n1056), .Z(n1049) );
NOR2_X1 U753 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
XNOR2_X1 U754 ( .A(n1057), .B(KEYINPUT35), .ZN(n1054) );
NOR3_X1 U755 ( .A1(n1058), .A2(n1034), .A3(n1028), .ZN(n1041) );
NOR3_X1 U756 ( .A1(n1059), .A2(n1060), .A3(n1061), .ZN(n1058) );
INV_X1 U757 ( .A(KEYINPUT62), .ZN(n1059) );
NAND2_X1 U758 ( .A1(n1062), .A2(n1063), .ZN(n1040) );
NAND3_X1 U759 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1062) );
NAND2_X1 U760 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U761 ( .A1(n1069), .A2(n1070), .ZN(n1065) );
NAND2_X1 U762 ( .A1(KEYINPUT62), .A2(G478), .ZN(n1070) );
INV_X1 U763 ( .A(n1071), .ZN(n1069) );
NAND2_X1 U764 ( .A1(n1072), .A2(n1073), .ZN(n1064) );
OR2_X1 U765 ( .A1(n1073), .A2(n1074), .ZN(n1039) );
XOR2_X1 U766 ( .A(G475), .B(KEYINPUT24), .Z(n1073) );
XNOR2_X1 U767 ( .A(KEYINPUT44), .B(n1004), .ZN(n1037) );
XOR2_X1 U768 ( .A(n1075), .B(n1076), .Z(G72) );
XOR2_X1 U769 ( .A(n1077), .B(n1078), .Z(n1076) );
NOR2_X1 U770 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
XNOR2_X1 U771 ( .A(G953), .B(KEYINPUT25), .ZN(n1080) );
AND2_X1 U772 ( .A1(G227), .A2(G900), .ZN(n1079) );
NAND2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1077) );
XNOR2_X1 U774 ( .A(KEYINPUT50), .B(n1010), .ZN(n1081) );
NAND3_X1 U775 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1075) );
XOR2_X1 U776 ( .A(n1086), .B(KEYINPUT33), .Z(n1085) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
INV_X1 U778 ( .A(n1089), .ZN(n1088) );
XNOR2_X1 U779 ( .A(n1090), .B(n1091), .ZN(n1087) );
INV_X1 U780 ( .A(n1092), .ZN(n1084) );
NAND2_X1 U781 ( .A1(n1093), .A2(n1089), .ZN(n1083) );
XOR2_X1 U782 ( .A(G140), .B(n1094), .Z(n1089) );
XNOR2_X1 U783 ( .A(n1095), .B(n1091), .ZN(n1093) );
XNOR2_X1 U784 ( .A(n1096), .B(KEYINPUT43), .ZN(n1091) );
NAND2_X1 U785 ( .A1(KEYINPUT6), .A2(n1097), .ZN(n1096) );
XOR2_X1 U786 ( .A(n1098), .B(n1099), .Z(G69) );
XOR2_X1 U787 ( .A(n1100), .B(n1101), .Z(n1099) );
NOR2_X1 U788 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U789 ( .A(n1104), .B(n1105), .Z(n1103) );
XOR2_X1 U790 ( .A(KEYINPUT42), .B(n1106), .Z(n1105) );
XNOR2_X1 U791 ( .A(n1107), .B(n1108), .ZN(n1104) );
NOR2_X1 U792 ( .A1(G953), .A2(n1109), .ZN(n1100) );
NOR2_X1 U793 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
XOR2_X1 U794 ( .A(n1112), .B(KEYINPUT28), .Z(n1110) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1010), .ZN(n1098) );
AND2_X1 U796 ( .A1(G224), .A2(G898), .ZN(n1113) );
NOR2_X1 U797 ( .A1(n1114), .A2(n1115), .ZN(G66) );
XOR2_X1 U798 ( .A(n1116), .B(n1067), .Z(n1115) );
NAND2_X1 U799 ( .A1(n1117), .A2(n1048), .ZN(n1116) );
INV_X1 U800 ( .A(n1068), .ZN(n1048) );
NOR2_X1 U801 ( .A1(n1114), .A2(n1118), .ZN(G63) );
NOR2_X1 U802 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1121), .B(KEYINPUT54), .Z(n1120) );
NAND2_X1 U804 ( .A1(n1122), .A2(n1071), .ZN(n1121) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1071), .ZN(n1119) );
NOR2_X1 U806 ( .A1(n1123), .A2(n1061), .ZN(n1122) );
NOR3_X1 U807 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(G60) );
NOR3_X1 U808 ( .A1(n1127), .A2(G952), .A3(n1128), .ZN(n1126) );
INV_X1 U809 ( .A(KEYINPUT63), .ZN(n1127) );
NOR2_X1 U810 ( .A1(KEYINPUT63), .A2(n1129), .ZN(n1125) );
XOR2_X1 U811 ( .A(n1130), .B(n1072), .Z(n1124) );
NAND2_X1 U812 ( .A1(n1117), .A2(G475), .ZN(n1130) );
XNOR2_X1 U813 ( .A(n1131), .B(n1132), .ZN(G6) );
NOR2_X1 U814 ( .A1(n1005), .A2(n1133), .ZN(n1132) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1135), .ZN(G57) );
XNOR2_X1 U816 ( .A(KEYINPUT55), .B(n1129), .ZN(n1135) );
XOR2_X1 U817 ( .A(n1136), .B(n1137), .Z(n1134) );
XOR2_X1 U818 ( .A(n1138), .B(n1139), .Z(n1137) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(n1136) );
NAND2_X1 U820 ( .A1(n1117), .A2(G472), .ZN(n1141) );
NAND2_X1 U821 ( .A1(KEYINPUT14), .A2(n1142), .ZN(n1140) );
XOR2_X1 U822 ( .A(KEYINPUT27), .B(n1143), .Z(n1142) );
NOR2_X1 U823 ( .A1(n1114), .A2(n1144), .ZN(G54) );
XOR2_X1 U824 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U825 ( .A(n1138), .B(n1147), .Z(n1146) );
XNOR2_X1 U826 ( .A(n1148), .B(n1149), .ZN(n1147) );
NOR3_X1 U827 ( .A1(n1123), .A2(KEYINPUT31), .A3(n1057), .ZN(n1148) );
INV_X1 U828 ( .A(n1117), .ZN(n1123) );
NOR2_X1 U829 ( .A1(n1063), .A2(n1150), .ZN(n1117) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1145) );
XOR2_X1 U831 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U832 ( .A1(KEYINPUT23), .A2(n1155), .ZN(n1154) );
XNOR2_X1 U833 ( .A(KEYINPUT34), .B(n1156), .ZN(n1155) );
XNOR2_X1 U834 ( .A(KEYINPUT40), .B(n1157), .ZN(n1151) );
NOR2_X1 U835 ( .A1(n1114), .A2(n1158), .ZN(G51) );
XOR2_X1 U836 ( .A(n1159), .B(n1160), .Z(n1158) );
XNOR2_X1 U837 ( .A(n1161), .B(n1162), .ZN(n1160) );
NAND3_X1 U838 ( .A1(n1163), .A2(n1164), .A3(G902), .ZN(n1161) );
XNOR2_X1 U839 ( .A(KEYINPUT3), .B(n1002), .ZN(n1164) );
INV_X1 U840 ( .A(n1150), .ZN(n1002) );
NOR4_X1 U841 ( .A1(n1112), .A2(n1111), .A3(n1165), .A4(n1166), .ZN(n1150) );
AND2_X1 U842 ( .A1(n1082), .A2(n1167), .ZN(n1166) );
NAND4_X1 U843 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1082) );
NOR4_X1 U844 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1171) );
NOR2_X1 U845 ( .A1(n1176), .A2(n1177), .ZN(n1170) );
INV_X1 U846 ( .A(n1178), .ZN(n1177) );
NOR2_X1 U847 ( .A1(n1167), .A2(n1176), .ZN(n1165) );
NOR2_X1 U848 ( .A1(n1179), .A2(n1180), .ZN(n1176) );
XNOR2_X1 U849 ( .A(n1181), .B(KEYINPUT10), .ZN(n1179) );
INV_X1 U850 ( .A(KEYINPUT20), .ZN(n1167) );
NAND4_X1 U851 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1111) );
NAND2_X1 U852 ( .A1(KEYINPUT32), .A2(n1186), .ZN(n1183) );
NOR2_X1 U853 ( .A1(n1187), .A2(n1188), .ZN(n1182) );
NOR2_X1 U854 ( .A1(n1005), .A2(n1189), .ZN(n1188) );
XOR2_X1 U855 ( .A(n1190), .B(KEYINPUT9), .Z(n1189) );
NOR4_X1 U856 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1187) );
NAND3_X1 U857 ( .A1(n1195), .A2(n1196), .A3(n1032), .ZN(n1192) );
INV_X1 U858 ( .A(KEYINPUT32), .ZN(n1196) );
NAND4_X1 U859 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n998), .ZN(n1112) );
NAND3_X1 U860 ( .A1(n1032), .A2(n1200), .A3(n1021), .ZN(n998) );
NAND2_X1 U861 ( .A1(n1201), .A2(n1191), .ZN(n1197) );
XOR2_X1 U862 ( .A(n1133), .B(KEYINPUT49), .Z(n1201) );
NAND4_X1 U863 ( .A1(n1031), .A2(n1021), .A3(n1026), .A4(n1195), .ZN(n1133) );
INV_X1 U864 ( .A(n1129), .ZN(n1114) );
NAND2_X1 U865 ( .A1(n1128), .A2(n1004), .ZN(n1129) );
INV_X1 U866 ( .A(G952), .ZN(n1004) );
XNOR2_X1 U867 ( .A(G953), .B(KEYINPUT61), .ZN(n1128) );
XNOR2_X1 U868 ( .A(G146), .B(n1168), .ZN(G48) );
NAND3_X1 U869 ( .A1(n1031), .A2(n1191), .A3(n1202), .ZN(n1168) );
XNOR2_X1 U870 ( .A(G143), .B(n1169), .ZN(G45) );
NAND4_X1 U871 ( .A1(n1203), .A2(n1204), .A3(n1191), .A4(n1205), .ZN(n1169) );
XNOR2_X1 U872 ( .A(n1156), .B(n1206), .ZN(G42) );
NOR2_X1 U873 ( .A1(n1207), .A2(n1180), .ZN(n1206) );
NAND4_X1 U874 ( .A1(n1011), .A2(n1031), .A3(n1019), .A4(n1026), .ZN(n1180) );
XOR2_X1 U875 ( .A(G137), .B(n1175), .Z(G39) );
AND3_X1 U876 ( .A1(n1011), .A2(n1016), .A3(n1202), .ZN(n1175) );
XOR2_X1 U877 ( .A(n1208), .B(n1209), .Z(G36) );
XOR2_X1 U878 ( .A(KEYINPUT60), .B(G134), .Z(n1209) );
NOR2_X1 U879 ( .A1(KEYINPUT2), .A2(n1178), .ZN(n1208) );
NAND3_X1 U880 ( .A1(n1011), .A2(n1032), .A3(n1204), .ZN(n1178) );
XOR2_X1 U881 ( .A(G131), .B(n1174), .Z(G33) );
AND3_X1 U882 ( .A1(n1011), .A2(n1031), .A3(n1204), .ZN(n1174) );
AND3_X1 U883 ( .A1(n1026), .A2(n1181), .A3(n1020), .ZN(n1204) );
AND2_X1 U884 ( .A1(n1210), .A2(n1033), .ZN(n1011) );
XNOR2_X1 U885 ( .A(n1034), .B(KEYINPUT56), .ZN(n1210) );
XNOR2_X1 U886 ( .A(n1211), .B(n1173), .ZN(G30) );
AND3_X1 U887 ( .A1(n1032), .A2(n1191), .A3(n1202), .ZN(n1173) );
AND4_X1 U888 ( .A1(n1026), .A2(n1212), .A3(n1213), .A4(n1181), .ZN(n1202) );
NAND2_X1 U889 ( .A1(n1214), .A2(n1215), .ZN(G3) );
NAND2_X1 U890 ( .A1(G101), .A2(n1198), .ZN(n1215) );
XOR2_X1 U891 ( .A(n1216), .B(KEYINPUT47), .Z(n1214) );
OR2_X1 U892 ( .A1(n1198), .A2(G101), .ZN(n1216) );
NAND3_X1 U893 ( .A1(n1016), .A2(n1200), .A3(n1020), .ZN(n1198) );
INV_X1 U894 ( .A(n1193), .ZN(n1020) );
NAND2_X1 U895 ( .A1(n1217), .A2(n1213), .ZN(n1193) );
XOR2_X1 U896 ( .A(G125), .B(n1172), .Z(G27) );
AND4_X1 U897 ( .A1(n1018), .A2(n1031), .A3(n1218), .A4(n1019), .ZN(n1172) );
NOR2_X1 U898 ( .A1(n1207), .A2(n1005), .ZN(n1218) );
INV_X1 U899 ( .A(n1181), .ZN(n1207) );
NAND2_X1 U900 ( .A1(n1036), .A2(n1219), .ZN(n1181) );
NAND3_X1 U901 ( .A1(G902), .A2(n1220), .A3(n1092), .ZN(n1219) );
NOR2_X1 U902 ( .A1(n1010), .A2(G900), .ZN(n1092) );
XOR2_X1 U903 ( .A(G122), .B(n1221), .Z(G24) );
NOR2_X1 U904 ( .A1(n1005), .A2(n1190), .ZN(n1221) );
NAND4_X1 U905 ( .A1(n1205), .A2(n1195), .A3(n1021), .A4(n1222), .ZN(n1190) );
NOR2_X1 U906 ( .A1(n1194), .A2(n1223), .ZN(n1222) );
NOR2_X1 U907 ( .A1(n1213), .A2(n1212), .ZN(n1021) );
INV_X1 U908 ( .A(n1191), .ZN(n1005) );
XOR2_X1 U909 ( .A(n1184), .B(n1224), .Z(G21) );
NOR2_X1 U910 ( .A1(G119), .A2(KEYINPUT26), .ZN(n1224) );
NAND3_X1 U911 ( .A1(n1016), .A2(n1212), .A3(n1225), .ZN(n1184) );
XOR2_X1 U912 ( .A(G116), .B(n1186), .Z(G18) );
AND3_X1 U913 ( .A1(n1217), .A2(n1032), .A3(n1225), .ZN(n1186) );
AND2_X1 U914 ( .A1(n1205), .A2(n1223), .ZN(n1032) );
XOR2_X1 U915 ( .A(n1226), .B(G113), .Z(G15) );
NAND2_X1 U916 ( .A1(KEYINPUT1), .A2(n1185), .ZN(n1226) );
NAND3_X1 U917 ( .A1(n1217), .A2(n1031), .A3(n1225), .ZN(n1185) );
AND4_X1 U918 ( .A1(n1018), .A2(n1191), .A3(n1213), .A4(n1195), .ZN(n1225) );
INV_X1 U919 ( .A(n1194), .ZN(n1018) );
NAND2_X1 U920 ( .A1(n1027), .A2(n1227), .ZN(n1194) );
NOR2_X1 U921 ( .A1(n1223), .A2(n1205), .ZN(n1031) );
XNOR2_X1 U922 ( .A(n1228), .B(n1199), .ZN(G12) );
NAND3_X1 U923 ( .A1(n1016), .A2(n1200), .A3(n1019), .ZN(n1199) );
NOR2_X1 U924 ( .A1(n1213), .A2(n1217), .ZN(n1019) );
INV_X1 U925 ( .A(n1212), .ZN(n1217) );
XOR2_X1 U926 ( .A(n1047), .B(n1068), .Z(n1212) );
NAND2_X1 U927 ( .A1(G217), .A2(n1229), .ZN(n1068) );
NAND2_X1 U928 ( .A1(n1067), .A2(n1063), .ZN(n1047) );
XNOR2_X1 U929 ( .A(n1230), .B(n1231), .ZN(n1067) );
XOR2_X1 U930 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U931 ( .A(n1234), .B(n1235), .ZN(n1233) );
NAND2_X1 U932 ( .A1(KEYINPUT7), .A2(n1211), .ZN(n1235) );
NAND2_X1 U933 ( .A1(KEYINPUT41), .A2(n1157), .ZN(n1234) );
NAND2_X1 U934 ( .A1(G221), .A2(n1236), .ZN(n1232) );
XOR2_X1 U935 ( .A(n1237), .B(n1238), .Z(n1230) );
NOR2_X1 U936 ( .A1(KEYINPUT36), .A2(n1239), .ZN(n1238) );
XOR2_X1 U937 ( .A(n1240), .B(n1241), .Z(n1239) );
XNOR2_X1 U938 ( .A(KEYINPUT59), .B(n1242), .ZN(n1241) );
XNOR2_X1 U939 ( .A(G140), .B(n1243), .ZN(n1240) );
NOR2_X1 U940 ( .A1(KEYINPUT16), .A2(n1094), .ZN(n1243) );
XNOR2_X1 U941 ( .A(G119), .B(G137), .ZN(n1237) );
XNOR2_X1 U942 ( .A(n1053), .B(G472), .ZN(n1213) );
NAND2_X1 U943 ( .A1(n1244), .A2(n1063), .ZN(n1053) );
XNOR2_X1 U944 ( .A(n1139), .B(n1245), .ZN(n1244) );
XOR2_X1 U945 ( .A(n1246), .B(n1143), .Z(n1245) );
XNOR2_X1 U946 ( .A(n1108), .B(KEYINPUT57), .ZN(n1143) );
NOR2_X1 U947 ( .A1(KEYINPUT46), .A2(n1138), .ZN(n1246) );
XOR2_X1 U948 ( .A(n1247), .B(n1248), .Z(n1139) );
NAND2_X1 U949 ( .A1(G210), .A2(n1249), .ZN(n1247) );
AND3_X1 U950 ( .A1(n1026), .A2(n1195), .A3(n1191), .ZN(n1200) );
NOR2_X1 U951 ( .A1(n1033), .A2(n1034), .ZN(n1191) );
AND2_X1 U952 ( .A1(G214), .A2(n1250), .ZN(n1034) );
XOR2_X1 U953 ( .A(n1251), .B(n1163), .Z(n1033) );
AND2_X1 U954 ( .A1(G210), .A2(n1250), .ZN(n1163) );
NAND2_X1 U955 ( .A1(n1252), .A2(n1063), .ZN(n1250) );
INV_X1 U956 ( .A(G237), .ZN(n1252) );
NAND2_X1 U957 ( .A1(n1253), .A2(n1063), .ZN(n1251) );
XNOR2_X1 U958 ( .A(n1254), .B(n1255), .ZN(n1253) );
INV_X1 U959 ( .A(n1162), .ZN(n1255) );
XNOR2_X1 U960 ( .A(n1256), .B(n1106), .ZN(n1162) );
XNOR2_X1 U961 ( .A(G122), .B(n1157), .ZN(n1106) );
NAND2_X1 U962 ( .A1(n1257), .A2(KEYINPUT51), .ZN(n1256) );
XNOR2_X1 U963 ( .A(n1258), .B(n1108), .ZN(n1257) );
XNOR2_X1 U964 ( .A(G113), .B(n1259), .ZN(n1108) );
XOR2_X1 U965 ( .A(G119), .B(G116), .Z(n1259) );
NAND2_X1 U966 ( .A1(KEYINPUT8), .A2(n1107), .ZN(n1258) );
XNOR2_X1 U967 ( .A(n1260), .B(n1248), .ZN(n1107) );
NAND3_X1 U968 ( .A1(n1261), .A2(n1262), .A3(n1263), .ZN(n1260) );
OR2_X1 U969 ( .A1(G107), .A2(KEYINPUT58), .ZN(n1263) );
NAND3_X1 U970 ( .A1(KEYINPUT58), .A2(G107), .A3(n1131), .ZN(n1262) );
NAND2_X1 U971 ( .A1(G104), .A2(n1264), .ZN(n1261) );
NAND2_X1 U972 ( .A1(KEYINPUT58), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U973 ( .A(KEYINPUT38), .B(n1266), .ZN(n1265) );
NOR2_X1 U974 ( .A1(KEYINPUT15), .A2(n1159), .ZN(n1254) );
XNOR2_X1 U975 ( .A(n1094), .B(n1267), .ZN(n1159) );
XNOR2_X1 U976 ( .A(n1268), .B(n1090), .ZN(n1267) );
AND2_X1 U977 ( .A1(n1010), .A2(G224), .ZN(n1268) );
NAND2_X1 U978 ( .A1(n1036), .A2(n1269), .ZN(n1195) );
NAND3_X1 U979 ( .A1(n1102), .A2(n1220), .A3(G902), .ZN(n1269) );
NOR2_X1 U980 ( .A1(n1010), .A2(G898), .ZN(n1102) );
NAND3_X1 U981 ( .A1(n1220), .A2(n1010), .A3(G952), .ZN(n1036) );
NAND2_X1 U982 ( .A1(G237), .A2(G234), .ZN(n1220) );
NOR2_X1 U983 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
INV_X1 U984 ( .A(n1227), .ZN(n1028) );
NAND2_X1 U985 ( .A1(G221), .A2(n1229), .ZN(n1227) );
NAND2_X1 U986 ( .A1(G234), .A2(n1063), .ZN(n1229) );
XNOR2_X1 U987 ( .A(n1055), .B(n1057), .ZN(n1027) );
INV_X1 U988 ( .A(G469), .ZN(n1057) );
NAND2_X1 U989 ( .A1(n1270), .A2(n1063), .ZN(n1055) );
XOR2_X1 U990 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U991 ( .A1(n1273), .A2(n1274), .ZN(n1272) );
NOR2_X1 U992 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NOR2_X1 U993 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
INV_X1 U994 ( .A(KEYINPUT37), .ZN(n1278) );
NOR2_X1 U995 ( .A1(G110), .A2(n1279), .ZN(n1277) );
XOR2_X1 U996 ( .A(n1280), .B(KEYINPUT53), .Z(n1279) );
AND2_X1 U997 ( .A1(KEYINPUT37), .A2(n1275), .ZN(n1273) );
NOR2_X1 U998 ( .A1(n1157), .A2(n1280), .ZN(n1275) );
XNOR2_X1 U999 ( .A(G140), .B(KEYINPUT29), .ZN(n1280) );
XOR2_X1 U1000 ( .A(n1281), .B(n1153), .Z(n1271) );
AND2_X1 U1001 ( .A1(G227), .A2(n1010), .ZN(n1153) );
NAND4_X1 U1002 ( .A1(KEYINPUT45), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1281) );
NAND2_X1 U1003 ( .A1(KEYINPUT19), .A2(n1285), .ZN(n1284) );
XNOR2_X1 U1004 ( .A(n1286), .B(n1097), .ZN(n1285) );
NAND2_X1 U1005 ( .A1(n1149), .A2(n1095), .ZN(n1286) );
NAND2_X1 U1006 ( .A1(n1287), .A2(n1288), .ZN(n1283) );
INV_X1 U1007 ( .A(KEYINPUT19), .ZN(n1288) );
NAND2_X1 U1008 ( .A1(n1289), .A2(n1290), .ZN(n1287) );
NAND2_X1 U1009 ( .A1(n1138), .A2(n1149), .ZN(n1290) );
XNOR2_X1 U1010 ( .A(n1097), .B(n1095), .ZN(n1138) );
OR3_X1 U1011 ( .A1(n1097), .A2(n1090), .A3(n1149), .ZN(n1289) );
INV_X1 U1012 ( .A(n1291), .ZN(n1149) );
NAND3_X1 U1013 ( .A1(n1097), .A2(n1291), .A3(n1090), .ZN(n1282) );
INV_X1 U1014 ( .A(n1095), .ZN(n1090) );
XOR2_X1 U1015 ( .A(G146), .B(n1292), .Z(n1095) );
XNOR2_X1 U1016 ( .A(n1293), .B(n1294), .ZN(n1291) );
XNOR2_X1 U1017 ( .A(n1266), .B(G104), .ZN(n1294) );
INV_X1 U1018 ( .A(G107), .ZN(n1266) );
NAND2_X1 U1019 ( .A1(KEYINPUT30), .A2(n1248), .ZN(n1293) );
INV_X1 U1020 ( .A(G101), .ZN(n1248) );
XNOR2_X1 U1021 ( .A(G131), .B(n1295), .ZN(n1097) );
XOR2_X1 U1022 ( .A(G137), .B(G134), .Z(n1295) );
NOR2_X1 U1023 ( .A1(n1205), .A2(n1203), .ZN(n1016) );
INV_X1 U1024 ( .A(n1223), .ZN(n1203) );
XOR2_X1 U1025 ( .A(G475), .B(n1296), .Z(n1223) );
NOR2_X1 U1026 ( .A1(n1074), .A2(KEYINPUT0), .ZN(n1296) );
AND2_X1 U1027 ( .A1(n1072), .A2(n1063), .ZN(n1074) );
INV_X1 U1028 ( .A(G902), .ZN(n1063) );
XOR2_X1 U1029 ( .A(n1297), .B(n1298), .Z(n1072) );
XOR2_X1 U1030 ( .A(n1299), .B(n1300), .Z(n1298) );
XNOR2_X1 U1031 ( .A(n1131), .B(n1301), .ZN(n1300) );
NOR2_X1 U1032 ( .A1(KEYINPUT18), .A2(n1302), .ZN(n1301) );
XOR2_X1 U1033 ( .A(n1303), .B(n1304), .Z(n1302) );
XOR2_X1 U1034 ( .A(G143), .B(G131), .Z(n1304) );
NAND2_X1 U1035 ( .A1(G214), .A2(n1249), .ZN(n1303) );
NOR2_X1 U1036 ( .A1(G953), .A2(G237), .ZN(n1249) );
INV_X1 U1037 ( .A(G104), .ZN(n1131) );
NOR2_X1 U1038 ( .A1(KEYINPUT52), .A2(n1305), .ZN(n1299) );
XNOR2_X1 U1039 ( .A(n1306), .B(n1156), .ZN(n1305) );
INV_X1 U1040 ( .A(G140), .ZN(n1156) );
NAND2_X1 U1041 ( .A1(KEYINPUT17), .A2(n1094), .ZN(n1306) );
XNOR2_X1 U1042 ( .A(G125), .B(KEYINPUT48), .ZN(n1094) );
XNOR2_X1 U1043 ( .A(G113), .B(n1307), .ZN(n1297) );
XNOR2_X1 U1044 ( .A(n1242), .B(G122), .ZN(n1307) );
INV_X1 U1045 ( .A(G146), .ZN(n1242) );
XNOR2_X1 U1046 ( .A(n1060), .B(n1061), .ZN(n1205) );
INV_X1 U1047 ( .A(G478), .ZN(n1061) );
NOR2_X1 U1048 ( .A1(n1071), .A2(G902), .ZN(n1060) );
XNOR2_X1 U1049 ( .A(n1308), .B(n1309), .ZN(n1071) );
XOR2_X1 U1050 ( .A(n1310), .B(n1311), .Z(n1309) );
NAND2_X1 U1051 ( .A1(n1236), .A2(G217), .ZN(n1311) );
AND2_X1 U1052 ( .A1(G234), .A2(n1010), .ZN(n1236) );
INV_X1 U1053 ( .A(G953), .ZN(n1010) );
NAND2_X1 U1054 ( .A1(n1312), .A2(KEYINPUT13), .ZN(n1310) );
XNOR2_X1 U1055 ( .A(G134), .B(n1292), .ZN(n1312) );
XNOR2_X1 U1056 ( .A(n1211), .B(G143), .ZN(n1292) );
INV_X1 U1057 ( .A(G128), .ZN(n1211) );
XNOR2_X1 U1058 ( .A(G107), .B(n1313), .ZN(n1308) );
XOR2_X1 U1059 ( .A(G122), .B(G116), .Z(n1313) );
NAND2_X1 U1060 ( .A1(KEYINPUT5), .A2(n1157), .ZN(n1228) );
INV_X1 U1061 ( .A(G110), .ZN(n1157) );
endmodule


