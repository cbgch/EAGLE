//Key = 0001111001101101100100111010111001000110000011011111010010101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354;

XOR2_X1 U735 ( .A(G107), .B(n1029), .Z(G9) );
NOR2_X1 U736 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR3_X1 U737 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1031) );
NOR3_X1 U738 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1033) );
NOR2_X1 U739 ( .A1(n1038), .A2(n1039), .ZN(n1037) );
NOR2_X1 U740 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
INV_X1 U741 ( .A(n1042), .ZN(n1041) );
NOR2_X1 U742 ( .A1(n1043), .A2(n1044), .ZN(n1040) );
NOR4_X1 U743 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1038) );
NOR2_X1 U744 ( .A1(n1049), .A2(n1050), .ZN(n1046) );
NOR2_X1 U745 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NOR2_X1 U746 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
NOR2_X1 U747 ( .A1(n1055), .A2(n1056), .ZN(n1053) );
NOR2_X1 U748 ( .A1(n1057), .A2(n1058), .ZN(n1049) );
NOR2_X1 U749 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND3_X1 U750 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1032) );
NAND3_X1 U751 ( .A1(n1064), .A2(n1065), .A3(n1042), .ZN(n1063) );
NOR4_X1 U752 ( .A1(n1048), .A2(n1058), .A3(n1052), .A4(n1045), .ZN(n1042) );
INV_X1 U753 ( .A(KEYINPUT60), .ZN(n1048) );
NAND2_X1 U754 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NAND2_X1 U755 ( .A1(n1036), .A2(n1068), .ZN(n1067) );
XOR2_X1 U756 ( .A(KEYINPUT6), .B(n1035), .Z(n1068) );
NOR3_X1 U757 ( .A1(n1069), .A2(G953), .A3(G952), .ZN(n1030) );
INV_X1 U758 ( .A(n1061), .ZN(n1069) );
NAND2_X1 U759 ( .A1(n1070), .A2(n1071), .ZN(n1061) );
NOR4_X1 U760 ( .A1(n1036), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1071) );
XOR2_X1 U761 ( .A(n1075), .B(n1076), .Z(n1073) );
NAND2_X1 U762 ( .A1(KEYINPUT53), .A2(n1077), .ZN(n1075) );
INV_X1 U763 ( .A(n1078), .ZN(n1036) );
NOR4_X1 U764 ( .A1(n1079), .A2(n1035), .A3(n1080), .A4(n1081), .ZN(n1070) );
XNOR2_X1 U765 ( .A(G469), .B(n1082), .ZN(n1081) );
XOR2_X1 U766 ( .A(n1083), .B(n1084), .Z(n1080) );
NAND2_X1 U767 ( .A1(KEYINPUT49), .A2(n1085), .ZN(n1084) );
XOR2_X1 U768 ( .A(n1086), .B(n1087), .Z(G72) );
XOR2_X1 U769 ( .A(n1088), .B(n1089), .Z(n1087) );
NAND2_X1 U770 ( .A1(G953), .A2(n1090), .ZN(n1089) );
NAND2_X1 U771 ( .A1(G900), .A2(G227), .ZN(n1090) );
NAND2_X1 U772 ( .A1(n1091), .A2(n1092), .ZN(n1088) );
NAND2_X1 U773 ( .A1(G953), .A2(n1093), .ZN(n1092) );
XOR2_X1 U774 ( .A(n1094), .B(n1095), .Z(n1091) );
XNOR2_X1 U775 ( .A(n1096), .B(n1097), .ZN(n1095) );
XOR2_X1 U776 ( .A(n1098), .B(n1099), .Z(n1097) );
NAND2_X1 U777 ( .A1(n1100), .A2(KEYINPUT48), .ZN(n1098) );
XOR2_X1 U778 ( .A(n1101), .B(G125), .Z(n1100) );
NAND2_X1 U779 ( .A1(n1102), .A2(KEYINPUT50), .ZN(n1101) );
XNOR2_X1 U780 ( .A(G140), .B(KEYINPUT29), .ZN(n1102) );
XOR2_X1 U781 ( .A(n1103), .B(n1104), .Z(n1094) );
XOR2_X1 U782 ( .A(G146), .B(G137), .Z(n1104) );
XOR2_X1 U783 ( .A(n1105), .B(G131), .Z(n1103) );
NAND2_X1 U784 ( .A1(n1106), .A2(KEYINPUT26), .ZN(n1105) );
XNOR2_X1 U785 ( .A(G134), .B(KEYINPUT41), .ZN(n1106) );
AND2_X1 U786 ( .A1(n1107), .A2(n1062), .ZN(n1086) );
NAND2_X1 U787 ( .A1(n1108), .A2(n1109), .ZN(G69) );
NAND2_X1 U788 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U789 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
NAND2_X1 U790 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
NAND2_X1 U791 ( .A1(KEYINPUT52), .A2(n1116), .ZN(n1115) );
OR2_X1 U792 ( .A1(n1110), .A2(KEYINPUT52), .ZN(n1114) );
NOR2_X1 U793 ( .A1(n1117), .A2(KEYINPUT2), .ZN(n1110) );
INV_X1 U794 ( .A(n1116), .ZN(n1117) );
NAND2_X1 U795 ( .A1(n1118), .A2(n1119), .ZN(n1116) );
NAND2_X1 U796 ( .A1(n1120), .A2(G898), .ZN(n1119) );
XNOR2_X1 U797 ( .A(G224), .B(KEYINPUT62), .ZN(n1120) );
XOR2_X1 U798 ( .A(n1062), .B(KEYINPUT45), .Z(n1118) );
INV_X1 U799 ( .A(n1111), .ZN(n1112) );
NAND2_X1 U800 ( .A1(n1121), .A2(n1122), .ZN(n1111) );
NAND3_X1 U801 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1122) );
NAND2_X1 U802 ( .A1(KEYINPUT54), .A2(n1126), .ZN(n1124) );
NAND2_X1 U803 ( .A1(G953), .A2(n1127), .ZN(n1126) );
NAND2_X1 U804 ( .A1(G898), .A2(n1128), .ZN(n1127) );
NAND2_X1 U805 ( .A1(n1129), .A2(n1130), .ZN(n1123) );
NAND2_X1 U806 ( .A1(n1131), .A2(n1062), .ZN(n1129) );
NAND2_X1 U807 ( .A1(n1128), .A2(n1132), .ZN(n1121) );
NAND2_X1 U808 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U809 ( .A1(G898), .A2(n1135), .ZN(n1134) );
NAND2_X1 U810 ( .A1(n1125), .A2(n1136), .ZN(n1135) );
NAND2_X1 U811 ( .A1(G953), .A2(n1130), .ZN(n1136) );
NAND2_X1 U812 ( .A1(n1137), .A2(n1062), .ZN(n1133) );
NAND2_X1 U813 ( .A1(n1130), .A2(n1125), .ZN(n1137) );
INV_X1 U814 ( .A(KEYINPUT54), .ZN(n1130) );
NOR2_X1 U815 ( .A1(n1138), .A2(n1139), .ZN(G66) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR3_X1 U817 ( .A1(n1142), .A2(KEYINPUT40), .A3(n1083), .ZN(n1140) );
NOR2_X1 U818 ( .A1(n1138), .A2(n1143), .ZN(G63) );
NOR3_X1 U819 ( .A1(n1076), .A2(n1144), .A3(n1145), .ZN(n1143) );
AND3_X1 U820 ( .A1(n1146), .A2(G478), .A3(n1147), .ZN(n1145) );
NOR2_X1 U821 ( .A1(n1148), .A2(n1146), .ZN(n1144) );
NOR2_X1 U822 ( .A1(n1149), .A2(n1077), .ZN(n1148) );
INV_X1 U823 ( .A(G478), .ZN(n1077) );
NOR2_X1 U824 ( .A1(n1150), .A2(n1151), .ZN(G60) );
XOR2_X1 U825 ( .A(KEYINPUT11), .B(n1138), .Z(n1151) );
XOR2_X1 U826 ( .A(n1152), .B(n1153), .Z(n1150) );
XOR2_X1 U827 ( .A(KEYINPUT22), .B(n1154), .Z(n1153) );
AND2_X1 U828 ( .A1(G475), .A2(n1147), .ZN(n1154) );
XNOR2_X1 U829 ( .A(G104), .B(n1155), .ZN(G6) );
NAND4_X1 U830 ( .A1(n1054), .A2(n1156), .A3(n1064), .A4(n1157), .ZN(n1155) );
NOR2_X1 U831 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U832 ( .A(KEYINPUT23), .B(n1160), .Z(n1159) );
NOR2_X1 U833 ( .A1(n1138), .A2(n1161), .ZN(G57) );
XOR2_X1 U834 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U835 ( .A(n1164), .B(n1165), .Z(n1163) );
AND2_X1 U836 ( .A1(G472), .A2(n1147), .ZN(n1165) );
NOR2_X1 U837 ( .A1(n1166), .A2(n1167), .ZN(n1164) );
XOR2_X1 U838 ( .A(n1168), .B(KEYINPUT30), .Z(n1167) );
NAND2_X1 U839 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U840 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
XOR2_X1 U841 ( .A(n1171), .B(G101), .Z(n1162) );
NOR2_X1 U842 ( .A1(n1138), .A2(n1172), .ZN(G54) );
XOR2_X1 U843 ( .A(n1173), .B(n1174), .Z(n1172) );
XNOR2_X1 U844 ( .A(n1175), .B(n1176), .ZN(n1173) );
NAND3_X1 U845 ( .A1(n1147), .A2(G469), .A3(KEYINPUT44), .ZN(n1175) );
INV_X1 U846 ( .A(n1142), .ZN(n1147) );
NOR2_X1 U847 ( .A1(n1062), .A2(G952), .ZN(n1138) );
NOR2_X1 U848 ( .A1(n1177), .A2(n1178), .ZN(G51) );
XOR2_X1 U849 ( .A(n1179), .B(n1180), .Z(n1178) );
XOR2_X1 U850 ( .A(n1131), .B(n1181), .Z(n1180) );
NOR2_X1 U851 ( .A1(n1182), .A2(n1142), .ZN(n1181) );
NAND2_X1 U852 ( .A1(G902), .A2(n1034), .ZN(n1142) );
INV_X1 U853 ( .A(n1149), .ZN(n1034) );
NOR2_X1 U854 ( .A1(n1107), .A2(n1125), .ZN(n1149) );
NAND2_X1 U855 ( .A1(n1183), .A2(n1184), .ZN(n1125) );
NOR4_X1 U856 ( .A1(n1029), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1184) );
NOR3_X1 U857 ( .A1(n1047), .A2(n1188), .A3(n1189), .ZN(n1029) );
NOR4_X1 U858 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1183) );
NOR2_X1 U859 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
INV_X1 U860 ( .A(KEYINPUT16), .ZN(n1195) );
NOR2_X1 U861 ( .A1(n1066), .A2(n1196), .ZN(n1192) );
NOR2_X1 U862 ( .A1(n1197), .A2(n1158), .ZN(n1191) );
NOR2_X1 U863 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR2_X1 U864 ( .A1(n1047), .A2(n1189), .ZN(n1199) );
INV_X1 U865 ( .A(n1064), .ZN(n1047) );
NOR4_X1 U866 ( .A1(KEYINPUT16), .A2(n1200), .A3(n1201), .A4(n1156), .ZN(n1198) );
NAND4_X1 U867 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1107) );
AND4_X1 U868 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205) );
INV_X1 U869 ( .A(n1210), .ZN(n1207) );
NOR4_X1 U870 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1204) );
NOR2_X1 U871 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
AND3_X1 U872 ( .A1(n1215), .A2(n1200), .A3(n1217), .ZN(n1213) );
INV_X1 U873 ( .A(KEYINPUT58), .ZN(n1215) );
NOR2_X1 U874 ( .A1(n1218), .A2(n1219), .ZN(n1212) );
INV_X1 U875 ( .A(KEYINPUT10), .ZN(n1218) );
NOR4_X1 U876 ( .A1(KEYINPUT10), .A2(n1220), .A3(n1221), .A4(n1058), .ZN(n1211) );
INV_X1 U877 ( .A(n1222), .ZN(n1058) );
NAND3_X1 U878 ( .A1(n1223), .A2(n1066), .A3(n1060), .ZN(n1220) );
OR3_X1 U879 ( .A1(n1224), .A2(n1225), .A3(n1052), .ZN(n1203) );
OR2_X1 U880 ( .A1(n1226), .A2(n1227), .ZN(n1202) );
XOR2_X1 U881 ( .A(n1228), .B(n1229), .Z(n1179) );
NOR2_X1 U882 ( .A1(KEYINPUT61), .A2(n1230), .ZN(n1229) );
XOR2_X1 U883 ( .A(n1231), .B(n1232), .Z(n1230) );
NOR2_X1 U884 ( .A1(KEYINPUT39), .A2(n1233), .ZN(n1232) );
NOR2_X1 U885 ( .A1(n1062), .A2(n1234), .ZN(n1177) );
XOR2_X1 U886 ( .A(KEYINPUT1), .B(G952), .Z(n1234) );
XNOR2_X1 U887 ( .A(G146), .B(n1209), .ZN(G48) );
NAND3_X1 U888 ( .A1(n1235), .A2(n1236), .A3(n1060), .ZN(n1209) );
XOR2_X1 U889 ( .A(G143), .B(n1237), .Z(G45) );
NOR3_X1 U890 ( .A1(n1226), .A2(KEYINPUT55), .A3(n1227), .ZN(n1237) );
NAND3_X1 U891 ( .A1(n1235), .A2(n1079), .A3(n1043), .ZN(n1226) );
XNOR2_X1 U892 ( .A(G140), .B(n1208), .ZN(G42) );
NAND2_X1 U893 ( .A1(n1044), .A2(n1217), .ZN(n1208) );
XOR2_X1 U894 ( .A(G137), .B(n1238), .Z(G39) );
NOR4_X1 U895 ( .A1(KEYINPUT34), .A2(n1225), .A3(n1224), .A4(n1052), .ZN(n1238) );
XNOR2_X1 U896 ( .A(G134), .B(n1239), .ZN(G36) );
NAND2_X1 U897 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
NAND2_X1 U898 ( .A1(KEYINPUT27), .A2(n1210), .ZN(n1241) );
OR2_X1 U899 ( .A1(KEYINPUT0), .A2(n1210), .ZN(n1240) );
NOR3_X1 U900 ( .A1(n1224), .A2(n1188), .A3(n1200), .ZN(n1210) );
XOR2_X1 U901 ( .A(n1216), .B(n1242), .Z(G33) );
XOR2_X1 U902 ( .A(KEYINPUT63), .B(G131), .Z(n1242) );
NAND2_X1 U903 ( .A1(n1217), .A2(n1043), .ZN(n1216) );
NOR2_X1 U904 ( .A1(n1158), .A2(n1224), .ZN(n1217) );
NAND4_X1 U905 ( .A1(n1243), .A2(n1054), .A3(n1223), .A4(n1078), .ZN(n1224) );
XNOR2_X1 U906 ( .A(G128), .B(n1206), .ZN(G30) );
NAND3_X1 U907 ( .A1(n1236), .A2(n1059), .A3(n1235), .ZN(n1206) );
AND3_X1 U908 ( .A1(n1054), .A2(n1223), .A3(n1160), .ZN(n1235) );
INV_X1 U909 ( .A(n1225), .ZN(n1236) );
XOR2_X1 U910 ( .A(G101), .B(n1190), .Z(G3) );
NOR3_X1 U911 ( .A1(n1200), .A2(n1189), .A3(n1052), .ZN(n1190) );
INV_X1 U912 ( .A(n1043), .ZN(n1200) );
XOR2_X1 U913 ( .A(n1233), .B(n1219), .Z(G27) );
NAND4_X1 U914 ( .A1(n1244), .A2(n1044), .A3(n1060), .A4(n1223), .ZN(n1219) );
NAND2_X1 U915 ( .A1(n1245), .A2(n1246), .ZN(n1223) );
NAND2_X1 U916 ( .A1(n1247), .A2(n1093), .ZN(n1246) );
INV_X1 U917 ( .A(G900), .ZN(n1093) );
INV_X1 U918 ( .A(n1221), .ZN(n1044) );
XOR2_X1 U919 ( .A(G122), .B(n1187), .Z(G24) );
AND4_X1 U920 ( .A1(n1248), .A2(n1064), .A3(n1249), .A4(n1079), .ZN(n1187) );
NOR2_X1 U921 ( .A1(n1074), .A2(n1250), .ZN(n1064) );
XOR2_X1 U922 ( .A(G119), .B(n1186), .Z(G21) );
NOR3_X1 U923 ( .A1(n1052), .A2(n1225), .A3(n1251), .ZN(n1186) );
NAND2_X1 U924 ( .A1(n1250), .A2(n1074), .ZN(n1225) );
INV_X1 U925 ( .A(n1252), .ZN(n1074) );
XOR2_X1 U926 ( .A(n1253), .B(n1254), .Z(G18) );
XOR2_X1 U927 ( .A(KEYINPUT51), .B(G116), .Z(n1254) );
NAND2_X1 U928 ( .A1(n1255), .A2(n1160), .ZN(n1253) );
XOR2_X1 U929 ( .A(n1196), .B(KEYINPUT12), .Z(n1255) );
NAND4_X1 U930 ( .A1(n1222), .A2(n1043), .A3(n1059), .A4(n1156), .ZN(n1196) );
INV_X1 U931 ( .A(n1188), .ZN(n1059) );
NAND2_X1 U932 ( .A1(n1249), .A2(n1256), .ZN(n1188) );
XNOR2_X1 U933 ( .A(G113), .B(n1194), .ZN(G15) );
NAND3_X1 U934 ( .A1(n1060), .A2(n1043), .A3(n1248), .ZN(n1194) );
INV_X1 U935 ( .A(n1251), .ZN(n1248) );
NAND2_X1 U936 ( .A1(n1244), .A2(n1156), .ZN(n1251) );
INV_X1 U937 ( .A(n1201), .ZN(n1244) );
NAND2_X1 U938 ( .A1(n1222), .A2(n1160), .ZN(n1201) );
NOR2_X1 U939 ( .A1(n1055), .A2(n1072), .ZN(n1222) );
INV_X1 U940 ( .A(n1056), .ZN(n1072) );
NOR2_X1 U941 ( .A1(n1250), .A2(n1252), .ZN(n1043) );
INV_X1 U942 ( .A(n1158), .ZN(n1060) );
NAND2_X1 U943 ( .A1(n1227), .A2(n1079), .ZN(n1158) );
XOR2_X1 U944 ( .A(G110), .B(n1185), .Z(G12) );
NOR3_X1 U945 ( .A1(n1221), .A2(n1189), .A3(n1052), .ZN(n1185) );
NAND2_X1 U946 ( .A1(n1227), .A2(n1256), .ZN(n1052) );
XOR2_X1 U947 ( .A(n1079), .B(KEYINPUT28), .Z(n1256) );
XNOR2_X1 U948 ( .A(n1257), .B(G475), .ZN(n1079) );
NAND2_X1 U949 ( .A1(n1152), .A2(n1258), .ZN(n1257) );
XNOR2_X1 U950 ( .A(n1259), .B(n1260), .ZN(n1152) );
XOR2_X1 U951 ( .A(G104), .B(n1261), .Z(n1260) );
NAND2_X1 U952 ( .A1(n1262), .A2(n1263), .ZN(n1259) );
NAND2_X1 U953 ( .A1(KEYINPUT13), .A2(n1264), .ZN(n1263) );
NAND2_X1 U954 ( .A1(KEYINPUT20), .A2(n1265), .ZN(n1262) );
INV_X1 U955 ( .A(n1264), .ZN(n1265) );
XOR2_X1 U956 ( .A(n1266), .B(n1267), .Z(n1264) );
NOR2_X1 U957 ( .A1(KEYINPUT32), .A2(n1268), .ZN(n1267) );
XOR2_X1 U958 ( .A(n1269), .B(n1270), .Z(n1268) );
NOR3_X1 U959 ( .A1(n1271), .A2(G237), .A3(n1272), .ZN(n1270) );
INV_X1 U960 ( .A(G214), .ZN(n1272) );
XOR2_X1 U961 ( .A(KEYINPUT35), .B(G953), .Z(n1271) );
XOR2_X1 U962 ( .A(n1273), .B(G143), .Z(n1269) );
INV_X1 U963 ( .A(G131), .ZN(n1273) );
INV_X1 U964 ( .A(n1249), .ZN(n1227) );
XOR2_X1 U965 ( .A(n1076), .B(G478), .Z(n1249) );
NOR2_X1 U966 ( .A1(n1146), .A2(G902), .ZN(n1076) );
XNOR2_X1 U967 ( .A(n1274), .B(n1275), .ZN(n1146) );
XOR2_X1 U968 ( .A(G134), .B(n1276), .Z(n1275) );
XOR2_X1 U969 ( .A(KEYINPUT18), .B(G143), .Z(n1276) );
XOR2_X1 U970 ( .A(n1277), .B(n1278), .Z(n1274) );
XNOR2_X1 U971 ( .A(G128), .B(n1279), .ZN(n1278) );
NAND2_X1 U972 ( .A1(n1280), .A2(KEYINPUT5), .ZN(n1279) );
XNOR2_X1 U973 ( .A(G107), .B(n1281), .ZN(n1280) );
XOR2_X1 U974 ( .A(G122), .B(G116), .Z(n1281) );
NAND2_X1 U975 ( .A1(n1282), .A2(G217), .ZN(n1277) );
INV_X1 U976 ( .A(n1283), .ZN(n1282) );
NAND3_X1 U977 ( .A1(n1054), .A2(n1156), .A3(n1160), .ZN(n1189) );
INV_X1 U978 ( .A(n1066), .ZN(n1160) );
NAND2_X1 U979 ( .A1(n1035), .A2(n1078), .ZN(n1066) );
NAND2_X1 U980 ( .A1(G214), .A2(n1284), .ZN(n1078) );
INV_X1 U981 ( .A(n1243), .ZN(n1035) );
XNOR2_X1 U982 ( .A(n1285), .B(n1182), .ZN(n1243) );
NAND2_X1 U983 ( .A1(G210), .A2(n1284), .ZN(n1182) );
NAND2_X1 U984 ( .A1(n1286), .A2(n1258), .ZN(n1284) );
NAND2_X1 U985 ( .A1(n1287), .A2(n1258), .ZN(n1285) );
XOR2_X1 U986 ( .A(n1288), .B(n1128), .Z(n1287) );
INV_X1 U987 ( .A(n1131), .ZN(n1128) );
XOR2_X1 U988 ( .A(n1289), .B(n1290), .Z(n1131) );
XNOR2_X1 U989 ( .A(n1261), .B(n1291), .ZN(n1290) );
XNOR2_X1 U990 ( .A(KEYINPUT21), .B(n1292), .ZN(n1291) );
NOR2_X1 U991 ( .A1(G104), .A2(KEYINPUT36), .ZN(n1292) );
XOR2_X1 U992 ( .A(G113), .B(G122), .Z(n1261) );
XOR2_X1 U993 ( .A(n1293), .B(n1294), .Z(n1289) );
NAND2_X1 U994 ( .A1(n1295), .A2(n1296), .ZN(n1288) );
NAND2_X1 U995 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
NAND2_X1 U996 ( .A1(n1299), .A2(n1300), .ZN(n1298) );
NAND2_X1 U997 ( .A1(KEYINPUT33), .A2(n1301), .ZN(n1300) );
INV_X1 U998 ( .A(n1228), .ZN(n1301) );
INV_X1 U999 ( .A(KEYINPUT42), .ZN(n1299) );
NAND2_X1 U1000 ( .A1(n1302), .A2(n1228), .ZN(n1295) );
NAND2_X1 U1001 ( .A1(n1303), .A2(n1062), .ZN(n1228) );
XOR2_X1 U1002 ( .A(KEYINPUT14), .B(G224), .Z(n1303) );
NAND2_X1 U1003 ( .A1(KEYINPUT33), .A2(n1304), .ZN(n1302) );
OR2_X1 U1004 ( .A1(n1297), .A2(KEYINPUT42), .ZN(n1304) );
XNOR2_X1 U1005 ( .A(n1231), .B(G125), .ZN(n1297) );
XOR2_X1 U1006 ( .A(n1305), .B(n1306), .Z(n1231) );
NAND2_X1 U1007 ( .A1(n1245), .A2(n1307), .ZN(n1156) );
NAND2_X1 U1008 ( .A1(n1247), .A2(n1308), .ZN(n1307) );
INV_X1 U1009 ( .A(G898), .ZN(n1308) );
NOR3_X1 U1010 ( .A1(n1258), .A2(n1045), .A3(n1062), .ZN(n1247) );
INV_X1 U1011 ( .A(n1309), .ZN(n1045) );
NAND3_X1 U1012 ( .A1(n1309), .A2(n1062), .A3(G952), .ZN(n1245) );
NAND2_X1 U1013 ( .A1(G237), .A2(G234), .ZN(n1309) );
AND2_X1 U1014 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NAND2_X1 U1015 ( .A1(G221), .A2(n1310), .ZN(n1056) );
XOR2_X1 U1016 ( .A(n1311), .B(G469), .Z(n1055) );
NAND2_X1 U1017 ( .A1(KEYINPUT15), .A2(n1082), .ZN(n1311) );
NAND2_X1 U1018 ( .A1(n1312), .A2(n1258), .ZN(n1082) );
XNOR2_X1 U1019 ( .A(n1174), .B(n1313), .ZN(n1312) );
XNOR2_X1 U1020 ( .A(n1314), .B(KEYINPUT57), .ZN(n1313) );
NAND2_X1 U1021 ( .A1(KEYINPUT24), .A2(n1176), .ZN(n1314) );
NAND2_X1 U1022 ( .A1(G227), .A2(n1062), .ZN(n1176) );
XNOR2_X1 U1023 ( .A(n1315), .B(n1316), .ZN(n1174) );
XOR2_X1 U1024 ( .A(n1317), .B(n1096), .Z(n1316) );
XNOR2_X1 U1025 ( .A(n1318), .B(KEYINPUT43), .ZN(n1096) );
INV_X1 U1026 ( .A(n1293), .ZN(n1317) );
XOR2_X1 U1027 ( .A(n1319), .B(n1320), .Z(n1293) );
XOR2_X1 U1028 ( .A(G110), .B(G107), .Z(n1320) );
XOR2_X1 U1029 ( .A(n1321), .B(n1322), .Z(n1315) );
XOR2_X1 U1030 ( .A(G104), .B(n1323), .Z(n1322) );
NAND2_X1 U1031 ( .A1(n1252), .A2(n1250), .ZN(n1221) );
XNOR2_X1 U1032 ( .A(n1085), .B(n1083), .ZN(n1250) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1310), .ZN(n1083) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1258), .ZN(n1310) );
NOR2_X1 U1035 ( .A1(n1141), .A2(G902), .ZN(n1085) );
XNOR2_X1 U1036 ( .A(n1324), .B(n1325), .ZN(n1141) );
XOR2_X1 U1037 ( .A(n1326), .B(n1327), .Z(n1325) );
XNOR2_X1 U1038 ( .A(KEYINPUT37), .B(KEYINPUT17), .ZN(n1327) );
XOR2_X1 U1039 ( .A(n1266), .B(n1328), .Z(n1324) );
XNOR2_X1 U1040 ( .A(n1329), .B(n1330), .ZN(n1328) );
NOR3_X1 U1041 ( .A1(n1283), .A2(KEYINPUT31), .A3(n1331), .ZN(n1330) );
INV_X1 U1042 ( .A(G221), .ZN(n1331) );
NAND2_X1 U1043 ( .A1(n1332), .A2(n1062), .ZN(n1283) );
XNOR2_X1 U1044 ( .A(G234), .B(KEYINPUT4), .ZN(n1332) );
NAND3_X1 U1045 ( .A1(n1333), .A2(n1334), .A3(KEYINPUT3), .ZN(n1329) );
NAND2_X1 U1046 ( .A1(n1335), .A2(n1336), .ZN(n1334) );
INV_X1 U1047 ( .A(G110), .ZN(n1336) );
XOR2_X1 U1048 ( .A(n1337), .B(KEYINPUT7), .Z(n1335) );
NAND2_X1 U1049 ( .A1(G110), .A2(n1338), .ZN(n1333) );
XOR2_X1 U1050 ( .A(n1337), .B(KEYINPUT9), .Z(n1338) );
XOR2_X1 U1051 ( .A(n1339), .B(G128), .Z(n1337) );
INV_X1 U1052 ( .A(G119), .ZN(n1339) );
XOR2_X1 U1053 ( .A(n1233), .B(n1323), .Z(n1266) );
XOR2_X1 U1054 ( .A(G140), .B(G146), .Z(n1323) );
INV_X1 U1055 ( .A(G125), .ZN(n1233) );
XOR2_X1 U1056 ( .A(n1340), .B(n1341), .Z(n1252) );
XOR2_X1 U1057 ( .A(KEYINPUT25), .B(G472), .Z(n1341) );
NAND2_X1 U1058 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
XOR2_X1 U1059 ( .A(n1344), .B(n1345), .Z(n1343) );
XOR2_X1 U1060 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1061 ( .A(KEYINPUT19), .B(n1171), .ZN(n1347) );
NAND3_X1 U1062 ( .A1(n1286), .A2(n1062), .A3(G210), .ZN(n1171) );
INV_X1 U1063 ( .A(G953), .ZN(n1062) );
INV_X1 U1064 ( .A(G237), .ZN(n1286) );
NOR2_X1 U1065 ( .A1(KEYINPUT59), .A2(n1319), .ZN(n1346) );
INV_X1 U1066 ( .A(G101), .ZN(n1319) );
XNOR2_X1 U1067 ( .A(n1169), .B(n1170), .ZN(n1344) );
XNOR2_X1 U1068 ( .A(n1294), .B(n1348), .ZN(n1170) );
NOR2_X1 U1069 ( .A1(G113), .A2(KEYINPUT8), .ZN(n1348) );
XOR2_X1 U1070 ( .A(G116), .B(G119), .Z(n1294) );
XNOR2_X1 U1071 ( .A(n1321), .B(n1305), .ZN(n1169) );
NAND2_X1 U1072 ( .A1(n1349), .A2(KEYINPUT56), .ZN(n1305) );
XOR2_X1 U1073 ( .A(n1318), .B(G146), .Z(n1349) );
INV_X1 U1074 ( .A(G143), .ZN(n1318) );
XOR2_X1 U1075 ( .A(n1350), .B(n1306), .Z(n1321) );
INV_X1 U1076 ( .A(n1099), .ZN(n1306) );
XNOR2_X1 U1077 ( .A(G128), .B(KEYINPUT47), .ZN(n1099) );
XOR2_X1 U1078 ( .A(n1351), .B(G131), .Z(n1350) );
NAND2_X1 U1079 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND2_X1 U1080 ( .A1(G134), .A2(n1326), .ZN(n1353) );
XOR2_X1 U1081 ( .A(KEYINPUT38), .B(n1354), .Z(n1352) );
NOR2_X1 U1082 ( .A1(G134), .A2(n1326), .ZN(n1354) );
INV_X1 U1083 ( .A(G137), .ZN(n1326) );
XOR2_X1 U1084 ( .A(n1258), .B(KEYINPUT46), .Z(n1342) );
INV_X1 U1085 ( .A(G902), .ZN(n1258) );
endmodule


