//Key = 0111111001001000110011110011011000101110110010010111010100010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348;

XNOR2_X1 U739 ( .A(G107), .B(n1024), .ZN(G9) );
NOR2_X1 U740 ( .A1(n1025), .A2(n1026), .ZN(G75) );
NOR3_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
INV_X1 U742 ( .A(n1030), .ZN(n1029) );
NOR2_X1 U743 ( .A1(n1031), .A2(n1032), .ZN(n1028) );
XOR2_X1 U744 ( .A(n1033), .B(KEYINPUT43), .Z(n1031) );
NAND3_X1 U745 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1027) );
NAND3_X1 U746 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NAND2_X1 U747 ( .A1(n1040), .A2(n1033), .ZN(n1038) );
NAND4_X1 U748 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1033) );
NAND2_X1 U749 ( .A1(n1045), .A2(n1046), .ZN(n1037) );
NAND4_X1 U750 ( .A1(n1047), .A2(n1048), .A3(n1041), .A4(n1049), .ZN(n1045) );
NOR2_X1 U751 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NOR2_X1 U753 ( .A1(n1043), .A2(n1054), .ZN(n1050) );
NOR3_X1 U754 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n1054) );
NOR2_X1 U755 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
INV_X1 U756 ( .A(n1060), .ZN(n1041) );
NAND2_X1 U757 ( .A1(n1057), .A2(n1055), .ZN(n1048) );
INV_X1 U758 ( .A(n1044), .ZN(n1057) );
NAND4_X1 U759 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1042), .ZN(n1047) );
NOR2_X1 U760 ( .A1(n1064), .A2(n1058), .ZN(n1063) );
NOR3_X1 U761 ( .A1(n1065), .A2(G953), .A3(G952), .ZN(n1025) );
INV_X1 U762 ( .A(n1034), .ZN(n1065) );
NAND4_X1 U763 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1034) );
XNOR2_X1 U764 ( .A(G478), .B(n1070), .ZN(n1069) );
NOR2_X1 U765 ( .A1(KEYINPUT28), .A2(n1071), .ZN(n1070) );
INV_X1 U766 ( .A(n1072), .ZN(n1071) );
NOR2_X1 U767 ( .A1(n1073), .A2(n1074), .ZN(n1068) );
XNOR2_X1 U768 ( .A(n1075), .B(KEYINPUT17), .ZN(n1074) );
XOR2_X1 U769 ( .A(n1076), .B(KEYINPUT32), .Z(n1073) );
NAND2_X1 U770 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U771 ( .A(n1079), .B(KEYINPUT11), .Z(n1077) );
NAND2_X1 U772 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XNOR2_X1 U773 ( .A(KEYINPUT25), .B(n1082), .ZN(n1080) );
XOR2_X1 U774 ( .A(n1083), .B(KEYINPUT6), .Z(n1067) );
NAND2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XNOR2_X1 U776 ( .A(n1086), .B(n1087), .ZN(n1085) );
XNOR2_X1 U777 ( .A(G469), .B(KEYINPUT51), .ZN(n1087) );
XNOR2_X1 U778 ( .A(n1088), .B(KEYINPUT35), .ZN(n1066) );
XOR2_X1 U779 ( .A(n1089), .B(n1090), .Z(G72) );
NOR2_X1 U780 ( .A1(n1091), .A2(n1035), .ZN(n1090) );
AND2_X1 U781 ( .A1(G227), .A2(G900), .ZN(n1091) );
NAND2_X1 U782 ( .A1(n1092), .A2(n1093), .ZN(n1089) );
NAND2_X1 U783 ( .A1(n1094), .A2(n1035), .ZN(n1093) );
XOR2_X1 U784 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND3_X1 U785 ( .A1(n1096), .A2(n1097), .A3(G953), .ZN(n1092) );
INV_X1 U786 ( .A(n1098), .ZN(n1097) );
AND2_X1 U787 ( .A1(n1099), .A2(KEYINPUT23), .ZN(n1096) );
XOR2_X1 U788 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U789 ( .A(G128), .B(n1102), .Z(n1101) );
NOR2_X1 U790 ( .A1(KEYINPUT15), .A2(n1103), .ZN(n1102) );
XNOR2_X1 U791 ( .A(G131), .B(n1104), .ZN(n1103) );
XOR2_X1 U792 ( .A(n1105), .B(n1106), .Z(n1100) );
NAND2_X1 U793 ( .A1(KEYINPUT9), .A2(n1107), .ZN(n1105) );
XOR2_X1 U794 ( .A(KEYINPUT40), .B(n1108), .Z(n1107) );
NAND2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(G69) );
NAND2_X1 U796 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1113), .A2(G953), .ZN(n1112) );
XNOR2_X1 U798 ( .A(G224), .B(KEYINPUT52), .ZN(n1113) );
NAND3_X1 U799 ( .A1(G953), .A2(n1114), .A3(n1115), .ZN(n1109) );
INV_X1 U800 ( .A(n1111), .ZN(n1115) );
XNOR2_X1 U801 ( .A(n1116), .B(n1117), .ZN(n1111) );
NOR2_X1 U802 ( .A1(n1118), .A2(G953), .ZN(n1117) );
NOR2_X1 U803 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U804 ( .A1(n1121), .A2(n1122), .ZN(n1116) );
NAND2_X1 U805 ( .A1(G953), .A2(n1123), .ZN(n1122) );
XNOR2_X1 U806 ( .A(n1124), .B(n1125), .ZN(n1121) );
NAND2_X1 U807 ( .A1(G898), .A2(n1126), .ZN(n1114) );
XOR2_X1 U808 ( .A(KEYINPUT52), .B(G224), .Z(n1126) );
NOR2_X1 U809 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XNOR2_X1 U810 ( .A(n1129), .B(KEYINPUT22), .ZN(n1128) );
NOR2_X1 U811 ( .A1(n1130), .A2(n1131), .ZN(n1127) );
XOR2_X1 U812 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U813 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND2_X1 U814 ( .A1(KEYINPUT50), .A2(n1136), .ZN(n1132) );
NOR2_X1 U815 ( .A1(KEYINPUT50), .A2(n1136), .ZN(n1130) );
NOR2_X1 U816 ( .A1(n1129), .A2(n1137), .ZN(G63) );
NOR3_X1 U817 ( .A1(n1072), .A2(n1138), .A3(n1139), .ZN(n1137) );
AND3_X1 U818 ( .A1(n1140), .A2(G478), .A3(n1141), .ZN(n1139) );
NOR2_X1 U819 ( .A1(n1142), .A2(n1140), .ZN(n1138) );
NOR2_X1 U820 ( .A1(n1030), .A2(n1143), .ZN(n1142) );
NOR2_X1 U821 ( .A1(n1129), .A2(n1144), .ZN(G60) );
XNOR2_X1 U822 ( .A(n1145), .B(n1146), .ZN(n1144) );
NOR2_X1 U823 ( .A1(n1082), .A2(n1135), .ZN(n1145) );
INV_X1 U824 ( .A(n1141), .ZN(n1135) );
XOR2_X1 U825 ( .A(G104), .B(n1147), .Z(G6) );
NOR2_X1 U826 ( .A1(n1032), .A2(n1148), .ZN(n1147) );
NOR2_X1 U827 ( .A1(n1129), .A2(n1149), .ZN(G57) );
XNOR2_X1 U828 ( .A(n1150), .B(n1151), .ZN(n1149) );
XNOR2_X1 U829 ( .A(n1152), .B(n1153), .ZN(n1151) );
AND2_X1 U830 ( .A1(G472), .A2(n1141), .ZN(n1152) );
NOR2_X1 U831 ( .A1(n1129), .A2(n1154), .ZN(G54) );
XOR2_X1 U832 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U833 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U834 ( .A(n1159), .B(n1160), .Z(n1155) );
NAND2_X1 U835 ( .A1(n1141), .A2(G469), .ZN(n1160) );
NAND2_X1 U836 ( .A1(KEYINPUT53), .A2(n1161), .ZN(n1159) );
NOR2_X1 U837 ( .A1(n1129), .A2(n1162), .ZN(G51) );
XOR2_X1 U838 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U839 ( .A(n1165), .B(n1166), .Z(n1164) );
NOR2_X1 U840 ( .A1(KEYINPUT13), .A2(n1167), .ZN(n1166) );
XNOR2_X1 U841 ( .A(n1168), .B(G125), .ZN(n1167) );
NAND2_X1 U842 ( .A1(n1141), .A2(G210), .ZN(n1165) );
NOR2_X1 U843 ( .A1(n1169), .A2(n1030), .ZN(n1141) );
NOR3_X1 U844 ( .A1(n1120), .A2(n1095), .A3(n1170), .ZN(n1030) );
XNOR2_X1 U845 ( .A(n1119), .B(KEYINPUT26), .ZN(n1170) );
NAND3_X1 U846 ( .A1(n1171), .A2(n1172), .A3(n1173), .ZN(n1119) );
NAND2_X1 U847 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
INV_X1 U848 ( .A(KEYINPUT8), .ZN(n1175) );
NAND3_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1042), .ZN(n1172) );
NAND2_X1 U850 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
NAND3_X1 U851 ( .A1(n1180), .A2(n1032), .A3(KEYINPUT18), .ZN(n1178) );
NAND2_X1 U852 ( .A1(n1181), .A2(n1182), .ZN(n1176) );
NAND2_X1 U853 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND2_X1 U854 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
NAND2_X1 U855 ( .A1(KEYINPUT8), .A2(n1187), .ZN(n1186) );
OR2_X1 U856 ( .A1(n1188), .A2(KEYINPUT12), .ZN(n1185) );
NAND2_X1 U857 ( .A1(n1189), .A2(n1190), .ZN(n1171) );
NAND3_X1 U858 ( .A1(n1191), .A2(n1192), .A3(n1193), .ZN(n1190) );
NAND2_X1 U859 ( .A1(n1180), .A2(n1194), .ZN(n1193) );
INV_X1 U860 ( .A(KEYINPUT18), .ZN(n1194) );
NAND2_X1 U861 ( .A1(KEYINPUT12), .A2(n1195), .ZN(n1191) );
INV_X1 U862 ( .A(n1188), .ZN(n1195) );
NAND2_X1 U863 ( .A1(n1196), .A2(n1197), .ZN(n1095) );
AND4_X1 U864 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1197) );
AND4_X1 U865 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1196) );
NAND4_X1 U866 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1024), .ZN(n1120) );
NAND4_X1 U867 ( .A1(n1209), .A2(n1044), .A3(n1059), .A4(n1179), .ZN(n1024) );
NAND4_X1 U868 ( .A1(n1064), .A2(n1043), .A3(n1209), .A4(n1179), .ZN(n1207) );
NAND2_X1 U869 ( .A1(n1210), .A2(n1183), .ZN(n1206) );
XOR2_X1 U870 ( .A(n1148), .B(KEYINPUT37), .Z(n1210) );
NAND3_X1 U871 ( .A1(n1058), .A2(n1044), .A3(n1211), .ZN(n1148) );
NOR3_X1 U872 ( .A1(n1052), .A2(n1212), .A3(n1181), .ZN(n1211) );
NOR2_X1 U873 ( .A1(n1035), .A2(G952), .ZN(n1129) );
XOR2_X1 U874 ( .A(n1205), .B(n1213), .Z(G48) );
NOR2_X1 U875 ( .A1(G146), .A2(KEYINPUT33), .ZN(n1213) );
NAND2_X1 U876 ( .A1(n1214), .A2(n1058), .ZN(n1205) );
XNOR2_X1 U877 ( .A(G143), .B(n1204), .ZN(G45) );
NAND3_X1 U878 ( .A1(n1215), .A2(n1209), .A3(n1216), .ZN(n1204) );
AND3_X1 U879 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1216) );
XNOR2_X1 U880 ( .A(G140), .B(n1203), .ZN(G42) );
NAND3_X1 U881 ( .A1(n1058), .A2(n1064), .A3(n1220), .ZN(n1203) );
XNOR2_X1 U882 ( .A(G137), .B(n1201), .ZN(G39) );
OR2_X1 U883 ( .A1(n1192), .A2(n1221), .ZN(n1201) );
NAND2_X1 U884 ( .A1(n1222), .A2(n1223), .ZN(G36) );
NAND2_X1 U885 ( .A1(G134), .A2(n1202), .ZN(n1223) );
XOR2_X1 U886 ( .A(n1224), .B(KEYINPUT0), .Z(n1222) );
OR2_X1 U887 ( .A1(n1202), .A2(G134), .ZN(n1224) );
NAND2_X1 U888 ( .A1(n1180), .A2(n1220), .ZN(n1202) );
XNOR2_X1 U889 ( .A(G131), .B(n1200), .ZN(G33) );
NAND2_X1 U890 ( .A1(n1187), .A2(n1220), .ZN(n1200) );
INV_X1 U891 ( .A(n1221), .ZN(n1220) );
NAND3_X1 U892 ( .A1(n1225), .A2(n1219), .A3(n1084), .ZN(n1221) );
NOR3_X1 U893 ( .A1(n1040), .A2(n1212), .A3(n1226), .ZN(n1084) );
XNOR2_X1 U894 ( .A(G128), .B(n1199), .ZN(G30) );
NAND2_X1 U895 ( .A1(n1214), .A2(n1059), .ZN(n1199) );
INV_X1 U896 ( .A(n1062), .ZN(n1059) );
AND4_X1 U897 ( .A1(n1209), .A2(n1088), .A3(n1075), .A4(n1219), .ZN(n1214) );
XNOR2_X1 U898 ( .A(G101), .B(n1208), .ZN(G3) );
NAND4_X1 U899 ( .A1(n1043), .A2(n1209), .A3(n1217), .A4(n1179), .ZN(n1208) );
XNOR2_X1 U900 ( .A(G125), .B(n1198), .ZN(G27) );
NAND4_X1 U901 ( .A1(n1183), .A2(n1219), .A3(n1064), .A4(n1227), .ZN(n1198) );
AND2_X1 U902 ( .A1(n1058), .A2(n1042), .ZN(n1227) );
NAND2_X1 U903 ( .A1(n1228), .A2(n1060), .ZN(n1219) );
XOR2_X1 U904 ( .A(n1229), .B(KEYINPUT45), .Z(n1228) );
NAND4_X1 U905 ( .A1(G953), .A2(G902), .A3(n1098), .A4(n1230), .ZN(n1229) );
XOR2_X1 U906 ( .A(G900), .B(KEYINPUT1), .Z(n1098) );
XOR2_X1 U907 ( .A(n1231), .B(n1232), .Z(G24) );
XNOR2_X1 U908 ( .A(KEYINPUT56), .B(n1233), .ZN(n1232) );
NOR3_X1 U909 ( .A1(n1234), .A2(KEYINPUT7), .A3(n1188), .ZN(n1231) );
NAND3_X1 U910 ( .A1(n1215), .A2(n1218), .A3(n1044), .ZN(n1188) );
XOR2_X1 U911 ( .A(G119), .B(n1235), .Z(G21) );
NOR3_X1 U912 ( .A1(n1234), .A2(KEYINPUT54), .A3(n1192), .ZN(n1235) );
NAND3_X1 U913 ( .A1(n1088), .A2(n1075), .A3(n1043), .ZN(n1192) );
INV_X1 U914 ( .A(n1189), .ZN(n1234) );
XNOR2_X1 U915 ( .A(G116), .B(n1236), .ZN(G18) );
NAND2_X1 U916 ( .A1(n1189), .A2(n1180), .ZN(n1236) );
NOR2_X1 U917 ( .A1(n1062), .A2(n1061), .ZN(n1180) );
INV_X1 U918 ( .A(n1217), .ZN(n1061) );
NAND2_X1 U919 ( .A1(n1237), .A2(n1215), .ZN(n1062) );
NAND2_X1 U920 ( .A1(n1238), .A2(n1239), .ZN(G15) );
NAND2_X1 U921 ( .A1(n1174), .A2(n1240), .ZN(n1239) );
XOR2_X1 U922 ( .A(KEYINPUT36), .B(n1241), .Z(n1238) );
NOR2_X1 U923 ( .A1(n1174), .A2(n1240), .ZN(n1241) );
AND2_X1 U924 ( .A1(n1189), .A2(n1187), .ZN(n1174) );
AND2_X1 U925 ( .A1(n1058), .A2(n1217), .ZN(n1187) );
NAND2_X1 U926 ( .A1(n1242), .A2(n1243), .ZN(n1217) );
NAND2_X1 U927 ( .A1(n1044), .A2(n1244), .ZN(n1243) );
NOR2_X1 U928 ( .A1(n1075), .A2(n1088), .ZN(n1044) );
OR3_X1 U929 ( .A1(n1245), .A2(n1088), .A3(n1244), .ZN(n1242) );
INV_X1 U930 ( .A(KEYINPUT20), .ZN(n1244) );
NOR2_X1 U931 ( .A1(n1215), .A2(n1237), .ZN(n1058) );
INV_X1 U932 ( .A(n1218), .ZN(n1237) );
NOR3_X1 U933 ( .A1(n1032), .A2(n1181), .A3(n1055), .ZN(n1189) );
INV_X1 U934 ( .A(n1042), .ZN(n1055) );
NOR2_X1 U935 ( .A1(n1225), .A2(n1212), .ZN(n1042) );
INV_X1 U936 ( .A(n1052), .ZN(n1225) );
INV_X1 U937 ( .A(n1179), .ZN(n1181) );
XNOR2_X1 U938 ( .A(G110), .B(n1246), .ZN(G12) );
NOR2_X1 U939 ( .A1(KEYINPUT42), .A2(n1247), .ZN(n1246) );
AND4_X1 U940 ( .A1(n1248), .A2(n1209), .A3(n1043), .A4(n1064), .ZN(n1247) );
AND2_X1 U941 ( .A1(n1245), .A2(n1088), .ZN(n1064) );
XOR2_X1 U942 ( .A(n1249), .B(n1134), .Z(n1088) );
NAND2_X1 U943 ( .A1(G217), .A2(n1250), .ZN(n1134) );
OR2_X1 U944 ( .A1(n1136), .A2(G902), .ZN(n1249) );
XNOR2_X1 U945 ( .A(n1251), .B(n1252), .ZN(n1136) );
XNOR2_X1 U946 ( .A(G137), .B(n1253), .ZN(n1252) );
NAND3_X1 U947 ( .A1(G234), .A2(n1254), .A3(G221), .ZN(n1253) );
XNOR2_X1 U948 ( .A(KEYINPUT47), .B(n1035), .ZN(n1254) );
NAND2_X1 U949 ( .A1(n1255), .A2(n1256), .ZN(n1251) );
NAND4_X1 U950 ( .A1(KEYINPUT5), .A2(n1257), .A3(n1258), .A4(n1259), .ZN(n1256) );
NAND2_X1 U951 ( .A1(G110), .A2(n1260), .ZN(n1259) );
NAND2_X1 U952 ( .A1(n1261), .A2(n1161), .ZN(n1258) );
NAND3_X1 U953 ( .A1(n1262), .A2(n1263), .A3(n1264), .ZN(n1255) );
NAND2_X1 U954 ( .A1(KEYINPUT5), .A2(n1257), .ZN(n1264) );
XOR2_X1 U955 ( .A(G128), .B(G119), .Z(n1257) );
NAND2_X1 U956 ( .A1(n1260), .A2(n1161), .ZN(n1263) );
INV_X1 U957 ( .A(G110), .ZN(n1161) );
NAND2_X1 U958 ( .A1(G110), .A2(n1261), .ZN(n1262) );
XNOR2_X1 U959 ( .A(n1265), .B(n1260), .ZN(n1261) );
XNOR2_X1 U960 ( .A(KEYINPUT38), .B(KEYINPUT19), .ZN(n1265) );
INV_X1 U961 ( .A(n1075), .ZN(n1245) );
XNOR2_X1 U962 ( .A(n1266), .B(G472), .ZN(n1075) );
NAND2_X1 U963 ( .A1(n1267), .A2(n1169), .ZN(n1266) );
XOR2_X1 U964 ( .A(n1268), .B(n1269), .Z(n1267) );
XNOR2_X1 U965 ( .A(KEYINPUT2), .B(n1270), .ZN(n1269) );
INV_X1 U966 ( .A(n1150), .ZN(n1270) );
XNOR2_X1 U967 ( .A(n1271), .B(n1272), .ZN(n1150) );
XNOR2_X1 U968 ( .A(G113), .B(n1273), .ZN(n1272) );
XOR2_X1 U969 ( .A(n1274), .B(n1275), .Z(n1271) );
NAND2_X1 U970 ( .A1(n1276), .A2(n1277), .ZN(n1268) );
NAND2_X1 U971 ( .A1(KEYINPUT59), .A2(n1153), .ZN(n1277) );
INV_X1 U972 ( .A(n1278), .ZN(n1153) );
NAND2_X1 U973 ( .A1(KEYINPUT48), .A2(n1278), .ZN(n1276) );
XOR2_X1 U974 ( .A(n1279), .B(n1280), .Z(n1278) );
INV_X1 U975 ( .A(G101), .ZN(n1280) );
NAND3_X1 U976 ( .A1(n1281), .A2(n1035), .A3(n1282), .ZN(n1279) );
XNOR2_X1 U977 ( .A(G210), .B(KEYINPUT30), .ZN(n1282) );
NOR2_X1 U978 ( .A1(n1218), .A2(n1215), .ZN(n1043) );
XNOR2_X1 U979 ( .A(n1072), .B(n1283), .ZN(n1215) );
XNOR2_X1 U980 ( .A(KEYINPUT44), .B(n1143), .ZN(n1283) );
INV_X1 U981 ( .A(G478), .ZN(n1143) );
NOR2_X1 U982 ( .A1(n1140), .A2(G902), .ZN(n1072) );
XNOR2_X1 U983 ( .A(n1284), .B(n1285), .ZN(n1140) );
XOR2_X1 U984 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U985 ( .A(G107), .B(n1288), .Z(n1287) );
AND3_X1 U986 ( .A1(G217), .A2(n1035), .A3(G234), .ZN(n1288) );
XNOR2_X1 U987 ( .A(n1233), .B(G116), .ZN(n1286) );
XOR2_X1 U988 ( .A(n1289), .B(n1290), .Z(n1284) );
XNOR2_X1 U989 ( .A(KEYINPUT3), .B(n1291), .ZN(n1290) );
XNOR2_X1 U990 ( .A(G134), .B(G128), .ZN(n1289) );
NAND2_X1 U991 ( .A1(n1078), .A2(n1292), .ZN(n1218) );
NAND2_X1 U992 ( .A1(G475), .A2(n1081), .ZN(n1292) );
NAND2_X1 U993 ( .A1(n1146), .A2(n1169), .ZN(n1081) );
NAND3_X1 U994 ( .A1(n1082), .A2(n1169), .A3(n1146), .ZN(n1078) );
XOR2_X1 U995 ( .A(n1293), .B(n1294), .Z(n1146) );
XOR2_X1 U996 ( .A(G131), .B(n1295), .Z(n1294) );
NOR2_X1 U997 ( .A1(KEYINPUT62), .A2(n1296), .ZN(n1295) );
XNOR2_X1 U998 ( .A(n1291), .B(n1297), .ZN(n1296) );
AND3_X1 U999 ( .A1(G214), .A2(n1035), .A3(n1281), .ZN(n1297) );
INV_X1 U1000 ( .A(G143), .ZN(n1291) );
XNOR2_X1 U1001 ( .A(n1298), .B(n1260), .ZN(n1293) );
XOR2_X1 U1002 ( .A(n1299), .B(n1108), .Z(n1260) );
XOR2_X1 U1003 ( .A(G140), .B(G125), .Z(n1108) );
NAND2_X1 U1004 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
NAND2_X1 U1005 ( .A1(n1302), .A2(G104), .ZN(n1301) );
XOR2_X1 U1006 ( .A(n1303), .B(KEYINPUT63), .Z(n1300) );
OR2_X1 U1007 ( .A1(n1302), .A2(G104), .ZN(n1303) );
XOR2_X1 U1008 ( .A(n1304), .B(G122), .Z(n1302) );
NAND2_X1 U1009 ( .A1(KEYINPUT29), .A2(n1240), .ZN(n1304) );
INV_X1 U1010 ( .A(G475), .ZN(n1082) );
NOR3_X1 U1011 ( .A1(n1052), .A2(n1212), .A3(n1032), .ZN(n1209) );
INV_X1 U1012 ( .A(n1183), .ZN(n1032) );
NOR2_X1 U1013 ( .A1(n1040), .A2(n1039), .ZN(n1183) );
INV_X1 U1014 ( .A(n1226), .ZN(n1039) );
NAND3_X1 U1015 ( .A1(n1305), .A2(n1306), .A3(n1307), .ZN(n1226) );
NAND2_X1 U1016 ( .A1(n1308), .A2(n1309), .ZN(n1307) );
OR3_X1 U1017 ( .A1(n1309), .A2(n1308), .A3(G902), .ZN(n1306) );
AND2_X1 U1018 ( .A1(G237), .A2(G210), .ZN(n1308) );
XOR2_X1 U1019 ( .A(n1310), .B(n1311), .Z(n1309) );
XOR2_X1 U1020 ( .A(n1163), .B(n1312), .Z(n1311) );
XOR2_X1 U1021 ( .A(n1313), .B(G125), .Z(n1312) );
NAND2_X1 U1022 ( .A1(KEYINPUT41), .A2(n1168), .ZN(n1313) );
XOR2_X1 U1023 ( .A(G128), .B(n1275), .Z(n1168) );
AND2_X1 U1024 ( .A1(n1314), .A2(n1315), .ZN(n1275) );
OR2_X1 U1025 ( .A1(n1106), .A2(KEYINPUT24), .ZN(n1315) );
NAND3_X1 U1026 ( .A1(G143), .A2(n1299), .A3(KEYINPUT24), .ZN(n1314) );
XOR2_X1 U1027 ( .A(n1316), .B(n1125), .Z(n1163) );
XNOR2_X1 U1028 ( .A(n1317), .B(n1318), .ZN(n1125) );
XOR2_X1 U1029 ( .A(n1319), .B(n1274), .Z(n1318) );
XNOR2_X1 U1030 ( .A(G116), .B(G119), .ZN(n1274) );
NAND2_X1 U1031 ( .A1(KEYINPUT27), .A2(n1233), .ZN(n1319) );
INV_X1 U1032 ( .A(G122), .ZN(n1233) );
XOR2_X1 U1033 ( .A(n1320), .B(n1321), .Z(n1317) );
NOR2_X1 U1034 ( .A1(KEYINPUT10), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U1035 ( .A(KEYINPUT31), .B(n1240), .ZN(n1322) );
INV_X1 U1036 ( .A(G113), .ZN(n1240) );
XNOR2_X1 U1037 ( .A(G110), .B(KEYINPUT55), .ZN(n1320) );
XOR2_X1 U1038 ( .A(n1323), .B(n1324), .Z(n1316) );
NOR2_X1 U1039 ( .A1(KEYINPUT46), .A2(n1124), .ZN(n1324) );
NAND2_X1 U1040 ( .A1(G224), .A2(n1035), .ZN(n1323) );
XOR2_X1 U1041 ( .A(n1325), .B(n1326), .Z(n1310) );
XOR2_X1 U1042 ( .A(KEYINPUT60), .B(KEYINPUT57), .Z(n1326) );
XNOR2_X1 U1043 ( .A(KEYINPUT21), .B(KEYINPUT14), .ZN(n1325) );
NAND2_X1 U1044 ( .A1(G902), .A2(G210), .ZN(n1305) );
INV_X1 U1045 ( .A(n1046), .ZN(n1040) );
NAND2_X1 U1046 ( .A1(G214), .A2(n1327), .ZN(n1046) );
NAND2_X1 U1047 ( .A1(n1281), .A2(n1169), .ZN(n1327) );
INV_X1 U1048 ( .A(G237), .ZN(n1281) );
INV_X1 U1049 ( .A(n1053), .ZN(n1212) );
NAND2_X1 U1050 ( .A1(G221), .A2(n1250), .ZN(n1053) );
NAND2_X1 U1051 ( .A1(G234), .A2(n1169), .ZN(n1250) );
NAND3_X1 U1052 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1052) );
OR2_X1 U1053 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
NAND3_X1 U1054 ( .A1(n1332), .A2(n1331), .A3(KEYINPUT4), .ZN(n1329) );
INV_X1 U1055 ( .A(G469), .ZN(n1331) );
NOR2_X1 U1056 ( .A1(n1086), .A2(KEYINPUT39), .ZN(n1332) );
INV_X1 U1057 ( .A(n1333), .ZN(n1086) );
OR2_X1 U1058 ( .A1(n1333), .A2(KEYINPUT4), .ZN(n1328) );
NAND3_X1 U1059 ( .A1(n1334), .A2(n1335), .A3(n1169), .ZN(n1333) );
INV_X1 U1060 ( .A(G902), .ZN(n1169) );
NAND2_X1 U1061 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
XOR2_X1 U1062 ( .A(n1338), .B(n1158), .Z(n1336) );
OR3_X1 U1063 ( .A1(n1338), .A2(n1158), .A3(n1337), .ZN(n1334) );
INV_X1 U1064 ( .A(KEYINPUT61), .ZN(n1337) );
XNOR2_X1 U1065 ( .A(n1124), .B(n1339), .ZN(n1158) );
XNOR2_X1 U1066 ( .A(n1273), .B(n1106), .ZN(n1339) );
XNOR2_X1 U1067 ( .A(G143), .B(n1299), .ZN(n1106) );
INV_X1 U1068 ( .A(G146), .ZN(n1299) );
XOR2_X1 U1069 ( .A(n1340), .B(n1341), .Z(n1273) );
XOR2_X1 U1070 ( .A(G131), .B(G128), .Z(n1341) );
NAND2_X1 U1071 ( .A1(n1342), .A2(n1343), .ZN(n1340) );
NAND2_X1 U1072 ( .A1(KEYINPUT34), .A2(n1104), .ZN(n1343) );
NAND2_X1 U1073 ( .A1(KEYINPUT58), .A2(n1344), .ZN(n1342) );
INV_X1 U1074 ( .A(n1104), .ZN(n1344) );
XNOR2_X1 U1075 ( .A(G137), .B(G134), .ZN(n1104) );
XNOR2_X1 U1076 ( .A(G101), .B(n1345), .ZN(n1124) );
XOR2_X1 U1077 ( .A(G107), .B(G104), .Z(n1345) );
XNOR2_X1 U1078 ( .A(G110), .B(n1157), .ZN(n1338) );
XOR2_X1 U1079 ( .A(G140), .B(n1346), .Z(n1157) );
AND2_X1 U1080 ( .A1(n1035), .A2(G227), .ZN(n1346) );
XNOR2_X1 U1081 ( .A(n1179), .B(KEYINPUT49), .ZN(n1248) );
NAND2_X1 U1082 ( .A1(n1060), .A2(n1347), .ZN(n1179) );
NAND4_X1 U1083 ( .A1(G953), .A2(G902), .A3(n1230), .A4(n1123), .ZN(n1347) );
INV_X1 U1084 ( .A(G898), .ZN(n1123) );
NAND3_X1 U1085 ( .A1(n1230), .A2(n1035), .A3(n1348), .ZN(n1060) );
XNOR2_X1 U1086 ( .A(G952), .B(KEYINPUT16), .ZN(n1348) );
INV_X1 U1087 ( .A(G953), .ZN(n1035) );
NAND2_X1 U1088 ( .A1(G234), .A2(G237), .ZN(n1230) );
endmodule


