//Key = 0001110010000001100000111001010011000100111010100000011111010000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320;

XNOR2_X1 U726 ( .A(G107), .B(n1005), .ZN(G9) );
NOR2_X1 U727 ( .A1(n1006), .A2(n1007), .ZN(G75) );
NOR4_X1 U728 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1007) );
AND3_X1 U729 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1010) );
OR2_X1 U730 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
XOR2_X1 U731 ( .A(n1017), .B(KEYINPUT8), .Z(n1016) );
NOR2_X1 U732 ( .A1(n1018), .A2(n1019), .ZN(n1015) );
NAND3_X1 U733 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n1008) );
NAND3_X1 U734 ( .A1(n1023), .A2(n1019), .A3(n1024), .ZN(n1022) );
NAND3_X1 U735 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1023) );
NAND4_X1 U736 ( .A1(n1028), .A2(n1029), .A3(n1014), .A4(n1030), .ZN(n1027) );
NAND2_X1 U737 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
INV_X1 U738 ( .A(n1033), .ZN(n1029) );
NOR2_X1 U739 ( .A1(n1034), .A2(n1035), .ZN(n1028) );
NOR3_X1 U740 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NOR2_X1 U741 ( .A1(n1039), .A2(n1040), .ZN(n1034) );
NAND2_X1 U742 ( .A1(KEYINPUT45), .A2(n1041), .ZN(n1026) );
NAND2_X1 U743 ( .A1(n1012), .A2(n1042), .ZN(n1041) );
NAND3_X1 U744 ( .A1(n1012), .A2(n1043), .A3(n1044), .ZN(n1025) );
INV_X1 U745 ( .A(KEYINPUT45), .ZN(n1044) );
OR2_X1 U746 ( .A1(n1042), .A2(n1045), .ZN(n1043) );
NOR3_X1 U747 ( .A1(n1036), .A2(n1046), .A3(n1033), .ZN(n1012) );
NOR3_X1 U748 ( .A1(n1047), .A2(G953), .A3(G952), .ZN(n1006) );
INV_X1 U749 ( .A(n1020), .ZN(n1047) );
NAND2_X1 U750 ( .A1(n1048), .A2(n1049), .ZN(n1020) );
NOR4_X1 U751 ( .A1(n1050), .A2(n1031), .A3(n1051), .A4(n1052), .ZN(n1049) );
XOR2_X1 U752 ( .A(n1053), .B(KEYINPUT28), .Z(n1052) );
NAND3_X1 U753 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
OR2_X1 U754 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U755 ( .A1(KEYINPUT12), .A2(n1059), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1060), .A2(n1057), .ZN(n1059) );
XNOR2_X1 U757 ( .A(n1058), .B(KEYINPUT29), .ZN(n1060) );
NAND2_X1 U758 ( .A1(n1061), .A2(n1062), .ZN(n1054) );
INV_X1 U759 ( .A(KEYINPUT12), .ZN(n1062) );
NAND2_X1 U760 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
OR2_X1 U761 ( .A1(n1058), .A2(KEYINPUT29), .ZN(n1064) );
NAND3_X1 U762 ( .A1(n1058), .A2(n1057), .A3(KEYINPUT29), .ZN(n1063) );
XOR2_X1 U763 ( .A(n1065), .B(n1066), .Z(n1051) );
NOR2_X1 U764 ( .A1(G472), .A2(KEYINPUT34), .ZN(n1066) );
INV_X1 U765 ( .A(n1019), .ZN(n1050) );
NOR4_X1 U766 ( .A1(n1067), .A2(n1068), .A3(n1018), .A4(n1069), .ZN(n1048) );
XNOR2_X1 U767 ( .A(G469), .B(n1070), .ZN(n1069) );
XOR2_X1 U768 ( .A(n1071), .B(n1072), .Z(G72) );
XOR2_X1 U769 ( .A(n1073), .B(n1074), .Z(n1072) );
NOR3_X1 U770 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
NOR2_X1 U771 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
XOR2_X1 U772 ( .A(n1080), .B(KEYINPUT42), .Z(n1075) );
NAND2_X1 U773 ( .A1(n1079), .A2(n1078), .ZN(n1080) );
XOR2_X1 U774 ( .A(n1081), .B(n1082), .Z(n1079) );
NOR2_X1 U775 ( .A1(G137), .A2(KEYINPUT18), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1021), .A2(n1011), .ZN(n1073) );
NAND2_X1 U777 ( .A1(G953), .A2(n1083), .ZN(n1071) );
NAND2_X1 U778 ( .A1(G900), .A2(G227), .ZN(n1083) );
XOR2_X1 U779 ( .A(n1084), .B(n1085), .Z(G69) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1085) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
XOR2_X1 U782 ( .A(n1021), .B(KEYINPUT58), .Z(n1089) );
NOR2_X1 U783 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR2_X1 U784 ( .A1(KEYINPUT14), .A2(n1092), .ZN(n1086) );
NOR2_X1 U785 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U786 ( .A(n1021), .B(KEYINPUT3), .Z(n1094) );
NAND2_X1 U787 ( .A1(n1095), .A2(n1096), .ZN(n1084) );
NAND2_X1 U788 ( .A1(G953), .A2(n1091), .ZN(n1096) );
XOR2_X1 U789 ( .A(n1097), .B(n1098), .Z(n1095) );
NOR3_X1 U790 ( .A1(n1099), .A2(n1100), .A3(n1101), .ZN(n1098) );
AND2_X1 U791 ( .A1(n1102), .A2(KEYINPUT52), .ZN(n1101) );
NOR3_X1 U792 ( .A1(KEYINPUT52), .A2(n1103), .A3(n1102), .ZN(n1100) );
INV_X1 U793 ( .A(n1104), .ZN(n1103) );
NOR2_X1 U794 ( .A1(n1105), .A2(n1104), .ZN(n1099) );
NOR2_X1 U795 ( .A1(KEYINPUT52), .A2(n1106), .ZN(n1105) );
XOR2_X1 U796 ( .A(n1102), .B(KEYINPUT19), .Z(n1106) );
NOR2_X1 U797 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XOR2_X1 U798 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
NOR2_X1 U800 ( .A1(n1107), .A2(n1113), .ZN(G63) );
XOR2_X1 U801 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U802 ( .A(n1116), .B(KEYINPUT17), .Z(n1115) );
NAND2_X1 U803 ( .A1(n1111), .A2(G478), .ZN(n1116) );
NOR2_X1 U804 ( .A1(n1107), .A2(n1117), .ZN(G60) );
NOR3_X1 U805 ( .A1(n1058), .A2(n1118), .A3(n1119), .ZN(n1117) );
AND3_X1 U806 ( .A1(n1120), .A2(G475), .A3(n1111), .ZN(n1119) );
NOR2_X1 U807 ( .A1(n1121), .A2(n1120), .ZN(n1118) );
NOR2_X1 U808 ( .A1(n1122), .A2(n1057), .ZN(n1121) );
INV_X1 U809 ( .A(G475), .ZN(n1057) );
XOR2_X1 U810 ( .A(G104), .B(n1123), .Z(G6) );
NOR2_X1 U811 ( .A1(n1124), .A2(n1125), .ZN(G57) );
XOR2_X1 U812 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U813 ( .A1(n1128), .A2(n1129), .ZN(n1126) );
NAND4_X1 U814 ( .A1(n1130), .A2(G472), .A3(n1131), .A4(n1132), .ZN(n1129) );
XOR2_X1 U815 ( .A(n1133), .B(KEYINPUT6), .Z(n1130) );
NAND2_X1 U816 ( .A1(n1134), .A2(n1135), .ZN(n1128) );
NAND3_X1 U817 ( .A1(n1131), .A2(n1132), .A3(G472), .ZN(n1135) );
NAND2_X1 U818 ( .A1(n1136), .A2(n1137), .ZN(n1132) );
INV_X1 U819 ( .A(KEYINPUT62), .ZN(n1137) );
NAND2_X1 U820 ( .A1(KEYINPUT62), .A2(n1138), .ZN(n1131) );
NAND2_X1 U821 ( .A1(n1122), .A2(G902), .ZN(n1138) );
XNOR2_X1 U822 ( .A(KEYINPUT6), .B(n1133), .ZN(n1134) );
NOR2_X1 U823 ( .A1(G952), .A2(n1139), .ZN(n1124) );
XOR2_X1 U824 ( .A(n1021), .B(KEYINPUT49), .Z(n1139) );
NOR2_X1 U825 ( .A1(n1107), .A2(n1140), .ZN(G54) );
XOR2_X1 U826 ( .A(n1141), .B(n1142), .Z(n1140) );
XOR2_X1 U827 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U828 ( .A(n1145), .B(n1146), .Z(n1141) );
XNOR2_X1 U829 ( .A(KEYINPUT43), .B(n1147), .ZN(n1146) );
NOR2_X1 U830 ( .A1(KEYINPUT60), .A2(n1148), .ZN(n1147) );
NAND2_X1 U831 ( .A1(n1111), .A2(G469), .ZN(n1145) );
NOR2_X1 U832 ( .A1(n1107), .A2(n1149), .ZN(G51) );
XOR2_X1 U833 ( .A(n1150), .B(n1151), .Z(n1149) );
XOR2_X1 U834 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U835 ( .A(KEYINPUT7), .B(KEYINPUT5), .Z(n1153) );
NOR2_X1 U836 ( .A1(KEYINPUT30), .A2(n1154), .ZN(n1152) );
XOR2_X1 U837 ( .A(n1155), .B(KEYINPUT22), .Z(n1154) );
XOR2_X1 U838 ( .A(n1156), .B(n1157), .Z(n1150) );
XNOR2_X1 U839 ( .A(n1158), .B(n1159), .ZN(n1157) );
NOR3_X1 U840 ( .A1(n1136), .A2(KEYINPUT47), .A3(n1160), .ZN(n1159) );
INV_X1 U841 ( .A(G210), .ZN(n1160) );
INV_X1 U842 ( .A(n1111), .ZN(n1136) );
NOR2_X1 U843 ( .A1(n1161), .A2(n1122), .ZN(n1111) );
AND2_X1 U844 ( .A1(n1093), .A2(n1162), .ZN(n1122) );
XNOR2_X1 U845 ( .A(KEYINPUT51), .B(n1011), .ZN(n1162) );
NAND4_X1 U846 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1011) );
NOR4_X1 U847 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
INV_X1 U848 ( .A(n1171), .ZN(n1168) );
NOR2_X1 U849 ( .A1(n1172), .A2(n1173), .ZN(n1165) );
NOR2_X1 U850 ( .A1(n1174), .A2(n1017), .ZN(n1173) );
XOR2_X1 U851 ( .A(n1175), .B(KEYINPUT1), .Z(n1174) );
NOR3_X1 U852 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1172) );
INV_X1 U853 ( .A(n1009), .ZN(n1093) );
NAND4_X1 U854 ( .A1(n1179), .A2(n1005), .A3(n1180), .A4(n1181), .ZN(n1009) );
NOR4_X1 U855 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1123), .ZN(n1181) );
AND3_X1 U856 ( .A1(n1185), .A2(n1014), .A3(n1037), .ZN(n1123) );
NOR2_X1 U857 ( .A1(n1186), .A2(n1187), .ZN(n1180) );
NOR3_X1 U858 ( .A1(n1188), .A2(n1046), .A3(n1189), .ZN(n1187) );
INV_X1 U859 ( .A(n1039), .ZN(n1046) );
XOR2_X1 U860 ( .A(KEYINPUT44), .B(n1190), .Z(n1188) );
INV_X1 U861 ( .A(n1191), .ZN(n1186) );
NAND3_X1 U862 ( .A1(n1038), .A2(n1014), .A3(n1185), .ZN(n1005) );
NAND2_X1 U863 ( .A1(KEYINPUT57), .A2(n1192), .ZN(n1158) );
NOR2_X1 U864 ( .A1(n1021), .A2(G952), .ZN(n1107) );
XOR2_X1 U865 ( .A(n1193), .B(n1163), .Z(G48) );
NAND2_X1 U866 ( .A1(n1194), .A2(n1037), .ZN(n1163) );
XOR2_X1 U867 ( .A(G143), .B(n1195), .Z(G45) );
NOR2_X1 U868 ( .A1(n1017), .A2(n1175), .ZN(n1195) );
NAND4_X1 U869 ( .A1(n1196), .A2(n1045), .A3(n1068), .A4(n1197), .ZN(n1175) );
XNOR2_X1 U870 ( .A(G140), .B(n1164), .ZN(G42) );
NAND3_X1 U871 ( .A1(n1037), .A2(n1042), .A3(n1198), .ZN(n1164) );
XOR2_X1 U872 ( .A(n1199), .B(n1170), .Z(G39) );
AND3_X1 U873 ( .A1(n1190), .A2(n1039), .A3(n1198), .ZN(n1170) );
NOR2_X1 U874 ( .A1(KEYINPUT36), .A2(n1200), .ZN(n1199) );
XOR2_X1 U875 ( .A(KEYINPUT23), .B(G137), .Z(n1200) );
XNOR2_X1 U876 ( .A(n1169), .B(n1201), .ZN(G36) );
XOR2_X1 U877 ( .A(n1202), .B(KEYINPUT50), .Z(n1201) );
AND3_X1 U878 ( .A1(n1045), .A2(n1038), .A3(n1198), .ZN(n1169) );
NAND2_X1 U879 ( .A1(n1203), .A2(n1204), .ZN(G33) );
NAND2_X1 U880 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U881 ( .A(KEYINPUT37), .B(n1207), .Z(n1203) );
NOR2_X1 U882 ( .A1(n1205), .A2(n1206), .ZN(n1207) );
INV_X1 U883 ( .A(G131), .ZN(n1206) );
AND3_X1 U884 ( .A1(n1037), .A2(n1208), .A3(n1198), .ZN(n1205) );
INV_X1 U885 ( .A(n1176), .ZN(n1198) );
NAND3_X1 U886 ( .A1(n1024), .A2(n1019), .A3(n1196), .ZN(n1176) );
INV_X1 U887 ( .A(n1018), .ZN(n1024) );
XOR2_X1 U888 ( .A(KEYINPUT63), .B(n1045), .Z(n1208) );
XOR2_X1 U889 ( .A(n1209), .B(n1171), .Z(G30) );
NAND2_X1 U890 ( .A1(n1194), .A2(n1038), .ZN(n1171) );
AND3_X1 U891 ( .A1(n1190), .A2(n1210), .A3(n1196), .ZN(n1194) );
NOR3_X1 U892 ( .A1(n1211), .A2(n1031), .A3(n1212), .ZN(n1196) );
INV_X1 U893 ( .A(n1213), .ZN(n1031) );
NAND2_X1 U894 ( .A1(n1214), .A2(n1215), .ZN(G3) );
NAND2_X1 U895 ( .A1(G101), .A2(n1191), .ZN(n1215) );
XOR2_X1 U896 ( .A(n1216), .B(KEYINPUT35), .Z(n1214) );
OR2_X1 U897 ( .A1(n1191), .A2(G101), .ZN(n1216) );
NAND3_X1 U898 ( .A1(n1039), .A2(n1185), .A3(n1045), .ZN(n1191) );
XOR2_X1 U899 ( .A(n1167), .B(n1217), .Z(G27) );
NOR2_X1 U900 ( .A1(KEYINPUT21), .A2(n1218), .ZN(n1217) );
AND4_X1 U901 ( .A1(n1037), .A2(n1040), .A3(n1219), .A4(n1042), .ZN(n1167) );
NOR2_X1 U902 ( .A1(n1211), .A2(n1017), .ZN(n1219) );
AND2_X1 U903 ( .A1(n1033), .A2(n1220), .ZN(n1211) );
NAND3_X1 U904 ( .A1(G902), .A2(n1221), .A3(n1076), .ZN(n1220) );
AND2_X1 U905 ( .A1(G953), .A2(n1222), .ZN(n1076) );
XOR2_X1 U906 ( .A(KEYINPUT54), .B(G900), .Z(n1222) );
INV_X1 U907 ( .A(n1178), .ZN(n1037) );
XNOR2_X1 U908 ( .A(G122), .B(n1179), .ZN(G24) );
NAND4_X1 U909 ( .A1(n1223), .A2(n1014), .A3(n1068), .A4(n1197), .ZN(n1179) );
NOR2_X1 U910 ( .A1(n1224), .A2(n1225), .ZN(n1014) );
NAND2_X1 U911 ( .A1(n1226), .A2(n1227), .ZN(G21) );
NAND2_X1 U912 ( .A1(G119), .A2(n1228), .ZN(n1227) );
XOR2_X1 U913 ( .A(n1229), .B(KEYINPUT39), .Z(n1226) );
OR2_X1 U914 ( .A1(n1228), .A2(G119), .ZN(n1229) );
NAND3_X1 U915 ( .A1(n1223), .A2(n1039), .A3(n1190), .ZN(n1228) );
AND2_X1 U916 ( .A1(n1225), .A2(n1224), .ZN(n1190) );
XOR2_X1 U917 ( .A(G116), .B(n1184), .Z(G18) );
AND3_X1 U918 ( .A1(n1223), .A2(n1038), .A3(n1045), .ZN(n1184) );
INV_X1 U919 ( .A(n1177), .ZN(n1045) );
NOR2_X1 U920 ( .A1(n1197), .A2(n1230), .ZN(n1038) );
INV_X1 U921 ( .A(n1189), .ZN(n1223) );
XOR2_X1 U922 ( .A(G113), .B(n1183), .Z(G15) );
NOR3_X1 U923 ( .A1(n1177), .A2(n1189), .A3(n1178), .ZN(n1183) );
NAND2_X1 U924 ( .A1(n1230), .A2(n1197), .ZN(n1178) );
NAND2_X1 U925 ( .A1(n1040), .A2(n1231), .ZN(n1189) );
INV_X1 U926 ( .A(n1036), .ZN(n1040) );
NAND2_X1 U927 ( .A1(n1212), .A2(n1213), .ZN(n1036) );
INV_X1 U928 ( .A(n1032), .ZN(n1212) );
NAND2_X1 U929 ( .A1(n1232), .A2(n1224), .ZN(n1177) );
XOR2_X1 U930 ( .A(G110), .B(n1182), .Z(G12) );
AND3_X1 U931 ( .A1(n1042), .A2(n1185), .A3(n1039), .ZN(n1182) );
NOR2_X1 U932 ( .A1(n1068), .A2(n1197), .ZN(n1039) );
XOR2_X1 U933 ( .A(n1058), .B(G475), .Z(n1197) );
NOR2_X1 U934 ( .A1(n1120), .A2(G902), .ZN(n1058) );
XNOR2_X1 U935 ( .A(n1233), .B(n1234), .ZN(n1120) );
XNOR2_X1 U936 ( .A(n1235), .B(n1236), .ZN(n1234) );
NAND2_X1 U937 ( .A1(n1237), .A2(G214), .ZN(n1235) );
XOR2_X1 U938 ( .A(n1238), .B(n1239), .Z(n1233) );
XNOR2_X1 U939 ( .A(n1240), .B(n1241), .ZN(n1239) );
NOR2_X1 U940 ( .A1(KEYINPUT13), .A2(G131), .ZN(n1241) );
NAND2_X1 U941 ( .A1(n1242), .A2(KEYINPUT16), .ZN(n1240) );
XOR2_X1 U942 ( .A(n1078), .B(KEYINPUT11), .Z(n1242) );
XOR2_X1 U943 ( .A(G140), .B(n1218), .Z(n1078) );
NAND2_X1 U944 ( .A1(n1243), .A2(KEYINPUT33), .ZN(n1238) );
XNOR2_X1 U945 ( .A(G104), .B(n1244), .ZN(n1243) );
XOR2_X1 U946 ( .A(G122), .B(G113), .Z(n1244) );
INV_X1 U947 ( .A(n1230), .ZN(n1068) );
XOR2_X1 U948 ( .A(n1245), .B(G478), .Z(n1230) );
NAND2_X1 U949 ( .A1(n1114), .A2(n1161), .ZN(n1245) );
XOR2_X1 U950 ( .A(n1246), .B(n1247), .Z(n1114) );
NOR2_X1 U951 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
AND2_X1 U952 ( .A1(KEYINPUT61), .A2(n1250), .ZN(n1249) );
NOR2_X1 U953 ( .A1(KEYINPUT0), .A2(n1250), .ZN(n1248) );
NAND3_X1 U954 ( .A1(G234), .A2(n1021), .A3(G217), .ZN(n1250) );
NAND2_X1 U955 ( .A1(n1251), .A2(n1252), .ZN(n1246) );
NAND2_X1 U956 ( .A1(n1253), .A2(n1254), .ZN(n1252) );
XOR2_X1 U957 ( .A(G143), .B(n1255), .Z(n1253) );
NAND2_X1 U958 ( .A1(n1256), .A2(n1257), .ZN(n1251) );
XOR2_X1 U959 ( .A(KEYINPUT24), .B(n1254), .Z(n1257) );
XOR2_X1 U960 ( .A(n1258), .B(n1202), .Z(n1254) );
INV_X1 U961 ( .A(G134), .ZN(n1202) );
NAND2_X1 U962 ( .A1(n1259), .A2(KEYINPUT32), .ZN(n1258) );
XOR2_X1 U963 ( .A(n1260), .B(n1261), .Z(n1259) );
XOR2_X1 U964 ( .A(n1262), .B(G122), .Z(n1260) );
NAND2_X1 U965 ( .A1(KEYINPUT53), .A2(n1263), .ZN(n1262) );
XOR2_X1 U966 ( .A(n1264), .B(n1255), .Z(n1256) );
NOR2_X1 U967 ( .A1(G128), .A2(KEYINPUT26), .ZN(n1255) );
AND3_X1 U968 ( .A1(n1032), .A2(n1213), .A3(n1231), .ZN(n1185) );
AND2_X1 U969 ( .A1(n1210), .A2(n1265), .ZN(n1231) );
NAND2_X1 U970 ( .A1(n1033), .A2(n1266), .ZN(n1265) );
NAND4_X1 U971 ( .A1(G953), .A2(G902), .A3(n1221), .A4(n1091), .ZN(n1266) );
INV_X1 U972 ( .A(G898), .ZN(n1091) );
NAND3_X1 U973 ( .A1(n1221), .A2(n1021), .A3(G952), .ZN(n1033) );
NAND2_X1 U974 ( .A1(G234), .A2(G237), .ZN(n1221) );
INV_X1 U975 ( .A(n1017), .ZN(n1210) );
NAND2_X1 U976 ( .A1(n1019), .A2(n1018), .ZN(n1017) );
NAND3_X1 U977 ( .A1(n1267), .A2(n1268), .A3(n1269), .ZN(n1018) );
NAND2_X1 U978 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
OR3_X1 U979 ( .A1(n1271), .A2(n1270), .A3(G902), .ZN(n1268) );
AND2_X1 U980 ( .A1(G237), .A2(G210), .ZN(n1270) );
XNOR2_X1 U981 ( .A(n1272), .B(n1273), .ZN(n1271) );
XOR2_X1 U982 ( .A(n1192), .B(n1274), .Z(n1273) );
INV_X1 U983 ( .A(n1156), .ZN(n1274) );
XOR2_X1 U984 ( .A(n1218), .B(n1275), .Z(n1156) );
NOR2_X1 U985 ( .A1(G953), .A2(n1090), .ZN(n1275) );
INV_X1 U986 ( .A(G224), .ZN(n1090) );
INV_X1 U987 ( .A(G125), .ZN(n1218) );
XOR2_X1 U988 ( .A(n1276), .B(n1104), .Z(n1192) );
XOR2_X1 U989 ( .A(n1277), .B(n1278), .Z(n1104) );
NOR2_X1 U990 ( .A1(KEYINPUT38), .A2(n1279), .ZN(n1278) );
INV_X1 U991 ( .A(G113), .ZN(n1279) );
XOR2_X1 U992 ( .A(n1263), .B(G119), .Z(n1277) );
INV_X1 U993 ( .A(G116), .ZN(n1263) );
XOR2_X1 U994 ( .A(n1102), .B(n1097), .Z(n1276) );
AND2_X1 U995 ( .A1(n1280), .A2(n1281), .ZN(n1097) );
NAND2_X1 U996 ( .A1(G122), .A2(n1282), .ZN(n1281) );
XOR2_X1 U997 ( .A(KEYINPUT41), .B(n1283), .Z(n1280) );
NOR2_X1 U998 ( .A1(G122), .A2(n1282), .ZN(n1283) );
XOR2_X1 U999 ( .A(KEYINPUT40), .B(n1284), .Z(n1282) );
NAND3_X1 U1000 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1102) );
NAND2_X1 U1001 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
OR3_X1 U1002 ( .A1(n1289), .A2(n1288), .A3(n1290), .ZN(n1286) );
XNOR2_X1 U1003 ( .A(n1291), .B(n1261), .ZN(n1288) );
XNOR2_X1 U1004 ( .A(G104), .B(KEYINPUT25), .ZN(n1291) );
OR2_X1 U1005 ( .A1(KEYINPUT10), .A2(n1292), .ZN(n1289) );
NAND2_X1 U1006 ( .A1(n1292), .A2(n1290), .ZN(n1285) );
INV_X1 U1007 ( .A(KEYINPUT59), .ZN(n1290) );
XOR2_X1 U1008 ( .A(n1155), .B(KEYINPUT46), .Z(n1272) );
NAND2_X1 U1009 ( .A1(G902), .A2(G210), .ZN(n1267) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1293), .ZN(n1019) );
OR2_X1 U1011 ( .A1(G237), .A2(G902), .ZN(n1293) );
NAND2_X1 U1012 ( .A1(G221), .A2(n1294), .ZN(n1213) );
XOR2_X1 U1013 ( .A(n1070), .B(n1295), .Z(n1032) );
NOR2_X1 U1014 ( .A1(G469), .A2(KEYINPUT20), .ZN(n1295) );
NAND2_X1 U1015 ( .A1(n1296), .A2(n1161), .ZN(n1070) );
XNOR2_X1 U1016 ( .A(n1144), .B(n1297), .ZN(n1296) );
XNOR2_X1 U1017 ( .A(n1148), .B(n1143), .ZN(n1297) );
NAND2_X1 U1018 ( .A1(G227), .A2(n1021), .ZN(n1148) );
XNOR2_X1 U1019 ( .A(n1298), .B(n1299), .ZN(n1144) );
XOR2_X1 U1020 ( .A(n1300), .B(n1292), .Z(n1298) );
NAND2_X1 U1021 ( .A1(n1301), .A2(n1302), .ZN(n1300) );
NAND2_X1 U1022 ( .A1(G104), .A2(n1261), .ZN(n1302) );
XOR2_X1 U1023 ( .A(KEYINPUT56), .B(n1303), .Z(n1301) );
NOR2_X1 U1024 ( .A1(G104), .A2(n1261), .ZN(n1303) );
XOR2_X1 U1025 ( .A(G107), .B(KEYINPUT15), .Z(n1261) );
NOR2_X1 U1026 ( .A1(n1232), .A2(n1224), .ZN(n1042) );
XNOR2_X1 U1027 ( .A(n1065), .B(G472), .ZN(n1224) );
NAND2_X1 U1028 ( .A1(n1304), .A2(n1305), .ZN(n1065) );
XNOR2_X1 U1029 ( .A(n1306), .B(n1127), .ZN(n1305) );
XNOR2_X1 U1030 ( .A(n1307), .B(n1292), .ZN(n1127) );
XOR2_X1 U1031 ( .A(G101), .B(KEYINPUT9), .Z(n1292) );
NAND2_X1 U1032 ( .A1(n1237), .A2(G210), .ZN(n1307) );
NOR2_X1 U1033 ( .A1(G953), .A2(G237), .ZN(n1237) );
NAND2_X1 U1034 ( .A1(KEYINPUT27), .A2(n1133), .ZN(n1306) );
XOR2_X1 U1035 ( .A(n1308), .B(n1309), .Z(n1133) );
XOR2_X1 U1036 ( .A(G119), .B(G113), .Z(n1309) );
XNOR2_X1 U1037 ( .A(n1299), .B(n1310), .ZN(n1308) );
NOR2_X1 U1038 ( .A1(G116), .A2(KEYINPUT48), .ZN(n1310) );
XNOR2_X1 U1039 ( .A(n1311), .B(n1312), .ZN(n1299) );
INV_X1 U1040 ( .A(n1081), .ZN(n1312) );
XOR2_X1 U1041 ( .A(n1155), .B(n1313), .Z(n1081) );
XOR2_X1 U1042 ( .A(G134), .B(G131), .Z(n1313) );
XOR2_X1 U1043 ( .A(n1209), .B(n1236), .Z(n1155) );
XOR2_X1 U1044 ( .A(n1193), .B(n1264), .Z(n1236) );
INV_X1 U1045 ( .A(G143), .ZN(n1264) );
INV_X1 U1046 ( .A(G146), .ZN(n1193) );
INV_X1 U1047 ( .A(G128), .ZN(n1209) );
XNOR2_X1 U1048 ( .A(G137), .B(KEYINPUT31), .ZN(n1311) );
XOR2_X1 U1049 ( .A(KEYINPUT4), .B(G902), .Z(n1304) );
INV_X1 U1050 ( .A(n1225), .ZN(n1232) );
XNOR2_X1 U1051 ( .A(n1067), .B(KEYINPUT55), .ZN(n1225) );
XNOR2_X1 U1052 ( .A(n1314), .B(n1112), .ZN(n1067) );
AND2_X1 U1053 ( .A1(G217), .A2(n1294), .ZN(n1112) );
NAND2_X1 U1054 ( .A1(G234), .A2(n1161), .ZN(n1294) );
NAND2_X1 U1055 ( .A1(n1110), .A2(n1161), .ZN(n1314) );
INV_X1 U1056 ( .A(G902), .ZN(n1161) );
XNOR2_X1 U1057 ( .A(n1315), .B(n1316), .ZN(n1110) );
XOR2_X1 U1058 ( .A(n1317), .B(n1318), .Z(n1316) );
XOR2_X1 U1059 ( .A(G128), .B(G125), .Z(n1318) );
XOR2_X1 U1060 ( .A(G146), .B(G137), .Z(n1317) );
XNOR2_X1 U1061 ( .A(n1143), .B(n1319), .ZN(n1315) );
XOR2_X1 U1062 ( .A(G119), .B(n1320), .Z(n1319) );
AND3_X1 U1063 ( .A1(G221), .A2(n1021), .A3(G234), .ZN(n1320) );
INV_X1 U1064 ( .A(G953), .ZN(n1021) );
XOR2_X1 U1065 ( .A(G140), .B(n1284), .Z(n1143) );
XOR2_X1 U1066 ( .A(G110), .B(KEYINPUT2), .Z(n1284) );
endmodule


