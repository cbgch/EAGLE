//Key = 0110101100000110101101100001111010100111010000101000110111000111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365;

XNOR2_X1 U756 ( .A(n1032), .B(n1033), .ZN(G9) );
NOR2_X1 U757 ( .A1(n1034), .A2(n1035), .ZN(G75) );
NOR3_X1 U758 ( .A1(n1036), .A2(n1037), .A3(n1038), .ZN(n1035) );
NAND3_X1 U759 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1036) );
NAND2_X1 U760 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U761 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U762 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NAND2_X1 U763 ( .A1(n1049), .A2(n1050), .ZN(n1047) );
NAND2_X1 U764 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
OR2_X1 U765 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U766 ( .A1(n1055), .A2(n1056), .ZN(n1049) );
NAND2_X1 U767 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND2_X1 U768 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
NAND3_X1 U769 ( .A1(n1051), .A2(n1061), .A3(n1055), .ZN(n1044) );
NAND2_X1 U770 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U771 ( .A1(n1048), .A2(n1064), .ZN(n1063) );
OR2_X1 U772 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U773 ( .A1(n1046), .A2(n1067), .ZN(n1062) );
NAND2_X1 U774 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U775 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
INV_X1 U776 ( .A(n1072), .ZN(n1042) );
NOR3_X1 U777 ( .A1(n1073), .A2(G953), .A3(G952), .ZN(n1034) );
INV_X1 U778 ( .A(n1039), .ZN(n1073) );
NAND4_X1 U779 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1039) );
NOR4_X1 U780 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1077) );
XOR2_X1 U781 ( .A(n1082), .B(KEYINPUT29), .Z(n1079) );
XNOR2_X1 U782 ( .A(n1083), .B(n1084), .ZN(n1078) );
NOR2_X1 U783 ( .A1(G475), .A2(KEYINPUT51), .ZN(n1084) );
NOR3_X1 U784 ( .A1(n1085), .A2(n1070), .A3(n1086), .ZN(n1076) );
NAND2_X1 U785 ( .A1(n1087), .A2(n1088), .ZN(n1075) );
NAND2_X1 U786 ( .A1(G472), .A2(n1089), .ZN(n1074) );
XOR2_X1 U787 ( .A(n1090), .B(n1091), .Z(G72) );
NOR2_X1 U788 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR3_X1 U789 ( .A1(n1040), .A2(n1094), .A3(n1095), .ZN(n1093) );
NOR2_X1 U790 ( .A1(G953), .A2(n1096), .ZN(n1092) );
XOR2_X1 U791 ( .A(n1037), .B(n1094), .Z(n1096) );
XNOR2_X1 U792 ( .A(n1097), .B(n1098), .ZN(n1094) );
XNOR2_X1 U793 ( .A(n1099), .B(n1100), .ZN(n1098) );
NAND2_X1 U794 ( .A1(KEYINPUT22), .A2(n1101), .ZN(n1099) );
INV_X1 U795 ( .A(G134), .ZN(n1101) );
XOR2_X1 U796 ( .A(n1102), .B(n1103), .Z(n1097) );
XNOR2_X1 U797 ( .A(KEYINPUT47), .B(n1104), .ZN(n1103) );
NOR2_X1 U798 ( .A1(KEYINPUT31), .A2(n1105), .ZN(n1090) );
NOR2_X1 U799 ( .A1(n1106), .A2(n1040), .ZN(n1105) );
AND2_X1 U800 ( .A1(G227), .A2(G900), .ZN(n1106) );
XOR2_X1 U801 ( .A(n1107), .B(n1108), .Z(G69) );
XOR2_X1 U802 ( .A(n1109), .B(n1110), .Z(n1108) );
NAND2_X1 U803 ( .A1(G953), .A2(n1111), .ZN(n1110) );
NAND2_X1 U804 ( .A1(G898), .A2(G224), .ZN(n1111) );
NAND2_X1 U805 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
NAND2_X1 U806 ( .A1(G953), .A2(n1114), .ZN(n1113) );
XNOR2_X1 U807 ( .A(n1115), .B(n1116), .ZN(n1112) );
XNOR2_X1 U808 ( .A(n1117), .B(n1118), .ZN(n1116) );
NOR2_X1 U809 ( .A1(KEYINPUT40), .A2(n1119), .ZN(n1118) );
NAND2_X1 U810 ( .A1(n1120), .A2(KEYINPUT52), .ZN(n1117) );
XNOR2_X1 U811 ( .A(n1121), .B(KEYINPUT34), .ZN(n1120) );
AND2_X1 U812 ( .A1(n1038), .A2(n1040), .ZN(n1107) );
NOR2_X1 U813 ( .A1(n1122), .A2(n1123), .ZN(G66) );
XOR2_X1 U814 ( .A(n1124), .B(n1125), .Z(n1123) );
NOR2_X1 U815 ( .A1(KEYINPUT45), .A2(n1126), .ZN(n1125) );
NAND2_X1 U816 ( .A1(n1127), .A2(n1087), .ZN(n1124) );
NOR2_X1 U817 ( .A1(n1122), .A2(n1128), .ZN(G63) );
XOR2_X1 U818 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U819 ( .A1(n1127), .A2(G478), .ZN(n1129) );
NOR2_X1 U820 ( .A1(n1122), .A2(n1131), .ZN(G60) );
NOR3_X1 U821 ( .A1(n1083), .A2(n1132), .A3(n1133), .ZN(n1131) );
NOR3_X1 U822 ( .A1(n1134), .A2(n1135), .A3(n1136), .ZN(n1133) );
NOR2_X1 U823 ( .A1(n1137), .A2(n1138), .ZN(n1132) );
NOR2_X1 U824 ( .A1(n1139), .A2(n1135), .ZN(n1137) );
NOR2_X1 U825 ( .A1(n1037), .A2(n1038), .ZN(n1139) );
XNOR2_X1 U826 ( .A(n1140), .B(n1141), .ZN(G6) );
NOR2_X1 U827 ( .A1(n1122), .A2(n1142), .ZN(G57) );
XOR2_X1 U828 ( .A(n1143), .B(n1144), .Z(n1142) );
XOR2_X1 U829 ( .A(n1145), .B(n1146), .Z(n1144) );
XOR2_X1 U830 ( .A(n1147), .B(n1148), .Z(n1143) );
XNOR2_X1 U831 ( .A(n1149), .B(KEYINPUT46), .ZN(n1148) );
NAND2_X1 U832 ( .A1(KEYINPUT48), .A2(n1150), .ZN(n1149) );
AND2_X1 U833 ( .A1(G472), .A2(n1127), .ZN(n1147) );
NOR2_X1 U834 ( .A1(n1122), .A2(n1151), .ZN(G54) );
XOR2_X1 U835 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U836 ( .A(n1154), .B(n1155), .Z(n1153) );
AND2_X1 U837 ( .A1(G469), .A2(n1127), .ZN(n1154) );
XOR2_X1 U838 ( .A(n1156), .B(n1157), .Z(n1152) );
NOR2_X1 U839 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U840 ( .A(n1160), .B(KEYINPUT27), .Z(n1159) );
NAND2_X1 U841 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NOR2_X1 U842 ( .A1(n1162), .A2(n1161), .ZN(n1158) );
XNOR2_X1 U843 ( .A(KEYINPUT12), .B(n1163), .ZN(n1161) );
XNOR2_X1 U844 ( .A(G128), .B(KEYINPUT62), .ZN(n1156) );
NOR2_X1 U845 ( .A1(n1122), .A2(n1164), .ZN(G51) );
XOR2_X1 U846 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U847 ( .A(n1167), .B(KEYINPUT20), .Z(n1166) );
NAND2_X1 U848 ( .A1(n1127), .A2(n1168), .ZN(n1167) );
INV_X1 U849 ( .A(n1136), .ZN(n1127) );
NAND2_X1 U850 ( .A1(G902), .A2(n1169), .ZN(n1136) );
OR2_X1 U851 ( .A1(n1038), .A2(n1037), .ZN(n1169) );
NAND4_X1 U852 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1037) );
AND4_X1 U853 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173) );
NAND2_X1 U854 ( .A1(n1178), .A2(n1179), .ZN(n1172) );
XNOR2_X1 U855 ( .A(KEYINPUT10), .B(n1180), .ZN(n1179) );
NAND2_X1 U856 ( .A1(n1048), .A2(n1181), .ZN(n1170) );
NAND2_X1 U857 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U858 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NAND2_X1 U859 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NAND2_X1 U860 ( .A1(KEYINPUT7), .A2(n1066), .ZN(n1187) );
OR2_X1 U861 ( .A1(n1188), .A2(KEYINPUT7), .ZN(n1182) );
NAND2_X1 U862 ( .A1(n1189), .A2(n1190), .ZN(n1038) );
NOR4_X1 U863 ( .A1(n1191), .A2(n1192), .A3(n1033), .A4(n1193), .ZN(n1190) );
AND3_X1 U864 ( .A1(n1194), .A2(n1054), .A3(n1046), .ZN(n1033) );
NOR4_X1 U865 ( .A1(n1141), .A2(n1195), .A3(n1196), .A4(n1197), .ZN(n1189) );
NOR2_X1 U866 ( .A1(n1198), .A2(n1199), .ZN(n1197) );
NOR2_X1 U867 ( .A1(n1200), .A2(n1201), .ZN(n1198) );
INV_X1 U868 ( .A(n1202), .ZN(n1201) );
NOR2_X1 U869 ( .A1(KEYINPUT58), .A2(n1203), .ZN(n1200) );
NOR3_X1 U870 ( .A1(n1186), .A2(n1204), .A3(n1205), .ZN(n1196) );
XNOR2_X1 U871 ( .A(n1055), .B(KEYINPUT5), .ZN(n1204) );
NOR3_X1 U872 ( .A1(n1206), .A2(n1203), .A3(n1207), .ZN(n1195) );
INV_X1 U873 ( .A(KEYINPUT58), .ZN(n1207) );
NAND3_X1 U874 ( .A1(n1208), .A2(n1068), .A3(n1051), .ZN(n1206) );
INV_X1 U875 ( .A(n1080), .ZN(n1051) );
AND3_X1 U876 ( .A1(n1046), .A2(n1194), .A3(n1053), .ZN(n1141) );
NOR2_X1 U877 ( .A1(n1040), .A2(G952), .ZN(n1122) );
XNOR2_X1 U878 ( .A(G146), .B(n1171), .ZN(G48) );
NAND3_X1 U879 ( .A1(n1209), .A2(n1178), .A3(n1184), .ZN(n1171) );
XNOR2_X1 U880 ( .A(G143), .B(n1177), .ZN(G45) );
NAND4_X1 U881 ( .A1(n1210), .A2(n1178), .A3(n1066), .A4(n1211), .ZN(n1177) );
AND3_X1 U882 ( .A1(n1212), .A2(n1213), .A3(n1081), .ZN(n1211) );
XNOR2_X1 U883 ( .A(G140), .B(n1214), .ZN(G42) );
NAND3_X1 U884 ( .A1(n1184), .A2(n1215), .A3(n1216), .ZN(n1214) );
XNOR2_X1 U885 ( .A(n1048), .B(KEYINPUT37), .ZN(n1216) );
XNOR2_X1 U886 ( .A(KEYINPUT0), .B(n1186), .ZN(n1215) );
XNOR2_X1 U887 ( .A(G137), .B(n1176), .ZN(G39) );
NAND3_X1 U888 ( .A1(n1055), .A2(n1209), .A3(n1217), .ZN(n1176) );
INV_X1 U889 ( .A(n1218), .ZN(n1217) );
XNOR2_X1 U890 ( .A(G134), .B(n1175), .ZN(G36) );
OR2_X1 U891 ( .A1(n1218), .A2(n1203), .ZN(n1175) );
NAND3_X1 U892 ( .A1(n1212), .A2(n1213), .A3(n1048), .ZN(n1218) );
XNOR2_X1 U893 ( .A(G131), .B(n1219), .ZN(G33) );
NAND2_X1 U894 ( .A1(n1188), .A2(n1048), .ZN(n1219) );
NOR2_X1 U895 ( .A1(n1220), .A2(n1221), .ZN(n1048) );
AND2_X1 U896 ( .A1(n1184), .A2(n1066), .ZN(n1188) );
AND3_X1 U897 ( .A1(n1212), .A2(n1213), .A3(n1053), .ZN(n1184) );
XNOR2_X1 U898 ( .A(n1222), .B(n1223), .ZN(G30) );
NOR2_X1 U899 ( .A1(n1068), .A2(n1180), .ZN(n1223) );
NAND4_X1 U900 ( .A1(n1209), .A2(n1054), .A3(n1224), .A4(n1213), .ZN(n1180) );
XNOR2_X1 U901 ( .A(n1225), .B(n1193), .ZN(G3) );
AND3_X1 U902 ( .A1(n1066), .A2(n1194), .A3(n1055), .ZN(n1193) );
INV_X1 U903 ( .A(n1205), .ZN(n1194) );
XNOR2_X1 U904 ( .A(G125), .B(n1174), .ZN(G27) );
NAND4_X1 U905 ( .A1(n1065), .A2(n1053), .A3(n1226), .A4(n1213), .ZN(n1174) );
NAND2_X1 U906 ( .A1(n1072), .A2(n1227), .ZN(n1213) );
NAND4_X1 U907 ( .A1(G953), .A2(G902), .A3(n1228), .A4(n1095), .ZN(n1227) );
INV_X1 U908 ( .A(G900), .ZN(n1095) );
INV_X1 U909 ( .A(n1186), .ZN(n1065) );
XOR2_X1 U910 ( .A(n1229), .B(n1230), .Z(G24) );
NOR2_X1 U911 ( .A1(KEYINPUT50), .A2(n1231), .ZN(n1230) );
NOR3_X1 U912 ( .A1(n1202), .A2(n1232), .A3(n1233), .ZN(n1229) );
NOR2_X1 U913 ( .A1(KEYINPUT30), .A2(n1234), .ZN(n1233) );
NOR2_X1 U914 ( .A1(n1235), .A2(n1208), .ZN(n1234) );
INV_X1 U915 ( .A(n1226), .ZN(n1235) );
AND2_X1 U916 ( .A1(n1199), .A2(KEYINPUT30), .ZN(n1232) );
NAND3_X1 U917 ( .A1(n1046), .A2(n1081), .A3(n1210), .ZN(n1202) );
AND2_X1 U918 ( .A1(n1236), .A2(n1237), .ZN(n1046) );
XOR2_X1 U919 ( .A(G119), .B(n1192), .Z(G21) );
AND3_X1 U920 ( .A1(n1209), .A2(n1238), .A3(n1055), .ZN(n1192) );
NOR2_X1 U921 ( .A1(n1236), .A2(n1237), .ZN(n1209) );
XNOR2_X1 U922 ( .A(n1239), .B(n1240), .ZN(G18) );
NOR2_X1 U923 ( .A1(n1199), .A2(n1203), .ZN(n1240) );
NAND2_X1 U924 ( .A1(n1066), .A2(n1054), .ZN(n1203) );
NOR2_X1 U925 ( .A1(n1241), .A2(n1210), .ZN(n1054) );
INV_X1 U926 ( .A(n1081), .ZN(n1241) );
XOR2_X1 U927 ( .A(G113), .B(n1191), .Z(G15) );
AND3_X1 U928 ( .A1(n1053), .A2(n1238), .A3(n1066), .ZN(n1191) );
NOR2_X1 U929 ( .A1(n1242), .A2(n1236), .ZN(n1066) );
INV_X1 U930 ( .A(n1199), .ZN(n1238) );
NAND2_X1 U931 ( .A1(n1226), .A2(n1208), .ZN(n1199) );
NOR2_X1 U932 ( .A1(n1080), .A2(n1068), .ZN(n1226) );
INV_X1 U933 ( .A(n1178), .ZN(n1068) );
NAND2_X1 U934 ( .A1(n1060), .A2(n1243), .ZN(n1080) );
NOR2_X1 U935 ( .A1(n1244), .A2(n1081), .ZN(n1053) );
XNOR2_X1 U936 ( .A(n1162), .B(n1245), .ZN(G12) );
NOR4_X1 U937 ( .A1(KEYINPUT3), .A2(n1205), .A3(n1246), .A4(n1186), .ZN(n1245) );
NAND2_X1 U938 ( .A1(n1236), .A2(n1242), .ZN(n1186) );
INV_X1 U939 ( .A(n1237), .ZN(n1242) );
NOR2_X1 U940 ( .A1(n1247), .A2(n1085), .ZN(n1237) );
NOR3_X1 U941 ( .A1(n1087), .A2(G902), .A3(n1126), .ZN(n1085) );
INV_X1 U942 ( .A(n1248), .ZN(n1126) );
AND2_X1 U943 ( .A1(n1249), .A2(n1088), .ZN(n1247) );
NAND2_X1 U944 ( .A1(n1248), .A2(n1250), .ZN(n1088) );
XNOR2_X1 U945 ( .A(n1251), .B(n1252), .ZN(n1248) );
XNOR2_X1 U946 ( .A(n1253), .B(n1254), .ZN(n1252) );
XNOR2_X1 U947 ( .A(n1255), .B(n1256), .ZN(n1254) );
NOR2_X1 U948 ( .A1(G110), .A2(KEYINPUT59), .ZN(n1256) );
NAND2_X1 U949 ( .A1(KEYINPUT14), .A2(G146), .ZN(n1255) );
INV_X1 U950 ( .A(n1100), .ZN(n1253) );
XNOR2_X1 U951 ( .A(n1257), .B(n1258), .ZN(n1100) );
XNOR2_X1 U952 ( .A(G125), .B(G137), .ZN(n1257) );
XOR2_X1 U953 ( .A(n1259), .B(n1260), .Z(n1251) );
XOR2_X1 U954 ( .A(KEYINPUT19), .B(G119), .Z(n1260) );
NAND2_X1 U955 ( .A1(G221), .A2(n1261), .ZN(n1259) );
XOR2_X1 U956 ( .A(n1262), .B(n1087), .Z(n1249) );
AND2_X1 U957 ( .A1(G217), .A2(n1263), .ZN(n1087) );
XNOR2_X1 U958 ( .A(KEYINPUT28), .B(KEYINPUT11), .ZN(n1262) );
NOR2_X1 U959 ( .A1(n1264), .A2(n1086), .ZN(n1236) );
NOR2_X1 U960 ( .A1(n1089), .A2(G472), .ZN(n1086) );
AND2_X1 U961 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
XOR2_X1 U962 ( .A(KEYINPUT25), .B(G472), .Z(n1266) );
XOR2_X1 U963 ( .A(n1089), .B(KEYINPUT24), .Z(n1265) );
NAND2_X1 U964 ( .A1(n1267), .A2(n1250), .ZN(n1089) );
XOR2_X1 U965 ( .A(n1268), .B(n1145), .Z(n1267) );
XNOR2_X1 U966 ( .A(n1269), .B(n1270), .ZN(n1145) );
XNOR2_X1 U967 ( .A(G101), .B(n1271), .ZN(n1270) );
NAND2_X1 U968 ( .A1(G210), .A2(n1272), .ZN(n1271) );
XNOR2_X1 U969 ( .A(n1150), .B(n1273), .ZN(n1268) );
NOR2_X1 U970 ( .A1(KEYINPUT23), .A2(n1146), .ZN(n1273) );
XOR2_X1 U971 ( .A(G113), .B(n1274), .Z(n1146) );
XNOR2_X1 U972 ( .A(n1275), .B(KEYINPUT55), .ZN(n1150) );
INV_X1 U973 ( .A(n1055), .ZN(n1246) );
NOR2_X1 U974 ( .A1(n1081), .A2(n1210), .ZN(n1055) );
INV_X1 U975 ( .A(n1244), .ZN(n1210) );
XOR2_X1 U976 ( .A(n1276), .B(n1135), .Z(n1244) );
INV_X1 U977 ( .A(G475), .ZN(n1135) );
NAND2_X1 U978 ( .A1(KEYINPUT32), .A2(n1277), .ZN(n1276) );
INV_X1 U979 ( .A(n1083), .ZN(n1277) );
NOR2_X1 U980 ( .A1(n1138), .A2(G902), .ZN(n1083) );
INV_X1 U981 ( .A(n1134), .ZN(n1138) );
XNOR2_X1 U982 ( .A(n1278), .B(n1279), .ZN(n1134) );
NOR2_X1 U983 ( .A1(KEYINPUT8), .A2(n1280), .ZN(n1279) );
XOR2_X1 U984 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR3_X1 U985 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1282) );
NOR2_X1 U986 ( .A1(n1286), .A2(n1104), .ZN(n1285) );
NOR3_X1 U987 ( .A1(G131), .A2(KEYINPUT26), .A3(n1287), .ZN(n1284) );
INV_X1 U988 ( .A(n1286), .ZN(n1287) );
NOR2_X1 U989 ( .A1(KEYINPUT35), .A2(n1288), .ZN(n1286) );
AND2_X1 U990 ( .A1(n1288), .A2(KEYINPUT26), .ZN(n1283) );
XOR2_X1 U991 ( .A(n1289), .B(n1290), .Z(n1288) );
NAND2_X1 U992 ( .A1(G214), .A2(n1272), .ZN(n1289) );
NOR2_X1 U993 ( .A1(G953), .A2(G237), .ZN(n1272) );
NOR2_X1 U994 ( .A1(KEYINPUT44), .A2(n1291), .ZN(n1281) );
XOR2_X1 U995 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U996 ( .A(n1163), .B(G125), .ZN(n1293) );
INV_X1 U997 ( .A(G140), .ZN(n1163) );
XOR2_X1 U998 ( .A(KEYINPUT41), .B(G146), .Z(n1292) );
XNOR2_X1 U999 ( .A(n1294), .B(n1140), .ZN(n1278) );
NAND3_X1 U1000 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
OR2_X1 U1001 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND3_X1 U1002 ( .A1(n1299), .A2(n1298), .A3(G122), .ZN(n1296) );
NAND2_X1 U1003 ( .A1(n1300), .A2(n1231), .ZN(n1295) );
NAND2_X1 U1004 ( .A1(n1301), .A2(n1298), .ZN(n1300) );
INV_X1 U1005 ( .A(KEYINPUT54), .ZN(n1298) );
XNOR2_X1 U1006 ( .A(n1299), .B(KEYINPUT61), .ZN(n1301) );
XOR2_X1 U1007 ( .A(G113), .B(KEYINPUT21), .Z(n1299) );
XNOR2_X1 U1008 ( .A(n1302), .B(G478), .ZN(n1081) );
NAND2_X1 U1009 ( .A1(n1130), .A2(n1250), .ZN(n1302) );
XNOR2_X1 U1010 ( .A(n1303), .B(n1304), .ZN(n1130) );
XOR2_X1 U1011 ( .A(n1305), .B(n1306), .Z(n1304) );
NAND2_X1 U1012 ( .A1(n1261), .A2(G217), .ZN(n1306) );
AND2_X1 U1013 ( .A1(G234), .A2(n1040), .ZN(n1261) );
NAND2_X1 U1014 ( .A1(KEYINPUT57), .A2(n1307), .ZN(n1305) );
XNOR2_X1 U1015 ( .A(n1222), .B(n1308), .ZN(n1307) );
XNOR2_X1 U1016 ( .A(n1290), .B(G134), .ZN(n1308) );
INV_X1 U1017 ( .A(G143), .ZN(n1290) );
NAND2_X1 U1018 ( .A1(n1309), .A2(n1310), .ZN(n1303) );
NAND2_X1 U1019 ( .A1(n1311), .A2(n1239), .ZN(n1310) );
NAND2_X1 U1020 ( .A1(n1312), .A2(n1313), .ZN(n1311) );
NAND2_X1 U1021 ( .A1(n1314), .A2(n1032), .ZN(n1313) );
NAND2_X1 U1022 ( .A1(n1315), .A2(n1316), .ZN(n1312) );
NAND2_X1 U1023 ( .A1(G116), .A2(n1317), .ZN(n1309) );
NAND2_X1 U1024 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND2_X1 U1025 ( .A1(n1316), .A2(n1032), .ZN(n1319) );
NAND2_X1 U1026 ( .A1(n1315), .A2(n1314), .ZN(n1318) );
INV_X1 U1027 ( .A(n1316), .ZN(n1314) );
NOR2_X1 U1028 ( .A1(KEYINPUT17), .A2(n1231), .ZN(n1316) );
XNOR2_X1 U1029 ( .A(n1320), .B(G107), .ZN(n1315) );
XNOR2_X1 U1030 ( .A(KEYINPUT53), .B(KEYINPUT2), .ZN(n1320) );
NAND3_X1 U1031 ( .A1(n1224), .A2(n1208), .A3(n1178), .ZN(n1205) );
NOR2_X1 U1032 ( .A1(n1071), .A2(n1220), .ZN(n1178) );
XOR2_X1 U1033 ( .A(n1070), .B(KEYINPUT49), .Z(n1220) );
AND2_X1 U1034 ( .A1(G214), .A2(n1321), .ZN(n1070) );
XOR2_X1 U1035 ( .A(KEYINPUT63), .B(n1322), .Z(n1321) );
INV_X1 U1036 ( .A(n1221), .ZN(n1071) );
XOR2_X1 U1037 ( .A(n1082), .B(KEYINPUT16), .Z(n1221) );
XOR2_X1 U1038 ( .A(n1323), .B(n1168), .Z(n1082) );
NOR2_X1 U1039 ( .A1(n1324), .A2(n1322), .ZN(n1168) );
NOR2_X1 U1040 ( .A1(G902), .A2(G237), .ZN(n1322) );
INV_X1 U1041 ( .A(G210), .ZN(n1324) );
NAND2_X1 U1042 ( .A1(n1325), .A2(n1250), .ZN(n1323) );
XOR2_X1 U1043 ( .A(n1165), .B(KEYINPUT60), .Z(n1325) );
XOR2_X1 U1044 ( .A(n1326), .B(n1327), .Z(n1165) );
XOR2_X1 U1045 ( .A(n1275), .B(n1328), .Z(n1327) );
XNOR2_X1 U1046 ( .A(G125), .B(n1329), .ZN(n1328) );
AND2_X1 U1047 ( .A1(n1040), .A2(G224), .ZN(n1329) );
NAND3_X1 U1048 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1275) );
OR2_X1 U1049 ( .A1(n1333), .A2(KEYINPUT13), .ZN(n1332) );
NAND3_X1 U1050 ( .A1(KEYINPUT13), .A2(n1333), .A3(n1222), .ZN(n1331) );
NAND2_X1 U1051 ( .A1(G128), .A2(n1334), .ZN(n1330) );
NAND2_X1 U1052 ( .A1(KEYINPUT13), .A2(n1335), .ZN(n1334) );
XOR2_X1 U1053 ( .A(KEYINPUT9), .B(n1333), .Z(n1335) );
XOR2_X1 U1054 ( .A(G146), .B(n1336), .Z(n1333) );
XNOR2_X1 U1055 ( .A(n1337), .B(n1338), .ZN(n1326) );
INV_X1 U1056 ( .A(n1121), .ZN(n1338) );
XNOR2_X1 U1057 ( .A(n1339), .B(n1340), .ZN(n1121) );
XNOR2_X1 U1058 ( .A(KEYINPUT43), .B(n1032), .ZN(n1340) );
XNOR2_X1 U1059 ( .A(G101), .B(G104), .ZN(n1339) );
XOR2_X1 U1060 ( .A(n1341), .B(n1119), .Z(n1337) );
XNOR2_X1 U1061 ( .A(n1231), .B(G110), .ZN(n1119) );
INV_X1 U1062 ( .A(G122), .ZN(n1231) );
NAND2_X1 U1063 ( .A1(KEYINPUT38), .A2(n1115), .ZN(n1341) );
XOR2_X1 U1064 ( .A(n1274), .B(n1342), .Z(n1115) );
NOR2_X1 U1065 ( .A1(G113), .A2(KEYINPUT15), .ZN(n1342) );
XNOR2_X1 U1066 ( .A(G119), .B(n1239), .ZN(n1274) );
INV_X1 U1067 ( .A(G116), .ZN(n1239) );
NAND2_X1 U1068 ( .A1(n1072), .A2(n1343), .ZN(n1208) );
NAND4_X1 U1069 ( .A1(G953), .A2(G902), .A3(n1228), .A4(n1114), .ZN(n1343) );
INV_X1 U1070 ( .A(G898), .ZN(n1114) );
NAND3_X1 U1071 ( .A1(n1228), .A2(n1040), .A3(G952), .ZN(n1072) );
NAND2_X1 U1072 ( .A1(G237), .A2(G234), .ZN(n1228) );
XNOR2_X1 U1073 ( .A(n1057), .B(KEYINPUT42), .ZN(n1224) );
INV_X1 U1074 ( .A(n1212), .ZN(n1057) );
NOR2_X1 U1075 ( .A1(n1060), .A2(n1059), .ZN(n1212) );
INV_X1 U1076 ( .A(n1243), .ZN(n1059) );
NAND2_X1 U1077 ( .A1(n1344), .A2(n1263), .ZN(n1243) );
NAND2_X1 U1078 ( .A1(G234), .A2(n1250), .ZN(n1263) );
XOR2_X1 U1079 ( .A(KEYINPUT36), .B(G221), .Z(n1344) );
XOR2_X1 U1080 ( .A(n1345), .B(G469), .Z(n1060) );
NAND2_X1 U1081 ( .A1(n1346), .A2(n1250), .ZN(n1345) );
INV_X1 U1082 ( .A(G902), .ZN(n1250) );
XNOR2_X1 U1083 ( .A(n1258), .B(n1347), .ZN(n1346) );
XNOR2_X1 U1084 ( .A(n1155), .B(G110), .ZN(n1347) );
XNOR2_X1 U1085 ( .A(n1348), .B(n1349), .ZN(n1155) );
XOR2_X1 U1086 ( .A(n1350), .B(n1269), .Z(n1349) );
XNOR2_X1 U1087 ( .A(n1351), .B(n1104), .ZN(n1269) );
INV_X1 U1088 ( .A(G131), .ZN(n1104) );
NAND2_X1 U1089 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
NAND2_X1 U1090 ( .A1(G134), .A2(n1354), .ZN(n1353) );
XOR2_X1 U1091 ( .A(KEYINPUT1), .B(n1355), .Z(n1352) );
NOR2_X1 U1092 ( .A1(G134), .A2(n1354), .ZN(n1355) );
INV_X1 U1093 ( .A(G137), .ZN(n1354) );
NAND2_X1 U1094 ( .A1(KEYINPUT6), .A2(n1225), .ZN(n1350) );
INV_X1 U1095 ( .A(G101), .ZN(n1225) );
XOR2_X1 U1096 ( .A(n1356), .B(n1357), .Z(n1348) );
XOR2_X1 U1097 ( .A(n1358), .B(n1102), .Z(n1357) );
NAND2_X1 U1098 ( .A1(KEYINPUT39), .A2(n1359), .ZN(n1102) );
XNOR2_X1 U1099 ( .A(n1360), .B(n1336), .ZN(n1359) );
XOR2_X1 U1100 ( .A(G143), .B(KEYINPUT56), .Z(n1336) );
NAND2_X1 U1101 ( .A1(KEYINPUT18), .A2(G146), .ZN(n1360) );
NAND3_X1 U1102 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1358) );
OR2_X1 U1103 ( .A1(n1032), .A2(KEYINPUT4), .ZN(n1363) );
NAND3_X1 U1104 ( .A1(KEYINPUT4), .A2(n1032), .A3(G104), .ZN(n1362) );
INV_X1 U1105 ( .A(G107), .ZN(n1032) );
NAND2_X1 U1106 ( .A1(n1364), .A2(n1140), .ZN(n1361) );
INV_X1 U1107 ( .A(G104), .ZN(n1140) );
NAND2_X1 U1108 ( .A1(n1365), .A2(KEYINPUT4), .ZN(n1364) );
XNOR2_X1 U1109 ( .A(G107), .B(KEYINPUT33), .ZN(n1365) );
NAND2_X1 U1110 ( .A1(G227), .A2(n1040), .ZN(n1356) );
INV_X1 U1111 ( .A(G953), .ZN(n1040) );
XNOR2_X1 U1112 ( .A(G140), .B(n1222), .ZN(n1258) );
INV_X1 U1113 ( .A(G128), .ZN(n1222) );
INV_X1 U1114 ( .A(G110), .ZN(n1162) );
endmodule


