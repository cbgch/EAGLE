//Key = 0110001000110000101001111000000111011100111101000111000011000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
n1365, n1366;

XNOR2_X1 U757 ( .A(n1045), .B(n1046), .ZN(G9) );
NAND4_X1 U758 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(G75) );
NOR3_X1 U759 ( .A1(n1051), .A2(G953), .A3(n1052), .ZN(n1050) );
NOR4_X1 U760 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NAND3_X1 U761 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1053) );
OR2_X1 U762 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND3_X1 U763 ( .A1(n1062), .A2(n1063), .A3(n1060), .ZN(n1057) );
NOR4_X1 U764 ( .A1(n1064), .A2(n1056), .A3(n1065), .A4(n1066), .ZN(n1051) );
NAND4_X1 U765 ( .A1(n1067), .A2(n1068), .A3(n1060), .A4(n1069), .ZN(n1064) );
XOR2_X1 U766 ( .A(n1070), .B(n1071), .Z(n1068) );
XNOR2_X1 U767 ( .A(G472), .B(KEYINPUT61), .ZN(n1071) );
XNOR2_X1 U768 ( .A(n1072), .B(n1073), .ZN(n1067) );
NOR2_X1 U769 ( .A1(n1074), .A2(KEYINPUT29), .ZN(n1073) );
NAND3_X1 U770 ( .A1(n1061), .A2(n1075), .A3(n1059), .ZN(n1048) );
INV_X1 U771 ( .A(n1076), .ZN(n1059) );
NAND2_X1 U772 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND3_X1 U773 ( .A1(n1079), .A2(n1080), .A3(n1081), .ZN(n1078) );
NAND3_X1 U774 ( .A1(n1082), .A2(n1060), .A3(n1083), .ZN(n1077) );
NAND2_X1 U775 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1081), .A2(n1086), .ZN(n1085) );
NAND2_X1 U777 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
OR2_X1 U778 ( .A1(n1066), .A2(n1069), .ZN(n1088) );
NAND2_X1 U779 ( .A1(n1079), .A2(n1089), .ZN(n1084) );
NAND2_X1 U780 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XOR2_X1 U781 ( .A(n1092), .B(n1093), .Z(G72) );
XOR2_X1 U782 ( .A(n1094), .B(n1095), .Z(n1093) );
NAND2_X1 U783 ( .A1(G953), .A2(n1096), .ZN(n1095) );
NAND2_X1 U784 ( .A1(G900), .A2(G227), .ZN(n1096) );
NAND2_X1 U785 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
NAND2_X1 U786 ( .A1(G953), .A2(n1099), .ZN(n1098) );
XOR2_X1 U787 ( .A(n1100), .B(n1101), .Z(n1097) );
XNOR2_X1 U788 ( .A(n1102), .B(n1103), .ZN(n1101) );
NOR2_X1 U789 ( .A1(KEYINPUT54), .A2(n1104), .ZN(n1103) );
NAND2_X1 U790 ( .A1(KEYINPUT50), .A2(n1105), .ZN(n1102) );
XNOR2_X1 U791 ( .A(n1106), .B(n1107), .ZN(n1105) );
NOR2_X1 U792 ( .A1(n1047), .A2(G953), .ZN(n1092) );
XOR2_X1 U793 ( .A(n1108), .B(n1109), .Z(G69) );
NOR2_X1 U794 ( .A1(n1049), .A2(G953), .ZN(n1109) );
NAND2_X1 U795 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NAND2_X1 U796 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NAND2_X1 U797 ( .A1(G953), .A2(n1114), .ZN(n1113) );
XNOR2_X1 U798 ( .A(KEYINPUT57), .B(n1115), .ZN(n1112) );
NAND2_X1 U799 ( .A1(G953), .A2(n1116), .ZN(n1110) );
NAND2_X1 U800 ( .A1(G898), .A2(n1117), .ZN(n1116) );
NAND2_X1 U801 ( .A1(n1118), .A2(n1114), .ZN(n1117) );
XOR2_X1 U802 ( .A(n1115), .B(KEYINPUT57), .Z(n1118) );
NAND3_X1 U803 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1115) );
NAND2_X1 U804 ( .A1(KEYINPUT39), .A2(n1122), .ZN(n1121) );
NAND3_X1 U805 ( .A1(n1123), .A2(n1124), .A3(n1125), .ZN(n1120) );
INV_X1 U806 ( .A(KEYINPUT39), .ZN(n1124) );
OR2_X1 U807 ( .A1(n1125), .A2(n1123), .ZN(n1119) );
NOR2_X1 U808 ( .A1(KEYINPUT60), .A2(n1122), .ZN(n1123) );
NOR2_X1 U809 ( .A1(n1126), .A2(n1127), .ZN(G66) );
XOR2_X1 U810 ( .A(KEYINPUT48), .B(n1128), .Z(n1127) );
XOR2_X1 U811 ( .A(n1129), .B(n1130), .Z(n1126) );
NOR2_X1 U812 ( .A1(KEYINPUT28), .A2(n1131), .ZN(n1130) );
XNOR2_X1 U813 ( .A(n1132), .B(n1133), .ZN(n1131) );
NAND3_X1 U814 ( .A1(n1134), .A2(G217), .A3(KEYINPUT49), .ZN(n1129) );
NOR2_X1 U815 ( .A1(n1128), .A2(n1135), .ZN(G63) );
XNOR2_X1 U816 ( .A(n1136), .B(n1137), .ZN(n1135) );
AND2_X1 U817 ( .A1(G478), .A2(n1134), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1128), .A2(n1138), .ZN(G60) );
XOR2_X1 U819 ( .A(n1139), .B(n1140), .Z(n1138) );
AND2_X1 U820 ( .A1(G475), .A2(n1134), .ZN(n1139) );
XOR2_X1 U821 ( .A(G104), .B(n1141), .Z(G6) );
NOR2_X1 U822 ( .A1(n1128), .A2(n1142), .ZN(G57) );
XOR2_X1 U823 ( .A(n1143), .B(n1144), .Z(n1142) );
NOR2_X1 U824 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
XOR2_X1 U825 ( .A(n1147), .B(KEYINPUT22), .Z(n1146) );
NAND3_X1 U826 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
XOR2_X1 U827 ( .A(KEYINPUT38), .B(n1151), .Z(n1150) );
NOR2_X1 U828 ( .A1(n1152), .A2(n1151), .ZN(n1145) );
NOR2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1151) );
INV_X1 U830 ( .A(G472), .ZN(n1153) );
AND2_X1 U831 ( .A1(n1149), .A2(n1148), .ZN(n1152) );
NAND2_X1 U832 ( .A1(n1155), .A2(n1156), .ZN(n1148) );
XOR2_X1 U833 ( .A(n1157), .B(n1158), .Z(n1155) );
NAND2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1149) );
XNOR2_X1 U835 ( .A(n1158), .B(n1157), .ZN(n1160) );
NOR2_X1 U836 ( .A1(KEYINPUT14), .A2(n1161), .ZN(n1158) );
XNOR2_X1 U837 ( .A(KEYINPUT25), .B(n1156), .ZN(n1159) );
XNOR2_X1 U838 ( .A(n1162), .B(G101), .ZN(n1143) );
NOR2_X1 U839 ( .A1(n1128), .A2(n1163), .ZN(G54) );
XOR2_X1 U840 ( .A(n1164), .B(n1165), .Z(n1163) );
XOR2_X1 U841 ( .A(G140), .B(G110), .Z(n1165) );
XOR2_X1 U842 ( .A(n1166), .B(n1167), .Z(n1164) );
NAND3_X1 U843 ( .A1(n1134), .A2(G469), .A3(KEYINPUT45), .ZN(n1166) );
INV_X1 U844 ( .A(n1154), .ZN(n1134) );
NOR2_X1 U845 ( .A1(n1128), .A2(n1168), .ZN(G51) );
XOR2_X1 U846 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U847 ( .A(n1171), .B(n1172), .Z(n1170) );
NOR2_X1 U848 ( .A1(KEYINPUT9), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U849 ( .A(n1174), .B(n1175), .ZN(n1173) );
NOR2_X1 U850 ( .A1(n1072), .A2(n1154), .ZN(n1169) );
NAND2_X1 U851 ( .A1(G902), .A2(n1176), .ZN(n1154) );
NAND2_X1 U852 ( .A1(n1047), .A2(n1177), .ZN(n1176) );
XOR2_X1 U853 ( .A(KEYINPUT47), .B(n1049), .Z(n1177) );
AND4_X1 U854 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1049) );
NOR4_X1 U855 ( .A1(n1182), .A2(n1183), .A3(n1141), .A4(n1184), .ZN(n1181) );
NOR4_X1 U856 ( .A1(n1185), .A2(n1186), .A3(n1062), .A4(n1090), .ZN(n1184) );
NOR2_X1 U857 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
INV_X1 U858 ( .A(KEYINPUT4), .ZN(n1188) );
NOR3_X1 U859 ( .A1(n1055), .A2(n1189), .A3(n1080), .ZN(n1187) );
NOR2_X1 U860 ( .A1(KEYINPUT4), .A2(n1190), .ZN(n1185) );
NOR3_X1 U861 ( .A1(n1191), .A2(n1192), .A3(n1090), .ZN(n1141) );
NOR3_X1 U862 ( .A1(n1056), .A2(n1191), .A3(n1063), .ZN(n1183) );
NOR2_X1 U863 ( .A1(n1046), .A2(n1193), .ZN(n1180) );
NOR3_X1 U864 ( .A1(n1091), .A2(n1192), .A3(n1191), .ZN(n1046) );
INV_X1 U865 ( .A(n1194), .ZN(n1191) );
NAND3_X1 U866 ( .A1(n1195), .A2(n1194), .A3(n1081), .ZN(n1178) );
AND4_X1 U867 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1047) );
NOR4_X1 U868 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199) );
NOR2_X1 U869 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
INV_X1 U870 ( .A(KEYINPUT21), .ZN(n1205) );
NOR2_X1 U871 ( .A1(KEYINPUT46), .A2(n1206), .ZN(n1202) );
NOR3_X1 U872 ( .A1(n1207), .A2(n1056), .A3(n1208), .ZN(n1201) );
NOR2_X1 U873 ( .A1(n1209), .A2(n1210), .ZN(n1200) );
NOR2_X1 U874 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
NOR4_X1 U875 ( .A1(KEYINPUT21), .A2(n1079), .A3(n1063), .A4(n1090), .ZN(n1212) );
NOR3_X1 U876 ( .A1(n1213), .A2(n1087), .A3(n1214), .ZN(n1211) );
INV_X1 U877 ( .A(KEYINPUT46), .ZN(n1214) );
NAND3_X1 U878 ( .A1(n1215), .A2(n1062), .A3(n1216), .ZN(n1213) );
NOR3_X1 U879 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1198) );
NOR2_X1 U880 ( .A1(n1220), .A2(G952), .ZN(n1128) );
XNOR2_X1 U881 ( .A(G146), .B(n1196), .ZN(G48) );
NAND3_X1 U882 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1196) );
NAND2_X1 U883 ( .A1(n1224), .A2(n1225), .ZN(G45) );
NAND2_X1 U884 ( .A1(n1226), .A2(n1206), .ZN(n1225) );
XOR2_X1 U885 ( .A(KEYINPUT10), .B(n1227), .Z(n1224) );
NOR2_X1 U886 ( .A1(n1206), .A2(n1226), .ZN(n1227) );
XNOR2_X1 U887 ( .A(KEYINPUT55), .B(n1106), .ZN(n1226) );
NAND3_X1 U888 ( .A1(n1228), .A2(n1195), .A3(n1229), .ZN(n1206) );
NOR3_X1 U889 ( .A1(n1087), .A2(n1230), .A3(n1231), .ZN(n1229) );
INV_X1 U890 ( .A(n1210), .ZN(n1228) );
XNOR2_X1 U891 ( .A(G140), .B(n1197), .ZN(G42) );
OR3_X1 U892 ( .A1(n1090), .A2(n1063), .A3(n1207), .ZN(n1197) );
INV_X1 U893 ( .A(n1232), .ZN(n1063) );
XOR2_X1 U894 ( .A(G137), .B(n1233), .Z(G39) );
NOR3_X1 U895 ( .A1(n1234), .A2(n1208), .A3(n1207), .ZN(n1233) );
XNOR2_X1 U896 ( .A(KEYINPUT42), .B(n1056), .ZN(n1234) );
NAND3_X1 U897 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(G36) );
NAND2_X1 U898 ( .A1(n1217), .A2(n1238), .ZN(n1237) );
NAND2_X1 U899 ( .A1(n1239), .A2(n1240), .ZN(n1236) );
INV_X1 U900 ( .A(KEYINPUT16), .ZN(n1240) );
NAND2_X1 U901 ( .A1(n1241), .A2(G134), .ZN(n1239) );
XNOR2_X1 U902 ( .A(KEYINPUT13), .B(n1217), .ZN(n1241) );
NAND2_X1 U903 ( .A1(KEYINPUT16), .A2(n1242), .ZN(n1235) );
NAND2_X1 U904 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
OR3_X1 U905 ( .A1(n1238), .A2(n1217), .A3(KEYINPUT13), .ZN(n1244) );
NAND2_X1 U906 ( .A1(KEYINPUT13), .A2(n1217), .ZN(n1243) );
NOR3_X1 U907 ( .A1(n1062), .A2(n1091), .A3(n1207), .ZN(n1217) );
XOR2_X1 U908 ( .A(G131), .B(n1219), .Z(G33) );
NOR3_X1 U909 ( .A1(n1090), .A2(n1062), .A3(n1207), .ZN(n1219) );
NAND4_X1 U910 ( .A1(n1083), .A2(n1222), .A3(n1245), .A4(n1060), .ZN(n1207) );
INV_X1 U911 ( .A(n1087), .ZN(n1222) );
INV_X1 U912 ( .A(n1054), .ZN(n1083) );
XOR2_X1 U913 ( .A(G128), .B(n1218), .Z(G30) );
NOR4_X1 U914 ( .A1(n1210), .A2(n1208), .A3(n1091), .A4(n1087), .ZN(n1218) );
XNOR2_X1 U915 ( .A(G101), .B(n1246), .ZN(G3) );
NAND4_X1 U916 ( .A1(KEYINPUT43), .A2(n1081), .A3(n1247), .A4(n1248), .ZN(n1246) );
NOR3_X1 U917 ( .A1(n1062), .A2(n1189), .A3(n1087), .ZN(n1248) );
XNOR2_X1 U918 ( .A(n1080), .B(KEYINPUT41), .ZN(n1247) );
XOR2_X1 U919 ( .A(n1204), .B(n1249), .Z(G27) );
NAND2_X1 U920 ( .A1(KEYINPUT33), .A2(G125), .ZN(n1249) );
NAND3_X1 U921 ( .A1(n1232), .A2(n1079), .A3(n1223), .ZN(n1204) );
NOR2_X1 U922 ( .A1(n1210), .A2(n1090), .ZN(n1223) );
NAND2_X1 U923 ( .A1(n1080), .A2(n1245), .ZN(n1210) );
NAND2_X1 U924 ( .A1(n1076), .A2(n1250), .ZN(n1245) );
NAND4_X1 U925 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1099), .ZN(n1250) );
INV_X1 U926 ( .A(G900), .ZN(n1099) );
INV_X1 U927 ( .A(n1252), .ZN(n1080) );
INV_X1 U928 ( .A(n1055), .ZN(n1079) );
XNOR2_X1 U929 ( .A(G122), .B(n1179), .ZN(G24) );
NAND4_X1 U930 ( .A1(n1190), .A2(n1061), .A3(n1216), .A4(n1215), .ZN(n1179) );
INV_X1 U931 ( .A(n1192), .ZN(n1061) );
NAND2_X1 U932 ( .A1(n1253), .A2(n1254), .ZN(n1192) );
XNOR2_X1 U933 ( .A(KEYINPUT12), .B(n1255), .ZN(n1254) );
XOR2_X1 U934 ( .A(G119), .B(n1193), .Z(G21) );
NOR3_X1 U935 ( .A1(n1056), .A2(n1256), .A3(n1208), .ZN(n1193) );
INV_X1 U936 ( .A(n1221), .ZN(n1208) );
NOR2_X1 U937 ( .A1(n1257), .A2(n1253), .ZN(n1221) );
XOR2_X1 U938 ( .A(G116), .B(n1182), .Z(G18) );
NOR3_X1 U939 ( .A1(n1062), .A2(n1091), .A3(n1256), .ZN(n1182) );
NAND2_X1 U940 ( .A1(n1230), .A2(n1216), .ZN(n1091) );
INV_X1 U941 ( .A(n1215), .ZN(n1230) );
XNOR2_X1 U942 ( .A(G113), .B(n1258), .ZN(G15) );
OR3_X1 U943 ( .A1(n1256), .A2(n1062), .A3(n1090), .ZN(n1258) );
NAND2_X1 U944 ( .A1(n1231), .A2(n1215), .ZN(n1090) );
INV_X1 U945 ( .A(n1216), .ZN(n1231) );
INV_X1 U946 ( .A(n1195), .ZN(n1062) );
NOR2_X1 U947 ( .A1(n1255), .A2(n1253), .ZN(n1195) );
INV_X1 U948 ( .A(n1259), .ZN(n1253) );
INV_X1 U949 ( .A(n1257), .ZN(n1255) );
INV_X1 U950 ( .A(n1190), .ZN(n1256) );
NOR3_X1 U951 ( .A1(n1252), .A2(n1189), .A3(n1055), .ZN(n1190) );
NAND2_X1 U952 ( .A1(n1260), .A2(n1261), .ZN(n1055) );
XNOR2_X1 U953 ( .A(n1066), .B(KEYINPUT8), .ZN(n1260) );
XNOR2_X1 U954 ( .A(G110), .B(n1262), .ZN(G12) );
NAND3_X1 U955 ( .A1(n1194), .A2(n1263), .A3(n1232), .ZN(n1262) );
NOR2_X1 U956 ( .A1(n1259), .A2(n1257), .ZN(n1232) );
XOR2_X1 U957 ( .A(n1065), .B(KEYINPUT24), .Z(n1257) );
XNOR2_X1 U958 ( .A(n1264), .B(n1265), .ZN(n1065) );
AND2_X1 U959 ( .A1(n1266), .A2(G217), .ZN(n1265) );
NAND2_X1 U960 ( .A1(n1267), .A2(n1268), .ZN(n1264) );
XNOR2_X1 U961 ( .A(n1133), .B(n1269), .ZN(n1267) );
INV_X1 U962 ( .A(n1132), .ZN(n1269) );
XNOR2_X1 U963 ( .A(n1270), .B(G137), .ZN(n1132) );
NAND2_X1 U964 ( .A1(n1271), .A2(G221), .ZN(n1270) );
XNOR2_X1 U965 ( .A(n1272), .B(n1273), .ZN(n1133) );
NOR3_X1 U966 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1273) );
NOR2_X1 U967 ( .A1(n1277), .A2(n1278), .ZN(n1276) );
NOR2_X1 U968 ( .A1(n1279), .A2(G110), .ZN(n1277) );
NOR2_X1 U969 ( .A1(n1280), .A2(n1281), .ZN(n1279) );
NOR4_X1 U970 ( .A1(KEYINPUT7), .A2(n1280), .A3(KEYINPUT3), .A4(G110), .ZN(n1275) );
INV_X1 U971 ( .A(n1282), .ZN(n1280) );
NOR2_X1 U972 ( .A1(n1283), .A2(n1282), .ZN(n1274) );
XNOR2_X1 U973 ( .A(n1284), .B(G128), .ZN(n1282) );
NAND2_X1 U974 ( .A1(KEYINPUT6), .A2(n1285), .ZN(n1284) );
XOR2_X1 U975 ( .A(KEYINPUT18), .B(G119), .Z(n1285) );
NOR3_X1 U976 ( .A1(n1286), .A2(n1287), .A3(n1288), .ZN(n1283) );
NOR2_X1 U977 ( .A1(n1289), .A2(n1290), .ZN(n1288) );
INV_X1 U978 ( .A(KEYINPUT2), .ZN(n1290) );
NOR2_X1 U979 ( .A1(n1291), .A2(G110), .ZN(n1289) );
NOR2_X1 U980 ( .A1(KEYINPUT7), .A2(n1281), .ZN(n1291) );
INV_X1 U981 ( .A(KEYINPUT3), .ZN(n1281) );
NOR2_X1 U982 ( .A1(KEYINPUT2), .A2(G110), .ZN(n1287) );
NOR2_X1 U983 ( .A1(KEYINPUT3), .A2(n1278), .ZN(n1286) );
INV_X1 U984 ( .A(KEYINPUT7), .ZN(n1278) );
NAND2_X1 U985 ( .A1(KEYINPUT37), .A2(n1292), .ZN(n1272) );
XOR2_X1 U986 ( .A(n1293), .B(n1104), .Z(n1292) );
XOR2_X1 U987 ( .A(G125), .B(G140), .Z(n1104) );
NOR2_X1 U988 ( .A1(KEYINPUT62), .A2(n1294), .ZN(n1293) );
NAND2_X1 U989 ( .A1(n1295), .A2(n1296), .ZN(n1259) );
NAND2_X1 U990 ( .A1(G472), .A2(n1070), .ZN(n1296) );
XOR2_X1 U991 ( .A(KEYINPUT56), .B(n1297), .Z(n1295) );
NOR2_X1 U992 ( .A1(G472), .A2(n1070), .ZN(n1297) );
NAND2_X1 U993 ( .A1(n1298), .A2(n1268), .ZN(n1070) );
XOR2_X1 U994 ( .A(n1299), .B(n1300), .Z(n1298) );
XOR2_X1 U995 ( .A(G101), .B(n1301), .Z(n1300) );
NOR2_X1 U996 ( .A1(KEYINPUT58), .A2(n1302), .ZN(n1301) );
XOR2_X1 U997 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U998 ( .A(n1305), .B(n1156), .ZN(n1299) );
NAND2_X1 U999 ( .A1(KEYINPUT23), .A2(n1162), .ZN(n1305) );
AND3_X1 U1000 ( .A1(n1306), .A2(n1220), .A3(G210), .ZN(n1162) );
XNOR2_X1 U1001 ( .A(KEYINPUT0), .B(n1056), .ZN(n1263) );
INV_X1 U1002 ( .A(n1081), .ZN(n1056) );
NOR2_X1 U1003 ( .A1(n1216), .A2(n1215), .ZN(n1081) );
XNOR2_X1 U1004 ( .A(n1307), .B(G475), .ZN(n1215) );
OR2_X1 U1005 ( .A1(n1140), .A2(G902), .ZN(n1307) );
XNOR2_X1 U1006 ( .A(n1308), .B(n1309), .ZN(n1140) );
XOR2_X1 U1007 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1008 ( .A(n1312), .B(n1313), .ZN(n1311) );
NOR2_X1 U1009 ( .A1(G140), .A2(KEYINPUT17), .ZN(n1313) );
NOR2_X1 U1010 ( .A1(KEYINPUT5), .A2(n1314), .ZN(n1312) );
XNOR2_X1 U1011 ( .A(n1315), .B(n1316), .ZN(n1314) );
NAND2_X1 U1012 ( .A1(KEYINPUT1), .A2(n1317), .ZN(n1315) );
NAND2_X1 U1013 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND2_X1 U1014 ( .A1(n1320), .A2(n1106), .ZN(n1319) );
XOR2_X1 U1015 ( .A(n1321), .B(KEYINPUT20), .Z(n1318) );
NAND2_X1 U1016 ( .A1(G143), .A2(n1322), .ZN(n1321) );
XNOR2_X1 U1017 ( .A(KEYINPUT53), .B(n1320), .ZN(n1322) );
NAND3_X1 U1018 ( .A1(n1306), .A2(n1220), .A3(G214), .ZN(n1320) );
XNOR2_X1 U1019 ( .A(G113), .B(G104), .ZN(n1310) );
XOR2_X1 U1020 ( .A(n1323), .B(n1324), .Z(n1308) );
XNOR2_X1 U1021 ( .A(KEYINPUT52), .B(n1294), .ZN(n1324) );
XNOR2_X1 U1022 ( .A(G122), .B(G125), .ZN(n1323) );
XNOR2_X1 U1023 ( .A(n1325), .B(G478), .ZN(n1216) );
NAND2_X1 U1024 ( .A1(n1136), .A2(n1268), .ZN(n1325) );
XNOR2_X1 U1025 ( .A(n1326), .B(n1327), .ZN(n1136) );
XOR2_X1 U1026 ( .A(n1328), .B(n1329), .Z(n1327) );
XOR2_X1 U1027 ( .A(G128), .B(G122), .Z(n1329) );
XNOR2_X1 U1028 ( .A(KEYINPUT63), .B(n1238), .ZN(n1328) );
INV_X1 U1029 ( .A(G134), .ZN(n1238) );
XOR2_X1 U1030 ( .A(n1330), .B(n1331), .Z(n1326) );
XOR2_X1 U1031 ( .A(n1332), .B(n1333), .Z(n1331) );
NAND2_X1 U1032 ( .A1(KEYINPUT35), .A2(G143), .ZN(n1333) );
NAND2_X1 U1033 ( .A1(G217), .A2(n1271), .ZN(n1332) );
AND2_X1 U1034 ( .A1(G234), .A2(n1220), .ZN(n1271) );
XNOR2_X1 U1035 ( .A(G116), .B(G107), .ZN(n1330) );
NOR3_X1 U1036 ( .A1(n1252), .A2(n1189), .A3(n1087), .ZN(n1194) );
NAND2_X1 U1037 ( .A1(n1066), .A2(n1261), .ZN(n1087) );
XNOR2_X1 U1038 ( .A(n1069), .B(KEYINPUT32), .ZN(n1261) );
NAND2_X1 U1039 ( .A1(G221), .A2(n1266), .ZN(n1069) );
NAND2_X1 U1040 ( .A1(G234), .A2(n1268), .ZN(n1266) );
XNOR2_X1 U1041 ( .A(n1334), .B(G469), .ZN(n1066) );
NAND2_X1 U1042 ( .A1(n1335), .A2(n1268), .ZN(n1334) );
XNOR2_X1 U1043 ( .A(n1167), .B(n1336), .ZN(n1335) );
XOR2_X1 U1044 ( .A(G140), .B(n1337), .Z(n1336) );
NOR2_X1 U1045 ( .A1(G110), .A2(KEYINPUT34), .ZN(n1337) );
XNOR2_X1 U1046 ( .A(n1338), .B(n1339), .ZN(n1167) );
XOR2_X1 U1047 ( .A(n1340), .B(n1341), .Z(n1339) );
XNOR2_X1 U1048 ( .A(n1045), .B(G104), .ZN(n1341) );
XNOR2_X1 U1049 ( .A(KEYINPUT19), .B(n1106), .ZN(n1340) );
XOR2_X1 U1050 ( .A(n1304), .B(n1342), .Z(n1338) );
XOR2_X1 U1051 ( .A(n1343), .B(n1344), .Z(n1342) );
NOR2_X1 U1052 ( .A1(G101), .A2(KEYINPUT59), .ZN(n1344) );
AND2_X1 U1053 ( .A1(n1220), .A2(G227), .ZN(n1343) );
XOR2_X1 U1054 ( .A(n1157), .B(n1107), .Z(n1304) );
XOR2_X1 U1055 ( .A(n1100), .B(KEYINPUT15), .Z(n1157) );
XOR2_X1 U1056 ( .A(n1345), .B(n1346), .Z(n1100) );
XOR2_X1 U1057 ( .A(KEYINPUT31), .B(G137), .Z(n1346) );
XNOR2_X1 U1058 ( .A(G134), .B(n1316), .ZN(n1345) );
XOR2_X1 U1059 ( .A(G131), .B(KEYINPUT26), .Z(n1316) );
AND2_X1 U1060 ( .A1(n1347), .A2(n1076), .ZN(n1189) );
NAND3_X1 U1061 ( .A1(n1251), .A2(n1220), .A3(G952), .ZN(n1076) );
INV_X1 U1062 ( .A(G953), .ZN(n1220) );
NAND4_X1 U1063 ( .A1(G953), .A2(G902), .A3(n1251), .A4(n1348), .ZN(n1347) );
INV_X1 U1064 ( .A(G898), .ZN(n1348) );
NAND2_X1 U1065 ( .A1(G237), .A2(G234), .ZN(n1251) );
NAND2_X1 U1066 ( .A1(n1054), .A2(n1060), .ZN(n1252) );
NAND2_X1 U1067 ( .A1(G214), .A2(n1349), .ZN(n1060) );
XNOR2_X1 U1068 ( .A(n1074), .B(n1072), .ZN(n1054) );
NAND2_X1 U1069 ( .A1(G210), .A2(n1349), .ZN(n1072) );
NAND2_X1 U1070 ( .A1(n1306), .A2(n1268), .ZN(n1349) );
INV_X1 U1071 ( .A(G237), .ZN(n1306) );
AND3_X1 U1072 ( .A1(n1350), .A2(n1268), .A3(n1351), .ZN(n1074) );
XOR2_X1 U1073 ( .A(KEYINPUT36), .B(n1352), .Z(n1351) );
NOR2_X1 U1074 ( .A1(n1171), .A2(n1353), .ZN(n1352) );
INV_X1 U1075 ( .A(G902), .ZN(n1268) );
NAND2_X1 U1076 ( .A1(n1171), .A2(n1353), .ZN(n1350) );
XNOR2_X1 U1077 ( .A(n1354), .B(KEYINPUT44), .ZN(n1353) );
NAND2_X1 U1078 ( .A1(n1355), .A2(n1356), .ZN(n1354) );
NAND2_X1 U1079 ( .A1(n1175), .A2(n1161), .ZN(n1356) );
INV_X1 U1080 ( .A(n1174), .ZN(n1161) );
NAND2_X1 U1081 ( .A1(n1357), .A2(n1174), .ZN(n1355) );
XNOR2_X1 U1082 ( .A(n1303), .B(n1107), .ZN(n1174) );
XNOR2_X1 U1083 ( .A(G128), .B(n1294), .ZN(n1107) );
INV_X1 U1084 ( .A(G146), .ZN(n1294) );
NAND2_X1 U1085 ( .A1(KEYINPUT51), .A2(n1106), .ZN(n1303) );
INV_X1 U1086 ( .A(G143), .ZN(n1106) );
XNOR2_X1 U1087 ( .A(KEYINPUT30), .B(n1175), .ZN(n1357) );
XNOR2_X1 U1088 ( .A(G125), .B(n1358), .ZN(n1175) );
NOR2_X1 U1089 ( .A1(G953), .A2(n1114), .ZN(n1358) );
INV_X1 U1090 ( .A(G224), .ZN(n1114) );
AND2_X1 U1091 ( .A1(n1359), .A2(n1360), .ZN(n1171) );
NAND2_X1 U1092 ( .A1(n1125), .A2(n1122), .ZN(n1360) );
XOR2_X1 U1093 ( .A(n1361), .B(KEYINPUT27), .Z(n1359) );
OR2_X1 U1094 ( .A1(n1122), .A2(n1125), .ZN(n1361) );
XNOR2_X1 U1095 ( .A(n1362), .B(n1363), .ZN(n1125) );
XNOR2_X1 U1096 ( .A(G104), .B(n1364), .ZN(n1363) );
NAND2_X1 U1097 ( .A1(KEYINPUT40), .A2(G101), .ZN(n1364) );
XNOR2_X1 U1098 ( .A(n1365), .B(n1156), .ZN(n1362) );
XNOR2_X1 U1099 ( .A(G113), .B(n1366), .ZN(n1156) );
XOR2_X1 U1100 ( .A(G119), .B(G116), .Z(n1366) );
NAND2_X1 U1101 ( .A1(KEYINPUT11), .A2(n1045), .ZN(n1365) );
INV_X1 U1102 ( .A(G107), .ZN(n1045) );
XOR2_X1 U1103 ( .A(G122), .B(G110), .Z(n1122) );
endmodule


