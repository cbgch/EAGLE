//Key = 1011101111111000000010110100010001111111001011111010101111110000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279;

XOR2_X1 U717 ( .A(n982), .B(n983), .Z(G9) );
XOR2_X1 U718 ( .A(KEYINPUT15), .B(G107), .Z(n983) );
NOR2_X1 U719 ( .A1(n984), .A2(n985), .ZN(G75) );
NOR4_X1 U720 ( .A1(G953), .A2(n986), .A3(n987), .A4(n988), .ZN(n985) );
NOR2_X1 U721 ( .A1(n989), .A2(n990), .ZN(n987) );
NOR2_X1 U722 ( .A1(n991), .A2(n992), .ZN(n989) );
NOR3_X1 U723 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n992) );
NOR2_X1 U724 ( .A1(n996), .A2(n997), .ZN(n995) );
NOR2_X1 U725 ( .A1(n998), .A2(n999), .ZN(n997) );
NOR2_X1 U726 ( .A1(n1000), .A2(n1001), .ZN(n998) );
NOR2_X1 U727 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
NOR2_X1 U728 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NOR2_X1 U729 ( .A1(n1006), .A2(n1007), .ZN(n1004) );
NOR2_X1 U730 ( .A1(n1008), .A2(n1009), .ZN(n1000) );
NOR2_X1 U731 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR3_X1 U732 ( .A1(n1009), .A2(n1012), .A3(n1003), .ZN(n996) );
NOR2_X1 U733 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
NOR4_X1 U734 ( .A1(n1015), .A2(n1003), .A3(n1009), .A4(n999), .ZN(n991) );
INV_X1 U735 ( .A(n1016), .ZN(n999) );
XNOR2_X1 U736 ( .A(n994), .B(n993), .ZN(n1015) );
NOR3_X1 U737 ( .A1(n986), .A2(G953), .A3(G952), .ZN(n984) );
AND4_X1 U738 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n986) );
NOR4_X1 U739 ( .A1(n1021), .A2(n1022), .A3(n1023), .A4(n994), .ZN(n1020) );
INV_X1 U740 ( .A(n1007), .ZN(n1023) );
NAND3_X1 U741 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1021) );
NAND2_X1 U742 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NOR3_X1 U743 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1019) );
XNOR2_X1 U744 ( .A(n993), .B(KEYINPUT36), .ZN(n1031) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
XOR2_X1 U746 ( .A(G472), .B(n1034), .Z(n1029) );
NOR2_X1 U747 ( .A1(KEYINPUT26), .A2(n1035), .ZN(n1034) );
XOR2_X1 U748 ( .A(n1036), .B(KEYINPUT32), .Z(n1018) );
OR2_X1 U749 ( .A1(n1028), .A2(n1027), .ZN(n1036) );
XNOR2_X1 U750 ( .A(n1037), .B(KEYINPUT63), .ZN(n1017) );
XOR2_X1 U751 ( .A(n1038), .B(n1039), .Z(G72) );
NOR2_X1 U752 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NOR3_X1 U753 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
NOR2_X1 U754 ( .A1(G953), .A2(n1045), .ZN(n1040) );
XNOR2_X1 U755 ( .A(n1046), .B(n1044), .ZN(n1045) );
NAND3_X1 U756 ( .A1(n1047), .A2(n1048), .A3(KEYINPUT29), .ZN(n1044) );
OR3_X1 U757 ( .A1(n1049), .A2(KEYINPUT41), .A3(n1050), .ZN(n1048) );
INV_X1 U758 ( .A(n1051), .ZN(n1049) );
NAND2_X1 U759 ( .A1(n1050), .A2(n1052), .ZN(n1047) );
NAND2_X1 U760 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
NAND2_X1 U761 ( .A1(n1051), .A2(n1055), .ZN(n1054) );
OR2_X1 U762 ( .A1(KEYINPUT41), .A2(KEYINPUT5), .ZN(n1055) );
OR2_X1 U763 ( .A1(n1051), .A2(KEYINPUT5), .ZN(n1053) );
XNOR2_X1 U764 ( .A(n1056), .B(n1057), .ZN(n1051) );
XNOR2_X1 U765 ( .A(G137), .B(n1058), .ZN(n1057) );
XOR2_X1 U766 ( .A(n1059), .B(n1060), .Z(n1056) );
NOR2_X1 U767 ( .A1(G131), .A2(KEYINPUT51), .ZN(n1060) );
XOR2_X1 U768 ( .A(n1061), .B(KEYINPUT22), .Z(n1050) );
NAND3_X1 U769 ( .A1(G953), .A2(n1062), .A3(KEYINPUT10), .ZN(n1038) );
NAND2_X1 U770 ( .A1(G900), .A2(G227), .ZN(n1062) );
NAND2_X1 U771 ( .A1(n1063), .A2(n1064), .ZN(G69) );
NAND2_X1 U772 ( .A1(G953), .A2(n1065), .ZN(n1064) );
NAND2_X1 U773 ( .A1(G898), .A2(n1066), .ZN(n1065) );
NAND2_X1 U774 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
XOR2_X1 U775 ( .A(n1069), .B(KEYINPUT60), .Z(n1063) );
NAND2_X1 U776 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
NAND2_X1 U777 ( .A1(G953), .A2(n1068), .ZN(n1071) );
XOR2_X1 U778 ( .A(n1072), .B(n1067), .Z(n1070) );
XOR2_X1 U779 ( .A(n1073), .B(n1074), .Z(n1067) );
NAND3_X1 U780 ( .A1(n1075), .A2(n1042), .A3(KEYINPUT0), .ZN(n1072) );
NAND2_X1 U781 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
NOR2_X1 U782 ( .A1(n1078), .A2(n1079), .ZN(G66) );
XOR2_X1 U783 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U784 ( .A1(n1033), .A2(n1082), .ZN(n1080) );
NOR2_X1 U785 ( .A1(n1083), .A2(n1084), .ZN(G63) );
XNOR2_X1 U786 ( .A(n1078), .B(KEYINPUT33), .ZN(n1084) );
XOR2_X1 U787 ( .A(n1085), .B(n1086), .Z(n1083) );
NAND3_X1 U788 ( .A1(n1087), .A2(n1088), .A3(G478), .ZN(n1085) );
NAND2_X1 U789 ( .A1(KEYINPUT54), .A2(n1082), .ZN(n1088) );
NAND2_X1 U790 ( .A1(n1089), .A2(n1090), .ZN(n1087) );
INV_X1 U791 ( .A(KEYINPUT54), .ZN(n1090) );
OR2_X1 U792 ( .A1(n988), .A2(n1091), .ZN(n1089) );
NOR2_X1 U793 ( .A1(n1078), .A2(n1092), .ZN(G60) );
XOR2_X1 U794 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U795 ( .A(KEYINPUT24), .B(n1095), .ZN(n1094) );
AND2_X1 U796 ( .A1(G475), .A2(n1096), .ZN(n1093) );
XNOR2_X1 U797 ( .A(n1097), .B(n1098), .ZN(G6) );
NOR2_X1 U798 ( .A1(KEYINPUT30), .A2(n1099), .ZN(n1097) );
XNOR2_X1 U799 ( .A(G104), .B(KEYINPUT28), .ZN(n1099) );
NOR2_X1 U800 ( .A1(n1078), .A2(n1100), .ZN(G57) );
XNOR2_X1 U801 ( .A(n1101), .B(n1102), .ZN(n1100) );
NAND2_X1 U802 ( .A1(KEYINPUT3), .A2(n1103), .ZN(n1101) );
NAND2_X1 U803 ( .A1(n1096), .A2(G472), .ZN(n1103) );
NOR2_X1 U804 ( .A1(n1078), .A2(n1104), .ZN(G54) );
XOR2_X1 U805 ( .A(n1105), .B(n1106), .Z(n1104) );
AND2_X1 U806 ( .A1(G469), .A2(n1096), .ZN(n1106) );
INV_X1 U807 ( .A(n1082), .ZN(n1096) );
NAND2_X1 U808 ( .A1(n1107), .A2(KEYINPUT38), .ZN(n1105) );
XOR2_X1 U809 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U810 ( .A1(KEYINPUT19), .A2(n1059), .ZN(n1109) );
NOR2_X1 U811 ( .A1(n1078), .A2(n1110), .ZN(G51) );
XOR2_X1 U812 ( .A(n1111), .B(n1112), .Z(n1110) );
XOR2_X1 U813 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U814 ( .A1(n1115), .A2(n1082), .ZN(n1114) );
NAND2_X1 U815 ( .A1(G902), .A2(n988), .ZN(n1082) );
NAND3_X1 U816 ( .A1(n1076), .A2(n1116), .A3(n1046), .ZN(n988) );
AND4_X1 U817 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1046) );
NOR4_X1 U818 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
NOR3_X1 U819 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1124) );
INV_X1 U820 ( .A(n1010), .ZN(n1127) );
XNOR2_X1 U821 ( .A(n1014), .B(KEYINPUT49), .ZN(n1126) );
NOR2_X1 U822 ( .A1(n1125), .A2(n1128), .ZN(n1123) );
NOR2_X1 U823 ( .A1(n1129), .A2(n1130), .ZN(n1119) );
XNOR2_X1 U824 ( .A(KEYINPUT55), .B(n1077), .ZN(n1116) );
AND4_X1 U825 ( .A1(n1098), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1076) );
NOR4_X1 U826 ( .A1(n982), .A2(n1134), .A3(n1135), .A4(n1136), .ZN(n1133) );
INV_X1 U827 ( .A(n1137), .ZN(n1135) );
AND3_X1 U828 ( .A1(n1013), .A2(n1138), .A3(n1139), .ZN(n982) );
NAND3_X1 U829 ( .A1(n1140), .A2(n1141), .A3(n1142), .ZN(n1132) );
NOR3_X1 U830 ( .A1(n993), .A2(n1143), .A3(n994), .ZN(n1142) );
INV_X1 U831 ( .A(n1128), .ZN(n1141) );
XNOR2_X1 U832 ( .A(n1005), .B(KEYINPUT4), .ZN(n1140) );
NAND3_X1 U833 ( .A1(n1139), .A2(n1138), .A3(n1014), .ZN(n1098) );
NAND2_X1 U834 ( .A1(KEYINPUT6), .A2(n1144), .ZN(n1113) );
NOR2_X1 U835 ( .A1(n1042), .A2(G952), .ZN(n1078) );
XNOR2_X1 U836 ( .A(n1145), .B(n1122), .ZN(G48) );
AND3_X1 U837 ( .A1(n1014), .A2(n1005), .A3(n1146), .ZN(n1122) );
XOR2_X1 U838 ( .A(G143), .B(n1121), .Z(G45) );
AND3_X1 U839 ( .A1(n1011), .A2(n1147), .A3(n1148), .ZN(n1121) );
NOR3_X1 U840 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
XOR2_X1 U841 ( .A(n1152), .B(n1153), .Z(G42) );
NOR2_X1 U842 ( .A1(KEYINPUT13), .A2(n1154), .ZN(n1153) );
NOR2_X1 U843 ( .A1(n1009), .A2(n1155), .ZN(n1152) );
XOR2_X1 U844 ( .A(KEYINPUT48), .B(n1156), .Z(n1155) );
AND3_X1 U845 ( .A1(n1147), .A2(n1010), .A3(n1014), .ZN(n1156) );
XNOR2_X1 U846 ( .A(G137), .B(n1117), .ZN(G39) );
NAND3_X1 U847 ( .A1(n1157), .A2(n1146), .A3(n1016), .ZN(n1117) );
XNOR2_X1 U848 ( .A(G134), .B(n1118), .ZN(G36) );
NAND3_X1 U849 ( .A1(n1158), .A2(n1013), .A3(n1011), .ZN(n1118) );
INV_X1 U850 ( .A(n1125), .ZN(n1158) );
NAND2_X1 U851 ( .A1(n1157), .A2(n1147), .ZN(n1125) );
INV_X1 U852 ( .A(n1009), .ZN(n1157) );
XOR2_X1 U853 ( .A(G131), .B(n1159), .Z(G33) );
NOR4_X1 U854 ( .A1(n1009), .A2(n1160), .A3(n1128), .A4(n1161), .ZN(n1159) );
XNOR2_X1 U855 ( .A(KEYINPUT40), .B(n1162), .ZN(n1161) );
NAND2_X1 U856 ( .A1(n993), .A2(n1163), .ZN(n1160) );
NAND2_X1 U857 ( .A1(n1164), .A2(n1165), .ZN(n1009) );
XOR2_X1 U858 ( .A(n1006), .B(KEYINPUT50), .Z(n1164) );
XOR2_X1 U859 ( .A(n1166), .B(KEYINPUT43), .Z(n1006) );
XNOR2_X1 U860 ( .A(n1167), .B(n1130), .ZN(G30) );
AND3_X1 U861 ( .A1(n1013), .A2(n1005), .A3(n1146), .ZN(n1130) );
AND3_X1 U862 ( .A1(n1168), .A2(n1169), .A3(n1147), .ZN(n1146) );
AND3_X1 U863 ( .A1(n1162), .A2(n1163), .A3(n993), .ZN(n1147) );
INV_X1 U864 ( .A(n1149), .ZN(n1005) );
XNOR2_X1 U865 ( .A(G101), .B(n1131), .ZN(G3) );
NAND3_X1 U866 ( .A1(n1011), .A2(n1139), .A3(n1016), .ZN(n1131) );
XNOR2_X1 U867 ( .A(n1129), .B(n1170), .ZN(G27) );
NAND2_X1 U868 ( .A1(KEYINPUT34), .A2(G125), .ZN(n1170) );
AND4_X1 U869 ( .A1(n1014), .A2(n1171), .A3(n1010), .A4(n1162), .ZN(n1129) );
NAND2_X1 U870 ( .A1(n990), .A2(n1172), .ZN(n1162) );
NAND4_X1 U871 ( .A1(G953), .A2(G902), .A3(n1173), .A4(n1043), .ZN(n1172) );
INV_X1 U872 ( .A(G900), .ZN(n1043) );
XNOR2_X1 U873 ( .A(n1174), .B(n1136), .ZN(G24) );
NOR4_X1 U874 ( .A1(n1175), .A2(n1003), .A3(n1151), .A4(n1150), .ZN(n1136) );
INV_X1 U875 ( .A(n1138), .ZN(n1003) );
NOR2_X1 U876 ( .A1(n1169), .A2(n1168), .ZN(n1138) );
NAND2_X1 U877 ( .A1(n1176), .A2(n1177), .ZN(G21) );
OR2_X1 U878 ( .A1(n1137), .A2(G119), .ZN(n1177) );
XOR2_X1 U879 ( .A(n1178), .B(KEYINPUT16), .Z(n1176) );
NAND2_X1 U880 ( .A1(G119), .A2(n1137), .ZN(n1178) );
NAND4_X1 U881 ( .A1(n1179), .A2(n1016), .A3(n1168), .A4(n1169), .ZN(n1137) );
XNOR2_X1 U882 ( .A(n1134), .B(n1180), .ZN(G18) );
XOR2_X1 U883 ( .A(KEYINPUT39), .B(G116), .Z(n1180) );
AND3_X1 U884 ( .A1(n1011), .A2(n1013), .A3(n1179), .ZN(n1134) );
INV_X1 U885 ( .A(n1175), .ZN(n1179) );
NOR2_X1 U886 ( .A1(n1037), .A2(n1150), .ZN(n1013) );
INV_X1 U887 ( .A(n1181), .ZN(n1150) );
XOR2_X1 U888 ( .A(G113), .B(n1182), .Z(G15) );
NOR2_X1 U889 ( .A1(n1128), .A2(n1175), .ZN(n1182) );
NAND2_X1 U890 ( .A1(n1171), .A2(n1183), .ZN(n1175) );
NOR3_X1 U891 ( .A1(n1149), .A2(n994), .A3(n993), .ZN(n1171) );
NAND2_X1 U892 ( .A1(n1011), .A2(n1014), .ZN(n1128) );
NOR2_X1 U893 ( .A1(n1181), .A2(n1151), .ZN(n1014) );
INV_X1 U894 ( .A(n1037), .ZN(n1151) );
AND2_X1 U895 ( .A1(n1184), .A2(n1168), .ZN(n1011) );
XNOR2_X1 U896 ( .A(G110), .B(n1077), .ZN(G12) );
NAND3_X1 U897 ( .A1(n1010), .A2(n1139), .A3(n1016), .ZN(n1077) );
NOR2_X1 U898 ( .A1(n1181), .A2(n1037), .ZN(n1016) );
XNOR2_X1 U899 ( .A(n1185), .B(G475), .ZN(n1037) );
NAND2_X1 U900 ( .A1(n1091), .A2(n1095), .ZN(n1185) );
NAND2_X1 U901 ( .A1(n1186), .A2(n1187), .ZN(n1095) );
NAND2_X1 U902 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
XOR2_X1 U903 ( .A(KEYINPUT62), .B(n1190), .Z(n1189) );
XOR2_X1 U904 ( .A(KEYINPUT31), .B(n1191), .Z(n1188) );
XOR2_X1 U905 ( .A(KEYINPUT44), .B(n1192), .Z(n1186) );
NOR2_X1 U906 ( .A1(n1190), .A2(n1191), .ZN(n1192) );
XNOR2_X1 U907 ( .A(n1193), .B(G104), .ZN(n1191) );
NAND2_X1 U908 ( .A1(KEYINPUT2), .A2(n1194), .ZN(n1193) );
XNOR2_X1 U909 ( .A(n1174), .B(G113), .ZN(n1194) );
XNOR2_X1 U910 ( .A(n1195), .B(n1196), .ZN(n1190) );
XNOR2_X1 U911 ( .A(n1197), .B(n1198), .ZN(n1196) );
NOR3_X1 U912 ( .A1(n1199), .A2(KEYINPUT17), .A3(n1200), .ZN(n1198) );
INV_X1 U913 ( .A(G214), .ZN(n1200) );
NAND2_X1 U914 ( .A1(n1201), .A2(KEYINPUT46), .ZN(n1197) );
XNOR2_X1 U915 ( .A(G146), .B(n1061), .ZN(n1201) );
XNOR2_X1 U916 ( .A(G131), .B(G143), .ZN(n1195) );
NAND3_X1 U917 ( .A1(n1202), .A2(n1203), .A3(n1024), .ZN(n1181) );
NAND2_X1 U918 ( .A1(n1204), .A2(n1205), .ZN(n1024) );
OR2_X1 U919 ( .A1(G478), .A2(KEYINPUT42), .ZN(n1203) );
NAND2_X1 U920 ( .A1(n1022), .A2(KEYINPUT42), .ZN(n1202) );
NOR2_X1 U921 ( .A1(n1205), .A2(n1204), .ZN(n1022) );
AND2_X1 U922 ( .A1(n1086), .A2(n1091), .ZN(n1204) );
AND3_X1 U923 ( .A1(n1206), .A2(n1207), .A3(n1208), .ZN(n1086) );
NAND2_X1 U924 ( .A1(KEYINPUT1), .A2(n1209), .ZN(n1208) );
NAND2_X1 U925 ( .A1(G217), .A2(n1210), .ZN(n1209) );
NAND2_X1 U926 ( .A1(n1211), .A2(n1212), .ZN(n1207) );
INV_X1 U927 ( .A(n1213), .ZN(n1212) );
AND4_X1 U928 ( .A1(n1214), .A2(n1210), .A3(G217), .A4(KEYINPUT25), .ZN(n1211) );
INV_X1 U929 ( .A(KEYINPUT1), .ZN(n1214) );
NAND2_X1 U930 ( .A1(n1213), .A2(n1215), .ZN(n1206) );
NAND3_X1 U931 ( .A1(G217), .A2(n1210), .A3(KEYINPUT25), .ZN(n1215) );
XNOR2_X1 U932 ( .A(n1216), .B(n1217), .ZN(n1213) );
XNOR2_X1 U933 ( .A(n1058), .B(G128), .ZN(n1217) );
INV_X1 U934 ( .A(G134), .ZN(n1058) );
XNOR2_X1 U935 ( .A(n1218), .B(n1219), .ZN(n1216) );
NAND2_X1 U936 ( .A1(KEYINPUT12), .A2(G143), .ZN(n1219) );
NAND2_X1 U937 ( .A1(n1220), .A2(KEYINPUT20), .ZN(n1218) );
XNOR2_X1 U938 ( .A(G107), .B(n1221), .ZN(n1220) );
XNOR2_X1 U939 ( .A(n1174), .B(G116), .ZN(n1221) );
INV_X1 U940 ( .A(G122), .ZN(n1174) );
INV_X1 U941 ( .A(G478), .ZN(n1205) );
NOR4_X1 U942 ( .A1(n1149), .A2(n1222), .A3(n994), .A4(n1143), .ZN(n1139) );
INV_X1 U943 ( .A(n1183), .ZN(n1143) );
NAND2_X1 U944 ( .A1(n1223), .A2(n990), .ZN(n1183) );
NAND3_X1 U945 ( .A1(n1173), .A2(n1042), .A3(G952), .ZN(n990) );
XOR2_X1 U946 ( .A(KEYINPUT37), .B(n1224), .Z(n1223) );
NOR4_X1 U947 ( .A1(G898), .A2(n1225), .A3(n1091), .A4(n1042), .ZN(n1224) );
INV_X1 U948 ( .A(n1173), .ZN(n1225) );
NAND2_X1 U949 ( .A1(G234), .A2(G237), .ZN(n1173) );
INV_X1 U950 ( .A(n1163), .ZN(n994) );
NAND2_X1 U951 ( .A1(G221), .A2(n1226), .ZN(n1163) );
INV_X1 U952 ( .A(n993), .ZN(n1222) );
XNOR2_X1 U953 ( .A(n1227), .B(G469), .ZN(n993) );
NAND2_X1 U954 ( .A1(n1228), .A2(n1091), .ZN(n1227) );
XOR2_X1 U955 ( .A(n1059), .B(n1229), .Z(n1228) );
XOR2_X1 U956 ( .A(n1108), .B(KEYINPUT57), .Z(n1229) );
XOR2_X1 U957 ( .A(n1230), .B(n1231), .Z(n1108) );
XOR2_X1 U958 ( .A(n1232), .B(n1233), .Z(n1231) );
XNOR2_X1 U959 ( .A(G101), .B(G140), .ZN(n1233) );
NAND2_X1 U960 ( .A1(n1234), .A2(KEYINPUT45), .ZN(n1232) );
XNOR2_X1 U961 ( .A(G104), .B(n1235), .ZN(n1234) );
NOR2_X1 U962 ( .A1(G107), .A2(KEYINPUT18), .ZN(n1235) );
XOR2_X1 U963 ( .A(n1236), .B(n1237), .Z(n1230) );
XOR2_X1 U964 ( .A(n1238), .B(n1239), .Z(n1236) );
AND2_X1 U965 ( .A1(n1042), .A2(G227), .ZN(n1239) );
XNOR2_X1 U966 ( .A(G146), .B(n1240), .ZN(n1059) );
NAND2_X1 U967 ( .A1(n1166), .A2(n1165), .ZN(n1149) );
XNOR2_X1 U968 ( .A(n1007), .B(KEYINPUT47), .ZN(n1165) );
NAND2_X1 U969 ( .A1(G214), .A2(n1241), .ZN(n1007) );
XOR2_X1 U970 ( .A(n1028), .B(n1242), .Z(n1166) );
NOR2_X1 U971 ( .A1(n1243), .A2(n1244), .ZN(n1242) );
XNOR2_X1 U972 ( .A(KEYINPUT8), .B(KEYINPUT14), .ZN(n1244) );
XNOR2_X1 U973 ( .A(n1027), .B(KEYINPUT9), .ZN(n1243) );
INV_X1 U974 ( .A(n1115), .ZN(n1027) );
NAND2_X1 U975 ( .A1(G210), .A2(n1241), .ZN(n1115) );
NAND2_X1 U976 ( .A1(n1245), .A2(n1091), .ZN(n1241) );
XOR2_X1 U977 ( .A(KEYINPUT58), .B(G237), .Z(n1245) );
NAND2_X1 U978 ( .A1(n1246), .A2(n1091), .ZN(n1028) );
XOR2_X1 U979 ( .A(n1111), .B(n1247), .Z(n1246) );
XNOR2_X1 U980 ( .A(n1144), .B(KEYINPUT56), .ZN(n1247) );
XNOR2_X1 U981 ( .A(n1248), .B(n1249), .ZN(n1144) );
XOR2_X1 U982 ( .A(G125), .B(n1250), .Z(n1249) );
NOR2_X1 U983 ( .A1(G953), .A2(n1068), .ZN(n1250) );
INV_X1 U984 ( .A(G224), .ZN(n1068) );
XNOR2_X1 U985 ( .A(n1074), .B(n1251), .ZN(n1111) );
NOR2_X1 U986 ( .A1(KEYINPUT21), .A2(n1073), .ZN(n1251) );
XOR2_X1 U987 ( .A(n1252), .B(n1253), .Z(n1073) );
XOR2_X1 U988 ( .A(KEYINPUT53), .B(G107), .Z(n1253) );
XNOR2_X1 U989 ( .A(n1254), .B(n1255), .ZN(n1252) );
INV_X1 U990 ( .A(G104), .ZN(n1255) );
XOR2_X1 U991 ( .A(G122), .B(n1237), .Z(n1074) );
NOR2_X1 U992 ( .A1(n1168), .A2(n1184), .ZN(n1010) );
INV_X1 U993 ( .A(n1169), .ZN(n1184) );
NAND3_X1 U994 ( .A1(n1256), .A2(n1257), .A3(n1026), .ZN(n1169) );
NAND2_X1 U995 ( .A1(n1032), .A2(n1033), .ZN(n1026) );
NAND2_X1 U996 ( .A1(n1033), .A2(n1258), .ZN(n1257) );
OR3_X1 U997 ( .A1(n1033), .A2(n1032), .A3(n1258), .ZN(n1256) );
INV_X1 U998 ( .A(KEYINPUT23), .ZN(n1258) );
NOR2_X1 U999 ( .A1(n1081), .A2(G902), .ZN(n1032) );
XNOR2_X1 U1000 ( .A(n1259), .B(n1260), .ZN(n1081) );
XNOR2_X1 U1001 ( .A(n1061), .B(n1261), .ZN(n1260) );
XNOR2_X1 U1002 ( .A(n1237), .B(n1262), .ZN(n1261) );
XOR2_X1 U1003 ( .A(G110), .B(KEYINPUT52), .Z(n1237) );
XNOR2_X1 U1004 ( .A(G125), .B(n1154), .ZN(n1061) );
INV_X1 U1005 ( .A(G140), .ZN(n1154) );
XOR2_X1 U1006 ( .A(n1263), .B(n1264), .Z(n1259) );
XOR2_X1 U1007 ( .A(n1265), .B(n1266), .Z(n1264) );
NAND2_X1 U1008 ( .A1(KEYINPUT35), .A2(n1167), .ZN(n1266) );
NAND2_X1 U1009 ( .A1(KEYINPUT59), .A2(n1145), .ZN(n1265) );
XOR2_X1 U1010 ( .A(n1267), .B(G137), .Z(n1263) );
NAND2_X1 U1011 ( .A1(n1210), .A2(G221), .ZN(n1267) );
AND2_X1 U1012 ( .A1(G234), .A2(n1042), .ZN(n1210) );
INV_X1 U1013 ( .A(G953), .ZN(n1042) );
NAND2_X1 U1014 ( .A1(G217), .A2(n1226), .ZN(n1033) );
NAND2_X1 U1015 ( .A1(G234), .A2(n1091), .ZN(n1226) );
XNOR2_X1 U1016 ( .A(n1035), .B(G472), .ZN(n1168) );
NAND2_X1 U1017 ( .A1(n1102), .A2(n1091), .ZN(n1035) );
INV_X1 U1018 ( .A(G902), .ZN(n1091) );
XNOR2_X1 U1019 ( .A(n1268), .B(n1269), .ZN(n1102) );
XOR2_X1 U1020 ( .A(n1238), .B(n1248), .Z(n1269) );
NAND2_X1 U1021 ( .A1(n1270), .A2(n1271), .ZN(n1248) );
NAND2_X1 U1022 ( .A1(n1272), .A2(n1145), .ZN(n1271) );
INV_X1 U1023 ( .A(G146), .ZN(n1145) );
XOR2_X1 U1024 ( .A(KEYINPUT7), .B(n1240), .Z(n1272) );
NAND2_X1 U1025 ( .A1(n1240), .A2(G146), .ZN(n1270) );
XNOR2_X1 U1026 ( .A(n1167), .B(G143), .ZN(n1240) );
INV_X1 U1027 ( .A(G128), .ZN(n1167) );
XOR2_X1 U1028 ( .A(n1273), .B(G131), .Z(n1238) );
NAND2_X1 U1029 ( .A1(n1274), .A2(KEYINPUT11), .ZN(n1273) );
XNOR2_X1 U1030 ( .A(G134), .B(n1275), .ZN(n1274) );
NOR2_X1 U1031 ( .A1(G137), .A2(KEYINPUT61), .ZN(n1275) );
XOR2_X1 U1032 ( .A(n1254), .B(n1276), .Z(n1268) );
NOR2_X1 U1033 ( .A1(n1277), .A2(n1199), .ZN(n1276) );
OR2_X1 U1034 ( .A1(G953), .A2(G237), .ZN(n1199) );
INV_X1 U1035 ( .A(G210), .ZN(n1277) );
XOR2_X1 U1036 ( .A(n1278), .B(n1279), .Z(n1254) );
XOR2_X1 U1037 ( .A(G116), .B(G113), .Z(n1279) );
XNOR2_X1 U1038 ( .A(G101), .B(n1262), .ZN(n1278) );
XOR2_X1 U1039 ( .A(G119), .B(KEYINPUT27), .Z(n1262) );
endmodule


