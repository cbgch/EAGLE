//Key = 0011110001101110111011001011000010111010101100100000001100101000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355;

XNOR2_X1 U744 ( .A(n1030), .B(n1031), .ZN(G9) );
NOR2_X1 U745 ( .A1(n1032), .A2(n1033), .ZN(G75) );
NOR4_X1 U746 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1033) );
XOR2_X1 U747 ( .A(KEYINPUT20), .B(n1038), .Z(n1035) );
NOR2_X1 U748 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NOR2_X1 U749 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NOR2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
XOR2_X1 U751 ( .A(KEYINPUT62), .B(n1045), .Z(n1044) );
NOR3_X1 U752 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1045) );
NOR3_X1 U753 ( .A1(n1049), .A2(n1050), .A3(n1051), .ZN(n1043) );
NOR2_X1 U754 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
AND2_X1 U755 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
AND2_X1 U756 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
NOR3_X1 U757 ( .A1(n1058), .A2(n1059), .A3(n1060), .ZN(n1039) );
NAND4_X1 U758 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n1034) );
NAND3_X1 U759 ( .A1(n1065), .A2(n1066), .A3(n1067), .ZN(n1062) );
NAND2_X1 U760 ( .A1(n1068), .A2(n1069), .ZN(n1066) );
NAND3_X1 U761 ( .A1(n1070), .A2(n1054), .A3(n1071), .ZN(n1069) );
NAND2_X1 U762 ( .A1(n1056), .A2(n1072), .ZN(n1068) );
NAND2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U764 ( .A1(n1054), .A2(n1075), .ZN(n1074) );
NAND2_X1 U765 ( .A1(n1076), .A2(n1070), .ZN(n1073) );
NAND2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1061) );
XNOR2_X1 U767 ( .A(KEYINPUT1), .B(n1060), .ZN(n1078) );
OR2_X1 U768 ( .A1(n1047), .A2(n1051), .ZN(n1060) );
INV_X1 U769 ( .A(n1070), .ZN(n1051) );
NAND3_X1 U770 ( .A1(n1054), .A2(n1056), .A3(n1067), .ZN(n1047) );
INV_X1 U771 ( .A(n1049), .ZN(n1067) );
NOR3_X1 U772 ( .A1(n1079), .A2(G953), .A3(G952), .ZN(n1032) );
INV_X1 U773 ( .A(n1063), .ZN(n1079) );
NAND4_X1 U774 ( .A1(n1080), .A2(n1065), .A3(n1081), .A4(n1082), .ZN(n1063) );
NOR4_X1 U775 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
XNOR2_X1 U776 ( .A(n1048), .B(KEYINPUT10), .ZN(n1086) );
XOR2_X1 U777 ( .A(n1087), .B(KEYINPUT50), .Z(n1085) );
NAND3_X1 U778 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1087) );
OR2_X1 U779 ( .A1(G475), .A2(KEYINPUT26), .ZN(n1089) );
NAND3_X1 U780 ( .A1(G475), .A2(n1091), .A3(KEYINPUT26), .ZN(n1088) );
XOR2_X1 U781 ( .A(n1092), .B(G472), .Z(n1084) );
NAND2_X1 U782 ( .A1(KEYINPUT35), .A2(n1093), .ZN(n1092) );
XOR2_X1 U783 ( .A(n1094), .B(n1095), .Z(n1081) );
XOR2_X1 U784 ( .A(n1096), .B(n1097), .Z(G72) );
XOR2_X1 U785 ( .A(n1098), .B(n1099), .Z(n1097) );
NOR2_X1 U786 ( .A1(n1100), .A2(n1064), .ZN(n1099) );
AND2_X1 U787 ( .A1(G227), .A2(G900), .ZN(n1100) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1102), .ZN(n1098) );
NAND2_X1 U789 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
XOR2_X1 U790 ( .A(n1105), .B(n1106), .Z(n1101) );
XOR2_X1 U791 ( .A(n1107), .B(n1108), .Z(n1106) );
XOR2_X1 U792 ( .A(n1109), .B(n1110), .Z(n1107) );
NOR2_X1 U793 ( .A1(KEYINPUT52), .A2(n1111), .ZN(n1110) );
NOR2_X1 U794 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
XOR2_X1 U795 ( .A(n1114), .B(G131), .Z(n1105) );
XNOR2_X1 U796 ( .A(KEYINPUT63), .B(KEYINPUT47), .ZN(n1114) );
NAND2_X1 U797 ( .A1(n1064), .A2(n1036), .ZN(n1096) );
XOR2_X1 U798 ( .A(n1115), .B(n1116), .Z(G69) );
NAND2_X1 U799 ( .A1(G953), .A2(n1117), .ZN(n1116) );
NAND2_X1 U800 ( .A1(G898), .A2(G224), .ZN(n1117) );
NAND2_X1 U801 ( .A1(KEYINPUT43), .A2(n1118), .ZN(n1115) );
XOR2_X1 U802 ( .A(n1119), .B(n1120), .Z(n1118) );
NOR3_X1 U803 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(n1120) );
NOR2_X1 U804 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U805 ( .A(KEYINPUT3), .B(n1126), .Z(n1124) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1126), .ZN(n1122) );
XNOR2_X1 U807 ( .A(n1128), .B(n1129), .ZN(n1126) );
NAND2_X1 U808 ( .A1(KEYINPUT18), .A2(n1130), .ZN(n1128) );
XOR2_X1 U809 ( .A(n1131), .B(n1132), .Z(n1130) );
NOR3_X1 U810 ( .A1(n1133), .A2(KEYINPUT41), .A3(G953), .ZN(n1119) );
INV_X1 U811 ( .A(n1037), .ZN(n1133) );
NOR2_X1 U812 ( .A1(n1134), .A2(n1135), .ZN(G66) );
XOR2_X1 U813 ( .A(n1136), .B(n1137), .Z(n1135) );
NAND2_X1 U814 ( .A1(n1138), .A2(G217), .ZN(n1136) );
NOR2_X1 U815 ( .A1(n1134), .A2(n1139), .ZN(G63) );
XOR2_X1 U816 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U817 ( .A1(n1138), .A2(G478), .ZN(n1140) );
NOR2_X1 U818 ( .A1(n1134), .A2(n1142), .ZN(G60) );
NOR2_X1 U819 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
XOR2_X1 U820 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U821 ( .A1(n1138), .A2(G475), .ZN(n1146) );
NAND2_X1 U822 ( .A1(n1147), .A2(n1148), .ZN(n1145) );
NOR2_X1 U823 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
INV_X1 U824 ( .A(KEYINPUT48), .ZN(n1148) );
XOR2_X1 U825 ( .A(G104), .B(n1149), .Z(G6) );
NOR2_X1 U826 ( .A1(n1150), .A2(n1151), .ZN(G57) );
XOR2_X1 U827 ( .A(KEYINPUT19), .B(n1134), .Z(n1151) );
XOR2_X1 U828 ( .A(n1152), .B(n1153), .Z(n1150) );
XNOR2_X1 U829 ( .A(n1154), .B(n1155), .ZN(n1153) );
XOR2_X1 U830 ( .A(n1156), .B(n1131), .Z(n1155) );
NAND2_X1 U831 ( .A1(KEYINPUT14), .A2(n1157), .ZN(n1156) );
XOR2_X1 U832 ( .A(n1158), .B(n1159), .Z(n1152) );
XOR2_X1 U833 ( .A(n1160), .B(KEYINPUT61), .Z(n1159) );
NAND2_X1 U834 ( .A1(n1138), .A2(G472), .ZN(n1160) );
NAND2_X1 U835 ( .A1(KEYINPUT13), .A2(n1161), .ZN(n1158) );
NOR2_X1 U836 ( .A1(n1134), .A2(n1162), .ZN(G54) );
XOR2_X1 U837 ( .A(n1163), .B(n1164), .Z(n1162) );
XOR2_X1 U838 ( .A(n1165), .B(n1166), .Z(n1164) );
NAND2_X1 U839 ( .A1(n1138), .A2(G469), .ZN(n1165) );
XOR2_X1 U840 ( .A(n1167), .B(n1168), .Z(n1163) );
XOR2_X1 U841 ( .A(KEYINPUT5), .B(KEYINPUT17), .Z(n1168) );
NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n1169), .ZN(n1167) );
XOR2_X1 U843 ( .A(n1170), .B(n1171), .Z(n1169) );
XNOR2_X1 U844 ( .A(n1172), .B(n1108), .ZN(n1171) );
XOR2_X1 U845 ( .A(n1173), .B(KEYINPUT8), .Z(n1170) );
NAND2_X1 U846 ( .A1(KEYINPUT54), .A2(n1174), .ZN(n1173) );
INV_X1 U847 ( .A(n1129), .ZN(n1174) );
NOR2_X1 U848 ( .A1(n1134), .A2(n1175), .ZN(G51) );
XOR2_X1 U849 ( .A(n1176), .B(n1177), .Z(n1175) );
XOR2_X1 U850 ( .A(n1178), .B(KEYINPUT59), .Z(n1177) );
NAND2_X1 U851 ( .A1(n1138), .A2(G210), .ZN(n1178) );
AND2_X1 U852 ( .A1(G902), .A2(n1179), .ZN(n1138) );
OR2_X1 U853 ( .A1(n1037), .A2(n1036), .ZN(n1179) );
NAND4_X1 U854 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1036) );
NOR3_X1 U855 ( .A1(n1184), .A2(n1185), .A3(n1186), .ZN(n1183) );
NAND3_X1 U856 ( .A1(n1076), .A2(n1187), .A3(n1188), .ZN(n1182) );
NAND2_X1 U857 ( .A1(n1189), .A2(n1190), .ZN(n1187) );
NAND2_X1 U858 ( .A1(n1065), .A2(n1055), .ZN(n1190) );
NAND2_X1 U859 ( .A1(n1191), .A2(n1077), .ZN(n1189) );
NAND4_X1 U860 ( .A1(n1057), .A2(n1071), .A3(n1192), .A4(n1193), .ZN(n1180) );
NAND2_X1 U861 ( .A1(n1194), .A2(n1195), .ZN(n1192) );
NAND2_X1 U862 ( .A1(n1065), .A2(n1196), .ZN(n1195) );
XOR2_X1 U863 ( .A(KEYINPUT22), .B(n1075), .Z(n1196) );
NAND2_X1 U864 ( .A1(n1197), .A2(n1070), .ZN(n1194) );
XNOR2_X1 U865 ( .A(n1077), .B(KEYINPUT60), .ZN(n1197) );
NAND4_X1 U866 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1037) );
NOR4_X1 U867 ( .A1(n1031), .A2(n1149), .A3(n1202), .A4(n1203), .ZN(n1201) );
INV_X1 U868 ( .A(n1204), .ZN(n1202) );
AND3_X1 U869 ( .A1(n1054), .A2(n1205), .A3(n1071), .ZN(n1149) );
AND3_X1 U870 ( .A1(n1054), .A2(n1205), .A3(n1055), .ZN(n1031) );
NOR2_X1 U871 ( .A1(n1206), .A2(n1207), .ZN(n1200) );
NOR3_X1 U872 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1207) );
NOR2_X1 U873 ( .A1(n1064), .A2(G952), .ZN(n1134) );
XNOR2_X1 U874 ( .A(G146), .B(n1181), .ZN(G48) );
NAND3_X1 U875 ( .A1(n1071), .A2(n1077), .A3(n1211), .ZN(n1181) );
XNOR2_X1 U876 ( .A(n1212), .B(n1213), .ZN(G45) );
NOR2_X1 U877 ( .A1(n1214), .A2(n1215), .ZN(n1213) );
XOR2_X1 U878 ( .A(KEYINPUT32), .B(n1216), .Z(n1215) );
NOR3_X1 U879 ( .A1(n1217), .A2(n1208), .A3(n1218), .ZN(n1216) );
XOR2_X1 U880 ( .A(KEYINPUT21), .B(n1191), .Z(n1217) );
XNOR2_X1 U881 ( .A(G140), .B(n1219), .ZN(G42) );
NAND4_X1 U882 ( .A1(n1188), .A2(n1057), .A3(n1220), .A4(n1071), .ZN(n1219) );
NOR2_X1 U883 ( .A1(KEYINPUT11), .A2(n1042), .ZN(n1220) );
XOR2_X1 U884 ( .A(G137), .B(n1184), .Z(G39) );
AND3_X1 U885 ( .A1(n1065), .A2(n1056), .A3(n1211), .ZN(n1184) );
XNOR2_X1 U886 ( .A(G134), .B(n1221), .ZN(G36) );
NAND3_X1 U887 ( .A1(n1222), .A2(n1055), .A3(KEYINPUT2), .ZN(n1221) );
XOR2_X1 U888 ( .A(G131), .B(n1186), .Z(G33) );
AND2_X1 U889 ( .A1(n1222), .A2(n1071), .ZN(n1186) );
NOR3_X1 U890 ( .A1(n1208), .A2(n1042), .A3(n1218), .ZN(n1222) );
INV_X1 U891 ( .A(n1065), .ZN(n1042) );
NOR2_X1 U892 ( .A1(n1059), .A2(n1223), .ZN(n1065) );
INV_X1 U893 ( .A(n1058), .ZN(n1223) );
XNOR2_X1 U894 ( .A(n1224), .B(n1185), .ZN(G30) );
AND3_X1 U895 ( .A1(n1055), .A2(n1077), .A3(n1211), .ZN(n1185) );
AND3_X1 U896 ( .A1(n1225), .A2(n1226), .A3(n1188), .ZN(n1211) );
INV_X1 U897 ( .A(n1218), .ZN(n1188) );
NAND2_X1 U898 ( .A1(n1075), .A2(n1193), .ZN(n1218) );
INV_X1 U899 ( .A(n1227), .ZN(n1055) );
XNOR2_X1 U900 ( .A(n1228), .B(n1206), .ZN(G3) );
AND3_X1 U901 ( .A1(n1205), .A2(n1056), .A3(n1076), .ZN(n1206) );
XNOR2_X1 U902 ( .A(n1229), .B(n1230), .ZN(G27) );
NOR4_X1 U903 ( .A1(n1231), .A2(n1214), .A3(KEYINPUT7), .A4(n1232), .ZN(n1230) );
INV_X1 U904 ( .A(n1193), .ZN(n1232) );
NAND2_X1 U905 ( .A1(n1049), .A2(n1233), .ZN(n1193) );
NAND4_X1 U906 ( .A1(n1103), .A2(G902), .A3(n1234), .A4(n1104), .ZN(n1233) );
INV_X1 U907 ( .A(G900), .ZN(n1104) );
INV_X1 U908 ( .A(n1235), .ZN(n1103) );
NAND3_X1 U909 ( .A1(n1071), .A2(n1070), .A3(n1057), .ZN(n1231) );
XNOR2_X1 U910 ( .A(G122), .B(n1198), .ZN(G24) );
NAND3_X1 U911 ( .A1(n1236), .A2(n1054), .A3(n1191), .ZN(n1198) );
AND2_X1 U912 ( .A1(n1237), .A2(n1238), .ZN(n1191) );
XNOR2_X1 U913 ( .A(KEYINPUT42), .B(n1239), .ZN(n1237) );
NOR2_X1 U914 ( .A1(n1226), .A2(n1240), .ZN(n1054) );
XNOR2_X1 U915 ( .A(G119), .B(n1199), .ZN(G21) );
NAND4_X1 U916 ( .A1(n1225), .A2(n1236), .A3(n1056), .A4(n1226), .ZN(n1199) );
INV_X1 U917 ( .A(n1210), .ZN(n1236) );
NAND2_X1 U918 ( .A1(n1241), .A2(n1242), .ZN(G18) );
NAND2_X1 U919 ( .A1(n1203), .A2(n1243), .ZN(n1242) );
XOR2_X1 U920 ( .A(n1244), .B(KEYINPUT53), .Z(n1241) );
OR2_X1 U921 ( .A1(n1243), .A2(n1203), .ZN(n1244) );
NOR3_X1 U922 ( .A1(n1210), .A2(n1227), .A3(n1208), .ZN(n1203) );
INV_X1 U923 ( .A(n1076), .ZN(n1208) );
NAND2_X1 U924 ( .A1(n1245), .A2(n1238), .ZN(n1227) );
XNOR2_X1 U925 ( .A(n1246), .B(KEYINPUT34), .ZN(n1245) );
NAND2_X1 U926 ( .A1(n1070), .A2(n1247), .ZN(n1210) );
XOR2_X1 U927 ( .A(n1248), .B(n1249), .Z(G15) );
NAND2_X1 U928 ( .A1(KEYINPUT55), .A2(G113), .ZN(n1249) );
NAND4_X1 U929 ( .A1(n1250), .A2(n1076), .A3(n1071), .A4(n1247), .ZN(n1248) );
NOR2_X1 U930 ( .A1(n1251), .A2(n1240), .ZN(n1076) );
INV_X1 U931 ( .A(n1252), .ZN(n1240) );
XNOR2_X1 U932 ( .A(n1070), .B(KEYINPUT16), .ZN(n1250) );
NOR2_X1 U933 ( .A1(n1048), .A2(n1083), .ZN(n1070) );
XOR2_X1 U934 ( .A(G110), .B(n1253), .Z(G12) );
NOR2_X1 U935 ( .A1(KEYINPUT31), .A2(n1204), .ZN(n1253) );
NAND3_X1 U936 ( .A1(n1205), .A2(n1056), .A3(n1057), .ZN(n1204) );
AND2_X1 U937 ( .A1(n1225), .A2(n1251), .ZN(n1057) );
INV_X1 U938 ( .A(n1226), .ZN(n1251) );
XNOR2_X1 U939 ( .A(n1093), .B(G472), .ZN(n1226) );
NAND2_X1 U940 ( .A1(n1254), .A2(n1255), .ZN(n1093) );
XNOR2_X1 U941 ( .A(n1256), .B(n1257), .ZN(n1254) );
INV_X1 U942 ( .A(n1154), .ZN(n1257) );
XOR2_X1 U943 ( .A(n1258), .B(n1259), .Z(n1154) );
INV_X1 U944 ( .A(n1172), .ZN(n1259) );
XNOR2_X1 U945 ( .A(n1260), .B(n1228), .ZN(n1258) );
INV_X1 U946 ( .A(G101), .ZN(n1228) );
NAND2_X1 U947 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
OR2_X1 U948 ( .A1(n1263), .A2(n1243), .ZN(n1262) );
XOR2_X1 U949 ( .A(n1264), .B(KEYINPUT37), .Z(n1261) );
NAND2_X1 U950 ( .A1(n1263), .A2(n1243), .ZN(n1264) );
INV_X1 U951 ( .A(G116), .ZN(n1243) );
XOR2_X1 U952 ( .A(G119), .B(KEYINPUT56), .Z(n1263) );
XNOR2_X1 U953 ( .A(n1157), .B(n1265), .ZN(n1256) );
AND3_X1 U954 ( .A1(n1266), .A2(n1064), .A3(G210), .ZN(n1157) );
XNOR2_X1 U955 ( .A(n1252), .B(KEYINPUT23), .ZN(n1225) );
XNOR2_X1 U956 ( .A(n1094), .B(n1267), .ZN(n1252) );
NOR2_X1 U957 ( .A1(n1095), .A2(KEYINPUT29), .ZN(n1267) );
AND2_X1 U958 ( .A1(n1137), .A2(n1255), .ZN(n1095) );
XOR2_X1 U959 ( .A(n1268), .B(n1269), .Z(n1137) );
XOR2_X1 U960 ( .A(n1270), .B(n1271), .Z(n1269) );
XOR2_X1 U961 ( .A(n1272), .B(n1273), .Z(n1271) );
NOR3_X1 U962 ( .A1(n1274), .A2(KEYINPUT15), .A3(n1275), .ZN(n1273) );
INV_X1 U963 ( .A(G221), .ZN(n1274) );
NOR3_X1 U964 ( .A1(n1113), .A2(n1276), .A3(n1277), .ZN(n1272) );
NOR2_X1 U965 ( .A1(n1229), .A2(n1278), .ZN(n1277) );
AND2_X1 U966 ( .A1(n1278), .A2(n1112), .ZN(n1276) );
INV_X1 U967 ( .A(KEYINPUT25), .ZN(n1278) );
INV_X1 U968 ( .A(n1279), .ZN(n1113) );
XNOR2_X1 U969 ( .A(n1280), .B(G110), .ZN(n1270) );
XOR2_X1 U970 ( .A(n1281), .B(n1282), .Z(n1268) );
XOR2_X1 U971 ( .A(KEYINPUT27), .B(G146), .Z(n1282) );
XNOR2_X1 U972 ( .A(G137), .B(G128), .ZN(n1281) );
NAND2_X1 U973 ( .A1(n1283), .A2(G217), .ZN(n1094) );
XOR2_X1 U974 ( .A(n1284), .B(KEYINPUT39), .Z(n1283) );
NAND2_X1 U975 ( .A1(n1285), .A2(n1286), .ZN(n1056) );
OR2_X1 U976 ( .A1(n1209), .A2(KEYINPUT34), .ZN(n1286) );
INV_X1 U977 ( .A(n1071), .ZN(n1209) );
NOR2_X1 U978 ( .A1(n1238), .A2(n1246), .ZN(n1071) );
NAND3_X1 U979 ( .A1(n1246), .A2(n1080), .A3(KEYINPUT34), .ZN(n1285) );
INV_X1 U980 ( .A(n1238), .ZN(n1080) );
XNOR2_X1 U981 ( .A(n1287), .B(G478), .ZN(n1238) );
NAND2_X1 U982 ( .A1(n1141), .A2(n1255), .ZN(n1287) );
XNOR2_X1 U983 ( .A(n1288), .B(n1289), .ZN(n1141) );
NOR2_X1 U984 ( .A1(n1275), .A2(n1290), .ZN(n1289) );
INV_X1 U985 ( .A(G217), .ZN(n1290) );
NAND2_X1 U986 ( .A1(G234), .A2(n1064), .ZN(n1275) );
NAND2_X1 U987 ( .A1(KEYINPUT58), .A2(n1291), .ZN(n1288) );
XOR2_X1 U988 ( .A(n1292), .B(n1293), .Z(n1291) );
XNOR2_X1 U989 ( .A(n1294), .B(n1295), .ZN(n1293) );
NAND3_X1 U990 ( .A1(n1296), .A2(n1297), .A3(n1298), .ZN(n1294) );
NAND2_X1 U991 ( .A1(KEYINPUT0), .A2(n1299), .ZN(n1298) );
NAND3_X1 U992 ( .A1(n1300), .A2(n1301), .A3(n1030), .ZN(n1297) );
INV_X1 U993 ( .A(KEYINPUT0), .ZN(n1301) );
OR2_X1 U994 ( .A1(n1030), .A2(n1300), .ZN(n1296) );
NOR2_X1 U995 ( .A1(KEYINPUT30), .A2(n1299), .ZN(n1300) );
XNOR2_X1 U996 ( .A(n1302), .B(G116), .ZN(n1299) );
NAND2_X1 U997 ( .A1(KEYINPUT40), .A2(n1303), .ZN(n1302) );
XNOR2_X1 U998 ( .A(n1212), .B(G128), .ZN(n1292) );
INV_X1 U999 ( .A(n1239), .ZN(n1246) );
NAND2_X1 U1000 ( .A1(n1090), .A2(n1304), .ZN(n1239) );
NAND2_X1 U1001 ( .A1(G475), .A2(n1091), .ZN(n1304) );
OR2_X1 U1002 ( .A1(n1091), .A2(G475), .ZN(n1090) );
NAND2_X1 U1003 ( .A1(n1147), .A2(n1255), .ZN(n1091) );
XNOR2_X1 U1004 ( .A(n1305), .B(n1306), .ZN(n1147) );
XNOR2_X1 U1005 ( .A(n1307), .B(n1308), .ZN(n1306) );
XOR2_X1 U1006 ( .A(n1309), .B(n1131), .Z(n1308) );
NAND3_X1 U1007 ( .A1(n1310), .A2(n1311), .A3(n1279), .ZN(n1309) );
NAND2_X1 U1008 ( .A1(G140), .A2(G125), .ZN(n1279) );
OR2_X1 U1009 ( .A1(n1229), .A2(KEYINPUT36), .ZN(n1311) );
NAND2_X1 U1010 ( .A1(n1112), .A2(KEYINPUT36), .ZN(n1310) );
NOR2_X1 U1011 ( .A1(G125), .A2(G140), .ZN(n1112) );
XOR2_X1 U1012 ( .A(n1312), .B(n1313), .Z(n1305) );
XNOR2_X1 U1013 ( .A(G131), .B(n1303), .ZN(n1313) );
XNOR2_X1 U1014 ( .A(G104), .B(n1314), .ZN(n1312) );
NOR2_X1 U1015 ( .A1(n1315), .A2(KEYINPUT6), .ZN(n1314) );
AND3_X1 U1016 ( .A1(G214), .A2(n1064), .A3(n1266), .ZN(n1315) );
AND2_X1 U1017 ( .A1(n1075), .A2(n1247), .ZN(n1205) );
AND2_X1 U1018 ( .A1(n1077), .A2(n1316), .ZN(n1247) );
NAND2_X1 U1019 ( .A1(n1049), .A2(n1317), .ZN(n1316) );
NAND3_X1 U1020 ( .A1(n1121), .A2(n1234), .A3(G902), .ZN(n1317) );
NOR2_X1 U1021 ( .A1(n1235), .A2(G898), .ZN(n1121) );
XOR2_X1 U1022 ( .A(G953), .B(KEYINPUT9), .Z(n1235) );
NAND3_X1 U1023 ( .A1(n1234), .A2(n1064), .A3(G952), .ZN(n1049) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1234) );
INV_X1 U1025 ( .A(n1214), .ZN(n1077) );
NAND2_X1 U1026 ( .A1(n1059), .A2(n1058), .ZN(n1214) );
NAND2_X1 U1027 ( .A1(G214), .A2(n1318), .ZN(n1058) );
NAND2_X1 U1028 ( .A1(n1266), .A2(n1255), .ZN(n1318) );
NAND2_X1 U1029 ( .A1(n1319), .A2(n1320), .ZN(n1059) );
NAND2_X1 U1030 ( .A1(G210), .A2(n1321), .ZN(n1320) );
NAND2_X1 U1031 ( .A1(n1255), .A2(n1322), .ZN(n1321) );
OR2_X1 U1032 ( .A1(n1266), .A2(n1323), .ZN(n1322) );
INV_X1 U1033 ( .A(G237), .ZN(n1266) );
NAND3_X1 U1034 ( .A1(n1324), .A2(n1255), .A3(n1323), .ZN(n1319) );
XOR2_X1 U1035 ( .A(n1176), .B(KEYINPUT28), .Z(n1323) );
XOR2_X1 U1036 ( .A(n1325), .B(n1326), .Z(n1176) );
XOR2_X1 U1037 ( .A(n1327), .B(n1328), .Z(n1326) );
XNOR2_X1 U1038 ( .A(n1229), .B(n1329), .ZN(n1328) );
NOR2_X1 U1039 ( .A1(n1127), .A2(KEYINPUT51), .ZN(n1329) );
INV_X1 U1040 ( .A(n1125), .ZN(n1127) );
NAND3_X1 U1041 ( .A1(n1330), .A2(n1331), .A3(n1332), .ZN(n1125) );
NAND2_X1 U1042 ( .A1(n1333), .A2(n1303), .ZN(n1332) );
OR3_X1 U1043 ( .A1(n1333), .A2(n1303), .A3(KEYINPUT57), .ZN(n1331) );
INV_X1 U1044 ( .A(G122), .ZN(n1303) );
NAND2_X1 U1045 ( .A1(KEYINPUT12), .A2(G110), .ZN(n1333) );
NAND2_X1 U1046 ( .A1(KEYINPUT57), .A2(n1334), .ZN(n1330) );
INV_X1 U1047 ( .A(G125), .ZN(n1229) );
AND2_X1 U1048 ( .A1(n1064), .A2(G224), .ZN(n1327) );
XOR2_X1 U1049 ( .A(n1335), .B(n1132), .Z(n1325) );
XNOR2_X1 U1050 ( .A(n1280), .B(G116), .ZN(n1132) );
INV_X1 U1051 ( .A(G119), .ZN(n1280) );
XNOR2_X1 U1052 ( .A(n1129), .B(n1265), .ZN(n1335) );
XOR2_X1 U1053 ( .A(n1131), .B(n1161), .Z(n1265) );
XNOR2_X1 U1054 ( .A(n1336), .B(G128), .ZN(n1161) );
NAND2_X1 U1055 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
NAND2_X1 U1056 ( .A1(n1339), .A2(n1340), .ZN(n1338) );
XNOR2_X1 U1057 ( .A(KEYINPUT44), .B(n1212), .ZN(n1340) );
INV_X1 U1058 ( .A(G143), .ZN(n1212) );
XNOR2_X1 U1059 ( .A(KEYINPUT49), .B(G146), .ZN(n1339) );
XOR2_X1 U1060 ( .A(n1341), .B(KEYINPUT45), .Z(n1337) );
NAND2_X1 U1061 ( .A1(n1342), .A2(n1343), .ZN(n1341) );
XOR2_X1 U1062 ( .A(KEYINPUT49), .B(G146), .Z(n1343) );
XNOR2_X1 U1063 ( .A(KEYINPUT44), .B(G143), .ZN(n1342) );
XOR2_X1 U1064 ( .A(G113), .B(KEYINPUT4), .Z(n1131) );
NAND2_X1 U1065 ( .A1(G237), .A2(G210), .ZN(n1324) );
NOR2_X1 U1066 ( .A1(n1344), .A2(n1083), .ZN(n1075) );
INV_X1 U1067 ( .A(n1046), .ZN(n1083) );
NAND2_X1 U1068 ( .A1(G221), .A2(n1284), .ZN(n1046) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1255), .ZN(n1284) );
INV_X1 U1070 ( .A(n1048), .ZN(n1344) );
XNOR2_X1 U1071 ( .A(n1345), .B(G469), .ZN(n1048) );
NAND2_X1 U1072 ( .A1(n1346), .A2(n1255), .ZN(n1345) );
INV_X1 U1073 ( .A(G902), .ZN(n1255) );
XOR2_X1 U1074 ( .A(n1347), .B(n1348), .Z(n1346) );
XNOR2_X1 U1075 ( .A(n1166), .B(n1108), .ZN(n1348) );
XOR2_X1 U1076 ( .A(n1349), .B(n1350), .Z(n1108) );
INV_X1 U1077 ( .A(n1307), .ZN(n1350) );
XOR2_X1 U1078 ( .A(G143), .B(G146), .Z(n1307) );
XOR2_X1 U1079 ( .A(n1351), .B(KEYINPUT44), .Z(n1349) );
NAND2_X1 U1080 ( .A1(KEYINPUT24), .A2(n1224), .ZN(n1351) );
INV_X1 U1081 ( .A(G128), .ZN(n1224) );
XOR2_X1 U1082 ( .A(n1352), .B(n1353), .Z(n1166) );
XNOR2_X1 U1083 ( .A(G140), .B(n1334), .ZN(n1353) );
INV_X1 U1084 ( .A(G110), .ZN(n1334) );
NAND2_X1 U1085 ( .A1(G227), .A2(n1064), .ZN(n1352) );
INV_X1 U1086 ( .A(G953), .ZN(n1064) );
XNOR2_X1 U1087 ( .A(n1172), .B(n1129), .ZN(n1347) );
XOR2_X1 U1088 ( .A(G101), .B(n1354), .Z(n1129) );
XNOR2_X1 U1089 ( .A(n1030), .B(G104), .ZN(n1354) );
INV_X1 U1090 ( .A(G107), .ZN(n1030) );
XNOR2_X1 U1091 ( .A(n1355), .B(G131), .ZN(n1172) );
NAND2_X1 U1092 ( .A1(KEYINPUT38), .A2(n1109), .ZN(n1355) );
XNOR2_X1 U1093 ( .A(G137), .B(n1295), .ZN(n1109) );
XOR2_X1 U1094 ( .A(G134), .B(KEYINPUT46), .Z(n1295) );
endmodule


