//Key = 0001010110100010010000000101000001001000011111101111100110111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356;

XOR2_X1 U735 ( .A(n1020), .B(n1021), .Z(G9) );
NOR2_X1 U736 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR3_X1 U737 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
INV_X1 U738 ( .A(KEYINPUT20), .ZN(n1024) );
NOR2_X1 U739 ( .A1(KEYINPUT20), .A2(n1027), .ZN(n1022) );
NOR2_X1 U740 ( .A1(n1028), .A2(n1029), .ZN(G75) );
NOR4_X1 U741 ( .A1(G953), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1029) );
NOR2_X1 U742 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR2_X1 U743 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NOR3_X1 U744 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
NOR3_X1 U745 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n1039) );
NOR2_X1 U746 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR2_X1 U747 ( .A1(n1045), .A2(n1046), .ZN(n1041) );
NOR2_X1 U748 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NOR2_X1 U749 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U750 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
XOR2_X1 U751 ( .A(KEYINPUT21), .B(n1053), .Z(n1052) );
NOR2_X1 U752 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR3_X1 U753 ( .A1(n1056), .A2(KEYINPUT14), .A3(n1043), .ZN(n1047) );
AND3_X1 U754 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1043) );
NAND2_X1 U755 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
NAND2_X1 U757 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
XOR2_X1 U758 ( .A(KEYINPUT45), .B(n1066), .Z(n1065) );
INV_X1 U759 ( .A(n1067), .ZN(n1064) );
NAND2_X1 U760 ( .A1(KEYINPUT14), .A2(n1068), .ZN(n1062) );
NAND2_X1 U761 ( .A1(n1069), .A2(n1070), .ZN(n1057) );
OR2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1038) );
AND2_X1 U764 ( .A1(n1075), .A2(n1073), .ZN(n1035) );
NOR3_X1 U765 ( .A1(n1044), .A2(n1050), .A3(n1046), .ZN(n1073) );
INV_X1 U766 ( .A(n1069), .ZN(n1050) );
NOR3_X1 U767 ( .A1(n1030), .A2(G953), .A3(G952), .ZN(n1028) );
AND4_X1 U768 ( .A1(n1076), .A2(n1067), .A3(n1077), .A4(n1078), .ZN(n1030) );
NOR4_X1 U769 ( .A1(n1079), .A2(n1044), .A3(n1080), .A4(n1066), .ZN(n1078) );
AND2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND3_X1 U771 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1079) );
XOR2_X1 U772 ( .A(n1086), .B(G472), .Z(n1085) );
OR2_X1 U773 ( .A1(G478), .A2(KEYINPUT62), .ZN(n1084) );
NAND3_X1 U774 ( .A1(G478), .A2(n1087), .A3(KEYINPUT62), .ZN(n1083) );
NOR3_X1 U775 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1077) );
NAND2_X1 U776 ( .A1(G475), .A2(n1091), .ZN(n1076) );
XOR2_X1 U777 ( .A(n1092), .B(n1093), .Z(G72) );
NOR2_X1 U778 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
AND2_X1 U779 ( .A1(G227), .A2(G900), .ZN(n1094) );
NOR2_X1 U780 ( .A1(KEYINPUT39), .A2(n1096), .ZN(n1092) );
NOR2_X1 U781 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U782 ( .A(KEYINPUT30), .B(n1099), .Z(n1098) );
NOR2_X1 U783 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
AND2_X1 U784 ( .A1(n1101), .A2(n1100), .ZN(n1097) );
AND2_X1 U785 ( .A1(n1102), .A2(n1103), .ZN(n1100) );
NAND2_X1 U786 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U787 ( .A(KEYINPUT3), .B(G953), .Z(n1102) );
NAND2_X1 U788 ( .A1(n1106), .A2(n1107), .ZN(n1101) );
NAND2_X1 U789 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
XOR2_X1 U790 ( .A(KEYINPUT34), .B(G953), .Z(n1108) );
XOR2_X1 U791 ( .A(n1110), .B(n1111), .Z(n1106) );
XOR2_X1 U792 ( .A(KEYINPUT23), .B(n1112), .Z(n1111) );
NOR2_X1 U793 ( .A1(n1113), .A2(n1114), .ZN(n1112) );
XOR2_X1 U794 ( .A(KEYINPUT11), .B(n1115), .Z(n1114) );
NOR2_X1 U795 ( .A1(G140), .A2(n1116), .ZN(n1115) );
NAND2_X1 U796 ( .A1(n1117), .A2(n1118), .ZN(G69) );
NAND2_X1 U797 ( .A1(n1119), .A2(n1095), .ZN(n1118) );
XNOR2_X1 U798 ( .A(n1120), .B(n1121), .ZN(n1119) );
NOR2_X1 U799 ( .A1(n1122), .A2(KEYINPUT57), .ZN(n1121) );
NAND2_X1 U800 ( .A1(n1123), .A2(G953), .ZN(n1117) );
XOR2_X1 U801 ( .A(n1120), .B(n1124), .Z(n1123) );
AND2_X1 U802 ( .A1(G224), .A2(G898), .ZN(n1124) );
NAND4_X1 U803 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1120) );
NAND2_X1 U804 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
INV_X1 U805 ( .A(KEYINPUT25), .ZN(n1130) );
XNOR2_X1 U806 ( .A(n1131), .B(n1132), .ZN(n1129) );
NAND2_X1 U807 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
NAND2_X1 U808 ( .A1(KEYINPUT25), .A2(n1135), .ZN(n1127) );
INV_X1 U809 ( .A(n1136), .ZN(n1126) );
NAND2_X1 U810 ( .A1(G953), .A2(n1137), .ZN(n1125) );
XOR2_X1 U811 ( .A(KEYINPUT44), .B(G898), .Z(n1137) );
NOR2_X1 U812 ( .A1(n1138), .A2(n1139), .ZN(G66) );
XOR2_X1 U813 ( .A(KEYINPUT29), .B(n1140), .Z(n1139) );
XOR2_X1 U814 ( .A(n1141), .B(n1142), .Z(n1138) );
NAND2_X1 U815 ( .A1(n1143), .A2(n1082), .ZN(n1141) );
NOR2_X1 U816 ( .A1(n1140), .A2(n1144), .ZN(G63) );
XOR2_X1 U817 ( .A(n1145), .B(n1146), .Z(n1144) );
NAND2_X1 U818 ( .A1(n1143), .A2(G478), .ZN(n1145) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1147), .ZN(G60) );
XOR2_X1 U820 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U821 ( .A1(n1143), .A2(G475), .ZN(n1148) );
XNOR2_X1 U822 ( .A(G104), .B(n1150), .ZN(G6) );
NOR2_X1 U823 ( .A1(n1140), .A2(n1151), .ZN(G57) );
NOR2_X1 U824 ( .A1(n1152), .A2(n1153), .ZN(n1151) );
XOR2_X1 U825 ( .A(n1154), .B(KEYINPUT43), .Z(n1153) );
NAND2_X1 U826 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U827 ( .A1(n1155), .A2(n1156), .ZN(n1152) );
XNOR2_X1 U828 ( .A(n1157), .B(n1158), .ZN(n1156) );
XNOR2_X1 U829 ( .A(n1159), .B(n1160), .ZN(n1157) );
NAND2_X1 U830 ( .A1(n1143), .A2(G472), .ZN(n1159) );
NOR2_X1 U831 ( .A1(n1140), .A2(n1161), .ZN(G54) );
XOR2_X1 U832 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND2_X1 U833 ( .A1(n1143), .A2(G469), .ZN(n1163) );
NAND2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1162) );
NAND2_X1 U835 ( .A1(n1166), .A2(n1167), .ZN(n1165) );
XOR2_X1 U836 ( .A(KEYINPUT48), .B(n1168), .Z(n1164) );
NOR2_X1 U837 ( .A1(n1167), .A2(n1166), .ZN(n1168) );
XNOR2_X1 U838 ( .A(n1169), .B(n1170), .ZN(n1166) );
NOR2_X1 U839 ( .A1(KEYINPUT19), .A2(n1171), .ZN(n1170) );
XOR2_X1 U840 ( .A(n1172), .B(n1173), .Z(n1171) );
XOR2_X1 U841 ( .A(n1174), .B(KEYINPUT18), .Z(n1173) );
NOR2_X1 U842 ( .A1(n1140), .A2(n1175), .ZN(G51) );
NOR2_X1 U843 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
XOR2_X1 U844 ( .A(KEYINPUT15), .B(n1178), .Z(n1177) );
NOR2_X1 U845 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
AND2_X1 U846 ( .A1(n1180), .A2(n1179), .ZN(n1176) );
XNOR2_X1 U847 ( .A(n1181), .B(n1182), .ZN(n1179) );
NAND2_X1 U848 ( .A1(n1183), .A2(n1184), .ZN(n1181) );
NAND2_X1 U849 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U850 ( .A(KEYINPUT55), .B(n1187), .Z(n1183) );
NOR2_X1 U851 ( .A1(n1186), .A2(n1185), .ZN(n1187) );
XNOR2_X1 U852 ( .A(n1188), .B(KEYINPUT13), .ZN(n1185) );
NAND2_X1 U853 ( .A1(n1143), .A2(G210), .ZN(n1180) );
AND2_X1 U854 ( .A1(G902), .A2(n1032), .ZN(n1143) );
NAND3_X1 U855 ( .A1(n1104), .A2(n1189), .A3(n1122), .ZN(n1032) );
AND4_X1 U856 ( .A1(n1190), .A2(n1150), .A3(n1191), .A4(n1192), .ZN(n1122) );
AND4_X1 U857 ( .A1(n1193), .A2(n1194), .A3(n1027), .A4(n1195), .ZN(n1192) );
NAND2_X1 U858 ( .A1(n1025), .A2(n1051), .ZN(n1027) );
AND2_X1 U859 ( .A1(n1071), .A2(n1196), .ZN(n1025) );
AND2_X1 U860 ( .A1(n1197), .A2(n1198), .ZN(n1191) );
NAND3_X1 U861 ( .A1(n1051), .A2(n1196), .A3(n1072), .ZN(n1150) );
AND4_X1 U862 ( .A1(n1068), .A2(n1074), .A3(n1199), .A4(n1200), .ZN(n1196) );
NAND2_X1 U863 ( .A1(n1201), .A2(n1202), .ZN(n1190) );
XOR2_X1 U864 ( .A(n1203), .B(KEYINPUT46), .Z(n1201) );
XNOR2_X1 U865 ( .A(KEYINPUT61), .B(n1105), .ZN(n1189) );
AND4_X1 U866 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1104) );
NOR4_X1 U867 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1207) );
INV_X1 U868 ( .A(n1212), .ZN(n1211) );
INV_X1 U869 ( .A(n1213), .ZN(n1209) );
NAND2_X1 U870 ( .A1(n1059), .A2(n1214), .ZN(n1206) );
XOR2_X1 U871 ( .A(KEYINPUT4), .B(n1215), .Z(n1214) );
NAND3_X1 U872 ( .A1(n1216), .A2(n1071), .A3(n1217), .ZN(n1204) );
AND2_X1 U873 ( .A1(G953), .A2(n1218), .ZN(n1140) );
XOR2_X1 U874 ( .A(KEYINPUT50), .B(G952), .Z(n1218) );
XNOR2_X1 U875 ( .A(n1205), .B(n1219), .ZN(G48) );
NOR2_X1 U876 ( .A1(KEYINPUT40), .A2(n1220), .ZN(n1219) );
NAND3_X1 U877 ( .A1(n1216), .A2(n1072), .A3(n1217), .ZN(n1205) );
XOR2_X1 U878 ( .A(G143), .B(n1221), .Z(G45) );
NOR2_X1 U879 ( .A1(KEYINPUT6), .A2(n1212), .ZN(n1221) );
NAND4_X1 U880 ( .A1(n1217), .A2(n1075), .A3(n1222), .A4(n1223), .ZN(n1212) );
XOR2_X1 U881 ( .A(n1224), .B(n1225), .Z(G42) );
NAND2_X1 U882 ( .A1(n1215), .A2(n1059), .ZN(n1225) );
AND2_X1 U883 ( .A1(n1226), .A2(n1068), .ZN(n1215) );
XNOR2_X1 U884 ( .A(G137), .B(n1227), .ZN(G39) );
NOR2_X1 U885 ( .A1(n1210), .A2(KEYINPUT47), .ZN(n1227) );
AND3_X1 U886 ( .A1(n1216), .A2(n1060), .A3(n1228), .ZN(n1210) );
XNOR2_X1 U887 ( .A(G134), .B(n1105), .ZN(G36) );
NAND3_X1 U888 ( .A1(n1075), .A2(n1071), .A3(n1228), .ZN(n1105) );
XOR2_X1 U889 ( .A(n1229), .B(n1213), .Z(G33) );
NAND3_X1 U890 ( .A1(n1072), .A2(n1075), .A3(n1228), .ZN(n1213) );
AND3_X1 U891 ( .A1(n1068), .A2(n1230), .A3(n1059), .ZN(n1228) );
INV_X1 U892 ( .A(n1044), .ZN(n1059) );
NAND2_X1 U893 ( .A1(n1231), .A2(n1055), .ZN(n1044) );
XOR2_X1 U894 ( .A(n1232), .B(n1233), .Z(G30) );
NAND3_X1 U895 ( .A1(n1071), .A2(n1234), .A3(n1217), .ZN(n1233) );
AND3_X1 U896 ( .A1(n1068), .A2(n1230), .A3(n1051), .ZN(n1217) );
XOR2_X1 U897 ( .A(KEYINPUT37), .B(n1216), .Z(n1234) );
XOR2_X1 U898 ( .A(G101), .B(n1235), .Z(G3) );
NOR3_X1 U899 ( .A1(n1203), .A2(KEYINPUT24), .A3(n1236), .ZN(n1235) );
XOR2_X1 U900 ( .A(G125), .B(n1208), .Z(G27) );
AND3_X1 U901 ( .A1(n1051), .A2(n1069), .A3(n1226), .ZN(n1208) );
AND4_X1 U902 ( .A1(n1072), .A2(n1199), .A3(n1230), .A4(n1040), .ZN(n1226) );
NAND2_X1 U903 ( .A1(n1237), .A2(n1238), .ZN(n1230) );
NAND4_X1 U904 ( .A1(G902), .A2(G953), .A3(n1239), .A4(n1109), .ZN(n1238) );
INV_X1 U905 ( .A(G900), .ZN(n1109) );
XNOR2_X1 U906 ( .A(KEYINPUT42), .B(n1034), .ZN(n1237) );
XNOR2_X1 U907 ( .A(G122), .B(n1198), .ZN(G24) );
NAND3_X1 U908 ( .A1(n1240), .A2(n1074), .A3(n1241), .ZN(n1198) );
NOR3_X1 U909 ( .A1(n1037), .A2(n1242), .A3(n1243), .ZN(n1241) );
XOR2_X1 U910 ( .A(n1244), .B(n1197), .Z(G21) );
NAND3_X1 U911 ( .A1(n1240), .A2(n1060), .A3(n1216), .ZN(n1197) );
NOR2_X1 U912 ( .A1(n1199), .A2(n1074), .ZN(n1216) );
XNOR2_X1 U913 ( .A(G116), .B(n1245), .ZN(G18) );
NAND2_X1 U914 ( .A1(KEYINPUT59), .A2(n1246), .ZN(n1245) );
INV_X1 U915 ( .A(n1194), .ZN(n1246) );
NAND3_X1 U916 ( .A1(n1075), .A2(n1071), .A3(n1240), .ZN(n1194) );
NOR2_X1 U917 ( .A1(n1222), .A2(n1242), .ZN(n1071) );
INV_X1 U918 ( .A(n1243), .ZN(n1222) );
XOR2_X1 U919 ( .A(n1247), .B(n1195), .Z(G15) );
NAND3_X1 U920 ( .A1(n1240), .A2(n1075), .A3(n1072), .ZN(n1195) );
NOR2_X1 U921 ( .A1(n1223), .A2(n1243), .ZN(n1072) );
INV_X1 U922 ( .A(n1242), .ZN(n1223) );
INV_X1 U923 ( .A(n1203), .ZN(n1075) );
NAND2_X1 U924 ( .A1(n1037), .A2(n1074), .ZN(n1203) );
INV_X1 U925 ( .A(n1040), .ZN(n1074) );
AND3_X1 U926 ( .A1(n1069), .A2(n1200), .A3(n1051), .ZN(n1240) );
NAND2_X1 U927 ( .A1(n1248), .A2(n1249), .ZN(n1069) );
OR2_X1 U928 ( .A1(n1056), .A2(KEYINPUT45), .ZN(n1249) );
NAND3_X1 U929 ( .A1(n1250), .A2(n1067), .A3(KEYINPUT45), .ZN(n1248) );
XNOR2_X1 U930 ( .A(G110), .B(n1193), .ZN(G12) );
NAND3_X1 U931 ( .A1(n1199), .A2(n1040), .A3(n1202), .ZN(n1193) );
INV_X1 U932 ( .A(n1236), .ZN(n1202) );
NAND4_X1 U933 ( .A1(n1060), .A2(n1051), .A3(n1068), .A4(n1200), .ZN(n1236) );
NAND2_X1 U934 ( .A1(n1034), .A2(n1251), .ZN(n1200) );
NAND4_X1 U935 ( .A1(G902), .A2(G953), .A3(n1239), .A4(n1252), .ZN(n1251) );
INV_X1 U936 ( .A(G898), .ZN(n1252) );
NAND3_X1 U937 ( .A1(n1239), .A2(n1095), .A3(G952), .ZN(n1034) );
NAND2_X1 U938 ( .A1(G234), .A2(G237), .ZN(n1239) );
INV_X1 U939 ( .A(n1056), .ZN(n1068) );
NAND2_X1 U940 ( .A1(n1066), .A2(n1067), .ZN(n1056) );
NAND2_X1 U941 ( .A1(G221), .A2(n1253), .ZN(n1067) );
INV_X1 U942 ( .A(n1250), .ZN(n1066) );
XOR2_X1 U943 ( .A(n1254), .B(G469), .Z(n1250) );
NAND2_X1 U944 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
XOR2_X1 U945 ( .A(n1257), .B(n1167), .Z(n1255) );
XOR2_X1 U946 ( .A(n1258), .B(n1259), .Z(n1167) );
XOR2_X1 U947 ( .A(G140), .B(G110), .Z(n1259) );
NAND2_X1 U948 ( .A1(G227), .A2(n1095), .ZN(n1258) );
NAND2_X1 U949 ( .A1(n1260), .A2(KEYINPUT36), .ZN(n1257) );
XOR2_X1 U950 ( .A(n1261), .B(n1110), .Z(n1260) );
XNOR2_X1 U951 ( .A(n1174), .B(n1169), .ZN(n1110) );
NAND2_X1 U952 ( .A1(n1262), .A2(n1263), .ZN(n1174) );
NAND2_X1 U953 ( .A1(G128), .A2(n1264), .ZN(n1263) );
XOR2_X1 U954 ( .A(n1265), .B(KEYINPUT0), .Z(n1262) );
NAND2_X1 U955 ( .A1(n1266), .A2(n1232), .ZN(n1265) );
XOR2_X1 U956 ( .A(n1172), .B(KEYINPUT5), .Z(n1261) );
XNOR2_X1 U957 ( .A(n1267), .B(n1268), .ZN(n1172) );
NOR2_X1 U958 ( .A1(KEYINPUT54), .A2(n1269), .ZN(n1268) );
INV_X1 U959 ( .A(n1026), .ZN(n1051) );
NAND2_X1 U960 ( .A1(n1270), .A2(n1055), .ZN(n1026) );
NAND2_X1 U961 ( .A1(G214), .A2(n1271), .ZN(n1055) );
OR2_X1 U962 ( .A1(G237), .A2(G902), .ZN(n1271) );
XNOR2_X1 U963 ( .A(n1231), .B(KEYINPUT16), .ZN(n1270) );
INV_X1 U964 ( .A(n1054), .ZN(n1231) );
NAND2_X1 U965 ( .A1(n1272), .A2(n1273), .ZN(n1054) );
NAND2_X1 U966 ( .A1(G210), .A2(n1274), .ZN(n1273) );
NAND2_X1 U967 ( .A1(n1256), .A2(n1275), .ZN(n1274) );
NAND2_X1 U968 ( .A1(G237), .A2(n1276), .ZN(n1275) );
INV_X1 U969 ( .A(n1277), .ZN(n1276) );
NAND3_X1 U970 ( .A1(n1278), .A2(n1256), .A3(n1277), .ZN(n1272) );
XNOR2_X1 U971 ( .A(n1279), .B(n1188), .ZN(n1277) );
XNOR2_X1 U972 ( .A(n1280), .B(n1116), .ZN(n1188) );
XOR2_X1 U973 ( .A(n1186), .B(n1182), .Z(n1279) );
NOR2_X1 U974 ( .A1(n1135), .A2(n1136), .ZN(n1182) );
NOR3_X1 U975 ( .A1(n1281), .A2(n1133), .A3(n1134), .ZN(n1136) );
NAND2_X1 U976 ( .A1(n1282), .A2(n1283), .ZN(n1135) );
OR3_X1 U977 ( .A1(n1132), .A2(n1284), .A3(n1134), .ZN(n1283) );
NAND2_X1 U978 ( .A1(n1285), .A2(n1134), .ZN(n1282) );
XNOR2_X1 U979 ( .A(n1286), .B(n1287), .ZN(n1134) );
XOR2_X1 U980 ( .A(G119), .B(n1288), .Z(n1287) );
NOR2_X1 U981 ( .A1(G113), .A2(KEYINPUT31), .ZN(n1288) );
NAND2_X1 U982 ( .A1(KEYINPUT41), .A2(n1289), .ZN(n1286) );
XOR2_X1 U983 ( .A(n1284), .B(n1132), .Z(n1285) );
INV_X1 U984 ( .A(n1281), .ZN(n1132) );
XNOR2_X1 U985 ( .A(G110), .B(G122), .ZN(n1281) );
INV_X1 U986 ( .A(n1133), .ZN(n1284) );
XNOR2_X1 U987 ( .A(n1269), .B(n1267), .ZN(n1133) );
XNOR2_X1 U988 ( .A(n1290), .B(KEYINPUT10), .ZN(n1267) );
XOR2_X1 U989 ( .A(G104), .B(G107), .Z(n1269) );
NAND2_X1 U990 ( .A1(G224), .A2(n1095), .ZN(n1186) );
NAND2_X1 U991 ( .A1(G210), .A2(G237), .ZN(n1278) );
INV_X1 U992 ( .A(n1046), .ZN(n1060) );
NAND2_X1 U993 ( .A1(n1242), .A2(n1243), .ZN(n1046) );
NOR2_X1 U994 ( .A1(n1291), .A2(n1090), .ZN(n1243) );
NOR3_X1 U995 ( .A1(G475), .A2(G902), .A3(n1292), .ZN(n1090) );
AND2_X1 U996 ( .A1(n1293), .A2(n1091), .ZN(n1291) );
NAND2_X1 U997 ( .A1(n1149), .A2(n1256), .ZN(n1091) );
INV_X1 U998 ( .A(n1292), .ZN(n1149) );
XNOR2_X1 U999 ( .A(n1294), .B(n1295), .ZN(n1292) );
XOR2_X1 U1000 ( .A(n1296), .B(n1297), .Z(n1295) );
XOR2_X1 U1001 ( .A(n1298), .B(n1299), .Z(n1297) );
AND2_X1 U1002 ( .A1(G214), .A2(n1300), .ZN(n1299) );
NAND2_X1 U1003 ( .A1(KEYINPUT7), .A2(n1247), .ZN(n1298) );
NAND2_X1 U1004 ( .A1(KEYINPUT49), .A2(n1229), .ZN(n1296) );
XOR2_X1 U1005 ( .A(n1301), .B(n1264), .Z(n1294) );
INV_X1 U1006 ( .A(n1266), .ZN(n1264) );
NAND3_X1 U1007 ( .A1(n1302), .A2(n1303), .A3(n1304), .ZN(n1301) );
NAND2_X1 U1008 ( .A1(n1305), .A2(n1224), .ZN(n1304) );
XOR2_X1 U1009 ( .A(G125), .B(n1306), .Z(n1305) );
NAND3_X1 U1010 ( .A1(G140), .A2(G125), .A3(n1306), .ZN(n1303) );
NAND2_X1 U1011 ( .A1(n1113), .A2(n1307), .ZN(n1302) );
INV_X1 U1012 ( .A(n1306), .ZN(n1307) );
XOR2_X1 U1013 ( .A(G104), .B(G122), .Z(n1306) );
NOR2_X1 U1014 ( .A1(n1224), .A2(G125), .ZN(n1113) );
INV_X1 U1015 ( .A(G140), .ZN(n1224) );
XNOR2_X1 U1016 ( .A(G475), .B(KEYINPUT56), .ZN(n1293) );
NOR2_X1 U1017 ( .A1(n1308), .A2(n1089), .ZN(n1242) );
NOR2_X1 U1018 ( .A1(n1087), .A2(G478), .ZN(n1089) );
AND2_X1 U1019 ( .A1(G478), .A2(n1087), .ZN(n1308) );
NAND2_X1 U1020 ( .A1(n1146), .A2(n1256), .ZN(n1087) );
XNOR2_X1 U1021 ( .A(n1309), .B(n1310), .ZN(n1146) );
XOR2_X1 U1022 ( .A(n1289), .B(n1311), .Z(n1310) );
XOR2_X1 U1023 ( .A(n1312), .B(n1313), .Z(n1311) );
NOR2_X1 U1024 ( .A1(KEYINPUT63), .A2(n1314), .ZN(n1313) );
XOR2_X1 U1025 ( .A(n1232), .B(n1315), .Z(n1314) );
INV_X1 U1026 ( .A(G128), .ZN(n1232) );
NAND3_X1 U1027 ( .A1(G217), .A2(n1095), .A3(G234), .ZN(n1312) );
XOR2_X1 U1028 ( .A(n1020), .B(n1316), .Z(n1309) );
XOR2_X1 U1029 ( .A(G134), .B(G122), .Z(n1316) );
INV_X1 U1030 ( .A(G107), .ZN(n1020) );
NAND3_X1 U1031 ( .A1(n1317), .A2(n1318), .A3(n1319), .ZN(n1040) );
INV_X1 U1032 ( .A(n1088), .ZN(n1319) );
NOR2_X1 U1033 ( .A1(n1081), .A2(n1082), .ZN(n1088) );
OR2_X1 U1034 ( .A1(n1082), .A2(KEYINPUT33), .ZN(n1318) );
NAND3_X1 U1035 ( .A1(n1082), .A2(n1081), .A3(KEYINPUT33), .ZN(n1317) );
NAND2_X1 U1036 ( .A1(n1142), .A2(n1256), .ZN(n1081) );
XNOR2_X1 U1037 ( .A(n1320), .B(n1321), .ZN(n1142) );
NOR2_X1 U1038 ( .A1(KEYINPUT35), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1039 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1040 ( .A(n1325), .B(n1326), .Z(n1324) );
NOR2_X1 U1041 ( .A1(KEYINPUT1), .A2(G140), .ZN(n1326) );
XOR2_X1 U1042 ( .A(G110), .B(n1244), .Z(n1325) );
XOR2_X1 U1043 ( .A(n1116), .B(n1327), .Z(n1323) );
XOR2_X1 U1044 ( .A(G146), .B(G128), .Z(n1327) );
INV_X1 U1045 ( .A(G125), .ZN(n1116) );
XNOR2_X1 U1046 ( .A(G137), .B(n1328), .ZN(n1320) );
NOR4_X1 U1047 ( .A1(KEYINPUT53), .A2(n1329), .A3(n1330), .A4(n1331), .ZN(n1328) );
INV_X1 U1048 ( .A(G221), .ZN(n1331) );
INV_X1 U1049 ( .A(G234), .ZN(n1330) );
XOR2_X1 U1050 ( .A(n1095), .B(KEYINPUT51), .Z(n1329) );
INV_X1 U1051 ( .A(G953), .ZN(n1095) );
AND2_X1 U1052 ( .A1(G217), .A2(n1253), .ZN(n1082) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1256), .ZN(n1253) );
INV_X1 U1054 ( .A(n1037), .ZN(n1199) );
XOR2_X1 U1055 ( .A(n1086), .B(n1332), .Z(n1037) );
NOR2_X1 U1056 ( .A1(G472), .A2(KEYINPUT32), .ZN(n1332) );
NAND2_X1 U1057 ( .A1(n1333), .A2(n1256), .ZN(n1086) );
INV_X1 U1058 ( .A(G902), .ZN(n1256) );
XOR2_X1 U1059 ( .A(n1334), .B(n1335), .Z(n1333) );
XOR2_X1 U1060 ( .A(n1336), .B(n1337), .Z(n1335) );
NAND2_X1 U1061 ( .A1(KEYINPUT17), .A2(n1160), .ZN(n1337) );
NAND3_X1 U1062 ( .A1(n1338), .A2(n1339), .A3(n1340), .ZN(n1160) );
OR2_X1 U1063 ( .A1(n1247), .A2(n1341), .ZN(n1340) );
NAND3_X1 U1064 ( .A1(n1341), .A2(n1247), .A3(KEYINPUT58), .ZN(n1339) );
INV_X1 U1065 ( .A(G113), .ZN(n1247) );
NOR2_X1 U1066 ( .A1(KEYINPUT22), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1067 ( .A1(n1342), .A2(n1343), .ZN(n1338) );
INV_X1 U1068 ( .A(KEYINPUT58), .ZN(n1343) );
XOR2_X1 U1069 ( .A(n1344), .B(n1289), .Z(n1342) );
XNOR2_X1 U1070 ( .A(G116), .B(KEYINPUT38), .ZN(n1289) );
XOR2_X1 U1071 ( .A(n1244), .B(KEYINPUT8), .Z(n1344) );
INV_X1 U1072 ( .A(G119), .ZN(n1244) );
NAND2_X1 U1073 ( .A1(KEYINPUT27), .A2(n1155), .ZN(n1336) );
AND2_X1 U1074 ( .A1(n1345), .A2(n1346), .ZN(n1155) );
NAND2_X1 U1075 ( .A1(n1347), .A2(n1290), .ZN(n1346) );
INV_X1 U1076 ( .A(G101), .ZN(n1290) );
NAND2_X1 U1077 ( .A1(n1300), .A2(G210), .ZN(n1347) );
NAND3_X1 U1078 ( .A1(n1300), .A2(G210), .A3(G101), .ZN(n1345) );
NOR2_X1 U1079 ( .A1(G953), .A2(G237), .ZN(n1300) );
NAND2_X1 U1080 ( .A1(n1348), .A2(n1349), .ZN(n1334) );
NAND2_X1 U1081 ( .A1(n1158), .A2(n1350), .ZN(n1349) );
INV_X1 U1082 ( .A(KEYINPUT2), .ZN(n1350) );
XOR2_X1 U1083 ( .A(n1351), .B(n1169), .Z(n1158) );
NAND3_X1 U1084 ( .A1(n1351), .A2(n1169), .A3(KEYINPUT2), .ZN(n1348) );
XNOR2_X1 U1085 ( .A(n1352), .B(n1353), .ZN(n1169) );
XOR2_X1 U1086 ( .A(KEYINPUT26), .B(G137), .Z(n1353) );
XOR2_X1 U1087 ( .A(n1229), .B(G134), .Z(n1352) );
INV_X1 U1088 ( .A(G131), .ZN(n1229) );
XNOR2_X1 U1089 ( .A(n1280), .B(KEYINPUT28), .ZN(n1351) );
XOR2_X1 U1090 ( .A(n1354), .B(G128), .Z(n1280) );
NAND2_X1 U1091 ( .A1(n1355), .A2(KEYINPUT52), .ZN(n1354) );
XOR2_X1 U1092 ( .A(n1266), .B(n1356), .Z(n1355) );
XOR2_X1 U1093 ( .A(KEYINPUT60), .B(KEYINPUT12), .Z(n1356) );
XOR2_X1 U1094 ( .A(n1220), .B(n1315), .Z(n1266) );
XOR2_X1 U1095 ( .A(G143), .B(KEYINPUT9), .Z(n1315) );
INV_X1 U1096 ( .A(G146), .ZN(n1220) );
endmodule


