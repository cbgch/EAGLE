//Key = 0101011011000011011000001000010011010100100010000111001100011001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
n1369, n1370, n1371, n1372, n1373, n1374, n1375;

XOR2_X1 U754 ( .A(G107), .B(n1049), .Z(G9) );
NOR2_X1 U755 ( .A1(n1050), .A2(n1051), .ZN(G75) );
NOR4_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1051) );
INV_X1 U757 ( .A(G952), .ZN(n1055) );
NOR2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NOR2_X1 U759 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR3_X1 U760 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1059) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
INV_X1 U762 ( .A(n1065), .ZN(n1061) );
NAND3_X1 U763 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1060) );
NAND2_X1 U764 ( .A1(n1069), .A2(n1070), .ZN(n1067) );
OR3_X1 U765 ( .A1(n1071), .A2(n1072), .A3(n1069), .ZN(n1066) );
NOR2_X1 U766 ( .A1(n1073), .A2(n1074), .ZN(n1058) );
NOR2_X1 U767 ( .A1(n1075), .A2(n1076), .ZN(n1073) );
NOR2_X1 U768 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
XOR2_X1 U769 ( .A(KEYINPUT6), .B(n1079), .Z(n1078) );
XOR2_X1 U770 ( .A(n1080), .B(KEYINPUT21), .Z(n1077) );
NAND3_X1 U771 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1052) );
NAND3_X1 U772 ( .A1(n1068), .A2(n1084), .A3(n1085), .ZN(n1083) );
INV_X1 U773 ( .A(n1074), .ZN(n1085) );
NAND3_X1 U774 ( .A1(n1086), .A2(n1065), .A3(n1087), .ZN(n1074) );
NAND2_X1 U775 ( .A1(n1088), .A2(n1089), .ZN(n1084) );
NOR3_X1 U776 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(n1050) );
NOR2_X1 U777 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
INV_X1 U778 ( .A(KEYINPUT40), .ZN(n1094) );
NOR2_X1 U779 ( .A1(G953), .A2(G952), .ZN(n1093) );
NOR2_X1 U780 ( .A1(KEYINPUT40), .A2(n1095), .ZN(n1091) );
INV_X1 U781 ( .A(n1081), .ZN(n1090) );
NAND4_X1 U782 ( .A1(n1096), .A2(n1097), .A3(n1098), .A4(n1099), .ZN(n1081) );
NOR4_X1 U783 ( .A1(n1100), .A2(n1101), .A3(n1069), .A4(n1102), .ZN(n1099) );
XNOR2_X1 U784 ( .A(G469), .B(n1103), .ZN(n1102) );
NOR3_X1 U785 ( .A1(n1104), .A2(n1105), .A3(n1106), .ZN(n1098) );
NOR2_X1 U786 ( .A1(n1107), .A2(n1108), .ZN(n1104) );
XOR2_X1 U787 ( .A(KEYINPUT38), .B(G475), .Z(n1108) );
NAND2_X1 U788 ( .A1(G478), .A2(n1109), .ZN(n1097) );
NAND2_X1 U789 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U790 ( .A1(KEYINPUT46), .A2(n1112), .ZN(n1111) );
NAND3_X1 U791 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1096) );
INV_X1 U792 ( .A(KEYINPUT46), .ZN(n1115) );
NAND2_X1 U793 ( .A1(n1116), .A2(n1112), .ZN(n1114) );
INV_X1 U794 ( .A(KEYINPUT45), .ZN(n1112) );
NAND2_X1 U795 ( .A1(n1110), .A2(n1117), .ZN(n1113) );
OR2_X1 U796 ( .A1(G478), .A2(KEYINPUT45), .ZN(n1117) );
XOR2_X1 U797 ( .A(n1118), .B(n1119), .Z(G72) );
XOR2_X1 U798 ( .A(n1120), .B(n1121), .Z(n1119) );
NAND4_X1 U799 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121) );
NAND2_X1 U800 ( .A1(KEYINPUT7), .A2(n1126), .ZN(n1125) );
NAND2_X1 U801 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XNOR2_X1 U802 ( .A(KEYINPUT20), .B(n1129), .ZN(n1128) );
NAND2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(n1124) );
INV_X1 U804 ( .A(KEYINPUT7), .ZN(n1131) );
NAND2_X1 U805 ( .A1(n1132), .A2(n1133), .ZN(n1130) );
NAND2_X1 U806 ( .A1(KEYINPUT20), .A2(n1129), .ZN(n1133) );
OR3_X1 U807 ( .A1(n1134), .A2(KEYINPUT20), .A3(n1129), .ZN(n1132) );
NAND2_X1 U808 ( .A1(n1129), .A2(n1134), .ZN(n1123) );
INV_X1 U809 ( .A(n1127), .ZN(n1134) );
XOR2_X1 U810 ( .A(n1135), .B(n1136), .Z(n1127) );
XOR2_X1 U811 ( .A(n1137), .B(n1138), .Z(n1129) );
XOR2_X1 U812 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U813 ( .A1(KEYINPUT33), .A2(n1141), .ZN(n1139) );
NAND2_X1 U814 ( .A1(G953), .A2(n1142), .ZN(n1122) );
NAND2_X1 U815 ( .A1(n1082), .A2(n1143), .ZN(n1120) );
NAND2_X1 U816 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U817 ( .A(n1146), .B(KEYINPUT12), .Z(n1144) );
NOR2_X1 U818 ( .A1(n1147), .A2(n1082), .ZN(n1118) );
NOR2_X1 U819 ( .A1(n1148), .A2(n1142), .ZN(n1147) );
XOR2_X1 U820 ( .A(n1149), .B(n1150), .Z(G69) );
XOR2_X1 U821 ( .A(n1151), .B(n1152), .Z(n1150) );
NAND2_X1 U822 ( .A1(G953), .A2(n1153), .ZN(n1152) );
NAND2_X1 U823 ( .A1(G898), .A2(G224), .ZN(n1153) );
NAND2_X1 U824 ( .A1(n1154), .A2(n1155), .ZN(n1151) );
NAND2_X1 U825 ( .A1(G953), .A2(n1156), .ZN(n1155) );
XOR2_X1 U826 ( .A(n1157), .B(n1158), .Z(n1154) );
NOR2_X1 U827 ( .A1(KEYINPUT56), .A2(n1159), .ZN(n1158) );
NOR2_X1 U828 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
XOR2_X1 U829 ( .A(n1162), .B(KEYINPUT32), .Z(n1161) );
NOR2_X1 U830 ( .A1(n1163), .A2(n1164), .ZN(n1160) );
NOR2_X1 U831 ( .A1(n1165), .A2(G953), .ZN(n1149) );
NOR2_X1 U832 ( .A1(n1095), .A2(n1166), .ZN(G66) );
NOR2_X1 U833 ( .A1(n1167), .A2(n1168), .ZN(n1166) );
XOR2_X1 U834 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U835 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
AND2_X1 U836 ( .A1(n1173), .A2(KEYINPUT49), .ZN(n1169) );
NOR2_X1 U837 ( .A1(KEYINPUT49), .A2(n1173), .ZN(n1167) );
NOR2_X1 U838 ( .A1(n1095), .A2(n1174), .ZN(G63) );
NOR3_X1 U839 ( .A1(n1175), .A2(n1110), .A3(n1176), .ZN(n1174) );
NOR2_X1 U840 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
AND2_X1 U841 ( .A1(n1053), .A2(G478), .ZN(n1177) );
XOR2_X1 U842 ( .A(KEYINPUT2), .B(n1179), .Z(n1175) );
AND3_X1 U843 ( .A1(n1180), .A2(n1178), .A3(G478), .ZN(n1179) );
NOR2_X1 U844 ( .A1(n1095), .A2(n1181), .ZN(G60) );
XNOR2_X1 U845 ( .A(n1182), .B(n1183), .ZN(n1181) );
AND2_X1 U846 ( .A1(G475), .A2(n1180), .ZN(n1183) );
XOR2_X1 U847 ( .A(n1184), .B(n1185), .Z(G6) );
NOR3_X1 U848 ( .A1(n1088), .A2(n1186), .A3(n1070), .ZN(n1185) );
NOR2_X1 U849 ( .A1(KEYINPUT22), .A2(n1187), .ZN(n1184) );
NOR2_X1 U850 ( .A1(n1095), .A2(n1188), .ZN(G57) );
XOR2_X1 U851 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U852 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
NOR2_X1 U853 ( .A1(n1193), .A2(n1194), .ZN(n1192) );
XNOR2_X1 U854 ( .A(KEYINPUT61), .B(n1195), .ZN(n1194) );
INV_X1 U855 ( .A(n1196), .ZN(n1193) );
NOR2_X1 U856 ( .A1(n1196), .A2(n1195), .ZN(n1191) );
NAND2_X1 U857 ( .A1(n1180), .A2(G472), .ZN(n1195) );
NAND3_X1 U858 ( .A1(n1197), .A2(n1198), .A3(n1199), .ZN(n1196) );
NAND2_X1 U859 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U860 ( .A1(n1202), .A2(n1203), .ZN(n1198) );
NAND2_X1 U861 ( .A1(KEYINPUT15), .A2(n1204), .ZN(n1203) );
XOR2_X1 U862 ( .A(n1200), .B(KEYINPUT50), .Z(n1204) );
OR3_X1 U863 ( .A1(n1201), .A2(n1200), .A3(n1202), .ZN(n1197) );
XOR2_X1 U864 ( .A(n1205), .B(n1206), .Z(n1202) );
INV_X1 U865 ( .A(KEYINPUT15), .ZN(n1201) );
XOR2_X1 U866 ( .A(n1207), .B(n1208), .Z(n1189) );
INV_X1 U867 ( .A(G101), .ZN(n1208) );
NOR2_X1 U868 ( .A1(n1209), .A2(n1210), .ZN(G54) );
XOR2_X1 U869 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U870 ( .A(n1213), .B(n1214), .Z(n1212) );
NAND2_X1 U871 ( .A1(n1215), .A2(KEYINPUT35), .ZN(n1213) );
XOR2_X1 U872 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U873 ( .A(n1218), .B(n1219), .Z(n1216) );
NAND2_X1 U874 ( .A1(KEYINPUT14), .A2(n1137), .ZN(n1218) );
XOR2_X1 U875 ( .A(KEYINPUT39), .B(n1220), .Z(n1211) );
AND2_X1 U876 ( .A1(G469), .A2(n1180), .ZN(n1220) );
INV_X1 U877 ( .A(n1172), .ZN(n1180) );
NOR2_X1 U878 ( .A1(n1082), .A2(n1221), .ZN(n1209) );
XOR2_X1 U879 ( .A(KEYINPUT31), .B(G952), .Z(n1221) );
NOR2_X1 U880 ( .A1(n1095), .A2(n1222), .ZN(G51) );
XOR2_X1 U881 ( .A(n1223), .B(n1224), .Z(n1222) );
XOR2_X1 U882 ( .A(n1225), .B(n1206), .Z(n1224) );
XOR2_X1 U883 ( .A(n1226), .B(n1227), .Z(n1223) );
NOR2_X1 U884 ( .A1(G125), .A2(KEYINPUT23), .ZN(n1227) );
XOR2_X1 U885 ( .A(n1228), .B(n1229), .Z(n1226) );
NOR2_X1 U886 ( .A1(n1230), .A2(n1172), .ZN(n1229) );
NAND2_X1 U887 ( .A1(G902), .A2(n1053), .ZN(n1172) );
NAND3_X1 U888 ( .A1(n1145), .A2(n1146), .A3(n1165), .ZN(n1053) );
AND4_X1 U889 ( .A1(n1231), .A2(n1232), .A3(n1233), .A4(n1234), .ZN(n1165) );
NOR4_X1 U890 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1049), .ZN(n1234) );
NOR3_X1 U891 ( .A1(n1070), .A2(n1186), .A3(n1089), .ZN(n1049) );
NOR4_X1 U892 ( .A1(n1238), .A2(n1239), .A3(n1070), .A4(n1088), .ZN(n1237) );
INV_X1 U893 ( .A(n1240), .ZN(n1088) );
INV_X1 U894 ( .A(n1086), .ZN(n1070) );
XOR2_X1 U895 ( .A(n1241), .B(KEYINPUT36), .Z(n1238) );
AND2_X1 U896 ( .A1(n1242), .A2(n1243), .ZN(n1233) );
AND4_X1 U897 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1145) );
NOR4_X1 U898 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1247) );
NOR2_X1 U899 ( .A1(n1082), .A2(G952), .ZN(n1095) );
XNOR2_X1 U900 ( .A(G146), .B(n1246), .ZN(G48) );
NAND4_X1 U901 ( .A1(n1252), .A2(n1240), .A3(n1076), .A4(n1253), .ZN(n1246) );
XOR2_X1 U902 ( .A(G143), .B(n1254), .Z(G45) );
NOR2_X1 U903 ( .A1(KEYINPUT11), .A2(n1244), .ZN(n1254) );
NAND4_X1 U904 ( .A1(n1072), .A2(n1076), .A3(n1255), .A4(n1256), .ZN(n1244) );
AND4_X1 U905 ( .A1(n1257), .A2(n1064), .A3(n1258), .A4(n1259), .ZN(n1256) );
NAND2_X1 U906 ( .A1(n1260), .A2(n1261), .ZN(G42) );
NAND2_X1 U907 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
XOR2_X1 U908 ( .A(KEYINPUT44), .B(n1264), .Z(n1260) );
NOR2_X1 U909 ( .A1(n1262), .A2(n1263), .ZN(n1264) );
INV_X1 U910 ( .A(G140), .ZN(n1263) );
INV_X1 U911 ( .A(n1245), .ZN(n1262) );
NAND3_X1 U912 ( .A1(n1240), .A2(n1071), .A3(n1265), .ZN(n1245) );
INV_X1 U913 ( .A(n1266), .ZN(n1071) );
XOR2_X1 U914 ( .A(G137), .B(n1251), .Z(G39) );
AND2_X1 U915 ( .A1(n1265), .A2(n1267), .ZN(n1251) );
XOR2_X1 U916 ( .A(G134), .B(n1250), .Z(G36) );
AND3_X1 U917 ( .A1(n1072), .A2(n1268), .A3(n1265), .ZN(n1250) );
XNOR2_X1 U918 ( .A(G131), .B(n1146), .ZN(G33) );
NAND3_X1 U919 ( .A1(n1072), .A2(n1240), .A3(n1265), .ZN(n1146) );
AND3_X1 U920 ( .A1(n1087), .A2(n1076), .A3(n1255), .ZN(n1265) );
INV_X1 U921 ( .A(n1069), .ZN(n1087) );
NAND2_X1 U922 ( .A1(n1063), .A2(n1064), .ZN(n1069) );
XOR2_X1 U923 ( .A(n1269), .B(n1270), .Z(G30) );
NAND2_X1 U924 ( .A1(KEYINPUT17), .A2(n1249), .ZN(n1270) );
AND4_X1 U925 ( .A1(n1252), .A2(n1268), .A3(n1253), .A4(n1271), .ZN(n1249) );
INV_X1 U926 ( .A(n1241), .ZN(n1271) );
XOR2_X1 U927 ( .A(G101), .B(n1272), .Z(G3) );
NOR2_X1 U928 ( .A1(KEYINPUT10), .A2(n1231), .ZN(n1272) );
NAND3_X1 U929 ( .A1(n1273), .A2(n1274), .A3(n1072), .ZN(n1231) );
XOR2_X1 U930 ( .A(n1248), .B(n1275), .Z(G27) );
NOR2_X1 U931 ( .A1(KEYINPUT48), .A2(n1135), .ZN(n1275) );
INV_X1 U932 ( .A(G125), .ZN(n1135) );
AND4_X1 U933 ( .A1(n1252), .A2(n1240), .A3(n1276), .A4(n1068), .ZN(n1248) );
AND4_X1 U934 ( .A1(n1255), .A2(n1100), .A3(n1259), .A4(n1064), .ZN(n1252) );
AND2_X1 U935 ( .A1(n1277), .A2(n1065), .ZN(n1255) );
NAND2_X1 U936 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
NAND3_X1 U937 ( .A1(G953), .A2(n1142), .A3(G902), .ZN(n1279) );
INV_X1 U938 ( .A(G900), .ZN(n1142) );
XOR2_X1 U939 ( .A(n1280), .B(G122), .Z(G24) );
NAND2_X1 U940 ( .A1(KEYINPUT54), .A2(n1232), .ZN(n1280) );
NAND4_X1 U941 ( .A1(n1281), .A2(n1086), .A3(n1258), .A4(n1257), .ZN(n1232) );
NOR2_X1 U942 ( .A1(n1253), .A2(n1100), .ZN(n1086) );
XOR2_X1 U943 ( .A(n1282), .B(n1243), .Z(G21) );
NAND2_X1 U944 ( .A1(n1267), .A2(n1281), .ZN(n1243) );
AND3_X1 U945 ( .A1(n1100), .A2(n1253), .A3(n1273), .ZN(n1267) );
INV_X1 U946 ( .A(n1276), .ZN(n1253) );
XNOR2_X1 U947 ( .A(G116), .B(n1242), .ZN(G18) );
NAND3_X1 U948 ( .A1(n1281), .A2(n1268), .A3(n1072), .ZN(n1242) );
INV_X1 U949 ( .A(n1089), .ZN(n1268) );
NAND2_X1 U950 ( .A1(n1283), .A2(n1258), .ZN(n1089) );
XOR2_X1 U951 ( .A(G113), .B(n1236), .Z(G15) );
AND3_X1 U952 ( .A1(n1240), .A2(n1281), .A3(n1072), .ZN(n1236) );
NOR2_X1 U953 ( .A1(n1100), .A2(n1276), .ZN(n1072) );
NOR2_X1 U954 ( .A1(n1239), .A2(n1284), .ZN(n1281) );
INV_X1 U955 ( .A(n1068), .ZN(n1284) );
NAND2_X1 U956 ( .A1(n1285), .A2(n1286), .ZN(n1068) );
NAND2_X1 U957 ( .A1(n1076), .A2(n1287), .ZN(n1286) );
INV_X1 U958 ( .A(KEYINPUT55), .ZN(n1287) );
NAND3_X1 U959 ( .A1(n1079), .A2(n1080), .A3(KEYINPUT55), .ZN(n1285) );
NOR2_X1 U960 ( .A1(n1258), .A2(n1283), .ZN(n1240) );
XOR2_X1 U961 ( .A(n1235), .B(n1288), .Z(G12) );
NOR2_X1 U962 ( .A1(KEYINPUT57), .A2(n1289), .ZN(n1288) );
NOR3_X1 U963 ( .A1(n1266), .A2(n1186), .A3(n1057), .ZN(n1235) );
INV_X1 U964 ( .A(n1273), .ZN(n1057) );
NOR2_X1 U965 ( .A1(n1258), .A2(n1257), .ZN(n1273) );
INV_X1 U966 ( .A(n1283), .ZN(n1257) );
NOR2_X1 U967 ( .A1(n1290), .A2(n1105), .ZN(n1283) );
AND2_X1 U968 ( .A1(G475), .A2(n1107), .ZN(n1105) );
NOR2_X1 U969 ( .A1(n1107), .A2(G475), .ZN(n1290) );
NAND2_X1 U970 ( .A1(n1182), .A2(n1291), .ZN(n1107) );
XNOR2_X1 U971 ( .A(n1292), .B(n1293), .ZN(n1182) );
XOR2_X1 U972 ( .A(n1294), .B(n1295), .Z(n1293) );
XOR2_X1 U973 ( .A(G122), .B(G113), .Z(n1295) );
XOR2_X1 U974 ( .A(KEYINPUT29), .B(G125), .Z(n1294) );
XOR2_X1 U975 ( .A(n1296), .B(n1297), .Z(n1292) );
XOR2_X1 U976 ( .A(n1298), .B(n1299), .Z(n1297) );
NOR2_X1 U977 ( .A1(KEYINPUT30), .A2(n1300), .ZN(n1299) );
NOR2_X1 U978 ( .A1(KEYINPUT58), .A2(n1136), .ZN(n1298) );
XOR2_X1 U979 ( .A(n1187), .B(n1301), .Z(n1296) );
NOR2_X1 U980 ( .A1(KEYINPUT52), .A2(n1302), .ZN(n1301) );
XOR2_X1 U981 ( .A(n1303), .B(n1304), .Z(n1302) );
XNOR2_X1 U982 ( .A(G131), .B(n1305), .ZN(n1304) );
AND3_X1 U983 ( .A1(G214), .A2(n1082), .A3(n1306), .ZN(n1305) );
NAND2_X1 U984 ( .A1(KEYINPUT37), .A2(n1307), .ZN(n1303) );
INV_X1 U985 ( .A(G104), .ZN(n1187) );
NAND2_X1 U986 ( .A1(n1308), .A2(n1309), .ZN(n1258) );
NAND2_X1 U987 ( .A1(G478), .A2(n1116), .ZN(n1309) );
XOR2_X1 U988 ( .A(KEYINPUT3), .B(n1310), .Z(n1308) );
NOR2_X1 U989 ( .A1(G478), .A2(n1116), .ZN(n1310) );
INV_X1 U990 ( .A(n1110), .ZN(n1116) );
NOR2_X1 U991 ( .A1(n1178), .A2(G902), .ZN(n1110) );
XNOR2_X1 U992 ( .A(n1311), .B(n1312), .ZN(n1178) );
XOR2_X1 U993 ( .A(n1313), .B(n1314), .Z(n1312) );
XOR2_X1 U994 ( .A(G128), .B(G122), .Z(n1314) );
XOR2_X1 U995 ( .A(KEYINPUT53), .B(G134), .Z(n1313) );
XOR2_X1 U996 ( .A(n1315), .B(n1316), .Z(n1311) );
XOR2_X1 U997 ( .A(G116), .B(G107), .Z(n1316) );
XOR2_X1 U998 ( .A(n1317), .B(n1307), .Z(n1315) );
NAND3_X1 U999 ( .A1(G217), .A2(n1082), .A3(G234), .ZN(n1317) );
INV_X1 U1000 ( .A(n1274), .ZN(n1186) );
NOR2_X1 U1001 ( .A1(n1239), .A2(n1241), .ZN(n1274) );
XNOR2_X1 U1002 ( .A(n1076), .B(KEYINPUT13), .ZN(n1241) );
NOR2_X1 U1003 ( .A1(n1079), .A2(n1106), .ZN(n1076) );
INV_X1 U1004 ( .A(n1080), .ZN(n1106) );
NAND2_X1 U1005 ( .A1(G221), .A2(n1318), .ZN(n1080) );
XNOR2_X1 U1006 ( .A(n1319), .B(n1320), .ZN(n1079) );
NOR2_X1 U1007 ( .A1(G469), .A2(KEYINPUT19), .ZN(n1320) );
XOR2_X1 U1008 ( .A(n1103), .B(KEYINPUT41), .Z(n1319) );
NAND2_X1 U1009 ( .A1(n1321), .A2(n1291), .ZN(n1103) );
XOR2_X1 U1010 ( .A(n1322), .B(n1323), .Z(n1321) );
XOR2_X1 U1011 ( .A(n1137), .B(n1205), .Z(n1323) );
XOR2_X1 U1012 ( .A(n1324), .B(n1325), .Z(n1137) );
XOR2_X1 U1013 ( .A(n1326), .B(G128), .Z(n1324) );
NAND2_X1 U1014 ( .A1(KEYINPUT63), .A2(n1307), .ZN(n1326) );
XNOR2_X1 U1015 ( .A(n1327), .B(n1328), .ZN(n1322) );
NOR2_X1 U1016 ( .A1(KEYINPUT0), .A2(n1214), .ZN(n1328) );
XOR2_X1 U1017 ( .A(n1329), .B(n1330), .Z(n1214) );
NOR2_X1 U1018 ( .A1(G953), .A2(n1148), .ZN(n1330) );
INV_X1 U1019 ( .A(G227), .ZN(n1148) );
NOR2_X1 U1020 ( .A1(KEYINPUT25), .A2(n1331), .ZN(n1327) );
XOR2_X1 U1021 ( .A(G101), .B(n1219), .Z(n1331) );
NAND4_X1 U1022 ( .A1(n1259), .A2(n1332), .A3(n1065), .A4(n1064), .ZN(n1239) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1333), .ZN(n1064) );
NAND2_X1 U1024 ( .A1(G237), .A2(G234), .ZN(n1065) );
NAND2_X1 U1025 ( .A1(n1334), .A2(n1278), .ZN(n1332) );
NAND2_X1 U1026 ( .A1(n1335), .A2(G952), .ZN(n1278) );
XOR2_X1 U1027 ( .A(n1082), .B(KEYINPUT16), .Z(n1335) );
NAND3_X1 U1028 ( .A1(G953), .A2(n1156), .A3(G902), .ZN(n1334) );
INV_X1 U1029 ( .A(G898), .ZN(n1156) );
INV_X1 U1030 ( .A(n1063), .ZN(n1259) );
XNOR2_X1 U1031 ( .A(n1336), .B(n1230), .ZN(n1063) );
NAND2_X1 U1032 ( .A1(G210), .A2(n1333), .ZN(n1230) );
NAND2_X1 U1033 ( .A1(n1306), .A2(n1291), .ZN(n1333) );
NAND2_X1 U1034 ( .A1(n1337), .A2(n1291), .ZN(n1336) );
XOR2_X1 U1035 ( .A(n1338), .B(n1339), .Z(n1337) );
XNOR2_X1 U1036 ( .A(n1228), .B(n1340), .ZN(n1339) );
NOR2_X1 U1037 ( .A1(KEYINPUT43), .A2(n1341), .ZN(n1340) );
XOR2_X1 U1038 ( .A(KEYINPUT34), .B(n1342), .Z(n1341) );
INV_X1 U1039 ( .A(n1225), .ZN(n1342) );
XOR2_X1 U1040 ( .A(n1343), .B(n1344), .Z(n1225) );
INV_X1 U1041 ( .A(n1157), .ZN(n1344) );
XOR2_X1 U1042 ( .A(n1345), .B(n1346), .Z(n1157) );
NOR2_X1 U1043 ( .A1(KEYINPUT62), .A2(n1289), .ZN(n1346) );
XNOR2_X1 U1044 ( .A(G122), .B(KEYINPUT9), .ZN(n1345) );
NAND2_X1 U1045 ( .A1(n1162), .A2(n1347), .ZN(n1343) );
OR2_X1 U1046 ( .A1(n1164), .A2(n1163), .ZN(n1347) );
NAND2_X1 U1047 ( .A1(n1163), .A2(n1164), .ZN(n1162) );
XNOR2_X1 U1048 ( .A(n1282), .B(n1348), .ZN(n1164) );
XNOR2_X1 U1049 ( .A(G101), .B(n1349), .ZN(n1163) );
NOR2_X1 U1050 ( .A1(KEYINPUT27), .A2(n1219), .ZN(n1349) );
XOR2_X1 U1051 ( .A(G104), .B(G107), .Z(n1219) );
NAND2_X1 U1052 ( .A1(G224), .A2(n1082), .ZN(n1228) );
NAND2_X1 U1053 ( .A1(KEYINPUT18), .A2(n1350), .ZN(n1338) );
XOR2_X1 U1054 ( .A(n1206), .B(G125), .Z(n1350) );
NAND2_X1 U1055 ( .A1(n1276), .A2(n1100), .ZN(n1266) );
XOR2_X1 U1056 ( .A(n1351), .B(n1171), .Z(n1100) );
NAND2_X1 U1057 ( .A1(G217), .A2(n1318), .ZN(n1171) );
NAND2_X1 U1058 ( .A1(G234), .A2(n1291), .ZN(n1318) );
NAND2_X1 U1059 ( .A1(n1173), .A2(n1291), .ZN(n1351) );
XOR2_X1 U1060 ( .A(n1352), .B(n1353), .Z(n1173) );
XOR2_X1 U1061 ( .A(n1354), .B(n1355), .Z(n1353) );
XOR2_X1 U1062 ( .A(G125), .B(G119), .Z(n1355) );
XOR2_X1 U1063 ( .A(KEYINPUT51), .B(G137), .Z(n1354) );
XOR2_X1 U1064 ( .A(n1356), .B(n1357), .Z(n1352) );
XOR2_X1 U1065 ( .A(n1358), .B(n1359), .Z(n1357) );
NAND2_X1 U1066 ( .A1(KEYINPUT60), .A2(n1269), .ZN(n1359) );
NAND3_X1 U1067 ( .A1(G234), .A2(n1082), .A3(G221), .ZN(n1358) );
XOR2_X1 U1068 ( .A(n1329), .B(n1360), .Z(n1356) );
NOR2_X1 U1069 ( .A1(KEYINPUT26), .A2(n1325), .ZN(n1360) );
XOR2_X1 U1070 ( .A(n1289), .B(n1136), .Z(n1329) );
XOR2_X1 U1071 ( .A(G140), .B(KEYINPUT4), .Z(n1136) );
INV_X1 U1072 ( .A(G110), .ZN(n1289) );
XNOR2_X1 U1073 ( .A(n1101), .B(KEYINPUT28), .ZN(n1276) );
XNOR2_X1 U1074 ( .A(n1361), .B(G472), .ZN(n1101) );
NAND2_X1 U1075 ( .A1(n1362), .A2(n1291), .ZN(n1361) );
INV_X1 U1076 ( .A(G902), .ZN(n1291) );
XOR2_X1 U1077 ( .A(n1363), .B(n1364), .Z(n1362) );
XNOR2_X1 U1078 ( .A(n1217), .B(n1200), .ZN(n1364) );
NAND2_X1 U1079 ( .A1(n1365), .A2(n1366), .ZN(n1200) );
NAND2_X1 U1080 ( .A1(n1367), .A2(n1282), .ZN(n1366) );
INV_X1 U1081 ( .A(G119), .ZN(n1282) );
XOR2_X1 U1082 ( .A(KEYINPUT1), .B(n1348), .Z(n1367) );
NAND2_X1 U1083 ( .A1(n1348), .A2(G119), .ZN(n1365) );
XOR2_X1 U1084 ( .A(G113), .B(G116), .Z(n1348) );
XOR2_X1 U1085 ( .A(n1205), .B(G101), .Z(n1217) );
XOR2_X1 U1086 ( .A(n1141), .B(n1140), .Z(n1205) );
XNOR2_X1 U1087 ( .A(G131), .B(G134), .ZN(n1140) );
INV_X1 U1088 ( .A(G137), .ZN(n1141) );
XOR2_X1 U1089 ( .A(n1206), .B(n1368), .Z(n1363) );
XNOR2_X1 U1090 ( .A(n1369), .B(KEYINPUT8), .ZN(n1368) );
NAND2_X1 U1091 ( .A1(KEYINPUT59), .A2(n1207), .ZN(n1369) );
AND3_X1 U1092 ( .A1(n1306), .A2(n1082), .A3(G210), .ZN(n1207) );
INV_X1 U1093 ( .A(G953), .ZN(n1082) );
INV_X1 U1094 ( .A(G237), .ZN(n1306) );
XOR2_X1 U1095 ( .A(n1269), .B(n1370), .Z(n1206) );
NOR2_X1 U1096 ( .A1(n1371), .A2(n1372), .ZN(n1370) );
NOR2_X1 U1097 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XOR2_X1 U1098 ( .A(KEYINPUT42), .B(n1325), .Z(n1374) );
NOR2_X1 U1099 ( .A1(n1307), .A2(n1375), .ZN(n1371) );
XOR2_X1 U1100 ( .A(KEYINPUT24), .B(n1325), .Z(n1375) );
INV_X1 U1101 ( .A(n1300), .ZN(n1325) );
XNOR2_X1 U1102 ( .A(G146), .B(KEYINPUT47), .ZN(n1300) );
INV_X1 U1103 ( .A(n1373), .ZN(n1307) );
XNOR2_X1 U1104 ( .A(G143), .B(KEYINPUT5), .ZN(n1373) );
INV_X1 U1105 ( .A(G128), .ZN(n1269) );
endmodule


