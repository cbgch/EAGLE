//Key = 0011011011000111010110010110100011001000100111001110010100111110


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340;

XNOR2_X1 U740 ( .A(G107), .B(n1028), .ZN(G9) );
NAND3_X1 U741 ( .A1(n1029), .A2(n1030), .A3(n1031), .ZN(n1028) );
XNOR2_X1 U742 ( .A(n1032), .B(KEYINPUT19), .ZN(n1031) );
NOR2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(G75) );
NOR3_X1 U744 ( .A1(n1035), .A2(G953), .A3(n1036), .ZN(n1034) );
INV_X1 U745 ( .A(n1037), .ZN(n1036) );
XNOR2_X1 U746 ( .A(G952), .B(KEYINPUT48), .ZN(n1035) );
NOR4_X1 U747 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1033) );
INV_X1 U748 ( .A(G952), .ZN(n1041) );
XOR2_X1 U749 ( .A(n1042), .B(KEYINPUT41), .Z(n1040) );
NAND2_X1 U750 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NAND3_X1 U751 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NAND3_X1 U752 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1046) );
NAND4_X1 U753 ( .A1(n1051), .A2(n1052), .A3(n1053), .A4(n1032), .ZN(n1050) );
NAND3_X1 U754 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1049) );
NAND3_X1 U755 ( .A1(n1053), .A2(n1057), .A3(n1058), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1059), .A2(n1030), .ZN(n1043) );
NAND4_X1 U757 ( .A1(n1037), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1038) );
NAND3_X1 U758 ( .A1(n1045), .A2(n1063), .A3(n1047), .ZN(n1061) );
NAND2_X1 U759 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NAND2_X1 U760 ( .A1(n1055), .A2(n1066), .ZN(n1065) );
NAND2_X1 U761 ( .A1(n1053), .A2(n1067), .ZN(n1064) );
NAND2_X1 U762 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
NAND2_X1 U763 ( .A1(n1070), .A2(n1032), .ZN(n1069) );
XNOR2_X1 U764 ( .A(n1071), .B(KEYINPUT60), .ZN(n1070) );
NAND2_X1 U765 ( .A1(n1072), .A2(n1073), .ZN(n1068) );
XNOR2_X1 U766 ( .A(n1058), .B(KEYINPUT59), .ZN(n1072) );
NAND2_X1 U767 ( .A1(n1059), .A2(n1074), .ZN(n1060) );
AND3_X1 U768 ( .A1(n1055), .A2(n1053), .A3(n1047), .ZN(n1059) );
INV_X1 U769 ( .A(n1075), .ZN(n1047) );
AND2_X1 U770 ( .A1(n1058), .A2(n1032), .ZN(n1055) );
NAND4_X1 U771 ( .A1(n1058), .A2(n1045), .A3(n1076), .A4(n1077), .ZN(n1037) );
NOR3_X1 U772 ( .A1(n1078), .A2(n1056), .A3(n1079), .ZN(n1077) );
XOR2_X1 U773 ( .A(n1080), .B(n1081), .Z(n1079) );
NOR2_X1 U774 ( .A1(G469), .A2(KEYINPUT30), .ZN(n1081) );
XNOR2_X1 U775 ( .A(n1082), .B(KEYINPUT56), .ZN(n1076) );
XOR2_X1 U776 ( .A(n1083), .B(n1084), .Z(G72) );
NOR2_X1 U777 ( .A1(n1085), .A2(n1062), .ZN(n1084) );
NOR2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U779 ( .A1(n1088), .A2(n1089), .ZN(n1083) );
NAND2_X1 U780 ( .A1(KEYINPUT46), .A2(n1090), .ZN(n1089) );
XOR2_X1 U781 ( .A(n1091), .B(n1092), .Z(n1088) );
NOR2_X1 U782 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
XOR2_X1 U783 ( .A(n1095), .B(n1096), .Z(n1094) );
XNOR2_X1 U784 ( .A(KEYINPUT45), .B(n1097), .ZN(n1096) );
XNOR2_X1 U785 ( .A(n1098), .B(n1099), .ZN(n1095) );
NAND2_X1 U786 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
OR2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U788 ( .A(n1104), .B(KEYINPUT52), .Z(n1100) );
NAND2_X1 U789 ( .A1(n1102), .A2(n1103), .ZN(n1104) );
XNOR2_X1 U790 ( .A(n1105), .B(G131), .ZN(n1102) );
NAND2_X1 U791 ( .A1(KEYINPUT61), .A2(n1106), .ZN(n1105) );
XNOR2_X1 U792 ( .A(n1107), .B(n1108), .ZN(n1106) );
NOR2_X1 U793 ( .A1(G900), .A2(n1109), .ZN(n1093) );
XNOR2_X1 U794 ( .A(KEYINPUT3), .B(n1062), .ZN(n1109) );
NOR2_X1 U795 ( .A1(n1090), .A2(KEYINPUT46), .ZN(n1091) );
AND2_X1 U796 ( .A1(n1062), .A2(n1110), .ZN(n1090) );
NAND2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
XNOR2_X1 U798 ( .A(KEYINPUT6), .B(n1113), .ZN(n1112) );
XOR2_X1 U799 ( .A(n1114), .B(n1115), .Z(G69) );
NOR2_X1 U800 ( .A1(n1116), .A2(n1062), .ZN(n1115) );
AND2_X1 U801 ( .A1(G224), .A2(G898), .ZN(n1116) );
NAND2_X1 U802 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NAND2_X1 U803 ( .A1(n1119), .A2(n1062), .ZN(n1118) );
XOR2_X1 U804 ( .A(n1120), .B(n1121), .Z(n1119) );
OR3_X1 U805 ( .A1(n1122), .A2(n1121), .A3(n1062), .ZN(n1117) );
XNOR2_X1 U806 ( .A(n1123), .B(n1124), .ZN(n1121) );
XNOR2_X1 U807 ( .A(n1125), .B(n1126), .ZN(n1123) );
NOR2_X1 U808 ( .A1(n1127), .A2(n1128), .ZN(G66) );
XOR2_X1 U809 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U810 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1133), .ZN(G63) );
XOR2_X1 U812 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U813 ( .A1(KEYINPUT54), .A2(n1136), .ZN(n1135) );
INV_X1 U814 ( .A(n1137), .ZN(n1136) );
NAND2_X1 U815 ( .A1(n1138), .A2(G478), .ZN(n1134) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1140), .ZN(G60) );
XNOR2_X1 U817 ( .A(n1127), .B(KEYINPUT8), .ZN(n1140) );
XNOR2_X1 U818 ( .A(n1141), .B(n1142), .ZN(n1139) );
AND2_X1 U819 ( .A1(G475), .A2(n1138), .ZN(n1142) );
XNOR2_X1 U820 ( .A(G104), .B(n1143), .ZN(G6) );
NAND2_X1 U821 ( .A1(KEYINPUT5), .A2(n1144), .ZN(n1143) );
INV_X1 U822 ( .A(n1145), .ZN(n1144) );
NOR2_X1 U823 ( .A1(n1127), .A2(n1146), .ZN(G57) );
XOR2_X1 U824 ( .A(n1147), .B(n1148), .Z(n1146) );
XNOR2_X1 U825 ( .A(n1126), .B(n1149), .ZN(n1148) );
XOR2_X1 U826 ( .A(n1150), .B(n1151), .Z(n1147) );
XOR2_X1 U827 ( .A(G101), .B(n1152), .Z(n1151) );
NOR3_X1 U828 ( .A1(n1132), .A2(KEYINPUT63), .A3(n1153), .ZN(n1150) );
NOR2_X1 U829 ( .A1(n1127), .A2(n1154), .ZN(G54) );
XOR2_X1 U830 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1156) );
XNOR2_X1 U832 ( .A(n1097), .B(G110), .ZN(n1158) );
AND2_X1 U833 ( .A1(G469), .A2(n1138), .ZN(n1157) );
INV_X1 U834 ( .A(n1132), .ZN(n1138) );
XNOR2_X1 U835 ( .A(n1159), .B(n1160), .ZN(n1155) );
NOR2_X1 U836 ( .A1(n1127), .A2(n1161), .ZN(G51) );
XOR2_X1 U837 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U838 ( .A(n1164), .B(n1165), .Z(n1162) );
NOR2_X1 U839 ( .A1(n1166), .A2(n1132), .ZN(n1165) );
NAND2_X1 U840 ( .A1(G902), .A2(n1039), .ZN(n1132) );
NAND3_X1 U841 ( .A1(n1111), .A2(n1113), .A3(n1120), .ZN(n1039) );
AND4_X1 U842 ( .A1(n1145), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1120) );
NOR4_X1 U843 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169) );
NOR2_X1 U844 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
AND3_X1 U845 ( .A1(n1029), .A2(n1032), .A3(n1030), .ZN(n1171) );
NOR2_X1 U846 ( .A1(n1176), .A2(n1177), .ZN(n1168) );
NAND3_X1 U847 ( .A1(n1029), .A2(n1032), .A3(n1074), .ZN(n1145) );
NAND3_X1 U848 ( .A1(n1178), .A2(n1071), .A3(n1179), .ZN(n1113) );
XNOR2_X1 U849 ( .A(n1053), .B(KEYINPUT36), .ZN(n1179) );
AND4_X1 U850 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1111) );
NOR4_X1 U851 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
INV_X1 U852 ( .A(n1188), .ZN(n1185) );
OR2_X1 U853 ( .A1(n1189), .A2(n1190), .ZN(n1182) );
NAND2_X1 U854 ( .A1(n1058), .A2(n1191), .ZN(n1181) );
NAND2_X1 U855 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NAND2_X1 U856 ( .A1(n1194), .A2(n1074), .ZN(n1193) );
NAND2_X1 U857 ( .A1(n1195), .A2(n1196), .ZN(n1192) );
NAND2_X1 U858 ( .A1(n1197), .A2(n1198), .ZN(n1195) );
NAND4_X1 U859 ( .A1(n1199), .A2(n1045), .A3(n1200), .A4(n1189), .ZN(n1198) );
INV_X1 U860 ( .A(KEYINPUT25), .ZN(n1189) );
NAND2_X1 U861 ( .A1(KEYINPUT7), .A2(n1178), .ZN(n1197) );
NAND2_X1 U862 ( .A1(n1201), .A2(n1202), .ZN(n1180) );
INV_X1 U863 ( .A(KEYINPUT7), .ZN(n1202) );
NAND2_X1 U864 ( .A1(KEYINPUT26), .A2(n1099), .ZN(n1164) );
NOR2_X1 U865 ( .A1(n1062), .A2(G952), .ZN(n1127) );
XOR2_X1 U866 ( .A(n1203), .B(n1187), .Z(G48) );
AND3_X1 U867 ( .A1(n1074), .A2(n1071), .A3(n1204), .ZN(n1187) );
XNOR2_X1 U868 ( .A(G146), .B(KEYINPUT55), .ZN(n1203) );
XOR2_X1 U869 ( .A(n1205), .B(n1186), .Z(G45) );
AND4_X1 U870 ( .A1(n1194), .A2(n1071), .A3(n1206), .A4(n1207), .ZN(n1186) );
NAND2_X1 U871 ( .A1(KEYINPUT14), .A2(n1208), .ZN(n1205) );
XOR2_X1 U872 ( .A(n1209), .B(n1201), .Z(G42) );
NOR3_X1 U873 ( .A1(n1210), .A2(n1196), .A3(n1211), .ZN(n1201) );
NAND2_X1 U874 ( .A1(KEYINPUT43), .A2(n1097), .ZN(n1209) );
INV_X1 U875 ( .A(G140), .ZN(n1097) );
XOR2_X1 U876 ( .A(n1190), .B(n1212), .Z(G39) );
XNOR2_X1 U877 ( .A(G137), .B(KEYINPUT27), .ZN(n1212) );
NAND3_X1 U878 ( .A1(n1204), .A2(n1045), .A3(n1058), .ZN(n1190) );
XNOR2_X1 U879 ( .A(G134), .B(n1188), .ZN(G36) );
NAND3_X1 U880 ( .A1(n1058), .A2(n1030), .A3(n1194), .ZN(n1188) );
AND3_X1 U881 ( .A1(n1066), .A2(n1200), .A3(n1073), .ZN(n1194) );
INV_X1 U882 ( .A(n1210), .ZN(n1058) );
XOR2_X1 U883 ( .A(G131), .B(n1213), .Z(G33) );
NOR3_X1 U884 ( .A1(n1214), .A2(n1210), .A3(n1215), .ZN(n1213) );
XNOR2_X1 U885 ( .A(KEYINPUT2), .B(n1196), .ZN(n1215) );
INV_X1 U886 ( .A(n1066), .ZN(n1196) );
NAND2_X1 U887 ( .A1(n1051), .A2(n1216), .ZN(n1210) );
NAND3_X1 U888 ( .A1(n1073), .A2(n1200), .A3(n1074), .ZN(n1214) );
XNOR2_X1 U889 ( .A(n1217), .B(n1184), .ZN(G30) );
AND3_X1 U890 ( .A1(n1030), .A2(n1071), .A3(n1204), .ZN(n1184) );
AND3_X1 U891 ( .A1(n1066), .A2(n1200), .A3(n1199), .ZN(n1204) );
XOR2_X1 U892 ( .A(G101), .B(n1172), .Z(G3) );
AND3_X1 U893 ( .A1(n1045), .A2(n1029), .A3(n1073), .ZN(n1172) );
XNOR2_X1 U894 ( .A(G125), .B(n1218), .ZN(G27) );
NAND2_X1 U895 ( .A1(n1071), .A2(n1219), .ZN(n1218) );
XOR2_X1 U896 ( .A(KEYINPUT22), .B(n1220), .Z(n1219) );
AND2_X1 U897 ( .A1(n1053), .A2(n1178), .ZN(n1220) );
INV_X1 U898 ( .A(n1211), .ZN(n1178) );
NAND3_X1 U899 ( .A1(n1057), .A2(n1200), .A3(n1074), .ZN(n1211) );
NAND2_X1 U900 ( .A1(n1075), .A2(n1221), .ZN(n1200) );
NAND4_X1 U901 ( .A1(G953), .A2(n1222), .A3(n1223), .A4(n1087), .ZN(n1221) );
INV_X1 U902 ( .A(G900), .ZN(n1087) );
XNOR2_X1 U903 ( .A(KEYINPUT51), .B(n1224), .ZN(n1222) );
XNOR2_X1 U904 ( .A(G122), .B(n1167), .ZN(G24) );
NAND4_X1 U905 ( .A1(n1225), .A2(n1032), .A3(n1206), .A4(n1207), .ZN(n1167) );
NOR2_X1 U906 ( .A1(n1078), .A2(n1082), .ZN(n1032) );
XNOR2_X1 U907 ( .A(n1226), .B(n1227), .ZN(G21) );
NOR2_X1 U908 ( .A1(n1228), .A2(n1174), .ZN(n1227) );
XOR2_X1 U909 ( .A(n1175), .B(KEYINPUT1), .Z(n1228) );
NAND3_X1 U910 ( .A1(n1229), .A2(n1045), .A3(n1199), .ZN(n1175) );
AND2_X1 U911 ( .A1(n1082), .A2(n1078), .ZN(n1199) );
XOR2_X1 U912 ( .A(n1230), .B(n1231), .Z(G18) );
NOR2_X1 U913 ( .A1(KEYINPUT11), .A2(n1232), .ZN(n1231) );
INV_X1 U914 ( .A(G116), .ZN(n1232) );
NAND2_X1 U915 ( .A1(n1233), .A2(n1234), .ZN(n1230) );
NAND4_X1 U916 ( .A1(n1030), .A2(n1174), .A3(n1235), .A4(n1236), .ZN(n1234) );
INV_X1 U917 ( .A(KEYINPUT44), .ZN(n1236) );
AND2_X1 U918 ( .A1(n1229), .A2(n1073), .ZN(n1235) );
INV_X1 U919 ( .A(n1237), .ZN(n1229) );
NAND2_X1 U920 ( .A1(n1170), .A2(KEYINPUT44), .ZN(n1233) );
AND3_X1 U921 ( .A1(n1225), .A2(n1030), .A3(n1073), .ZN(n1170) );
NOR2_X1 U922 ( .A1(n1207), .A2(n1238), .ZN(n1030) );
XOR2_X1 U923 ( .A(G113), .B(n1177), .Z(G15) );
AND3_X1 U924 ( .A1(n1073), .A2(n1225), .A3(n1074), .ZN(n1177) );
AND2_X1 U925 ( .A1(n1238), .A2(n1207), .ZN(n1074) );
INV_X1 U926 ( .A(n1206), .ZN(n1238) );
NOR2_X1 U927 ( .A1(n1237), .A2(n1174), .ZN(n1225) );
INV_X1 U928 ( .A(n1071), .ZN(n1174) );
NAND2_X1 U929 ( .A1(n1053), .A2(n1239), .ZN(n1237) );
NOR2_X1 U930 ( .A1(n1240), .A2(n1056), .ZN(n1053) );
NOR2_X1 U931 ( .A1(n1082), .A2(n1241), .ZN(n1073) );
XOR2_X1 U932 ( .A(n1176), .B(n1242), .Z(G12) );
NOR2_X1 U933 ( .A1(KEYINPUT21), .A2(n1243), .ZN(n1242) );
AND3_X1 U934 ( .A1(n1057), .A2(n1029), .A3(n1045), .ZN(n1176) );
NOR2_X1 U935 ( .A1(n1206), .A2(n1207), .ZN(n1045) );
XNOR2_X1 U936 ( .A(n1244), .B(G475), .ZN(n1207) );
NAND2_X1 U937 ( .A1(n1141), .A2(n1224), .ZN(n1244) );
XNOR2_X1 U938 ( .A(n1245), .B(n1246), .ZN(n1141) );
XOR2_X1 U939 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U940 ( .A(n1249), .B(n1250), .Z(n1248) );
AND2_X1 U941 ( .A1(G214), .A2(n1251), .ZN(n1250) );
NAND2_X1 U942 ( .A1(KEYINPUT13), .A2(n1252), .ZN(n1249) );
XOR2_X1 U943 ( .A(n1253), .B(n1254), .Z(n1252) );
XNOR2_X1 U944 ( .A(n1255), .B(G125), .ZN(n1254) );
NOR2_X1 U945 ( .A1(G140), .A2(KEYINPUT24), .ZN(n1253) );
XNOR2_X1 U946 ( .A(G104), .B(G113), .ZN(n1247) );
XOR2_X1 U947 ( .A(n1256), .B(n1257), .Z(n1245) );
XNOR2_X1 U948 ( .A(KEYINPUT53), .B(n1208), .ZN(n1257) );
XNOR2_X1 U949 ( .A(G122), .B(G131), .ZN(n1256) );
XNOR2_X1 U950 ( .A(n1258), .B(G478), .ZN(n1206) );
NAND2_X1 U951 ( .A1(n1259), .A2(n1137), .ZN(n1258) );
XNOR2_X1 U952 ( .A(n1260), .B(n1261), .ZN(n1137) );
NOR2_X1 U953 ( .A1(n1262), .A2(n1131), .ZN(n1261) );
NAND2_X1 U954 ( .A1(n1263), .A2(KEYINPUT49), .ZN(n1260) );
XOR2_X1 U955 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U956 ( .A(n1266), .B(n1267), .ZN(n1265) );
XNOR2_X1 U957 ( .A(KEYINPUT62), .B(n1107), .ZN(n1267) );
INV_X1 U958 ( .A(G122), .ZN(n1266) );
XOR2_X1 U959 ( .A(n1268), .B(n1269), .Z(n1264) );
NOR2_X1 U960 ( .A1(KEYINPUT39), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U961 ( .A(G128), .B(n1271), .ZN(n1270) );
NAND2_X1 U962 ( .A1(n1272), .A2(n1208), .ZN(n1271) );
XNOR2_X1 U963 ( .A(KEYINPUT18), .B(KEYINPUT12), .ZN(n1272) );
XNOR2_X1 U964 ( .A(G116), .B(G107), .ZN(n1268) );
XNOR2_X1 U965 ( .A(KEYINPUT28), .B(n1224), .ZN(n1259) );
AND3_X1 U966 ( .A1(n1071), .A2(n1239), .A3(n1066), .ZN(n1029) );
NOR2_X1 U967 ( .A1(n1054), .A2(n1056), .ZN(n1066) );
AND2_X1 U968 ( .A1(G221), .A2(n1273), .ZN(n1056) );
INV_X1 U969 ( .A(n1240), .ZN(n1054) );
XNOR2_X1 U970 ( .A(n1080), .B(G469), .ZN(n1240) );
NAND2_X1 U971 ( .A1(n1274), .A2(n1224), .ZN(n1080) );
XOR2_X1 U972 ( .A(n1160), .B(n1275), .Z(n1274) );
XNOR2_X1 U973 ( .A(n1276), .B(n1277), .ZN(n1275) );
NOR2_X1 U974 ( .A1(KEYINPUT47), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U975 ( .A(n1243), .B(n1279), .ZN(n1278) );
NOR2_X1 U976 ( .A1(G140), .A2(KEYINPUT38), .ZN(n1279) );
NAND2_X1 U977 ( .A1(KEYINPUT23), .A2(n1280), .ZN(n1276) );
XNOR2_X1 U978 ( .A(KEYINPUT29), .B(n1281), .ZN(n1280) );
INV_X1 U979 ( .A(n1159), .ZN(n1281) );
XNOR2_X1 U980 ( .A(n1282), .B(n1283), .ZN(n1159) );
XOR2_X1 U981 ( .A(n1284), .B(n1103), .Z(n1283) );
XNOR2_X1 U982 ( .A(G128), .B(n1285), .ZN(n1103) );
XOR2_X1 U983 ( .A(n1286), .B(n1287), .Z(n1282) );
NOR2_X1 U984 ( .A1(G107), .A2(KEYINPUT31), .ZN(n1287) );
NOR2_X1 U985 ( .A1(n1086), .A2(G953), .ZN(n1160) );
INV_X1 U986 ( .A(G227), .ZN(n1086) );
NAND2_X1 U987 ( .A1(n1075), .A2(n1288), .ZN(n1239) );
NAND4_X1 U988 ( .A1(G953), .A2(G902), .A3(n1223), .A4(n1122), .ZN(n1288) );
INV_X1 U989 ( .A(G898), .ZN(n1122) );
NAND3_X1 U990 ( .A1(n1223), .A2(n1062), .A3(G952), .ZN(n1075) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1223) );
NOR2_X1 U992 ( .A1(n1051), .A2(n1052), .ZN(n1071) );
INV_X1 U993 ( .A(n1216), .ZN(n1052) );
NAND2_X1 U994 ( .A1(G214), .A2(n1289), .ZN(n1216) );
XNOR2_X1 U995 ( .A(n1290), .B(n1166), .ZN(n1051) );
NAND2_X1 U996 ( .A1(G210), .A2(n1289), .ZN(n1166) );
NAND2_X1 U997 ( .A1(n1291), .A2(n1224), .ZN(n1289) );
INV_X1 U998 ( .A(G237), .ZN(n1291) );
NAND2_X1 U999 ( .A1(n1292), .A2(n1224), .ZN(n1290) );
XOR2_X1 U1000 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U1001 ( .A(n1099), .B(n1163), .ZN(n1294) );
XNOR2_X1 U1002 ( .A(n1295), .B(n1296), .ZN(n1163) );
XOR2_X1 U1003 ( .A(n1297), .B(n1124), .Z(n1296) );
XNOR2_X1 U1004 ( .A(n1243), .B(G122), .ZN(n1124) );
INV_X1 U1005 ( .A(G110), .ZN(n1243) );
XOR2_X1 U1006 ( .A(n1298), .B(n1299), .Z(n1295) );
NOR2_X1 U1007 ( .A1(KEYINPUT10), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1008 ( .A(n1125), .B(n1301), .Z(n1300) );
XNOR2_X1 U1009 ( .A(n1302), .B(KEYINPUT42), .ZN(n1301) );
NAND2_X1 U1010 ( .A1(KEYINPUT17), .A2(n1126), .ZN(n1302) );
XNOR2_X1 U1011 ( .A(G107), .B(n1284), .ZN(n1125) );
XOR2_X1 U1012 ( .A(G104), .B(G101), .Z(n1284) );
NAND2_X1 U1013 ( .A1(G224), .A2(n1062), .ZN(n1298) );
INV_X1 U1014 ( .A(G125), .ZN(n1099) );
XOR2_X1 U1015 ( .A(KEYINPUT40), .B(KEYINPUT16), .Z(n1293) );
AND2_X1 U1016 ( .A1(n1241), .A2(n1082), .ZN(n1057) );
XNOR2_X1 U1017 ( .A(n1303), .B(n1304), .ZN(n1082) );
NOR2_X1 U1018 ( .A1(n1131), .A2(n1305), .ZN(n1304) );
XNOR2_X1 U1019 ( .A(KEYINPUT35), .B(n1273), .ZN(n1305) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1224), .ZN(n1273) );
INV_X1 U1021 ( .A(G217), .ZN(n1131) );
OR2_X1 U1022 ( .A1(n1130), .A2(G902), .ZN(n1303) );
XNOR2_X1 U1023 ( .A(n1306), .B(n1307), .ZN(n1130) );
XOR2_X1 U1024 ( .A(n1308), .B(n1309), .Z(n1307) );
NAND2_X1 U1025 ( .A1(n1310), .A2(KEYINPUT50), .ZN(n1309) );
XNOR2_X1 U1026 ( .A(n1108), .B(KEYINPUT33), .ZN(n1310) );
NAND3_X1 U1027 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1308) );
OR2_X1 U1028 ( .A1(n1314), .A2(KEYINPUT15), .ZN(n1313) );
NAND3_X1 U1029 ( .A1(KEYINPUT15), .A2(n1314), .A3(n1315), .ZN(n1312) );
NAND2_X1 U1030 ( .A1(n1316), .A2(n1317), .ZN(n1311) );
NAND2_X1 U1031 ( .A1(n1318), .A2(KEYINPUT15), .ZN(n1317) );
XOR2_X1 U1032 ( .A(KEYINPUT57), .B(n1314), .Z(n1318) );
XNOR2_X1 U1033 ( .A(n1255), .B(n1319), .ZN(n1314) );
NOR2_X1 U1034 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NOR2_X1 U1035 ( .A1(G140), .A2(n1322), .ZN(n1321) );
XOR2_X1 U1036 ( .A(KEYINPUT37), .B(n1323), .Z(n1322) );
AND2_X1 U1037 ( .A1(G140), .A2(n1323), .ZN(n1320) );
XOR2_X1 U1038 ( .A(G125), .B(KEYINPUT4), .Z(n1323) );
INV_X1 U1039 ( .A(n1315), .ZN(n1316) );
XNOR2_X1 U1040 ( .A(n1324), .B(n1325), .ZN(n1315) );
XNOR2_X1 U1041 ( .A(KEYINPUT32), .B(n1217), .ZN(n1325) );
XNOR2_X1 U1042 ( .A(G119), .B(G110), .ZN(n1324) );
NAND2_X1 U1043 ( .A1(n1326), .A2(G221), .ZN(n1306) );
INV_X1 U1044 ( .A(n1262), .ZN(n1326) );
NAND2_X1 U1045 ( .A1(G234), .A2(n1062), .ZN(n1262) );
INV_X1 U1046 ( .A(G953), .ZN(n1062) );
INV_X1 U1047 ( .A(n1078), .ZN(n1241) );
XOR2_X1 U1048 ( .A(n1327), .B(n1153), .Z(n1078) );
INV_X1 U1049 ( .A(G472), .ZN(n1153) );
NAND2_X1 U1050 ( .A1(n1328), .A2(n1224), .ZN(n1327) );
INV_X1 U1051 ( .A(G902), .ZN(n1224) );
XOR2_X1 U1052 ( .A(n1329), .B(n1330), .Z(n1328) );
XNOR2_X1 U1053 ( .A(G101), .B(n1331), .ZN(n1330) );
NAND2_X1 U1054 ( .A1(KEYINPUT20), .A2(n1152), .ZN(n1331) );
AND2_X1 U1055 ( .A1(n1251), .A2(G210), .ZN(n1152) );
NOR2_X1 U1056 ( .A1(G953), .A2(G237), .ZN(n1251) );
XNOR2_X1 U1057 ( .A(n1332), .B(n1126), .ZN(n1329) );
XNOR2_X1 U1058 ( .A(G113), .B(n1333), .ZN(n1126) );
XNOR2_X1 U1059 ( .A(n1226), .B(G116), .ZN(n1333) );
INV_X1 U1060 ( .A(G119), .ZN(n1226) );
NAND2_X1 U1061 ( .A1(n1334), .A2(n1335), .ZN(n1332) );
OR2_X1 U1062 ( .A1(n1336), .A2(n1149), .ZN(n1335) );
XNOR2_X1 U1063 ( .A(n1286), .B(n1297), .ZN(n1149) );
NAND3_X1 U1064 ( .A1(n1297), .A2(n1286), .A3(n1336), .ZN(n1334) );
INV_X1 U1065 ( .A(KEYINPUT9), .ZN(n1336) );
XNOR2_X1 U1066 ( .A(n1337), .B(n1338), .ZN(n1286) );
INV_X1 U1067 ( .A(n1108), .ZN(n1338) );
XOR2_X1 U1068 ( .A(G137), .B(KEYINPUT0), .Z(n1108) );
XOR2_X1 U1069 ( .A(n1339), .B(G131), .Z(n1337) );
NAND2_X1 U1070 ( .A1(KEYINPUT58), .A2(n1107), .ZN(n1339) );
INV_X1 U1071 ( .A(G134), .ZN(n1107) );
XNOR2_X1 U1072 ( .A(n1217), .B(n1340), .ZN(n1297) );
NOR2_X1 U1073 ( .A1(KEYINPUT34), .A2(n1285), .ZN(n1340) );
XNOR2_X1 U1074 ( .A(n1208), .B(n1255), .ZN(n1285) );
INV_X1 U1075 ( .A(G146), .ZN(n1255) );
INV_X1 U1076 ( .A(G143), .ZN(n1208) );
INV_X1 U1077 ( .A(G128), .ZN(n1217) );
endmodule


