//Key = 0010111110010110010001001111010100000100011101000011110110110001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317;

XOR2_X1 U728 ( .A(n1007), .B(n1008), .Z(G9) );
NAND4_X1 U729 ( .A1(KEYINPUT45), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1008) );
NOR2_X1 U730 ( .A1(n1012), .A2(n1013), .ZN(G75) );
NOR4_X1 U731 ( .A1(n1014), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1013) );
INV_X1 U732 ( .A(G952), .ZN(n1017) );
NOR2_X1 U733 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
INV_X1 U734 ( .A(n1020), .ZN(n1018) );
NAND3_X1 U735 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n1014) );
NAND3_X1 U736 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1023) );
NAND2_X1 U737 ( .A1(n1027), .A2(n1028), .ZN(n1025) );
NAND2_X1 U738 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
NAND2_X1 U739 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND3_X1 U740 ( .A1(n1011), .A2(n1033), .A3(n1034), .ZN(n1032) );
NAND2_X1 U741 ( .A1(n1035), .A2(n1036), .ZN(n1033) );
NAND2_X1 U742 ( .A1(n1037), .A2(n1038), .ZN(n1031) );
NAND2_X1 U743 ( .A1(n1039), .A2(n1040), .ZN(n1038) );
NAND2_X1 U744 ( .A1(n1011), .A2(n1041), .ZN(n1040) );
NAND2_X1 U745 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND2_X1 U746 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
INV_X1 U747 ( .A(n1046), .ZN(n1042) );
NAND2_X1 U748 ( .A1(n1034), .A2(n1047), .ZN(n1039) );
NAND2_X1 U749 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NAND2_X1 U750 ( .A1(n1050), .A2(n1051), .ZN(n1024) );
XOR2_X1 U751 ( .A(n1019), .B(KEYINPUT44), .Z(n1051) );
NAND4_X1 U752 ( .A1(n1029), .A2(n1034), .A3(n1037), .A4(n1011), .ZN(n1019) );
INV_X1 U753 ( .A(n1052), .ZN(n1029) );
NOR3_X1 U754 ( .A1(n1053), .A2(G953), .A3(n1054), .ZN(n1012) );
INV_X1 U755 ( .A(n1021), .ZN(n1054) );
NAND4_X1 U756 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1021) );
NOR4_X1 U757 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1058) );
XOR2_X1 U758 ( .A(KEYINPUT61), .B(n1063), .Z(n1062) );
NOR2_X1 U759 ( .A1(G472), .A2(n1064), .ZN(n1063) );
INV_X1 U760 ( .A(n1037), .ZN(n1061) );
XOR2_X1 U761 ( .A(n1045), .B(KEYINPUT14), .Z(n1060) );
XOR2_X1 U762 ( .A(n1065), .B(n1066), .Z(n1059) );
XNOR2_X1 U763 ( .A(KEYINPUT37), .B(n1067), .ZN(n1066) );
NAND2_X1 U764 ( .A1(KEYINPUT43), .A2(n1068), .ZN(n1065) );
XNOR2_X1 U765 ( .A(KEYINPUT10), .B(n1069), .ZN(n1068) );
NOR3_X1 U766 ( .A1(n1050), .A2(n1044), .A3(n1070), .ZN(n1057) );
NAND2_X1 U767 ( .A1(G472), .A2(n1064), .ZN(n1055) );
XOR2_X1 U768 ( .A(n1071), .B(G952), .Z(n1053) );
XNOR2_X1 U769 ( .A(KEYINPUT7), .B(KEYINPUT62), .ZN(n1071) );
XOR2_X1 U770 ( .A(n1072), .B(n1073), .Z(G72) );
XOR2_X1 U771 ( .A(n1074), .B(n1075), .Z(n1073) );
NOR2_X1 U772 ( .A1(G953), .A2(n1076), .ZN(n1075) );
NOR2_X1 U773 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U774 ( .A(KEYINPUT18), .B(n1079), .Z(n1078) );
NOR2_X1 U775 ( .A1(KEYINPUT35), .A2(n1080), .ZN(n1074) );
NOR2_X1 U776 ( .A1(n1081), .A2(n1022), .ZN(n1080) );
NOR2_X1 U777 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NAND2_X1 U778 ( .A1(n1084), .A2(n1085), .ZN(n1072) );
NAND2_X1 U779 ( .A1(G953), .A2(n1083), .ZN(n1085) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1084) );
XOR2_X1 U781 ( .A(n1088), .B(n1089), .Z(n1087) );
XOR2_X1 U782 ( .A(n1090), .B(n1091), .Z(n1086) );
NOR2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XOR2_X1 U784 ( .A(n1094), .B(KEYINPUT24), .Z(n1093) );
NAND2_X1 U785 ( .A1(G134), .A2(n1095), .ZN(n1094) );
NOR2_X1 U786 ( .A1(G134), .A2(n1095), .ZN(n1092) );
INV_X1 U787 ( .A(G137), .ZN(n1095) );
NOR2_X1 U788 ( .A1(KEYINPUT15), .A2(G125), .ZN(n1090) );
NAND2_X1 U789 ( .A1(n1096), .A2(n1097), .ZN(G69) );
NAND2_X1 U790 ( .A1(n1098), .A2(n1022), .ZN(n1097) );
XOR2_X1 U791 ( .A(n1099), .B(n1100), .Z(n1098) );
NAND2_X1 U792 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
XOR2_X1 U793 ( .A(n1103), .B(KEYINPUT41), .Z(n1101) );
NAND2_X1 U794 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U795 ( .A1(n1106), .A2(G953), .ZN(n1096) );
XOR2_X1 U796 ( .A(n1100), .B(n1107), .Z(n1106) );
NAND2_X1 U797 ( .A1(G898), .A2(G224), .ZN(n1107) );
NAND2_X1 U798 ( .A1(KEYINPUT56), .A2(n1108), .ZN(n1100) );
NAND2_X1 U799 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U800 ( .A1(G953), .A2(n1111), .ZN(n1110) );
XOR2_X1 U801 ( .A(n1112), .B(n1113), .Z(n1109) );
XNOR2_X1 U802 ( .A(n1114), .B(KEYINPUT8), .ZN(n1112) );
NOR2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XOR2_X1 U804 ( .A(n1117), .B(n1118), .Z(n1116) );
NOR2_X1 U805 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
NOR2_X1 U806 ( .A1(n1115), .A2(n1121), .ZN(G63) );
XOR2_X1 U807 ( .A(n1122), .B(n1123), .Z(n1121) );
AND2_X1 U808 ( .A1(G478), .A2(n1124), .ZN(n1122) );
NOR2_X1 U809 ( .A1(n1115), .A2(n1125), .ZN(G60) );
XOR2_X1 U810 ( .A(n1126), .B(n1127), .Z(n1125) );
NAND2_X1 U811 ( .A1(n1124), .A2(n1128), .ZN(n1126) );
XOR2_X1 U812 ( .A(KEYINPUT54), .B(G475), .Z(n1128) );
XOR2_X1 U813 ( .A(n1129), .B(n1130), .Z(G6) );
NOR2_X1 U814 ( .A1(n1131), .A2(n1132), .ZN(G57) );
XOR2_X1 U815 ( .A(n1133), .B(n1134), .Z(n1132) );
XNOR2_X1 U816 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U817 ( .A(n1137), .B(n1138), .Z(n1133) );
NOR2_X1 U818 ( .A1(KEYINPUT49), .A2(n1139), .ZN(n1138) );
XOR2_X1 U819 ( .A(n1140), .B(n1141), .Z(n1139) );
NAND2_X1 U820 ( .A1(KEYINPUT25), .A2(n1142), .ZN(n1140) );
XNOR2_X1 U821 ( .A(KEYINPUT36), .B(n1143), .ZN(n1142) );
NAND2_X1 U822 ( .A1(n1124), .A2(G472), .ZN(n1137) );
NOR2_X1 U823 ( .A1(G952), .A2(n1144), .ZN(n1131) );
XOR2_X1 U824 ( .A(n1022), .B(KEYINPUT9), .Z(n1144) );
NOR2_X1 U825 ( .A1(n1115), .A2(n1145), .ZN(G54) );
XOR2_X1 U826 ( .A(n1146), .B(n1147), .Z(n1145) );
XOR2_X1 U827 ( .A(n1148), .B(n1149), .Z(n1146) );
NOR2_X1 U828 ( .A1(KEYINPUT47), .A2(n1143), .ZN(n1149) );
NAND2_X1 U829 ( .A1(n1124), .A2(G469), .ZN(n1148) );
INV_X1 U830 ( .A(n1120), .ZN(n1124) );
NOR2_X1 U831 ( .A1(n1115), .A2(n1150), .ZN(G51) );
XOR2_X1 U832 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U833 ( .A1(n1069), .A2(n1120), .ZN(n1152) );
NAND2_X1 U834 ( .A1(G902), .A2(n1015), .ZN(n1120) );
NAND4_X1 U835 ( .A1(n1153), .A2(n1102), .A3(n1154), .A4(n1104), .ZN(n1015) );
AND3_X1 U836 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1104) );
NOR2_X1 U837 ( .A1(n1079), .A2(n1158), .ZN(n1154) );
XOR2_X1 U838 ( .A(n1105), .B(KEYINPUT26), .Z(n1158) );
AND4_X1 U839 ( .A1(n1159), .A2(n1130), .A3(n1160), .A4(n1161), .ZN(n1102) );
NAND3_X1 U840 ( .A1(n1009), .A2(n1011), .A3(n1162), .ZN(n1130) );
NAND3_X1 U841 ( .A1(n1010), .A2(n1011), .A3(n1009), .ZN(n1159) );
INV_X1 U842 ( .A(n1077), .ZN(n1153) );
NAND4_X1 U843 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1077) );
NOR4_X1 U844 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1166) );
INV_X1 U845 ( .A(n1171), .ZN(n1168) );
INV_X1 U846 ( .A(n1172), .ZN(n1167) );
NAND3_X1 U847 ( .A1(n1173), .A2(n1010), .A3(n1174), .ZN(n1165) );
XOR2_X1 U848 ( .A(n1048), .B(KEYINPUT6), .Z(n1174) );
NOR3_X1 U849 ( .A1(n1175), .A2(KEYINPUT22), .A3(n1176), .ZN(n1151) );
NOR2_X1 U850 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U851 ( .A(KEYINPUT2), .B(n1179), .Z(n1178) );
INV_X1 U852 ( .A(n1180), .ZN(n1177) );
XOR2_X1 U853 ( .A(KEYINPUT12), .B(n1181), .Z(n1175) );
NOR2_X1 U854 ( .A1(n1180), .A2(n1179), .ZN(n1181) );
XOR2_X1 U855 ( .A(n1182), .B(n1141), .Z(n1179) );
XOR2_X1 U856 ( .A(n1183), .B(n1184), .Z(n1182) );
NOR2_X1 U857 ( .A1(n1022), .A2(G952), .ZN(n1115) );
NAND2_X1 U858 ( .A1(n1185), .A2(n1186), .ZN(G48) );
NAND2_X1 U859 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
XOR2_X1 U860 ( .A(KEYINPUT17), .B(G146), .Z(n1188) );
XOR2_X1 U861 ( .A(KEYINPUT63), .B(n1189), .Z(n1185) );
NOR2_X1 U862 ( .A1(n1187), .A2(n1190), .ZN(n1189) );
XOR2_X1 U863 ( .A(n1191), .B(KEYINPUT20), .Z(n1190) );
INV_X1 U864 ( .A(n1163), .ZN(n1187) );
NAND3_X1 U865 ( .A1(n1192), .A2(n1162), .A3(n1193), .ZN(n1163) );
XOR2_X1 U866 ( .A(n1164), .B(n1194), .Z(G45) );
NOR2_X1 U867 ( .A1(G143), .A2(KEYINPUT40), .ZN(n1194) );
NAND3_X1 U868 ( .A1(n1192), .A2(n1195), .A3(n1196), .ZN(n1164) );
XOR2_X1 U869 ( .A(G140), .B(n1170), .Z(G42) );
NOR3_X1 U870 ( .A1(n1035), .A2(n1197), .A3(n1049), .ZN(n1170) );
XOR2_X1 U871 ( .A(G137), .B(n1169), .Z(G39) );
AND2_X1 U872 ( .A1(n1198), .A2(n1173), .ZN(n1169) );
INV_X1 U873 ( .A(n1197), .ZN(n1173) );
XOR2_X1 U874 ( .A(G134), .B(n1199), .Z(G36) );
NOR3_X1 U875 ( .A1(n1048), .A2(n1036), .A3(n1197), .ZN(n1199) );
INV_X1 U876 ( .A(n1010), .ZN(n1036) );
XOR2_X1 U877 ( .A(G131), .B(n1079), .Z(G33) );
NOR3_X1 U878 ( .A1(n1035), .A2(n1197), .A3(n1048), .ZN(n1079) );
INV_X1 U879 ( .A(n1195), .ZN(n1048) );
NAND4_X1 U880 ( .A1(n1026), .A2(n1046), .A3(n1200), .A4(n1028), .ZN(n1197) );
XOR2_X1 U881 ( .A(n1201), .B(n1171), .Z(G30) );
NAND3_X1 U882 ( .A1(n1192), .A2(n1010), .A3(n1193), .ZN(n1171) );
AND3_X1 U883 ( .A1(n1046), .A2(n1200), .A3(n1020), .ZN(n1192) );
XNOR2_X1 U884 ( .A(G101), .B(n1160), .ZN(G3) );
NAND3_X1 U885 ( .A1(n1037), .A2(n1009), .A3(n1195), .ZN(n1160) );
XOR2_X1 U886 ( .A(n1183), .B(n1172), .Z(G27) );
NAND4_X1 U887 ( .A1(n1020), .A2(n1200), .A3(n1162), .A4(n1202), .ZN(n1172) );
AND2_X1 U888 ( .A1(n1203), .A2(n1034), .ZN(n1202) );
NAND2_X1 U889 ( .A1(n1052), .A2(n1204), .ZN(n1200) );
NAND4_X1 U890 ( .A1(G953), .A2(G902), .A3(n1205), .A4(n1083), .ZN(n1204) );
INV_X1 U891 ( .A(G900), .ZN(n1083) );
XOR2_X1 U892 ( .A(n1206), .B(G122), .Z(G24) );
NAND2_X1 U893 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
OR2_X1 U894 ( .A1(n1157), .A2(KEYINPUT28), .ZN(n1208) );
NAND3_X1 U895 ( .A1(n1196), .A2(n1011), .A3(n1209), .ZN(n1157) );
INV_X1 U896 ( .A(n1210), .ZN(n1196) );
NAND4_X1 U897 ( .A1(n1011), .A2(n1210), .A3(n1209), .A4(KEYINPUT28), .ZN(n1207) );
NAND2_X1 U898 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
NOR2_X1 U899 ( .A1(n1213), .A2(n1214), .ZN(n1011) );
XOR2_X1 U900 ( .A(n1215), .B(n1216), .Z(G21) );
NOR2_X1 U901 ( .A1(KEYINPUT0), .A2(n1217), .ZN(n1216) );
NAND2_X1 U902 ( .A1(n1218), .A2(n1219), .ZN(n1215) );
OR2_X1 U903 ( .A1(n1105), .A2(KEYINPUT33), .ZN(n1219) );
NAND2_X1 U904 ( .A1(n1209), .A2(n1198), .ZN(n1105) );
NAND3_X1 U905 ( .A1(n1020), .A2(n1220), .A3(KEYINPUT33), .ZN(n1218) );
NAND3_X1 U906 ( .A1(n1034), .A2(n1221), .A3(n1198), .ZN(n1220) );
AND2_X1 U907 ( .A1(n1193), .A2(n1037), .ZN(n1198) );
AND2_X1 U908 ( .A1(n1214), .A2(n1213), .ZN(n1193) );
INV_X1 U909 ( .A(n1222), .ZN(n1214) );
XNOR2_X1 U910 ( .A(G116), .B(n1155), .ZN(G18) );
NAND3_X1 U911 ( .A1(n1195), .A2(n1010), .A3(n1209), .ZN(n1155) );
NOR2_X1 U912 ( .A1(n1211), .A2(n1223), .ZN(n1010) );
XNOR2_X1 U913 ( .A(G113), .B(n1156), .ZN(G15) );
NAND3_X1 U914 ( .A1(n1195), .A2(n1162), .A3(n1209), .ZN(n1156) );
AND3_X1 U915 ( .A1(n1020), .A2(n1221), .A3(n1034), .ZN(n1209) );
NOR2_X1 U916 ( .A1(n1224), .A2(n1044), .ZN(n1034) );
INV_X1 U917 ( .A(n1045), .ZN(n1224) );
INV_X1 U918 ( .A(n1035), .ZN(n1162) );
NAND2_X1 U919 ( .A1(n1223), .A2(n1211), .ZN(n1035) );
NOR2_X1 U920 ( .A1(n1213), .A2(n1222), .ZN(n1195) );
XOR2_X1 U921 ( .A(n1161), .B(n1225), .Z(G12) );
XOR2_X1 U922 ( .A(n1226), .B(KEYINPUT39), .Z(n1225) );
NAND3_X1 U923 ( .A1(n1037), .A2(n1009), .A3(n1203), .ZN(n1161) );
INV_X1 U924 ( .A(n1049), .ZN(n1203) );
NAND2_X1 U925 ( .A1(n1222), .A2(n1213), .ZN(n1049) );
NAND2_X1 U926 ( .A1(n1227), .A2(n1056), .ZN(n1213) );
NAND2_X1 U927 ( .A1(n1228), .A2(n1229), .ZN(n1056) );
OR2_X1 U928 ( .A1(n1118), .A2(G902), .ZN(n1229) );
XOR2_X1 U929 ( .A(KEYINPUT55), .B(n1070), .Z(n1227) );
NOR3_X1 U930 ( .A1(n1228), .A2(G902), .A3(n1118), .ZN(n1070) );
XNOR2_X1 U931 ( .A(n1230), .B(G125), .ZN(n1118) );
XOR2_X1 U932 ( .A(n1231), .B(n1232), .Z(n1230) );
XOR2_X1 U933 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U934 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U935 ( .A1(KEYINPUT38), .A2(n1191), .ZN(n1236) );
NAND2_X1 U936 ( .A1(n1237), .A2(G221), .ZN(n1235) );
XOR2_X1 U937 ( .A(n1238), .B(G110), .Z(n1233) );
NAND2_X1 U938 ( .A1(KEYINPUT59), .A2(n1239), .ZN(n1238) );
XOR2_X1 U939 ( .A(KEYINPUT5), .B(G128), .Z(n1239) );
XOR2_X1 U940 ( .A(n1240), .B(n1241), .Z(n1231) );
XOR2_X1 U941 ( .A(KEYINPUT19), .B(G140), .Z(n1241) );
XOR2_X1 U942 ( .A(n1217), .B(G137), .Z(n1240) );
INV_X1 U943 ( .A(G119), .ZN(n1217) );
INV_X1 U944 ( .A(n1119), .ZN(n1228) );
NAND2_X1 U945 ( .A1(G217), .A2(n1242), .ZN(n1119) );
XOR2_X1 U946 ( .A(n1064), .B(G472), .Z(n1222) );
NAND2_X1 U947 ( .A1(n1243), .A2(n1244), .ZN(n1064) );
XOR2_X1 U948 ( .A(n1245), .B(n1246), .Z(n1243) );
XOR2_X1 U949 ( .A(n1141), .B(n1143), .Z(n1246) );
XOR2_X1 U950 ( .A(n1247), .B(n1248), .Z(n1245) );
XNOR2_X1 U951 ( .A(n1249), .B(KEYINPUT13), .ZN(n1248) );
NAND2_X1 U952 ( .A1(KEYINPUT42), .A2(n1136), .ZN(n1249) );
XNOR2_X1 U953 ( .A(n1250), .B(G113), .ZN(n1136) );
NAND2_X1 U954 ( .A1(KEYINPUT51), .A2(n1251), .ZN(n1250) );
NAND2_X1 U955 ( .A1(KEYINPUT4), .A2(n1135), .ZN(n1247) );
XNOR2_X1 U956 ( .A(n1252), .B(n1253), .ZN(n1135) );
NAND2_X1 U957 ( .A1(n1254), .A2(G210), .ZN(n1252) );
AND3_X1 U958 ( .A1(n1046), .A2(n1221), .A3(n1020), .ZN(n1009) );
NOR2_X1 U959 ( .A1(n1026), .A2(n1050), .ZN(n1020) );
INV_X1 U960 ( .A(n1028), .ZN(n1050) );
NAND2_X1 U961 ( .A1(n1255), .A2(n1256), .ZN(n1028) );
XNOR2_X1 U962 ( .A(G214), .B(KEYINPUT53), .ZN(n1255) );
XNOR2_X1 U963 ( .A(n1067), .B(n1069), .ZN(n1026) );
NAND2_X1 U964 ( .A1(G210), .A2(n1256), .ZN(n1069) );
NAND2_X1 U965 ( .A1(n1257), .A2(n1244), .ZN(n1256) );
INV_X1 U966 ( .A(G237), .ZN(n1257) );
NAND2_X1 U967 ( .A1(n1258), .A2(n1244), .ZN(n1067) );
XOR2_X1 U968 ( .A(n1180), .B(n1259), .Z(n1258) );
NOR2_X1 U969 ( .A1(KEYINPUT48), .A2(n1260), .ZN(n1259) );
XNOR2_X1 U970 ( .A(n1184), .B(n1261), .ZN(n1260) );
NAND2_X1 U971 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND2_X1 U972 ( .A1(G125), .A2(n1264), .ZN(n1263) );
INV_X1 U973 ( .A(n1141), .ZN(n1264) );
XOR2_X1 U974 ( .A(n1265), .B(KEYINPUT30), .Z(n1262) );
NAND2_X1 U975 ( .A1(n1141), .A2(n1183), .ZN(n1265) );
XOR2_X1 U976 ( .A(n1201), .B(n1266), .Z(n1141) );
NOR2_X1 U977 ( .A1(KEYINPUT1), .A2(n1267), .ZN(n1266) );
XOR2_X1 U978 ( .A(G146), .B(G143), .Z(n1267) );
AND2_X1 U979 ( .A1(G224), .A2(n1022), .ZN(n1184) );
NAND2_X1 U980 ( .A1(n1268), .A2(n1269), .ZN(n1180) );
NAND2_X1 U981 ( .A1(n1113), .A2(n1114), .ZN(n1269) );
XOR2_X1 U982 ( .A(n1270), .B(KEYINPUT34), .Z(n1268) );
OR2_X1 U983 ( .A1(n1114), .A2(n1113), .ZN(n1270) );
XNOR2_X1 U984 ( .A(n1226), .B(G122), .ZN(n1113) );
INV_X1 U985 ( .A(G110), .ZN(n1226) );
XNOR2_X1 U986 ( .A(n1271), .B(n1272), .ZN(n1114) );
XOR2_X1 U987 ( .A(G113), .B(n1273), .Z(n1272) );
NOR2_X1 U988 ( .A1(KEYINPUT16), .A2(n1274), .ZN(n1273) );
XOR2_X1 U989 ( .A(n1129), .B(G107), .Z(n1274) );
XOR2_X1 U990 ( .A(n1251), .B(n1253), .Z(n1271) );
XNOR2_X1 U991 ( .A(G116), .B(n1275), .ZN(n1251) );
XOR2_X1 U992 ( .A(KEYINPUT58), .B(G119), .Z(n1275) );
NAND2_X1 U993 ( .A1(n1052), .A2(n1276), .ZN(n1221) );
NAND4_X1 U994 ( .A1(G953), .A2(G902), .A3(n1205), .A4(n1111), .ZN(n1276) );
INV_X1 U995 ( .A(G898), .ZN(n1111) );
NAND3_X1 U996 ( .A1(n1205), .A2(n1022), .A3(G952), .ZN(n1052) );
NAND2_X1 U997 ( .A1(G237), .A2(G234), .ZN(n1205) );
NOR2_X1 U998 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
AND2_X1 U999 ( .A1(G221), .A2(n1242), .ZN(n1044) );
NAND2_X1 U1000 ( .A1(n1277), .A2(G234), .ZN(n1242) );
XOR2_X1 U1001 ( .A(n1244), .B(KEYINPUT3), .Z(n1277) );
XOR2_X1 U1002 ( .A(n1278), .B(G469), .Z(n1045) );
NAND2_X1 U1003 ( .A1(n1279), .A2(n1244), .ZN(n1278) );
XOR2_X1 U1004 ( .A(n1280), .B(n1147), .Z(n1279) );
XNOR2_X1 U1005 ( .A(n1281), .B(n1282), .ZN(n1147) );
XOR2_X1 U1006 ( .A(n1283), .B(n1284), .Z(n1282) );
XOR2_X1 U1007 ( .A(G110), .B(n1285), .Z(n1284) );
NOR2_X1 U1008 ( .A1(KEYINPUT23), .A2(n1286), .ZN(n1285) );
XOR2_X1 U1009 ( .A(n1007), .B(n1287), .Z(n1286) );
NOR2_X1 U1010 ( .A1(KEYINPUT60), .A2(n1129), .ZN(n1287) );
INV_X1 U1011 ( .A(G107), .ZN(n1007) );
NOR2_X1 U1012 ( .A1(G953), .A2(n1082), .ZN(n1283) );
INV_X1 U1013 ( .A(G227), .ZN(n1082) );
XNOR2_X1 U1014 ( .A(n1089), .B(n1288), .ZN(n1281) );
XOR2_X1 U1015 ( .A(n1253), .B(n1289), .Z(n1288) );
XOR2_X1 U1016 ( .A(G101), .B(KEYINPUT46), .Z(n1253) );
XNOR2_X1 U1017 ( .A(n1290), .B(G143), .ZN(n1089) );
NAND2_X1 U1018 ( .A1(KEYINPUT11), .A2(n1201), .ZN(n1290) );
INV_X1 U1019 ( .A(G128), .ZN(n1201) );
XOR2_X1 U1020 ( .A(n1143), .B(KEYINPUT21), .Z(n1280) );
XOR2_X1 U1021 ( .A(n1291), .B(n1292), .Z(n1143) );
XOR2_X1 U1022 ( .A(G137), .B(G131), .Z(n1292) );
NAND2_X1 U1023 ( .A1(KEYINPUT50), .A2(n1293), .ZN(n1291) );
INV_X1 U1024 ( .A(G134), .ZN(n1293) );
NOR2_X1 U1025 ( .A1(n1212), .A2(n1211), .ZN(n1037) );
XNOR2_X1 U1026 ( .A(n1294), .B(G475), .ZN(n1211) );
NAND2_X1 U1027 ( .A1(n1127), .A2(n1244), .ZN(n1294) );
INV_X1 U1028 ( .A(G902), .ZN(n1244) );
XNOR2_X1 U1029 ( .A(n1295), .B(n1296), .ZN(n1127) );
XOR2_X1 U1030 ( .A(n1297), .B(n1088), .Z(n1296) );
XOR2_X1 U1031 ( .A(G131), .B(n1289), .Z(n1088) );
XNOR2_X1 U1032 ( .A(G140), .B(n1191), .ZN(n1289) );
INV_X1 U1033 ( .A(G146), .ZN(n1191) );
AND2_X1 U1034 ( .A1(G214), .A2(n1254), .ZN(n1297) );
NOR2_X1 U1035 ( .A1(G953), .A2(G237), .ZN(n1254) );
XOR2_X1 U1036 ( .A(n1298), .B(n1299), .Z(n1295) );
XOR2_X1 U1037 ( .A(n1183), .B(n1300), .Z(n1299) );
NAND3_X1 U1038 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1300) );
NAND2_X1 U1039 ( .A1(n1304), .A2(n1305), .ZN(n1303) );
INV_X1 U1040 ( .A(KEYINPUT52), .ZN(n1305) );
NAND3_X1 U1041 ( .A1(KEYINPUT52), .A2(n1306), .A3(n1129), .ZN(n1302) );
OR2_X1 U1042 ( .A1(n1129), .A2(n1306), .ZN(n1301) );
NOR2_X1 U1043 ( .A1(KEYINPUT32), .A2(n1304), .ZN(n1306) );
XOR2_X1 U1044 ( .A(G113), .B(n1307), .Z(n1304) );
XOR2_X1 U1045 ( .A(KEYINPUT29), .B(G122), .Z(n1307) );
INV_X1 U1046 ( .A(G104), .ZN(n1129) );
INV_X1 U1047 ( .A(G125), .ZN(n1183) );
NAND2_X1 U1048 ( .A1(KEYINPUT31), .A2(n1308), .ZN(n1298) );
INV_X1 U1049 ( .A(G143), .ZN(n1308) );
INV_X1 U1050 ( .A(n1223), .ZN(n1212) );
XOR2_X1 U1051 ( .A(n1309), .B(G478), .Z(n1223) );
OR2_X1 U1052 ( .A1(n1123), .A2(G902), .ZN(n1309) );
XNOR2_X1 U1053 ( .A(n1310), .B(n1311), .ZN(n1123) );
XOR2_X1 U1054 ( .A(n1312), .B(n1313), .Z(n1311) );
XOR2_X1 U1055 ( .A(G116), .B(G107), .Z(n1313) );
XOR2_X1 U1056 ( .A(G143), .B(G134), .Z(n1312) );
XOR2_X1 U1057 ( .A(n1314), .B(n1315), .Z(n1310) );
XNOR2_X1 U1058 ( .A(n1316), .B(n1317), .ZN(n1315) );
NOR2_X1 U1059 ( .A1(G122), .A2(KEYINPUT57), .ZN(n1317) );
NAND2_X1 U1060 ( .A1(KEYINPUT27), .A2(G128), .ZN(n1316) );
NAND2_X1 U1061 ( .A1(G217), .A2(n1237), .ZN(n1314) );
AND2_X1 U1062 ( .A1(G234), .A2(n1022), .ZN(n1237) );
INV_X1 U1063 ( .A(G953), .ZN(n1022) );
endmodule


