//Key = 0101000001110001010110111000011101000111001010110001011001001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;

XOR2_X1 U742 ( .A(n1020), .B(n1021), .Z(G9) );
NOR2_X1 U743 ( .A1(KEYINPUT12), .A2(n1022), .ZN(n1021) );
NOR2_X1 U744 ( .A1(n1023), .A2(n1024), .ZN(G75) );
NOR3_X1 U745 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1024) );
NOR3_X1 U746 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n1026) );
NOR3_X1 U747 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1030) );
NOR2_X1 U748 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U749 ( .A1(n1036), .A2(n1037), .ZN(n1034) );
NOR2_X1 U750 ( .A1(n1038), .A2(KEYINPUT24), .ZN(n1032) );
NOR3_X1 U751 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1038) );
NOR3_X1 U752 ( .A1(n1040), .A2(n1042), .A3(n1043), .ZN(n1031) );
NOR4_X1 U753 ( .A1(n1039), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1043) );
AND2_X1 U754 ( .A1(n1047), .A2(KEYINPUT54), .ZN(n1046) );
NOR2_X1 U755 ( .A1(n1048), .A2(n1049), .ZN(n1045) );
INV_X1 U756 ( .A(n1050), .ZN(n1049) );
NOR2_X1 U757 ( .A1(n1051), .A2(n1052), .ZN(n1048) );
NOR2_X1 U758 ( .A1(n1053), .A2(n1054), .ZN(n1051) );
AND2_X1 U759 ( .A1(n1055), .A2(KEYINPUT24), .ZN(n1044) );
NOR2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1042) );
NOR2_X1 U761 ( .A1(KEYINPUT54), .A2(n1058), .ZN(n1057) );
INV_X1 U762 ( .A(n1059), .ZN(n1040) );
NAND3_X1 U763 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1025) );
NAND3_X1 U764 ( .A1(n1059), .A2(n1063), .A3(n1064), .ZN(n1062) );
INV_X1 U765 ( .A(n1035), .ZN(n1064) );
NAND3_X1 U766 ( .A1(n1065), .A2(n1050), .A3(n1056), .ZN(n1035) );
INV_X1 U767 ( .A(n1039), .ZN(n1056) );
NAND2_X1 U768 ( .A1(n1066), .A2(n1067), .ZN(n1063) );
NAND2_X1 U769 ( .A1(n1068), .A2(n1029), .ZN(n1067) );
INV_X1 U770 ( .A(n1069), .ZN(n1029) );
AND3_X1 U771 ( .A1(n1060), .A2(n1061), .A3(n1070), .ZN(n1023) );
NAND4_X1 U772 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1060) );
NOR4_X1 U773 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1074) );
XOR2_X1 U774 ( .A(KEYINPUT5), .B(n1079), .Z(n1078) );
XNOR2_X1 U775 ( .A(n1080), .B(n1081), .ZN(n1077) );
XOR2_X1 U776 ( .A(n1082), .B(G472), .Z(n1075) );
NAND2_X1 U777 ( .A1(KEYINPUT22), .A2(n1083), .ZN(n1082) );
AND3_X1 U778 ( .A1(n1069), .A2(n1084), .A3(n1054), .ZN(n1073) );
OR2_X1 U779 ( .A1(n1085), .A2(n1086), .ZN(n1072) );
XOR2_X1 U780 ( .A(n1087), .B(n1088), .Z(n1071) );
NAND2_X1 U781 ( .A1(KEYINPUT42), .A2(n1089), .ZN(n1088) );
XOR2_X1 U782 ( .A(n1090), .B(n1091), .Z(G72) );
NOR2_X1 U783 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NOR3_X1 U784 ( .A1(n1061), .A2(KEYINPUT61), .A3(n1094), .ZN(n1093) );
XOR2_X1 U785 ( .A(KEYINPUT32), .B(n1095), .Z(n1094) );
NOR2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
XNOR2_X1 U787 ( .A(KEYINPUT51), .B(n1098), .ZN(n1097) );
NOR2_X1 U788 ( .A1(G953), .A2(n1099), .ZN(n1092) );
NAND2_X1 U789 ( .A1(n1100), .A2(n1101), .ZN(n1090) );
NAND2_X1 U790 ( .A1(G953), .A2(n1098), .ZN(n1101) );
XOR2_X1 U791 ( .A(n1102), .B(n1103), .Z(n1100) );
XNOR2_X1 U792 ( .A(n1104), .B(n1105), .ZN(n1103) );
XOR2_X1 U793 ( .A(n1106), .B(n1107), .Z(n1102) );
NAND3_X1 U794 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1106) );
OR2_X1 U795 ( .A1(n1111), .A2(G137), .ZN(n1110) );
NAND2_X1 U796 ( .A1(n1112), .A2(n1113), .ZN(n1109) );
INV_X1 U797 ( .A(KEYINPUT3), .ZN(n1113) );
NAND2_X1 U798 ( .A1(n1114), .A2(G137), .ZN(n1112) );
XNOR2_X1 U799 ( .A(KEYINPUT55), .B(G134), .ZN(n1114) );
NAND2_X1 U800 ( .A1(KEYINPUT3), .A2(n1115), .ZN(n1108) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND3_X1 U802 ( .A1(G137), .A2(n1111), .A3(n1118), .ZN(n1117) );
INV_X1 U803 ( .A(KEYINPUT55), .ZN(n1118) );
NAND2_X1 U804 ( .A1(KEYINPUT55), .A2(G134), .ZN(n1116) );
XOR2_X1 U805 ( .A(n1119), .B(n1120), .Z(G69) );
XOR2_X1 U806 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U807 ( .A1(n1123), .A2(G953), .ZN(n1122) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1121) );
XNOR2_X1 U809 ( .A(n1126), .B(n1127), .ZN(n1125) );
XNOR2_X1 U810 ( .A(n1128), .B(KEYINPUT18), .ZN(n1126) );
NOR2_X1 U811 ( .A1(G898), .A2(n1061), .ZN(n1124) );
NOR2_X1 U812 ( .A1(n1129), .A2(n1061), .ZN(n1119) );
NOR2_X1 U813 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NOR2_X1 U814 ( .A1(n1132), .A2(n1133), .ZN(G66) );
NOR3_X1 U815 ( .A1(n1080), .A2(n1134), .A3(n1135), .ZN(n1133) );
AND3_X1 U816 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(n1135) );
INV_X1 U817 ( .A(n1081), .ZN(n1137) );
NOR2_X1 U818 ( .A1(n1139), .A2(n1136), .ZN(n1134) );
NOR2_X1 U819 ( .A1(n1140), .A2(n1081), .ZN(n1139) );
NOR3_X1 U820 ( .A1(n1132), .A2(n1141), .A3(n1142), .ZN(G63) );
NOR2_X1 U821 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
NOR2_X1 U822 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NOR2_X1 U823 ( .A1(KEYINPUT30), .A2(n1147), .ZN(n1146) );
NOR3_X1 U824 ( .A1(n1148), .A2(KEYINPUT6), .A3(n1149), .ZN(n1145) );
INV_X1 U825 ( .A(KEYINPUT30), .ZN(n1149) );
NOR2_X1 U826 ( .A1(n1150), .A2(n1151), .ZN(n1141) );
INV_X1 U827 ( .A(n1143), .ZN(n1151) );
NOR2_X1 U828 ( .A1(KEYINPUT6), .A2(n1148), .ZN(n1150) );
INV_X1 U829 ( .A(n1147), .ZN(n1148) );
NAND2_X1 U830 ( .A1(n1138), .A2(G478), .ZN(n1147) );
NOR2_X1 U831 ( .A1(n1132), .A2(n1152), .ZN(G60) );
XOR2_X1 U832 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U833 ( .A1(KEYINPUT46), .A2(n1155), .ZN(n1153) );
NAND2_X1 U834 ( .A1(n1138), .A2(G475), .ZN(n1155) );
XNOR2_X1 U835 ( .A(n1156), .B(n1157), .ZN(G6) );
NOR2_X1 U836 ( .A1(n1158), .A2(n1066), .ZN(n1157) );
XOR2_X1 U837 ( .A(n1159), .B(KEYINPUT36), .Z(n1158) );
NOR2_X1 U838 ( .A1(n1132), .A2(n1160), .ZN(G57) );
XOR2_X1 U839 ( .A(n1161), .B(n1162), .Z(n1160) );
XNOR2_X1 U840 ( .A(n1163), .B(n1164), .ZN(n1162) );
NAND2_X1 U841 ( .A1(KEYINPUT62), .A2(n1165), .ZN(n1163) );
XOR2_X1 U842 ( .A(n1166), .B(n1167), .Z(n1161) );
NAND2_X1 U843 ( .A1(KEYINPUT10), .A2(n1168), .ZN(n1167) );
NAND2_X1 U844 ( .A1(n1138), .A2(G472), .ZN(n1166) );
NOR2_X1 U845 ( .A1(n1132), .A2(n1169), .ZN(G54) );
XOR2_X1 U846 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U847 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U848 ( .A1(n1174), .A2(n1175), .ZN(n1173) );
NOR2_X1 U849 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
NOR2_X1 U850 ( .A1(KEYINPUT58), .A2(G110), .ZN(n1177) );
NOR2_X1 U851 ( .A1(G140), .A2(n1178), .ZN(n1176) );
NOR2_X1 U852 ( .A1(KEYINPUT39), .A2(n1179), .ZN(n1178) );
NOR4_X1 U853 ( .A1(KEYINPUT58), .A2(G140), .A3(G110), .A4(n1180), .ZN(n1174) );
INV_X1 U854 ( .A(KEYINPUT39), .ZN(n1180) );
NAND2_X1 U855 ( .A1(n1138), .A2(G469), .ZN(n1172) );
NOR3_X1 U856 ( .A1(n1181), .A2(n1182), .A3(n1183), .ZN(G51) );
AND2_X1 U857 ( .A1(KEYINPUT15), .A2(n1132), .ZN(n1183) );
NOR2_X1 U858 ( .A1(n1061), .A2(G952), .ZN(n1132) );
NOR3_X1 U859 ( .A1(KEYINPUT15), .A2(n1061), .A3(n1070), .ZN(n1182) );
XOR2_X1 U860 ( .A(n1184), .B(n1185), .Z(n1181) );
XOR2_X1 U861 ( .A(n1186), .B(n1187), .Z(n1184) );
NOR2_X1 U862 ( .A1(KEYINPUT40), .A2(n1188), .ZN(n1187) );
XOR2_X1 U863 ( .A(n1189), .B(n1190), .Z(n1188) );
NOR2_X1 U864 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U865 ( .A(n1193), .B(KEYINPUT23), .Z(n1192) );
NAND2_X1 U866 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NAND2_X1 U867 ( .A1(n1138), .A2(n1196), .ZN(n1186) );
INV_X1 U868 ( .A(n1089), .ZN(n1196) );
NOR2_X1 U869 ( .A1(n1197), .A2(n1140), .ZN(n1138) );
INV_X1 U870 ( .A(n1027), .ZN(n1140) );
NAND2_X1 U871 ( .A1(n1099), .A2(n1123), .ZN(n1027) );
AND4_X1 U872 ( .A1(n1198), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1123) );
NOR4_X1 U873 ( .A1(n1020), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1201) );
AND4_X1 U874 ( .A1(n1050), .A2(n1036), .A3(n1205), .A4(n1206), .ZN(n1020) );
NOR2_X1 U875 ( .A1(n1207), .A2(n1208), .ZN(n1200) );
NAND2_X1 U876 ( .A1(n1209), .A2(n1210), .ZN(n1199) );
NAND2_X1 U877 ( .A1(n1159), .A2(n1211), .ZN(n1210) );
NAND2_X1 U878 ( .A1(KEYINPUT63), .A2(n1212), .ZN(n1211) );
NAND4_X1 U879 ( .A1(n1037), .A2(n1050), .A3(n1205), .A4(n1213), .ZN(n1159) );
OR3_X1 U880 ( .A1(n1214), .A2(KEYINPUT63), .A3(n1209), .ZN(n1198) );
AND2_X1 U881 ( .A1(n1215), .A2(n1216), .ZN(n1099) );
NOR4_X1 U882 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
NOR4_X1 U883 ( .A1(n1221), .A2(n1222), .A3(n1223), .A4(n1224), .ZN(n1215) );
AND4_X1 U884 ( .A1(n1225), .A2(n1205), .A3(n1036), .A4(n1226), .ZN(n1224) );
XOR2_X1 U885 ( .A(n1223), .B(n1227), .Z(G48) );
NOR2_X1 U886 ( .A1(KEYINPUT41), .A2(n1228), .ZN(n1227) );
AND4_X1 U887 ( .A1(n1052), .A2(n1226), .A3(n1037), .A4(n1225), .ZN(n1223) );
XNOR2_X1 U888 ( .A(n1222), .B(n1229), .ZN(G45) );
NAND2_X1 U889 ( .A1(KEYINPUT29), .A2(G143), .ZN(n1229) );
AND3_X1 U890 ( .A1(n1052), .A2(n1226), .A3(n1230), .ZN(n1222) );
AND3_X1 U891 ( .A1(n1231), .A2(n1232), .A3(n1076), .ZN(n1230) );
XNOR2_X1 U892 ( .A(n1233), .B(n1221), .ZN(G42) );
AND3_X1 U893 ( .A1(n1037), .A2(n1234), .A3(n1235), .ZN(n1221) );
XOR2_X1 U894 ( .A(G137), .B(n1220), .Z(G39) );
AND3_X1 U895 ( .A1(n1235), .A2(n1225), .A3(n1059), .ZN(n1220) );
XNOR2_X1 U896 ( .A(n1111), .B(n1219), .ZN(G36) );
AND3_X1 U897 ( .A1(n1036), .A2(n1231), .A3(n1235), .ZN(n1219) );
XOR2_X1 U898 ( .A(G131), .B(n1218), .Z(G33) );
AND3_X1 U899 ( .A1(n1037), .A2(n1231), .A3(n1235), .ZN(n1218) );
AND4_X1 U900 ( .A1(n1052), .A2(n1068), .A3(n1236), .A4(n1069), .ZN(n1235) );
INV_X1 U901 ( .A(n1028), .ZN(n1068) );
XOR2_X1 U902 ( .A(n1237), .B(KEYINPUT60), .Z(n1052) );
XOR2_X1 U903 ( .A(n1238), .B(n1239), .Z(G30) );
NOR2_X1 U904 ( .A1(KEYINPUT8), .A2(n1240), .ZN(n1239) );
NOR4_X1 U905 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1238) );
XNOR2_X1 U906 ( .A(KEYINPUT34), .B(n1236), .ZN(n1244) );
INV_X1 U907 ( .A(n1036), .ZN(n1243) );
NAND2_X1 U908 ( .A1(n1209), .A2(n1225), .ZN(n1242) );
XOR2_X1 U909 ( .A(G101), .B(n1208), .Z(G3) );
AND2_X1 U910 ( .A1(n1245), .A2(n1231), .ZN(n1208) );
XNOR2_X1 U911 ( .A(n1217), .B(n1246), .ZN(G27) );
NAND2_X1 U912 ( .A1(KEYINPUT31), .A2(n1247), .ZN(n1246) );
XNOR2_X1 U913 ( .A(KEYINPUT21), .B(n1195), .ZN(n1247) );
AND3_X1 U914 ( .A1(n1047), .A2(n1037), .A3(n1226), .ZN(n1217) );
AND2_X1 U915 ( .A1(n1209), .A2(n1236), .ZN(n1226) );
NAND2_X1 U916 ( .A1(n1039), .A2(n1248), .ZN(n1236) );
NAND4_X1 U917 ( .A1(G953), .A2(G902), .A3(n1249), .A4(n1098), .ZN(n1248) );
INV_X1 U918 ( .A(G900), .ZN(n1098) );
INV_X1 U919 ( .A(n1058), .ZN(n1047) );
NAND2_X1 U920 ( .A1(n1065), .A2(n1234), .ZN(n1058) );
XOR2_X1 U921 ( .A(G122), .B(n1207), .Z(G24) );
AND4_X1 U922 ( .A1(n1250), .A2(n1050), .A3(n1076), .A4(n1232), .ZN(n1207) );
XOR2_X1 U923 ( .A(G119), .B(n1204), .Z(G21) );
AND3_X1 U924 ( .A1(n1059), .A2(n1225), .A3(n1250), .ZN(n1204) );
NAND2_X1 U925 ( .A1(n1251), .A2(n1252), .ZN(n1225) );
NAND2_X1 U926 ( .A1(n1234), .A2(n1253), .ZN(n1252) );
NAND3_X1 U927 ( .A1(n1254), .A2(n1255), .A3(KEYINPUT57), .ZN(n1251) );
XOR2_X1 U928 ( .A(G116), .B(n1203), .Z(G18) );
AND3_X1 U929 ( .A1(n1036), .A2(n1231), .A3(n1250), .ZN(n1203) );
AND2_X1 U930 ( .A1(n1065), .A2(n1206), .ZN(n1250) );
NOR2_X1 U931 ( .A1(n1232), .A2(n1256), .ZN(n1036) );
XOR2_X1 U932 ( .A(G113), .B(n1257), .Z(G15) );
NOR2_X1 U933 ( .A1(n1258), .A2(n1066), .ZN(n1257) );
XNOR2_X1 U934 ( .A(n1212), .B(KEYINPUT56), .ZN(n1258) );
INV_X1 U935 ( .A(n1214), .ZN(n1212) );
NAND3_X1 U936 ( .A1(n1037), .A2(n1213), .A3(n1055), .ZN(n1214) );
INV_X1 U937 ( .A(n1041), .ZN(n1055) );
NAND2_X1 U938 ( .A1(n1065), .A2(n1231), .ZN(n1041) );
NAND2_X1 U939 ( .A1(n1259), .A2(n1260), .ZN(n1231) );
NAND2_X1 U940 ( .A1(n1050), .A2(n1253), .ZN(n1260) );
INV_X1 U941 ( .A(KEYINPUT57), .ZN(n1253) );
NOR2_X1 U942 ( .A1(n1255), .A2(n1254), .ZN(n1050) );
NAND3_X1 U943 ( .A1(n1261), .A2(n1254), .A3(KEYINPUT57), .ZN(n1259) );
NOR2_X1 U944 ( .A1(n1053), .A2(n1262), .ZN(n1065) );
INV_X1 U945 ( .A(n1054), .ZN(n1262) );
AND2_X1 U946 ( .A1(n1256), .A2(n1232), .ZN(n1037) );
INV_X1 U947 ( .A(n1076), .ZN(n1256) );
NAND2_X1 U948 ( .A1(n1263), .A2(n1264), .ZN(G12) );
NAND2_X1 U949 ( .A1(n1202), .A2(n1179), .ZN(n1264) );
XOR2_X1 U950 ( .A(KEYINPUT38), .B(n1265), .Z(n1263) );
NOR2_X1 U951 ( .A1(n1202), .A2(n1179), .ZN(n1265) );
AND2_X1 U952 ( .A1(n1245), .A2(n1234), .ZN(n1202) );
NOR2_X1 U953 ( .A1(n1254), .A2(n1261), .ZN(n1234) );
INV_X1 U954 ( .A(n1255), .ZN(n1261) );
XOR2_X1 U955 ( .A(n1081), .B(n1266), .Z(n1255) );
NOR2_X1 U956 ( .A1(n1267), .A2(n1268), .ZN(n1266) );
NOR2_X1 U957 ( .A1(KEYINPUT44), .A2(n1080), .ZN(n1268) );
NOR2_X1 U958 ( .A1(KEYINPUT14), .A2(n1269), .ZN(n1267) );
INV_X1 U959 ( .A(n1080), .ZN(n1269) );
NOR2_X1 U960 ( .A1(n1136), .A2(G902), .ZN(n1080) );
XOR2_X1 U961 ( .A(n1270), .B(n1105), .Z(n1136) );
INV_X1 U962 ( .A(n1271), .ZN(n1105) );
XOR2_X1 U963 ( .A(n1272), .B(n1273), .Z(n1270) );
XOR2_X1 U964 ( .A(n1274), .B(n1275), .Z(n1273) );
XNOR2_X1 U965 ( .A(n1228), .B(G137), .ZN(n1275) );
XOR2_X1 U966 ( .A(KEYINPUT43), .B(KEYINPUT20), .Z(n1274) );
XOR2_X1 U967 ( .A(n1276), .B(n1277), .Z(n1272) );
XNOR2_X1 U968 ( .A(n1240), .B(G119), .ZN(n1277) );
XOR2_X1 U969 ( .A(n1278), .B(n1279), .Z(n1276) );
NOR2_X1 U970 ( .A1(KEYINPUT2), .A2(n1179), .ZN(n1279) );
NAND2_X1 U971 ( .A1(G221), .A2(n1280), .ZN(n1278) );
NAND2_X1 U972 ( .A1(G217), .A2(n1281), .ZN(n1081) );
XNOR2_X1 U973 ( .A(n1083), .B(G472), .ZN(n1254) );
NAND2_X1 U974 ( .A1(n1282), .A2(n1197), .ZN(n1083) );
XNOR2_X1 U975 ( .A(n1283), .B(n1165), .ZN(n1282) );
XNOR2_X1 U976 ( .A(n1284), .B(n1285), .ZN(n1165) );
NAND2_X1 U977 ( .A1(G210), .A2(n1286), .ZN(n1284) );
XNOR2_X1 U978 ( .A(n1168), .B(n1127), .ZN(n1283) );
XOR2_X1 U979 ( .A(n1287), .B(n1288), .Z(n1168) );
AND3_X1 U980 ( .A1(n1205), .A2(n1206), .A3(n1059), .ZN(n1245) );
NOR2_X1 U981 ( .A1(n1076), .A2(n1232), .ZN(n1059) );
NAND3_X1 U982 ( .A1(n1289), .A2(n1290), .A3(n1084), .ZN(n1232) );
NAND2_X1 U983 ( .A1(n1086), .A2(n1085), .ZN(n1084) );
OR3_X1 U984 ( .A1(n1085), .A2(n1086), .A3(KEYINPUT48), .ZN(n1290) );
NOR2_X1 U985 ( .A1(n1154), .A2(G902), .ZN(n1086) );
XNOR2_X1 U986 ( .A(n1291), .B(n1292), .ZN(n1154) );
XOR2_X1 U987 ( .A(n1293), .B(n1294), .Z(n1292) );
XNOR2_X1 U988 ( .A(n1295), .B(n1156), .ZN(n1294) );
NAND2_X1 U989 ( .A1(G214), .A2(n1286), .ZN(n1295) );
NOR2_X1 U990 ( .A1(G953), .A2(G237), .ZN(n1286) );
XNOR2_X1 U991 ( .A(G113), .B(G131), .ZN(n1293) );
XNOR2_X1 U992 ( .A(n1271), .B(n1296), .ZN(n1291) );
XOR2_X1 U993 ( .A(n1297), .B(n1298), .Z(n1296) );
NOR2_X1 U994 ( .A1(G146), .A2(KEYINPUT45), .ZN(n1297) );
XNOR2_X1 U995 ( .A(G125), .B(n1233), .ZN(n1271) );
INV_X1 U996 ( .A(G140), .ZN(n1233) );
NAND2_X1 U997 ( .A1(KEYINPUT48), .A2(n1085), .ZN(n1289) );
INV_X1 U998 ( .A(G475), .ZN(n1085) );
XNOR2_X1 U999 ( .A(n1299), .B(n1300), .ZN(n1076) );
XOR2_X1 U1000 ( .A(KEYINPUT25), .B(G478), .Z(n1300) );
NAND2_X1 U1001 ( .A1(n1143), .A2(n1197), .ZN(n1299) );
XNOR2_X1 U1002 ( .A(n1301), .B(n1302), .ZN(n1143) );
XOR2_X1 U1003 ( .A(G116), .B(n1303), .Z(n1302) );
XNOR2_X1 U1004 ( .A(n1111), .B(G128), .ZN(n1303) );
INV_X1 U1005 ( .A(G134), .ZN(n1111) );
XOR2_X1 U1006 ( .A(n1304), .B(n1298), .Z(n1301) );
XOR2_X1 U1007 ( .A(G122), .B(G143), .Z(n1298) );
XNOR2_X1 U1008 ( .A(n1305), .B(n1022), .ZN(n1304) );
NAND2_X1 U1009 ( .A1(n1280), .A2(G217), .ZN(n1305) );
AND2_X1 U1010 ( .A1(G234), .A2(n1061), .ZN(n1280) );
AND2_X1 U1011 ( .A1(n1209), .A2(n1213), .ZN(n1206) );
NAND2_X1 U1012 ( .A1(n1039), .A2(n1306), .ZN(n1213) );
NAND4_X1 U1013 ( .A1(G953), .A2(G902), .A3(n1249), .A4(n1131), .ZN(n1306) );
INV_X1 U1014 ( .A(G898), .ZN(n1131) );
NAND3_X1 U1015 ( .A1(n1249), .A2(n1061), .A3(n1307), .ZN(n1039) );
XNOR2_X1 U1016 ( .A(KEYINPUT16), .B(n1070), .ZN(n1307) );
INV_X1 U1017 ( .A(G952), .ZN(n1070) );
INV_X1 U1018 ( .A(G953), .ZN(n1061) );
NAND2_X1 U1019 ( .A1(G237), .A2(G234), .ZN(n1249) );
INV_X1 U1020 ( .A(n1066), .ZN(n1209) );
NAND2_X1 U1021 ( .A1(n1308), .A2(n1028), .ZN(n1066) );
XNOR2_X1 U1022 ( .A(n1087), .B(n1309), .ZN(n1028) );
XOR2_X1 U1023 ( .A(KEYINPUT26), .B(n1310), .Z(n1309) );
NOR2_X1 U1024 ( .A1(KEYINPUT52), .A2(n1089), .ZN(n1310) );
NAND2_X1 U1025 ( .A1(G210), .A2(n1311), .ZN(n1089) );
NAND2_X1 U1026 ( .A1(n1312), .A2(n1197), .ZN(n1087) );
XNOR2_X1 U1027 ( .A(n1185), .B(n1313), .ZN(n1312) );
NOR2_X1 U1028 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
XNOR2_X1 U1029 ( .A(n1189), .B(n1316), .ZN(n1315) );
XOR2_X1 U1030 ( .A(n1317), .B(KEYINPUT47), .Z(n1316) );
NAND2_X1 U1031 ( .A1(n1318), .A2(n1319), .ZN(n1317) );
NAND2_X1 U1032 ( .A1(n1320), .A2(n1195), .ZN(n1319) );
OR2_X1 U1033 ( .A1(n1194), .A2(KEYINPUT7), .ZN(n1320) );
NAND2_X1 U1034 ( .A1(n1191), .A2(n1321), .ZN(n1318) );
INV_X1 U1035 ( .A(KEYINPUT7), .ZN(n1321) );
NOR2_X1 U1036 ( .A1(n1195), .A2(n1194), .ZN(n1191) );
XNOR2_X1 U1037 ( .A(n1287), .B(n1240), .ZN(n1194) );
INV_X1 U1038 ( .A(G128), .ZN(n1240) );
XOR2_X1 U1039 ( .A(n1322), .B(G143), .Z(n1287) );
NAND2_X1 U1040 ( .A1(KEYINPUT53), .A2(n1228), .ZN(n1322) );
INV_X1 U1041 ( .A(G146), .ZN(n1228) );
INV_X1 U1042 ( .A(G125), .ZN(n1195) );
NOR2_X1 U1043 ( .A1(n1130), .A2(G953), .ZN(n1189) );
INV_X1 U1044 ( .A(G224), .ZN(n1130) );
XOR2_X1 U1045 ( .A(KEYINPUT49), .B(KEYINPUT35), .Z(n1314) );
XOR2_X1 U1046 ( .A(n1323), .B(n1324), .Z(n1185) );
INV_X1 U1047 ( .A(n1128), .ZN(n1324) );
XNOR2_X1 U1048 ( .A(n1325), .B(n1326), .ZN(n1128) );
XNOR2_X1 U1049 ( .A(G122), .B(n1179), .ZN(n1326) );
XNOR2_X1 U1050 ( .A(n1327), .B(n1285), .ZN(n1325) );
NAND3_X1 U1051 ( .A1(n1328), .A2(n1329), .A3(n1330), .ZN(n1327) );
NAND2_X1 U1052 ( .A1(G104), .A2(n1022), .ZN(n1330) );
NAND2_X1 U1053 ( .A1(KEYINPUT50), .A2(n1331), .ZN(n1329) );
NAND2_X1 U1054 ( .A1(n1332), .A2(n1156), .ZN(n1331) );
XNOR2_X1 U1055 ( .A(KEYINPUT59), .B(n1022), .ZN(n1332) );
NAND2_X1 U1056 ( .A1(n1333), .A2(n1334), .ZN(n1328) );
INV_X1 U1057 ( .A(KEYINPUT50), .ZN(n1334) );
NAND2_X1 U1058 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
OR3_X1 U1059 ( .A1(n1022), .A2(G104), .A3(KEYINPUT59), .ZN(n1336) );
NAND2_X1 U1060 ( .A1(KEYINPUT59), .A2(n1022), .ZN(n1335) );
NAND2_X1 U1061 ( .A1(KEYINPUT9), .A2(n1127), .ZN(n1323) );
INV_X1 U1062 ( .A(n1164), .ZN(n1127) );
XOR2_X1 U1063 ( .A(G113), .B(n1337), .Z(n1164) );
XOR2_X1 U1064 ( .A(G119), .B(G116), .Z(n1337) );
XNOR2_X1 U1065 ( .A(KEYINPUT33), .B(n1069), .ZN(n1308) );
NAND2_X1 U1066 ( .A1(G214), .A2(n1311), .ZN(n1069) );
NAND2_X1 U1067 ( .A1(n1338), .A2(n1339), .ZN(n1311) );
INV_X1 U1068 ( .A(G237), .ZN(n1339) );
XNOR2_X1 U1069 ( .A(KEYINPUT37), .B(n1197), .ZN(n1338) );
INV_X1 U1070 ( .A(n1241), .ZN(n1205) );
XNOR2_X1 U1071 ( .A(n1237), .B(KEYINPUT17), .ZN(n1241) );
NAND2_X1 U1072 ( .A1(n1053), .A2(n1054), .ZN(n1237) );
NAND2_X1 U1073 ( .A1(G221), .A2(n1281), .ZN(n1054) );
NAND2_X1 U1074 ( .A1(n1340), .A2(n1197), .ZN(n1281) );
XNOR2_X1 U1075 ( .A(G234), .B(KEYINPUT11), .ZN(n1340) );
XNOR2_X1 U1076 ( .A(n1079), .B(KEYINPUT1), .ZN(n1053) );
XNOR2_X1 U1077 ( .A(n1341), .B(G469), .ZN(n1079) );
NAND2_X1 U1078 ( .A1(n1342), .A2(n1197), .ZN(n1341) );
INV_X1 U1079 ( .A(G902), .ZN(n1197) );
XOR2_X1 U1080 ( .A(n1343), .B(n1344), .Z(n1342) );
XNOR2_X1 U1081 ( .A(G140), .B(n1345), .ZN(n1344) );
XNOR2_X1 U1082 ( .A(KEYINPUT4), .B(KEYINPUT0), .ZN(n1345) );
XNOR2_X1 U1083 ( .A(n1170), .B(n1179), .ZN(n1343) );
INV_X1 U1084 ( .A(G110), .ZN(n1179) );
XOR2_X1 U1085 ( .A(n1346), .B(n1347), .Z(n1170) );
XNOR2_X1 U1086 ( .A(n1288), .B(n1348), .ZN(n1347) );
INV_X1 U1087 ( .A(n1104), .ZN(n1348) );
XOR2_X1 U1088 ( .A(G146), .B(n1349), .Z(n1104) );
NOR2_X1 U1089 ( .A1(G143), .A2(KEYINPUT27), .ZN(n1349) );
XNOR2_X1 U1090 ( .A(n1350), .B(n1107), .ZN(n1288) );
XOR2_X1 U1091 ( .A(G131), .B(G128), .Z(n1107) );
XNOR2_X1 U1092 ( .A(G134), .B(G137), .ZN(n1350) );
XOR2_X1 U1093 ( .A(n1351), .B(n1352), .Z(n1346) );
NOR2_X1 U1094 ( .A1(G953), .A2(n1096), .ZN(n1352) );
INV_X1 U1095 ( .A(G227), .ZN(n1096) );
NAND2_X1 U1096 ( .A1(n1353), .A2(n1354), .ZN(n1351) );
OR2_X1 U1097 ( .A1(n1355), .A2(n1285), .ZN(n1354) );
XOR2_X1 U1098 ( .A(n1356), .B(KEYINPUT28), .Z(n1353) );
NAND2_X1 U1099 ( .A1(n1285), .A2(n1355), .ZN(n1356) );
XOR2_X1 U1100 ( .A(n1357), .B(n1022), .Z(n1355) );
INV_X1 U1101 ( .A(G107), .ZN(n1022) );
NAND2_X1 U1102 ( .A1(KEYINPUT19), .A2(n1156), .ZN(n1357) );
INV_X1 U1103 ( .A(G104), .ZN(n1156) );
XNOR2_X1 U1104 ( .A(G101), .B(KEYINPUT13), .ZN(n1285) );
endmodule


