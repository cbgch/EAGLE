//Key = 0001011011110010110001100110000111100000100100111001010111111100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246;

XOR2_X1 U688 ( .A(n948), .B(n949), .Z(G9) );
NAND2_X1 U689 ( .A1(n950), .A2(n951), .ZN(n949) );
XNOR2_X1 U690 ( .A(n952), .B(KEYINPUT51), .ZN(n950) );
NOR2_X1 U691 ( .A1(n953), .A2(n954), .ZN(G75) );
NOR4_X1 U692 ( .A1(n955), .A2(n956), .A3(n957), .A4(n958), .ZN(n954) );
NOR2_X1 U693 ( .A1(n959), .A2(n960), .ZN(n958) );
XOR2_X1 U694 ( .A(n961), .B(KEYINPUT63), .Z(n960) );
NOR3_X1 U695 ( .A1(n961), .A2(n962), .A3(n963), .ZN(n957) );
XNOR2_X1 U696 ( .A(n964), .B(KEYINPUT20), .ZN(n963) );
NAND4_X1 U697 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(n961) );
AND2_X1 U698 ( .A1(n969), .A2(KEYINPUT43), .ZN(n968) );
NAND3_X1 U699 ( .A1(n970), .A2(n971), .A3(n972), .ZN(n955) );
NAND4_X1 U700 ( .A1(KEYINPUT43), .A2(n973), .A3(n974), .A4(n966), .ZN(n972) );
NAND2_X1 U701 ( .A1(n975), .A2(n976), .ZN(n974) );
NAND3_X1 U702 ( .A1(n965), .A2(n977), .A3(n967), .ZN(n976) );
OR2_X1 U703 ( .A1(n978), .A2(n979), .ZN(n977) );
NAND2_X1 U704 ( .A1(n969), .A2(n980), .ZN(n975) );
NAND2_X1 U705 ( .A1(n981), .A2(n982), .ZN(n980) );
NAND2_X1 U706 ( .A1(n965), .A2(n983), .ZN(n982) );
NAND2_X1 U707 ( .A1(n984), .A2(n985), .ZN(n983) );
NAND2_X1 U708 ( .A1(n986), .A2(n987), .ZN(n985) );
NAND2_X1 U709 ( .A1(n967), .A2(n988), .ZN(n981) );
OR2_X1 U710 ( .A1(n989), .A2(n990), .ZN(n988) );
NOR3_X1 U711 ( .A1(n991), .A2(G953), .A3(G952), .ZN(n953) );
INV_X1 U712 ( .A(n970), .ZN(n991) );
NAND4_X1 U713 ( .A1(n992), .A2(n993), .A3(n994), .A4(n995), .ZN(n970) );
NOR4_X1 U714 ( .A1(n964), .A2(n986), .A3(n996), .A4(n997), .ZN(n995) );
XOR2_X1 U715 ( .A(n998), .B(n999), .Z(n997) );
XNOR2_X1 U716 ( .A(n1000), .B(KEYINPUT11), .ZN(n998) );
XNOR2_X1 U717 ( .A(n1001), .B(n1002), .ZN(n996) );
NAND2_X1 U718 ( .A1(KEYINPUT58), .A2(n1003), .ZN(n1001) );
NOR2_X1 U719 ( .A1(n1004), .A2(n1005), .ZN(n994) );
XOR2_X1 U720 ( .A(KEYINPUT28), .B(n1006), .Z(n1005) );
XOR2_X1 U721 ( .A(G475), .B(n1007), .Z(n1004) );
XOR2_X1 U722 ( .A(n1008), .B(n1009), .Z(n993) );
XOR2_X1 U723 ( .A(KEYINPUT31), .B(n1010), .Z(n992) );
XOR2_X1 U724 ( .A(n1011), .B(n1012), .Z(G72) );
XOR2_X1 U725 ( .A(n1013), .B(n1014), .Z(n1012) );
NOR2_X1 U726 ( .A1(G953), .A2(n1015), .ZN(n1014) );
XOR2_X1 U727 ( .A(n1016), .B(KEYINPUT26), .Z(n1015) );
NAND2_X1 U728 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
XNOR2_X1 U729 ( .A(KEYINPUT57), .B(n1019), .ZN(n1018) );
NAND2_X1 U730 ( .A1(n1020), .A2(n1021), .ZN(n1013) );
OR2_X1 U731 ( .A1(n971), .A2(G900), .ZN(n1021) );
XOR2_X1 U732 ( .A(n1022), .B(n1023), .Z(n1020) );
NOR2_X1 U733 ( .A1(KEYINPUT38), .A2(n1024), .ZN(n1023) );
XOR2_X1 U734 ( .A(G137), .B(n1025), .Z(n1024) );
NAND2_X1 U735 ( .A1(n1026), .A2(n1027), .ZN(n1022) );
NAND2_X1 U736 ( .A1(G125), .A2(n1028), .ZN(n1027) );
XOR2_X1 U737 ( .A(n1029), .B(KEYINPUT7), .Z(n1026) );
NAND2_X1 U738 ( .A1(G140), .A2(n1030), .ZN(n1029) );
NAND2_X1 U739 ( .A1(G953), .A2(n1031), .ZN(n1011) );
NAND2_X1 U740 ( .A1(G900), .A2(G227), .ZN(n1031) );
XOR2_X1 U741 ( .A(n1032), .B(n1033), .Z(G69) );
XOR2_X1 U742 ( .A(n1034), .B(n1035), .Z(n1033) );
NOR2_X1 U743 ( .A1(n1036), .A2(n971), .ZN(n1035) );
NOR2_X1 U744 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND2_X1 U745 ( .A1(n1039), .A2(n1040), .ZN(n1034) );
NAND2_X1 U746 ( .A1(G953), .A2(n1038), .ZN(n1040) );
XOR2_X1 U747 ( .A(n1041), .B(n1042), .Z(n1039) );
NAND2_X1 U748 ( .A1(n971), .A2(n1043), .ZN(n1032) );
NAND2_X1 U749 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U750 ( .A1(n1046), .A2(n1047), .ZN(G66) );
NOR3_X1 U751 ( .A1(n1000), .A2(n1048), .A3(n1049), .ZN(n1047) );
AND3_X1 U752 ( .A1(n1050), .A2(n999), .A3(n1051), .ZN(n1049) );
NOR2_X1 U753 ( .A1(n1052), .A2(n1050), .ZN(n1048) );
AND2_X1 U754 ( .A1(n956), .A2(n999), .ZN(n1052) );
NOR2_X1 U755 ( .A1(n1046), .A2(n1053), .ZN(G63) );
XOR2_X1 U756 ( .A(n1054), .B(n1055), .Z(n1053) );
NOR2_X1 U757 ( .A1(KEYINPUT45), .A2(n1056), .ZN(n1055) );
NAND2_X1 U758 ( .A1(n1051), .A2(G478), .ZN(n1054) );
NOR2_X1 U759 ( .A1(n1046), .A2(n1057), .ZN(G60) );
NOR3_X1 U760 ( .A1(n1007), .A2(n1058), .A3(n1059), .ZN(n1057) );
AND3_X1 U761 ( .A1(n1060), .A2(G475), .A3(n1051), .ZN(n1059) );
NOR2_X1 U762 ( .A1(n1061), .A2(n1060), .ZN(n1058) );
AND2_X1 U763 ( .A1(n956), .A2(G475), .ZN(n1061) );
XNOR2_X1 U764 ( .A(G104), .B(n1062), .ZN(G6) );
NOR2_X1 U765 ( .A1(n1046), .A2(n1063), .ZN(G57) );
XOR2_X1 U766 ( .A(n1064), .B(n1065), .Z(n1063) );
XOR2_X1 U767 ( .A(G101), .B(n1066), .Z(n1065) );
AND2_X1 U768 ( .A1(G472), .A2(n1051), .ZN(n1066) );
NOR2_X1 U769 ( .A1(n1046), .A2(n1067), .ZN(G54) );
XOR2_X1 U770 ( .A(n1068), .B(n1069), .Z(n1067) );
AND2_X1 U771 ( .A1(G469), .A2(n1051), .ZN(n1069) );
INV_X1 U772 ( .A(n1070), .ZN(n1051) );
NAND2_X1 U773 ( .A1(n1071), .A2(KEYINPUT14), .ZN(n1068) );
XOR2_X1 U774 ( .A(n1072), .B(n1073), .Z(n1071) );
XOR2_X1 U775 ( .A(n1074), .B(n1075), .Z(n1073) );
XOR2_X1 U776 ( .A(n1028), .B(n1076), .Z(n1075) );
NAND2_X1 U777 ( .A1(KEYINPUT16), .A2(n1077), .ZN(n1074) );
XOR2_X1 U778 ( .A(n1078), .B(n1042), .Z(n1072) );
NOR2_X1 U779 ( .A1(n1046), .A2(n1079), .ZN(G51) );
XOR2_X1 U780 ( .A(n1080), .B(n1081), .Z(n1079) );
XOR2_X1 U781 ( .A(n1030), .B(n1082), .Z(n1080) );
NOR2_X1 U782 ( .A1(n1003), .A2(n1070), .ZN(n1082) );
NAND2_X1 U783 ( .A1(G902), .A2(n956), .ZN(n1070) );
NAND4_X1 U784 ( .A1(n1044), .A2(n1017), .A3(n1083), .A4(n1019), .ZN(n956) );
XNOR2_X1 U785 ( .A(KEYINPUT59), .B(n1045), .ZN(n1083) );
AND4_X1 U786 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1087), .ZN(n1017) );
NOR4_X1 U787 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1087) );
INV_X1 U788 ( .A(n1092), .ZN(n1091) );
INV_X1 U789 ( .A(n1093), .ZN(n1090) );
AND4_X1 U790 ( .A1(n1062), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1044) );
AND4_X1 U791 ( .A1(n1097), .A2(n1098), .A3(n1099), .A4(n1100), .ZN(n1096) );
NAND2_X1 U792 ( .A1(n951), .A2(n952), .ZN(n1095) );
AND4_X1 U793 ( .A1(n979), .A2(n965), .A3(n1101), .A4(n1102), .ZN(n952) );
INV_X1 U794 ( .A(n1103), .ZN(n951) );
NAND3_X1 U795 ( .A1(n978), .A2(n965), .A3(n1104), .ZN(n1062) );
NOR2_X1 U796 ( .A1(n971), .A2(G952), .ZN(n1046) );
XNOR2_X1 U797 ( .A(n1105), .B(n1086), .ZN(G48) );
NAND3_X1 U798 ( .A1(n978), .A2(n1106), .A3(n1107), .ZN(n1086) );
NOR2_X1 U799 ( .A1(KEYINPUT42), .A2(n1108), .ZN(n1105) );
XOR2_X1 U800 ( .A(KEYINPUT46), .B(G146), .Z(n1108) );
XOR2_X1 U801 ( .A(n1084), .B(n1109), .Z(G45) );
NOR2_X1 U802 ( .A1(G143), .A2(KEYINPUT15), .ZN(n1109) );
NAND4_X1 U803 ( .A1(n1110), .A2(n1106), .A3(n1111), .A4(n1112), .ZN(n1084) );
XOR2_X1 U804 ( .A(n1028), .B(n1085), .Z(G42) );
NAND4_X1 U805 ( .A1(n990), .A2(n978), .A3(n973), .A4(n1113), .ZN(n1085) );
NAND2_X1 U806 ( .A1(n1114), .A2(n1115), .ZN(G39) );
NAND2_X1 U807 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
NAND2_X1 U808 ( .A1(n1118), .A2(G137), .ZN(n1114) );
NAND2_X1 U809 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U810 ( .A1(KEYINPUT18), .A2(n1089), .ZN(n1120) );
OR2_X1 U811 ( .A1(n1116), .A2(KEYINPUT18), .ZN(n1119) );
AND2_X1 U812 ( .A1(KEYINPUT17), .A2(n1089), .ZN(n1116) );
AND3_X1 U813 ( .A1(n969), .A2(n973), .A3(n1107), .ZN(n1089) );
XOR2_X1 U814 ( .A(n1019), .B(n1121), .Z(G36) );
XOR2_X1 U815 ( .A(KEYINPUT34), .B(G134), .Z(n1121) );
NAND3_X1 U816 ( .A1(n1110), .A2(n979), .A3(n973), .ZN(n1019) );
XOR2_X1 U817 ( .A(n1122), .B(n1092), .Z(G33) );
NAND3_X1 U818 ( .A1(n973), .A2(n1110), .A3(n978), .ZN(n1092) );
AND2_X1 U819 ( .A1(n989), .A2(n1113), .ZN(n1110) );
NOR2_X1 U820 ( .A1(n1123), .A2(n962), .ZN(n973) );
INV_X1 U821 ( .A(n1124), .ZN(n1123) );
XOR2_X1 U822 ( .A(n1088), .B(n1125), .Z(G30) );
NOR2_X1 U823 ( .A1(KEYINPUT54), .A2(n1126), .ZN(n1125) );
AND3_X1 U824 ( .A1(n979), .A2(n1106), .A3(n1107), .ZN(n1088) );
AND3_X1 U825 ( .A1(n1113), .A2(n1127), .A3(n1128), .ZN(n1107) );
NOR2_X1 U826 ( .A1(n984), .A2(n1129), .ZN(n1113) );
XNOR2_X1 U827 ( .A(G101), .B(n1094), .ZN(G3) );
NAND3_X1 U828 ( .A1(n969), .A2(n989), .A3(n1104), .ZN(n1094) );
XOR2_X1 U829 ( .A(n1030), .B(n1093), .Z(G27) );
NAND4_X1 U830 ( .A1(n990), .A2(n978), .A3(n1130), .A4(n967), .ZN(n1093) );
NOR2_X1 U831 ( .A1(n1129), .A2(n959), .ZN(n1130) );
AND2_X1 U832 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NAND2_X1 U833 ( .A1(n1133), .A2(n1134), .ZN(n1131) );
XNOR2_X1 U834 ( .A(G900), .B(KEYINPUT49), .ZN(n1133) );
XNOR2_X1 U835 ( .A(G122), .B(n1100), .ZN(G24) );
NAND4_X1 U836 ( .A1(n1135), .A2(n965), .A3(n1111), .A4(n1112), .ZN(n1100) );
NOR2_X1 U837 ( .A1(n1010), .A2(n1128), .ZN(n965) );
NAND3_X1 U838 ( .A1(n1136), .A2(n1137), .A3(n1138), .ZN(G21) );
OR2_X1 U839 ( .A1(n1099), .A2(G119), .ZN(n1138) );
NAND2_X1 U840 ( .A1(n1139), .A2(n1140), .ZN(n1137) );
INV_X1 U841 ( .A(KEYINPUT40), .ZN(n1140) );
NAND2_X1 U842 ( .A1(G119), .A2(n1141), .ZN(n1139) );
XNOR2_X1 U843 ( .A(KEYINPUT53), .B(n1099), .ZN(n1141) );
NAND2_X1 U844 ( .A1(KEYINPUT40), .A2(n1142), .ZN(n1136) );
NAND2_X1 U845 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
OR2_X1 U846 ( .A1(n1099), .A2(KEYINPUT53), .ZN(n1144) );
NAND3_X1 U847 ( .A1(G119), .A2(n1099), .A3(KEYINPUT53), .ZN(n1143) );
NAND4_X1 U848 ( .A1(n1128), .A2(n969), .A3(n1135), .A4(n1127), .ZN(n1099) );
XNOR2_X1 U849 ( .A(G116), .B(n1098), .ZN(G18) );
NAND3_X1 U850 ( .A1(n989), .A2(n979), .A3(n1135), .ZN(n1098) );
AND3_X1 U851 ( .A1(n1106), .A2(n1102), .A3(n967), .ZN(n1135) );
INV_X1 U852 ( .A(n959), .ZN(n1106) );
XOR2_X1 U853 ( .A(n1103), .B(KEYINPUT62), .Z(n959) );
NOR2_X1 U854 ( .A1(n1111), .A2(n1145), .ZN(n979) );
XNOR2_X1 U855 ( .A(G113), .B(n1097), .ZN(G15) );
NAND4_X1 U856 ( .A1(n978), .A2(n967), .A3(n1146), .A4(n989), .ZN(n1097) );
AND2_X1 U857 ( .A1(n1127), .A2(n1147), .ZN(n989) );
XOR2_X1 U858 ( .A(n1010), .B(KEYINPUT29), .Z(n1127) );
NOR2_X1 U859 ( .A1(n1148), .A2(n1103), .ZN(n1146) );
NOR2_X1 U860 ( .A1(n1006), .A2(n986), .ZN(n967) );
INV_X1 U861 ( .A(n987), .ZN(n1006) );
AND2_X1 U862 ( .A1(n1145), .A2(n1111), .ZN(n978) );
INV_X1 U863 ( .A(n1112), .ZN(n1145) );
XOR2_X1 U864 ( .A(n1045), .B(n1149), .Z(G12) );
XOR2_X1 U865 ( .A(n1077), .B(KEYINPUT12), .Z(n1149) );
NAND3_X1 U866 ( .A1(n1104), .A2(n969), .A3(n990), .ZN(n1045) );
NOR2_X1 U867 ( .A1(n1147), .A2(n1010), .ZN(n990) );
XNOR2_X1 U868 ( .A(n1150), .B(G472), .ZN(n1010) );
NAND2_X1 U869 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
XOR2_X1 U870 ( .A(n1153), .B(n1064), .Z(n1151) );
XNOR2_X1 U871 ( .A(n1154), .B(n1155), .ZN(n1064) );
XOR2_X1 U872 ( .A(n1078), .B(n1156), .Z(n1154) );
AND3_X1 U873 ( .A1(G210), .A2(n971), .A3(n1157), .ZN(n1156) );
XNOR2_X1 U874 ( .A(n1158), .B(n1025), .ZN(n1078) );
XNOR2_X1 U875 ( .A(n1159), .B(n1160), .ZN(n1025) );
NOR2_X1 U876 ( .A1(G101), .A2(KEYINPUT30), .ZN(n1153) );
INV_X1 U877 ( .A(n1128), .ZN(n1147) );
XNOR2_X1 U878 ( .A(n1000), .B(n1161), .ZN(n1128) );
NOR2_X1 U879 ( .A1(n999), .A2(KEYINPUT27), .ZN(n1161) );
AND2_X1 U880 ( .A1(G217), .A2(n1162), .ZN(n999) );
NOR2_X1 U881 ( .A1(n1050), .A2(G902), .ZN(n1000) );
XNOR2_X1 U882 ( .A(n1163), .B(n1164), .ZN(n1050) );
XOR2_X1 U883 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U884 ( .A(G119), .B(G110), .Z(n1166) );
XOR2_X1 U885 ( .A(KEYINPUT19), .B(G146), .Z(n1165) );
XOR2_X1 U886 ( .A(n1167), .B(n1168), .Z(n1163) );
XOR2_X1 U887 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U888 ( .A1(KEYINPUT37), .A2(n1126), .ZN(n1170) );
AND3_X1 U889 ( .A1(n1171), .A2(G234), .A3(G221), .ZN(n1169) );
XOR2_X1 U890 ( .A(KEYINPUT35), .B(n971), .Z(n1171) );
XNOR2_X1 U891 ( .A(n1172), .B(n1173), .ZN(n1167) );
NOR2_X1 U892 ( .A1(G137), .A2(KEYINPUT52), .ZN(n1173) );
NOR2_X1 U893 ( .A1(n1112), .A2(n1111), .ZN(n969) );
XNOR2_X1 U894 ( .A(n1174), .B(n1175), .ZN(n1111) );
NOR2_X1 U895 ( .A1(KEYINPUT4), .A2(G475), .ZN(n1175) );
XNOR2_X1 U896 ( .A(n1007), .B(KEYINPUT5), .ZN(n1174) );
NOR2_X1 U897 ( .A1(n1060), .A2(G902), .ZN(n1007) );
XNOR2_X1 U898 ( .A(n1176), .B(n1177), .ZN(n1060) );
XNOR2_X1 U899 ( .A(n1178), .B(n1179), .ZN(n1177) );
NAND3_X1 U900 ( .A1(n1180), .A2(n1181), .A3(n1182), .ZN(n1178) );
NAND2_X1 U901 ( .A1(G104), .A2(n1183), .ZN(n1182) );
OR3_X1 U902 ( .A1(n1183), .A2(G104), .A3(n1184), .ZN(n1181) );
INV_X1 U903 ( .A(KEYINPUT3), .ZN(n1184) );
NAND2_X1 U904 ( .A1(KEYINPUT55), .A2(n1185), .ZN(n1183) );
OR2_X1 U905 ( .A1(n1185), .A2(KEYINPUT3), .ZN(n1180) );
XNOR2_X1 U906 ( .A(n1186), .B(G122), .ZN(n1185) );
NAND2_X1 U907 ( .A1(KEYINPUT56), .A2(G113), .ZN(n1186) );
XOR2_X1 U908 ( .A(n1187), .B(n1188), .Z(n1176) );
XOR2_X1 U909 ( .A(n1122), .B(n1189), .Z(n1188) );
NAND2_X1 U910 ( .A1(KEYINPUT48), .A2(n1172), .ZN(n1189) );
XOR2_X1 U911 ( .A(n1030), .B(n1028), .Z(n1172) );
INV_X1 U912 ( .A(G125), .ZN(n1030) );
INV_X1 U913 ( .A(G131), .ZN(n1122) );
NAND4_X1 U914 ( .A1(KEYINPUT6), .A2(G214), .A3(n1157), .A4(n971), .ZN(n1187) );
NAND2_X1 U915 ( .A1(n1190), .A2(n1191), .ZN(n1112) );
NAND2_X1 U916 ( .A1(n1192), .A2(n1009), .ZN(n1191) );
XOR2_X1 U917 ( .A(KEYINPUT0), .B(n1008), .Z(n1192) );
XOR2_X1 U918 ( .A(KEYINPUT22), .B(n1193), .Z(n1190) );
NOR2_X1 U919 ( .A1(n1008), .A2(n1194), .ZN(n1193) );
XOR2_X1 U920 ( .A(KEYINPUT50), .B(n1009), .Z(n1194) );
XOR2_X1 U921 ( .A(G478), .B(KEYINPUT21), .Z(n1009) );
NOR2_X1 U922 ( .A1(n1056), .A2(G902), .ZN(n1008) );
AND2_X1 U923 ( .A1(n1195), .A2(n1196), .ZN(n1056) );
NAND2_X1 U924 ( .A1(n1197), .A2(n1198), .ZN(n1196) );
NAND3_X1 U925 ( .A1(n1199), .A2(G217), .A3(G234), .ZN(n1198) );
INV_X1 U926 ( .A(n1200), .ZN(n1197) );
NAND4_X1 U927 ( .A1(n1199), .A2(G217), .A3(G234), .A4(n1200), .ZN(n1195) );
NAND3_X1 U928 ( .A1(n1201), .A2(n1202), .A3(n1203), .ZN(n1200) );
NAND2_X1 U929 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
OR3_X1 U930 ( .A1(n1205), .A2(n1204), .A3(n1206), .ZN(n1202) );
INV_X1 U931 ( .A(KEYINPUT61), .ZN(n1206) );
XNOR2_X1 U932 ( .A(n948), .B(n1207), .ZN(n1204) );
XOR2_X1 U933 ( .A(G122), .B(G116), .Z(n1207) );
INV_X1 U934 ( .A(G107), .ZN(n948) );
NAND2_X1 U935 ( .A1(KEYINPUT8), .A2(n1208), .ZN(n1205) );
OR2_X1 U936 ( .A1(n1208), .A2(KEYINPUT61), .ZN(n1201) );
XNOR2_X1 U937 ( .A(n1209), .B(n1210), .ZN(n1208) );
XOR2_X1 U938 ( .A(G143), .B(G134), .Z(n1210) );
NAND2_X1 U939 ( .A1(KEYINPUT33), .A2(n1126), .ZN(n1209) );
XOR2_X1 U940 ( .A(n971), .B(KEYINPUT2), .Z(n1199) );
NOR3_X1 U941 ( .A1(n984), .A2(n1148), .A3(n1103), .ZN(n1104) );
NAND2_X1 U942 ( .A1(n962), .A2(n1124), .ZN(n1103) );
XNOR2_X1 U943 ( .A(n964), .B(KEYINPUT44), .ZN(n1124) );
AND2_X1 U944 ( .A1(G214), .A2(n1211), .ZN(n964) );
XNOR2_X1 U945 ( .A(n1212), .B(n1003), .ZN(n962) );
NAND2_X1 U946 ( .A1(G210), .A2(n1211), .ZN(n1003) );
NAND2_X1 U947 ( .A1(n1157), .A2(n1152), .ZN(n1211) );
INV_X1 U948 ( .A(G237), .ZN(n1157) );
XOR2_X1 U949 ( .A(n1002), .B(KEYINPUT32), .Z(n1212) );
NAND2_X1 U950 ( .A1(n1213), .A2(n1152), .ZN(n1002) );
XNOR2_X1 U951 ( .A(n1081), .B(n1214), .ZN(n1213) );
XOR2_X1 U952 ( .A(KEYINPUT36), .B(n1215), .Z(n1214) );
NOR2_X1 U953 ( .A1(G125), .A2(KEYINPUT13), .ZN(n1215) );
XNOR2_X1 U954 ( .A(n1216), .B(n1217), .ZN(n1081) );
INV_X1 U955 ( .A(n1041), .ZN(n1217) );
XOR2_X1 U956 ( .A(n1218), .B(n1219), .Z(n1041) );
XOR2_X1 U957 ( .A(KEYINPUT25), .B(G122), .Z(n1219) );
XOR2_X1 U958 ( .A(n1077), .B(n1155), .Z(n1218) );
XNOR2_X1 U959 ( .A(n1220), .B(n1221), .ZN(n1155) );
XOR2_X1 U960 ( .A(KEYINPUT60), .B(G119), .Z(n1221) );
XNOR2_X1 U961 ( .A(G113), .B(G116), .ZN(n1220) );
XOR2_X1 U962 ( .A(n1222), .B(n1223), .Z(n1216) );
NOR2_X1 U963 ( .A1(G953), .A2(n1037), .ZN(n1223) );
INV_X1 U964 ( .A(G224), .ZN(n1037) );
INV_X1 U965 ( .A(n1102), .ZN(n1148) );
NAND2_X1 U966 ( .A1(n1224), .A2(n1132), .ZN(n1102) );
NAND3_X1 U967 ( .A1(n966), .A2(n971), .A3(G952), .ZN(n1132) );
NAND2_X1 U968 ( .A1(n1134), .A2(n1038), .ZN(n1224) );
INV_X1 U969 ( .A(G898), .ZN(n1038) );
AND3_X1 U970 ( .A1(G953), .A2(n966), .A3(G902), .ZN(n1134) );
NAND2_X1 U971 ( .A1(G237), .A2(G234), .ZN(n966) );
INV_X1 U972 ( .A(n1101), .ZN(n984) );
NOR2_X1 U973 ( .A1(n987), .A2(n986), .ZN(n1101) );
AND2_X1 U974 ( .A1(G221), .A2(n1162), .ZN(n986) );
NAND2_X1 U975 ( .A1(G234), .A2(n1152), .ZN(n1162) );
XOR2_X1 U976 ( .A(n1225), .B(n1226), .Z(n987) );
XOR2_X1 U977 ( .A(KEYINPUT23), .B(G469), .Z(n1226) );
NAND2_X1 U978 ( .A1(n1227), .A2(n1228), .ZN(n1225) );
XOR2_X1 U979 ( .A(n1229), .B(n1230), .Z(n1228) );
XOR2_X1 U980 ( .A(n1231), .B(n1222), .Z(n1230) );
XOR2_X1 U981 ( .A(n1159), .B(n1042), .Z(n1222) );
XOR2_X1 U982 ( .A(G101), .B(n1232), .Z(n1042) );
XOR2_X1 U983 ( .A(G107), .B(G104), .Z(n1232) );
XOR2_X1 U984 ( .A(n1126), .B(n1179), .Z(n1159) );
XOR2_X1 U985 ( .A(G143), .B(G146), .Z(n1179) );
INV_X1 U986 ( .A(G128), .ZN(n1126) );
NAND2_X1 U987 ( .A1(KEYINPUT10), .A2(n1233), .ZN(n1231) );
XOR2_X1 U988 ( .A(n1158), .B(n1160), .Z(n1233) );
XOR2_X1 U989 ( .A(G131), .B(G134), .Z(n1160) );
NOR2_X1 U990 ( .A1(KEYINPUT1), .A2(n1117), .ZN(n1158) );
INV_X1 U991 ( .A(G137), .ZN(n1117) );
XNOR2_X1 U992 ( .A(n1076), .B(n1234), .ZN(n1229) );
NAND2_X1 U993 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND2_X1 U994 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
NAND2_X1 U995 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
NAND2_X1 U996 ( .A1(n1241), .A2(n1242), .ZN(n1239) );
XOR2_X1 U997 ( .A(KEYINPUT47), .B(G140), .Z(n1241) );
XOR2_X1 U998 ( .A(KEYINPUT9), .B(G110), .Z(n1237) );
NAND2_X1 U999 ( .A1(n1243), .A2(n1244), .ZN(n1235) );
NAND2_X1 U1000 ( .A1(n1245), .A2(n1242), .ZN(n1244) );
INV_X1 U1001 ( .A(KEYINPUT39), .ZN(n1242) );
NAND2_X1 U1002 ( .A1(n1246), .A2(n1240), .ZN(n1245) );
INV_X1 U1003 ( .A(KEYINPUT41), .ZN(n1240) );
XOR2_X1 U1004 ( .A(KEYINPUT9), .B(n1077), .Z(n1246) );
INV_X1 U1005 ( .A(G110), .ZN(n1077) );
XOR2_X1 U1006 ( .A(KEYINPUT47), .B(n1028), .Z(n1243) );
INV_X1 U1007 ( .A(G140), .ZN(n1028) );
AND2_X1 U1008 ( .A1(G227), .A2(n971), .ZN(n1076) );
INV_X1 U1009 ( .A(G953), .ZN(n971) );
XOR2_X1 U1010 ( .A(n1152), .B(KEYINPUT24), .Z(n1227) );
INV_X1 U1011 ( .A(G902), .ZN(n1152) );
endmodule


