//Key = 1011100110010111110110101110100001000010100100110101100100101011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296;

NAND2_X1 U728 ( .A1(n994), .A2(n995), .ZN(G9) );
NAND2_X1 U729 ( .A1(G107), .A2(n996), .ZN(n995) );
XOR2_X1 U730 ( .A(KEYINPUT51), .B(n997), .Z(n994) );
NOR2_X1 U731 ( .A1(G107), .A2(n996), .ZN(n997) );
NOR2_X1 U732 ( .A1(n998), .A2(n999), .ZN(G75) );
XOR2_X1 U733 ( .A(n1000), .B(KEYINPUT0), .Z(n999) );
NAND3_X1 U734 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n1000) );
NAND2_X1 U735 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NAND2_X1 U736 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NAND3_X1 U737 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NAND2_X1 U738 ( .A1(n1011), .A2(n1012), .ZN(n1009) );
NAND2_X1 U739 ( .A1(n1013), .A2(n1014), .ZN(n1012) );
OR2_X1 U740 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U741 ( .A1(n1017), .A2(n1018), .ZN(n1011) );
NAND2_X1 U742 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
NAND3_X1 U743 ( .A1(n1013), .A2(n1021), .A3(n1017), .ZN(n1006) );
NAND2_X1 U744 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U745 ( .A1(n1010), .A2(n1024), .ZN(n1023) );
NAND2_X1 U746 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
NAND2_X1 U747 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
XOR2_X1 U748 ( .A(KEYINPUT14), .B(n1029), .Z(n1028) );
NAND2_X1 U749 ( .A1(n1008), .A2(n1030), .ZN(n1022) );
NAND2_X1 U750 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
OR2_X1 U751 ( .A1(n1033), .A2(n1034), .ZN(n1032) );
INV_X1 U752 ( .A(n1035), .ZN(n1004) );
INV_X1 U753 ( .A(n1036), .ZN(n1001) );
NOR2_X1 U754 ( .A1(G952), .A2(n1036), .ZN(n998) );
NAND2_X1 U755 ( .A1(n1037), .A2(n1038), .ZN(n1036) );
NAND4_X1 U756 ( .A1(n1039), .A2(n1008), .A3(n1040), .A4(n1041), .ZN(n1038) );
NOR4_X1 U757 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1041) );
XNOR2_X1 U758 ( .A(n1046), .B(n1047), .ZN(n1044) );
XNOR2_X1 U759 ( .A(n1048), .B(KEYINPUT63), .ZN(n1046) );
XOR2_X1 U760 ( .A(n1049), .B(n1050), .Z(n1043) );
XNOR2_X1 U761 ( .A(KEYINPUT10), .B(n1051), .ZN(n1050) );
NAND2_X1 U762 ( .A1(n1052), .A2(n1053), .ZN(n1049) );
XOR2_X1 U763 ( .A(KEYINPUT34), .B(KEYINPUT22), .Z(n1052) );
XNOR2_X1 U764 ( .A(n1054), .B(G475), .ZN(n1040) );
XNOR2_X1 U765 ( .A(n1055), .B(KEYINPUT48), .ZN(n1039) );
XOR2_X1 U766 ( .A(n1056), .B(n1057), .Z(G72) );
XOR2_X1 U767 ( .A(n1058), .B(n1059), .Z(n1057) );
NOR2_X1 U768 ( .A1(n1060), .A2(G953), .ZN(n1059) );
NOR3_X1 U769 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NOR2_X1 U770 ( .A1(n1064), .A2(n1065), .ZN(n1058) );
XOR2_X1 U771 ( .A(n1066), .B(n1067), .Z(n1065) );
XOR2_X1 U772 ( .A(n1068), .B(n1069), .Z(n1067) );
NOR2_X1 U773 ( .A1(KEYINPUT30), .A2(n1070), .ZN(n1068) );
XOR2_X1 U774 ( .A(n1071), .B(n1072), .Z(n1066) );
NOR2_X1 U775 ( .A1(KEYINPUT9), .A2(n1073), .ZN(n1072) );
XNOR2_X1 U776 ( .A(G125), .B(G140), .ZN(n1073) );
XNOR2_X1 U777 ( .A(G131), .B(KEYINPUT37), .ZN(n1071) );
NOR2_X1 U778 ( .A1(n1074), .A2(n1075), .ZN(n1056) );
INV_X1 U779 ( .A(n1076), .ZN(n1075) );
AND2_X1 U780 ( .A1(G227), .A2(G900), .ZN(n1074) );
XOR2_X1 U781 ( .A(n1077), .B(n1078), .Z(G69) );
XOR2_X1 U782 ( .A(n1079), .B(n1080), .Z(n1078) );
NAND2_X1 U783 ( .A1(n1076), .A2(n1081), .ZN(n1080) );
NAND2_X1 U784 ( .A1(G898), .A2(G224), .ZN(n1081) );
XOR2_X1 U785 ( .A(G953), .B(KEYINPUT18), .Z(n1076) );
NAND2_X1 U786 ( .A1(n1082), .A2(n1083), .ZN(n1079) );
NAND2_X1 U787 ( .A1(G953), .A2(n1084), .ZN(n1083) );
XOR2_X1 U788 ( .A(n1085), .B(n1086), .Z(n1082) );
NAND2_X1 U789 ( .A1(n1087), .A2(KEYINPUT55), .ZN(n1085) );
XOR2_X1 U790 ( .A(n1088), .B(KEYINPUT17), .Z(n1087) );
AND2_X1 U791 ( .A1(n1089), .A2(n1037), .ZN(n1077) );
NOR3_X1 U792 ( .A1(n1090), .A2(n1091), .A3(n1092), .ZN(G66) );
AND3_X1 U793 ( .A1(KEYINPUT29), .A2(G953), .A3(G952), .ZN(n1092) );
NOR2_X1 U794 ( .A1(KEYINPUT29), .A2(n1093), .ZN(n1091) );
INV_X1 U795 ( .A(n1094), .ZN(n1093) );
XNOR2_X1 U796 ( .A(n1095), .B(n1096), .ZN(n1090) );
NOR2_X1 U797 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U798 ( .A1(n1094), .A2(n1099), .ZN(G63) );
XNOR2_X1 U799 ( .A(n1100), .B(n1101), .ZN(n1099) );
NOR2_X1 U800 ( .A1(n1102), .A2(n1098), .ZN(n1101) );
NOR2_X1 U801 ( .A1(n1094), .A2(n1103), .ZN(G60) );
NOR3_X1 U802 ( .A1(n1054), .A2(n1104), .A3(n1105), .ZN(n1103) );
NOR3_X1 U803 ( .A1(n1106), .A2(n1107), .A3(n1098), .ZN(n1105) );
INV_X1 U804 ( .A(n1108), .ZN(n1106) );
NOR2_X1 U805 ( .A1(n1109), .A2(n1108), .ZN(n1104) );
NOR2_X1 U806 ( .A1(n1003), .A2(n1107), .ZN(n1109) );
XNOR2_X1 U807 ( .A(G104), .B(n1110), .ZN(G6) );
NOR2_X1 U808 ( .A1(n1094), .A2(n1111), .ZN(G57) );
XOR2_X1 U809 ( .A(n1112), .B(n1113), .Z(n1111) );
XNOR2_X1 U810 ( .A(n1114), .B(n1115), .ZN(n1113) );
XOR2_X1 U811 ( .A(n1116), .B(n1117), .Z(n1112) );
NOR2_X1 U812 ( .A1(n1051), .A2(n1098), .ZN(n1117) );
NAND2_X1 U813 ( .A1(KEYINPUT20), .A2(n1118), .ZN(n1116) );
NOR3_X1 U814 ( .A1(n1094), .A2(n1119), .A3(n1120), .ZN(G54) );
NOR2_X1 U815 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
XOR2_X1 U816 ( .A(n1123), .B(KEYINPUT57), .Z(n1122) );
INV_X1 U817 ( .A(n1124), .ZN(n1121) );
NOR2_X1 U818 ( .A1(n1124), .A2(n1125), .ZN(n1119) );
XOR2_X1 U819 ( .A(n1123), .B(KEYINPUT60), .Z(n1125) );
XOR2_X1 U820 ( .A(n1126), .B(n1127), .Z(n1123) );
XOR2_X1 U821 ( .A(KEYINPUT19), .B(n1128), .Z(n1127) );
NOR2_X1 U822 ( .A1(n1098), .A2(n1129), .ZN(n1128) );
XOR2_X1 U823 ( .A(KEYINPUT33), .B(G469), .Z(n1129) );
XOR2_X1 U824 ( .A(n1130), .B(n1131), .Z(n1126) );
NAND2_X1 U825 ( .A1(KEYINPUT47), .A2(n1132), .ZN(n1130) );
XNOR2_X1 U826 ( .A(n1133), .B(n1134), .ZN(n1124) );
XNOR2_X1 U827 ( .A(G140), .B(n1135), .ZN(n1134) );
NOR2_X1 U828 ( .A1(n1094), .A2(n1136), .ZN(G51) );
XOR2_X1 U829 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U830 ( .A1(n1047), .A2(n1098), .ZN(n1138) );
OR2_X1 U831 ( .A1(n1139), .A2(n1003), .ZN(n1098) );
NOR4_X1 U832 ( .A1(n1140), .A2(n1089), .A3(n1061), .A4(n1063), .ZN(n1003) );
NAND4_X1 U833 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1063) );
NAND2_X1 U834 ( .A1(n1145), .A2(n1146), .ZN(n1061) );
NAND2_X1 U835 ( .A1(n1010), .A2(n1147), .ZN(n1146) );
NAND2_X1 U836 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NAND2_X1 U837 ( .A1(n1150), .A2(n1016), .ZN(n1149) );
NAND2_X1 U838 ( .A1(n1151), .A2(n1017), .ZN(n1148) );
NAND2_X1 U839 ( .A1(n1152), .A2(n1153), .ZN(n1145) );
NAND4_X1 U840 ( .A1(n1154), .A2(n996), .A3(n1155), .A4(n1156), .ZN(n1089) );
NOR4_X1 U841 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
NOR3_X1 U842 ( .A1(n1020), .A2(n1161), .A3(n1162), .ZN(n1160) );
XNOR2_X1 U843 ( .A(n1017), .B(KEYINPUT54), .ZN(n1161) );
INV_X1 U844 ( .A(n1163), .ZN(n1159) );
AND2_X1 U845 ( .A1(n1164), .A2(n1110), .ZN(n1155) );
NAND3_X1 U846 ( .A1(n1013), .A2(n1165), .A3(n1015), .ZN(n1110) );
NAND3_X1 U847 ( .A1(n1013), .A2(n1165), .A3(n1016), .ZN(n996) );
XOR2_X1 U848 ( .A(n1062), .B(KEYINPUT61), .Z(n1140) );
NOR2_X1 U849 ( .A1(n1166), .A2(n1167), .ZN(n1137) );
XOR2_X1 U850 ( .A(n1168), .B(KEYINPUT16), .Z(n1167) );
NAND2_X1 U851 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
NOR2_X1 U852 ( .A1(n1170), .A2(n1169), .ZN(n1166) );
XOR2_X1 U853 ( .A(n1171), .B(n1172), .Z(n1169) );
NAND2_X1 U854 ( .A1(KEYINPUT52), .A2(n1173), .ZN(n1171) );
NOR2_X1 U855 ( .A1(n1037), .A2(G952), .ZN(n1094) );
XNOR2_X1 U856 ( .A(n1142), .B(n1174), .ZN(G48) );
NOR2_X1 U857 ( .A1(KEYINPUT42), .A2(n1175), .ZN(n1174) );
NAND3_X1 U858 ( .A1(n1015), .A2(n1176), .A3(n1151), .ZN(n1142) );
XOR2_X1 U859 ( .A(G143), .B(n1062), .Z(G45) );
AND4_X1 U860 ( .A1(n1150), .A2(n1176), .A3(n1177), .A4(n1055), .ZN(n1062) );
NOR3_X1 U861 ( .A1(n1025), .A2(n1178), .A3(n1020), .ZN(n1150) );
INV_X1 U862 ( .A(n1179), .ZN(n1020) );
XOR2_X1 U863 ( .A(G140), .B(n1180), .Z(G42) );
NOR2_X1 U864 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XNOR2_X1 U865 ( .A(n1153), .B(KEYINPUT53), .ZN(n1181) );
XNOR2_X1 U866 ( .A(G137), .B(n1183), .ZN(G39) );
NAND4_X1 U867 ( .A1(n1017), .A2(n1184), .A3(n1010), .A4(n1185), .ZN(n1183) );
NOR4_X1 U868 ( .A1(KEYINPUT50), .A2(n1178), .A3(n1186), .A4(n1187), .ZN(n1185) );
XNOR2_X1 U869 ( .A(KEYINPUT45), .B(n1025), .ZN(n1184) );
XNOR2_X1 U870 ( .A(G134), .B(n1188), .ZN(G36) );
NAND2_X1 U871 ( .A1(n1189), .A2(n1010), .ZN(n1188) );
XOR2_X1 U872 ( .A(n1190), .B(KEYINPUT62), .Z(n1189) );
NAND4_X1 U873 ( .A1(n1179), .A2(n1016), .A3(n1191), .A4(n1192), .ZN(n1190) );
XNOR2_X1 U874 ( .A(KEYINPUT36), .B(n1025), .ZN(n1191) );
XOR2_X1 U875 ( .A(n1141), .B(n1193), .Z(G33) );
NAND2_X1 U876 ( .A1(KEYINPUT26), .A2(G131), .ZN(n1193) );
NAND2_X1 U877 ( .A1(n1152), .A2(n1179), .ZN(n1141) );
INV_X1 U878 ( .A(n1182), .ZN(n1152) );
NAND4_X1 U879 ( .A1(n1010), .A2(n1015), .A3(n1194), .A4(n1192), .ZN(n1182) );
NOR2_X1 U880 ( .A1(n1033), .A2(n1042), .ZN(n1010) );
INV_X1 U881 ( .A(n1034), .ZN(n1042) );
XNOR2_X1 U882 ( .A(G128), .B(n1143), .ZN(G30) );
NAND3_X1 U883 ( .A1(n1016), .A2(n1176), .A3(n1151), .ZN(n1143) );
NOR4_X1 U884 ( .A1(n1025), .A2(n1187), .A3(n1186), .A4(n1178), .ZN(n1151) );
INV_X1 U885 ( .A(n1192), .ZN(n1178) );
XNOR2_X1 U886 ( .A(G101), .B(n1195), .ZN(G3) );
NAND2_X1 U887 ( .A1(n1179), .A2(n1196), .ZN(n1195) );
XNOR2_X1 U888 ( .A(G125), .B(n1144), .ZN(G27) );
NAND3_X1 U889 ( .A1(n1153), .A2(n1015), .A3(n1197), .ZN(n1144) );
AND3_X1 U890 ( .A1(n1008), .A2(n1192), .A3(n1176), .ZN(n1197) );
NAND2_X1 U891 ( .A1(n1035), .A2(n1198), .ZN(n1192) );
NAND3_X1 U892 ( .A1(G902), .A2(n1199), .A3(n1064), .ZN(n1198) );
NOR2_X1 U893 ( .A1(n1037), .A2(G900), .ZN(n1064) );
XNOR2_X1 U894 ( .A(G122), .B(n1163), .ZN(G24) );
NAND4_X1 U895 ( .A1(n1200), .A2(n1013), .A3(n1177), .A4(n1055), .ZN(n1163) );
AND2_X1 U896 ( .A1(n1187), .A2(n1201), .ZN(n1013) );
INV_X1 U897 ( .A(n1045), .ZN(n1187) );
XOR2_X1 U898 ( .A(n1164), .B(n1202), .Z(G21) );
NOR2_X1 U899 ( .A1(G119), .A2(KEYINPUT32), .ZN(n1202) );
NAND4_X1 U900 ( .A1(n1017), .A2(n1200), .A3(n1045), .A4(n1203), .ZN(n1164) );
XNOR2_X1 U901 ( .A(n1158), .B(n1204), .ZN(G18) );
NAND2_X1 U902 ( .A1(KEYINPUT3), .A2(G116), .ZN(n1204) );
AND3_X1 U903 ( .A1(n1200), .A2(n1016), .A3(n1179), .ZN(n1158) );
NOR2_X1 U904 ( .A1(n1205), .A2(n1206), .ZN(n1016) );
XNOR2_X1 U905 ( .A(n1207), .B(n1157), .ZN(G15) );
AND3_X1 U906 ( .A1(n1015), .A2(n1200), .A3(n1179), .ZN(n1157) );
NOR2_X1 U907 ( .A1(n1045), .A2(n1186), .ZN(n1179) );
AND3_X1 U908 ( .A1(n1176), .A2(n1208), .A3(n1008), .ZN(n1200) );
NOR2_X1 U909 ( .A1(n1029), .A2(n1027), .ZN(n1008) );
INV_X1 U910 ( .A(n1209), .ZN(n1027) );
AND2_X1 U911 ( .A1(n1206), .A2(n1177), .ZN(n1015) );
XNOR2_X1 U912 ( .A(n1205), .B(KEYINPUT38), .ZN(n1177) );
INV_X1 U913 ( .A(n1055), .ZN(n1206) );
XNOR2_X1 U914 ( .A(G110), .B(n1154), .ZN(G12) );
NAND2_X1 U915 ( .A1(n1153), .A2(n1196), .ZN(n1154) );
AND2_X1 U916 ( .A1(n1017), .A2(n1165), .ZN(n1196) );
INV_X1 U917 ( .A(n1162), .ZN(n1165) );
NAND3_X1 U918 ( .A1(n1194), .A2(n1208), .A3(n1176), .ZN(n1162) );
INV_X1 U919 ( .A(n1031), .ZN(n1176) );
NAND2_X1 U920 ( .A1(n1210), .A2(n1033), .ZN(n1031) );
NAND2_X1 U921 ( .A1(n1211), .A2(n1212), .ZN(n1033) );
NAND2_X1 U922 ( .A1(n1048), .A2(n1047), .ZN(n1212) );
XOR2_X1 U923 ( .A(KEYINPUT46), .B(n1213), .Z(n1211) );
NOR2_X1 U924 ( .A1(n1048), .A2(n1047), .ZN(n1213) );
NAND2_X1 U925 ( .A1(G210), .A2(n1214), .ZN(n1047) );
AND2_X1 U926 ( .A1(n1215), .A2(n1139), .ZN(n1048) );
XOR2_X1 U927 ( .A(n1170), .B(n1216), .Z(n1215) );
XOR2_X1 U928 ( .A(n1172), .B(n1217), .Z(n1216) );
NOR2_X1 U929 ( .A1(KEYINPUT6), .A2(n1218), .ZN(n1217) );
INV_X1 U930 ( .A(n1173), .ZN(n1218) );
XOR2_X1 U931 ( .A(G125), .B(n1219), .Z(n1173) );
AND2_X1 U932 ( .A1(G224), .A2(n1037), .ZN(n1172) );
XNOR2_X1 U933 ( .A(n1086), .B(n1088), .ZN(n1170) );
NAND3_X1 U934 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1088) );
OR2_X1 U935 ( .A1(n1223), .A2(KEYINPUT28), .ZN(n1222) );
NAND3_X1 U936 ( .A1(KEYINPUT28), .A2(n1223), .A3(G110), .ZN(n1221) );
NAND2_X1 U937 ( .A1(n1224), .A2(n1135), .ZN(n1220) );
NAND2_X1 U938 ( .A1(KEYINPUT28), .A2(n1225), .ZN(n1224) );
XNOR2_X1 U939 ( .A(KEYINPUT40), .B(n1223), .ZN(n1225) );
INV_X1 U940 ( .A(G122), .ZN(n1223) );
XOR2_X1 U941 ( .A(n1226), .B(n1227), .Z(n1086) );
XOR2_X1 U942 ( .A(n1228), .B(n1229), .Z(n1227) );
XNOR2_X1 U943 ( .A(G113), .B(G119), .ZN(n1226) );
XNOR2_X1 U944 ( .A(KEYINPUT58), .B(n1034), .ZN(n1210) );
NAND2_X1 U945 ( .A1(G214), .A2(n1214), .ZN(n1034) );
NAND2_X1 U946 ( .A1(n1230), .A2(n1139), .ZN(n1214) );
INV_X1 U947 ( .A(G237), .ZN(n1230) );
NAND2_X1 U948 ( .A1(n1035), .A2(n1231), .ZN(n1208) );
NAND4_X1 U949 ( .A1(G953), .A2(G902), .A3(n1199), .A4(n1084), .ZN(n1231) );
INV_X1 U950 ( .A(G898), .ZN(n1084) );
NAND3_X1 U951 ( .A1(n1199), .A2(n1037), .A3(G952), .ZN(n1035) );
NAND2_X1 U952 ( .A1(G237), .A2(G234), .ZN(n1199) );
INV_X1 U953 ( .A(n1025), .ZN(n1194) );
NAND2_X1 U954 ( .A1(n1029), .A2(n1209), .ZN(n1025) );
NAND2_X1 U955 ( .A1(G221), .A2(n1232), .ZN(n1209) );
XNOR2_X1 U956 ( .A(n1233), .B(G469), .ZN(n1029) );
NAND2_X1 U957 ( .A1(n1234), .A2(n1139), .ZN(n1233) );
XOR2_X1 U958 ( .A(n1235), .B(n1131), .Z(n1234) );
XNOR2_X1 U959 ( .A(n1236), .B(n1069), .ZN(n1131) );
XNOR2_X1 U960 ( .A(n1237), .B(n1238), .ZN(n1069) );
NOR2_X1 U961 ( .A1(KEYINPUT44), .A2(n1239), .ZN(n1238) );
XNOR2_X1 U962 ( .A(G143), .B(KEYINPUT43), .ZN(n1239) );
XNOR2_X1 U963 ( .A(n1240), .B(n1241), .ZN(n1236) );
INV_X1 U964 ( .A(G101), .ZN(n1241) );
NAND2_X1 U965 ( .A1(n1242), .A2(KEYINPUT25), .ZN(n1240) );
XNOR2_X1 U966 ( .A(n1228), .B(KEYINPUT2), .ZN(n1242) );
XOR2_X1 U967 ( .A(G104), .B(G107), .Z(n1228) );
XNOR2_X1 U968 ( .A(n1132), .B(n1243), .ZN(n1235) );
NOR2_X1 U969 ( .A1(KEYINPUT39), .A2(n1244), .ZN(n1243) );
XOR2_X1 U970 ( .A(n1133), .B(n1245), .Z(n1244) );
NOR2_X1 U971 ( .A1(KEYINPUT41), .A2(n1246), .ZN(n1245) );
XNOR2_X1 U972 ( .A(n1135), .B(n1247), .ZN(n1246) );
NOR2_X1 U973 ( .A1(G140), .A2(KEYINPUT27), .ZN(n1247) );
INV_X1 U974 ( .A(G110), .ZN(n1135) );
NAND2_X1 U975 ( .A1(G227), .A2(n1037), .ZN(n1133) );
NOR2_X1 U976 ( .A1(n1055), .A2(n1205), .ZN(n1017) );
XOR2_X1 U977 ( .A(n1248), .B(n1054), .Z(n1205) );
NOR2_X1 U978 ( .A1(n1108), .A2(G902), .ZN(n1054) );
XNOR2_X1 U979 ( .A(n1249), .B(n1250), .ZN(n1108) );
XOR2_X1 U980 ( .A(n1251), .B(n1252), .Z(n1250) );
XNOR2_X1 U981 ( .A(G131), .B(n1207), .ZN(n1252) );
XOR2_X1 U982 ( .A(KEYINPUT13), .B(G140), .Z(n1251) );
XOR2_X1 U983 ( .A(n1253), .B(n1254), .Z(n1249) );
XOR2_X1 U984 ( .A(n1255), .B(n1256), .Z(n1254) );
XNOR2_X1 U985 ( .A(n1257), .B(n1258), .ZN(n1253) );
INV_X1 U986 ( .A(G104), .ZN(n1258) );
NAND2_X1 U987 ( .A1(G214), .A2(n1259), .ZN(n1257) );
NAND2_X1 U988 ( .A1(KEYINPUT15), .A2(n1107), .ZN(n1248) );
INV_X1 U989 ( .A(G475), .ZN(n1107) );
XOR2_X1 U990 ( .A(n1260), .B(n1102), .Z(n1055) );
INV_X1 U991 ( .A(G478), .ZN(n1102) );
NAND2_X1 U992 ( .A1(n1100), .A2(n1139), .ZN(n1260) );
XNOR2_X1 U993 ( .A(n1261), .B(n1262), .ZN(n1100) );
XOR2_X1 U994 ( .A(G107), .B(n1263), .Z(n1262) );
XNOR2_X1 U995 ( .A(n1264), .B(G116), .ZN(n1263) );
INV_X1 U996 ( .A(G134), .ZN(n1264) );
XNOR2_X1 U997 ( .A(n1256), .B(n1265), .ZN(n1261) );
XOR2_X1 U998 ( .A(n1266), .B(n1267), .Z(n1265) );
NAND2_X1 U999 ( .A1(KEYINPUT49), .A2(G128), .ZN(n1267) );
NAND2_X1 U1000 ( .A1(G217), .A2(n1268), .ZN(n1266) );
XOR2_X1 U1001 ( .A(G122), .B(G143), .Z(n1256) );
INV_X1 U1002 ( .A(n1019), .ZN(n1153) );
NAND2_X1 U1003 ( .A1(n1269), .A2(n1045), .ZN(n1019) );
XOR2_X1 U1004 ( .A(n1270), .B(n1097), .Z(n1045) );
NAND2_X1 U1005 ( .A1(G217), .A2(n1232), .ZN(n1097) );
NAND2_X1 U1006 ( .A1(G234), .A2(n1139), .ZN(n1232) );
NAND2_X1 U1007 ( .A1(n1095), .A2(n1139), .ZN(n1270) );
XNOR2_X1 U1008 ( .A(n1271), .B(n1272), .ZN(n1095) );
XOR2_X1 U1009 ( .A(n1273), .B(n1274), .Z(n1272) );
XNOR2_X1 U1010 ( .A(n1275), .B(G110), .ZN(n1274) );
XOR2_X1 U1011 ( .A(KEYINPUT21), .B(G137), .Z(n1273) );
XOR2_X1 U1012 ( .A(n1276), .B(n1277), .Z(n1271) );
XOR2_X1 U1013 ( .A(n1278), .B(n1255), .Z(n1277) );
XNOR2_X1 U1014 ( .A(n1175), .B(G125), .ZN(n1255) );
INV_X1 U1015 ( .A(G146), .ZN(n1175) );
NOR2_X1 U1016 ( .A1(G140), .A2(KEYINPUT5), .ZN(n1278) );
XOR2_X1 U1017 ( .A(n1279), .B(n1280), .Z(n1276) );
NOR2_X1 U1018 ( .A1(G128), .A2(KEYINPUT23), .ZN(n1280) );
NAND2_X1 U1019 ( .A1(G221), .A2(n1268), .ZN(n1279) );
AND2_X1 U1020 ( .A1(G234), .A2(n1037), .ZN(n1268) );
INV_X1 U1021 ( .A(G953), .ZN(n1037) );
XOR2_X1 U1022 ( .A(KEYINPUT1), .B(n1201), .Z(n1269) );
XNOR2_X1 U1023 ( .A(n1186), .B(KEYINPUT4), .ZN(n1201) );
INV_X1 U1024 ( .A(n1203), .ZN(n1186) );
XOR2_X1 U1025 ( .A(n1053), .B(n1051), .Z(n1203) );
INV_X1 U1026 ( .A(G472), .ZN(n1051) );
NAND2_X1 U1027 ( .A1(n1281), .A2(n1139), .ZN(n1053) );
INV_X1 U1028 ( .A(G902), .ZN(n1139) );
XOR2_X1 U1029 ( .A(n1115), .B(n1282), .Z(n1281) );
XNOR2_X1 U1030 ( .A(n1283), .B(KEYINPUT7), .ZN(n1282) );
NAND2_X1 U1031 ( .A1(n1284), .A2(KEYINPUT11), .ZN(n1283) );
XNOR2_X1 U1032 ( .A(n1132), .B(n1285), .ZN(n1284) );
NOR2_X1 U1033 ( .A1(n1219), .A2(n1286), .ZN(n1285) );
XNOR2_X1 U1034 ( .A(KEYINPUT31), .B(KEYINPUT24), .ZN(n1286) );
INV_X1 U1035 ( .A(n1114), .ZN(n1219) );
XNOR2_X1 U1036 ( .A(n1237), .B(n1287), .ZN(n1114) );
NOR2_X1 U1037 ( .A1(G143), .A2(KEYINPUT59), .ZN(n1287) );
XNOR2_X1 U1038 ( .A(G146), .B(G128), .ZN(n1237) );
INV_X1 U1039 ( .A(n1118), .ZN(n1132) );
NAND2_X1 U1040 ( .A1(n1288), .A2(n1289), .ZN(n1118) );
OR2_X1 U1041 ( .A1(n1290), .A2(G131), .ZN(n1289) );
XOR2_X1 U1042 ( .A(n1291), .B(KEYINPUT35), .Z(n1288) );
NAND2_X1 U1043 ( .A1(G131), .A2(n1290), .ZN(n1291) );
XNOR2_X1 U1044 ( .A(n1070), .B(KEYINPUT12), .ZN(n1290) );
XNOR2_X1 U1045 ( .A(G134), .B(G137), .ZN(n1070) );
XNOR2_X1 U1046 ( .A(n1292), .B(n1293), .ZN(n1115) );
XOR2_X1 U1047 ( .A(n1294), .B(n1295), .Z(n1293) );
NAND2_X1 U1048 ( .A1(KEYINPUT8), .A2(n1275), .ZN(n1295) );
INV_X1 U1049 ( .A(G119), .ZN(n1275) );
NAND2_X1 U1050 ( .A1(G210), .A2(n1259), .ZN(n1294) );
NOR2_X1 U1051 ( .A1(G953), .A2(G237), .ZN(n1259) );
XNOR2_X1 U1052 ( .A(n1229), .B(n1296), .ZN(n1292) );
NOR2_X1 U1053 ( .A1(KEYINPUT56), .A2(n1207), .ZN(n1296) );
INV_X1 U1054 ( .A(G113), .ZN(n1207) );
XOR2_X1 U1055 ( .A(G101), .B(G116), .Z(n1229) );
endmodule


