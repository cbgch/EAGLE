//Key = 0100001111000000100010010111100101010111110100101010010101110010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378;

XNOR2_X1 U752 ( .A(G107), .B(n1054), .ZN(G9) );
NOR2_X1 U753 ( .A1(n1055), .A2(n1056), .ZN(G75) );
NOR4_X1 U754 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1056) );
NOR2_X1 U755 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NOR3_X1 U756 ( .A1(n1063), .A2(n1064), .A3(n1065), .ZN(n1061) );
NOR2_X1 U757 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
NOR4_X1 U758 ( .A1(n1068), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1064) );
NOR3_X1 U759 ( .A1(n1072), .A2(n1073), .A3(n1074), .ZN(n1068) );
NOR3_X1 U760 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1074) );
NOR2_X1 U761 ( .A1(n1078), .A2(n1079), .ZN(n1072) );
NOR2_X1 U762 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
XOR2_X1 U763 ( .A(n1082), .B(KEYINPUT37), .Z(n1063) );
NAND2_X1 U764 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U765 ( .A1(n1085), .A2(n1086), .ZN(n1059) );
XNOR2_X1 U766 ( .A(n1087), .B(KEYINPUT14), .ZN(n1085) );
NAND3_X1 U767 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1057) );
NAND3_X1 U768 ( .A1(n1091), .A2(n1087), .A3(n1092), .ZN(n1090) );
NOR3_X1 U769 ( .A1(n1069), .A2(n1070), .A3(n1067), .ZN(n1087) );
INV_X1 U770 ( .A(n1083), .ZN(n1067) );
NOR3_X1 U771 ( .A1(n1079), .A2(n1076), .A3(n1071), .ZN(n1083) );
NOR3_X1 U772 ( .A1(n1093), .A2(G953), .A3(G952), .ZN(n1055) );
INV_X1 U773 ( .A(n1088), .ZN(n1093) );
NAND4_X1 U774 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1088) );
NOR4_X1 U775 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XNOR2_X1 U776 ( .A(n1102), .B(KEYINPUT35), .ZN(n1101) );
XNOR2_X1 U777 ( .A(n1069), .B(KEYINPUT59), .ZN(n1100) );
NOR2_X1 U778 ( .A1(n1103), .A2(n1104), .ZN(n1099) );
NOR2_X1 U779 ( .A1(n1105), .A2(G469), .ZN(n1104) );
NOR2_X1 U780 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
AND2_X1 U781 ( .A1(n1108), .A2(KEYINPUT9), .ZN(n1106) );
NOR2_X1 U782 ( .A1(n1109), .A2(n1108), .ZN(n1103) );
NOR2_X1 U783 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
INV_X1 U784 ( .A(KEYINPUT9), .ZN(n1111) );
NOR2_X1 U785 ( .A1(n1112), .A2(n1107), .ZN(n1110) );
INV_X1 U786 ( .A(KEYINPUT50), .ZN(n1107) );
XNOR2_X1 U787 ( .A(n1113), .B(KEYINPUT4), .ZN(n1096) );
XOR2_X1 U788 ( .A(n1114), .B(n1115), .Z(G72) );
NOR2_X1 U789 ( .A1(n1116), .A2(n1089), .ZN(n1115) );
AND2_X1 U790 ( .A1(G227), .A2(G900), .ZN(n1116) );
NAND2_X1 U791 ( .A1(n1117), .A2(n1118), .ZN(n1114) );
NAND3_X1 U792 ( .A1(n1119), .A2(n1120), .A3(n1121), .ZN(n1118) );
NAND2_X1 U793 ( .A1(G953), .A2(n1122), .ZN(n1120) );
OR2_X1 U794 ( .A1(n1119), .A2(n1121), .ZN(n1117) );
NAND2_X1 U795 ( .A1(n1089), .A2(n1123), .ZN(n1121) );
NAND2_X1 U796 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U797 ( .A(KEYINPUT2), .B(n1126), .Z(n1125) );
INV_X1 U798 ( .A(n1127), .ZN(n1124) );
XOR2_X1 U799 ( .A(n1128), .B(n1129), .Z(n1119) );
XNOR2_X1 U800 ( .A(n1130), .B(n1131), .ZN(n1129) );
XNOR2_X1 U801 ( .A(n1132), .B(G131), .ZN(n1131) );
XOR2_X1 U802 ( .A(n1133), .B(n1134), .Z(n1128) );
NAND2_X1 U803 ( .A1(KEYINPUT58), .A2(n1135), .ZN(n1133) );
XOR2_X1 U804 ( .A(n1136), .B(n1137), .Z(G69) );
NOR2_X1 U805 ( .A1(n1138), .A2(G953), .ZN(n1137) );
NOR3_X1 U806 ( .A1(n1139), .A2(n1140), .A3(n1141), .ZN(n1138) );
XOR2_X1 U807 ( .A(n1142), .B(n1143), .Z(n1136) );
NOR2_X1 U808 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
NOR2_X1 U809 ( .A1(G224), .A2(n1089), .ZN(n1144) );
NAND2_X1 U810 ( .A1(n1146), .A2(n1147), .ZN(n1142) );
XOR2_X1 U811 ( .A(KEYINPUT40), .B(n1148), .Z(n1147) );
XOR2_X1 U812 ( .A(KEYINPUT6), .B(n1145), .Z(n1146) );
NOR2_X1 U813 ( .A1(n1149), .A2(n1150), .ZN(G66) );
XOR2_X1 U814 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U815 ( .A1(KEYINPUT13), .A2(n1153), .ZN(n1152) );
INV_X1 U816 ( .A(n1154), .ZN(n1153) );
NAND2_X1 U817 ( .A1(n1155), .A2(G217), .ZN(n1151) );
NOR2_X1 U818 ( .A1(n1149), .A2(n1156), .ZN(G63) );
XOR2_X1 U819 ( .A(n1157), .B(n1158), .Z(n1156) );
AND2_X1 U820 ( .A1(G478), .A2(n1155), .ZN(n1157) );
NOR2_X1 U821 ( .A1(n1149), .A2(n1159), .ZN(G60) );
XOR2_X1 U822 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND3_X1 U823 ( .A1(n1162), .A2(n1058), .A3(G475), .ZN(n1160) );
XNOR2_X1 U824 ( .A(KEYINPUT10), .B(n1163), .ZN(n1162) );
XNOR2_X1 U825 ( .A(n1164), .B(n1165), .ZN(G6) );
NOR2_X1 U826 ( .A1(KEYINPUT0), .A2(n1166), .ZN(n1165) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1167), .ZN(G57) );
XOR2_X1 U828 ( .A(n1168), .B(n1169), .Z(n1167) );
NAND2_X1 U829 ( .A1(n1170), .A2(KEYINPUT39), .ZN(n1169) );
XOR2_X1 U830 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U831 ( .A(n1173), .B(n1174), .Z(n1172) );
NOR2_X1 U832 ( .A1(KEYINPUT19), .A2(n1175), .ZN(n1174) );
AND2_X1 U833 ( .A1(G472), .A2(n1155), .ZN(n1173) );
INV_X1 U834 ( .A(n1176), .ZN(n1155) );
XNOR2_X1 U835 ( .A(n1177), .B(n1178), .ZN(n1171) );
NAND2_X1 U836 ( .A1(n1179), .A2(n1180), .ZN(n1168) );
NAND2_X1 U837 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
XOR2_X1 U838 ( .A(KEYINPUT43), .B(n1183), .Z(n1179) );
NOR2_X1 U839 ( .A1(n1182), .A2(n1181), .ZN(n1183) );
INV_X1 U840 ( .A(G101), .ZN(n1182) );
NOR2_X1 U841 ( .A1(n1149), .A2(n1184), .ZN(G54) );
XOR2_X1 U842 ( .A(n1185), .B(n1186), .Z(n1184) );
XNOR2_X1 U843 ( .A(n1187), .B(n1188), .ZN(n1186) );
NAND2_X1 U844 ( .A1(KEYINPUT25), .A2(n1189), .ZN(n1187) );
XOR2_X1 U845 ( .A(n1190), .B(n1191), .Z(n1185) );
XOR2_X1 U846 ( .A(G110), .B(n1192), .Z(n1191) );
NOR2_X1 U847 ( .A1(n1112), .A2(n1176), .ZN(n1192) );
NOR2_X1 U848 ( .A1(n1193), .A2(n1194), .ZN(n1190) );
XOR2_X1 U849 ( .A(n1195), .B(KEYINPUT8), .Z(n1194) );
NAND2_X1 U850 ( .A1(n1135), .A2(n1196), .ZN(n1195) );
NOR2_X1 U851 ( .A1(n1135), .A2(n1196), .ZN(n1193) );
NOR2_X1 U852 ( .A1(n1149), .A2(n1197), .ZN(G51) );
XOR2_X1 U853 ( .A(n1198), .B(n1199), .Z(n1197) );
XNOR2_X1 U854 ( .A(n1200), .B(n1201), .ZN(n1199) );
NOR3_X1 U855 ( .A1(n1202), .A2(KEYINPUT56), .A3(n1176), .ZN(n1201) );
NAND2_X1 U856 ( .A1(G902), .A2(n1058), .ZN(n1176) );
NAND3_X1 U857 ( .A1(n1203), .A2(n1126), .A3(n1204), .ZN(n1058) );
NOR3_X1 U858 ( .A1(n1139), .A2(n1205), .A3(n1127), .ZN(n1204) );
NAND4_X1 U859 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1127) );
XNOR2_X1 U860 ( .A(n1140), .B(KEYINPUT23), .ZN(n1205) );
NAND4_X1 U861 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1054), .ZN(n1139) );
NAND3_X1 U862 ( .A1(n1213), .A2(n1214), .A3(n1080), .ZN(n1054) );
NAND4_X1 U863 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1212) );
OR2_X1 U864 ( .A1(n1219), .A2(KEYINPUT45), .ZN(n1218) );
NAND2_X1 U865 ( .A1(KEYINPUT45), .A2(n1220), .ZN(n1217) );
NAND3_X1 U866 ( .A1(n1221), .A2(n1222), .A3(n1223), .ZN(n1220) );
NAND2_X1 U867 ( .A1(n1224), .A2(n1225), .ZN(n1211) );
NAND2_X1 U868 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND2_X1 U869 ( .A1(KEYINPUT16), .A2(n1081), .ZN(n1227) );
INV_X1 U870 ( .A(n1228), .ZN(n1224) );
NAND2_X1 U871 ( .A1(n1229), .A2(n1230), .ZN(n1210) );
NAND2_X1 U872 ( .A1(n1231), .A2(n1232), .ZN(n1230) );
OR4_X1 U873 ( .A1(n1233), .A2(n1234), .A3(n1223), .A4(KEYINPUT16), .ZN(n1232) );
NAND2_X1 U874 ( .A1(n1073), .A2(n1235), .ZN(n1231) );
NAND2_X1 U875 ( .A1(n1066), .A2(n1233), .ZN(n1235) );
INV_X1 U876 ( .A(n1236), .ZN(n1066) );
AND4_X1 U877 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1126) );
XNOR2_X1 U878 ( .A(n1141), .B(KEYINPUT44), .ZN(n1203) );
INV_X1 U879 ( .A(n1164), .ZN(n1141) );
NAND3_X1 U880 ( .A1(n1213), .A2(n1214), .A3(n1081), .ZN(n1164) );
XNOR2_X1 U881 ( .A(KEYINPUT53), .B(n1241), .ZN(n1202) );
NAND2_X1 U882 ( .A1(n1242), .A2(n1243), .ZN(n1198) );
NAND2_X1 U883 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
INV_X1 U884 ( .A(n1246), .ZN(n1245) );
XNOR2_X1 U885 ( .A(G125), .B(KEYINPUT3), .ZN(n1244) );
NAND2_X1 U886 ( .A1(n1247), .A2(n1246), .ZN(n1242) );
XOR2_X1 U887 ( .A(n1178), .B(KEYINPUT26), .Z(n1246) );
XNOR2_X1 U888 ( .A(KEYINPUT21), .B(n1130), .ZN(n1247) );
INV_X1 U889 ( .A(G125), .ZN(n1130) );
NOR2_X1 U890 ( .A1(n1089), .A2(G952), .ZN(n1149) );
XNOR2_X1 U891 ( .A(n1237), .B(n1248), .ZN(G48) );
NOR2_X1 U892 ( .A1(KEYINPUT36), .A2(n1249), .ZN(n1248) );
NAND3_X1 U893 ( .A1(n1250), .A2(n1222), .A3(n1081), .ZN(n1237) );
XNOR2_X1 U894 ( .A(G143), .B(n1238), .ZN(G45) );
NAND4_X1 U895 ( .A1(n1251), .A2(n1222), .A3(n1102), .A4(n1113), .ZN(n1238) );
XNOR2_X1 U896 ( .A(G140), .B(n1239), .ZN(G42) );
NAND3_X1 U897 ( .A1(n1094), .A2(n1214), .A3(n1252), .ZN(n1239) );
XNOR2_X1 U898 ( .A(G137), .B(n1240), .ZN(G39) );
NAND3_X1 U899 ( .A1(n1250), .A2(n1094), .A3(n1215), .ZN(n1240) );
XNOR2_X1 U900 ( .A(G134), .B(n1209), .ZN(G36) );
NAND3_X1 U901 ( .A1(n1094), .A2(n1080), .A3(n1251), .ZN(n1209) );
XNOR2_X1 U902 ( .A(G131), .B(n1206), .ZN(G33) );
NAND3_X1 U903 ( .A1(n1081), .A2(n1094), .A3(n1251), .ZN(n1206) );
AND3_X1 U904 ( .A1(n1214), .A2(n1253), .A3(n1084), .ZN(n1251) );
INV_X1 U905 ( .A(n1062), .ZN(n1094) );
NAND2_X1 U906 ( .A1(n1091), .A2(n1254), .ZN(n1062) );
INV_X1 U907 ( .A(n1092), .ZN(n1254) );
XNOR2_X1 U908 ( .A(G128), .B(n1207), .ZN(G30) );
NAND3_X1 U909 ( .A1(n1080), .A2(n1222), .A3(n1250), .ZN(n1207) );
AND3_X1 U910 ( .A1(n1214), .A2(n1253), .A3(n1216), .ZN(n1250) );
XNOR2_X1 U911 ( .A(G101), .B(n1255), .ZN(G3) );
NAND4_X1 U912 ( .A1(n1256), .A2(n1073), .A3(n1084), .A4(n1257), .ZN(n1255) );
XNOR2_X1 U913 ( .A(n1222), .B(KEYINPUT7), .ZN(n1256) );
XNOR2_X1 U914 ( .A(G125), .B(n1258), .ZN(G27) );
NOR2_X1 U915 ( .A1(n1259), .A2(KEYINPUT61), .ZN(n1258) );
INV_X1 U916 ( .A(n1208), .ZN(n1259) );
NAND3_X1 U917 ( .A1(n1252), .A2(n1222), .A3(n1223), .ZN(n1208) );
AND3_X1 U918 ( .A1(n1081), .A2(n1253), .A3(n1236), .ZN(n1252) );
NAND2_X1 U919 ( .A1(n1071), .A2(n1260), .ZN(n1253) );
NAND4_X1 U920 ( .A1(G902), .A2(G953), .A3(n1261), .A4(n1122), .ZN(n1260) );
INV_X1 U921 ( .A(G900), .ZN(n1122) );
INV_X1 U922 ( .A(n1234), .ZN(n1081) );
XNOR2_X1 U923 ( .A(G122), .B(n1262), .ZN(G24) );
NAND3_X1 U924 ( .A1(n1263), .A2(n1264), .A3(KEYINPUT31), .ZN(n1262) );
OR2_X1 U925 ( .A1(n1140), .A2(KEYINPUT30), .ZN(n1264) );
AND4_X1 U926 ( .A1(n1223), .A2(n1213), .A3(n1102), .A4(n1113), .ZN(n1140) );
NAND2_X1 U927 ( .A1(KEYINPUT30), .A2(n1265), .ZN(n1263) );
NAND3_X1 U928 ( .A1(n1213), .A2(n1266), .A3(n1223), .ZN(n1265) );
NAND2_X1 U929 ( .A1(n1102), .A2(n1113), .ZN(n1266) );
AND3_X1 U930 ( .A1(n1267), .A2(n1095), .A3(n1229), .ZN(n1213) );
XNOR2_X1 U931 ( .A(n1268), .B(n1269), .ZN(G21) );
NAND2_X1 U932 ( .A1(KEYINPUT62), .A2(n1270), .ZN(n1268) );
NAND3_X1 U933 ( .A1(n1216), .A2(n1271), .A3(n1219), .ZN(n1270) );
XNOR2_X1 U934 ( .A(KEYINPUT60), .B(n1076), .ZN(n1271) );
INV_X1 U935 ( .A(n1215), .ZN(n1076) );
NOR2_X1 U936 ( .A1(n1267), .A2(n1095), .ZN(n1216) );
XOR2_X1 U937 ( .A(G116), .B(n1272), .Z(G18) );
NOR3_X1 U938 ( .A1(n1228), .A2(KEYINPUT51), .A3(n1226), .ZN(n1272) );
INV_X1 U939 ( .A(n1080), .ZN(n1226) );
NOR2_X1 U940 ( .A1(n1113), .A2(n1273), .ZN(n1080) );
XNOR2_X1 U941 ( .A(G113), .B(n1274), .ZN(G15) );
NOR2_X1 U942 ( .A1(n1275), .A2(n1276), .ZN(n1274) );
NOR3_X1 U943 ( .A1(n1277), .A2(n1278), .A3(n1086), .ZN(n1276) );
NOR4_X1 U944 ( .A1(n1221), .A2(n1234), .A3(n1233), .A4(n1079), .ZN(n1278) );
INV_X1 U945 ( .A(n1223), .ZN(n1079) );
INV_X1 U946 ( .A(n1084), .ZN(n1233) );
INV_X1 U947 ( .A(KEYINPUT42), .ZN(n1277) );
NOR3_X1 U948 ( .A1(KEYINPUT42), .A2(n1234), .A3(n1228), .ZN(n1275) );
NAND2_X1 U949 ( .A1(n1219), .A2(n1084), .ZN(n1228) );
NOR2_X1 U950 ( .A1(n1070), .A2(n1267), .ZN(n1084) );
INV_X1 U951 ( .A(n1069), .ZN(n1267) );
AND2_X1 U952 ( .A1(n1223), .A2(n1229), .ZN(n1219) );
NOR2_X1 U953 ( .A1(n1086), .A2(n1221), .ZN(n1229) );
INV_X1 U954 ( .A(n1257), .ZN(n1221) );
INV_X1 U955 ( .A(n1222), .ZN(n1086) );
NOR2_X1 U956 ( .A1(n1077), .A2(n1098), .ZN(n1223) );
INV_X1 U957 ( .A(n1075), .ZN(n1098) );
NAND2_X1 U958 ( .A1(n1273), .A2(n1113), .ZN(n1234) );
INV_X1 U959 ( .A(n1102), .ZN(n1273) );
XOR2_X1 U960 ( .A(n1279), .B(n1280), .Z(G12) );
NAND2_X1 U961 ( .A1(KEYINPUT46), .A2(G110), .ZN(n1280) );
NAND4_X1 U962 ( .A1(n1281), .A2(n1073), .A3(n1236), .A4(n1257), .ZN(n1279) );
NAND2_X1 U963 ( .A1(n1071), .A2(n1282), .ZN(n1257) );
NAND3_X1 U964 ( .A1(n1145), .A2(n1261), .A3(G902), .ZN(n1282) );
NOR2_X1 U965 ( .A1(G898), .A2(n1089), .ZN(n1145) );
NAND3_X1 U966 ( .A1(n1261), .A2(n1089), .A3(G952), .ZN(n1071) );
NAND2_X1 U967 ( .A1(G234), .A2(G237), .ZN(n1261) );
NOR2_X1 U968 ( .A1(n1069), .A2(n1095), .ZN(n1236) );
INV_X1 U969 ( .A(n1070), .ZN(n1095) );
NAND3_X1 U970 ( .A1(n1283), .A2(n1284), .A3(n1285), .ZN(n1070) );
NAND2_X1 U971 ( .A1(G902), .A2(G217), .ZN(n1285) );
NAND3_X1 U972 ( .A1(n1154), .A2(n1163), .A3(n1286), .ZN(n1284) );
OR2_X1 U973 ( .A1(n1286), .A2(n1154), .ZN(n1283) );
XNOR2_X1 U974 ( .A(n1287), .B(n1288), .ZN(n1154) );
XOR2_X1 U975 ( .A(n1134), .B(n1289), .Z(n1288) );
XNOR2_X1 U976 ( .A(n1290), .B(G140), .ZN(n1134) );
INV_X1 U977 ( .A(G137), .ZN(n1290) );
XOR2_X1 U978 ( .A(n1291), .B(n1292), .Z(n1287) );
NOR4_X1 U979 ( .A1(KEYINPUT17), .A2(G953), .A3(n1293), .A4(n1294), .ZN(n1292) );
INV_X1 U980 ( .A(G221), .ZN(n1294) );
NAND2_X1 U981 ( .A1(n1295), .A2(n1296), .ZN(n1291) );
NAND2_X1 U982 ( .A1(n1297), .A2(n1298), .ZN(n1296) );
XOR2_X1 U983 ( .A(n1299), .B(KEYINPUT12), .Z(n1295) );
OR2_X1 U984 ( .A1(n1298), .A2(n1297), .ZN(n1299) );
AND2_X1 U985 ( .A1(n1300), .A2(n1301), .ZN(n1297) );
NAND2_X1 U986 ( .A1(G119), .A2(n1302), .ZN(n1301) );
XOR2_X1 U987 ( .A(n1303), .B(KEYINPUT52), .Z(n1300) );
NAND2_X1 U988 ( .A1(G128), .A2(n1269), .ZN(n1303) );
XOR2_X1 U989 ( .A(G110), .B(KEYINPUT48), .Z(n1298) );
NAND2_X1 U990 ( .A1(G217), .A2(n1293), .ZN(n1286) );
INV_X1 U991 ( .A(G234), .ZN(n1293) );
XNOR2_X1 U992 ( .A(n1304), .B(G472), .ZN(n1069) );
NAND2_X1 U993 ( .A1(n1305), .A2(n1163), .ZN(n1304) );
XOR2_X1 U994 ( .A(n1306), .B(n1307), .Z(n1305) );
XNOR2_X1 U995 ( .A(n1308), .B(n1175), .ZN(n1307) );
INV_X1 U996 ( .A(n1309), .ZN(n1175) );
NOR2_X1 U997 ( .A1(KEYINPUT47), .A2(n1181), .ZN(n1308) );
OR2_X1 U998 ( .A1(n1241), .A2(n1310), .ZN(n1181) );
XOR2_X1 U999 ( .A(n1311), .B(n1312), .Z(n1306) );
NOR2_X1 U1000 ( .A1(KEYINPUT29), .A2(n1313), .ZN(n1312) );
XNOR2_X1 U1001 ( .A(n1314), .B(n1178), .ZN(n1313) );
NAND2_X1 U1002 ( .A1(KEYINPUT27), .A2(n1315), .ZN(n1314) );
XNOR2_X1 U1003 ( .A(G101), .B(KEYINPUT28), .ZN(n1311) );
AND2_X1 U1004 ( .A1(n1215), .A2(n1214), .ZN(n1073) );
AND2_X1 U1005 ( .A1(n1077), .A2(n1075), .ZN(n1214) );
NAND2_X1 U1006 ( .A1(G221), .A2(n1316), .ZN(n1075) );
NAND2_X1 U1007 ( .A1(G234), .A2(n1163), .ZN(n1316) );
XOR2_X1 U1008 ( .A(n1108), .B(n1112), .Z(n1077) );
INV_X1 U1009 ( .A(G469), .ZN(n1112) );
NAND2_X1 U1010 ( .A1(n1317), .A2(n1163), .ZN(n1108) );
XOR2_X1 U1011 ( .A(n1318), .B(n1319), .Z(n1317) );
XNOR2_X1 U1012 ( .A(n1189), .B(n1320), .ZN(n1319) );
NOR2_X1 U1013 ( .A1(KEYINPUT15), .A2(n1321), .ZN(n1320) );
XOR2_X1 U1014 ( .A(n1135), .B(n1196), .Z(n1321) );
XOR2_X1 U1015 ( .A(G107), .B(n1322), .Z(n1196) );
AND2_X1 U1016 ( .A1(n1323), .A2(n1324), .ZN(n1135) );
NAND2_X1 U1017 ( .A1(n1325), .A2(G128), .ZN(n1324) );
XOR2_X1 U1018 ( .A(n1326), .B(KEYINPUT11), .Z(n1323) );
NAND2_X1 U1019 ( .A1(n1327), .A2(n1302), .ZN(n1326) );
INV_X1 U1020 ( .A(G128), .ZN(n1302) );
XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n1325), .ZN(n1327) );
XNOR2_X1 U1022 ( .A(n1328), .B(KEYINPUT57), .ZN(n1325) );
XNOR2_X1 U1023 ( .A(n1329), .B(n1330), .ZN(n1318) );
INV_X1 U1024 ( .A(n1188), .ZN(n1330) );
XOR2_X1 U1025 ( .A(n1331), .B(n1315), .Z(n1188) );
INV_X1 U1026 ( .A(n1177), .ZN(n1315) );
XNOR2_X1 U1027 ( .A(n1332), .B(n1333), .ZN(n1177) );
NOR2_X1 U1028 ( .A1(KEYINPUT5), .A2(n1132), .ZN(n1333) );
XNOR2_X1 U1029 ( .A(G137), .B(G131), .ZN(n1332) );
NAND2_X1 U1030 ( .A1(G227), .A2(n1089), .ZN(n1331) );
NAND2_X1 U1031 ( .A1(KEYINPUT41), .A2(G110), .ZN(n1329) );
NOR2_X1 U1032 ( .A1(n1102), .A2(n1113), .ZN(n1215) );
XNOR2_X1 U1033 ( .A(n1334), .B(G475), .ZN(n1113) );
NAND2_X1 U1034 ( .A1(n1161), .A2(n1163), .ZN(n1334) );
XNOR2_X1 U1035 ( .A(G113), .B(n1335), .ZN(n1161) );
XOR2_X1 U1036 ( .A(n1336), .B(n1337), .Z(n1335) );
XOR2_X1 U1037 ( .A(n1338), .B(n1339), .Z(n1337) );
XOR2_X1 U1038 ( .A(n1340), .B(n1341), .Z(n1339) );
NOR2_X1 U1039 ( .A1(G143), .A2(KEYINPUT34), .ZN(n1341) );
NOR2_X1 U1040 ( .A1(n1310), .A2(n1342), .ZN(n1340) );
NAND2_X1 U1041 ( .A1(n1343), .A2(n1089), .ZN(n1310) );
XNOR2_X1 U1042 ( .A(G237), .B(KEYINPUT54), .ZN(n1343) );
XOR2_X1 U1043 ( .A(n1344), .B(n1289), .Z(n1338) );
XNOR2_X1 U1044 ( .A(n1249), .B(G125), .ZN(n1289) );
INV_X1 U1045 ( .A(G146), .ZN(n1249) );
NAND2_X1 U1046 ( .A1(KEYINPUT20), .A2(n1189), .ZN(n1344) );
INV_X1 U1047 ( .A(G140), .ZN(n1189) );
XOR2_X1 U1048 ( .A(n1345), .B(n1346), .Z(n1336) );
XOR2_X1 U1049 ( .A(KEYINPUT55), .B(G131), .Z(n1346) );
XNOR2_X1 U1050 ( .A(G104), .B(G122), .ZN(n1345) );
XNOR2_X1 U1051 ( .A(n1347), .B(G478), .ZN(n1102) );
OR2_X1 U1052 ( .A1(n1158), .A2(G902), .ZN(n1347) );
XNOR2_X1 U1053 ( .A(n1348), .B(n1349), .ZN(n1158) );
XOR2_X1 U1054 ( .A(G107), .B(n1350), .Z(n1349) );
XNOR2_X1 U1055 ( .A(n1132), .B(G128), .ZN(n1350) );
INV_X1 U1056 ( .A(G134), .ZN(n1132) );
XOR2_X1 U1057 ( .A(n1351), .B(n1352), .Z(n1348) );
XOR2_X1 U1058 ( .A(n1353), .B(n1354), .Z(n1352) );
NAND2_X1 U1059 ( .A1(KEYINPUT1), .A2(n1355), .ZN(n1354) );
INV_X1 U1060 ( .A(G143), .ZN(n1355) );
NAND3_X1 U1061 ( .A1(n1356), .A2(n1357), .A3(n1358), .ZN(n1353) );
NAND2_X1 U1062 ( .A1(KEYINPUT18), .A2(G116), .ZN(n1358) );
NAND3_X1 U1063 ( .A1(n1359), .A2(n1360), .A3(n1361), .ZN(n1357) );
INV_X1 U1064 ( .A(KEYINPUT18), .ZN(n1360) );
OR2_X1 U1065 ( .A1(n1361), .A2(n1359), .ZN(n1356) );
NOR2_X1 U1066 ( .A1(G116), .A2(KEYINPUT22), .ZN(n1359) );
NAND3_X1 U1067 ( .A1(G217), .A2(n1089), .A3(G234), .ZN(n1351) );
XNOR2_X1 U1068 ( .A(n1222), .B(KEYINPUT38), .ZN(n1281) );
NOR2_X1 U1069 ( .A1(n1091), .A2(n1092), .ZN(n1222) );
NOR2_X1 U1070 ( .A1(n1342), .A2(n1362), .ZN(n1092) );
INV_X1 U1071 ( .A(G214), .ZN(n1342) );
XOR2_X1 U1072 ( .A(n1363), .B(n1364), .Z(n1091) );
NOR2_X1 U1073 ( .A1(n1362), .A2(n1241), .ZN(n1364) );
INV_X1 U1074 ( .A(G210), .ZN(n1241) );
NOR2_X1 U1075 ( .A1(G902), .A2(G237), .ZN(n1362) );
NAND2_X1 U1076 ( .A1(n1365), .A2(n1163), .ZN(n1363) );
INV_X1 U1077 ( .A(G902), .ZN(n1163) );
XNOR2_X1 U1078 ( .A(n1366), .B(n1367), .ZN(n1365) );
INV_X1 U1079 ( .A(n1200), .ZN(n1367) );
XOR2_X1 U1080 ( .A(n1148), .B(n1368), .Z(n1200) );
AND2_X1 U1081 ( .A1(n1089), .A2(G224), .ZN(n1368) );
INV_X1 U1082 ( .A(G953), .ZN(n1089) );
XNOR2_X1 U1083 ( .A(n1369), .B(n1370), .ZN(n1148) );
XOR2_X1 U1084 ( .A(n1371), .B(n1372), .Z(n1370) );
NOR2_X1 U1085 ( .A1(n1373), .A2(n1374), .ZN(n1372) );
XOR2_X1 U1086 ( .A(n1375), .B(KEYINPUT33), .Z(n1374) );
NAND2_X1 U1087 ( .A1(G110), .A2(n1361), .ZN(n1375) );
NOR2_X1 U1088 ( .A1(G110), .A2(n1361), .ZN(n1373) );
INV_X1 U1089 ( .A(G122), .ZN(n1361) );
NOR2_X1 U1090 ( .A1(G107), .A2(KEYINPUT32), .ZN(n1371) );
XNOR2_X1 U1091 ( .A(n1309), .B(n1322), .ZN(n1369) );
XNOR2_X1 U1092 ( .A(n1166), .B(G101), .ZN(n1322) );
INV_X1 U1093 ( .A(G104), .ZN(n1166) );
XOR2_X1 U1094 ( .A(G113), .B(n1376), .Z(n1309) );
XNOR2_X1 U1095 ( .A(n1269), .B(G116), .ZN(n1376) );
INV_X1 U1096 ( .A(G119), .ZN(n1269) );
NOR2_X1 U1097 ( .A1(KEYINPUT63), .A2(n1377), .ZN(n1366) );
XNOR2_X1 U1098 ( .A(G125), .B(n1178), .ZN(n1377) );
XNOR2_X1 U1099 ( .A(n1378), .B(n1328), .ZN(n1178) );
XOR2_X1 U1100 ( .A(G146), .B(G143), .Z(n1328) );
XNOR2_X1 U1101 ( .A(G128), .B(KEYINPUT24), .ZN(n1378) );
endmodule


