//Key = 0100011110111010101010010100010100111001101011010000101101010010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
n1311, n1312, n1313;

XOR2_X1 U714 ( .A(G107), .B(n990), .Z(G9) );
NOR2_X1 U715 ( .A1(n991), .A2(n992), .ZN(G75) );
NOR4_X1 U716 ( .A1(G953), .A2(n993), .A3(n994), .A4(n995), .ZN(n992) );
NOR2_X1 U717 ( .A1(n996), .A2(n997), .ZN(n994) );
NOR2_X1 U718 ( .A1(n998), .A2(n999), .ZN(n996) );
NOR2_X1 U719 ( .A1(n1000), .A2(n1001), .ZN(n999) );
NOR2_X1 U720 ( .A1(n1002), .A2(n1003), .ZN(n1000) );
NOR2_X1 U721 ( .A1(n1004), .A2(n1005), .ZN(n1002) );
NOR3_X1 U722 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n998) );
NOR2_X1 U723 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR3_X1 U724 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1009) );
NOR3_X1 U725 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1012) );
NOR2_X1 U726 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U727 ( .A1(n1018), .A2(n1019), .ZN(n1014) );
NOR2_X1 U728 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
AND2_X1 U729 ( .A1(n1001), .A2(n1013), .ZN(n1011) );
NOR3_X1 U730 ( .A1(n1001), .A2(n1016), .A3(n1013), .ZN(n1008) );
NOR3_X1 U731 ( .A1(n1022), .A2(n1010), .A3(n1023), .ZN(n1016) );
NAND2_X1 U732 ( .A1(n1024), .A2(n1025), .ZN(n1001) );
NOR3_X1 U733 ( .A1(n993), .A2(G953), .A3(G952), .ZN(n991) );
AND4_X1 U734 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n993) );
NOR4_X1 U735 ( .A1(n1030), .A2(n1031), .A3(n1010), .A4(n1013), .ZN(n1029) );
NOR2_X1 U736 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NOR2_X1 U737 ( .A1(G469), .A2(KEYINPUT0), .ZN(n1033) );
NAND2_X1 U738 ( .A1(n1034), .A2(n1035), .ZN(n1030) );
NAND2_X1 U739 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
NAND4_X1 U740 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1036) );
NAND3_X1 U741 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1041) );
INV_X1 U742 ( .A(KEYINPUT0), .ZN(n1043) );
NAND2_X1 U743 ( .A1(n1045), .A2(n1046), .ZN(n1040) );
NAND2_X1 U744 ( .A1(n1047), .A2(n1048), .ZN(n1039) );
NAND2_X1 U745 ( .A1(n1049), .A2(n1050), .ZN(n1038) );
OR2_X1 U746 ( .A1(n1048), .A2(n1051), .ZN(n1034) );
NOR3_X1 U747 ( .A1(n1052), .A2(n1053), .A3(n1054), .ZN(n1028) );
NOR3_X1 U748 ( .A1(n1055), .A2(n1056), .A3(n1050), .ZN(n1054) );
AND2_X1 U749 ( .A1(n1055), .A2(n1050), .ZN(n1053) );
INV_X1 U750 ( .A(KEYINPUT45), .ZN(n1055) );
OR2_X1 U751 ( .A1(n1046), .A2(n1057), .ZN(n1027) );
XOR2_X1 U752 ( .A(n1058), .B(n1059), .Z(G72) );
NAND2_X1 U753 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
OR3_X1 U754 ( .A1(n1062), .A2(G227), .A3(n1063), .ZN(n1061) );
NAND2_X1 U755 ( .A1(n1064), .A2(n1063), .ZN(n1060) );
NAND2_X1 U756 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
XNOR2_X1 U757 ( .A(n1067), .B(n1068), .ZN(n1065) );
NAND2_X1 U758 ( .A1(KEYINPUT34), .A2(n1069), .ZN(n1067) );
XOR2_X1 U759 ( .A(n1070), .B(n1071), .Z(n1069) );
XNOR2_X1 U760 ( .A(n1072), .B(n1073), .ZN(n1071) );
XNOR2_X1 U761 ( .A(G131), .B(n1074), .ZN(n1070) );
NOR2_X1 U762 ( .A1(KEYINPUT3), .A2(n1075), .ZN(n1074) );
XNOR2_X1 U763 ( .A(n1076), .B(n1077), .ZN(n1075) );
NOR2_X1 U764 ( .A1(G137), .A2(KEYINPUT41), .ZN(n1077) );
NAND2_X1 U765 ( .A1(G953), .A2(n1078), .ZN(n1064) );
NAND2_X1 U766 ( .A1(G900), .A2(G227), .ZN(n1078) );
NAND2_X1 U767 ( .A1(n1062), .A2(n1079), .ZN(n1058) );
NAND2_X1 U768 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XNOR2_X1 U769 ( .A(KEYINPUT42), .B(n1082), .ZN(n1081) );
XOR2_X1 U770 ( .A(n1083), .B(n1084), .Z(G69) );
NOR2_X1 U771 ( .A1(n1085), .A2(n1062), .ZN(n1084) );
NOR2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U773 ( .A1(n1088), .A2(n1089), .ZN(n1083) );
NAND2_X1 U774 ( .A1(n1090), .A2(n1062), .ZN(n1089) );
XOR2_X1 U775 ( .A(n1091), .B(n1092), .Z(n1090) );
OR3_X1 U776 ( .A1(n1091), .A2(n1087), .A3(n1062), .ZN(n1088) );
NAND2_X1 U777 ( .A1(n1093), .A2(KEYINPUT40), .ZN(n1091) );
XOR2_X1 U778 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U779 ( .A1(n1096), .A2(n1097), .ZN(G66) );
XNOR2_X1 U780 ( .A(n1049), .B(n1098), .ZN(n1097) );
NOR2_X1 U781 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
NOR2_X1 U782 ( .A1(n1096), .A2(n1101), .ZN(G63) );
XOR2_X1 U783 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U784 ( .A1(KEYINPUT60), .A2(n1104), .ZN(n1103) );
XOR2_X1 U785 ( .A(KEYINPUT18), .B(n1105), .Z(n1104) );
NAND2_X1 U786 ( .A1(n1106), .A2(G478), .ZN(n1102) );
NOR2_X1 U787 ( .A1(n1096), .A2(n1107), .ZN(G60) );
XNOR2_X1 U788 ( .A(n1045), .B(n1108), .ZN(n1107) );
NOR2_X1 U789 ( .A1(n1046), .A2(n1100), .ZN(n1108) );
INV_X1 U790 ( .A(G475), .ZN(n1046) );
XNOR2_X1 U791 ( .A(n1109), .B(n1110), .ZN(G6) );
XOR2_X1 U792 ( .A(KEYINPUT53), .B(G104), .Z(n1110) );
NOR2_X1 U793 ( .A1(n1096), .A2(n1111), .ZN(G57) );
XOR2_X1 U794 ( .A(n1112), .B(n1113), .Z(n1111) );
XOR2_X1 U795 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U796 ( .A(n1116), .B(n1117), .Z(n1115) );
AND2_X1 U797 ( .A1(G472), .A2(n1106), .ZN(n1116) );
INV_X1 U798 ( .A(n1100), .ZN(n1106) );
XOR2_X1 U799 ( .A(n1118), .B(n1119), .Z(n1112) );
XNOR2_X1 U800 ( .A(KEYINPUT25), .B(KEYINPUT2), .ZN(n1119) );
NOR2_X1 U801 ( .A1(n1096), .A2(n1120), .ZN(G54) );
XOR2_X1 U802 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U803 ( .A(n1123), .B(n1124), .Z(n1122) );
NAND2_X1 U804 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
INV_X1 U805 ( .A(n1127), .ZN(n1126) );
NAND2_X1 U806 ( .A1(n1128), .A2(n1129), .ZN(n1123) );
NAND2_X1 U807 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U808 ( .A(n1132), .B(G101), .Z(n1131) );
XNOR2_X1 U809 ( .A(KEYINPUT22), .B(n1133), .ZN(n1130) );
XOR2_X1 U810 ( .A(n1134), .B(KEYINPUT51), .Z(n1128) );
NAND2_X1 U811 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
XNOR2_X1 U812 ( .A(G101), .B(n1132), .ZN(n1136) );
XOR2_X1 U813 ( .A(KEYINPUT22), .B(n1133), .Z(n1135) );
NOR2_X1 U814 ( .A1(n1042), .A2(n1100), .ZN(n1121) );
NOR2_X1 U815 ( .A1(n1096), .A2(n1137), .ZN(G51) );
NOR2_X1 U816 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
XOR2_X1 U817 ( .A(KEYINPUT24), .B(n1140), .Z(n1139) );
AND2_X1 U818 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
NOR2_X1 U819 ( .A1(n1142), .A2(n1141), .ZN(n1138) );
XOR2_X1 U820 ( .A(n1047), .B(KEYINPUT1), .Z(n1141) );
NOR2_X1 U821 ( .A1(n1100), .A2(n1048), .ZN(n1142) );
NAND2_X1 U822 ( .A1(G902), .A2(n995), .ZN(n1100) );
NAND3_X1 U823 ( .A1(n1080), .A2(n1082), .A3(n1092), .ZN(n995) );
AND4_X1 U824 ( .A1(n1143), .A2(n1109), .A3(n1144), .A4(n1145), .ZN(n1092) );
NOR4_X1 U825 ( .A1(n1146), .A2(n1147), .A3(n990), .A4(n1148), .ZN(n1145) );
AND2_X1 U826 ( .A1(n1020), .A2(n1149), .ZN(n990) );
INV_X1 U827 ( .A(n1150), .ZN(n1147) );
NOR2_X1 U828 ( .A1(n1151), .A2(n1152), .ZN(n1144) );
NOR2_X1 U829 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
XNOR2_X1 U830 ( .A(KEYINPUT6), .B(n1155), .ZN(n1154) );
INV_X1 U831 ( .A(n1156), .ZN(n1151) );
NAND2_X1 U832 ( .A1(n1021), .A2(n1149), .ZN(n1109) );
AND3_X1 U833 ( .A1(n1025), .A2(n1157), .A3(n1158), .ZN(n1149) );
NAND4_X1 U834 ( .A1(n1159), .A2(n1022), .A3(n1024), .A4(n1158), .ZN(n1143) );
XOR2_X1 U835 ( .A(n1157), .B(KEYINPUT13), .Z(n1159) );
AND4_X1 U836 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1080) );
AND4_X1 U837 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163) );
NAND2_X1 U838 ( .A1(n1168), .A2(n1169), .ZN(n1162) );
INV_X1 U839 ( .A(KEYINPUT30), .ZN(n1169) );
NAND2_X1 U840 ( .A1(n1022), .A2(n1170), .ZN(n1160) );
NAND2_X1 U841 ( .A1(n1171), .A2(n1172), .ZN(n1170) );
NAND3_X1 U842 ( .A1(n1173), .A2(n1174), .A3(KEYINPUT30), .ZN(n1172) );
NAND2_X1 U843 ( .A1(n1175), .A2(n1020), .ZN(n1171) );
NOR2_X1 U844 ( .A1(n1062), .A2(G952), .ZN(n1096) );
NAND2_X1 U845 ( .A1(n1176), .A2(n1177), .ZN(G48) );
NAND2_X1 U846 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U847 ( .A(KEYINPUT29), .B(n1180), .Z(n1176) );
NOR2_X1 U848 ( .A1(n1178), .A2(n1179), .ZN(n1180) );
INV_X1 U849 ( .A(G146), .ZN(n1179) );
INV_X1 U850 ( .A(n1161), .ZN(n1178) );
NAND3_X1 U851 ( .A1(n1181), .A2(n1021), .A3(n1173), .ZN(n1161) );
NAND2_X1 U852 ( .A1(n1182), .A2(n1183), .ZN(G45) );
NAND2_X1 U853 ( .A1(n1168), .A2(n1184), .ZN(n1183) );
XOR2_X1 U854 ( .A(KEYINPUT20), .B(n1185), .Z(n1182) );
NOR2_X1 U855 ( .A1(n1168), .A2(n1184), .ZN(n1185) );
AND3_X1 U856 ( .A1(n1022), .A2(n1186), .A3(n1173), .ZN(n1168) );
XOR2_X1 U857 ( .A(n1167), .B(n1187), .Z(G42) );
XNOR2_X1 U858 ( .A(G140), .B(KEYINPUT38), .ZN(n1187) );
NAND3_X1 U859 ( .A1(n1021), .A2(n1023), .A3(n1175), .ZN(n1167) );
XNOR2_X1 U860 ( .A(G137), .B(n1166), .ZN(G39) );
NAND3_X1 U861 ( .A1(n1181), .A2(n1024), .A3(n1175), .ZN(n1166) );
XOR2_X1 U862 ( .A(n1188), .B(n1189), .Z(G36) );
XNOR2_X1 U863 ( .A(KEYINPUT57), .B(n1076), .ZN(n1189) );
NAND3_X1 U864 ( .A1(n1020), .A2(n1190), .A3(n1175), .ZN(n1188) );
XNOR2_X1 U865 ( .A(KEYINPUT50), .B(n1191), .ZN(n1190) );
XNOR2_X1 U866 ( .A(n1192), .B(n1193), .ZN(G33) );
NOR2_X1 U867 ( .A1(KEYINPUT9), .A2(n1082), .ZN(n1193) );
NAND3_X1 U868 ( .A1(n1021), .A2(n1022), .A3(n1175), .ZN(n1082) );
NOR3_X1 U869 ( .A1(n1004), .A2(n1194), .A3(n1005), .ZN(n1175) );
INV_X1 U870 ( .A(n1195), .ZN(n1194) );
XNOR2_X1 U871 ( .A(G128), .B(n1165), .ZN(G30) );
NAND3_X1 U872 ( .A1(n1181), .A2(n1020), .A3(n1173), .ZN(n1165) );
AND2_X1 U873 ( .A1(n1158), .A2(n1195), .ZN(n1173) );
INV_X1 U874 ( .A(n1155), .ZN(n1181) );
XOR2_X1 U875 ( .A(G101), .B(n1196), .Z(G3) );
NOR3_X1 U876 ( .A1(n1191), .A2(KEYINPUT26), .A3(n1197), .ZN(n1196) );
NAND2_X1 U877 ( .A1(n1198), .A2(n1199), .ZN(G27) );
NAND2_X1 U878 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
XOR2_X1 U879 ( .A(KEYINPUT31), .B(n1202), .Z(n1198) );
NOR2_X1 U880 ( .A1(n1200), .A2(n1201), .ZN(n1202) );
XNOR2_X1 U881 ( .A(KEYINPUT23), .B(n1203), .ZN(n1201) );
INV_X1 U882 ( .A(n1164), .ZN(n1200) );
NAND4_X1 U883 ( .A1(n1021), .A2(n1003), .A3(n1023), .A4(n1195), .ZN(n1164) );
NAND2_X1 U884 ( .A1(n1204), .A2(n997), .ZN(n1195) );
XOR2_X1 U885 ( .A(KEYINPUT52), .B(n1205), .Z(n1204) );
NOR3_X1 U886 ( .A1(n1066), .A2(n1206), .A3(n1037), .ZN(n1205) );
OR2_X1 U887 ( .A1(n1062), .A2(G900), .ZN(n1066) );
INV_X1 U888 ( .A(n1207), .ZN(n1023) );
XNOR2_X1 U889 ( .A(G122), .B(n1150), .ZN(G24) );
NAND3_X1 U890 ( .A1(n1186), .A2(n1025), .A3(n1208), .ZN(n1150) );
INV_X1 U891 ( .A(n1019), .ZN(n1025) );
NAND2_X1 U892 ( .A1(n1209), .A2(n1210), .ZN(n1019) );
INV_X1 U893 ( .A(n1174), .ZN(n1186) );
NAND2_X1 U894 ( .A1(n1211), .A2(n1212), .ZN(n1174) );
XOR2_X1 U895 ( .A(G119), .B(n1213), .Z(G21) );
NOR2_X1 U896 ( .A1(n1155), .A2(n1153), .ZN(n1213) );
NAND2_X1 U897 ( .A1(n1208), .A2(n1024), .ZN(n1153) );
NAND2_X1 U898 ( .A1(n1214), .A2(n1215), .ZN(n1155) );
XOR2_X1 U899 ( .A(G116), .B(n1216), .Z(G18) );
NOR2_X1 U900 ( .A1(KEYINPUT19), .A2(n1156), .ZN(n1216) );
NAND3_X1 U901 ( .A1(n1208), .A2(n1020), .A3(n1022), .ZN(n1156) );
AND2_X1 U902 ( .A1(n1217), .A2(n1218), .ZN(n1020) );
XOR2_X1 U903 ( .A(KEYINPUT21), .B(n1212), .Z(n1217) );
XOR2_X1 U904 ( .A(n1219), .B(KEYINPUT5), .Z(n1212) );
XOR2_X1 U905 ( .A(G113), .B(n1148), .Z(G15) );
AND3_X1 U906 ( .A1(n1022), .A2(n1208), .A3(n1021), .ZN(n1148) );
AND2_X1 U907 ( .A1(n1211), .A2(n1219), .ZN(n1021) );
INV_X1 U908 ( .A(n1218), .ZN(n1211) );
AND2_X1 U909 ( .A1(n1003), .A2(n1157), .ZN(n1208) );
NOR4_X1 U910 ( .A1(n1007), .A2(n1220), .A3(n1013), .A4(n1010), .ZN(n1003) );
INV_X1 U911 ( .A(n1221), .ZN(n1010) );
INV_X1 U912 ( .A(n1222), .ZN(n1013) );
INV_X1 U913 ( .A(n1191), .ZN(n1022) );
NAND2_X1 U914 ( .A1(n1215), .A2(n1210), .ZN(n1191) );
XNOR2_X1 U915 ( .A(n1223), .B(KEYINPUT54), .ZN(n1215) );
XOR2_X1 U916 ( .A(G110), .B(n1146), .Z(G12) );
NOR2_X1 U917 ( .A1(n1197), .A2(n1207), .ZN(n1146) );
NAND2_X1 U918 ( .A1(n1214), .A2(n1209), .ZN(n1207) );
XOR2_X1 U919 ( .A(n1223), .B(KEYINPUT36), .Z(n1209) );
XNOR2_X1 U920 ( .A(n1052), .B(KEYINPUT16), .ZN(n1223) );
XNOR2_X1 U921 ( .A(n1224), .B(G472), .ZN(n1052) );
NAND2_X1 U922 ( .A1(n1225), .A2(n1037), .ZN(n1224) );
XNOR2_X1 U923 ( .A(n1133), .B(n1226), .ZN(n1225) );
XOR2_X1 U924 ( .A(n1227), .B(n1117), .Z(n1226) );
NAND2_X1 U925 ( .A1(KEYINPUT44), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U926 ( .A(G101), .B(n1118), .ZN(n1228) );
NAND3_X1 U927 ( .A1(n1229), .A2(n1062), .A3(G210), .ZN(n1118) );
INV_X1 U928 ( .A(n1210), .ZN(n1214) );
XNOR2_X1 U929 ( .A(n1050), .B(n1230), .ZN(n1210) );
NOR2_X1 U930 ( .A1(n1056), .A2(KEYINPUT15), .ZN(n1230) );
NOR2_X1 U931 ( .A1(n1231), .A2(G902), .ZN(n1056) );
INV_X1 U932 ( .A(n1049), .ZN(n1231) );
XNOR2_X1 U933 ( .A(n1232), .B(n1233), .ZN(n1049) );
XOR2_X1 U934 ( .A(n1234), .B(n1235), .Z(n1233) );
NAND2_X1 U935 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
OR2_X1 U936 ( .A1(n1238), .A2(n1072), .ZN(n1237) );
XOR2_X1 U937 ( .A(n1239), .B(KEYINPUT28), .Z(n1236) );
NAND2_X1 U938 ( .A1(n1072), .A2(n1238), .ZN(n1239) );
NAND2_X1 U939 ( .A1(n1240), .A2(n1241), .ZN(n1238) );
NAND2_X1 U940 ( .A1(G140), .A2(n1203), .ZN(n1241) );
INV_X1 U941 ( .A(G125), .ZN(n1203) );
XOR2_X1 U942 ( .A(n1242), .B(KEYINPUT43), .Z(n1240) );
NAND2_X1 U943 ( .A1(G125), .A2(n1243), .ZN(n1242) );
INV_X1 U944 ( .A(G140), .ZN(n1243) );
NAND3_X1 U945 ( .A1(n1244), .A2(n1245), .A3(n1246), .ZN(n1234) );
NAND2_X1 U946 ( .A1(n1247), .A2(n1248), .ZN(n1246) );
NAND3_X1 U947 ( .A1(G234), .A2(n1062), .A3(G221), .ZN(n1248) );
NAND2_X1 U948 ( .A1(KEYINPUT62), .A2(n1249), .ZN(n1247) );
NAND4_X1 U949 ( .A1(KEYINPUT62), .A2(G221), .A3(n1250), .A4(n1251), .ZN(n1245) );
INV_X1 U950 ( .A(KEYINPUT17), .ZN(n1251) );
NOR3_X1 U951 ( .A1(n1252), .A2(G953), .A3(n1253), .ZN(n1250) );
NAND2_X1 U952 ( .A1(KEYINPUT17), .A2(n1253), .ZN(n1244) );
INV_X1 U953 ( .A(n1249), .ZN(n1253) );
XOR2_X1 U954 ( .A(G137), .B(KEYINPUT10), .Z(n1249) );
XOR2_X1 U955 ( .A(n1254), .B(n1255), .Z(n1232) );
NOR2_X1 U956 ( .A1(KEYINPUT56), .A2(n1256), .ZN(n1255) );
XOR2_X1 U957 ( .A(KEYINPUT4), .B(n1257), .Z(n1256) );
XNOR2_X1 U958 ( .A(G110), .B(G128), .ZN(n1254) );
NAND2_X1 U959 ( .A1(n1258), .A2(G217), .ZN(n1050) );
XOR2_X1 U960 ( .A(n1259), .B(KEYINPUT58), .Z(n1258) );
NAND3_X1 U961 ( .A1(n1158), .A2(n1157), .A3(n1024), .ZN(n1197) );
INV_X1 U962 ( .A(n1017), .ZN(n1024) );
NAND2_X1 U963 ( .A1(n1219), .A2(n1218), .ZN(n1017) );
XOR2_X1 U964 ( .A(G475), .B(n1260), .Z(n1218) );
NOR2_X1 U965 ( .A1(n1057), .A2(KEYINPUT37), .ZN(n1260) );
NOR2_X1 U966 ( .A1(n1261), .A2(G902), .ZN(n1057) );
INV_X1 U967 ( .A(n1045), .ZN(n1261) );
XNOR2_X1 U968 ( .A(n1262), .B(n1263), .ZN(n1045) );
XOR2_X1 U969 ( .A(n1264), .B(n1265), .Z(n1263) );
XNOR2_X1 U970 ( .A(n1192), .B(G113), .ZN(n1265) );
XNOR2_X1 U971 ( .A(KEYINPUT7), .B(n1184), .ZN(n1264) );
INV_X1 U972 ( .A(G143), .ZN(n1184) );
XOR2_X1 U973 ( .A(n1266), .B(n1267), .Z(n1262) );
XOR2_X1 U974 ( .A(n1268), .B(n1269), .Z(n1267) );
NOR2_X1 U975 ( .A1(G122), .A2(KEYINPUT33), .ZN(n1269) );
NOR3_X1 U976 ( .A1(n1270), .A2(G953), .A3(G237), .ZN(n1268) );
XOR2_X1 U977 ( .A(KEYINPUT14), .B(G214), .Z(n1270) );
XOR2_X1 U978 ( .A(n1271), .B(n1068), .Z(n1266) );
XOR2_X1 U979 ( .A(G140), .B(G125), .Z(n1068) );
XNOR2_X1 U980 ( .A(n1026), .B(KEYINPUT47), .ZN(n1219) );
XOR2_X1 U981 ( .A(n1272), .B(G478), .Z(n1026) );
NAND2_X1 U982 ( .A1(n1105), .A2(n1037), .ZN(n1272) );
XNOR2_X1 U983 ( .A(n1273), .B(n1274), .ZN(n1105) );
NOR3_X1 U984 ( .A1(n1252), .A2(G953), .A3(n1099), .ZN(n1274) );
INV_X1 U985 ( .A(G217), .ZN(n1099) );
NAND2_X1 U986 ( .A1(KEYINPUT35), .A2(n1275), .ZN(n1273) );
XOR2_X1 U987 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U988 ( .A(n1278), .B(n1279), .ZN(n1277) );
XOR2_X1 U989 ( .A(n1280), .B(G116), .Z(n1278) );
NAND2_X1 U990 ( .A1(KEYINPUT11), .A2(G107), .ZN(n1280) );
XNOR2_X1 U991 ( .A(G122), .B(n1281), .ZN(n1276) );
XNOR2_X1 U992 ( .A(KEYINPUT27), .B(n1076), .ZN(n1281) );
INV_X1 U993 ( .A(G134), .ZN(n1076) );
NAND2_X1 U994 ( .A1(n997), .A2(n1282), .ZN(n1157) );
NAND4_X1 U995 ( .A1(G953), .A2(G902), .A3(n1283), .A4(n1087), .ZN(n1282) );
INV_X1 U996 ( .A(G898), .ZN(n1087) );
NAND3_X1 U997 ( .A1(n1283), .A2(n1062), .A3(G952), .ZN(n997) );
INV_X1 U998 ( .A(n1206), .ZN(n1283) );
NOR2_X1 U999 ( .A1(n1229), .A2(n1252), .ZN(n1206) );
INV_X1 U1000 ( .A(G234), .ZN(n1252) );
INV_X1 U1001 ( .A(G237), .ZN(n1229) );
NOR2_X1 U1002 ( .A1(n1004), .A2(n1220), .ZN(n1158) );
INV_X1 U1003 ( .A(n1005), .ZN(n1220) );
XOR2_X1 U1004 ( .A(n1284), .B(n1048), .Z(n1005) );
NAND2_X1 U1005 ( .A1(G210), .A2(n1285), .ZN(n1048) );
NAND2_X1 U1006 ( .A1(KEYINPUT12), .A2(n1051), .ZN(n1284) );
NOR2_X1 U1007 ( .A1(n1286), .A2(G902), .ZN(n1051) );
INV_X1 U1008 ( .A(n1047), .ZN(n1286) );
XNOR2_X1 U1009 ( .A(n1287), .B(n1288), .ZN(n1047) );
XOR2_X1 U1010 ( .A(n1117), .B(n1095), .Z(n1288) );
XNOR2_X1 U1011 ( .A(n1289), .B(n1290), .ZN(n1095) );
XNOR2_X1 U1012 ( .A(n1291), .B(G110), .ZN(n1290) );
INV_X1 U1013 ( .A(G122), .ZN(n1291) );
NAND2_X1 U1014 ( .A1(n1292), .A2(n1293), .ZN(n1289) );
NAND2_X1 U1015 ( .A1(G101), .A2(n1294), .ZN(n1293) );
XOR2_X1 U1016 ( .A(n1295), .B(KEYINPUT32), .Z(n1292) );
OR2_X1 U1017 ( .A1(n1294), .A2(G101), .ZN(n1295) );
XOR2_X1 U1018 ( .A(G104), .B(G107), .Z(n1294) );
XNOR2_X1 U1019 ( .A(n1094), .B(n1296), .ZN(n1117) );
XOR2_X1 U1020 ( .A(G128), .B(n1297), .Z(n1296) );
NOR2_X1 U1021 ( .A1(KEYINPUT48), .A2(n1298), .ZN(n1297) );
XNOR2_X1 U1022 ( .A(G143), .B(n1072), .ZN(n1298) );
XOR2_X1 U1023 ( .A(n1299), .B(n1257), .Z(n1094) );
XOR2_X1 U1024 ( .A(G119), .B(KEYINPUT61), .Z(n1257) );
XNOR2_X1 U1025 ( .A(G113), .B(G116), .ZN(n1299) );
XNOR2_X1 U1026 ( .A(G125), .B(n1300), .ZN(n1287) );
NOR2_X1 U1027 ( .A1(G953), .A2(n1086), .ZN(n1300) );
INV_X1 U1028 ( .A(G224), .ZN(n1086) );
NAND3_X1 U1029 ( .A1(n1222), .A2(n1221), .A3(n1007), .ZN(n1004) );
XNOR2_X1 U1030 ( .A(n1032), .B(n1042), .ZN(n1007) );
INV_X1 U1031 ( .A(G469), .ZN(n1042) );
AND2_X1 U1032 ( .A1(n1044), .A2(n1037), .ZN(n1032) );
XNOR2_X1 U1033 ( .A(n1301), .B(n1302), .ZN(n1044) );
XNOR2_X1 U1034 ( .A(n1132), .B(n1114), .ZN(n1302) );
XOR2_X1 U1035 ( .A(G101), .B(n1133), .Z(n1114) );
XNOR2_X1 U1036 ( .A(n1303), .B(n1304), .ZN(n1133) );
NOR2_X1 U1037 ( .A1(KEYINPUT63), .A2(n1192), .ZN(n1304) );
INV_X1 U1038 ( .A(G131), .ZN(n1192) );
XNOR2_X1 U1039 ( .A(G134), .B(G137), .ZN(n1303) );
XOR2_X1 U1040 ( .A(n1305), .B(n1306), .Z(n1132) );
XOR2_X1 U1041 ( .A(KEYINPUT8), .B(G107), .Z(n1306) );
XOR2_X1 U1042 ( .A(n1271), .B(n1073), .Z(n1305) );
XNOR2_X1 U1043 ( .A(n1279), .B(KEYINPUT59), .ZN(n1073) );
XNOR2_X1 U1044 ( .A(G128), .B(G143), .ZN(n1279) );
XNOR2_X1 U1045 ( .A(G104), .B(n1072), .ZN(n1271) );
XOR2_X1 U1046 ( .A(G146), .B(KEYINPUT49), .Z(n1072) );
XOR2_X1 U1047 ( .A(n1307), .B(KEYINPUT55), .Z(n1301) );
NAND3_X1 U1048 ( .A1(n1308), .A2(n1309), .A3(n1125), .ZN(n1307) );
NAND2_X1 U1049 ( .A1(n1310), .A2(n1311), .ZN(n1125) );
NAND2_X1 U1050 ( .A1(n1310), .A2(n1312), .ZN(n1309) );
INV_X1 U1051 ( .A(KEYINPUT39), .ZN(n1312) );
NAND2_X1 U1052 ( .A1(n1127), .A2(KEYINPUT39), .ZN(n1308) );
NOR2_X1 U1053 ( .A1(n1311), .A2(n1310), .ZN(n1127) );
AND2_X1 U1054 ( .A1(G227), .A2(n1062), .ZN(n1310) );
INV_X1 U1055 ( .A(G953), .ZN(n1062) );
XNOR2_X1 U1056 ( .A(G110), .B(G140), .ZN(n1311) );
NAND2_X1 U1057 ( .A1(G214), .A2(n1285), .ZN(n1221) );
NAND2_X1 U1058 ( .A1(n1313), .A2(n1037), .ZN(n1285) );
XNOR2_X1 U1059 ( .A(G237), .B(KEYINPUT46), .ZN(n1313) );
NAND2_X1 U1060 ( .A1(G221), .A2(n1259), .ZN(n1222) );
NAND2_X1 U1061 ( .A1(G234), .A2(n1037), .ZN(n1259) );
INV_X1 U1062 ( .A(G902), .ZN(n1037) );
endmodule


