//Key = 1111101110101111110010011001010000010101010100000100001110111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
n1437, n1438, n1439, n1440, n1441, n1442;

XOR2_X1 U793 ( .A(G107), .B(n1097), .Z(G9) );
NOR2_X1 U794 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
NOR2_X1 U795 ( .A1(n1100), .A2(n1101), .ZN(G75) );
NOR3_X1 U796 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
NAND3_X1 U797 ( .A1(n1105), .A2(n1106), .A3(n1107), .ZN(n1102) );
NAND3_X1 U798 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1107) );
NAND2_X1 U799 ( .A1(n1111), .A2(n1112), .ZN(n1109) );
NAND3_X1 U800 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NAND2_X1 U801 ( .A1(n1116), .A2(n1117), .ZN(n1114) );
NAND2_X1 U802 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND3_X1 U803 ( .A1(n1120), .A2(n1121), .A3(n1119), .ZN(n1111) );
NAND3_X1 U804 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1120) );
NAND2_X1 U805 ( .A1(n1113), .A2(n1125), .ZN(n1124) );
OR2_X1 U806 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND3_X1 U807 ( .A1(n1128), .A2(n1115), .A3(n1129), .ZN(n1122) );
NAND4_X1 U808 ( .A1(n1119), .A2(n1121), .A3(n1130), .A4(n1131), .ZN(n1105) );
NAND2_X1 U809 ( .A1(KEYINPUT0), .A2(n1132), .ZN(n1131) );
NAND4_X1 U810 ( .A1(n1115), .A2(n1113), .A3(n1110), .A4(n1133), .ZN(n1132) );
NAND2_X1 U811 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NAND4_X1 U812 ( .A1(n1113), .A2(n1110), .A3(n1136), .A4(n1137), .ZN(n1130) );
INV_X1 U813 ( .A(KEYINPUT0), .ZN(n1137) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1138), .ZN(n1136) );
INV_X1 U815 ( .A(n1139), .ZN(n1110) );
NOR3_X1 U816 ( .A1(n1103), .A2(G952), .A3(n1140), .ZN(n1100) );
INV_X1 U817 ( .A(n1106), .ZN(n1140) );
NAND4_X1 U818 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1106) );
NOR4_X1 U819 ( .A1(n1145), .A2(n1118), .A3(n1146), .A4(n1147), .ZN(n1144) );
XOR2_X1 U820 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U821 ( .A1(KEYINPUT24), .A2(n1150), .ZN(n1148) );
NOR2_X1 U822 ( .A1(n1151), .A2(n1152), .ZN(n1146) );
XNOR2_X1 U823 ( .A(KEYINPUT16), .B(n1153), .ZN(n1152) );
INV_X1 U824 ( .A(n1154), .ZN(n1145) );
NOR3_X1 U825 ( .A1(n1155), .A2(n1156), .A3(n1157), .ZN(n1143) );
NOR2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
INV_X1 U827 ( .A(KEYINPUT48), .ZN(n1159) );
NOR3_X1 U828 ( .A1(n1160), .A2(n1161), .A3(n1129), .ZN(n1158) );
NOR2_X1 U829 ( .A1(KEYINPUT48), .A2(n1113), .ZN(n1156) );
XOR2_X1 U830 ( .A(n1162), .B(n1163), .Z(n1155) );
XOR2_X1 U831 ( .A(n1164), .B(n1165), .Z(G72) );
XOR2_X1 U832 ( .A(n1166), .B(n1167), .Z(n1165) );
NOR2_X1 U833 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
AND2_X1 U834 ( .A1(G227), .A2(G900), .ZN(n1168) );
NAND2_X1 U835 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
NAND2_X1 U836 ( .A1(G953), .A2(n1172), .ZN(n1171) );
XOR2_X1 U837 ( .A(n1173), .B(n1174), .Z(n1170) );
XOR2_X1 U838 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U839 ( .A1(KEYINPUT56), .A2(n1177), .ZN(n1176) );
XOR2_X1 U840 ( .A(n1178), .B(n1179), .Z(n1177) );
XOR2_X1 U841 ( .A(n1180), .B(G137), .Z(n1179) );
INV_X1 U842 ( .A(G134), .ZN(n1180) );
NAND2_X1 U843 ( .A1(KEYINPUT55), .A2(n1181), .ZN(n1178) );
XOR2_X1 U844 ( .A(n1182), .B(n1183), .Z(n1173) );
NAND2_X1 U845 ( .A1(KEYINPUT37), .A2(n1184), .ZN(n1182) );
NAND2_X1 U846 ( .A1(n1169), .A2(n1185), .ZN(n1164) );
NAND2_X1 U847 ( .A1(n1186), .A2(n1187), .ZN(G69) );
NAND2_X1 U848 ( .A1(n1188), .A2(n1169), .ZN(n1187) );
XNOR2_X1 U849 ( .A(n1189), .B(n1190), .ZN(n1188) );
NAND2_X1 U850 ( .A1(n1191), .A2(G953), .ZN(n1186) );
NAND2_X1 U851 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
NAND2_X1 U852 ( .A1(n1189), .A2(n1194), .ZN(n1193) );
INV_X1 U853 ( .A(G224), .ZN(n1194) );
NAND2_X1 U854 ( .A1(G224), .A2(n1195), .ZN(n1192) );
NAND2_X1 U855 ( .A1(G898), .A2(n1189), .ZN(n1195) );
NAND2_X1 U856 ( .A1(n1196), .A2(n1197), .ZN(n1189) );
NAND2_X1 U857 ( .A1(G953), .A2(n1198), .ZN(n1197) );
XOR2_X1 U858 ( .A(n1199), .B(n1200), .Z(n1196) );
XNOR2_X1 U859 ( .A(n1201), .B(n1202), .ZN(n1199) );
NOR2_X1 U860 ( .A1(n1203), .A2(n1204), .ZN(G66) );
XOR2_X1 U861 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U862 ( .A1(n1153), .A2(n1207), .ZN(n1205) );
NOR2_X1 U863 ( .A1(n1203), .A2(n1208), .ZN(G63) );
NOR3_X1 U864 ( .A1(n1149), .A2(n1209), .A3(n1210), .ZN(n1208) );
AND3_X1 U865 ( .A1(n1211), .A2(G478), .A3(n1212), .ZN(n1210) );
NOR2_X1 U866 ( .A1(n1213), .A2(n1211), .ZN(n1209) );
NOR2_X1 U867 ( .A1(n1214), .A2(n1150), .ZN(n1213) );
INV_X1 U868 ( .A(G478), .ZN(n1150) );
NOR2_X1 U869 ( .A1(n1203), .A2(n1215), .ZN(G60) );
XOR2_X1 U870 ( .A(n1216), .B(n1217), .Z(n1215) );
XOR2_X1 U871 ( .A(KEYINPUT2), .B(n1218), .Z(n1217) );
AND2_X1 U872 ( .A1(G475), .A2(n1212), .ZN(n1218) );
NAND2_X1 U873 ( .A1(n1219), .A2(n1220), .ZN(G6) );
NAND2_X1 U874 ( .A1(n1221), .A2(n1222), .ZN(n1220) );
NAND2_X1 U875 ( .A1(n1223), .A2(G104), .ZN(n1219) );
NAND2_X1 U876 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
NAND2_X1 U877 ( .A1(KEYINPUT28), .A2(n1226), .ZN(n1225) );
OR2_X1 U878 ( .A1(n1221), .A2(KEYINPUT28), .ZN(n1224) );
AND2_X1 U879 ( .A1(KEYINPUT20), .A2(n1226), .ZN(n1221) );
NOR2_X1 U880 ( .A1(n1203), .A2(n1227), .ZN(G57) );
XOR2_X1 U881 ( .A(n1228), .B(n1229), .Z(n1227) );
XOR2_X1 U882 ( .A(n1230), .B(n1231), .Z(n1229) );
XOR2_X1 U883 ( .A(n1232), .B(n1233), .Z(n1230) );
AND2_X1 U884 ( .A1(G472), .A2(n1212), .ZN(n1233) );
NAND2_X1 U885 ( .A1(n1234), .A2(KEYINPUT7), .ZN(n1232) );
XOR2_X1 U886 ( .A(n1235), .B(n1236), .Z(n1234) );
NOR2_X1 U887 ( .A1(KEYINPUT9), .A2(n1183), .ZN(n1236) );
XOR2_X1 U888 ( .A(n1237), .B(n1238), .Z(n1228) );
XOR2_X1 U889 ( .A(n1239), .B(KEYINPUT36), .Z(n1237) );
NOR2_X1 U890 ( .A1(n1203), .A2(n1240), .ZN(G54) );
XOR2_X1 U891 ( .A(n1241), .B(n1242), .Z(n1240) );
NOR2_X1 U892 ( .A1(n1160), .A2(n1207), .ZN(n1242) );
INV_X1 U893 ( .A(G469), .ZN(n1160) );
NOR3_X1 U894 ( .A1(n1243), .A2(n1244), .A3(n1245), .ZN(n1241) );
NOR2_X1 U895 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
AND3_X1 U896 ( .A1(n1247), .A2(n1246), .A3(n1248), .ZN(n1244) );
INV_X1 U897 ( .A(KEYINPUT44), .ZN(n1247) );
NOR2_X1 U898 ( .A1(n1249), .A2(n1248), .ZN(n1243) );
XNOR2_X1 U899 ( .A(n1250), .B(n1251), .ZN(n1248) );
NOR2_X1 U900 ( .A1(KEYINPUT44), .A2(n1252), .ZN(n1249) );
XOR2_X1 U901 ( .A(KEYINPUT15), .B(n1246), .Z(n1252) );
XNOR2_X1 U902 ( .A(n1253), .B(n1254), .ZN(n1246) );
NOR3_X1 U903 ( .A1(KEYINPUT52), .A2(n1255), .A3(n1256), .ZN(n1254) );
NOR2_X1 U904 ( .A1(n1175), .A2(n1257), .ZN(n1256) );
XOR2_X1 U905 ( .A(n1258), .B(KEYINPUT60), .Z(n1257) );
NOR2_X1 U906 ( .A1(G140), .A2(n1259), .ZN(n1255) );
XOR2_X1 U907 ( .A(n1258), .B(KEYINPUT30), .Z(n1259) );
NOR2_X1 U908 ( .A1(n1203), .A2(n1260), .ZN(G51) );
XOR2_X1 U909 ( .A(n1261), .B(n1262), .Z(n1260) );
XOR2_X1 U910 ( .A(n1263), .B(n1264), .Z(n1262) );
NAND3_X1 U911 ( .A1(n1212), .A2(n1265), .A3(KEYINPUT23), .ZN(n1263) );
INV_X1 U912 ( .A(n1207), .ZN(n1212) );
NAND2_X1 U913 ( .A1(G902), .A2(n1104), .ZN(n1207) );
INV_X1 U914 ( .A(n1214), .ZN(n1104) );
NOR2_X1 U915 ( .A1(n1185), .A2(n1190), .ZN(n1214) );
OR4_X1 U916 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1269), .ZN(n1190) );
OR4_X1 U917 ( .A1(n1270), .A2(n1271), .A3(n1272), .A4(n1226), .ZN(n1269) );
AND3_X1 U918 ( .A1(n1273), .A2(n1274), .A3(n1126), .ZN(n1226) );
NOR3_X1 U919 ( .A1(n1274), .A2(n1275), .A3(n1276), .ZN(n1271) );
INV_X1 U920 ( .A(KEYINPUT19), .ZN(n1276) );
NOR2_X1 U921 ( .A1(n1277), .A2(n1098), .ZN(n1270) );
NOR3_X1 U922 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
NOR2_X1 U923 ( .A1(KEYINPUT19), .A2(n1275), .ZN(n1280) );
NOR3_X1 U924 ( .A1(n1123), .A2(n1281), .A3(n1134), .ZN(n1279) );
INV_X1 U925 ( .A(n1282), .ZN(n1134) );
XNOR2_X1 U926 ( .A(KEYINPUT42), .B(n1099), .ZN(n1278) );
NAND2_X1 U927 ( .A1(n1127), .A2(n1273), .ZN(n1099) );
AND3_X1 U928 ( .A1(n1108), .A2(n1283), .A3(n1284), .ZN(n1273) );
NAND4_X1 U929 ( .A1(n1285), .A2(n1286), .A3(n1287), .A4(n1288), .ZN(n1185) );
NOR4_X1 U930 ( .A1(n1289), .A2(n1290), .A3(n1291), .A4(n1292), .ZN(n1288) );
NOR2_X1 U931 ( .A1(n1293), .A2(n1294), .ZN(n1287) );
NOR3_X1 U932 ( .A1(n1295), .A2(n1296), .A3(n1297), .ZN(n1294) );
XOR2_X1 U933 ( .A(n1298), .B(n1299), .Z(n1261) );
NAND2_X1 U934 ( .A1(KEYINPUT17), .A2(n1300), .ZN(n1299) );
INV_X1 U935 ( .A(n1301), .ZN(n1300) );
NOR2_X1 U936 ( .A1(n1169), .A2(G952), .ZN(n1203) );
XNOR2_X1 U937 ( .A(G146), .B(n1302), .ZN(G48) );
NOR2_X1 U938 ( .A1(KEYINPUT45), .A2(n1303), .ZN(n1302) );
NOR3_X1 U939 ( .A1(n1304), .A2(n1296), .A3(n1295), .ZN(n1303) );
INV_X1 U940 ( .A(n1305), .ZN(n1296) );
XOR2_X1 U941 ( .A(KEYINPUT41), .B(n1284), .Z(n1304) );
XNOR2_X1 U942 ( .A(G143), .B(n1285), .ZN(G45) );
NAND4_X1 U943 ( .A1(n1306), .A2(n1282), .A3(n1307), .A4(n1308), .ZN(n1285) );
XOR2_X1 U944 ( .A(n1175), .B(n1286), .Z(G42) );
NAND3_X1 U945 ( .A1(n1126), .A2(n1309), .A3(n1310), .ZN(n1286) );
XOR2_X1 U946 ( .A(G137), .B(n1292), .Z(G39) );
AND3_X1 U947 ( .A1(n1115), .A2(n1305), .A3(n1310), .ZN(n1292) );
XOR2_X1 U948 ( .A(G134), .B(n1291), .Z(G36) );
AND3_X1 U949 ( .A1(n1127), .A2(n1282), .A3(n1310), .ZN(n1291) );
XOR2_X1 U950 ( .A(G131), .B(n1290), .Z(G33) );
AND3_X1 U951 ( .A1(n1126), .A2(n1282), .A3(n1310), .ZN(n1290) );
AND4_X1 U952 ( .A1(n1284), .A2(n1119), .A3(n1311), .A4(n1121), .ZN(n1310) );
XOR2_X1 U953 ( .A(G128), .B(n1289), .Z(G30) );
AND3_X1 U954 ( .A1(n1127), .A2(n1305), .A3(n1306), .ZN(n1289) );
AND3_X1 U955 ( .A1(n1284), .A2(n1311), .A3(n1312), .ZN(n1306) );
XOR2_X1 U956 ( .A(n1313), .B(n1314), .Z(G3) );
NAND2_X1 U957 ( .A1(KEYINPUT3), .A2(G101), .ZN(n1314) );
NAND4_X1 U958 ( .A1(n1274), .A2(n1283), .A3(n1282), .A4(n1315), .ZN(n1313) );
NOR2_X1 U959 ( .A1(n1316), .A2(n1138), .ZN(n1315) );
INV_X1 U960 ( .A(n1115), .ZN(n1138) );
XOR2_X1 U961 ( .A(n1297), .B(KEYINPUT50), .Z(n1316) );
INV_X1 U962 ( .A(n1284), .ZN(n1297) );
INV_X1 U963 ( .A(n1098), .ZN(n1274) );
XOR2_X1 U964 ( .A(G125), .B(n1293), .Z(G27) );
NOR3_X1 U965 ( .A1(n1135), .A2(n1317), .A3(n1295), .ZN(n1293) );
NAND3_X1 U966 ( .A1(n1312), .A2(n1311), .A3(n1126), .ZN(n1295) );
NAND2_X1 U967 ( .A1(n1139), .A2(n1318), .ZN(n1311) );
NAND4_X1 U968 ( .A1(G953), .A2(G902), .A3(n1319), .A4(n1172), .ZN(n1318) );
INV_X1 U969 ( .A(G900), .ZN(n1172) );
XOR2_X1 U970 ( .A(G122), .B(n1272), .Z(G24) );
AND4_X1 U971 ( .A1(n1320), .A2(n1108), .A3(n1307), .A4(n1308), .ZN(n1272) );
XOR2_X1 U972 ( .A(G119), .B(n1268), .Z(G21) );
AND3_X1 U973 ( .A1(n1115), .A2(n1305), .A3(n1320), .ZN(n1268) );
NAND2_X1 U974 ( .A1(n1321), .A2(n1322), .ZN(n1305) );
NAND3_X1 U975 ( .A1(n1323), .A2(n1324), .A3(n1325), .ZN(n1322) );
INV_X1 U976 ( .A(KEYINPUT26), .ZN(n1325) );
NAND2_X1 U977 ( .A1(KEYINPUT26), .A2(n1309), .ZN(n1321) );
INV_X1 U978 ( .A(n1135), .ZN(n1309) );
XOR2_X1 U979 ( .A(G116), .B(n1266), .Z(G18) );
AND3_X1 U980 ( .A1(n1127), .A2(n1282), .A3(n1320), .ZN(n1266) );
NOR3_X1 U981 ( .A1(n1116), .A2(n1281), .A3(n1317), .ZN(n1320) );
AND2_X1 U982 ( .A1(n1141), .A2(n1308), .ZN(n1127) );
XOR2_X1 U983 ( .A(G113), .B(n1326), .Z(G15) );
NOR2_X1 U984 ( .A1(n1098), .A2(n1275), .ZN(n1326) );
NAND4_X1 U985 ( .A1(n1126), .A2(n1113), .A3(n1282), .A4(n1283), .ZN(n1275) );
NAND2_X1 U986 ( .A1(n1327), .A2(n1328), .ZN(n1282) );
OR3_X1 U987 ( .A1(n1324), .A2(n1142), .A3(KEYINPUT26), .ZN(n1328) );
NAND2_X1 U988 ( .A1(KEYINPUT26), .A2(n1108), .ZN(n1327) );
NOR2_X1 U989 ( .A1(n1324), .A2(n1323), .ZN(n1108) );
INV_X1 U990 ( .A(n1142), .ZN(n1323) );
INV_X1 U991 ( .A(n1317), .ZN(n1113) );
NAND2_X1 U992 ( .A1(n1128), .A2(n1329), .ZN(n1317) );
NOR2_X1 U993 ( .A1(n1308), .A2(n1141), .ZN(n1126) );
NAND2_X1 U994 ( .A1(n1330), .A2(n1331), .ZN(G12) );
NAND2_X1 U995 ( .A1(n1267), .A2(n1258), .ZN(n1331) );
XOR2_X1 U996 ( .A(KEYINPUT10), .B(n1332), .Z(n1330) );
NOR2_X1 U997 ( .A1(n1267), .A2(n1258), .ZN(n1332) );
NOR4_X1 U998 ( .A1(n1123), .A2(n1135), .A3(n1098), .A4(n1281), .ZN(n1267) );
INV_X1 U999 ( .A(n1283), .ZN(n1281) );
NAND2_X1 U1000 ( .A1(n1139), .A2(n1333), .ZN(n1283) );
NAND4_X1 U1001 ( .A1(G953), .A2(G902), .A3(n1319), .A4(n1198), .ZN(n1333) );
INV_X1 U1002 ( .A(G898), .ZN(n1198) );
NAND3_X1 U1003 ( .A1(n1334), .A2(n1319), .A3(G952), .ZN(n1139) );
NAND2_X1 U1004 ( .A1(G237), .A2(G234), .ZN(n1319) );
INV_X1 U1005 ( .A(n1103), .ZN(n1334) );
XOR2_X1 U1006 ( .A(n1169), .B(KEYINPUT6), .Z(n1103) );
XOR2_X1 U1007 ( .A(n1116), .B(KEYINPUT33), .Z(n1098) );
INV_X1 U1008 ( .A(n1312), .ZN(n1116) );
NOR2_X1 U1009 ( .A1(n1119), .A2(n1118), .ZN(n1312) );
INV_X1 U1010 ( .A(n1121), .ZN(n1118) );
NAND2_X1 U1011 ( .A1(G214), .A2(n1335), .ZN(n1121) );
XNOR2_X1 U1012 ( .A(n1336), .B(n1265), .ZN(n1119) );
INV_X1 U1013 ( .A(n1162), .ZN(n1265) );
NAND2_X1 U1014 ( .A1(G210), .A2(n1335), .ZN(n1162) );
NAND2_X1 U1015 ( .A1(n1337), .A2(n1338), .ZN(n1335) );
INV_X1 U1016 ( .A(G237), .ZN(n1337) );
NAND2_X1 U1017 ( .A1(KEYINPUT59), .A2(n1163), .ZN(n1336) );
NAND4_X1 U1018 ( .A1(n1339), .A2(n1338), .A3(n1340), .A4(n1341), .ZN(n1163) );
NAND2_X1 U1019 ( .A1(KEYINPUT53), .A2(n1342), .ZN(n1341) );
NAND2_X1 U1020 ( .A1(n1343), .A2(n1298), .ZN(n1342) );
XNOR2_X1 U1021 ( .A(KEYINPUT54), .B(n1344), .ZN(n1343) );
NAND2_X1 U1022 ( .A1(n1345), .A2(n1346), .ZN(n1340) );
INV_X1 U1023 ( .A(KEYINPUT53), .ZN(n1346) );
NAND2_X1 U1024 ( .A1(n1347), .A2(n1348), .ZN(n1345) );
OR2_X1 U1025 ( .A1(n1344), .A2(KEYINPUT54), .ZN(n1348) );
NAND3_X1 U1026 ( .A1(n1344), .A2(n1298), .A3(KEYINPUT54), .ZN(n1347) );
OR2_X1 U1027 ( .A1(n1298), .A2(n1344), .ZN(n1339) );
XNOR2_X1 U1028 ( .A(n1264), .B(n1349), .ZN(n1344) );
NOR2_X1 U1029 ( .A1(KEYINPUT18), .A2(n1301), .ZN(n1349) );
NAND2_X1 U1030 ( .A1(G224), .A2(n1169), .ZN(n1301) );
XOR2_X1 U1031 ( .A(n1184), .B(n1183), .Z(n1264) );
NAND2_X1 U1032 ( .A1(n1350), .A2(n1351), .ZN(n1298) );
NAND2_X1 U1033 ( .A1(n1200), .A2(n1352), .ZN(n1351) );
XOR2_X1 U1034 ( .A(KEYINPUT39), .B(n1353), .Z(n1350) );
NOR2_X1 U1035 ( .A1(n1200), .A2(n1352), .ZN(n1353) );
NAND2_X1 U1036 ( .A1(n1354), .A2(n1355), .ZN(n1352) );
NAND2_X1 U1037 ( .A1(n1202), .A2(n1201), .ZN(n1355) );
XOR2_X1 U1038 ( .A(KEYINPUT63), .B(n1356), .Z(n1354) );
NOR2_X1 U1039 ( .A1(n1201), .A2(n1202), .ZN(n1356) );
AND2_X1 U1040 ( .A1(n1357), .A2(n1358), .ZN(n1202) );
NAND2_X1 U1041 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
XOR2_X1 U1042 ( .A(KEYINPUT62), .B(n1361), .Z(n1357) );
NOR2_X1 U1043 ( .A1(n1359), .A2(n1360), .ZN(n1361) );
INV_X1 U1044 ( .A(G113), .ZN(n1360) );
AND2_X1 U1045 ( .A1(n1362), .A2(n1363), .ZN(n1359) );
OR2_X1 U1046 ( .A1(n1364), .A2(G119), .ZN(n1363) );
XOR2_X1 U1047 ( .A(n1365), .B(KEYINPUT40), .Z(n1362) );
NAND2_X1 U1048 ( .A1(G119), .A2(n1364), .ZN(n1365) );
AND2_X1 U1049 ( .A1(n1366), .A2(n1367), .ZN(n1201) );
NAND2_X1 U1050 ( .A1(n1368), .A2(n1239), .ZN(n1367) );
XNOR2_X1 U1051 ( .A(n1369), .B(n1370), .ZN(n1368) );
XOR2_X1 U1052 ( .A(n1371), .B(KEYINPUT32), .Z(n1366) );
NAND2_X1 U1053 ( .A1(n1372), .A2(G101), .ZN(n1371) );
XOR2_X1 U1054 ( .A(n1369), .B(n1370), .Z(n1372) );
NAND2_X1 U1055 ( .A1(KEYINPUT61), .A2(G104), .ZN(n1369) );
XNOR2_X1 U1056 ( .A(n1373), .B(n1374), .ZN(n1200) );
NAND2_X1 U1057 ( .A1(KEYINPUT1), .A2(n1258), .ZN(n1373) );
NAND2_X1 U1058 ( .A1(n1142), .A2(n1324), .ZN(n1135) );
NAND2_X1 U1059 ( .A1(n1375), .A2(n1154), .ZN(n1324) );
NAND2_X1 U1060 ( .A1(n1151), .A2(n1153), .ZN(n1154) );
OR2_X1 U1061 ( .A1(n1153), .A2(n1151), .ZN(n1375) );
NOR2_X1 U1062 ( .A1(n1206), .A2(G902), .ZN(n1151) );
XNOR2_X1 U1063 ( .A(n1376), .B(n1377), .ZN(n1206) );
XOR2_X1 U1064 ( .A(n1378), .B(n1379), .Z(n1377) );
XOR2_X1 U1065 ( .A(G137), .B(G119), .Z(n1379) );
XOR2_X1 U1066 ( .A(KEYINPUT49), .B(KEYINPUT25), .Z(n1378) );
XOR2_X1 U1067 ( .A(n1380), .B(n1381), .Z(n1376) );
XOR2_X1 U1068 ( .A(n1258), .B(n1382), .Z(n1381) );
NAND3_X1 U1069 ( .A1(G234), .A2(n1169), .A3(G221), .ZN(n1382) );
XNOR2_X1 U1070 ( .A(n1383), .B(n1384), .ZN(n1380) );
NAND2_X1 U1071 ( .A1(G217), .A2(n1385), .ZN(n1153) );
XOR2_X1 U1072 ( .A(n1386), .B(G472), .Z(n1142) );
NAND2_X1 U1073 ( .A1(n1387), .A2(n1338), .ZN(n1386) );
XOR2_X1 U1074 ( .A(n1388), .B(n1389), .Z(n1387) );
XOR2_X1 U1075 ( .A(n1390), .B(n1231), .Z(n1389) );
XOR2_X1 U1076 ( .A(G113), .B(n1391), .Z(n1231) );
XOR2_X1 U1077 ( .A(G119), .B(G116), .Z(n1391) );
NOR2_X1 U1078 ( .A1(KEYINPUT34), .A2(n1392), .ZN(n1390) );
XNOR2_X1 U1079 ( .A(n1251), .B(n1393), .ZN(n1388) );
NOR2_X1 U1080 ( .A1(n1394), .A2(n1395), .ZN(n1393) );
NOR2_X1 U1081 ( .A1(KEYINPUT27), .A2(n1238), .ZN(n1395) );
AND2_X1 U1082 ( .A1(KEYINPUT4), .A2(n1238), .ZN(n1394) );
AND2_X1 U1083 ( .A1(G210), .A2(n1396), .ZN(n1238) );
XNOR2_X1 U1084 ( .A(n1239), .B(n1183), .ZN(n1251) );
NAND2_X1 U1085 ( .A1(n1115), .A2(n1284), .ZN(n1123) );
NOR2_X1 U1086 ( .A1(n1128), .A2(n1129), .ZN(n1284) );
INV_X1 U1087 ( .A(n1329), .ZN(n1129) );
NAND2_X1 U1088 ( .A1(G221), .A2(n1385), .ZN(n1329) );
NAND2_X1 U1089 ( .A1(G234), .A2(n1338), .ZN(n1385) );
XNOR2_X1 U1090 ( .A(n1161), .B(G469), .ZN(n1128) );
AND2_X1 U1091 ( .A1(n1338), .A2(n1397), .ZN(n1161) );
NAND2_X1 U1092 ( .A1(n1398), .A2(n1399), .ZN(n1397) );
NAND2_X1 U1093 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
XOR2_X1 U1094 ( .A(n1402), .B(n1403), .Z(n1401) );
INV_X1 U1095 ( .A(n1250), .ZN(n1402) );
XOR2_X1 U1096 ( .A(n1253), .B(n1404), .Z(n1400) );
XOR2_X1 U1097 ( .A(n1405), .B(KEYINPUT46), .Z(n1398) );
NAND2_X1 U1098 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
XNOR2_X1 U1099 ( .A(n1404), .B(n1253), .ZN(n1407) );
NAND2_X1 U1100 ( .A1(G227), .A2(n1169), .ZN(n1253) );
NOR2_X1 U1101 ( .A1(KEYINPUT57), .A2(n1408), .ZN(n1404) );
XOR2_X1 U1102 ( .A(n1258), .B(n1409), .Z(n1408) );
XOR2_X1 U1103 ( .A(KEYINPUT51), .B(G140), .Z(n1409) );
INV_X1 U1104 ( .A(G110), .ZN(n1258) );
XOR2_X1 U1105 ( .A(n1250), .B(n1403), .Z(n1406) );
XOR2_X1 U1106 ( .A(n1410), .B(n1239), .Z(n1403) );
INV_X1 U1107 ( .A(G101), .ZN(n1239) );
NAND2_X1 U1108 ( .A1(KEYINPUT29), .A2(n1183), .ZN(n1410) );
XOR2_X1 U1109 ( .A(G143), .B(n1383), .Z(n1183) );
XNOR2_X1 U1110 ( .A(G128), .B(n1411), .ZN(n1383) );
XOR2_X1 U1111 ( .A(n1412), .B(n1392), .Z(n1250) );
INV_X1 U1112 ( .A(n1235), .ZN(n1392) );
XOR2_X1 U1113 ( .A(n1413), .B(n1414), .Z(n1235) );
XOR2_X1 U1114 ( .A(G134), .B(n1415), .Z(n1414) );
NOR2_X1 U1115 ( .A1(KEYINPUT31), .A2(n1416), .ZN(n1415) );
INV_X1 U1116 ( .A(G137), .ZN(n1416) );
NAND2_X1 U1117 ( .A1(KEYINPUT12), .A2(n1181), .ZN(n1413) );
NAND2_X1 U1118 ( .A1(n1417), .A2(n1418), .ZN(n1412) );
NAND2_X1 U1119 ( .A1(n1419), .A2(n1222), .ZN(n1418) );
XOR2_X1 U1120 ( .A(KEYINPUT8), .B(n1420), .Z(n1417) );
NOR2_X1 U1121 ( .A1(n1419), .A2(n1222), .ZN(n1420) );
INV_X1 U1122 ( .A(G104), .ZN(n1222) );
XNOR2_X1 U1123 ( .A(KEYINPUT21), .B(n1370), .ZN(n1419) );
NOR2_X1 U1124 ( .A1(n1308), .A2(n1307), .ZN(n1115) );
INV_X1 U1125 ( .A(n1141), .ZN(n1307) );
XOR2_X1 U1126 ( .A(n1421), .B(G475), .Z(n1141) );
NAND2_X1 U1127 ( .A1(n1216), .A2(n1338), .ZN(n1421) );
INV_X1 U1128 ( .A(G902), .ZN(n1338) );
XOR2_X1 U1129 ( .A(n1422), .B(n1423), .Z(n1216) );
XOR2_X1 U1130 ( .A(n1424), .B(n1425), .Z(n1423) );
NOR2_X1 U1131 ( .A1(G113), .A2(KEYINPUT22), .ZN(n1425) );
AND2_X1 U1132 ( .A1(n1396), .A2(G214), .ZN(n1424) );
AND2_X1 U1133 ( .A1(n1426), .A2(n1169), .ZN(n1396) );
INV_X1 U1134 ( .A(G953), .ZN(n1169) );
XOR2_X1 U1135 ( .A(KEYINPUT14), .B(G237), .Z(n1426) );
XOR2_X1 U1136 ( .A(n1427), .B(n1428), .Z(n1422) );
NOR2_X1 U1137 ( .A1(KEYINPUT5), .A2(n1411), .ZN(n1428) );
XNOR2_X1 U1138 ( .A(G146), .B(KEYINPUT47), .ZN(n1411) );
XOR2_X1 U1139 ( .A(n1429), .B(n1430), .Z(n1427) );
XOR2_X1 U1140 ( .A(G104), .B(n1431), .Z(n1430) );
XOR2_X1 U1141 ( .A(KEYINPUT35), .B(G143), .Z(n1431) );
XNOR2_X1 U1142 ( .A(n1384), .B(n1432), .ZN(n1429) );
XOR2_X1 U1143 ( .A(n1433), .B(n1374), .Z(n1432) );
NOR2_X1 U1144 ( .A1(KEYINPUT11), .A2(n1181), .ZN(n1433) );
INV_X1 U1145 ( .A(G131), .ZN(n1181) );
XOR2_X1 U1146 ( .A(n1184), .B(n1175), .Z(n1384) );
INV_X1 U1147 ( .A(G140), .ZN(n1175) );
INV_X1 U1148 ( .A(G125), .ZN(n1184) );
XOR2_X1 U1149 ( .A(n1149), .B(G478), .Z(n1308) );
NOR2_X1 U1150 ( .A1(n1211), .A2(G902), .ZN(n1149) );
XNOR2_X1 U1151 ( .A(n1434), .B(n1435), .ZN(n1211) );
XOR2_X1 U1152 ( .A(G128), .B(n1436), .Z(n1435) );
XOR2_X1 U1153 ( .A(G143), .B(G134), .Z(n1436) );
XOR2_X1 U1154 ( .A(n1437), .B(n1370), .Z(n1434) );
XOR2_X1 U1155 ( .A(G107), .B(KEYINPUT13), .Z(n1370) );
XOR2_X1 U1156 ( .A(n1438), .B(n1439), .Z(n1437) );
NOR3_X1 U1157 ( .A1(n1440), .A2(G953), .A3(n1441), .ZN(n1439) );
XNOR2_X1 U1158 ( .A(G234), .B(KEYINPUT38), .ZN(n1441) );
INV_X1 U1159 ( .A(G217), .ZN(n1440) );
NAND2_X1 U1160 ( .A1(n1442), .A2(KEYINPUT58), .ZN(n1438) );
XOR2_X1 U1161 ( .A(n1364), .B(n1374), .Z(n1442) );
XOR2_X1 U1162 ( .A(G122), .B(KEYINPUT43), .Z(n1374) );
INV_X1 U1163 ( .A(G116), .ZN(n1364) );
endmodule


