//Key = 1110001100100100110001100001001100001101101011100011010111100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334;

XOR2_X1 U737 ( .A(n1024), .B(n1025), .Z(G9) );
NOR2_X1 U738 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR4_X1 U739 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1027) );
NOR2_X1 U740 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
AND4_X1 U741 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1032) );
NAND4_X1 U742 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1028) );
NAND3_X1 U743 ( .A1(n1034), .A2(n1042), .A3(n1036), .ZN(n1039) );
NAND2_X1 U744 ( .A1(n1035), .A2(n1043), .ZN(n1038) );
NAND2_X1 U745 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U746 ( .A1(n1046), .A2(n1047), .A3(n1036), .ZN(n1045) );
NOR3_X1 U747 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n1036) );
NAND2_X1 U748 ( .A1(n1037), .A2(n1051), .ZN(n1047) );
NAND2_X1 U749 ( .A1(n1034), .A2(n1033), .ZN(n1051) );
INV_X1 U750 ( .A(KEYINPUT11), .ZN(n1033) );
OR3_X1 U751 ( .A1(n1052), .A2(n1053), .A3(n1037), .ZN(n1046) );
NAND4_X1 U752 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1044) );
NOR3_X1 U753 ( .A1(n1050), .A2(n1058), .A3(n1059), .ZN(n1057) );
NOR2_X1 U754 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NAND2_X1 U755 ( .A1(n1048), .A2(n1049), .ZN(n1056) );
OR4_X1 U756 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1060), .ZN(n1054) );
NOR3_X1 U757 ( .A1(n1065), .A2(G953), .A3(G952), .ZN(n1026) );
INV_X1 U758 ( .A(n1040), .ZN(n1065) );
NAND4_X1 U759 ( .A1(n1066), .A2(n1067), .A3(n1068), .A4(n1069), .ZN(n1040) );
NOR4_X1 U760 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1069) );
XOR2_X1 U761 ( .A(G478), .B(n1074), .Z(n1073) );
XNOR2_X1 U762 ( .A(n1075), .B(n1076), .ZN(n1072) );
XOR2_X1 U763 ( .A(n1077), .B(KEYINPUT62), .Z(n1076) );
XOR2_X1 U764 ( .A(n1078), .B(n1079), .Z(n1071) );
NOR2_X1 U765 ( .A1(KEYINPUT19), .A2(n1080), .ZN(n1079) );
XOR2_X1 U766 ( .A(n1081), .B(G475), .Z(n1070) );
NAND2_X1 U767 ( .A1(KEYINPUT1), .A2(n1082), .ZN(n1081) );
INV_X1 U768 ( .A(n1083), .ZN(n1082) );
NOR2_X1 U769 ( .A1(n1064), .A2(n1037), .ZN(n1068) );
XNOR2_X1 U770 ( .A(n1084), .B(n1085), .ZN(n1066) );
NOR2_X1 U771 ( .A1(n1086), .A2(KEYINPUT43), .ZN(n1085) );
XOR2_X1 U772 ( .A(n1087), .B(n1088), .Z(G72) );
XOR2_X1 U773 ( .A(n1089), .B(n1090), .Z(n1088) );
NOR2_X1 U774 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U775 ( .A(n1041), .B(KEYINPUT16), .Z(n1092) );
NOR2_X1 U776 ( .A1(n1093), .A2(n1094), .ZN(n1091) );
NAND2_X1 U777 ( .A1(n1095), .A2(n1096), .ZN(n1089) );
NAND2_X1 U778 ( .A1(G953), .A2(n1097), .ZN(n1096) );
XOR2_X1 U779 ( .A(n1098), .B(n1099), .Z(n1095) );
XOR2_X1 U780 ( .A(n1100), .B(n1101), .Z(n1099) );
XOR2_X1 U781 ( .A(n1102), .B(n1103), .Z(n1098) );
NOR2_X1 U782 ( .A1(G131), .A2(KEYINPUT49), .ZN(n1103) );
XOR2_X1 U783 ( .A(n1104), .B(KEYINPUT45), .Z(n1102) );
NAND2_X1 U784 ( .A1(G953), .A2(n1105), .ZN(n1087) );
NAND2_X1 U785 ( .A1(G900), .A2(G227), .ZN(n1105) );
XOR2_X1 U786 ( .A(n1106), .B(n1107), .Z(G69) );
XOR2_X1 U787 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U788 ( .A1(KEYINPUT32), .A2(n1110), .ZN(n1109) );
NOR2_X1 U789 ( .A1(n1111), .A2(n1041), .ZN(n1110) );
AND2_X1 U790 ( .A1(G224), .A2(G898), .ZN(n1111) );
NOR2_X1 U791 ( .A1(n1112), .A2(n1113), .ZN(n1108) );
XOR2_X1 U792 ( .A(KEYINPUT18), .B(G953), .Z(n1113) );
NOR2_X1 U793 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NAND2_X1 U794 ( .A1(n1116), .A2(n1117), .ZN(n1106) );
NAND2_X1 U795 ( .A1(G953), .A2(n1118), .ZN(n1117) );
XOR2_X1 U796 ( .A(KEYINPUT2), .B(G898), .Z(n1118) );
XNOR2_X1 U797 ( .A(n1119), .B(n1120), .ZN(n1116) );
NOR3_X1 U798 ( .A1(n1121), .A2(n1122), .A3(n1123), .ZN(G66) );
NOR3_X1 U799 ( .A1(n1124), .A2(n1125), .A3(n1080), .ZN(n1123) );
NOR2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1121) );
XNOR2_X1 U801 ( .A(KEYINPUT3), .B(n1125), .ZN(n1127) );
NOR2_X1 U802 ( .A1(n1080), .A2(n1124), .ZN(n1126) );
NOR2_X1 U803 ( .A1(n1122), .A2(n1128), .ZN(G63) );
XOR2_X1 U804 ( .A(n1129), .B(n1130), .Z(n1128) );
NOR2_X1 U805 ( .A1(n1131), .A2(KEYINPUT60), .ZN(n1129) );
NOR2_X1 U806 ( .A1(n1132), .A2(n1124), .ZN(n1131) );
NOR2_X1 U807 ( .A1(n1122), .A2(n1133), .ZN(G60) );
XOR2_X1 U808 ( .A(n1134), .B(n1135), .Z(n1133) );
XOR2_X1 U809 ( .A(KEYINPUT35), .B(n1136), .Z(n1135) );
NOR2_X1 U810 ( .A1(n1137), .A2(n1124), .ZN(n1136) );
INV_X1 U811 ( .A(G475), .ZN(n1137) );
XOR2_X1 U812 ( .A(G104), .B(n1138), .Z(G6) );
NOR3_X1 U813 ( .A1(n1139), .A2(n1059), .A3(n1140), .ZN(n1138) );
INV_X1 U814 ( .A(n1034), .ZN(n1059) );
XOR2_X1 U815 ( .A(KEYINPUT6), .B(n1062), .Z(n1139) );
NOR3_X1 U816 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(G57) );
NOR3_X1 U817 ( .A1(n1144), .A2(G953), .A3(G952), .ZN(n1143) );
AND2_X1 U818 ( .A1(n1144), .A2(n1122), .ZN(n1142) );
INV_X1 U819 ( .A(KEYINPUT23), .ZN(n1144) );
XOR2_X1 U820 ( .A(n1145), .B(n1146), .Z(n1141) );
XOR2_X1 U821 ( .A(n1147), .B(n1148), .Z(n1146) );
NAND2_X1 U822 ( .A1(KEYINPUT27), .A2(G101), .ZN(n1147) );
XNOR2_X1 U823 ( .A(n1149), .B(n1150), .ZN(n1145) );
XOR2_X1 U824 ( .A(n1151), .B(n1152), .Z(n1150) );
NOR2_X1 U825 ( .A1(n1153), .A2(n1124), .ZN(n1152) );
INV_X1 U826 ( .A(G472), .ZN(n1153) );
NOR2_X1 U827 ( .A1(KEYINPUT47), .A2(n1154), .ZN(n1151) );
XOR2_X1 U828 ( .A(n1155), .B(n1156), .Z(n1154) );
NOR2_X1 U829 ( .A1(KEYINPUT61), .A2(n1157), .ZN(n1155) );
NOR2_X1 U830 ( .A1(n1122), .A2(n1158), .ZN(G54) );
XOR2_X1 U831 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U832 ( .A(n1161), .B(n1156), .Z(n1160) );
NAND2_X1 U833 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
NAND2_X1 U834 ( .A1(n1164), .A2(n1165), .ZN(n1163) );
NAND2_X1 U835 ( .A1(KEYINPUT36), .A2(n1166), .ZN(n1165) );
NAND3_X1 U836 ( .A1(KEYINPUT36), .A2(n1166), .A3(n1167), .ZN(n1162) );
XOR2_X1 U837 ( .A(n1168), .B(n1169), .Z(n1159) );
NOR2_X1 U838 ( .A1(n1077), .A2(n1124), .ZN(n1169) );
NAND4_X1 U839 ( .A1(KEYINPUT51), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(n1168) );
NAND3_X1 U840 ( .A1(KEYINPUT57), .A2(n1173), .A3(n1104), .ZN(n1172) );
NAND2_X1 U841 ( .A1(n1174), .A2(n1175), .ZN(n1171) );
NAND2_X1 U842 ( .A1(KEYINPUT57), .A2(n1176), .ZN(n1175) );
XOR2_X1 U843 ( .A(KEYINPUT28), .B(n1173), .Z(n1176) );
INV_X1 U844 ( .A(n1104), .ZN(n1174) );
OR2_X1 U845 ( .A1(n1173), .A2(KEYINPUT57), .ZN(n1170) );
NOR2_X1 U846 ( .A1(n1122), .A2(n1177), .ZN(G51) );
XOR2_X1 U847 ( .A(n1178), .B(n1179), .Z(n1177) );
XNOR2_X1 U848 ( .A(n1180), .B(n1181), .ZN(n1179) );
NOR2_X1 U849 ( .A1(n1084), .A2(n1124), .ZN(n1181) );
NAND2_X1 U850 ( .A1(G902), .A2(n1182), .ZN(n1124) );
OR2_X1 U851 ( .A1(n1029), .A2(n1031), .ZN(n1182) );
XOR2_X1 U852 ( .A(n1115), .B(KEYINPUT15), .Z(n1031) );
NAND4_X1 U853 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1115) );
OR3_X1 U854 ( .A1(n1094), .A2(n1114), .A3(n1187), .ZN(n1029) );
XOR2_X1 U855 ( .A(n1093), .B(KEYINPUT8), .Z(n1187) );
NAND4_X1 U856 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1025), .ZN(n1114) );
NAND3_X1 U857 ( .A1(n1034), .A2(n1063), .A3(n1191), .ZN(n1025) );
NAND3_X1 U858 ( .A1(n1191), .A2(n1034), .A3(n1062), .ZN(n1188) );
NAND4_X1 U859 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1094) );
NOR4_X1 U860 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1195) );
INV_X1 U861 ( .A(n1200), .ZN(n1199) );
NAND3_X1 U862 ( .A1(n1063), .A2(n1060), .A3(n1201), .ZN(n1194) );
XOR2_X1 U863 ( .A(n1202), .B(n1203), .Z(n1178) );
XOR2_X1 U864 ( .A(n1157), .B(G125), .Z(n1202) );
NOR2_X1 U865 ( .A1(n1041), .A2(G952), .ZN(n1122) );
XNOR2_X1 U866 ( .A(G146), .B(n1192), .ZN(G48) );
NAND3_X1 U867 ( .A1(n1062), .A2(n1060), .A3(n1201), .ZN(n1192) );
XOR2_X1 U868 ( .A(n1204), .B(n1193), .Z(G45) );
NAND4_X1 U869 ( .A1(n1205), .A2(n1053), .A3(n1206), .A4(n1060), .ZN(n1193) );
NOR2_X1 U870 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U871 ( .A(n1198), .B(n1209), .Z(G42) );
XOR2_X1 U872 ( .A(KEYINPUT26), .B(G140), .Z(n1209) );
AND3_X1 U873 ( .A1(n1052), .A2(n1210), .A3(n1062), .ZN(n1198) );
XOR2_X1 U874 ( .A(G137), .B(n1197), .Z(G39) );
AND4_X1 U875 ( .A1(n1211), .A2(n1210), .A3(n1212), .A4(n1213), .ZN(n1197) );
XOR2_X1 U876 ( .A(G134), .B(n1196), .Z(G36) );
AND3_X1 U877 ( .A1(n1210), .A2(n1063), .A3(n1053), .ZN(n1196) );
XOR2_X1 U878 ( .A(G131), .B(n1093), .Z(G33) );
AND3_X1 U879 ( .A1(n1053), .A2(n1210), .A3(n1062), .ZN(n1093) );
AND4_X1 U880 ( .A1(n1035), .A2(n1060), .A3(n1214), .A4(n1055), .ZN(n1210) );
XOR2_X1 U881 ( .A(n1215), .B(n1216), .Z(G30) );
XOR2_X1 U882 ( .A(n1217), .B(KEYINPUT48), .Z(n1216) );
NAND3_X1 U883 ( .A1(n1201), .A2(n1063), .A3(n1218), .ZN(n1215) );
XNOR2_X1 U884 ( .A(n1060), .B(KEYINPUT46), .ZN(n1218) );
AND3_X1 U885 ( .A1(n1212), .A2(n1213), .A3(n1205), .ZN(n1201) );
XOR2_X1 U886 ( .A(n1189), .B(n1219), .Z(G3) );
NAND2_X1 U887 ( .A1(KEYINPUT22), .A2(G101), .ZN(n1219) );
NAND3_X1 U888 ( .A1(n1053), .A2(n1191), .A3(n1211), .ZN(n1189) );
XOR2_X1 U889 ( .A(n1220), .B(n1200), .Z(G27) );
NAND4_X1 U890 ( .A1(n1221), .A2(n1205), .A3(n1062), .A4(n1052), .ZN(n1200) );
AND2_X1 U891 ( .A1(n1042), .A2(n1214), .ZN(n1205) );
NAND2_X1 U892 ( .A1(n1222), .A2(n1050), .ZN(n1214) );
XOR2_X1 U893 ( .A(n1223), .B(KEYINPUT24), .Z(n1222) );
NAND4_X1 U894 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1097), .ZN(n1223) );
INV_X1 U895 ( .A(G900), .ZN(n1097) );
XNOR2_X1 U896 ( .A(n1183), .B(n1225), .ZN(G24) );
NOR2_X1 U897 ( .A1(KEYINPUT4), .A2(n1226), .ZN(n1225) );
NAND4_X1 U898 ( .A1(n1227), .A2(n1034), .A3(n1228), .A4(n1229), .ZN(n1183) );
NOR2_X1 U899 ( .A1(n1213), .A2(n1212), .ZN(n1034) );
XNOR2_X1 U900 ( .A(G119), .B(n1184), .ZN(G21) );
NAND4_X1 U901 ( .A1(n1227), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1184) );
XNOR2_X1 U902 ( .A(n1185), .B(n1230), .ZN(G18) );
XOR2_X1 U903 ( .A(KEYINPUT41), .B(G116), .Z(n1230) );
NAND3_X1 U904 ( .A1(n1053), .A2(n1063), .A3(n1227), .ZN(n1185) );
NOR2_X1 U905 ( .A1(n1229), .A2(n1208), .ZN(n1063) );
INV_X1 U906 ( .A(n1207), .ZN(n1229) );
XNOR2_X1 U907 ( .A(n1231), .B(n1186), .ZN(G15) );
NAND3_X1 U908 ( .A1(n1062), .A2(n1053), .A3(n1227), .ZN(n1186) );
AND3_X1 U909 ( .A1(n1042), .A2(n1232), .A3(n1221), .ZN(n1227) );
INV_X1 U910 ( .A(n1048), .ZN(n1221) );
NAND2_X1 U911 ( .A1(n1061), .A2(n1233), .ZN(n1048) );
NOR2_X1 U912 ( .A1(n1067), .A2(n1213), .ZN(n1053) );
NOR2_X1 U913 ( .A1(n1228), .A2(n1207), .ZN(n1062) );
INV_X1 U914 ( .A(n1208), .ZN(n1228) );
XOR2_X1 U915 ( .A(n1234), .B(KEYINPUT30), .Z(n1231) );
XNOR2_X1 U916 ( .A(G110), .B(n1190), .ZN(G12) );
NAND3_X1 U917 ( .A1(n1211), .A2(n1191), .A3(n1052), .ZN(n1190) );
AND2_X1 U918 ( .A1(n1067), .A2(n1213), .ZN(n1052) );
XNOR2_X1 U919 ( .A(n1078), .B(n1080), .ZN(n1213) );
NAND2_X1 U920 ( .A1(G217), .A2(n1235), .ZN(n1080) );
NOR2_X1 U921 ( .A1(n1125), .A2(G902), .ZN(n1078) );
XOR2_X1 U922 ( .A(n1236), .B(n1237), .Z(n1125) );
XNOR2_X1 U923 ( .A(n1101), .B(n1238), .ZN(n1237) );
XOR2_X1 U924 ( .A(n1239), .B(n1240), .Z(n1238) );
NAND2_X1 U925 ( .A1(n1241), .A2(G221), .ZN(n1239) );
XOR2_X1 U926 ( .A(n1220), .B(n1242), .Z(n1101) );
XOR2_X1 U927 ( .A(n1243), .B(n1244), .Z(n1236) );
XOR2_X1 U928 ( .A(G137), .B(G128), .Z(n1244) );
XNOR2_X1 U929 ( .A(G119), .B(G110), .ZN(n1243) );
INV_X1 U930 ( .A(n1212), .ZN(n1067) );
XOR2_X1 U931 ( .A(n1245), .B(n1246), .Z(n1212) );
XOR2_X1 U932 ( .A(KEYINPUT0), .B(G472), .Z(n1246) );
NAND2_X1 U933 ( .A1(n1247), .A2(n1248), .ZN(n1245) );
XOR2_X1 U934 ( .A(n1249), .B(n1250), .Z(n1247) );
XOR2_X1 U935 ( .A(n1148), .B(n1251), .Z(n1250) );
XOR2_X1 U936 ( .A(n1149), .B(n1156), .Z(n1251) );
NAND3_X1 U937 ( .A1(n1252), .A2(n1041), .A3(G210), .ZN(n1149) );
XOR2_X1 U938 ( .A(n1234), .B(n1253), .Z(n1148) );
XOR2_X1 U939 ( .A(n1157), .B(n1254), .Z(n1249) );
XOR2_X1 U940 ( .A(KEYINPUT21), .B(G101), .Z(n1254) );
INV_X1 U941 ( .A(n1140), .ZN(n1191) );
NAND3_X1 U942 ( .A1(n1042), .A2(n1232), .A3(n1060), .ZN(n1140) );
NOR2_X1 U943 ( .A1(n1061), .A2(n1064), .ZN(n1060) );
INV_X1 U944 ( .A(n1233), .ZN(n1064) );
NAND2_X1 U945 ( .A1(G221), .A2(n1235), .ZN(n1233) );
NAND2_X1 U946 ( .A1(n1255), .A2(n1248), .ZN(n1235) );
NAND3_X1 U947 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1061) );
NAND2_X1 U948 ( .A1(KEYINPUT29), .A2(n1075), .ZN(n1258) );
NAND3_X1 U949 ( .A1(n1259), .A2(n1260), .A3(n1077), .ZN(n1257) );
INV_X1 U950 ( .A(KEYINPUT29), .ZN(n1260) );
OR2_X1 U951 ( .A1(n1077), .A2(n1259), .ZN(n1256) );
NOR2_X1 U952 ( .A1(n1075), .A2(KEYINPUT25), .ZN(n1259) );
AND2_X1 U953 ( .A1(n1261), .A2(n1248), .ZN(n1075) );
XOR2_X1 U954 ( .A(n1262), .B(n1263), .Z(n1261) );
XOR2_X1 U955 ( .A(n1264), .B(n1173), .Z(n1263) );
XNOR2_X1 U956 ( .A(n1265), .B(n1266), .ZN(n1173) );
NOR2_X1 U957 ( .A1(G107), .A2(KEYINPUT33), .ZN(n1266) );
XOR2_X1 U958 ( .A(n1164), .B(n1156), .Z(n1264) );
XNOR2_X1 U959 ( .A(n1267), .B(n1100), .ZN(n1156) );
XOR2_X1 U960 ( .A(G134), .B(G137), .Z(n1100) );
XNOR2_X1 U961 ( .A(G131), .B(KEYINPUT38), .ZN(n1267) );
INV_X1 U962 ( .A(n1167), .ZN(n1164) );
XOR2_X1 U963 ( .A(G110), .B(G140), .Z(n1167) );
XNOR2_X1 U964 ( .A(n1268), .B(n1166), .ZN(n1262) );
NAND2_X1 U965 ( .A1(G227), .A2(n1041), .ZN(n1166) );
XOR2_X1 U966 ( .A(n1104), .B(KEYINPUT55), .Z(n1268) );
NAND2_X1 U967 ( .A1(n1269), .A2(n1270), .ZN(n1104) );
NAND3_X1 U968 ( .A1(KEYINPUT7), .A2(n1271), .A3(n1272), .ZN(n1270) );
XOR2_X1 U969 ( .A(n1217), .B(n1273), .Z(n1272) );
NOR2_X1 U970 ( .A1(G143), .A2(n1274), .ZN(n1273) );
NAND4_X1 U971 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1269) );
NAND2_X1 U972 ( .A1(G128), .A2(n1274), .ZN(n1278) );
INV_X1 U973 ( .A(KEYINPUT53), .ZN(n1274) );
NAND2_X1 U974 ( .A1(n1279), .A2(KEYINPUT53), .ZN(n1277) );
NAND2_X1 U975 ( .A1(KEYINPUT7), .A2(n1271), .ZN(n1275) );
XOR2_X1 U976 ( .A(KEYINPUT14), .B(n1240), .Z(n1271) );
INV_X1 U977 ( .A(G469), .ZN(n1077) );
NAND2_X1 U978 ( .A1(n1050), .A2(n1280), .ZN(n1232) );
NAND4_X1 U979 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1281), .ZN(n1280) );
INV_X1 U980 ( .A(G898), .ZN(n1281) );
NAND3_X1 U981 ( .A1(n1224), .A2(n1041), .A3(G952), .ZN(n1050) );
NAND2_X1 U982 ( .A1(G237), .A2(n1255), .ZN(n1224) );
XOR2_X1 U983 ( .A(G234), .B(KEYINPUT5), .Z(n1255) );
NOR2_X1 U984 ( .A1(n1035), .A2(n1037), .ZN(n1042) );
INV_X1 U985 ( .A(n1055), .ZN(n1037) );
NAND2_X1 U986 ( .A1(G214), .A2(n1282), .ZN(n1055) );
XOR2_X1 U987 ( .A(n1086), .B(n1084), .Z(n1035) );
NAND2_X1 U988 ( .A1(G210), .A2(n1282), .ZN(n1084) );
NAND2_X1 U989 ( .A1(n1252), .A2(n1248), .ZN(n1282) );
AND2_X1 U990 ( .A1(n1283), .A2(n1248), .ZN(n1086) );
XOR2_X1 U991 ( .A(n1284), .B(n1285), .Z(n1283) );
NOR2_X1 U992 ( .A1(KEYINPUT20), .A2(n1180), .ZN(n1285) );
XOR2_X1 U993 ( .A(n1119), .B(n1286), .Z(n1180) );
NOR2_X1 U994 ( .A1(KEYINPUT59), .A2(n1120), .ZN(n1286) );
XOR2_X1 U995 ( .A(n1287), .B(n1253), .Z(n1120) );
XOR2_X1 U996 ( .A(G116), .B(G119), .Z(n1253) );
NAND2_X1 U997 ( .A1(KEYINPUT42), .A2(n1234), .ZN(n1287) );
XNOR2_X1 U998 ( .A(n1288), .B(n1289), .ZN(n1119) );
XNOR2_X1 U999 ( .A(n1290), .B(n1265), .ZN(n1289) );
XNOR2_X1 U1000 ( .A(G104), .B(G101), .ZN(n1265) );
NOR2_X1 U1001 ( .A1(KEYINPUT34), .A2(n1024), .ZN(n1290) );
INV_X1 U1002 ( .A(G107), .ZN(n1024) );
XNOR2_X1 U1003 ( .A(G110), .B(n1291), .ZN(n1288) );
NOR2_X1 U1004 ( .A1(KEYINPUT12), .A2(n1226), .ZN(n1291) );
INV_X1 U1005 ( .A(G122), .ZN(n1226) );
NAND2_X1 U1006 ( .A1(n1292), .A2(n1293), .ZN(n1284) );
NAND2_X1 U1007 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XNOR2_X1 U1008 ( .A(n1157), .B(n1296), .ZN(n1294) );
XOR2_X1 U1009 ( .A(n1297), .B(KEYINPUT52), .Z(n1292) );
NAND2_X1 U1010 ( .A1(n1203), .A2(n1298), .ZN(n1297) );
XOR2_X1 U1011 ( .A(n1157), .B(n1296), .Z(n1298) );
NAND2_X1 U1012 ( .A1(KEYINPUT17), .A2(n1220), .ZN(n1296) );
INV_X1 U1013 ( .A(G125), .ZN(n1220) );
NAND3_X1 U1014 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1157) );
XOR2_X1 U1015 ( .A(n1302), .B(KEYINPUT37), .Z(n1301) );
NAND2_X1 U1016 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND3_X1 U1017 ( .A1(G143), .A2(G128), .A3(n1305), .ZN(n1304) );
OR2_X1 U1018 ( .A1(n1276), .A2(n1305), .ZN(n1303) );
NAND3_X1 U1019 ( .A1(n1217), .A2(n1204), .A3(n1305), .ZN(n1300) );
NAND2_X1 U1020 ( .A1(n1240), .A2(n1279), .ZN(n1299) );
INV_X1 U1021 ( .A(n1306), .ZN(n1279) );
INV_X1 U1022 ( .A(n1295), .ZN(n1203) );
NAND2_X1 U1023 ( .A1(G224), .A2(n1041), .ZN(n1295) );
INV_X1 U1024 ( .A(n1049), .ZN(n1211) );
NAND2_X1 U1025 ( .A1(n1208), .A2(n1207), .ZN(n1049) );
XOR2_X1 U1026 ( .A(n1307), .B(G475), .Z(n1207) );
NAND2_X1 U1027 ( .A1(KEYINPUT13), .A2(n1083), .ZN(n1307) );
NOR2_X1 U1028 ( .A1(n1134), .A2(G902), .ZN(n1083) );
XNOR2_X1 U1029 ( .A(n1308), .B(n1309), .ZN(n1134) );
XOR2_X1 U1030 ( .A(n1310), .B(n1311), .Z(n1309) );
XNOR2_X1 U1031 ( .A(n1312), .B(n1313), .ZN(n1311) );
NAND2_X1 U1032 ( .A1(n1314), .A2(KEYINPUT58), .ZN(n1313) );
XOR2_X1 U1033 ( .A(n1315), .B(G143), .Z(n1314) );
NAND3_X1 U1034 ( .A1(n1252), .A2(n1041), .A3(n1316), .ZN(n1315) );
XNOR2_X1 U1035 ( .A(G214), .B(KEYINPUT50), .ZN(n1316) );
INV_X1 U1036 ( .A(G237), .ZN(n1252) );
NAND2_X1 U1037 ( .A1(KEYINPUT44), .A2(n1317), .ZN(n1312) );
XOR2_X1 U1038 ( .A(KEYINPUT56), .B(n1240), .Z(n1317) );
INV_X1 U1039 ( .A(n1305), .ZN(n1240) );
XNOR2_X1 U1040 ( .A(G146), .B(KEYINPUT54), .ZN(n1305) );
XOR2_X1 U1041 ( .A(n1318), .B(G104), .Z(n1310) );
NAND2_X1 U1042 ( .A1(KEYINPUT39), .A2(n1242), .ZN(n1318) );
INV_X1 U1043 ( .A(G140), .ZN(n1242) );
XOR2_X1 U1044 ( .A(n1319), .B(n1320), .Z(n1308) );
XOR2_X1 U1045 ( .A(G131), .B(G125), .Z(n1320) );
XOR2_X1 U1046 ( .A(n1234), .B(G122), .Z(n1319) );
INV_X1 U1047 ( .A(G113), .ZN(n1234) );
XNOR2_X1 U1048 ( .A(n1074), .B(n1321), .ZN(n1208) );
NOR2_X1 U1049 ( .A1(KEYINPUT63), .A2(n1132), .ZN(n1321) );
INV_X1 U1050 ( .A(G478), .ZN(n1132) );
AND2_X1 U1051 ( .A1(n1130), .A2(n1248), .ZN(n1074) );
INV_X1 U1052 ( .A(G902), .ZN(n1248) );
XNOR2_X1 U1053 ( .A(n1322), .B(n1323), .ZN(n1130) );
AND2_X1 U1054 ( .A1(n1241), .A2(G217), .ZN(n1323) );
AND2_X1 U1055 ( .A1(G234), .A2(n1041), .ZN(n1241) );
INV_X1 U1056 ( .A(G953), .ZN(n1041) );
NAND2_X1 U1057 ( .A1(KEYINPUT40), .A2(n1324), .ZN(n1322) );
XOR2_X1 U1058 ( .A(n1325), .B(n1326), .Z(n1324) );
XOR2_X1 U1059 ( .A(n1327), .B(G107), .Z(n1326) );
NAND2_X1 U1060 ( .A1(KEYINPUT31), .A2(n1328), .ZN(n1327) );
XOR2_X1 U1061 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1062 ( .A(n1331), .B(KEYINPUT10), .Z(n1330) );
INV_X1 U1063 ( .A(G134), .ZN(n1331) );
NAND3_X1 U1064 ( .A1(n1332), .A2(n1333), .A3(n1306), .ZN(n1329) );
NAND2_X1 U1065 ( .A1(G143), .A2(n1217), .ZN(n1306) );
NAND2_X1 U1066 ( .A1(KEYINPUT9), .A2(n1217), .ZN(n1333) );
INV_X1 U1067 ( .A(G128), .ZN(n1217) );
OR2_X1 U1068 ( .A1(n1276), .A2(KEYINPUT9), .ZN(n1332) );
NAND2_X1 U1069 ( .A1(G128), .A2(n1204), .ZN(n1276) );
INV_X1 U1070 ( .A(G143), .ZN(n1204) );
XOR2_X1 U1071 ( .A(n1334), .B(G122), .Z(n1325) );
INV_X1 U1072 ( .A(G116), .ZN(n1334) );
endmodule


