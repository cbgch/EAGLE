//Key = 0011111100000010111111001110001101100001001110101000111001101010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;

XOR2_X1 U683 ( .A(G107), .B(n937), .Z(G9) );
NOR2_X1 U684 ( .A1(n938), .A2(n939), .ZN(G75) );
NOR4_X1 U685 ( .A1(n940), .A2(n941), .A3(n942), .A4(n943), .ZN(n939) );
INV_X1 U686 ( .A(G952), .ZN(n942) );
NAND4_X1 U687 ( .A1(n944), .A2(n945), .A3(n946), .A4(n947), .ZN(n940) );
NAND4_X1 U688 ( .A1(n948), .A2(n949), .A3(n950), .A4(n951), .ZN(n945) );
NAND2_X1 U689 ( .A1(KEYINPUT26), .A2(n952), .ZN(n950) );
NOR2_X1 U690 ( .A1(n953), .A2(n954), .ZN(n948) );
NOR2_X1 U691 ( .A1(n955), .A2(n956), .ZN(n954) );
NOR2_X1 U692 ( .A1(n957), .A2(n952), .ZN(n955) );
NOR2_X1 U693 ( .A1(n958), .A2(n959), .ZN(n957) );
NOR2_X1 U694 ( .A1(n960), .A2(n961), .ZN(n953) );
NOR2_X1 U695 ( .A1(n962), .A2(n963), .ZN(n960) );
NOR2_X1 U696 ( .A1(KEYINPUT26), .A2(n952), .ZN(n962) );
NAND4_X1 U697 ( .A1(n964), .A2(n965), .A3(n966), .A4(n967), .ZN(n944) );
NOR2_X1 U698 ( .A1(n963), .A2(n956), .ZN(n967) );
INV_X1 U699 ( .A(n952), .ZN(n966) );
NAND2_X1 U700 ( .A1(n968), .A2(n969), .ZN(n965) );
NAND3_X1 U701 ( .A1(n970), .A2(n971), .A3(n951), .ZN(n964) );
NAND2_X1 U702 ( .A1(n972), .A2(n973), .ZN(n971) );
NAND2_X1 U703 ( .A1(n974), .A2(n975), .ZN(n973) );
OR2_X1 U704 ( .A1(n976), .A2(n977), .ZN(n975) );
NAND2_X1 U705 ( .A1(n978), .A2(n979), .ZN(n970) );
OR2_X1 U706 ( .A1(n980), .A2(n981), .ZN(n979) );
NOR3_X1 U707 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n938) );
NOR2_X1 U708 ( .A1(KEYINPUT9), .A2(n985), .ZN(n984) );
NOR2_X1 U709 ( .A1(G953), .A2(G952), .ZN(n985) );
NOR2_X1 U710 ( .A1(n986), .A2(n987), .ZN(n983) );
INV_X1 U711 ( .A(KEYINPUT9), .ZN(n987) );
INV_X1 U712 ( .A(n946), .ZN(n982) );
NAND4_X1 U713 ( .A1(n988), .A2(n989), .A3(n990), .A4(n991), .ZN(n946) );
NOR3_X1 U714 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n991) );
XNOR2_X1 U715 ( .A(n968), .B(KEYINPUT62), .ZN(n994) );
NOR2_X1 U716 ( .A1(n995), .A2(n996), .ZN(n993) );
NAND3_X1 U717 ( .A1(n997), .A2(n976), .A3(n998), .ZN(n992) );
NOR3_X1 U718 ( .A1(n999), .A2(n1000), .A3(n1001), .ZN(n990) );
XNOR2_X1 U719 ( .A(n956), .B(KEYINPUT16), .ZN(n1001) );
XOR2_X1 U720 ( .A(n1002), .B(n1003), .Z(n1000) );
NOR2_X1 U721 ( .A1(G478), .A2(KEYINPUT40), .ZN(n1003) );
XOR2_X1 U722 ( .A(n1004), .B(KEYINPUT41), .Z(n988) );
NAND2_X1 U723 ( .A1(n995), .A2(n996), .ZN(n1004) );
XOR2_X1 U724 ( .A(n1005), .B(n1006), .Z(G72) );
XOR2_X1 U725 ( .A(n1007), .B(n1008), .Z(n1006) );
NOR2_X1 U726 ( .A1(n1009), .A2(n947), .ZN(n1008) );
AND2_X1 U727 ( .A1(G227), .A2(G900), .ZN(n1009) );
NAND2_X1 U728 ( .A1(n1010), .A2(n1011), .ZN(n1007) );
NAND2_X1 U729 ( .A1(G953), .A2(n1012), .ZN(n1011) );
XOR2_X1 U730 ( .A(n1013), .B(n1014), .Z(n1010) );
XOR2_X1 U731 ( .A(n1015), .B(n1016), .Z(n1014) );
XNOR2_X1 U732 ( .A(n1017), .B(n1018), .ZN(n1015) );
XNOR2_X1 U733 ( .A(G134), .B(n1019), .ZN(n1013) );
XOR2_X1 U734 ( .A(G140), .B(G137), .Z(n1019) );
NAND2_X1 U735 ( .A1(n947), .A2(n943), .ZN(n1005) );
XOR2_X1 U736 ( .A(n1020), .B(n1021), .Z(G69) );
NAND2_X1 U737 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U738 ( .A1(n941), .A2(n947), .ZN(n1023) );
NAND2_X1 U739 ( .A1(G953), .A2(n1024), .ZN(n1022) );
NAND2_X1 U740 ( .A1(n1025), .A2(G224), .ZN(n1024) );
XNOR2_X1 U741 ( .A(G898), .B(KEYINPUT48), .ZN(n1025) );
NAND2_X1 U742 ( .A1(KEYINPUT57), .A2(n1026), .ZN(n1020) );
NAND3_X1 U743 ( .A1(n1027), .A2(n1028), .A3(n1029), .ZN(n1026) );
XOR2_X1 U744 ( .A(KEYINPUT7), .B(n1030), .Z(n1029) );
NOR2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U746 ( .A1(n1031), .A2(n1032), .ZN(n1028) );
XOR2_X1 U747 ( .A(n1033), .B(n1034), .Z(n1032) );
NAND2_X1 U748 ( .A1(G953), .A2(n1035), .ZN(n1027) );
NOR2_X1 U749 ( .A1(n986), .A2(n1036), .ZN(G66) );
XOR2_X1 U750 ( .A(n1037), .B(n1038), .Z(n1036) );
NAND2_X1 U751 ( .A1(n1039), .A2(n1040), .ZN(n1037) );
NOR2_X1 U752 ( .A1(n986), .A2(n1041), .ZN(G63) );
XOR2_X1 U753 ( .A(n1042), .B(n1043), .Z(n1041) );
NAND2_X1 U754 ( .A1(n1039), .A2(G478), .ZN(n1042) );
NOR2_X1 U755 ( .A1(n986), .A2(n1044), .ZN(G60) );
XOR2_X1 U756 ( .A(n1045), .B(n1046), .Z(n1044) );
NAND2_X1 U757 ( .A1(n1039), .A2(G475), .ZN(n1045) );
XOR2_X1 U758 ( .A(G104), .B(n1047), .Z(G6) );
NOR2_X1 U759 ( .A1(n986), .A2(n1048), .ZN(G57) );
XOR2_X1 U760 ( .A(n1049), .B(n1050), .Z(n1048) );
XNOR2_X1 U761 ( .A(n1051), .B(n1052), .ZN(n1050) );
XOR2_X1 U762 ( .A(n1053), .B(n1054), .Z(n1049) );
NOR2_X1 U763 ( .A1(KEYINPUT47), .A2(n1055), .ZN(n1054) );
XOR2_X1 U764 ( .A(n1056), .B(n1057), .Z(n1053) );
NOR2_X1 U765 ( .A1(KEYINPUT35), .A2(n1058), .ZN(n1057) );
XOR2_X1 U766 ( .A(n1059), .B(n1060), .Z(n1058) );
NAND2_X1 U767 ( .A1(n1039), .A2(G472), .ZN(n1056) );
NOR2_X1 U768 ( .A1(n986), .A2(n1061), .ZN(G54) );
XOR2_X1 U769 ( .A(n1062), .B(n1063), .Z(n1061) );
XOR2_X1 U770 ( .A(n1064), .B(n1065), .Z(n1063) );
NAND2_X1 U771 ( .A1(n1039), .A2(G469), .ZN(n1064) );
INV_X1 U772 ( .A(n1066), .ZN(n1039) );
XNOR2_X1 U773 ( .A(KEYINPUT22), .B(n1067), .ZN(n1062) );
NOR2_X1 U774 ( .A1(KEYINPUT56), .A2(n1068), .ZN(n1067) );
NOR2_X1 U775 ( .A1(n986), .A2(n1069), .ZN(G51) );
XOR2_X1 U776 ( .A(n1070), .B(n1071), .Z(n1069) );
NOR2_X1 U777 ( .A1(n1066), .A2(n1072), .ZN(n1071) );
XOR2_X1 U778 ( .A(KEYINPUT54), .B(n1073), .Z(n1072) );
NAND2_X1 U779 ( .A1(G902), .A2(n1074), .ZN(n1066) );
OR2_X1 U780 ( .A1(n941), .A2(n943), .ZN(n1074) );
NAND4_X1 U781 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n943) );
NOR4_X1 U782 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1078) );
NOR2_X1 U783 ( .A1(n1083), .A2(n1084), .ZN(n1077) );
NOR3_X1 U784 ( .A1(n1085), .A2(n1086), .A3(n1087), .ZN(n1084) );
NAND4_X1 U785 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n941) );
NOR4_X1 U786 ( .A1(n1092), .A2(n1093), .A3(n937), .A4(n1094), .ZN(n1091) );
INV_X1 U787 ( .A(n1095), .ZN(n1094) );
AND3_X1 U788 ( .A1(n959), .A2(n972), .A3(n1096), .ZN(n937) );
NOR3_X1 U789 ( .A1(n1047), .A2(n1097), .A3(n1098), .ZN(n1090) );
NOR2_X1 U790 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
INV_X1 U791 ( .A(KEYINPUT46), .ZN(n1099) );
NOR4_X1 U792 ( .A1(KEYINPUT46), .A2(n1101), .A3(n969), .A4(n1102), .ZN(n1097) );
AND3_X1 U793 ( .A1(n1096), .A2(n972), .A3(n958), .ZN(n1047) );
NAND2_X1 U794 ( .A1(KEYINPUT3), .A2(n1103), .ZN(n1070) );
XOR2_X1 U795 ( .A(n1104), .B(n1105), .Z(n1103) );
NOR2_X1 U796 ( .A1(n1106), .A2(n1107), .ZN(n1105) );
XOR2_X1 U797 ( .A(KEYINPUT29), .B(n1108), .Z(n1107) );
AND2_X1 U798 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NOR2_X1 U799 ( .A1(n1109), .A2(n1110), .ZN(n1106) );
XNOR2_X1 U800 ( .A(n1111), .B(KEYINPUT53), .ZN(n1110) );
NOR2_X1 U801 ( .A1(KEYINPUT37), .A2(n1112), .ZN(n1104) );
XOR2_X1 U802 ( .A(n1113), .B(KEYINPUT31), .Z(n1112) );
NOR2_X1 U803 ( .A1(n947), .A2(G952), .ZN(n986) );
XOR2_X1 U804 ( .A(G146), .B(n1083), .Z(G48) );
AND4_X1 U805 ( .A1(n1114), .A2(n958), .A3(n1115), .A4(n1116), .ZN(n1083) );
XOR2_X1 U806 ( .A(n1076), .B(n1117), .Z(G45) );
NOR2_X1 U807 ( .A1(G143), .A2(KEYINPUT63), .ZN(n1117) );
NAND4_X1 U808 ( .A1(n1118), .A2(n980), .A3(n1115), .A4(n1119), .ZN(n1076) );
INV_X1 U809 ( .A(n1101), .ZN(n1118) );
NAND3_X1 U810 ( .A1(n999), .A2(n1120), .A3(n1121), .ZN(n1101) );
XOR2_X1 U811 ( .A(G140), .B(n1082), .Z(G42) );
AND3_X1 U812 ( .A1(n958), .A2(n981), .A3(n1122), .ZN(n1082) );
XOR2_X1 U813 ( .A(n1081), .B(n1123), .Z(G39) );
XOR2_X1 U814 ( .A(KEYINPUT49), .B(G137), .Z(n1123) );
AND2_X1 U815 ( .A1(n1122), .A2(n1124), .ZN(n1081) );
XNOR2_X1 U816 ( .A(n1125), .B(n1126), .ZN(G36) );
NOR4_X1 U817 ( .A1(n1127), .A2(n1086), .A3(n1087), .A4(n1085), .ZN(n1126) );
INV_X1 U818 ( .A(n980), .ZN(n1087) );
INV_X1 U819 ( .A(n959), .ZN(n1086) );
XNOR2_X1 U820 ( .A(KEYINPUT39), .B(KEYINPUT28), .ZN(n1127) );
XNOR2_X1 U821 ( .A(n1018), .B(n1080), .ZN(G33) );
AND3_X1 U822 ( .A1(n958), .A2(n980), .A3(n1122), .ZN(n1080) );
INV_X1 U823 ( .A(n1085), .ZN(n1122) );
NAND4_X1 U824 ( .A1(n961), .A2(n1115), .A3(n1119), .A4(n951), .ZN(n1085) );
INV_X1 U825 ( .A(n974), .ZN(n1115) );
XOR2_X1 U826 ( .A(G128), .B(n1128), .Z(G30) );
NOR2_X1 U827 ( .A1(KEYINPUT10), .A2(n1075), .ZN(n1128) );
NAND4_X1 U828 ( .A1(n1114), .A2(n959), .A3(n1129), .A4(n1116), .ZN(n1075) );
XOR2_X1 U829 ( .A(n1088), .B(n1130), .Z(G3) );
XOR2_X1 U830 ( .A(KEYINPUT2), .B(G101), .Z(n1130) );
NAND3_X1 U831 ( .A1(n980), .A2(n1096), .A3(n1131), .ZN(n1088) );
XOR2_X1 U832 ( .A(G125), .B(n1079), .Z(G27) );
AND4_X1 U833 ( .A1(n1114), .A2(n958), .A3(n978), .A4(n1132), .ZN(n1079) );
AND3_X1 U834 ( .A1(n1133), .A2(n1119), .A3(n1121), .ZN(n1114) );
NAND2_X1 U835 ( .A1(n952), .A2(n1134), .ZN(n1119) );
NAND4_X1 U836 ( .A1(G953), .A2(G902), .A3(n1135), .A4(n1012), .ZN(n1134) );
INV_X1 U837 ( .A(G900), .ZN(n1012) );
XNOR2_X1 U838 ( .A(G122), .B(n1100), .ZN(G24) );
NAND4_X1 U839 ( .A1(n949), .A2(n1136), .A3(n999), .A4(n1120), .ZN(n1100) );
INV_X1 U840 ( .A(n969), .ZN(n949) );
NAND2_X1 U841 ( .A1(n978), .A2(n972), .ZN(n969) );
NAND2_X1 U842 ( .A1(n1137), .A2(n1138), .ZN(n972) );
OR3_X1 U843 ( .A1(n1116), .A2(n1133), .A3(KEYINPUT11), .ZN(n1138) );
NAND2_X1 U844 ( .A1(KEYINPUT11), .A2(n981), .ZN(n1137) );
NAND2_X1 U845 ( .A1(n1139), .A2(n1140), .ZN(G21) );
NAND2_X1 U846 ( .A1(n1093), .A2(n1141), .ZN(n1140) );
XOR2_X1 U847 ( .A(KEYINPUT30), .B(n1142), .Z(n1139) );
NOR2_X1 U848 ( .A1(n1093), .A2(n1141), .ZN(n1142) );
AND3_X1 U849 ( .A1(n978), .A2(n1136), .A3(n1124), .ZN(n1093) );
NOR3_X1 U850 ( .A1(n989), .A2(n1132), .A3(n963), .ZN(n1124) );
INV_X1 U851 ( .A(n1131), .ZN(n963) );
XNOR2_X1 U852 ( .A(G116), .B(n1143), .ZN(G18) );
NAND2_X1 U853 ( .A1(KEYINPUT24), .A2(n1092), .ZN(n1143) );
AND4_X1 U854 ( .A1(n978), .A2(n980), .A3(n959), .A4(n1136), .ZN(n1092) );
NOR2_X1 U855 ( .A1(n999), .A2(n1144), .ZN(n959) );
XNOR2_X1 U856 ( .A(G113), .B(n1089), .ZN(G15) );
NAND4_X1 U857 ( .A1(n958), .A2(n978), .A3(n980), .A4(n1136), .ZN(n1089) );
NOR2_X1 U858 ( .A1(n1133), .A2(n1132), .ZN(n980) );
INV_X1 U859 ( .A(n1116), .ZN(n1132) );
NOR2_X1 U860 ( .A1(n977), .A2(n1145), .ZN(n978) );
INV_X1 U861 ( .A(n976), .ZN(n1145) );
AND2_X1 U862 ( .A1(n1144), .A2(n999), .ZN(n958) );
INV_X1 U863 ( .A(n1120), .ZN(n1144) );
XOR2_X1 U864 ( .A(n1146), .B(G110), .Z(G12) );
NAND2_X1 U865 ( .A1(KEYINPUT5), .A2(n1095), .ZN(n1146) );
NAND3_X1 U866 ( .A1(n1096), .A2(n981), .A3(n1131), .ZN(n1095) );
NOR2_X1 U867 ( .A1(n1120), .A2(n999), .ZN(n1131) );
XNOR2_X1 U868 ( .A(n1147), .B(G475), .ZN(n999) );
NAND2_X1 U869 ( .A1(n1046), .A2(n1148), .ZN(n1147) );
XOR2_X1 U870 ( .A(n1149), .B(n1150), .Z(n1046) );
XOR2_X1 U871 ( .A(n1151), .B(n1152), .Z(n1150) );
XNOR2_X1 U872 ( .A(G125), .B(n1153), .ZN(n1152) );
NOR2_X1 U873 ( .A1(KEYINPUT12), .A2(n1154), .ZN(n1153) );
XOR2_X1 U874 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U875 ( .A(n1157), .B(G104), .ZN(n1156) );
XOR2_X1 U876 ( .A(n1158), .B(G122), .Z(n1155) );
XNOR2_X1 U877 ( .A(KEYINPUT60), .B(KEYINPUT15), .ZN(n1158) );
NAND2_X1 U878 ( .A1(n1159), .A2(n1160), .ZN(n1151) );
NAND2_X1 U879 ( .A1(n1161), .A2(n1018), .ZN(n1160) );
XOR2_X1 U880 ( .A(KEYINPUT25), .B(n1162), .Z(n1159) );
NOR2_X1 U881 ( .A1(n1161), .A2(n1018), .ZN(n1162) );
INV_X1 U882 ( .A(G131), .ZN(n1018) );
XNOR2_X1 U883 ( .A(n1163), .B(n1164), .ZN(n1161) );
AND3_X1 U884 ( .A1(n1165), .A2(n1166), .A3(G214), .ZN(n1164) );
INV_X1 U885 ( .A(KEYINPUT23), .ZN(n1166) );
XNOR2_X1 U886 ( .A(G140), .B(n1167), .ZN(n1149) );
XOR2_X1 U887 ( .A(KEYINPUT44), .B(G146), .Z(n1167) );
NAND2_X1 U888 ( .A1(n1168), .A2(n1169), .ZN(n1120) );
OR2_X1 U889 ( .A1(n1002), .A2(G478), .ZN(n1169) );
XOR2_X1 U890 ( .A(n1170), .B(KEYINPUT27), .Z(n1168) );
NAND2_X1 U891 ( .A1(G478), .A2(n1002), .ZN(n1170) );
NAND2_X1 U892 ( .A1(n1171), .A2(n1043), .ZN(n1002) );
XNOR2_X1 U893 ( .A(n1172), .B(n1173), .ZN(n1043) );
XOR2_X1 U894 ( .A(n1174), .B(n1175), .Z(n1173) );
XNOR2_X1 U895 ( .A(n1125), .B(G128), .ZN(n1175) );
INV_X1 U896 ( .A(G134), .ZN(n1125) );
XNOR2_X1 U897 ( .A(KEYINPUT43), .B(n1163), .ZN(n1174) );
XOR2_X1 U898 ( .A(n1176), .B(n1177), .Z(n1172) );
XOR2_X1 U899 ( .A(G116), .B(G107), .Z(n1177) );
XOR2_X1 U900 ( .A(n1178), .B(n1179), .Z(n1176) );
NOR2_X1 U901 ( .A1(KEYINPUT51), .A2(G122), .ZN(n1179) );
NAND2_X1 U902 ( .A1(G217), .A2(n1180), .ZN(n1178) );
XNOR2_X1 U903 ( .A(G902), .B(KEYINPUT32), .ZN(n1171) );
NOR2_X1 U904 ( .A1(n1116), .A2(n989), .ZN(n981) );
INV_X1 U905 ( .A(n1133), .ZN(n989) );
XNOR2_X1 U906 ( .A(n1181), .B(n1040), .ZN(n1133) );
AND2_X1 U907 ( .A1(G217), .A2(n1182), .ZN(n1040) );
NAND2_X1 U908 ( .A1(n1038), .A2(n1148), .ZN(n1181) );
XNOR2_X1 U909 ( .A(n1183), .B(n1184), .ZN(n1038) );
XNOR2_X1 U910 ( .A(G119), .B(n1185), .ZN(n1184) );
NAND2_X1 U911 ( .A1(n1186), .A2(KEYINPUT58), .ZN(n1185) );
XOR2_X1 U912 ( .A(n1187), .B(G137), .Z(n1186) );
NAND2_X1 U913 ( .A1(n1180), .A2(G221), .ZN(n1187) );
AND2_X1 U914 ( .A1(G234), .A2(n947), .ZN(n1180) );
XOR2_X1 U915 ( .A(n1017), .B(n1188), .Z(n1183) );
NAND2_X1 U916 ( .A1(n1189), .A2(n998), .ZN(n1116) );
NAND3_X1 U917 ( .A1(n1190), .A2(n1148), .A3(n1191), .ZN(n998) );
XNOR2_X1 U918 ( .A(G472), .B(KEYINPUT59), .ZN(n1191) );
XNOR2_X1 U919 ( .A(KEYINPUT6), .B(n997), .ZN(n1189) );
NAND2_X1 U920 ( .A1(n1192), .A2(n1193), .ZN(n997) );
NAND2_X1 U921 ( .A1(n1190), .A2(n1148), .ZN(n1193) );
XNOR2_X1 U922 ( .A(n1194), .B(n1195), .ZN(n1190) );
XOR2_X1 U923 ( .A(n1196), .B(n1197), .Z(n1195) );
XNOR2_X1 U924 ( .A(KEYINPUT14), .B(n1059), .ZN(n1197) );
XNOR2_X1 U925 ( .A(n1055), .B(n1198), .ZN(n1194) );
INV_X1 U926 ( .A(n1051), .ZN(n1198) );
XNOR2_X1 U927 ( .A(n1199), .B(G101), .ZN(n1051) );
NAND2_X1 U928 ( .A1(n1165), .A2(G210), .ZN(n1199) );
NOR2_X1 U929 ( .A1(G953), .A2(G237), .ZN(n1165) );
XNOR2_X1 U930 ( .A(G113), .B(n1200), .ZN(n1055) );
XOR2_X1 U931 ( .A(KEYINPUT59), .B(G472), .Z(n1192) );
AND2_X1 U932 ( .A1(n1136), .A2(n1129), .ZN(n1096) );
XNOR2_X1 U933 ( .A(KEYINPUT36), .B(n974), .ZN(n1129) );
NAND2_X1 U934 ( .A1(n977), .A2(n976), .ZN(n974) );
NAND2_X1 U935 ( .A1(G221), .A2(n1182), .ZN(n976) );
NAND2_X1 U936 ( .A1(G234), .A2(n1201), .ZN(n1182) );
XNOR2_X1 U937 ( .A(KEYINPUT19), .B(n1148), .ZN(n1201) );
XNOR2_X1 U938 ( .A(n995), .B(n996), .ZN(n977) );
INV_X1 U939 ( .A(G469), .ZN(n996) );
AND2_X1 U940 ( .A1(n1202), .A2(n1148), .ZN(n995) );
XOR2_X1 U941 ( .A(n1065), .B(n1203), .Z(n1202) );
XNOR2_X1 U942 ( .A(KEYINPUT42), .B(n1068), .ZN(n1203) );
NAND2_X1 U943 ( .A1(G227), .A2(n947), .ZN(n1068) );
XOR2_X1 U944 ( .A(n1204), .B(n1205), .Z(n1065) );
XOR2_X1 U945 ( .A(n1206), .B(n1207), .Z(n1205) );
XOR2_X1 U946 ( .A(KEYINPUT55), .B(G101), .Z(n1207) );
NOR2_X1 U947 ( .A1(KEYINPUT45), .A2(n1208), .ZN(n1206) );
XOR2_X1 U948 ( .A(KEYINPUT4), .B(n1209), .Z(n1208) );
XNOR2_X1 U949 ( .A(n1016), .B(n1210), .ZN(n1204) );
XOR2_X1 U950 ( .A(n1188), .B(n1196), .Z(n1210) );
XOR2_X1 U951 ( .A(n1060), .B(n1052), .Z(n1196) );
XNOR2_X1 U952 ( .A(n1211), .B(n1212), .ZN(n1052) );
XOR2_X1 U953 ( .A(n1213), .B(n1214), .Z(n1212) );
NOR2_X1 U954 ( .A1(G134), .A2(KEYINPUT1), .ZN(n1214) );
NOR2_X1 U955 ( .A1(G131), .A2(n1215), .ZN(n1213) );
XNOR2_X1 U956 ( .A(KEYINPUT18), .B(KEYINPUT13), .ZN(n1215) );
XNOR2_X1 U957 ( .A(G137), .B(KEYINPUT38), .ZN(n1211) );
XOR2_X1 U958 ( .A(G140), .B(n1216), .Z(n1188) );
XOR2_X1 U959 ( .A(G143), .B(KEYINPUT34), .Z(n1016) );
AND2_X1 U960 ( .A1(n1121), .A2(n1102), .ZN(n1136) );
NAND2_X1 U961 ( .A1(n952), .A2(n1217), .ZN(n1102) );
NAND4_X1 U962 ( .A1(G953), .A2(G902), .A3(n1135), .A4(n1035), .ZN(n1217) );
INV_X1 U963 ( .A(G898), .ZN(n1035) );
NAND3_X1 U964 ( .A1(n1135), .A2(n947), .A3(G952), .ZN(n952) );
NAND2_X1 U965 ( .A1(G237), .A2(G234), .ZN(n1135) );
NOR2_X1 U966 ( .A1(n961), .A2(n968), .ZN(n1121) );
INV_X1 U967 ( .A(n951), .ZN(n968) );
NAND2_X1 U968 ( .A1(G214), .A2(n1218), .ZN(n951) );
INV_X1 U969 ( .A(n956), .ZN(n961) );
XNOR2_X1 U970 ( .A(n1219), .B(n1073), .ZN(n956) );
AND2_X1 U971 ( .A1(G210), .A2(n1218), .ZN(n1073) );
NAND2_X1 U972 ( .A1(n1220), .A2(n1148), .ZN(n1218) );
INV_X1 U973 ( .A(G237), .ZN(n1220) );
NAND2_X1 U974 ( .A1(n1221), .A2(n1148), .ZN(n1219) );
INV_X1 U975 ( .A(G902), .ZN(n1148) );
XOR2_X1 U976 ( .A(n1113), .B(n1222), .Z(n1221) );
XNOR2_X1 U977 ( .A(n1223), .B(n1109), .ZN(n1222) );
NAND2_X1 U978 ( .A1(G224), .A2(n947), .ZN(n1109) );
INV_X1 U979 ( .A(G953), .ZN(n947) );
NAND2_X1 U980 ( .A1(KEYINPUT52), .A2(n1111), .ZN(n1223) );
XNOR2_X1 U981 ( .A(n1017), .B(n1059), .ZN(n1111) );
NAND2_X1 U982 ( .A1(KEYINPUT21), .A2(n1163), .ZN(n1059) );
INV_X1 U983 ( .A(G143), .ZN(n1163) );
XNOR2_X1 U984 ( .A(G125), .B(n1060), .ZN(n1017) );
XOR2_X1 U985 ( .A(G128), .B(G146), .Z(n1060) );
XOR2_X1 U986 ( .A(n1033), .B(n1224), .Z(n1113) );
XNOR2_X1 U987 ( .A(n1225), .B(n1031), .ZN(n1224) );
XNOR2_X1 U988 ( .A(G122), .B(n1226), .ZN(n1031) );
NOR2_X1 U989 ( .A1(KEYINPUT0), .A2(n1227), .ZN(n1226) );
XNOR2_X1 U990 ( .A(n1216), .B(KEYINPUT20), .ZN(n1227) );
XOR2_X1 U991 ( .A(G110), .B(KEYINPUT17), .Z(n1216) );
NOR2_X1 U992 ( .A1(KEYINPUT8), .A2(n1034), .ZN(n1225) );
XOR2_X1 U993 ( .A(n1228), .B(n1200), .Z(n1034) );
XNOR2_X1 U994 ( .A(G116), .B(n1141), .ZN(n1200) );
INV_X1 U995 ( .A(G119), .ZN(n1141) );
NAND2_X1 U996 ( .A1(KEYINPUT33), .A2(n1157), .ZN(n1228) );
INV_X1 U997 ( .A(G113), .ZN(n1157) );
XNOR2_X1 U998 ( .A(n1209), .B(n1229), .ZN(n1033) );
NOR2_X1 U999 ( .A1(KEYINPUT50), .A2(n1230), .ZN(n1229) );
XOR2_X1 U1000 ( .A(KEYINPUT61), .B(G101), .Z(n1230) );
XOR2_X1 U1001 ( .A(G104), .B(G107), .Z(n1209) );
endmodule


