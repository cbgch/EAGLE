//Key = 1101111110100111110001101001100011011011001010111101010100001011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
n1358, n1359, n1360, n1361;

XOR2_X1 U748 ( .A(n1038), .B(n1039), .Z(G9) );
NAND4_X1 U749 ( .A1(n1040), .A2(KEYINPUT0), .A3(n1041), .A4(n1042), .ZN(n1039) );
XOR2_X1 U750 ( .A(n1043), .B(KEYINPUT7), .Z(n1040) );
NOR2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(G75) );
NOR4_X1 U752 ( .A1(G953), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1045) );
NOR3_X1 U753 ( .A1(n1049), .A2(KEYINPUT54), .A3(n1050), .ZN(n1047) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR4_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052) );
NOR2_X1 U756 ( .A1(n1057), .A2(n1058), .ZN(n1053) );
XNOR2_X1 U757 ( .A(n1059), .B(KEYINPUT38), .ZN(n1058) );
NOR3_X1 U758 ( .A1(n1060), .A2(n1061), .A3(n1062), .ZN(n1051) );
NOR2_X1 U759 ( .A1(n1063), .A2(n1064), .ZN(n1061) );
NOR2_X1 U760 ( .A1(n1065), .A2(n1056), .ZN(n1064) );
NOR3_X1 U761 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1065) );
NOR3_X1 U762 ( .A1(n1069), .A2(KEYINPUT36), .A3(n1070), .ZN(n1068) );
NOR3_X1 U763 ( .A1(n1071), .A2(n1072), .A3(n1054), .ZN(n1066) );
NOR2_X1 U764 ( .A1(n1070), .A2(n1055), .ZN(n1063) );
AND3_X1 U765 ( .A1(n1073), .A2(n1074), .A3(n1075), .ZN(n1070) );
INV_X1 U766 ( .A(n1055), .ZN(n1075) );
NAND2_X1 U767 ( .A1(n1076), .A2(n1077), .ZN(n1074) );
NAND2_X1 U768 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U769 ( .A1(n1080), .A2(n1081), .ZN(n1079) );
XOR2_X1 U770 ( .A(n1082), .B(n1083), .Z(n1081) );
NAND2_X1 U771 ( .A1(KEYINPUT36), .A2(n1084), .ZN(n1078) );
NAND2_X1 U772 ( .A1(n1085), .A2(n1086), .ZN(n1073) );
NAND2_X1 U773 ( .A1(n1087), .A2(n1088), .ZN(n1086) );
NOR3_X1 U774 ( .A1(n1046), .A2(G953), .A3(G952), .ZN(n1044) );
AND4_X1 U775 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1046) );
NOR3_X1 U776 ( .A1(n1093), .A2(n1060), .A3(n1094), .ZN(n1092) );
XOR2_X1 U777 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND3_X1 U778 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1093) );
XOR2_X1 U779 ( .A(n1100), .B(KEYINPUT40), .Z(n1099) );
NAND2_X1 U780 ( .A1(KEYINPUT20), .A2(n1101), .ZN(n1098) );
NAND3_X1 U781 ( .A1(n1102), .A2(n1103), .A3(G478), .ZN(n1097) );
INV_X1 U782 ( .A(KEYINPUT20), .ZN(n1103) );
NOR3_X1 U783 ( .A1(n1104), .A2(n1105), .A3(n1080), .ZN(n1091) );
INV_X1 U784 ( .A(n1071), .ZN(n1105) );
NOR3_X1 U785 ( .A1(n1106), .A2(KEYINPUT58), .A3(n1107), .ZN(n1104) );
NAND2_X1 U786 ( .A1(n1108), .A2(n1109), .ZN(n1090) );
NAND2_X1 U787 ( .A1(n1110), .A2(n1111), .ZN(n1108) );
NAND2_X1 U788 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
OR2_X1 U789 ( .A1(n1106), .A2(KEYINPUT58), .ZN(n1113) );
NAND2_X1 U790 ( .A1(n1114), .A2(n1101), .ZN(n1110) );
INV_X1 U791 ( .A(G478), .ZN(n1101) );
XNOR2_X1 U792 ( .A(G469), .B(n1115), .ZN(n1089) );
NAND2_X1 U793 ( .A1(KEYINPUT21), .A2(n1116), .ZN(n1115) );
XOR2_X1 U794 ( .A(n1117), .B(n1118), .Z(G72) );
NOR2_X1 U795 ( .A1(n1119), .A2(G953), .ZN(n1118) );
NAND2_X1 U796 ( .A1(n1120), .A2(n1121), .ZN(n1117) );
NAND2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
INV_X1 U798 ( .A(n1124), .ZN(n1122) );
NAND2_X1 U799 ( .A1(n1125), .A2(n1124), .ZN(n1120) );
NAND2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1124) );
XNOR2_X1 U801 ( .A(n1128), .B(n1129), .ZN(n1126) );
NOR2_X1 U802 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U803 ( .A(n1132), .B(KEYINPUT14), .Z(n1131) );
NAND2_X1 U804 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U805 ( .A1(n1133), .A2(n1134), .ZN(n1130) );
XOR2_X1 U806 ( .A(G137), .B(n1135), .Z(n1134) );
NAND2_X1 U807 ( .A1(n1127), .A2(n1123), .ZN(n1125) );
NAND2_X1 U808 ( .A1(G953), .A2(n1136), .ZN(n1123) );
INV_X1 U809 ( .A(n1137), .ZN(n1127) );
NAND3_X1 U810 ( .A1(n1138), .A2(n1139), .A3(n1140), .ZN(G69) );
NAND2_X1 U811 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
OR3_X1 U812 ( .A1(n1142), .A2(n1141), .A3(n1143), .ZN(n1139) );
INV_X1 U813 ( .A(KEYINPUT6), .ZN(n1142) );
NAND2_X1 U814 ( .A1(n1143), .A2(n1144), .ZN(n1138) );
NAND2_X1 U815 ( .A1(KEYINPUT6), .A2(n1145), .ZN(n1144) );
XNOR2_X1 U816 ( .A(KEYINPUT29), .B(n1141), .ZN(n1145) );
NAND2_X1 U817 ( .A1(G953), .A2(n1146), .ZN(n1141) );
NAND2_X1 U818 ( .A1(G898), .A2(G224), .ZN(n1146) );
NAND2_X1 U819 ( .A1(n1147), .A2(n1148), .ZN(n1143) );
NAND2_X1 U820 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
XNOR2_X1 U821 ( .A(n1151), .B(n1152), .ZN(n1149) );
NOR3_X1 U822 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
XOR2_X1 U823 ( .A(KEYINPUT43), .B(n1156), .Z(n1153) );
NAND3_X1 U824 ( .A1(G898), .A2(n1151), .A3(G953), .ZN(n1147) );
XNOR2_X1 U825 ( .A(n1157), .B(KEYINPUT19), .ZN(n1151) );
NOR2_X1 U826 ( .A1(n1158), .A2(n1159), .ZN(G66) );
XOR2_X1 U827 ( .A(n1160), .B(n1161), .Z(n1159) );
NAND2_X1 U828 ( .A1(KEYINPUT39), .A2(n1162), .ZN(n1161) );
NAND2_X1 U829 ( .A1(n1163), .A2(G217), .ZN(n1160) );
NOR2_X1 U830 ( .A1(n1158), .A2(n1164), .ZN(G63) );
XOR2_X1 U831 ( .A(n1114), .B(n1165), .Z(n1164) );
NAND2_X1 U832 ( .A1(n1163), .A2(G478), .ZN(n1165) );
NOR2_X1 U833 ( .A1(n1158), .A2(n1166), .ZN(G60) );
XNOR2_X1 U834 ( .A(n1167), .B(n1168), .ZN(n1166) );
XOR2_X1 U835 ( .A(n1169), .B(KEYINPUT3), .Z(n1168) );
NAND2_X1 U836 ( .A1(n1163), .A2(G475), .ZN(n1169) );
XOR2_X1 U837 ( .A(G104), .B(n1170), .Z(G6) );
NOR3_X1 U838 ( .A1(n1087), .A2(n1043), .A3(n1171), .ZN(n1170) );
NOR2_X1 U839 ( .A1(n1158), .A2(n1172), .ZN(G57) );
XOR2_X1 U840 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U841 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U842 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
NAND2_X1 U843 ( .A1(n1179), .A2(G101), .ZN(n1178) );
NAND2_X1 U844 ( .A1(n1180), .A2(n1181), .ZN(n1177) );
XNOR2_X1 U845 ( .A(n1179), .B(KEYINPUT59), .ZN(n1180) );
XOR2_X1 U846 ( .A(n1182), .B(n1183), .Z(n1173) );
NOR2_X1 U847 ( .A1(KEYINPUT37), .A2(n1184), .ZN(n1183) );
NAND2_X1 U848 ( .A1(n1163), .A2(G472), .ZN(n1182) );
NOR2_X1 U849 ( .A1(n1158), .A2(n1185), .ZN(G54) );
XOR2_X1 U850 ( .A(n1186), .B(n1187), .Z(n1185) );
NAND2_X1 U851 ( .A1(n1163), .A2(G469), .ZN(n1187) );
NAND2_X1 U852 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
NAND2_X1 U853 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
XOR2_X1 U854 ( .A(KEYINPUT33), .B(n1192), .Z(n1188) );
NOR2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1192) );
XOR2_X1 U856 ( .A(n1193), .B(n1194), .Z(n1191) );
XOR2_X1 U857 ( .A(n1195), .B(KEYINPUT60), .Z(n1193) );
XOR2_X1 U858 ( .A(n1196), .B(n1197), .Z(n1190) );
XOR2_X1 U859 ( .A(G110), .B(n1198), .Z(n1197) );
XOR2_X1 U860 ( .A(n1199), .B(KEYINPUT9), .Z(n1196) );
INV_X1 U861 ( .A(G140), .ZN(n1199) );
NOR2_X1 U862 ( .A1(n1158), .A2(n1200), .ZN(G51) );
XOR2_X1 U863 ( .A(n1157), .B(n1201), .Z(n1200) );
XOR2_X1 U864 ( .A(n1202), .B(n1203), .Z(n1201) );
NAND2_X1 U865 ( .A1(KEYINPUT15), .A2(n1204), .ZN(n1203) );
NAND2_X1 U866 ( .A1(n1163), .A2(n1205), .ZN(n1202) );
AND2_X1 U867 ( .A1(G902), .A2(n1048), .ZN(n1163) );
NAND3_X1 U868 ( .A1(n1206), .A2(n1207), .A3(n1119), .ZN(n1048) );
AND4_X1 U869 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1119) );
NOR4_X1 U870 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1211) );
NOR2_X1 U871 ( .A1(n1216), .A2(n1217), .ZN(n1210) );
INV_X1 U872 ( .A(n1218), .ZN(n1217) );
XOR2_X1 U873 ( .A(KEYINPUT30), .B(n1219), .Z(n1207) );
NOR2_X1 U874 ( .A1(n1156), .A2(n1154), .ZN(n1219) );
NAND3_X1 U875 ( .A1(n1220), .A2(n1221), .A3(n1222), .ZN(n1154) );
NAND3_X1 U876 ( .A1(n1223), .A2(n1042), .A3(n1224), .ZN(n1222) );
XOR2_X1 U877 ( .A(n1043), .B(KEYINPUT8), .Z(n1224) );
INV_X1 U878 ( .A(n1171), .ZN(n1042) );
NOR3_X1 U879 ( .A1(n1171), .A2(n1043), .A3(n1088), .ZN(n1156) );
NAND4_X1 U880 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1171) );
INV_X1 U881 ( .A(n1155), .ZN(n1206) );
NAND4_X1 U882 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1155) );
NAND4_X1 U883 ( .A1(n1233), .A2(n1067), .A3(n1057), .A4(n1223), .ZN(n1230) );
XOR2_X1 U884 ( .A(n1228), .B(KEYINPUT31), .Z(n1233) );
NAND2_X1 U885 ( .A1(n1234), .A2(n1235), .ZN(n1229) );
NOR2_X1 U886 ( .A1(n1150), .A2(G952), .ZN(n1158) );
XNOR2_X1 U887 ( .A(G146), .B(n1209), .ZN(G48) );
NAND3_X1 U888 ( .A1(n1084), .A2(n1223), .A3(n1236), .ZN(n1209) );
XOR2_X1 U889 ( .A(n1237), .B(n1218), .Z(G45) );
NAND4_X1 U890 ( .A1(n1084), .A2(n1238), .A3(n1057), .A4(n1239), .ZN(n1218) );
NOR3_X1 U891 ( .A1(n1100), .A2(n1240), .A3(n1241), .ZN(n1239) );
XOR2_X1 U892 ( .A(G140), .B(n1215), .Z(G42) );
AND3_X1 U893 ( .A1(n1242), .A2(n1223), .A3(n1059), .ZN(n1215) );
XOR2_X1 U894 ( .A(G137), .B(n1214), .Z(G39) );
AND2_X1 U895 ( .A1(n1235), .A2(n1242), .ZN(n1214) );
XOR2_X1 U896 ( .A(n1243), .B(n1213), .Z(G36) );
AND3_X1 U897 ( .A1(n1242), .A2(n1041), .A3(n1057), .ZN(n1213) );
XNOR2_X1 U898 ( .A(G134), .B(KEYINPUT51), .ZN(n1243) );
XOR2_X1 U899 ( .A(G131), .B(n1212), .Z(G33) );
AND3_X1 U900 ( .A1(n1242), .A2(n1223), .A3(n1057), .ZN(n1212) );
NOR3_X1 U901 ( .A1(n1069), .A2(n1240), .A3(n1055), .ZN(n1242) );
NAND2_X1 U902 ( .A1(n1071), .A2(n1244), .ZN(n1055) );
INV_X1 U903 ( .A(n1084), .ZN(n1069) );
XNOR2_X1 U904 ( .A(n1225), .B(KEYINPUT62), .ZN(n1084) );
XNOR2_X1 U905 ( .A(G128), .B(n1245), .ZN(G30) );
NAND2_X1 U906 ( .A1(n1246), .A2(n1216), .ZN(n1245) );
AND3_X1 U907 ( .A1(n1041), .A2(n1225), .A3(n1236), .ZN(n1216) );
NOR4_X1 U908 ( .A1(n1227), .A2(n1043), .A3(n1240), .A4(n1226), .ZN(n1236) );
INV_X1 U909 ( .A(n1247), .ZN(n1240) );
INV_X1 U910 ( .A(n1088), .ZN(n1041) );
XNOR2_X1 U911 ( .A(KEYINPUT56), .B(KEYINPUT34), .ZN(n1246) );
XOR2_X1 U912 ( .A(n1181), .B(n1220), .Z(G3) );
NAND2_X1 U913 ( .A1(n1248), .A2(n1057), .ZN(n1220) );
INV_X1 U914 ( .A(G101), .ZN(n1181) );
NAND3_X1 U915 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(G27) );
NAND2_X1 U916 ( .A1(n1208), .A2(n1252), .ZN(n1251) );
OR3_X1 U917 ( .A1(n1252), .A2(n1208), .A3(G125), .ZN(n1250) );
INV_X1 U918 ( .A(KEYINPUT49), .ZN(n1252) );
NAND2_X1 U919 ( .A1(G125), .A2(n1253), .ZN(n1249) );
NAND2_X1 U920 ( .A1(KEYINPUT49), .A2(n1254), .ZN(n1253) );
XNOR2_X1 U921 ( .A(KEYINPUT57), .B(n1208), .ZN(n1254) );
NAND4_X1 U922 ( .A1(n1067), .A2(n1059), .A3(n1223), .A4(n1247), .ZN(n1208) );
NAND2_X1 U923 ( .A1(n1255), .A2(n1256), .ZN(n1247) );
NAND3_X1 U924 ( .A1(G902), .A2(n1257), .A3(n1137), .ZN(n1256) );
NOR2_X1 U925 ( .A1(G900), .A2(n1150), .ZN(n1137) );
INV_X1 U926 ( .A(n1087), .ZN(n1223) );
XOR2_X1 U927 ( .A(n1231), .B(n1258), .Z(G24) );
NAND2_X1 U928 ( .A1(KEYINPUT63), .A2(G122), .ZN(n1258) );
NAND3_X1 U929 ( .A1(n1234), .A2(n1226), .A3(n1259), .ZN(n1231) );
NOR3_X1 U930 ( .A1(n1062), .A2(n1241), .A3(n1100), .ZN(n1259) );
XNOR2_X1 U931 ( .A(G119), .B(n1260), .ZN(G21) );
NAND3_X1 U932 ( .A1(n1234), .A2(n1235), .A3(KEYINPUT10), .ZN(n1260) );
NOR3_X1 U933 ( .A1(n1227), .A2(n1226), .A3(n1056), .ZN(n1235) );
XNOR2_X1 U934 ( .A(G116), .B(n1232), .ZN(G18) );
OR2_X1 U935 ( .A1(n1261), .A2(n1088), .ZN(n1232) );
NAND2_X1 U936 ( .A1(n1100), .A2(n1262), .ZN(n1088) );
INV_X1 U937 ( .A(n1241), .ZN(n1262) );
XOR2_X1 U938 ( .A(G113), .B(n1263), .Z(G15) );
NOR2_X1 U939 ( .A1(n1087), .A2(n1261), .ZN(n1263) );
NAND2_X1 U940 ( .A1(n1234), .A2(n1057), .ZN(n1261) );
NOR2_X1 U941 ( .A1(n1227), .A2(n1060), .ZN(n1057) );
INV_X1 U942 ( .A(n1062), .ZN(n1227) );
AND2_X1 U943 ( .A1(n1067), .A2(n1228), .ZN(n1234) );
NOR2_X1 U944 ( .A1(n1043), .A2(n1054), .ZN(n1067) );
INV_X1 U945 ( .A(n1085), .ZN(n1054) );
NAND2_X1 U946 ( .A1(n1264), .A2(n1265), .ZN(n1085) );
NAND2_X1 U947 ( .A1(n1225), .A2(n1082), .ZN(n1265) );
INV_X1 U948 ( .A(KEYINPUT22), .ZN(n1082) );
NAND3_X1 U949 ( .A1(n1083), .A2(n1266), .A3(KEYINPUT22), .ZN(n1264) );
NAND2_X1 U950 ( .A1(n1241), .A2(n1267), .ZN(n1087) );
INV_X1 U951 ( .A(n1100), .ZN(n1267) );
XOR2_X1 U952 ( .A(n1268), .B(n1221), .Z(G12) );
NAND2_X1 U953 ( .A1(n1248), .A2(n1059), .ZN(n1221) );
NOR2_X1 U954 ( .A1(n1062), .A2(n1226), .ZN(n1059) );
INV_X1 U955 ( .A(n1060), .ZN(n1226) );
NAND3_X1 U956 ( .A1(n1269), .A2(n1270), .A3(n1271), .ZN(n1060) );
NAND2_X1 U957 ( .A1(G902), .A2(G217), .ZN(n1271) );
OR3_X1 U958 ( .A1(n1162), .A2(G902), .A3(n1272), .ZN(n1270) );
NAND2_X1 U959 ( .A1(n1272), .A2(n1162), .ZN(n1269) );
XNOR2_X1 U960 ( .A(n1273), .B(n1274), .ZN(n1162) );
XOR2_X1 U961 ( .A(n1275), .B(n1276), .Z(n1274) );
XOR2_X1 U962 ( .A(G110), .B(n1277), .Z(n1276) );
NOR2_X1 U963 ( .A1(G146), .A2(n1278), .ZN(n1277) );
XNOR2_X1 U964 ( .A(KEYINPUT52), .B(KEYINPUT46), .ZN(n1278) );
XOR2_X1 U965 ( .A(G137), .B(G119), .Z(n1275) );
XNOR2_X1 U966 ( .A(n1128), .B(n1279), .ZN(n1273) );
XOR2_X1 U967 ( .A(n1280), .B(n1281), .Z(n1279) );
NAND2_X1 U968 ( .A1(KEYINPUT4), .A2(G128), .ZN(n1281) );
NAND3_X1 U969 ( .A1(n1282), .A2(n1150), .A3(G221), .ZN(n1280) );
NOR2_X1 U970 ( .A1(n1283), .A2(G234), .ZN(n1272) );
INV_X1 U971 ( .A(G217), .ZN(n1283) );
XNOR2_X1 U972 ( .A(n1284), .B(n1096), .ZN(n1062) );
NAND2_X1 U973 ( .A1(n1285), .A2(n1109), .ZN(n1096) );
XOR2_X1 U974 ( .A(n1286), .B(n1287), .Z(n1285) );
XOR2_X1 U975 ( .A(G101), .B(n1179), .Z(n1287) );
AND3_X1 U976 ( .A1(n1288), .A2(n1150), .A3(G210), .ZN(n1179) );
XNOR2_X1 U977 ( .A(n1289), .B(n1184), .ZN(n1286) );
XOR2_X1 U978 ( .A(n1290), .B(G113), .Z(n1184) );
NAND2_X1 U979 ( .A1(KEYINPUT32), .A2(n1291), .ZN(n1290) );
NAND2_X1 U980 ( .A1(n1292), .A2(n1176), .ZN(n1289) );
XNOR2_X1 U981 ( .A(n1194), .B(n1293), .ZN(n1176) );
XNOR2_X1 U982 ( .A(KEYINPUT41), .B(KEYINPUT26), .ZN(n1292) );
NAND2_X1 U983 ( .A1(KEYINPUT5), .A2(n1095), .ZN(n1284) );
INV_X1 U984 ( .A(G472), .ZN(n1095) );
AND4_X1 U985 ( .A1(n1076), .A2(n1238), .A3(n1225), .A4(n1228), .ZN(n1248) );
NAND2_X1 U986 ( .A1(n1255), .A2(n1294), .ZN(n1228) );
OR4_X1 U987 ( .A1(n1150), .A2(n1109), .A3(n1050), .A4(G898), .ZN(n1294) );
INV_X1 U988 ( .A(n1257), .ZN(n1050) );
NAND3_X1 U989 ( .A1(n1257), .A2(n1150), .A3(G952), .ZN(n1255) );
NAND2_X1 U990 ( .A1(G237), .A2(G234), .ZN(n1257) );
NOR2_X1 U991 ( .A1(n1083), .A2(n1080), .ZN(n1225) );
INV_X1 U992 ( .A(n1266), .ZN(n1080) );
NAND2_X1 U993 ( .A1(G221), .A2(n1295), .ZN(n1266) );
NAND2_X1 U994 ( .A1(G234), .A2(n1109), .ZN(n1295) );
XOR2_X1 U995 ( .A(n1116), .B(G469), .Z(n1083) );
NAND2_X1 U996 ( .A1(n1296), .A2(n1109), .ZN(n1116) );
XOR2_X1 U997 ( .A(n1297), .B(n1298), .Z(n1296) );
XOR2_X1 U998 ( .A(n1299), .B(n1195), .Z(n1298) );
XOR2_X1 U999 ( .A(n1300), .B(n1301), .Z(n1195) );
XOR2_X1 U1000 ( .A(G107), .B(G104), .Z(n1301) );
XOR2_X1 U1001 ( .A(n1133), .B(n1302), .Z(n1300) );
NOR2_X1 U1002 ( .A1(KEYINPUT11), .A2(n1303), .ZN(n1302) );
XNOR2_X1 U1003 ( .A(n1293), .B(KEYINPUT13), .ZN(n1133) );
NAND2_X1 U1004 ( .A1(n1304), .A2(KEYINPUT55), .ZN(n1299) );
XOR2_X1 U1005 ( .A(n1268), .B(n1305), .Z(n1304) );
NOR2_X1 U1006 ( .A1(G140), .A2(KEYINPUT61), .ZN(n1305) );
XOR2_X1 U1007 ( .A(n1306), .B(n1307), .Z(n1297) );
XNOR2_X1 U1008 ( .A(n1198), .B(KEYINPUT25), .ZN(n1307) );
NOR2_X1 U1009 ( .A1(n1136), .A2(G953), .ZN(n1198) );
INV_X1 U1010 ( .A(G227), .ZN(n1136) );
NAND2_X1 U1011 ( .A1(KEYINPUT53), .A2(n1194), .ZN(n1306) );
NAND2_X1 U1012 ( .A1(n1308), .A2(n1309), .ZN(n1194) );
NAND2_X1 U1013 ( .A1(n1135), .A2(n1310), .ZN(n1309) );
INV_X1 U1014 ( .A(G137), .ZN(n1310) );
NAND2_X1 U1015 ( .A1(n1311), .A2(G137), .ZN(n1308) );
XOR2_X1 U1016 ( .A(KEYINPUT47), .B(n1135), .Z(n1311) );
XOR2_X1 U1017 ( .A(G131), .B(G134), .Z(n1135) );
INV_X1 U1018 ( .A(n1043), .ZN(n1238) );
NAND2_X1 U1019 ( .A1(n1072), .A2(n1071), .ZN(n1043) );
NAND2_X1 U1020 ( .A1(G214), .A2(n1312), .ZN(n1071) );
INV_X1 U1021 ( .A(n1244), .ZN(n1072) );
NAND3_X1 U1022 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1244) );
NAND2_X1 U1023 ( .A1(KEYINPUT50), .A2(n1205), .ZN(n1315) );
INV_X1 U1024 ( .A(n1106), .ZN(n1205) );
OR3_X1 U1025 ( .A1(n1316), .A2(KEYINPUT50), .A3(n1107), .ZN(n1314) );
NAND2_X1 U1026 ( .A1(n1107), .A2(n1316), .ZN(n1313) );
NAND2_X1 U1027 ( .A1(KEYINPUT24), .A2(n1106), .ZN(n1316) );
NAND2_X1 U1028 ( .A1(G210), .A2(n1312), .ZN(n1106) );
NAND2_X1 U1029 ( .A1(n1288), .A2(n1109), .ZN(n1312) );
AND2_X1 U1030 ( .A1(n1112), .A2(n1109), .ZN(n1107) );
XNOR2_X1 U1031 ( .A(n1157), .B(n1317), .ZN(n1112) );
XNOR2_X1 U1032 ( .A(KEYINPUT16), .B(n1204), .ZN(n1317) );
XNOR2_X1 U1033 ( .A(n1293), .B(n1318), .ZN(n1204) );
XOR2_X1 U1034 ( .A(G125), .B(n1319), .Z(n1318) );
AND2_X1 U1035 ( .A1(n1150), .A2(G224), .ZN(n1319) );
XOR2_X1 U1036 ( .A(G128), .B(n1320), .Z(n1293) );
XOR2_X1 U1037 ( .A(G146), .B(G143), .Z(n1320) );
XOR2_X1 U1038 ( .A(n1321), .B(n1322), .Z(n1157) );
XOR2_X1 U1039 ( .A(n1323), .B(n1324), .Z(n1322) );
XNOR2_X1 U1040 ( .A(G113), .B(KEYINPUT45), .ZN(n1324) );
NAND3_X1 U1041 ( .A1(n1325), .A2(n1326), .A3(n1327), .ZN(n1323) );
NAND2_X1 U1042 ( .A1(KEYINPUT18), .A2(n1328), .ZN(n1327) );
NAND3_X1 U1043 ( .A1(G122), .A2(n1329), .A3(n1268), .ZN(n1326) );
NAND2_X1 U1044 ( .A1(G110), .A2(n1330), .ZN(n1325) );
NAND2_X1 U1045 ( .A1(n1331), .A2(n1329), .ZN(n1330) );
INV_X1 U1046 ( .A(KEYINPUT18), .ZN(n1329) );
XOR2_X1 U1047 ( .A(n1328), .B(KEYINPUT28), .Z(n1331) );
XOR2_X1 U1048 ( .A(n1332), .B(n1291), .Z(n1321) );
XOR2_X1 U1049 ( .A(G116), .B(G119), .Z(n1291) );
XNOR2_X1 U1050 ( .A(n1333), .B(n1303), .ZN(n1332) );
XNOR2_X1 U1051 ( .A(G101), .B(KEYINPUT48), .ZN(n1303) );
NAND2_X1 U1052 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
NAND2_X1 U1053 ( .A1(G104), .A2(n1038), .ZN(n1335) );
XOR2_X1 U1054 ( .A(KEYINPUT44), .B(n1336), .Z(n1334) );
NOR2_X1 U1055 ( .A1(G104), .A2(n1038), .ZN(n1336) );
INV_X1 U1056 ( .A(G107), .ZN(n1038) );
INV_X1 U1057 ( .A(n1056), .ZN(n1076) );
NAND2_X1 U1058 ( .A1(n1241), .A2(n1100), .ZN(n1056) );
XOR2_X1 U1059 ( .A(n1337), .B(G475), .Z(n1100) );
NAND2_X1 U1060 ( .A1(n1167), .A2(n1109), .ZN(n1337) );
XNOR2_X1 U1061 ( .A(n1338), .B(n1339), .ZN(n1167) );
XOR2_X1 U1062 ( .A(n1340), .B(n1341), .Z(n1339) );
XOR2_X1 U1063 ( .A(n1342), .B(n1128), .Z(n1341) );
XOR2_X1 U1064 ( .A(G125), .B(G140), .Z(n1128) );
NAND3_X1 U1065 ( .A1(n1288), .A2(n1150), .A3(G214), .ZN(n1342) );
INV_X1 U1066 ( .A(G237), .ZN(n1288) );
XOR2_X1 U1067 ( .A(n1343), .B(n1344), .Z(n1340) );
NOR2_X1 U1068 ( .A1(KEYINPUT12), .A2(n1237), .ZN(n1344) );
INV_X1 U1069 ( .A(G143), .ZN(n1237) );
NAND2_X1 U1070 ( .A1(n1345), .A2(n1346), .ZN(n1343) );
NAND2_X1 U1071 ( .A1(G113), .A2(n1328), .ZN(n1346) );
XOR2_X1 U1072 ( .A(n1347), .B(KEYINPUT2), .Z(n1345) );
OR2_X1 U1073 ( .A1(n1328), .A2(G113), .ZN(n1347) );
INV_X1 U1074 ( .A(G122), .ZN(n1328) );
XOR2_X1 U1075 ( .A(n1348), .B(n1349), .Z(n1338) );
XOR2_X1 U1076 ( .A(KEYINPUT27), .B(G146), .Z(n1349) );
XNOR2_X1 U1077 ( .A(G131), .B(G104), .ZN(n1348) );
XOR2_X1 U1078 ( .A(n1102), .B(G478), .Z(n1241) );
NAND2_X1 U1079 ( .A1(n1109), .A2(n1114), .ZN(n1102) );
NAND2_X1 U1080 ( .A1(n1350), .A2(n1351), .ZN(n1114) );
NAND2_X1 U1081 ( .A1(n1352), .A2(n1353), .ZN(n1351) );
XOR2_X1 U1082 ( .A(KEYINPUT17), .B(n1354), .Z(n1350) );
NOR2_X1 U1083 ( .A1(n1352), .A2(n1353), .ZN(n1354) );
NAND3_X1 U1084 ( .A1(n1282), .A2(n1150), .A3(G217), .ZN(n1353) );
INV_X1 U1085 ( .A(G953), .ZN(n1150) );
XNOR2_X1 U1086 ( .A(G234), .B(KEYINPUT42), .ZN(n1282) );
XNOR2_X1 U1087 ( .A(n1355), .B(n1356), .ZN(n1352) );
XOR2_X1 U1088 ( .A(G134), .B(n1357), .Z(n1356) );
XOR2_X1 U1089 ( .A(KEYINPUT1), .B(G143), .Z(n1357) );
XOR2_X1 U1090 ( .A(n1358), .B(n1359), .Z(n1355) );
NOR2_X1 U1091 ( .A1(G128), .A2(KEYINPUT23), .ZN(n1359) );
XOR2_X1 U1092 ( .A(n1360), .B(G107), .Z(n1358) );
NAND2_X1 U1093 ( .A1(KEYINPUT35), .A2(n1361), .ZN(n1360) );
XOR2_X1 U1094 ( .A(G122), .B(G116), .Z(n1361) );
INV_X1 U1095 ( .A(G902), .ZN(n1109) );
INV_X1 U1096 ( .A(G110), .ZN(n1268) );
endmodule


