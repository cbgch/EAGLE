//Key = 1001010111010011111111100001011000101011001110100100001001111101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398;

XOR2_X1 U753 ( .A(G107), .B(n1054), .Z(G9) );
NOR2_X1 U754 ( .A1(n1055), .A2(n1056), .ZN(G75) );
NOR4_X1 U755 ( .A1(G953), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1056) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U757 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR3_X1 U758 ( .A1(n1064), .A2(n1065), .A3(n1066), .ZN(n1063) );
NOR2_X1 U759 ( .A1(n1067), .A2(n1068), .ZN(n1065) );
NOR2_X1 U760 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
NOR2_X1 U761 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
NOR2_X1 U762 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NOR3_X1 U763 ( .A1(n1075), .A2(n1076), .A3(n1077), .ZN(n1073) );
NOR3_X1 U764 ( .A1(n1078), .A2(n1079), .A3(n1080), .ZN(n1077) );
INV_X1 U765 ( .A(KEYINPUT27), .ZN(n1078) );
NOR2_X1 U766 ( .A1(KEYINPUT27), .A2(n1081), .ZN(n1076) );
NOR2_X1 U767 ( .A1(n1082), .A2(n1081), .ZN(n1071) );
NOR2_X1 U768 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U769 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NOR3_X1 U770 ( .A1(n1074), .A2(n1087), .A3(n1081), .ZN(n1067) );
NOR2_X1 U771 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
NOR4_X1 U772 ( .A1(n1090), .A2(n1081), .A3(n1074), .A4(n1070), .ZN(n1062) );
INV_X1 U773 ( .A(n1091), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1092), .A2(n1093), .ZN(n1090) );
NOR3_X1 U775 ( .A1(n1057), .A2(G953), .A3(G952), .ZN(n1055) );
AND4_X1 U776 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1057) );
NOR4_X1 U777 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097) );
XOR2_X1 U778 ( .A(n1102), .B(n1103), .Z(n1101) );
NAND2_X1 U779 ( .A1(KEYINPUT39), .A2(n1104), .ZN(n1102) );
XOR2_X1 U780 ( .A(n1105), .B(n1106), .Z(n1100) );
NOR2_X1 U781 ( .A1(G475), .A2(KEYINPUT33), .ZN(n1106) );
XOR2_X1 U782 ( .A(n1107), .B(n1108), .Z(n1099) );
NAND2_X1 U783 ( .A1(KEYINPUT43), .A2(n1109), .ZN(n1107) );
XOR2_X1 U784 ( .A(n1110), .B(G469), .Z(n1096) );
XOR2_X1 U785 ( .A(n1111), .B(n1112), .Z(G72) );
XOR2_X1 U786 ( .A(n1113), .B(n1114), .Z(n1112) );
NOR2_X1 U787 ( .A1(n1115), .A2(n1116), .ZN(n1114) );
NOR2_X1 U788 ( .A1(n1117), .A2(n1118), .ZN(n1115) );
NAND2_X1 U789 ( .A1(n1119), .A2(n1120), .ZN(n1113) );
NAND2_X1 U790 ( .A1(G953), .A2(n1118), .ZN(n1120) );
XOR2_X1 U791 ( .A(n1121), .B(n1122), .Z(n1119) );
XOR2_X1 U792 ( .A(n1123), .B(n1124), .Z(n1122) );
XOR2_X1 U793 ( .A(G137), .B(G134), .Z(n1124) );
XOR2_X1 U794 ( .A(KEYINPUT45), .B(KEYINPUT44), .Z(n1123) );
XOR2_X1 U795 ( .A(n1125), .B(n1126), .Z(n1121) );
XNOR2_X1 U796 ( .A(G131), .B(n1127), .ZN(n1125) );
NAND2_X1 U797 ( .A1(n1116), .A2(n1128), .ZN(n1111) );
NAND2_X1 U798 ( .A1(n1129), .A2(n1130), .ZN(G69) );
NAND2_X1 U799 ( .A1(G953), .A2(n1131), .ZN(n1130) );
XOR2_X1 U800 ( .A(n1132), .B(n1133), .Z(n1129) );
NOR2_X1 U801 ( .A1(n1134), .A2(n1135), .ZN(n1133) );
NOR2_X1 U802 ( .A1(n1116), .A2(n1136), .ZN(n1135) );
NOR3_X1 U803 ( .A1(G953), .A2(n1137), .A3(n1138), .ZN(n1134) );
XOR2_X1 U804 ( .A(n1139), .B(KEYINPUT24), .Z(n1137) );
NAND4_X1 U805 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1139) );
XNOR2_X1 U806 ( .A(KEYINPUT5), .B(n1144), .ZN(n1140) );
NAND2_X1 U807 ( .A1(n1145), .A2(KEYINPUT42), .ZN(n1132) );
XOR2_X1 U808 ( .A(n1146), .B(n1147), .Z(n1145) );
NAND3_X1 U809 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1146) );
OR2_X1 U810 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
NAND2_X1 U811 ( .A1(KEYINPUT50), .A2(n1153), .ZN(n1149) );
NAND2_X1 U812 ( .A1(n1154), .A2(n1152), .ZN(n1153) );
XNOR2_X1 U813 ( .A(KEYINPUT34), .B(n1151), .ZN(n1154) );
NAND2_X1 U814 ( .A1(n1155), .A2(n1156), .ZN(n1148) );
INV_X1 U815 ( .A(KEYINPUT50), .ZN(n1156) );
NAND2_X1 U816 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
OR2_X1 U817 ( .A1(n1151), .A2(KEYINPUT34), .ZN(n1158) );
NAND3_X1 U818 ( .A1(n1152), .A2(n1151), .A3(KEYINPUT34), .ZN(n1157) );
NOR2_X1 U819 ( .A1(n1159), .A2(n1160), .ZN(G66) );
XOR2_X1 U820 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U821 ( .A(KEYINPUT52), .B(n1163), .Z(n1162) );
NOR2_X1 U822 ( .A1(n1109), .A2(n1164), .ZN(n1163) );
NOR2_X1 U823 ( .A1(n1159), .A2(n1165), .ZN(G63) );
NOR3_X1 U824 ( .A1(n1103), .A2(n1166), .A3(n1167), .ZN(n1165) );
NOR3_X1 U825 ( .A1(n1168), .A2(n1104), .A3(n1164), .ZN(n1167) );
NOR2_X1 U826 ( .A1(n1169), .A2(n1170), .ZN(n1166) );
NOR2_X1 U827 ( .A1(n1171), .A2(n1104), .ZN(n1170) );
INV_X1 U828 ( .A(G478), .ZN(n1104) );
NOR2_X1 U829 ( .A1(n1159), .A2(n1172), .ZN(G60) );
NOR3_X1 U830 ( .A1(n1173), .A2(n1174), .A3(n1175), .ZN(n1172) );
NOR3_X1 U831 ( .A1(n1176), .A2(n1177), .A3(n1164), .ZN(n1175) );
NOR2_X1 U832 ( .A1(n1178), .A2(n1179), .ZN(n1174) );
INV_X1 U833 ( .A(n1176), .ZN(n1179) );
NOR2_X1 U834 ( .A1(n1171), .A2(n1177), .ZN(n1178) );
INV_X1 U835 ( .A(G475), .ZN(n1177) );
XOR2_X1 U836 ( .A(n1180), .B(n1181), .Z(G6) );
NOR3_X1 U837 ( .A1(n1159), .A2(n1182), .A3(n1183), .ZN(G57) );
NOR2_X1 U838 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
NOR2_X1 U839 ( .A1(n1186), .A2(n1187), .ZN(n1185) );
NOR2_X1 U840 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
NOR2_X1 U841 ( .A1(n1190), .A2(n1191), .ZN(n1186) );
NOR2_X1 U842 ( .A1(n1192), .A2(n1193), .ZN(n1182) );
NOR2_X1 U843 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
NOR2_X1 U844 ( .A1(n1189), .A2(n1191), .ZN(n1195) );
XOR2_X1 U845 ( .A(n1190), .B(KEYINPUT29), .Z(n1189) );
NOR2_X1 U846 ( .A1(n1188), .A2(n1190), .ZN(n1194) );
XNOR2_X1 U847 ( .A(n1196), .B(n1197), .ZN(n1190) );
XNOR2_X1 U848 ( .A(n1198), .B(n1199), .ZN(n1197) );
XOR2_X1 U849 ( .A(n1200), .B(n1201), .Z(n1196) );
NOR2_X1 U850 ( .A1(n1202), .A2(n1164), .ZN(n1201) );
INV_X1 U851 ( .A(G472), .ZN(n1202) );
NAND2_X1 U852 ( .A1(KEYINPUT22), .A2(n1203), .ZN(n1200) );
INV_X1 U853 ( .A(n1191), .ZN(n1188) );
NOR2_X1 U854 ( .A1(n1159), .A2(n1204), .ZN(G54) );
XOR2_X1 U855 ( .A(n1205), .B(n1206), .Z(n1204) );
NOR2_X1 U856 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
XOR2_X1 U857 ( .A(n1209), .B(KEYINPUT54), .Z(n1208) );
NAND2_X1 U858 ( .A1(n1210), .A2(n1211), .ZN(n1209) );
NOR2_X1 U859 ( .A1(n1210), .A2(n1211), .ZN(n1207) );
AND2_X1 U860 ( .A1(n1212), .A2(n1213), .ZN(n1210) );
XOR2_X1 U861 ( .A(n1214), .B(KEYINPUT28), .Z(n1212) );
NAND2_X1 U862 ( .A1(n1215), .A2(n1116), .ZN(n1214) );
NOR2_X1 U863 ( .A1(n1216), .A2(n1164), .ZN(n1205) );
INV_X1 U864 ( .A(G469), .ZN(n1216) );
NOR2_X1 U865 ( .A1(n1159), .A2(n1217), .ZN(G51) );
XOR2_X1 U866 ( .A(n1218), .B(n1219), .Z(n1217) );
XOR2_X1 U867 ( .A(n1220), .B(n1221), .Z(n1219) );
NOR2_X1 U868 ( .A1(n1222), .A2(n1164), .ZN(n1220) );
NAND2_X1 U869 ( .A1(G902), .A2(n1059), .ZN(n1164) );
INV_X1 U870 ( .A(n1171), .ZN(n1059) );
NOR4_X1 U871 ( .A1(n1138), .A2(n1223), .A3(n1128), .A4(n1224), .ZN(n1171) );
NAND3_X1 U872 ( .A1(n1142), .A2(n1144), .A3(n1143), .ZN(n1224) );
NAND4_X1 U873 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1128) );
AND4_X1 U874 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
NAND3_X1 U875 ( .A1(n1233), .A2(n1234), .A3(n1075), .ZN(n1227) );
NAND2_X1 U876 ( .A1(n1235), .A2(n1236), .ZN(n1233) );
NAND4_X1 U877 ( .A1(n1092), .A2(n1084), .A3(n1237), .A4(n1238), .ZN(n1236) );
NAND3_X1 U878 ( .A1(n1089), .A2(n1091), .A3(n1093), .ZN(n1235) );
INV_X1 U879 ( .A(n1141), .ZN(n1223) );
NAND2_X1 U880 ( .A1(n1239), .A2(n1075), .ZN(n1141) );
XOR2_X1 U881 ( .A(n1240), .B(KEYINPUT60), .Z(n1239) );
NAND4_X1 U882 ( .A1(n1241), .A2(n1242), .A3(n1181), .A4(n1243), .ZN(n1138) );
NOR2_X1 U883 ( .A1(n1054), .A2(n1244), .ZN(n1243) );
INV_X1 U884 ( .A(n1245), .ZN(n1244) );
AND2_X1 U885 ( .A1(n1088), .A2(n1246), .ZN(n1054) );
NAND2_X1 U886 ( .A1(n1089), .A2(n1246), .ZN(n1181) );
AND4_X1 U887 ( .A1(n1084), .A2(n1247), .A3(n1094), .A4(n1248), .ZN(n1246) );
NAND2_X1 U888 ( .A1(n1249), .A2(n1250), .ZN(n1242) );
INV_X1 U889 ( .A(KEYINPUT51), .ZN(n1250) );
NAND3_X1 U890 ( .A1(n1075), .A2(n1251), .A3(KEYINPUT51), .ZN(n1241) );
XNOR2_X1 U891 ( .A(G210), .B(KEYINPUT26), .ZN(n1222) );
NOR2_X1 U892 ( .A1(n1116), .A2(G952), .ZN(n1159) );
XNOR2_X1 U893 ( .A(n1225), .B(n1252), .ZN(G48) );
NOR2_X1 U894 ( .A1(KEYINPUT10), .A2(n1253), .ZN(n1252) );
NAND3_X1 U895 ( .A1(n1089), .A2(n1075), .A3(n1254), .ZN(n1225) );
XOR2_X1 U896 ( .A(n1255), .B(n1256), .Z(G45) );
NAND4_X1 U897 ( .A1(n1238), .A2(n1234), .A3(n1237), .A4(n1257), .ZN(n1256) );
NOR3_X1 U898 ( .A1(n1258), .A2(n1259), .A3(n1260), .ZN(n1257) );
XOR2_X1 U899 ( .A(KEYINPUT38), .B(n1084), .Z(n1258) );
INV_X1 U900 ( .A(n1261), .ZN(n1237) );
XNOR2_X1 U901 ( .A(G140), .B(n1226), .ZN(G42) );
NAND3_X1 U902 ( .A1(n1262), .A2(n1089), .A3(n1093), .ZN(n1226) );
XOR2_X1 U903 ( .A(n1232), .B(n1263), .Z(G39) );
NAND2_X1 U904 ( .A1(KEYINPUT57), .A2(G137), .ZN(n1263) );
NAND3_X1 U905 ( .A1(n1264), .A2(n1095), .A3(n1254), .ZN(n1232) );
XOR2_X1 U906 ( .A(n1265), .B(n1231), .Z(G36) );
NAND3_X1 U907 ( .A1(n1092), .A2(n1088), .A3(n1262), .ZN(n1231) );
XNOR2_X1 U908 ( .A(G131), .B(n1230), .ZN(G33) );
NAND3_X1 U909 ( .A1(n1089), .A2(n1092), .A3(n1262), .ZN(n1230) );
AND3_X1 U910 ( .A1(n1084), .A2(n1234), .A3(n1095), .ZN(n1262) );
INV_X1 U911 ( .A(n1081), .ZN(n1095) );
NAND2_X1 U912 ( .A1(n1266), .A2(n1080), .ZN(n1081) );
XOR2_X1 U913 ( .A(n1267), .B(n1229), .Z(G30) );
NAND3_X1 U914 ( .A1(n1088), .A2(n1075), .A3(n1254), .ZN(n1229) );
AND4_X1 U915 ( .A1(n1084), .A2(n1066), .A3(n1064), .A4(n1234), .ZN(n1254) );
NAND2_X1 U916 ( .A1(n1268), .A2(n1269), .ZN(G3) );
NAND2_X1 U917 ( .A1(n1270), .A2(n1271), .ZN(n1269) );
XNOR2_X1 U918 ( .A(n1249), .B(KEYINPUT21), .ZN(n1270) );
NAND2_X1 U919 ( .A1(G101), .A2(n1272), .ZN(n1268) );
XNOR2_X1 U920 ( .A(n1249), .B(KEYINPUT53), .ZN(n1272) );
NOR2_X1 U921 ( .A1(n1251), .A2(n1259), .ZN(n1249) );
NAND4_X1 U922 ( .A1(n1264), .A2(n1092), .A3(n1084), .A4(n1273), .ZN(n1251) );
XNOR2_X1 U923 ( .A(G125), .B(n1274), .ZN(G27) );
NAND4_X1 U924 ( .A1(n1093), .A2(n1091), .A3(n1275), .A4(n1075), .ZN(n1274) );
NOR2_X1 U925 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U926 ( .A(n1089), .B(KEYINPUT55), .ZN(n1277) );
INV_X1 U927 ( .A(n1234), .ZN(n1276) );
NAND2_X1 U928 ( .A1(n1061), .A2(n1278), .ZN(n1234) );
NAND4_X1 U929 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1118), .ZN(n1278) );
INV_X1 U930 ( .A(G900), .ZN(n1118) );
XOR2_X1 U931 ( .A(n1142), .B(n1280), .Z(G24) );
XOR2_X1 U932 ( .A(KEYINPUT17), .B(G122), .Z(n1280) );
NAND4_X1 U933 ( .A1(n1094), .A2(n1281), .A3(n1282), .A4(n1248), .ZN(n1142) );
NOR2_X1 U934 ( .A1(n1283), .A2(n1261), .ZN(n1282) );
XNOR2_X1 U935 ( .A(G119), .B(n1143), .ZN(G21) );
NAND4_X1 U936 ( .A1(n1264), .A2(n1281), .A3(n1066), .A4(n1064), .ZN(n1143) );
INV_X1 U937 ( .A(n1248), .ZN(n1066) );
XOR2_X1 U938 ( .A(G116), .B(n1284), .Z(G18) );
NOR2_X1 U939 ( .A1(n1259), .A2(n1240), .ZN(n1284) );
NAND4_X1 U940 ( .A1(n1092), .A2(n1091), .A3(n1088), .A4(n1273), .ZN(n1240) );
AND2_X1 U941 ( .A1(n1285), .A2(n1238), .ZN(n1088) );
XNOR2_X1 U942 ( .A(KEYINPUT36), .B(n1286), .ZN(n1285) );
XNOR2_X1 U943 ( .A(n1287), .B(n1144), .ZN(G15) );
NAND3_X1 U944 ( .A1(n1092), .A2(n1281), .A3(n1089), .ZN(n1144) );
NOR2_X1 U945 ( .A1(n1238), .A2(n1261), .ZN(n1089) );
XOR2_X1 U946 ( .A(n1286), .B(KEYINPUT6), .Z(n1261) );
AND2_X1 U947 ( .A1(n1091), .A2(n1247), .ZN(n1281) );
NOR2_X1 U948 ( .A1(n1085), .A2(n1098), .ZN(n1091) );
INV_X1 U949 ( .A(n1086), .ZN(n1098) );
INV_X1 U950 ( .A(n1260), .ZN(n1092) );
NAND2_X1 U951 ( .A1(n1248), .A2(n1064), .ZN(n1260) );
NAND2_X1 U952 ( .A1(KEYINPUT0), .A2(n1288), .ZN(n1287) );
XOR2_X1 U953 ( .A(n1289), .B(n1245), .Z(G12) );
NAND4_X1 U954 ( .A1(n1093), .A2(n1264), .A3(n1084), .A4(n1247), .ZN(n1245) );
AND2_X1 U955 ( .A1(n1075), .A2(n1273), .ZN(n1247) );
NAND2_X1 U956 ( .A1(n1061), .A2(n1290), .ZN(n1273) );
NAND4_X1 U957 ( .A1(G953), .A2(G902), .A3(n1279), .A4(n1131), .ZN(n1290) );
INV_X1 U958 ( .A(G898), .ZN(n1131) );
NAND3_X1 U959 ( .A1(n1279), .A2(n1116), .A3(G952), .ZN(n1061) );
NAND2_X1 U960 ( .A1(G237), .A2(G234), .ZN(n1279) );
INV_X1 U961 ( .A(n1259), .ZN(n1075) );
NAND2_X1 U962 ( .A1(n1079), .A2(n1080), .ZN(n1259) );
NAND2_X1 U963 ( .A1(G214), .A2(n1291), .ZN(n1080) );
INV_X1 U964 ( .A(n1266), .ZN(n1079) );
XOR2_X1 U965 ( .A(n1292), .B(n1293), .Z(n1266) );
AND2_X1 U966 ( .A1(n1291), .A2(G210), .ZN(n1293) );
NAND2_X1 U967 ( .A1(n1294), .A2(n1295), .ZN(n1291) );
NAND2_X1 U968 ( .A1(n1296), .A2(n1294), .ZN(n1292) );
XOR2_X1 U969 ( .A(n1297), .B(n1221), .Z(n1296) );
XNOR2_X1 U970 ( .A(n1298), .B(n1151), .ZN(n1221) );
XNOR2_X1 U971 ( .A(n1180), .B(n1299), .ZN(n1151) );
XNOR2_X1 U972 ( .A(n1152), .B(n1147), .ZN(n1298) );
XOR2_X1 U973 ( .A(G110), .B(G122), .Z(n1147) );
NAND2_X1 U974 ( .A1(KEYINPUT16), .A2(n1218), .ZN(n1297) );
XOR2_X1 U975 ( .A(n1203), .B(n1300), .Z(n1218) );
XOR2_X1 U976 ( .A(n1301), .B(n1302), .Z(n1300) );
NOR2_X1 U977 ( .A1(G953), .A2(n1136), .ZN(n1301) );
INV_X1 U978 ( .A(G224), .ZN(n1136) );
AND2_X1 U979 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NAND2_X1 U980 ( .A1(G221), .A2(n1303), .ZN(n1086) );
XOR2_X1 U981 ( .A(n1110), .B(n1304), .Z(n1085) );
NOR2_X1 U982 ( .A1(G469), .A2(KEYINPUT13), .ZN(n1304) );
NAND2_X1 U983 ( .A1(n1305), .A2(n1294), .ZN(n1110) );
XOR2_X1 U984 ( .A(n1211), .B(n1306), .Z(n1305) );
XOR2_X1 U985 ( .A(KEYINPUT14), .B(n1307), .Z(n1306) );
NOR3_X1 U986 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1307) );
AND2_X1 U987 ( .A1(n1311), .A2(KEYINPUT25), .ZN(n1310) );
NOR2_X1 U988 ( .A1(KEYINPUT25), .A2(n1312), .ZN(n1309) );
INV_X1 U989 ( .A(n1215), .ZN(n1312) );
NOR2_X1 U990 ( .A1(n1311), .A2(n1117), .ZN(n1215) );
INV_X1 U991 ( .A(G227), .ZN(n1117) );
INV_X1 U992 ( .A(n1213), .ZN(n1308) );
NAND2_X1 U993 ( .A1(n1311), .A2(n1313), .ZN(n1213) );
NAND2_X1 U994 ( .A1(G227), .A2(n1116), .ZN(n1313) );
XNOR2_X1 U995 ( .A(n1289), .B(G140), .ZN(n1311) );
XNOR2_X1 U996 ( .A(n1314), .B(n1315), .ZN(n1211) );
XOR2_X1 U997 ( .A(n1299), .B(n1127), .Z(n1315) );
XNOR2_X1 U998 ( .A(n1316), .B(n1317), .ZN(n1127) );
XOR2_X1 U999 ( .A(n1253), .B(KEYINPUT59), .Z(n1316) );
XOR2_X1 U1000 ( .A(n1318), .B(n1184), .Z(n1299) );
XNOR2_X1 U1001 ( .A(n1198), .B(n1319), .ZN(n1314) );
NOR2_X1 U1002 ( .A1(G104), .A2(KEYINPUT31), .ZN(n1319) );
INV_X1 U1003 ( .A(n1070), .ZN(n1264) );
NAND2_X1 U1004 ( .A1(n1283), .A2(n1286), .ZN(n1070) );
NAND3_X1 U1005 ( .A1(n1320), .A2(n1321), .A3(n1322), .ZN(n1286) );
NAND2_X1 U1006 ( .A1(KEYINPUT48), .A2(n1173), .ZN(n1322) );
INV_X1 U1007 ( .A(n1105), .ZN(n1173) );
OR3_X1 U1008 ( .A1(n1323), .A2(KEYINPUT48), .A3(G475), .ZN(n1321) );
NAND2_X1 U1009 ( .A1(G475), .A2(n1323), .ZN(n1320) );
NAND2_X1 U1010 ( .A1(KEYINPUT8), .A2(n1105), .ZN(n1323) );
NAND2_X1 U1011 ( .A1(n1176), .A2(n1294), .ZN(n1105) );
XOR2_X1 U1012 ( .A(n1324), .B(n1325), .Z(n1176) );
XOR2_X1 U1013 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1014 ( .A(n1288), .B(G122), .Z(n1327) );
NAND2_X1 U1015 ( .A1(KEYINPUT30), .A2(n1328), .ZN(n1326) );
XOR2_X1 U1016 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1017 ( .A(n1255), .B(G131), .Z(n1330) );
INV_X1 U1018 ( .A(G143), .ZN(n1255) );
NAND4_X1 U1019 ( .A1(KEYINPUT18), .A2(G214), .A3(n1295), .A4(n1116), .ZN(n1329) );
XNOR2_X1 U1020 ( .A(n1126), .B(n1331), .ZN(n1324) );
XOR2_X1 U1021 ( .A(n1332), .B(n1333), .Z(n1331) );
NOR2_X1 U1022 ( .A1(G146), .A2(KEYINPUT37), .ZN(n1333) );
NOR2_X1 U1023 ( .A1(KEYINPUT41), .A2(n1180), .ZN(n1332) );
INV_X1 U1024 ( .A(G104), .ZN(n1180) );
XOR2_X1 U1025 ( .A(G140), .B(n1302), .Z(n1126) );
INV_X1 U1026 ( .A(n1238), .ZN(n1283) );
XOR2_X1 U1027 ( .A(n1103), .B(G478), .Z(n1238) );
NOR2_X1 U1028 ( .A1(n1169), .A2(G902), .ZN(n1103) );
INV_X1 U1029 ( .A(n1168), .ZN(n1169) );
NAND3_X1 U1030 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1168) );
NAND2_X1 U1031 ( .A1(KEYINPUT56), .A2(n1337), .ZN(n1336) );
OR3_X1 U1032 ( .A1(n1337), .A2(KEYINPUT56), .A3(n1338), .ZN(n1335) );
NAND2_X1 U1033 ( .A1(n1339), .A2(n1338), .ZN(n1334) );
NAND3_X1 U1034 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1338) );
NAND2_X1 U1035 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
NAND2_X1 U1036 ( .A1(KEYINPUT32), .A2(n1345), .ZN(n1341) );
NAND2_X1 U1037 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
XOR2_X1 U1038 ( .A(n1344), .B(KEYINPUT9), .Z(n1346) );
NAND2_X1 U1039 ( .A1(n1348), .A2(n1349), .ZN(n1340) );
INV_X1 U1040 ( .A(KEYINPUT32), .ZN(n1349) );
NAND2_X1 U1041 ( .A1(n1350), .A2(n1351), .ZN(n1348) );
NAND2_X1 U1042 ( .A1(n1344), .A2(n1352), .ZN(n1351) );
OR3_X1 U1043 ( .A1(n1344), .A2(n1343), .A3(n1352), .ZN(n1350) );
INV_X1 U1044 ( .A(KEYINPUT9), .ZN(n1352) );
INV_X1 U1045 ( .A(n1347), .ZN(n1343) );
NAND3_X1 U1046 ( .A1(n1353), .A2(n1354), .A3(n1355), .ZN(n1347) );
NAND2_X1 U1047 ( .A1(KEYINPUT40), .A2(n1317), .ZN(n1355) );
NAND3_X1 U1048 ( .A1(n1356), .A2(n1357), .A3(n1265), .ZN(n1354) );
INV_X1 U1049 ( .A(G134), .ZN(n1265) );
INV_X1 U1050 ( .A(n1317), .ZN(n1356) );
NAND2_X1 U1051 ( .A1(G134), .A2(n1358), .ZN(n1353) );
NAND2_X1 U1052 ( .A1(n1359), .A2(n1357), .ZN(n1358) );
INV_X1 U1053 ( .A(KEYINPUT40), .ZN(n1357) );
XOR2_X1 U1054 ( .A(KEYINPUT11), .B(n1317), .Z(n1359) );
NAND2_X1 U1055 ( .A1(n1360), .A2(n1361), .ZN(n1344) );
NAND2_X1 U1056 ( .A1(n1362), .A2(n1318), .ZN(n1361) );
INV_X1 U1057 ( .A(G107), .ZN(n1318) );
XOR2_X1 U1058 ( .A(n1363), .B(G122), .Z(n1362) );
INV_X1 U1059 ( .A(G116), .ZN(n1363) );
XOR2_X1 U1060 ( .A(n1364), .B(KEYINPUT23), .Z(n1360) );
NAND2_X1 U1061 ( .A1(G107), .A2(n1365), .ZN(n1364) );
XOR2_X1 U1062 ( .A(G122), .B(G116), .Z(n1365) );
NAND2_X1 U1063 ( .A1(n1366), .A2(n1367), .ZN(n1339) );
INV_X1 U1064 ( .A(KEYINPUT56), .ZN(n1367) );
XOR2_X1 U1065 ( .A(n1337), .B(KEYINPUT46), .Z(n1366) );
NAND2_X1 U1066 ( .A1(G217), .A2(n1368), .ZN(n1337) );
NOR2_X1 U1067 ( .A1(n1064), .A2(n1248), .ZN(n1093) );
XOR2_X1 U1068 ( .A(n1108), .B(n1109), .Z(n1248) );
NAND2_X1 U1069 ( .A1(G217), .A2(n1303), .ZN(n1109) );
NAND2_X1 U1070 ( .A1(G234), .A2(n1294), .ZN(n1303) );
NOR2_X1 U1071 ( .A1(n1161), .A2(G902), .ZN(n1108) );
XNOR2_X1 U1072 ( .A(n1369), .B(n1370), .ZN(n1161) );
AND2_X1 U1073 ( .A1(n1368), .A2(G221), .ZN(n1370) );
AND2_X1 U1074 ( .A1(G234), .A2(n1116), .ZN(n1368) );
XOR2_X1 U1075 ( .A(n1371), .B(G137), .Z(n1369) );
NAND3_X1 U1076 ( .A1(n1372), .A2(n1373), .A3(KEYINPUT3), .ZN(n1371) );
NAND2_X1 U1077 ( .A1(n1374), .A2(n1375), .ZN(n1373) );
XOR2_X1 U1078 ( .A(KEYINPUT19), .B(n1376), .Z(n1375) );
XNOR2_X1 U1079 ( .A(n1377), .B(KEYINPUT35), .ZN(n1374) );
NAND2_X1 U1080 ( .A1(n1378), .A2(n1377), .ZN(n1372) );
XNOR2_X1 U1081 ( .A(n1379), .B(n1302), .ZN(n1377) );
XOR2_X1 U1082 ( .A(G125), .B(KEYINPUT4), .Z(n1302) );
XOR2_X1 U1083 ( .A(n1380), .B(G146), .Z(n1379) );
NAND2_X1 U1084 ( .A1(KEYINPUT58), .A2(G140), .ZN(n1380) );
XOR2_X1 U1085 ( .A(KEYINPUT12), .B(n1376), .Z(n1378) );
XNOR2_X1 U1086 ( .A(n1381), .B(n1382), .ZN(n1376) );
XOR2_X1 U1087 ( .A(n1383), .B(G128), .Z(n1381) );
NAND2_X1 U1088 ( .A1(KEYINPUT7), .A2(G110), .ZN(n1383) );
INV_X1 U1089 ( .A(n1094), .ZN(n1064) );
XOR2_X1 U1090 ( .A(n1384), .B(G472), .Z(n1094) );
NAND2_X1 U1091 ( .A1(n1385), .A2(n1294), .ZN(n1384) );
INV_X1 U1092 ( .A(G902), .ZN(n1294) );
XOR2_X1 U1093 ( .A(n1386), .B(n1387), .Z(n1385) );
XOR2_X1 U1094 ( .A(n1388), .B(n1389), .Z(n1387) );
XOR2_X1 U1095 ( .A(n1191), .B(n1390), .Z(n1389) );
NOR2_X1 U1096 ( .A1(KEYINPUT2), .A2(n1198), .ZN(n1390) );
XNOR2_X1 U1097 ( .A(n1391), .B(G131), .ZN(n1198) );
NAND2_X1 U1098 ( .A1(KEYINPUT61), .A2(n1392), .ZN(n1391) );
XOR2_X1 U1099 ( .A(G137), .B(n1393), .Z(n1392) );
NOR2_X1 U1100 ( .A1(G134), .A2(KEYINPUT62), .ZN(n1393) );
NAND3_X1 U1101 ( .A1(n1295), .A2(n1116), .A3(G210), .ZN(n1191) );
INV_X1 U1102 ( .A(G953), .ZN(n1116) );
INV_X1 U1103 ( .A(G237), .ZN(n1295) );
NAND2_X1 U1104 ( .A1(KEYINPUT49), .A2(n1192), .ZN(n1388) );
INV_X1 U1105 ( .A(n1184), .ZN(n1192) );
XOR2_X1 U1106 ( .A(n1271), .B(KEYINPUT63), .Z(n1184) );
INV_X1 U1107 ( .A(G101), .ZN(n1271) );
XOR2_X1 U1108 ( .A(n1199), .B(n1203), .Z(n1386) );
AND2_X1 U1109 ( .A1(n1394), .A2(n1395), .ZN(n1203) );
NAND2_X1 U1110 ( .A1(n1317), .A2(n1253), .ZN(n1395) );
INV_X1 U1111 ( .A(G146), .ZN(n1253) );
NAND2_X1 U1112 ( .A1(n1396), .A2(G146), .ZN(n1394) );
XOR2_X1 U1113 ( .A(KEYINPUT20), .B(n1317), .Z(n1396) );
XNOR2_X1 U1114 ( .A(n1267), .B(G143), .ZN(n1317) );
INV_X1 U1115 ( .A(G128), .ZN(n1267) );
XNOR2_X1 U1116 ( .A(n1152), .B(KEYINPUT1), .ZN(n1199) );
XNOR2_X1 U1117 ( .A(n1397), .B(n1398), .ZN(n1152) );
XOR2_X1 U1118 ( .A(KEYINPUT47), .B(G116), .Z(n1398) );
XOR2_X1 U1119 ( .A(n1288), .B(n1382), .Z(n1397) );
XOR2_X1 U1120 ( .A(G119), .B(KEYINPUT15), .Z(n1382) );
INV_X1 U1121 ( .A(G113), .ZN(n1288) );
INV_X1 U1122 ( .A(G110), .ZN(n1289) );
endmodule


