//Key = 1010000101001000111000011101110000111000101101011000001000010001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
n1422;

XNOR2_X1 U782 ( .A(G107), .B(n1082), .ZN(G9) );
NOR2_X1 U783 ( .A1(n1083), .A2(n1084), .ZN(G75) );
AND3_X1 U784 ( .A1(n1085), .A2(G952), .A3(n1086), .ZN(n1084) );
AND3_X1 U785 ( .A1(n1087), .A2(n1088), .A3(n1089), .ZN(n1085) );
NAND2_X1 U786 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
NAND2_X1 U787 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
NAND4_X1 U788 ( .A1(n1094), .A2(n1095), .A3(n1096), .A4(n1097), .ZN(n1093) );
NAND2_X1 U789 ( .A1(n1098), .A2(n1099), .ZN(n1092) );
NAND2_X1 U790 ( .A1(n1100), .A2(n1101), .ZN(n1099) );
NAND3_X1 U791 ( .A1(n1096), .A2(n1102), .A3(n1094), .ZN(n1101) );
NAND2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NAND2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
NAND2_X1 U794 ( .A1(n1095), .A2(n1107), .ZN(n1100) );
NAND2_X1 U795 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
NAND2_X1 U796 ( .A1(n1096), .A2(n1110), .ZN(n1109) );
NAND2_X1 U797 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND3_X1 U798 ( .A1(G214), .A2(n1113), .A3(n1114), .ZN(n1112) );
NAND2_X1 U799 ( .A1(n1094), .A2(n1115), .ZN(n1108) );
NAND3_X1 U800 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1115) );
INV_X1 U801 ( .A(n1119), .ZN(n1118) );
NAND3_X1 U802 ( .A1(n1120), .A2(KEYINPUT29), .A3(n1121), .ZN(n1117) );
NAND2_X1 U803 ( .A1(n1122), .A2(n1123), .ZN(n1116) );
INV_X1 U804 ( .A(n1124), .ZN(n1090) );
NOR3_X1 U805 ( .A1(n1125), .A2(G953), .A3(n1126), .ZN(n1083) );
INV_X1 U806 ( .A(n1087), .ZN(n1126) );
NAND4_X1 U807 ( .A1(n1127), .A2(n1094), .A3(n1128), .A4(n1129), .ZN(n1087) );
NOR4_X1 U808 ( .A1(n1120), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1129) );
XOR2_X1 U809 ( .A(n1133), .B(G469), .Z(n1132) );
NAND2_X1 U810 ( .A1(KEYINPUT27), .A2(n1134), .ZN(n1133) );
XOR2_X1 U811 ( .A(n1135), .B(n1136), .Z(n1131) );
NAND2_X1 U812 ( .A1(KEYINPUT7), .A2(n1137), .ZN(n1135) );
NOR2_X1 U813 ( .A1(n1138), .A2(n1139), .ZN(n1130) );
NOR2_X1 U814 ( .A1(n1140), .A2(n1141), .ZN(n1128) );
XOR2_X1 U815 ( .A(n1142), .B(KEYINPUT59), .Z(n1141) );
XNOR2_X1 U816 ( .A(n1143), .B(n1144), .ZN(n1140) );
NOR2_X1 U817 ( .A1(KEYINPUT10), .A2(n1145), .ZN(n1144) );
XNOR2_X1 U818 ( .A(KEYINPUT50), .B(n1146), .ZN(n1145) );
XOR2_X1 U819 ( .A(n1147), .B(G472), .Z(n1127) );
XOR2_X1 U820 ( .A(KEYINPUT33), .B(G952), .Z(n1125) );
XOR2_X1 U821 ( .A(n1148), .B(n1149), .Z(G72) );
NOR2_X1 U822 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
XOR2_X1 U823 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U824 ( .A(KEYINPUT0), .B(G137), .Z(n1153) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1152) );
NAND2_X1 U826 ( .A1(n1156), .A2(n1157), .ZN(n1148) );
NAND2_X1 U827 ( .A1(n1158), .A2(n1088), .ZN(n1157) );
XOR2_X1 U828 ( .A(KEYINPUT25), .B(n1159), .Z(n1156) );
NOR2_X1 U829 ( .A1(n1088), .A2(n1160), .ZN(n1159) );
XOR2_X1 U830 ( .A(KEYINPUT53), .B(n1161), .Z(n1160) );
AND2_X1 U831 ( .A1(G227), .A2(G900), .ZN(n1161) );
XOR2_X1 U832 ( .A(n1162), .B(n1163), .Z(G69) );
XOR2_X1 U833 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND2_X1 U834 ( .A1(G953), .A2(n1166), .ZN(n1165) );
NAND2_X1 U835 ( .A1(G898), .A2(G224), .ZN(n1166) );
NAND2_X1 U836 ( .A1(n1167), .A2(n1168), .ZN(n1164) );
NAND2_X1 U837 ( .A1(n1169), .A2(n1170), .ZN(n1168) );
XOR2_X1 U838 ( .A(n1171), .B(n1172), .Z(n1167) );
XNOR2_X1 U839 ( .A(n1173), .B(n1174), .ZN(n1171) );
AND2_X1 U840 ( .A1(n1175), .A2(n1088), .ZN(n1162) );
NOR2_X1 U841 ( .A1(n1176), .A2(n1177), .ZN(G66) );
NOR3_X1 U842 ( .A1(n1143), .A2(n1178), .A3(n1179), .ZN(n1177) );
NOR3_X1 U843 ( .A1(n1180), .A2(n1146), .A3(n1181), .ZN(n1179) );
INV_X1 U844 ( .A(n1182), .ZN(n1180) );
NOR2_X1 U845 ( .A1(n1183), .A2(n1182), .ZN(n1178) );
NOR2_X1 U846 ( .A1(n1086), .A2(n1146), .ZN(n1183) );
NOR2_X1 U847 ( .A1(n1176), .A2(n1184), .ZN(G63) );
NOR3_X1 U848 ( .A1(n1136), .A2(n1185), .A3(n1186), .ZN(n1184) );
AND3_X1 U849 ( .A1(n1187), .A2(n1188), .A3(G478), .ZN(n1186) );
NOR2_X1 U850 ( .A1(n1189), .A2(n1187), .ZN(n1185) );
NOR2_X1 U851 ( .A1(n1086), .A2(n1137), .ZN(n1189) );
INV_X1 U852 ( .A(G478), .ZN(n1137) );
NOR2_X1 U853 ( .A1(n1176), .A2(n1190), .ZN(G60) );
NOR2_X1 U854 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
XOR2_X1 U855 ( .A(KEYINPUT4), .B(n1193), .Z(n1192) );
NOR3_X1 U856 ( .A1(n1194), .A2(n1139), .A3(n1181), .ZN(n1193) );
XNOR2_X1 U857 ( .A(KEYINPUT57), .B(n1195), .ZN(n1194) );
NOR2_X1 U858 ( .A1(n1196), .A2(n1195), .ZN(n1191) );
NOR2_X1 U859 ( .A1(n1139), .A2(n1181), .ZN(n1196) );
INV_X1 U860 ( .A(n1188), .ZN(n1181) );
XNOR2_X1 U861 ( .A(G104), .B(n1197), .ZN(G6) );
NOR2_X1 U862 ( .A1(n1176), .A2(n1198), .ZN(G57) );
NOR2_X1 U863 ( .A1(n1199), .A2(n1200), .ZN(n1198) );
XOR2_X1 U864 ( .A(KEYINPUT5), .B(n1201), .Z(n1200) );
NOR2_X1 U865 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
AND2_X1 U866 ( .A1(n1203), .A2(n1202), .ZN(n1199) );
XNOR2_X1 U867 ( .A(n1204), .B(n1205), .ZN(n1203) );
NOR4_X1 U868 ( .A1(n1206), .A2(n1207), .A3(KEYINPUT61), .A4(n1208), .ZN(n1205) );
NOR2_X1 U869 ( .A1(n1209), .A2(n1173), .ZN(n1208) );
NOR2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(n1207) );
XNOR2_X1 U871 ( .A(n1212), .B(n1213), .ZN(n1210) );
AND3_X1 U872 ( .A1(n1211), .A2(n1173), .A3(n1209), .ZN(n1206) );
NOR2_X1 U873 ( .A1(KEYINPUT11), .A2(n1214), .ZN(n1209) );
XNOR2_X1 U874 ( .A(n1212), .B(n1215), .ZN(n1214) );
INV_X1 U875 ( .A(KEYINPUT55), .ZN(n1211) );
NAND2_X1 U876 ( .A1(n1188), .A2(G472), .ZN(n1204) );
NOR2_X1 U877 ( .A1(n1176), .A2(n1216), .ZN(G54) );
NOR2_X1 U878 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
XOR2_X1 U879 ( .A(n1219), .B(n1220), .Z(n1218) );
AND2_X1 U880 ( .A1(G469), .A2(n1188), .ZN(n1220) );
NOR2_X1 U881 ( .A1(KEYINPUT14), .A2(n1221), .ZN(n1219) );
XOR2_X1 U882 ( .A(n1222), .B(n1223), .Z(n1221) );
NOR2_X1 U883 ( .A1(n1224), .A2(n1225), .ZN(n1217) );
INV_X1 U884 ( .A(KEYINPUT14), .ZN(n1225) );
XNOR2_X1 U885 ( .A(n1223), .B(n1222), .ZN(n1224) );
NAND3_X1 U886 ( .A1(n1226), .A2(n1227), .A3(n1228), .ZN(n1222) );
NAND2_X1 U887 ( .A1(KEYINPUT39), .A2(n1229), .ZN(n1228) );
NAND2_X1 U888 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
NAND2_X1 U889 ( .A1(G110), .A2(n1232), .ZN(n1231) );
NAND4_X1 U890 ( .A1(n1230), .A2(n1233), .A3(KEYINPUT40), .A4(G110), .ZN(n1227) );
NAND2_X1 U891 ( .A1(n1234), .A2(n1235), .ZN(n1226) );
NAND3_X1 U892 ( .A1(n1236), .A2(n1237), .A3(n1238), .ZN(n1234) );
NAND2_X1 U893 ( .A1(KEYINPUT40), .A2(KEYINPUT39), .ZN(n1238) );
NAND2_X1 U894 ( .A1(KEYINPUT26), .A2(n1230), .ZN(n1237) );
NAND2_X1 U895 ( .A1(n1239), .A2(n1240), .ZN(n1236) );
INV_X1 U896 ( .A(KEYINPUT26), .ZN(n1240) );
NAND2_X1 U897 ( .A1(n1230), .A2(n1241), .ZN(n1239) );
NAND2_X1 U898 ( .A1(n1233), .A2(n1232), .ZN(n1241) );
INV_X1 U899 ( .A(KEYINPUT40), .ZN(n1232) );
INV_X1 U900 ( .A(KEYINPUT39), .ZN(n1233) );
NOR3_X1 U901 ( .A1(n1176), .A2(n1242), .A3(n1243), .ZN(G51) );
NOR2_X1 U902 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
INV_X1 U903 ( .A(n1246), .ZN(n1245) );
NOR2_X1 U904 ( .A1(n1247), .A2(n1248), .ZN(n1244) );
NOR3_X1 U905 ( .A1(n1249), .A2(n1250), .A3(n1251), .ZN(n1248) );
AND2_X1 U906 ( .A1(n1249), .A2(n1250), .ZN(n1247) );
INV_X1 U907 ( .A(KEYINPUT45), .ZN(n1249) );
NOR2_X1 U908 ( .A1(n1252), .A2(n1246), .ZN(n1242) );
XNOR2_X1 U909 ( .A(n1253), .B(n1254), .ZN(n1246) );
XOR2_X1 U910 ( .A(n1255), .B(n1256), .Z(n1254) );
NOR2_X1 U911 ( .A1(KEYINPUT3), .A2(n1257), .ZN(n1256) );
NOR2_X1 U912 ( .A1(n1258), .A2(n1259), .ZN(n1255) );
XOR2_X1 U913 ( .A(n1260), .B(KEYINPUT18), .Z(n1259) );
NAND2_X1 U914 ( .A1(n1215), .A2(n1261), .ZN(n1260) );
NOR2_X1 U915 ( .A1(n1215), .A2(n1261), .ZN(n1258) );
NOR2_X1 U916 ( .A1(n1250), .A2(n1251), .ZN(n1252) );
INV_X1 U917 ( .A(KEYINPUT63), .ZN(n1251) );
NAND2_X1 U918 ( .A1(n1188), .A2(n1262), .ZN(n1250) );
NOR2_X1 U919 ( .A1(n1263), .A2(n1086), .ZN(n1188) );
NOR2_X1 U920 ( .A1(n1175), .A2(n1158), .ZN(n1086) );
NAND4_X1 U921 ( .A1(n1264), .A2(n1265), .A3(n1266), .A4(n1267), .ZN(n1158) );
AND4_X1 U922 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1267) );
NAND3_X1 U923 ( .A1(n1094), .A2(n1097), .A3(n1272), .ZN(n1266) );
NAND2_X1 U924 ( .A1(n1273), .A2(n1274), .ZN(n1097) );
NAND2_X1 U925 ( .A1(n1275), .A2(n1276), .ZN(n1175) );
AND4_X1 U926 ( .A1(n1082), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1276) );
NAND3_X1 U927 ( .A1(n1280), .A2(n1095), .A3(n1281), .ZN(n1082) );
AND4_X1 U928 ( .A1(n1282), .A2(n1283), .A3(n1197), .A4(n1284), .ZN(n1275) );
NAND3_X1 U929 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1284) );
NAND3_X1 U930 ( .A1(n1281), .A2(n1095), .A3(n1285), .ZN(n1197) );
NOR2_X1 U931 ( .A1(n1088), .A2(G952), .ZN(n1176) );
XNOR2_X1 U932 ( .A(G146), .B(n1264), .ZN(G48) );
NAND3_X1 U933 ( .A1(n1285), .A2(n1288), .A3(n1289), .ZN(n1264) );
XNOR2_X1 U934 ( .A(G143), .B(n1265), .ZN(G45) );
NAND4_X1 U935 ( .A1(n1290), .A2(n1272), .A3(n1288), .A4(n1291), .ZN(n1265) );
INV_X1 U936 ( .A(n1292), .ZN(n1272) );
NAND2_X1 U937 ( .A1(n1293), .A2(n1294), .ZN(G42) );
NAND2_X1 U938 ( .A1(n1295), .A2(n1230), .ZN(n1294) );
XOR2_X1 U939 ( .A(KEYINPUT24), .B(n1296), .Z(n1293) );
NOR2_X1 U940 ( .A1(n1295), .A2(n1230), .ZN(n1296) );
INV_X1 U941 ( .A(G140), .ZN(n1230) );
INV_X1 U942 ( .A(n1271), .ZN(n1295) );
NAND3_X1 U943 ( .A1(n1094), .A2(n1119), .A3(n1297), .ZN(n1271) );
XNOR2_X1 U944 ( .A(G137), .B(n1270), .ZN(G39) );
NAND3_X1 U945 ( .A1(n1094), .A2(n1098), .A3(n1289), .ZN(n1270) );
INV_X1 U946 ( .A(n1298), .ZN(n1094) );
XOR2_X1 U947 ( .A(G134), .B(n1299), .Z(G36) );
NOR2_X1 U948 ( .A1(n1298), .A2(n1300), .ZN(n1299) );
XOR2_X1 U949 ( .A(KEYINPUT42), .B(n1301), .Z(n1300) );
NOR2_X1 U950 ( .A1(n1273), .A2(n1292), .ZN(n1301) );
XOR2_X1 U951 ( .A(n1302), .B(n1303), .Z(G33) );
NOR2_X1 U952 ( .A1(KEYINPUT46), .A2(n1304), .ZN(n1303) );
INV_X1 U953 ( .A(G131), .ZN(n1304) );
NOR3_X1 U954 ( .A1(n1305), .A2(n1274), .A3(n1292), .ZN(n1302) );
NAND3_X1 U955 ( .A1(n1119), .A2(n1306), .A3(n1287), .ZN(n1292) );
XNOR2_X1 U956 ( .A(KEYINPUT9), .B(n1298), .ZN(n1305) );
NAND2_X1 U957 ( .A1(n1114), .A2(n1307), .ZN(n1298) );
NAND2_X1 U958 ( .A1(G214), .A2(n1113), .ZN(n1307) );
XNOR2_X1 U959 ( .A(G128), .B(n1269), .ZN(G30) );
NAND3_X1 U960 ( .A1(n1280), .A2(n1288), .A3(n1289), .ZN(n1269) );
AND4_X1 U961 ( .A1(n1119), .A2(n1106), .A3(n1308), .A4(n1306), .ZN(n1289) );
XNOR2_X1 U962 ( .A(G101), .B(n1283), .ZN(G3) );
NAND3_X1 U963 ( .A1(n1281), .A2(n1098), .A3(n1287), .ZN(n1283) );
XNOR2_X1 U964 ( .A(G125), .B(n1268), .ZN(G27) );
NAND3_X1 U965 ( .A1(n1288), .A2(n1096), .A3(n1297), .ZN(n1268) );
AND4_X1 U966 ( .A1(n1105), .A2(n1285), .A3(n1106), .A4(n1306), .ZN(n1297) );
NAND2_X1 U967 ( .A1(n1124), .A2(n1309), .ZN(n1306) );
NAND3_X1 U968 ( .A1(G902), .A2(n1310), .A3(n1150), .ZN(n1309) );
NOR2_X1 U969 ( .A1(n1311), .A2(G900), .ZN(n1150) );
INV_X1 U970 ( .A(n1274), .ZN(n1285) );
XNOR2_X1 U971 ( .A(G122), .B(n1282), .ZN(G24) );
NAND4_X1 U972 ( .A1(n1286), .A2(n1095), .A3(n1290), .A4(n1291), .ZN(n1282) );
NOR2_X1 U973 ( .A1(n1308), .A2(n1106), .ZN(n1095) );
XNOR2_X1 U974 ( .A(G119), .B(n1279), .ZN(G21) );
NAND4_X1 U975 ( .A1(n1286), .A2(n1098), .A3(n1106), .A4(n1308), .ZN(n1279) );
XNOR2_X1 U976 ( .A(G116), .B(n1278), .ZN(G18) );
NAND3_X1 U977 ( .A1(n1286), .A2(n1280), .A3(n1287), .ZN(n1278) );
AND3_X1 U978 ( .A1(n1096), .A2(n1312), .A3(n1288), .ZN(n1286) );
XOR2_X1 U979 ( .A(n1313), .B(n1314), .Z(G15) );
NOR2_X1 U980 ( .A1(G113), .A2(KEYINPUT52), .ZN(n1314) );
NAND4_X1 U981 ( .A1(n1315), .A2(n1096), .A3(n1316), .A4(n1317), .ZN(n1313) );
NOR2_X1 U982 ( .A1(n1103), .A2(n1274), .ZN(n1317) );
NAND2_X1 U983 ( .A1(n1318), .A2(n1291), .ZN(n1274) );
XNOR2_X1 U984 ( .A(KEYINPUT32), .B(n1290), .ZN(n1318) );
INV_X1 U985 ( .A(n1287), .ZN(n1103) );
NOR2_X1 U986 ( .A1(n1106), .A2(n1105), .ZN(n1287) );
XNOR2_X1 U987 ( .A(KEYINPUT43), .B(n1312), .ZN(n1316) );
NAND2_X1 U988 ( .A1(n1319), .A2(n1320), .ZN(n1096) );
NAND2_X1 U989 ( .A1(n1119), .A2(n1123), .ZN(n1320) );
INV_X1 U990 ( .A(KEYINPUT29), .ZN(n1123) );
NAND3_X1 U991 ( .A1(n1121), .A2(n1321), .A3(KEYINPUT29), .ZN(n1319) );
XNOR2_X1 U992 ( .A(KEYINPUT56), .B(n1111), .ZN(n1315) );
INV_X1 U993 ( .A(n1288), .ZN(n1111) );
XNOR2_X1 U994 ( .A(G110), .B(n1277), .ZN(G12) );
NAND4_X1 U995 ( .A1(n1105), .A2(n1281), .A3(n1098), .A4(n1106), .ZN(n1277) );
XNOR2_X1 U996 ( .A(n1143), .B(n1146), .ZN(n1106) );
NAND2_X1 U997 ( .A1(G217), .A2(n1322), .ZN(n1146) );
NOR2_X1 U998 ( .A1(n1182), .A2(G902), .ZN(n1143) );
XNOR2_X1 U999 ( .A(n1323), .B(n1324), .ZN(n1182) );
XNOR2_X1 U1000 ( .A(n1235), .B(n1325), .ZN(n1324) );
XOR2_X1 U1001 ( .A(G137), .B(G119), .Z(n1325) );
XOR2_X1 U1002 ( .A(n1326), .B(n1327), .Z(n1323) );
XNOR2_X1 U1003 ( .A(n1328), .B(n1329), .ZN(n1327) );
NOR2_X1 U1004 ( .A1(KEYINPUT19), .A2(n1330), .ZN(n1329) );
INV_X1 U1005 ( .A(G128), .ZN(n1330) );
NAND2_X1 U1006 ( .A1(KEYINPUT23), .A2(n1331), .ZN(n1328) );
NAND2_X1 U1007 ( .A1(n1332), .A2(n1333), .ZN(n1331) );
NAND2_X1 U1008 ( .A1(n1334), .A2(n1335), .ZN(n1333) );
XOR2_X1 U1009 ( .A(n1336), .B(KEYINPUT30), .Z(n1332) );
OR2_X1 U1010 ( .A1(n1334), .A2(n1335), .ZN(n1336) );
INV_X1 U1011 ( .A(G146), .ZN(n1335) );
XNOR2_X1 U1012 ( .A(n1337), .B(n1261), .ZN(n1334) );
NAND2_X1 U1013 ( .A1(KEYINPUT2), .A2(G140), .ZN(n1337) );
NAND2_X1 U1014 ( .A1(n1338), .A2(G221), .ZN(n1326) );
NAND2_X1 U1015 ( .A1(n1339), .A2(n1340), .ZN(n1098) );
OR3_X1 U1016 ( .A1(n1291), .A2(n1290), .A3(KEYINPUT32), .ZN(n1340) );
NAND2_X1 U1017 ( .A1(KEYINPUT32), .A2(n1280), .ZN(n1339) );
INV_X1 U1018 ( .A(n1273), .ZN(n1280) );
NAND2_X1 U1019 ( .A1(n1341), .A2(n1290), .ZN(n1273) );
XNOR2_X1 U1020 ( .A(n1136), .B(n1342), .ZN(n1290) );
NOR2_X1 U1021 ( .A1(G478), .A2(KEYINPUT22), .ZN(n1342) );
NOR2_X1 U1022 ( .A1(n1187), .A2(G902), .ZN(n1136) );
XOR2_X1 U1023 ( .A(n1343), .B(n1344), .Z(n1187) );
NOR2_X1 U1024 ( .A1(KEYINPUT60), .A2(n1345), .ZN(n1344) );
XOR2_X1 U1025 ( .A(n1346), .B(n1347), .Z(n1345) );
XNOR2_X1 U1026 ( .A(n1348), .B(n1349), .ZN(n1347) );
NAND2_X1 U1027 ( .A1(KEYINPUT54), .A2(n1350), .ZN(n1348) );
XNOR2_X1 U1028 ( .A(n1351), .B(G107), .ZN(n1346) );
NAND2_X1 U1029 ( .A1(G217), .A2(n1338), .ZN(n1343) );
AND2_X1 U1030 ( .A1(G234), .A2(n1088), .ZN(n1338) );
INV_X1 U1031 ( .A(n1291), .ZN(n1341) );
NAND2_X1 U1032 ( .A1(n1142), .A2(n1352), .ZN(n1291) );
OR2_X1 U1033 ( .A1(n1139), .A2(n1138), .ZN(n1352) );
NAND2_X1 U1034 ( .A1(n1138), .A2(n1139), .ZN(n1142) );
INV_X1 U1035 ( .A(G475), .ZN(n1139) );
NOR2_X1 U1036 ( .A1(n1195), .A2(G902), .ZN(n1138) );
XOR2_X1 U1037 ( .A(n1353), .B(n1354), .Z(n1195) );
XNOR2_X1 U1038 ( .A(n1155), .B(n1355), .ZN(n1354) );
XOR2_X1 U1039 ( .A(n1356), .B(n1357), .Z(n1355) );
NOR2_X1 U1040 ( .A1(G146), .A2(KEYINPUT37), .ZN(n1357) );
NAND2_X1 U1041 ( .A1(KEYINPUT34), .A2(n1358), .ZN(n1356) );
XNOR2_X1 U1042 ( .A(n1359), .B(n1261), .ZN(n1155) );
XNOR2_X1 U1043 ( .A(G131), .B(G140), .ZN(n1359) );
XOR2_X1 U1044 ( .A(n1360), .B(n1361), .Z(n1353) );
XOR2_X1 U1045 ( .A(n1362), .B(n1363), .Z(n1361) );
NOR2_X1 U1046 ( .A1(G113), .A2(KEYINPUT51), .ZN(n1363) );
AND3_X1 U1047 ( .A1(G214), .A2(n1088), .A3(n1364), .ZN(n1362) );
XNOR2_X1 U1048 ( .A(G122), .B(G143), .ZN(n1360) );
AND3_X1 U1049 ( .A1(n1288), .A2(n1312), .A3(n1119), .ZN(n1281) );
NOR2_X1 U1050 ( .A1(n1121), .A2(n1120), .ZN(n1119) );
INV_X1 U1051 ( .A(n1321), .ZN(n1120) );
NAND2_X1 U1052 ( .A1(G221), .A2(n1322), .ZN(n1321) );
NAND2_X1 U1053 ( .A1(G234), .A2(n1365), .ZN(n1322) );
INV_X1 U1054 ( .A(n1122), .ZN(n1121) );
XNOR2_X1 U1055 ( .A(n1134), .B(G469), .ZN(n1122) );
NAND2_X1 U1056 ( .A1(n1366), .A2(n1263), .ZN(n1134) );
XOR2_X1 U1057 ( .A(n1223), .B(n1367), .Z(n1366) );
XNOR2_X1 U1058 ( .A(G110), .B(G140), .ZN(n1367) );
XOR2_X1 U1059 ( .A(n1368), .B(n1369), .Z(n1223) );
XOR2_X1 U1060 ( .A(n1370), .B(n1371), .Z(n1369) );
XNOR2_X1 U1061 ( .A(n1372), .B(n1373), .ZN(n1371) );
NAND2_X1 U1062 ( .A1(n1374), .A2(n1375), .ZN(n1372) );
NAND2_X1 U1063 ( .A1(G104), .A2(n1376), .ZN(n1375) );
XOR2_X1 U1064 ( .A(KEYINPUT28), .B(n1377), .Z(n1374) );
NOR2_X1 U1065 ( .A1(G104), .A2(n1376), .ZN(n1377) );
NAND2_X1 U1066 ( .A1(G227), .A2(n1088), .ZN(n1370) );
XOR2_X1 U1067 ( .A(n1154), .B(n1378), .Z(n1368) );
XOR2_X1 U1068 ( .A(n1350), .B(n1379), .Z(n1154) );
NOR2_X1 U1069 ( .A1(G146), .A2(KEYINPUT44), .ZN(n1379) );
XNOR2_X1 U1070 ( .A(G128), .B(n1380), .ZN(n1350) );
XOR2_X1 U1071 ( .A(G143), .B(G134), .Z(n1380) );
NAND2_X1 U1072 ( .A1(n1124), .A2(n1381), .ZN(n1312) );
NAND4_X1 U1073 ( .A1(n1169), .A2(n1170), .A3(G902), .A4(n1310), .ZN(n1381) );
INV_X1 U1074 ( .A(n1311), .ZN(n1170) );
XOR2_X1 U1075 ( .A(G953), .B(KEYINPUT36), .Z(n1311) );
XNOR2_X1 U1076 ( .A(G898), .B(KEYINPUT62), .ZN(n1169) );
NAND3_X1 U1077 ( .A1(n1310), .A2(n1088), .A3(G952), .ZN(n1124) );
NAND2_X1 U1078 ( .A1(G237), .A2(G234), .ZN(n1310) );
NOR2_X1 U1079 ( .A1(n1114), .A2(n1382), .ZN(n1288) );
AND2_X1 U1080 ( .A1(G214), .A2(n1113), .ZN(n1382) );
XOR2_X1 U1081 ( .A(n1383), .B(n1262), .Z(n1114) );
AND2_X1 U1082 ( .A1(G210), .A2(n1113), .ZN(n1262) );
NAND2_X1 U1083 ( .A1(n1365), .A2(n1364), .ZN(n1113) );
XNOR2_X1 U1084 ( .A(n1263), .B(KEYINPUT35), .ZN(n1365) );
NAND2_X1 U1085 ( .A1(n1384), .A2(n1263), .ZN(n1383) );
XOR2_X1 U1086 ( .A(n1385), .B(n1386), .Z(n1384) );
XNOR2_X1 U1087 ( .A(n1257), .B(n1261), .ZN(n1386) );
XOR2_X1 U1088 ( .A(G125), .B(KEYINPUT12), .Z(n1261) );
NAND2_X1 U1089 ( .A1(G224), .A2(n1088), .ZN(n1257) );
XNOR2_X1 U1090 ( .A(n1253), .B(n1215), .ZN(n1385) );
XOR2_X1 U1091 ( .A(n1387), .B(n1174), .Z(n1253) );
XNOR2_X1 U1092 ( .A(n1235), .B(n1388), .ZN(n1174) );
XNOR2_X1 U1093 ( .A(KEYINPUT48), .B(n1351), .ZN(n1388) );
INV_X1 U1094 ( .A(G122), .ZN(n1351) );
INV_X1 U1095 ( .A(G110), .ZN(n1235) );
NAND2_X1 U1096 ( .A1(KEYINPUT16), .A2(n1389), .ZN(n1387) );
XOR2_X1 U1097 ( .A(n1390), .B(n1172), .Z(n1389) );
XNOR2_X1 U1098 ( .A(n1391), .B(n1392), .ZN(n1172) );
XNOR2_X1 U1099 ( .A(KEYINPUT38), .B(n1373), .ZN(n1392) );
NAND3_X1 U1100 ( .A1(n1393), .A2(n1394), .A3(n1395), .ZN(n1391) );
NAND2_X1 U1101 ( .A1(KEYINPUT20), .A2(n1396), .ZN(n1395) );
NAND2_X1 U1102 ( .A1(n1376), .A2(n1397), .ZN(n1396) );
NAND2_X1 U1103 ( .A1(KEYINPUT49), .A2(G104), .ZN(n1397) );
NAND4_X1 U1104 ( .A1(n1398), .A2(n1399), .A3(n1376), .A4(G104), .ZN(n1394) );
NAND2_X1 U1105 ( .A1(n1400), .A2(n1358), .ZN(n1393) );
INV_X1 U1106 ( .A(G104), .ZN(n1358) );
NAND3_X1 U1107 ( .A1(n1401), .A2(n1402), .A3(n1403), .ZN(n1400) );
NAND2_X1 U1108 ( .A1(KEYINPUT20), .A2(n1399), .ZN(n1403) );
INV_X1 U1109 ( .A(KEYINPUT49), .ZN(n1399) );
NAND2_X1 U1110 ( .A1(KEYINPUT41), .A2(n1376), .ZN(n1402) );
NAND2_X1 U1111 ( .A1(n1404), .A2(n1405), .ZN(n1401) );
INV_X1 U1112 ( .A(KEYINPUT41), .ZN(n1405) );
NAND2_X1 U1113 ( .A1(n1376), .A2(n1406), .ZN(n1404) );
NAND2_X1 U1114 ( .A1(KEYINPUT49), .A2(n1398), .ZN(n1406) );
INV_X1 U1115 ( .A(KEYINPUT20), .ZN(n1398) );
INV_X1 U1116 ( .A(G107), .ZN(n1376) );
NOR2_X1 U1117 ( .A1(KEYINPUT13), .A2(n1407), .ZN(n1390) );
XNOR2_X1 U1118 ( .A(n1173), .B(KEYINPUT17), .ZN(n1407) );
INV_X1 U1119 ( .A(n1308), .ZN(n1105) );
XOR2_X1 U1120 ( .A(G472), .B(n1408), .Z(n1308) );
NOR2_X1 U1121 ( .A1(KEYINPUT15), .A2(n1147), .ZN(n1408) );
NAND2_X1 U1122 ( .A1(n1409), .A2(n1410), .ZN(n1147) );
XOR2_X1 U1123 ( .A(n1411), .B(n1412), .Z(n1410) );
XNOR2_X1 U1124 ( .A(n1215), .B(n1202), .ZN(n1412) );
AND2_X1 U1125 ( .A1(n1413), .A2(n1414), .ZN(n1202) );
NAND2_X1 U1126 ( .A1(n1415), .A2(n1373), .ZN(n1414) );
INV_X1 U1127 ( .A(G101), .ZN(n1373) );
NAND3_X1 U1128 ( .A1(n1364), .A2(n1088), .A3(G210), .ZN(n1415) );
NAND4_X1 U1129 ( .A1(n1364), .A2(n1088), .A3(G210), .A4(G101), .ZN(n1413) );
INV_X1 U1130 ( .A(G953), .ZN(n1088) );
INV_X1 U1131 ( .A(G237), .ZN(n1364) );
INV_X1 U1132 ( .A(n1213), .ZN(n1215) );
XNOR2_X1 U1133 ( .A(n1416), .B(n1417), .ZN(n1213) );
NOR2_X1 U1134 ( .A1(KEYINPUT8), .A2(G128), .ZN(n1417) );
XNOR2_X1 U1135 ( .A(G143), .B(G146), .ZN(n1416) );
XNOR2_X1 U1136 ( .A(n1173), .B(n1418), .ZN(n1411) );
NOR2_X1 U1137 ( .A1(KEYINPUT21), .A2(n1212), .ZN(n1418) );
XNOR2_X1 U1138 ( .A(n1378), .B(G134), .ZN(n1212) );
XOR2_X1 U1139 ( .A(n1419), .B(n1420), .Z(n1378) );
NOR2_X1 U1140 ( .A1(G131), .A2(KEYINPUT58), .ZN(n1420) );
NOR2_X1 U1141 ( .A1(G137), .A2(KEYINPUT31), .ZN(n1419) );
XNOR2_X1 U1142 ( .A(n1421), .B(n1422), .ZN(n1173) );
XOR2_X1 U1143 ( .A(KEYINPUT1), .B(G119), .Z(n1422) );
XNOR2_X1 U1144 ( .A(G113), .B(n1349), .ZN(n1421) );
XOR2_X1 U1145 ( .A(G116), .B(KEYINPUT6), .Z(n1349) );
XNOR2_X1 U1146 ( .A(KEYINPUT47), .B(n1263), .ZN(n1409) );
INV_X1 U1147 ( .A(G902), .ZN(n1263) );
endmodule


