//Key = 0010010000001110001001001111110001011011000011111110010110011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385;

NAND2_X1 U760 ( .A1(n1047), .A2(n1048), .ZN(G9) );
NAND2_X1 U761 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
XOR2_X1 U762 ( .A(n1051), .B(KEYINPUT34), .Z(n1047) );
NAND2_X1 U763 ( .A1(G107), .A2(n1052), .ZN(n1051) );
NAND4_X1 U764 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(G75) );
NOR2_X1 U765 ( .A1(n1057), .A2(n1058), .ZN(n1056) );
NAND4_X1 U766 ( .A1(n1059), .A2(n1060), .A3(n1061), .A4(n1062), .ZN(n1055) );
NOR4_X1 U767 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062) );
AND2_X1 U768 ( .A1(n1067), .A2(G478), .ZN(n1065) );
NOR2_X1 U769 ( .A1(n1068), .A2(n1069), .ZN(n1061) );
XOR2_X1 U770 ( .A(n1070), .B(n1071), .Z(n1069) );
XOR2_X1 U771 ( .A(n1072), .B(KEYINPUT16), .Z(n1071) );
OR2_X1 U772 ( .A1(n1073), .A2(KEYINPUT3), .ZN(n1060) );
NAND2_X1 U773 ( .A1(KEYINPUT3), .A2(n1074), .ZN(n1059) );
NAND3_X1 U774 ( .A1(n1075), .A2(n1076), .A3(G469), .ZN(n1074) );
NAND2_X1 U775 ( .A1(n1077), .A2(n1078), .ZN(n1053) );
NAND2_X1 U776 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
OR3_X1 U777 ( .A1(n1081), .A2(n1068), .A3(n1082), .ZN(n1080) );
INV_X1 U778 ( .A(n1083), .ZN(n1068) );
NAND2_X1 U779 ( .A1(n1084), .A2(n1085), .ZN(n1079) );
NAND2_X1 U780 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND3_X1 U781 ( .A1(n1083), .A2(n1088), .A3(n1089), .ZN(n1087) );
NAND2_X1 U782 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
OR2_X1 U783 ( .A1(n1075), .A2(n1092), .ZN(n1091) );
NAND2_X1 U784 ( .A1(n1073), .A2(n1093), .ZN(n1086) );
NAND2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1093) );
NAND2_X1 U786 ( .A1(n1089), .A2(n1096), .ZN(n1095) );
OR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U788 ( .A1(n1083), .A2(n1099), .ZN(n1094) );
NAND3_X1 U789 ( .A1(n1100), .A2(n1101), .A3(n1102), .ZN(n1099) );
OR2_X1 U790 ( .A1(n1103), .A2(KEYINPUT28), .ZN(n1101) );
NAND3_X1 U791 ( .A1(n1064), .A2(n1104), .A3(KEYINPUT28), .ZN(n1100) );
INV_X1 U792 ( .A(n1105), .ZN(n1077) );
NAND3_X1 U793 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(G72) );
XOR2_X1 U794 ( .A(n1109), .B(KEYINPUT31), .Z(n1108) );
NAND3_X1 U795 ( .A1(n1110), .A2(n1111), .A3(G953), .ZN(n1109) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1110) );
NAND2_X1 U797 ( .A1(n1112), .A2(n1054), .ZN(n1107) );
XNOR2_X1 U798 ( .A(n1058), .B(n1111), .ZN(n1112) );
NAND4_X1 U799 ( .A1(G900), .A2(G227), .A3(n1113), .A4(G953), .ZN(n1106) );
INV_X1 U800 ( .A(n1111), .ZN(n1113) );
NAND2_X1 U801 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NAND2_X1 U802 ( .A1(n1116), .A2(G953), .ZN(n1115) );
XNOR2_X1 U803 ( .A(G900), .B(KEYINPUT58), .ZN(n1116) );
XOR2_X1 U804 ( .A(n1117), .B(n1118), .Z(n1114) );
XNOR2_X1 U805 ( .A(n1119), .B(n1120), .ZN(n1118) );
XNOR2_X1 U806 ( .A(KEYINPUT1), .B(n1121), .ZN(n1120) );
XNOR2_X1 U807 ( .A(n1122), .B(n1123), .ZN(n1117) );
NAND2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(G69) );
NAND2_X1 U809 ( .A1(n1126), .A2(n1054), .ZN(n1125) );
XNOR2_X1 U810 ( .A(n1127), .B(n1057), .ZN(n1126) );
NAND2_X1 U811 ( .A1(n1128), .A2(G953), .ZN(n1124) );
NAND2_X1 U812 ( .A1(n1129), .A2(n1130), .ZN(n1128) );
NAND2_X1 U813 ( .A1(n1127), .A2(n1131), .ZN(n1130) );
NAND2_X1 U814 ( .A1(G224), .A2(n1132), .ZN(n1129) );
NAND2_X1 U815 ( .A1(G898), .A2(n1127), .ZN(n1132) );
NAND2_X1 U816 ( .A1(n1133), .A2(n1134), .ZN(n1127) );
NAND2_X1 U817 ( .A1(G953), .A2(n1135), .ZN(n1134) );
XOR2_X1 U818 ( .A(n1136), .B(n1137), .Z(n1133) );
NAND2_X1 U819 ( .A1(n1138), .A2(n1139), .ZN(n1136) );
OR2_X1 U820 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U821 ( .A(n1142), .B(KEYINPUT20), .Z(n1138) );
NAND2_X1 U822 ( .A1(n1141), .A2(n1140), .ZN(n1142) );
XOR2_X1 U823 ( .A(n1143), .B(KEYINPUT38), .Z(n1140) );
NOR2_X1 U824 ( .A1(n1144), .A2(n1145), .ZN(G66) );
XOR2_X1 U825 ( .A(n1146), .B(n1147), .Z(n1145) );
NOR2_X1 U826 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
NOR2_X1 U827 ( .A1(n1144), .A2(n1150), .ZN(G63) );
XNOR2_X1 U828 ( .A(n1151), .B(n1152), .ZN(n1150) );
NOR2_X1 U829 ( .A1(n1153), .A2(n1149), .ZN(n1152) );
INV_X1 U830 ( .A(G478), .ZN(n1153) );
NOR2_X1 U831 ( .A1(n1144), .A2(n1154), .ZN(G60) );
XNOR2_X1 U832 ( .A(n1155), .B(n1156), .ZN(n1154) );
NOR2_X1 U833 ( .A1(n1157), .A2(n1149), .ZN(n1156) );
XNOR2_X1 U834 ( .A(G104), .B(n1158), .ZN(G6) );
NOR2_X1 U835 ( .A1(n1144), .A2(n1159), .ZN(G57) );
NOR3_X1 U836 ( .A1(n1160), .A2(n1161), .A3(n1162), .ZN(n1159) );
NOR2_X1 U837 ( .A1(KEYINPUT49), .A2(n1163), .ZN(n1162) );
NOR3_X1 U838 ( .A1(n1164), .A2(n1165), .A3(n1166), .ZN(n1161) );
NOR2_X1 U839 ( .A1(n1167), .A2(n1168), .ZN(n1160) );
NOR2_X1 U840 ( .A1(n1166), .A2(n1169), .ZN(n1167) );
XNOR2_X1 U841 ( .A(KEYINPUT54), .B(n1163), .ZN(n1169) );
INV_X1 U842 ( .A(n1164), .ZN(n1163) );
XNOR2_X1 U843 ( .A(n1170), .B(n1171), .ZN(n1164) );
NOR2_X1 U844 ( .A1(n1172), .A2(n1149), .ZN(n1171) );
NAND2_X1 U845 ( .A1(n1173), .A2(KEYINPUT53), .ZN(n1170) );
XOR2_X1 U846 ( .A(n1174), .B(n1175), .Z(n1173) );
INV_X1 U847 ( .A(KEYINPUT49), .ZN(n1166) );
NOR2_X1 U848 ( .A1(n1144), .A2(n1176), .ZN(G54) );
NOR2_X1 U849 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
XOR2_X1 U850 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U851 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NOR2_X1 U852 ( .A1(n1183), .A2(n1149), .ZN(n1179) );
AND2_X1 U853 ( .A1(n1182), .A2(n1181), .ZN(n1177) );
XNOR2_X1 U854 ( .A(n1184), .B(n1185), .ZN(n1181) );
XNOR2_X1 U855 ( .A(G110), .B(n1186), .ZN(n1185) );
NAND2_X1 U856 ( .A1(KEYINPUT24), .A2(n1187), .ZN(n1186) );
XNOR2_X1 U857 ( .A(n1188), .B(n1189), .ZN(n1184) );
INV_X1 U858 ( .A(KEYINPUT14), .ZN(n1182) );
NOR2_X1 U859 ( .A1(n1144), .A2(n1190), .ZN(G51) );
XOR2_X1 U860 ( .A(n1191), .B(n1192), .Z(n1190) );
XOR2_X1 U861 ( .A(n1193), .B(n1194), .Z(n1192) );
NOR2_X1 U862 ( .A1(KEYINPUT23), .A2(n1195), .ZN(n1194) );
NOR2_X1 U863 ( .A1(n1070), .A2(n1149), .ZN(n1193) );
NAND2_X1 U864 ( .A1(G902), .A2(n1196), .ZN(n1149) );
OR2_X1 U865 ( .A1(n1058), .A2(n1057), .ZN(n1196) );
NAND2_X1 U866 ( .A1(n1197), .A2(n1198), .ZN(n1057) );
NOR4_X1 U867 ( .A1(n1049), .A2(n1199), .A3(n1200), .A4(n1201), .ZN(n1198) );
INV_X1 U868 ( .A(n1202), .ZN(n1201) );
INV_X1 U869 ( .A(n1052), .ZN(n1049) );
NAND3_X1 U870 ( .A1(n1203), .A2(n1204), .A3(n1083), .ZN(n1052) );
AND4_X1 U871 ( .A1(n1205), .A2(n1206), .A3(n1158), .A4(n1207), .ZN(n1197) );
OR2_X1 U872 ( .A1(n1102), .A2(n1208), .ZN(n1207) );
INV_X1 U873 ( .A(n1209), .ZN(n1102) );
NAND3_X1 U874 ( .A1(n1083), .A2(n1204), .A3(n1210), .ZN(n1158) );
NAND3_X1 U875 ( .A1(n1211), .A2(n1212), .A3(n1213), .ZN(n1058) );
AND3_X1 U876 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1213) );
NAND2_X1 U877 ( .A1(n1217), .A2(n1218), .ZN(n1211) );
NAND2_X1 U878 ( .A1(n1219), .A2(n1220), .ZN(n1218) );
NAND4_X1 U879 ( .A1(n1073), .A2(n1098), .A3(n1210), .A4(n1209), .ZN(n1220) );
NAND3_X1 U880 ( .A1(n1221), .A2(n1222), .A3(n1097), .ZN(n1219) );
NAND2_X1 U881 ( .A1(n1082), .A2(n1223), .ZN(n1222) );
NAND3_X1 U882 ( .A1(n1224), .A2(n1225), .A3(n1209), .ZN(n1223) );
NAND2_X1 U883 ( .A1(n1089), .A2(n1226), .ZN(n1082) );
OR2_X1 U884 ( .A1(n1210), .A2(n1203), .ZN(n1226) );
NOR2_X1 U885 ( .A1(n1054), .A2(G952), .ZN(n1144) );
XNOR2_X1 U886 ( .A(G146), .B(n1212), .ZN(G48) );
NAND3_X1 U887 ( .A1(n1227), .A2(n1209), .A3(n1210), .ZN(n1212) );
XNOR2_X1 U888 ( .A(G143), .B(n1228), .ZN(G45) );
NAND4_X1 U889 ( .A1(n1097), .A2(n1221), .A3(n1229), .A4(n1230), .ZN(n1228) );
AND3_X1 U890 ( .A1(n1224), .A2(n1225), .A3(n1217), .ZN(n1230) );
XNOR2_X1 U891 ( .A(n1209), .B(KEYINPUT59), .ZN(n1229) );
XNOR2_X1 U892 ( .A(n1231), .B(n1232), .ZN(G42) );
NOR2_X1 U893 ( .A1(KEYINPUT37), .A2(n1214), .ZN(n1232) );
NAND3_X1 U894 ( .A1(n1233), .A2(n1217), .A3(n1098), .ZN(n1214) );
XOR2_X1 U895 ( .A(n1216), .B(n1234), .Z(G39) );
NAND2_X1 U896 ( .A1(KEYINPUT39), .A2(G137), .ZN(n1234) );
NAND3_X1 U897 ( .A1(n1227), .A2(n1084), .A3(n1089), .ZN(n1216) );
XNOR2_X1 U898 ( .A(G134), .B(n1235), .ZN(G36) );
NAND3_X1 U899 ( .A1(n1236), .A2(n1097), .A3(n1237), .ZN(n1235) );
AND3_X1 U900 ( .A1(n1089), .A2(n1217), .A3(n1203), .ZN(n1237) );
INV_X1 U901 ( .A(n1103), .ZN(n1089) );
XNOR2_X1 U902 ( .A(n1221), .B(KEYINPUT2), .ZN(n1236) );
XNOR2_X1 U903 ( .A(G131), .B(n1238), .ZN(G33) );
NAND3_X1 U904 ( .A1(n1233), .A2(n1239), .A3(n1097), .ZN(n1238) );
XNOR2_X1 U905 ( .A(KEYINPUT56), .B(n1217), .ZN(n1239) );
NOR3_X1 U906 ( .A1(n1103), .A2(n1090), .A3(n1240), .ZN(n1233) );
NAND2_X1 U907 ( .A1(n1104), .A2(n1241), .ZN(n1103) );
XNOR2_X1 U908 ( .A(G128), .B(n1242), .ZN(G30) );
NOR2_X1 U909 ( .A1(n1243), .A2(KEYINPUT19), .ZN(n1242) );
INV_X1 U910 ( .A(n1215), .ZN(n1243) );
NAND3_X1 U911 ( .A1(n1203), .A2(n1209), .A3(n1227), .ZN(n1215) );
AND4_X1 U912 ( .A1(n1221), .A2(n1244), .A3(n1217), .A4(n1245), .ZN(n1227) );
NAND2_X1 U913 ( .A1(n1246), .A2(n1247), .ZN(G3) );
OR2_X1 U914 ( .A1(n1206), .A2(G101), .ZN(n1247) );
XOR2_X1 U915 ( .A(n1248), .B(KEYINPUT63), .Z(n1246) );
NAND2_X1 U916 ( .A1(G101), .A2(n1206), .ZN(n1248) );
NAND3_X1 U917 ( .A1(n1204), .A2(n1084), .A3(n1097), .ZN(n1206) );
AND3_X1 U918 ( .A1(n1221), .A2(n1249), .A3(n1209), .ZN(n1204) );
XNOR2_X1 U919 ( .A(G125), .B(n1250), .ZN(G27) );
NAND4_X1 U920 ( .A1(n1209), .A2(n1217), .A3(n1098), .A4(n1251), .ZN(n1250) );
NOR2_X1 U921 ( .A1(n1081), .A2(n1252), .ZN(n1251) );
XNOR2_X1 U922 ( .A(KEYINPUT18), .B(n1240), .ZN(n1252) );
INV_X1 U923 ( .A(n1073), .ZN(n1081) );
NAND2_X1 U924 ( .A1(n1105), .A2(n1253), .ZN(n1217) );
NAND4_X1 U925 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1255), .ZN(n1253) );
INV_X1 U926 ( .A(G900), .ZN(n1255) );
XOR2_X1 U927 ( .A(n1256), .B(G122), .Z(G24) );
NAND2_X1 U928 ( .A1(KEYINPUT33), .A2(n1205), .ZN(n1256) );
NAND4_X1 U929 ( .A1(n1257), .A2(n1083), .A3(n1224), .A4(n1225), .ZN(n1205) );
NOR2_X1 U930 ( .A1(n1245), .A2(n1244), .ZN(n1083) );
XOR2_X1 U931 ( .A(G119), .B(n1258), .Z(G21) );
NOR2_X1 U932 ( .A1(KEYINPUT43), .A2(n1202), .ZN(n1258) );
NAND4_X1 U933 ( .A1(n1257), .A2(n1084), .A3(n1244), .A4(n1245), .ZN(n1202) );
XNOR2_X1 U934 ( .A(n1259), .B(n1200), .ZN(G18) );
AND3_X1 U935 ( .A1(n1097), .A2(n1203), .A3(n1257), .ZN(n1200) );
NAND2_X1 U936 ( .A1(n1260), .A2(n1261), .ZN(G15) );
NAND2_X1 U937 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NAND2_X1 U938 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
NAND2_X1 U939 ( .A1(KEYINPUT32), .A2(n1266), .ZN(n1265) );
OR2_X1 U940 ( .A1(n1267), .A2(KEYINPUT32), .ZN(n1264) );
NAND2_X1 U941 ( .A1(G113), .A2(n1267), .ZN(n1260) );
NOR2_X1 U942 ( .A1(n1199), .A2(KEYINPUT17), .ZN(n1267) );
INV_X1 U943 ( .A(n1266), .ZN(n1199) );
NAND3_X1 U944 ( .A1(n1097), .A2(n1210), .A3(n1257), .ZN(n1266) );
AND3_X1 U945 ( .A1(n1209), .A2(n1249), .A3(n1073), .ZN(n1257) );
NOR2_X1 U946 ( .A1(n1092), .A2(n1268), .ZN(n1073) );
INV_X1 U947 ( .A(n1075), .ZN(n1268) );
INV_X1 U948 ( .A(n1240), .ZN(n1210) );
NAND2_X1 U949 ( .A1(n1269), .A2(n1224), .ZN(n1240) );
XNOR2_X1 U950 ( .A(KEYINPUT22), .B(n1225), .ZN(n1269) );
NOR2_X1 U951 ( .A1(n1245), .A2(n1270), .ZN(n1097) );
XOR2_X1 U952 ( .A(n1271), .B(n1272), .Z(G12) );
XNOR2_X1 U953 ( .A(KEYINPUT62), .B(n1273), .ZN(n1272) );
NAND2_X1 U954 ( .A1(n1274), .A2(n1209), .ZN(n1271) );
NOR2_X1 U955 ( .A1(n1104), .A2(n1064), .ZN(n1209) );
INV_X1 U956 ( .A(n1241), .ZN(n1064) );
NAND2_X1 U957 ( .A1(G214), .A2(n1275), .ZN(n1241) );
XOR2_X1 U958 ( .A(n1276), .B(n1072), .Z(n1104) );
NAND2_X1 U959 ( .A1(n1277), .A2(n1278), .ZN(n1072) );
XNOR2_X1 U960 ( .A(n1279), .B(n1195), .ZN(n1277) );
XOR2_X1 U961 ( .A(n1280), .B(n1281), .Z(n1195) );
XNOR2_X1 U962 ( .A(G125), .B(G128), .ZN(n1280) );
XNOR2_X1 U963 ( .A(n1191), .B(KEYINPUT42), .ZN(n1279) );
XNOR2_X1 U964 ( .A(n1282), .B(n1283), .ZN(n1191) );
XOR2_X1 U965 ( .A(n1284), .B(n1137), .Z(n1283) );
XNOR2_X1 U966 ( .A(n1273), .B(n1285), .ZN(n1137) );
XOR2_X1 U967 ( .A(KEYINPUT7), .B(G122), .Z(n1285) );
NOR2_X1 U968 ( .A1(G953), .A2(n1131), .ZN(n1284) );
INV_X1 U969 ( .A(G224), .ZN(n1131) );
XNOR2_X1 U970 ( .A(n1141), .B(n1143), .ZN(n1282) );
XNOR2_X1 U971 ( .A(n1286), .B(n1287), .ZN(n1143) );
XNOR2_X1 U972 ( .A(G116), .B(KEYINPUT4), .ZN(n1286) );
AND2_X1 U973 ( .A1(n1288), .A2(n1289), .ZN(n1141) );
NAND2_X1 U974 ( .A1(n1290), .A2(n1050), .ZN(n1289) );
XNOR2_X1 U975 ( .A(n1291), .B(n1292), .ZN(n1290) );
XNOR2_X1 U976 ( .A(KEYINPUT45), .B(KEYINPUT15), .ZN(n1292) );
NAND2_X1 U977 ( .A1(n1291), .A2(G107), .ZN(n1288) );
XOR2_X1 U978 ( .A(n1293), .B(n1294), .Z(n1291) );
INV_X1 U979 ( .A(G104), .ZN(n1294) );
NAND2_X1 U980 ( .A1(KEYINPUT48), .A2(n1295), .ZN(n1293) );
NAND2_X1 U981 ( .A1(KEYINPUT13), .A2(n1070), .ZN(n1276) );
NAND2_X1 U982 ( .A1(G210), .A2(n1275), .ZN(n1070) );
NAND2_X1 U983 ( .A1(n1296), .A2(n1278), .ZN(n1275) );
INV_X1 U984 ( .A(G237), .ZN(n1296) );
XOR2_X1 U985 ( .A(n1208), .B(KEYINPUT44), .Z(n1274) );
NAND4_X1 U986 ( .A1(n1098), .A2(n1221), .A3(n1084), .A4(n1249), .ZN(n1208) );
NAND2_X1 U987 ( .A1(n1105), .A2(n1297), .ZN(n1249) );
NAND4_X1 U988 ( .A1(G953), .A2(G902), .A3(n1254), .A4(n1135), .ZN(n1297) );
INV_X1 U989 ( .A(G898), .ZN(n1135) );
NAND3_X1 U990 ( .A1(n1254), .A2(n1054), .A3(G952), .ZN(n1105) );
NAND2_X1 U991 ( .A1(G237), .A2(G234), .ZN(n1254) );
NAND2_X1 U992 ( .A1(n1298), .A2(n1299), .ZN(n1084) );
OR3_X1 U993 ( .A1(n1225), .A2(n1224), .A3(KEYINPUT22), .ZN(n1299) );
NAND2_X1 U994 ( .A1(KEYINPUT22), .A2(n1203), .ZN(n1298) );
NOR2_X1 U995 ( .A1(n1224), .A2(n1300), .ZN(n1203) );
INV_X1 U996 ( .A(n1225), .ZN(n1300) );
NAND2_X1 U997 ( .A1(n1301), .A2(n1302), .ZN(n1225) );
NAND2_X1 U998 ( .A1(G478), .A2(n1067), .ZN(n1302) );
XNOR2_X1 U999 ( .A(n1063), .B(KEYINPUT57), .ZN(n1301) );
NOR2_X1 U1000 ( .A1(n1067), .A2(G478), .ZN(n1063) );
NAND2_X1 U1001 ( .A1(n1151), .A2(n1278), .ZN(n1067) );
XNOR2_X1 U1002 ( .A(n1303), .B(n1304), .ZN(n1151) );
XOR2_X1 U1003 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1004 ( .A(G134), .B(G107), .ZN(n1306) );
NAND2_X1 U1005 ( .A1(KEYINPUT25), .A2(n1307), .ZN(n1305) );
XNOR2_X1 U1006 ( .A(n1259), .B(n1308), .ZN(n1307) );
XOR2_X1 U1007 ( .A(KEYINPUT10), .B(G122), .Z(n1308) );
XOR2_X1 U1008 ( .A(n1309), .B(n1310), .Z(n1303) );
AND2_X1 U1009 ( .A1(G217), .A2(n1311), .ZN(n1310) );
NAND2_X1 U1010 ( .A1(n1312), .A2(n1313), .ZN(n1309) );
NAND2_X1 U1011 ( .A1(n1314), .A2(n1119), .ZN(n1313) );
XNOR2_X1 U1012 ( .A(n1315), .B(n1316), .ZN(n1314) );
XNOR2_X1 U1013 ( .A(KEYINPUT41), .B(KEYINPUT0), .ZN(n1315) );
NAND2_X1 U1014 ( .A1(n1317), .A2(n1318), .ZN(n1312) );
XNOR2_X1 U1015 ( .A(G128), .B(KEYINPUT5), .ZN(n1318) );
XOR2_X1 U1016 ( .A(n1066), .B(KEYINPUT30), .Z(n1224) );
XOR2_X1 U1017 ( .A(n1319), .B(n1157), .Z(n1066) );
INV_X1 U1018 ( .A(G475), .ZN(n1157) );
NAND2_X1 U1019 ( .A1(n1155), .A2(n1278), .ZN(n1319) );
XNOR2_X1 U1020 ( .A(n1320), .B(n1321), .ZN(n1155) );
XOR2_X1 U1021 ( .A(n1322), .B(n1323), .Z(n1321) );
XNOR2_X1 U1022 ( .A(n1121), .B(G122), .ZN(n1323) );
XNOR2_X1 U1023 ( .A(n1231), .B(G131), .ZN(n1322) );
INV_X1 U1024 ( .A(G140), .ZN(n1231) );
XOR2_X1 U1025 ( .A(n1324), .B(n1325), .Z(n1320) );
XOR2_X1 U1026 ( .A(n1326), .B(n1327), .Z(n1325) );
NAND2_X1 U1027 ( .A1(KEYINPUT50), .A2(n1328), .ZN(n1327) );
NAND2_X1 U1028 ( .A1(G214), .A2(n1329), .ZN(n1326) );
XOR2_X1 U1029 ( .A(n1330), .B(n1331), .Z(n1324) );
NOR2_X1 U1030 ( .A1(G113), .A2(KEYINPUT61), .ZN(n1331) );
INV_X1 U1031 ( .A(n1090), .ZN(n1221) );
NAND2_X1 U1032 ( .A1(n1092), .A2(n1075), .ZN(n1090) );
NAND2_X1 U1033 ( .A1(G221), .A2(n1332), .ZN(n1075) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1278), .ZN(n1332) );
XOR2_X1 U1035 ( .A(n1076), .B(n1183), .Z(n1092) );
INV_X1 U1036 ( .A(G469), .ZN(n1183) );
NAND2_X1 U1037 ( .A1(n1333), .A2(n1278), .ZN(n1076) );
XNOR2_X1 U1038 ( .A(n1334), .B(n1335), .ZN(n1333) );
XOR2_X1 U1039 ( .A(n1188), .B(n1336), .Z(n1335) );
NOR2_X1 U1040 ( .A1(n1337), .A2(n1338), .ZN(n1336) );
XOR2_X1 U1041 ( .A(KEYINPUT11), .B(n1339), .Z(n1338) );
NOR2_X1 U1042 ( .A1(n1340), .A2(n1341), .ZN(n1339) );
AND2_X1 U1043 ( .A1(n1341), .A2(n1340), .ZN(n1337) );
XOR2_X1 U1044 ( .A(n1187), .B(KEYINPUT27), .Z(n1340) );
AND2_X1 U1045 ( .A1(G227), .A2(n1054), .ZN(n1187) );
XNOR2_X1 U1046 ( .A(G140), .B(n1273), .ZN(n1341) );
XOR2_X1 U1047 ( .A(n1342), .B(n1343), .Z(n1188) );
XNOR2_X1 U1048 ( .A(n1295), .B(n1344), .ZN(n1343) );
XNOR2_X1 U1049 ( .A(KEYINPUT1), .B(n1050), .ZN(n1344) );
INV_X1 U1050 ( .A(G107), .ZN(n1050) );
XNOR2_X1 U1051 ( .A(n1330), .B(n1345), .ZN(n1342) );
INV_X1 U1052 ( .A(n1346), .ZN(n1345) );
XNOR2_X1 U1053 ( .A(G104), .B(n1317), .ZN(n1330) );
AND2_X1 U1054 ( .A1(n1270), .A2(n1245), .ZN(n1098) );
NAND3_X1 U1055 ( .A1(n1347), .A2(n1348), .A3(n1349), .ZN(n1245) );
NAND2_X1 U1056 ( .A1(n1350), .A2(n1146), .ZN(n1349) );
OR3_X1 U1057 ( .A1(n1146), .A2(n1350), .A3(G902), .ZN(n1348) );
NOR2_X1 U1058 ( .A1(n1148), .A2(G234), .ZN(n1350) );
INV_X1 U1059 ( .A(G217), .ZN(n1148) );
NAND3_X1 U1060 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1146) );
NAND2_X1 U1061 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
OR3_X1 U1062 ( .A1(n1355), .A2(n1354), .A3(KEYINPUT40), .ZN(n1352) );
XOR2_X1 U1063 ( .A(n1356), .B(G137), .Z(n1354) );
NAND2_X1 U1064 ( .A1(G221), .A2(n1311), .ZN(n1356) );
AND2_X1 U1065 ( .A1(G234), .A2(n1054), .ZN(n1311) );
INV_X1 U1066 ( .A(G953), .ZN(n1054) );
NAND2_X1 U1067 ( .A1(KEYINPUT29), .A2(n1357), .ZN(n1355) );
NAND2_X1 U1068 ( .A1(KEYINPUT40), .A2(n1358), .ZN(n1351) );
INV_X1 U1069 ( .A(n1357), .ZN(n1358) );
XOR2_X1 U1070 ( .A(n1359), .B(n1360), .Z(n1357) );
NOR2_X1 U1071 ( .A1(n1361), .A2(n1362), .ZN(n1360) );
NOR2_X1 U1072 ( .A1(n1363), .A2(n1273), .ZN(n1362) );
INV_X1 U1073 ( .A(G110), .ZN(n1273) );
NOR2_X1 U1074 ( .A1(n1364), .A2(n1365), .ZN(n1361) );
XNOR2_X1 U1075 ( .A(G110), .B(KEYINPUT12), .ZN(n1365) );
INV_X1 U1076 ( .A(n1363), .ZN(n1364) );
NAND2_X1 U1077 ( .A1(n1366), .A2(n1367), .ZN(n1363) );
NAND2_X1 U1078 ( .A1(G119), .A2(n1316), .ZN(n1367) );
XOR2_X1 U1079 ( .A(KEYINPUT46), .B(n1368), .Z(n1366) );
NOR2_X1 U1080 ( .A1(G119), .A2(n1316), .ZN(n1368) );
INV_X1 U1081 ( .A(G128), .ZN(n1316) );
NAND2_X1 U1082 ( .A1(n1369), .A2(KEYINPUT26), .ZN(n1359) );
XNOR2_X1 U1083 ( .A(n1370), .B(n1189), .ZN(n1369) );
INV_X1 U1084 ( .A(n1122), .ZN(n1189) );
XNOR2_X1 U1085 ( .A(G140), .B(n1328), .ZN(n1122) );
INV_X1 U1086 ( .A(n1334), .ZN(n1328) );
NAND2_X1 U1087 ( .A1(KEYINPUT35), .A2(n1121), .ZN(n1370) );
INV_X1 U1088 ( .A(G125), .ZN(n1121) );
NAND2_X1 U1089 ( .A1(G902), .A2(G217), .ZN(n1347) );
INV_X1 U1090 ( .A(n1244), .ZN(n1270) );
XOR2_X1 U1091 ( .A(n1371), .B(n1172), .Z(n1244) );
INV_X1 U1092 ( .A(G472), .ZN(n1172) );
NAND3_X1 U1093 ( .A1(n1372), .A2(n1373), .A3(n1278), .ZN(n1371) );
INV_X1 U1094 ( .A(G902), .ZN(n1278) );
OR3_X1 U1095 ( .A1(n1165), .A2(n1374), .A3(KEYINPUT36), .ZN(n1373) );
NAND2_X1 U1096 ( .A1(n1375), .A2(KEYINPUT36), .ZN(n1372) );
XNOR2_X1 U1097 ( .A(n1374), .B(n1168), .ZN(n1375) );
INV_X1 U1098 ( .A(n1165), .ZN(n1168) );
XOR2_X1 U1099 ( .A(n1376), .B(n1295), .Z(n1165) );
INV_X1 U1100 ( .A(G101), .ZN(n1295) );
NAND2_X1 U1101 ( .A1(G210), .A2(n1329), .ZN(n1376) );
NOR2_X1 U1102 ( .A1(G953), .A2(G237), .ZN(n1329) );
XNOR2_X1 U1103 ( .A(n1174), .B(n1377), .ZN(n1374) );
XOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1378), .Z(n1377) );
NOR2_X1 U1105 ( .A1(KEYINPUT9), .A2(n1175), .ZN(n1378) );
XNOR2_X1 U1106 ( .A(n1379), .B(n1287), .ZN(n1175) );
XNOR2_X1 U1107 ( .A(n1263), .B(G119), .ZN(n1287) );
INV_X1 U1108 ( .A(G113), .ZN(n1263) );
NAND2_X1 U1109 ( .A1(KEYINPUT55), .A2(n1259), .ZN(n1379) );
INV_X1 U1110 ( .A(G116), .ZN(n1259) );
XNOR2_X1 U1111 ( .A(n1346), .B(n1281), .ZN(n1174) );
NOR2_X1 U1112 ( .A1(KEYINPUT6), .A2(n1380), .ZN(n1281) );
XNOR2_X1 U1113 ( .A(n1119), .B(n1381), .ZN(n1380) );
XNOR2_X1 U1114 ( .A(n1382), .B(KEYINPUT60), .ZN(n1381) );
NAND2_X1 U1115 ( .A1(KEYINPUT21), .A2(n1334), .ZN(n1382) );
XOR2_X1 U1116 ( .A(G146), .B(KEYINPUT51), .Z(n1334) );
INV_X1 U1117 ( .A(n1317), .ZN(n1119) );
XOR2_X1 U1118 ( .A(G143), .B(KEYINPUT8), .Z(n1317) );
XOR2_X1 U1119 ( .A(n1123), .B(KEYINPUT47), .Z(n1346) );
XNOR2_X1 U1120 ( .A(n1383), .B(n1384), .ZN(n1123) );
XNOR2_X1 U1121 ( .A(G137), .B(n1385), .ZN(n1384) );
INV_X1 U1122 ( .A(G134), .ZN(n1385) );
XNOR2_X1 U1123 ( .A(G131), .B(G128), .ZN(n1383) );
endmodule


