//Key = 1111010000000011110000101110110110010101100010100001101000010100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;

XOR2_X1 U748 ( .A(n1045), .B(n1046), .Z(G9) );
NAND2_X1 U749 ( .A1(KEYINPUT16), .A2(G107), .ZN(n1046) );
NOR2_X1 U750 ( .A1(n1047), .A2(n1048), .ZN(G75) );
NOR4_X1 U751 ( .A1(G953), .A2(n1049), .A3(n1050), .A4(n1051), .ZN(n1048) );
NOR2_X1 U752 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U753 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
NOR2_X1 U754 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR2_X1 U755 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NOR2_X1 U756 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U757 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR2_X1 U758 ( .A1(n1064), .A2(n1065), .ZN(n1063) );
NOR3_X1 U759 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1064) );
NOR3_X1 U760 ( .A1(n1069), .A2(n1070), .A3(n1071), .ZN(n1068) );
INV_X1 U761 ( .A(KEYINPUT28), .ZN(n1069) );
NOR2_X1 U762 ( .A1(KEYINPUT28), .A2(n1072), .ZN(n1067) );
NOR2_X1 U763 ( .A1(n1073), .A2(n1072), .ZN(n1062) );
NOR2_X1 U764 ( .A1(n1074), .A2(n1075), .ZN(n1073) );
NOR3_X1 U765 ( .A1(n1072), .A2(n1076), .A3(n1065), .ZN(n1058) );
NOR2_X1 U766 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR2_X1 U767 ( .A1(n1079), .A2(n1080), .ZN(n1077) );
NOR4_X1 U768 ( .A1(n1081), .A2(n1065), .A3(n1061), .A4(n1072), .ZN(n1054) );
NOR2_X1 U769 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
NOR3_X1 U770 ( .A1(n1049), .A2(G953), .A3(G952), .ZN(n1047) );
AND4_X1 U771 ( .A1(n1084), .A2(n1085), .A3(n1086), .A4(n1071), .ZN(n1049) );
XNOR2_X1 U772 ( .A(n1087), .B(n1088), .ZN(n1086) );
NAND2_X1 U773 ( .A1(KEYINPUT25), .A2(n1089), .ZN(n1088) );
XOR2_X1 U774 ( .A(KEYINPUT19), .B(n1090), .Z(n1085) );
NOR4_X1 U775 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1090) );
NAND2_X1 U776 ( .A1(n1095), .A2(n1096), .ZN(n1092) );
XOR2_X1 U777 ( .A(n1097), .B(n1098), .Z(G72) );
XOR2_X1 U778 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U779 ( .A1(n1101), .A2(n1102), .ZN(n1100) );
XOR2_X1 U780 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U781 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U782 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
NOR3_X1 U783 ( .A1(KEYINPUT44), .A2(G137), .A3(n1109), .ZN(n1108) );
INV_X1 U784 ( .A(G134), .ZN(n1109) );
NOR2_X1 U785 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
INV_X1 U786 ( .A(KEYINPUT44), .ZN(n1111) );
XOR2_X1 U787 ( .A(n1112), .B(n1113), .Z(n1103) );
XNOR2_X1 U788 ( .A(G131), .B(KEYINPUT17), .ZN(n1113) );
NAND2_X1 U789 ( .A1(n1114), .A2(n1115), .ZN(n1112) );
NAND2_X1 U790 ( .A1(KEYINPUT52), .A2(n1116), .ZN(n1115) );
NAND2_X1 U791 ( .A1(G140), .A2(n1117), .ZN(n1114) );
NAND2_X1 U792 ( .A1(KEYINPUT52), .A2(n1118), .ZN(n1117) );
NOR2_X1 U793 ( .A1(G900), .A2(n1119), .ZN(n1101) );
NAND3_X1 U794 ( .A1(n1120), .A2(n1119), .A3(KEYINPUT29), .ZN(n1099) );
NAND2_X1 U795 ( .A1(G953), .A2(n1121), .ZN(n1097) );
NAND2_X1 U796 ( .A1(G900), .A2(G227), .ZN(n1121) );
NAND2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(G69) );
NAND2_X1 U798 ( .A1(n1124), .A2(n1119), .ZN(n1123) );
XNOR2_X1 U799 ( .A(n1125), .B(n1126), .ZN(n1124) );
NOR2_X1 U800 ( .A1(n1127), .A2(KEYINPUT36), .ZN(n1126) );
NOR2_X1 U801 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U802 ( .A1(n1130), .A2(G953), .ZN(n1122) );
XOR2_X1 U803 ( .A(n1125), .B(n1131), .Z(n1130) );
NOR2_X1 U804 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
NAND2_X1 U805 ( .A1(n1134), .A2(n1135), .ZN(n1125) );
NAND2_X1 U806 ( .A1(G953), .A2(n1133), .ZN(n1135) );
XOR2_X1 U807 ( .A(n1136), .B(n1137), .Z(n1134) );
NOR2_X1 U808 ( .A1(n1138), .A2(n1139), .ZN(G66) );
XOR2_X1 U809 ( .A(n1140), .B(n1141), .Z(n1139) );
NOR2_X1 U810 ( .A1(n1142), .A2(n1143), .ZN(n1140) );
NOR2_X1 U811 ( .A1(n1138), .A2(n1144), .ZN(G63) );
XOR2_X1 U812 ( .A(n1145), .B(n1146), .Z(n1144) );
NOR2_X1 U813 ( .A1(n1147), .A2(n1143), .ZN(n1145) );
INV_X1 U814 ( .A(G478), .ZN(n1147) );
NOR3_X1 U815 ( .A1(n1138), .A2(n1148), .A3(n1149), .ZN(G60) );
NOR4_X1 U816 ( .A1(n1150), .A2(n1151), .A3(n1152), .A4(n1143), .ZN(n1149) );
INV_X1 U817 ( .A(KEYINPUT51), .ZN(n1151) );
NOR2_X1 U818 ( .A1(n1153), .A2(n1154), .ZN(n1148) );
NOR3_X1 U819 ( .A1(n1143), .A2(n1155), .A3(n1152), .ZN(n1154) );
INV_X1 U820 ( .A(G475), .ZN(n1152) );
NOR2_X1 U821 ( .A1(KEYINPUT51), .A2(n1156), .ZN(n1155) );
INV_X1 U822 ( .A(n1150), .ZN(n1153) );
NAND2_X1 U823 ( .A1(KEYINPUT31), .A2(n1156), .ZN(n1150) );
XOR2_X1 U824 ( .A(G104), .B(n1157), .Z(G6) );
NOR2_X1 U825 ( .A1(n1158), .A2(n1159), .ZN(n1157) );
XOR2_X1 U826 ( .A(n1160), .B(KEYINPUT7), .Z(n1158) );
NOR2_X1 U827 ( .A1(n1138), .A2(n1161), .ZN(G57) );
XOR2_X1 U828 ( .A(n1162), .B(n1163), .Z(n1161) );
XOR2_X1 U829 ( .A(n1164), .B(n1165), .Z(n1163) );
NAND3_X1 U830 ( .A1(n1166), .A2(n1167), .A3(n1168), .ZN(n1164) );
XNOR2_X1 U831 ( .A(KEYINPUT50), .B(KEYINPUT12), .ZN(n1168) );
NAND2_X1 U832 ( .A1(n1169), .A2(n1170), .ZN(n1167) );
INV_X1 U833 ( .A(n1171), .ZN(n1170) );
XNOR2_X1 U834 ( .A(n1172), .B(KEYINPUT0), .ZN(n1169) );
NAND2_X1 U835 ( .A1(n1171), .A2(n1173), .ZN(n1166) );
XNOR2_X1 U836 ( .A(n1172), .B(KEYINPUT43), .ZN(n1173) );
XOR2_X1 U837 ( .A(KEYINPUT21), .B(n1174), .Z(n1162) );
NOR2_X1 U838 ( .A1(n1175), .A2(n1143), .ZN(n1174) );
INV_X1 U839 ( .A(G472), .ZN(n1175) );
NOR2_X1 U840 ( .A1(n1138), .A2(n1176), .ZN(G54) );
XOR2_X1 U841 ( .A(n1177), .B(n1178), .Z(n1176) );
XOR2_X1 U842 ( .A(n1179), .B(n1180), .Z(n1178) );
NOR2_X1 U843 ( .A1(n1181), .A2(n1143), .ZN(n1180) );
INV_X1 U844 ( .A(G469), .ZN(n1181) );
NOR2_X1 U845 ( .A1(KEYINPUT57), .A2(n1182), .ZN(n1179) );
XOR2_X1 U846 ( .A(n1183), .B(n1184), .Z(n1177) );
XNOR2_X1 U847 ( .A(KEYINPUT42), .B(n1185), .ZN(n1183) );
NOR2_X1 U848 ( .A1(KEYINPUT6), .A2(n1186), .ZN(n1185) );
XNOR2_X1 U849 ( .A(n1187), .B(n1188), .ZN(n1186) );
NOR2_X1 U850 ( .A1(KEYINPUT13), .A2(n1172), .ZN(n1187) );
NOR2_X1 U851 ( .A1(n1138), .A2(n1189), .ZN(G51) );
NOR3_X1 U852 ( .A1(n1087), .A2(n1190), .A3(n1191), .ZN(n1189) );
NOR4_X1 U853 ( .A1(n1192), .A2(n1143), .A3(KEYINPUT8), .A4(n1089), .ZN(n1191) );
NAND2_X1 U854 ( .A1(G902), .A2(n1051), .ZN(n1143) );
INV_X1 U855 ( .A(n1193), .ZN(n1051) );
NOR2_X1 U856 ( .A1(n1194), .A2(n1195), .ZN(n1190) );
NOR3_X1 U857 ( .A1(n1089), .A2(KEYINPUT8), .A3(n1193), .ZN(n1194) );
NOR3_X1 U858 ( .A1(n1129), .A2(n1196), .A3(n1120), .ZN(n1193) );
NAND4_X1 U859 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1120) );
NOR4_X1 U860 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1200) );
NOR2_X1 U861 ( .A1(n1205), .A2(n1206), .ZN(n1204) );
XOR2_X1 U862 ( .A(n1207), .B(KEYINPUT30), .Z(n1205) );
NOR3_X1 U863 ( .A1(n1208), .A2(n1209), .A3(n1210), .ZN(n1203) );
INV_X1 U864 ( .A(n1211), .ZN(n1201) );
AND2_X1 U865 ( .A1(n1212), .A2(n1213), .ZN(n1199) );
XNOR2_X1 U866 ( .A(KEYINPUT5), .B(n1128), .ZN(n1196) );
NAND4_X1 U867 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1129) );
AND3_X1 U868 ( .A1(n1045), .A2(n1218), .A3(n1219), .ZN(n1217) );
NAND4_X1 U869 ( .A1(n1220), .A2(n1082), .A3(n1221), .A4(n1222), .ZN(n1045) );
OR2_X1 U870 ( .A1(n1160), .A2(n1159), .ZN(n1216) );
NAND4_X1 U871 ( .A1(n1083), .A2(n1221), .A3(n1078), .A4(n1222), .ZN(n1160) );
NAND2_X1 U872 ( .A1(n1223), .A2(n1074), .ZN(n1215) );
NAND2_X1 U873 ( .A1(n1224), .A2(n1225), .ZN(n1214) );
NAND2_X1 U874 ( .A1(n1226), .A2(n1227), .ZN(n1225) );
NAND2_X1 U875 ( .A1(n1221), .A2(n1228), .ZN(n1227) );
NAND2_X1 U876 ( .A1(n1075), .A2(n1083), .ZN(n1226) );
NOR2_X1 U877 ( .A1(n1119), .A2(G952), .ZN(n1138) );
XOR2_X1 U878 ( .A(G146), .B(n1229), .Z(G48) );
NOR2_X1 U879 ( .A1(n1206), .A2(n1207), .ZN(n1229) );
INV_X1 U880 ( .A(n1083), .ZN(n1207) );
XNOR2_X1 U881 ( .A(n1202), .B(n1230), .ZN(G45) );
NAND2_X1 U882 ( .A1(n1231), .A2(KEYINPUT35), .ZN(n1230) );
XOR2_X1 U883 ( .A(n1232), .B(KEYINPUT59), .Z(n1231) );
AND4_X1 U884 ( .A1(n1075), .A2(n1220), .A3(n1228), .A4(n1233), .ZN(n1202) );
XOR2_X1 U885 ( .A(n1234), .B(n1211), .Z(G42) );
NAND2_X1 U886 ( .A1(n1235), .A2(n1236), .ZN(n1211) );
XNOR2_X1 U887 ( .A(G137), .B(n1213), .ZN(G39) );
NAND4_X1 U888 ( .A1(n1237), .A2(n1235), .A3(n1093), .A4(n1238), .ZN(n1213) );
XOR2_X1 U889 ( .A(G134), .B(n1239), .Z(G36) );
NOR4_X1 U890 ( .A1(n1209), .A2(n1240), .A3(n1072), .A4(n1210), .ZN(n1239) );
NAND2_X1 U891 ( .A1(n1241), .A2(n1233), .ZN(n1240) );
XOR2_X1 U892 ( .A(KEYINPUT49), .B(n1078), .Z(n1241) );
NAND2_X1 U893 ( .A1(n1242), .A2(n1243), .ZN(G33) );
NAND2_X1 U894 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
INV_X1 U895 ( .A(n1212), .ZN(n1245) );
XNOR2_X1 U896 ( .A(G131), .B(KEYINPUT34), .ZN(n1244) );
NAND2_X1 U897 ( .A1(n1246), .A2(n1247), .ZN(n1242) );
XOR2_X1 U898 ( .A(n1212), .B(KEYINPUT41), .Z(n1247) );
NAND3_X1 U899 ( .A1(n1075), .A2(n1083), .A3(n1235), .ZN(n1212) );
INV_X1 U900 ( .A(n1208), .ZN(n1235) );
NAND3_X1 U901 ( .A1(n1078), .A2(n1233), .A3(n1248), .ZN(n1208) );
INV_X1 U902 ( .A(n1072), .ZN(n1248) );
NAND2_X1 U903 ( .A1(n1249), .A2(n1071), .ZN(n1072) );
INV_X1 U904 ( .A(n1070), .ZN(n1249) );
XNOR2_X1 U905 ( .A(G131), .B(KEYINPUT24), .ZN(n1246) );
XNOR2_X1 U906 ( .A(n1250), .B(n1198), .ZN(G30) );
OR2_X1 U907 ( .A1(n1206), .A2(n1209), .ZN(n1198) );
NAND4_X1 U908 ( .A1(n1220), .A2(n1093), .A3(n1233), .A4(n1238), .ZN(n1206) );
XOR2_X1 U909 ( .A(n1251), .B(KEYINPUT1), .Z(n1250) );
XOR2_X1 U910 ( .A(n1219), .B(n1252), .Z(G3) );
XOR2_X1 U911 ( .A(KEYINPUT54), .B(G101), .Z(n1252) );
NAND2_X1 U912 ( .A1(n1223), .A2(n1075), .ZN(n1219) );
XOR2_X1 U913 ( .A(n1118), .B(n1197), .Z(G27) );
NAND4_X1 U914 ( .A1(n1236), .A2(n1084), .A3(n1066), .A4(n1233), .ZN(n1197) );
NAND2_X1 U915 ( .A1(n1253), .A2(n1254), .ZN(n1233) );
NAND4_X1 U916 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1256), .ZN(n1254) );
INV_X1 U917 ( .A(G900), .ZN(n1256) );
XNOR2_X1 U918 ( .A(KEYINPUT32), .B(n1053), .ZN(n1253) );
AND2_X1 U919 ( .A1(n1083), .A2(n1074), .ZN(n1236) );
XNOR2_X1 U920 ( .A(G122), .B(n1257), .ZN(G24) );
NAND3_X1 U921 ( .A1(n1224), .A2(n1221), .A3(n1258), .ZN(n1257) );
XNOR2_X1 U922 ( .A(KEYINPUT22), .B(n1228), .ZN(n1258) );
NAND2_X1 U923 ( .A1(n1259), .A2(n1260), .ZN(n1228) );
OR3_X1 U924 ( .A1(n1261), .A2(n1262), .A3(KEYINPUT60), .ZN(n1260) );
NAND2_X1 U925 ( .A1(KEYINPUT60), .A2(n1083), .ZN(n1259) );
INV_X1 U926 ( .A(n1065), .ZN(n1221) );
NAND2_X1 U927 ( .A1(n1263), .A2(n1264), .ZN(n1065) );
XNOR2_X1 U928 ( .A(n1128), .B(n1265), .ZN(G21) );
NOR2_X1 U929 ( .A1(G119), .A2(KEYINPUT9), .ZN(n1265) );
AND4_X1 U930 ( .A1(n1224), .A2(n1237), .A3(n1093), .A4(n1238), .ZN(n1128) );
XNOR2_X1 U931 ( .A(G116), .B(n1218), .ZN(G18) );
NAND3_X1 U932 ( .A1(n1075), .A2(n1082), .A3(n1224), .ZN(n1218) );
INV_X1 U933 ( .A(n1209), .ZN(n1082) );
NAND2_X1 U934 ( .A1(n1262), .A2(n1266), .ZN(n1209) );
XOR2_X1 U935 ( .A(KEYINPUT20), .B(n1094), .Z(n1266) );
INV_X1 U936 ( .A(n1210), .ZN(n1075) );
XOR2_X1 U937 ( .A(n1267), .B(G113), .Z(G15) );
NAND2_X1 U938 ( .A1(n1268), .A2(n1269), .ZN(n1267) );
NAND4_X1 U939 ( .A1(n1270), .A2(n1083), .A3(n1224), .A4(n1271), .ZN(n1269) );
INV_X1 U940 ( .A(KEYINPUT23), .ZN(n1271) );
AND3_X1 U941 ( .A1(n1066), .A2(n1222), .A3(n1084), .ZN(n1224) );
NAND3_X1 U942 ( .A1(n1066), .A2(n1272), .A3(KEYINPUT23), .ZN(n1268) );
NAND4_X1 U943 ( .A1(n1270), .A2(n1083), .A3(n1084), .A4(n1222), .ZN(n1272) );
INV_X1 U944 ( .A(n1061), .ZN(n1084) );
NAND2_X1 U945 ( .A1(n1273), .A2(n1080), .ZN(n1061) );
INV_X1 U946 ( .A(n1079), .ZN(n1273) );
NOR2_X1 U947 ( .A1(n1094), .A2(n1262), .ZN(n1083) );
XOR2_X1 U948 ( .A(n1210), .B(KEYINPUT15), .Z(n1270) );
NAND2_X1 U949 ( .A1(n1264), .A2(n1238), .ZN(n1210) );
XNOR2_X1 U950 ( .A(n1093), .B(KEYINPUT27), .ZN(n1264) );
XOR2_X1 U951 ( .A(n1274), .B(n1275), .Z(G12) );
NAND3_X1 U952 ( .A1(n1223), .A2(n1074), .A3(KEYINPUT61), .ZN(n1275) );
AND2_X1 U953 ( .A1(n1263), .A2(n1093), .ZN(n1074) );
XOR2_X1 U954 ( .A(n1276), .B(n1142), .Z(n1093) );
NAND2_X1 U955 ( .A1(G217), .A2(n1277), .ZN(n1142) );
OR2_X1 U956 ( .A1(n1141), .A2(G902), .ZN(n1276) );
XNOR2_X1 U957 ( .A(n1278), .B(n1279), .ZN(n1141) );
XOR2_X1 U958 ( .A(G137), .B(n1280), .Z(n1279) );
NOR2_X1 U959 ( .A1(KEYINPUT56), .A2(n1281), .ZN(n1280) );
XOR2_X1 U960 ( .A(n1282), .B(n1283), .Z(n1281) );
XOR2_X1 U961 ( .A(n1284), .B(n1285), .Z(n1283) );
NAND2_X1 U962 ( .A1(n1286), .A2(n1287), .ZN(n1284) );
NAND2_X1 U963 ( .A1(G125), .A2(n1288), .ZN(n1287) );
NAND2_X1 U964 ( .A1(KEYINPUT2), .A2(n1234), .ZN(n1288) );
NAND2_X1 U965 ( .A1(KEYINPUT2), .A2(n1116), .ZN(n1286) );
XOR2_X1 U966 ( .A(G119), .B(G110), .Z(n1282) );
NAND3_X1 U967 ( .A1(G234), .A2(n1119), .A3(G221), .ZN(n1278) );
INV_X1 U968 ( .A(n1238), .ZN(n1263) );
NAND2_X1 U969 ( .A1(n1289), .A2(n1095), .ZN(n1238) );
NAND2_X1 U970 ( .A1(G472), .A2(n1290), .ZN(n1095) );
XOR2_X1 U971 ( .A(n1096), .B(KEYINPUT38), .Z(n1289) );
OR2_X1 U972 ( .A1(n1290), .A2(G472), .ZN(n1096) );
NAND2_X1 U973 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U974 ( .A(n1171), .B(n1293), .Z(n1291) );
XNOR2_X1 U975 ( .A(n1172), .B(n1165), .ZN(n1293) );
XOR2_X1 U976 ( .A(n1294), .B(n1295), .Z(n1165) );
XOR2_X1 U977 ( .A(n1296), .B(n1297), .Z(n1295) );
NAND3_X1 U978 ( .A1(n1298), .A2(n1119), .A3(G210), .ZN(n1297) );
NAND2_X1 U979 ( .A1(n1299), .A2(n1300), .ZN(n1294) );
NAND2_X1 U980 ( .A1(G113), .A2(n1301), .ZN(n1300) );
XOR2_X1 U981 ( .A(n1302), .B(KEYINPUT10), .Z(n1299) );
OR2_X1 U982 ( .A1(n1301), .A2(G113), .ZN(n1302) );
AND3_X1 U983 ( .A1(n1220), .A2(n1222), .A3(n1237), .ZN(n1223) );
INV_X1 U984 ( .A(n1057), .ZN(n1237) );
NAND2_X1 U985 ( .A1(n1262), .A2(n1303), .ZN(n1057) );
XOR2_X1 U986 ( .A(KEYINPUT46), .B(n1094), .Z(n1303) );
INV_X1 U987 ( .A(n1261), .ZN(n1094) );
XOR2_X1 U988 ( .A(n1304), .B(G478), .Z(n1261) );
OR2_X1 U989 ( .A1(n1146), .A2(G902), .ZN(n1304) );
XNOR2_X1 U990 ( .A(n1305), .B(n1306), .ZN(n1146) );
XOR2_X1 U991 ( .A(G128), .B(n1307), .Z(n1306) );
XOR2_X1 U992 ( .A(G143), .B(G134), .Z(n1307) );
XOR2_X1 U993 ( .A(n1308), .B(n1309), .Z(n1305) );
XOR2_X1 U994 ( .A(G107), .B(n1310), .Z(n1309) );
NOR2_X1 U995 ( .A1(KEYINPUT63), .A2(n1311), .ZN(n1310) );
XNOR2_X1 U996 ( .A(G116), .B(n1312), .ZN(n1311) );
NOR2_X1 U997 ( .A1(KEYINPUT48), .A2(n1313), .ZN(n1312) );
NAND3_X1 U998 ( .A1(G217), .A2(G234), .A3(n1314), .ZN(n1308) );
XOR2_X1 U999 ( .A(n1119), .B(KEYINPUT18), .Z(n1314) );
XNOR2_X1 U1000 ( .A(n1091), .B(KEYINPUT47), .ZN(n1262) );
XNOR2_X1 U1001 ( .A(n1315), .B(G475), .ZN(n1091) );
NAND2_X1 U1002 ( .A1(n1156), .A2(n1292), .ZN(n1315) );
XNOR2_X1 U1003 ( .A(n1316), .B(n1317), .ZN(n1156) );
XOR2_X1 U1004 ( .A(n1318), .B(n1319), .Z(n1317) );
XOR2_X1 U1005 ( .A(n1320), .B(n1321), .Z(n1319) );
NAND2_X1 U1006 ( .A1(n1322), .A2(n1323), .ZN(n1321) );
OR2_X1 U1007 ( .A1(n1324), .A2(G104), .ZN(n1323) );
XOR2_X1 U1008 ( .A(n1325), .B(KEYINPUT55), .Z(n1322) );
NAND2_X1 U1009 ( .A1(G104), .A2(n1324), .ZN(n1325) );
NAND2_X1 U1010 ( .A1(n1326), .A2(n1327), .ZN(n1324) );
OR2_X1 U1011 ( .A1(n1328), .A2(G113), .ZN(n1327) );
XOR2_X1 U1012 ( .A(n1329), .B(KEYINPUT62), .Z(n1326) );
NAND2_X1 U1013 ( .A1(n1328), .A2(G113), .ZN(n1329) );
NAND3_X1 U1014 ( .A1(n1298), .A2(n1119), .A3(G214), .ZN(n1320) );
XOR2_X1 U1015 ( .A(G237), .B(KEYINPUT40), .Z(n1298) );
NOR2_X1 U1016 ( .A1(n1330), .A2(n1331), .ZN(n1318) );
AND2_X1 U1017 ( .A1(KEYINPUT14), .A2(n1116), .ZN(n1331) );
NOR2_X1 U1018 ( .A1(G125), .A2(G140), .ZN(n1116) );
NOR2_X1 U1019 ( .A1(n1332), .A2(n1118), .ZN(n1330) );
INV_X1 U1020 ( .A(G125), .ZN(n1118) );
AND2_X1 U1021 ( .A1(n1234), .A2(KEYINPUT14), .ZN(n1332) );
INV_X1 U1022 ( .A(G140), .ZN(n1234) );
XNOR2_X1 U1023 ( .A(G131), .B(n1333), .ZN(n1316) );
XOR2_X1 U1024 ( .A(G146), .B(G143), .Z(n1333) );
NAND2_X1 U1025 ( .A1(n1053), .A2(n1334), .ZN(n1222) );
NAND4_X1 U1026 ( .A1(G953), .A2(G902), .A3(n1255), .A4(n1133), .ZN(n1334) );
INV_X1 U1027 ( .A(G898), .ZN(n1133) );
NAND3_X1 U1028 ( .A1(n1255), .A2(n1119), .A3(G952), .ZN(n1053) );
NAND2_X1 U1029 ( .A1(G237), .A2(G234), .ZN(n1255) );
AND2_X1 U1030 ( .A1(n1066), .A2(n1078), .ZN(n1220) );
AND2_X1 U1031 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
NAND2_X1 U1032 ( .A1(G221), .A2(n1277), .ZN(n1080) );
NAND2_X1 U1033 ( .A1(G234), .A2(n1292), .ZN(n1277) );
XNOR2_X1 U1034 ( .A(n1335), .B(G469), .ZN(n1079) );
NAND2_X1 U1035 ( .A1(n1336), .A2(n1292), .ZN(n1335) );
XOR2_X1 U1036 ( .A(n1337), .B(n1338), .Z(n1336) );
XNOR2_X1 U1037 ( .A(n1339), .B(n1340), .ZN(n1338) );
NOR2_X1 U1038 ( .A1(KEYINPUT11), .A2(n1188), .ZN(n1340) );
XNOR2_X1 U1039 ( .A(n1341), .B(n1342), .ZN(n1188) );
XOR2_X1 U1040 ( .A(n1296), .B(n1105), .Z(n1341) );
XOR2_X1 U1041 ( .A(n1343), .B(n1344), .Z(n1105) );
NOR2_X1 U1042 ( .A1(G143), .A2(KEYINPUT45), .ZN(n1344) );
NAND2_X1 U1043 ( .A1(KEYINPUT3), .A2(n1184), .ZN(n1339) );
AND2_X1 U1044 ( .A1(G227), .A2(n1119), .ZN(n1184) );
INV_X1 U1045 ( .A(G953), .ZN(n1119) );
XNOR2_X1 U1046 ( .A(n1172), .B(n1182), .ZN(n1337) );
XOR2_X1 U1047 ( .A(G110), .B(G140), .Z(n1182) );
XOR2_X1 U1048 ( .A(G131), .B(n1110), .Z(n1172) );
XOR2_X1 U1049 ( .A(G134), .B(G137), .Z(n1110) );
INV_X1 U1050 ( .A(n1159), .ZN(n1066) );
NAND2_X1 U1051 ( .A1(n1070), .A2(n1071), .ZN(n1159) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1345), .ZN(n1071) );
NAND2_X1 U1053 ( .A1(n1346), .A2(n1347), .ZN(n1070) );
NAND2_X1 U1054 ( .A1(n1087), .A2(n1089), .ZN(n1347) );
XOR2_X1 U1055 ( .A(KEYINPUT37), .B(n1348), .Z(n1346) );
NOR2_X1 U1056 ( .A1(n1087), .A2(n1089), .ZN(n1348) );
NAND2_X1 U1057 ( .A1(G210), .A2(n1345), .ZN(n1089) );
NAND2_X1 U1058 ( .A1(n1349), .A2(n1292), .ZN(n1345) );
INV_X1 U1059 ( .A(G902), .ZN(n1292) );
INV_X1 U1060 ( .A(G237), .ZN(n1349) );
NOR2_X1 U1061 ( .A1(n1195), .A2(G902), .ZN(n1087) );
INV_X1 U1062 ( .A(n1192), .ZN(n1195) );
XOR2_X1 U1063 ( .A(n1350), .B(n1351), .Z(n1192) );
XOR2_X1 U1064 ( .A(n1352), .B(n1353), .Z(n1351) );
XOR2_X1 U1065 ( .A(G125), .B(n1354), .Z(n1353) );
NOR2_X1 U1066 ( .A1(KEYINPUT53), .A2(n1136), .ZN(n1354) );
NAND3_X1 U1067 ( .A1(n1355), .A2(n1356), .A3(n1357), .ZN(n1136) );
NAND2_X1 U1068 ( .A1(KEYINPUT58), .A2(n1296), .ZN(n1357) );
OR3_X1 U1069 ( .A1(n1296), .A2(KEYINPUT58), .A3(n1342), .ZN(n1356) );
NAND2_X1 U1070 ( .A1(n1342), .A2(n1358), .ZN(n1355) );
NAND2_X1 U1071 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
INV_X1 U1072 ( .A(KEYINPUT58), .ZN(n1360) );
XOR2_X1 U1073 ( .A(n1296), .B(KEYINPUT39), .Z(n1359) );
INV_X1 U1074 ( .A(G101), .ZN(n1296) );
XNOR2_X1 U1075 ( .A(G107), .B(G104), .ZN(n1342) );
NOR2_X1 U1076 ( .A1(G953), .A2(n1132), .ZN(n1352) );
INV_X1 U1077 ( .A(G224), .ZN(n1132) );
XOR2_X1 U1078 ( .A(n1137), .B(n1171), .Z(n1350) );
XNOR2_X1 U1079 ( .A(n1232), .B(n1343), .ZN(n1171) );
INV_X1 U1080 ( .A(n1285), .ZN(n1343) );
XOR2_X1 U1081 ( .A(n1251), .B(G146), .Z(n1285) );
INV_X1 U1082 ( .A(G128), .ZN(n1251) );
INV_X1 U1083 ( .A(G143), .ZN(n1232) );
XOR2_X1 U1084 ( .A(n1361), .B(n1362), .Z(n1137) );
XNOR2_X1 U1085 ( .A(G113), .B(n1363), .ZN(n1362) );
XNOR2_X1 U1086 ( .A(KEYINPUT4), .B(KEYINPUT26), .ZN(n1363) );
XOR2_X1 U1087 ( .A(n1364), .B(n1313), .Z(n1361) );
INV_X1 U1088 ( .A(n1328), .ZN(n1313) );
XNOR2_X1 U1089 ( .A(G122), .B(KEYINPUT33), .ZN(n1328) );
XOR2_X1 U1090 ( .A(n1274), .B(n1301), .Z(n1364) );
XOR2_X1 U1091 ( .A(G116), .B(G119), .Z(n1301) );
INV_X1 U1092 ( .A(G110), .ZN(n1274) );
endmodule


