//Key = 0011111010100111101100111110110001011100011001111110101110111111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
n1353, n1354, n1355, n1356, n1357, n1358;

NAND2_X1 U743 ( .A1(n1033), .A2(n1034), .ZN(G9) );
NAND2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
XOR2_X1 U745 ( .A(KEYINPUT29), .B(n1037), .Z(n1033) );
NOR2_X1 U746 ( .A1(n1035), .A2(n1036), .ZN(n1037) );
AND3_X1 U747 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1035) );
XNOR2_X1 U748 ( .A(n1041), .B(KEYINPUT59), .ZN(n1040) );
NOR2_X1 U749 ( .A1(n1042), .A2(n1043), .ZN(G75) );
NOR3_X1 U750 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND3_X1 U751 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1044) );
NAND2_X1 U752 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NAND2_X1 U753 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND3_X1 U754 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1053) );
NAND2_X1 U755 ( .A1(n1057), .A2(n1058), .ZN(n1055) );
NAND2_X1 U756 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
OR2_X1 U757 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND2_X1 U758 ( .A1(n1063), .A2(n1064), .ZN(n1057) );
NAND2_X1 U759 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NAND2_X1 U760 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND3_X1 U761 ( .A1(n1063), .A2(n1069), .A3(n1059), .ZN(n1052) );
NAND3_X1 U762 ( .A1(n1070), .A2(n1071), .A3(n1072), .ZN(n1069) );
NAND2_X1 U763 ( .A1(n1054), .A2(n1073), .ZN(n1072) );
OR2_X1 U764 ( .A1(n1038), .A2(n1074), .ZN(n1073) );
NAND3_X1 U765 ( .A1(n1056), .A2(n1075), .A3(n1076), .ZN(n1070) );
NOR3_X1 U766 ( .A1(n1077), .A2(G953), .A3(G952), .ZN(n1042) );
INV_X1 U767 ( .A(n1047), .ZN(n1077) );
NAND4_X1 U768 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1047) );
NOR4_X1 U769 ( .A1(n1082), .A2(n1083), .A3(n1067), .A4(n1084), .ZN(n1081) );
INV_X1 U770 ( .A(n1085), .ZN(n1084) );
NAND2_X1 U771 ( .A1(n1086), .A2(n1087), .ZN(n1082) );
NAND2_X1 U772 ( .A1(n1088), .A2(n1089), .ZN(n1086) );
XNOR2_X1 U773 ( .A(KEYINPUT31), .B(n1090), .ZN(n1088) );
NOR3_X1 U774 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(n1080) );
XNOR2_X1 U775 ( .A(n1094), .B(n1095), .ZN(n1092) );
NOR2_X1 U776 ( .A1(G475), .A2(KEYINPUT30), .ZN(n1095) );
XOR2_X1 U777 ( .A(n1096), .B(KEYINPUT11), .Z(n1078) );
XOR2_X1 U778 ( .A(n1097), .B(n1098), .Z(G72) );
NAND2_X1 U779 ( .A1(G953), .A2(n1099), .ZN(n1098) );
NAND2_X1 U780 ( .A1(G900), .A2(G227), .ZN(n1099) );
NAND3_X1 U781 ( .A1(n1100), .A2(n1101), .A3(KEYINPUT2), .ZN(n1097) );
NAND2_X1 U782 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
NAND2_X1 U783 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NAND2_X1 U784 ( .A1(G953), .A2(n1106), .ZN(n1105) );
XNOR2_X1 U785 ( .A(n1107), .B(n1108), .ZN(n1104) );
NAND2_X1 U786 ( .A1(n1109), .A2(n1045), .ZN(n1100) );
NAND2_X1 U787 ( .A1(n1110), .A2(n1048), .ZN(n1109) );
XNOR2_X1 U788 ( .A(n1107), .B(n1111), .ZN(n1110) );
NAND2_X1 U789 ( .A1(KEYINPUT49), .A2(n1112), .ZN(n1107) );
XOR2_X1 U790 ( .A(n1113), .B(n1114), .Z(n1112) );
NAND2_X1 U791 ( .A1(KEYINPUT55), .A2(n1115), .ZN(n1113) );
XOR2_X1 U792 ( .A(n1116), .B(n1117), .Z(n1115) );
XOR2_X1 U793 ( .A(G137), .B(G131), .Z(n1117) );
NOR2_X1 U794 ( .A1(G134), .A2(KEYINPUT20), .ZN(n1116) );
XOR2_X1 U795 ( .A(n1118), .B(n1119), .Z(G69) );
XOR2_X1 U796 ( .A(n1120), .B(n1121), .Z(n1119) );
NOR2_X1 U797 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
XNOR2_X1 U798 ( .A(G953), .B(KEYINPUT35), .ZN(n1123) );
NAND3_X1 U799 ( .A1(n1124), .A2(n1125), .A3(KEYINPUT5), .ZN(n1120) );
NAND2_X1 U800 ( .A1(G953), .A2(n1126), .ZN(n1125) );
XOR2_X1 U801 ( .A(n1127), .B(n1128), .Z(n1124) );
XOR2_X1 U802 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U803 ( .A(n1131), .B(n1132), .Z(n1127) );
NOR2_X1 U804 ( .A1(KEYINPUT38), .A2(n1133), .ZN(n1132) );
XNOR2_X1 U805 ( .A(KEYINPUT54), .B(KEYINPUT23), .ZN(n1131) );
NAND2_X1 U806 ( .A1(G953), .A2(n1134), .ZN(n1118) );
NAND2_X1 U807 ( .A1(G898), .A2(G224), .ZN(n1134) );
NOR2_X1 U808 ( .A1(n1135), .A2(n1136), .ZN(G66) );
XNOR2_X1 U809 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U810 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NOR2_X1 U811 ( .A1(n1135), .A2(n1141), .ZN(G63) );
XNOR2_X1 U812 ( .A(n1142), .B(n1143), .ZN(n1141) );
NOR3_X1 U813 ( .A1(n1140), .A2(KEYINPUT17), .A3(n1144), .ZN(n1142) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1145), .ZN(G60) );
NOR3_X1 U815 ( .A1(n1094), .A2(n1146), .A3(n1147), .ZN(n1145) );
NOR4_X1 U816 ( .A1(n1148), .A2(n1140), .A3(KEYINPUT0), .A4(n1149), .ZN(n1147) );
INV_X1 U817 ( .A(n1150), .ZN(n1148) );
NOR2_X1 U818 ( .A1(n1151), .A2(n1150), .ZN(n1146) );
NOR3_X1 U819 ( .A1(n1149), .A2(KEYINPUT0), .A3(n1152), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1045), .A2(n1046), .ZN(n1152) );
XOR2_X1 U821 ( .A(n1153), .B(n1154), .Z(G6) );
NAND2_X1 U822 ( .A1(KEYINPUT36), .A2(G104), .ZN(n1154) );
NOR2_X1 U823 ( .A1(n1135), .A2(n1155), .ZN(G57) );
XOR2_X1 U824 ( .A(n1156), .B(n1157), .Z(n1155) );
XOR2_X1 U825 ( .A(n1158), .B(n1159), .Z(n1157) );
NOR2_X1 U826 ( .A1(n1160), .A2(n1140), .ZN(n1158) );
XOR2_X1 U827 ( .A(KEYINPUT47), .B(n1161), .Z(n1156) );
NOR3_X1 U828 ( .A1(n1162), .A2(n1163), .A3(n1164), .ZN(n1161) );
NOR3_X1 U829 ( .A1(n1165), .A2(n1166), .A3(n1167), .ZN(n1162) );
NOR2_X1 U830 ( .A1(n1135), .A2(n1168), .ZN(G54) );
XOR2_X1 U831 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U832 ( .A(n1171), .B(n1172), .Z(n1169) );
NOR2_X1 U833 ( .A1(n1090), .A2(n1140), .ZN(n1172) );
INV_X1 U834 ( .A(G469), .ZN(n1090) );
NAND2_X1 U835 ( .A1(n1173), .A2(n1174), .ZN(n1171) );
NAND2_X1 U836 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
XOR2_X1 U837 ( .A(KEYINPUT18), .B(n1177), .Z(n1173) );
NOR2_X1 U838 ( .A1(n1175), .A2(n1176), .ZN(n1177) );
XNOR2_X1 U839 ( .A(n1114), .B(n1178), .ZN(n1176) );
NOR2_X1 U840 ( .A1(n1135), .A2(n1179), .ZN(G51) );
XOR2_X1 U841 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U842 ( .A1(n1182), .A2(n1140), .ZN(n1181) );
NAND2_X1 U843 ( .A1(G902), .A2(n1183), .ZN(n1140) );
NAND2_X1 U844 ( .A1(n1122), .A2(n1102), .ZN(n1183) );
INV_X1 U845 ( .A(n1045), .ZN(n1102) );
NAND2_X1 U846 ( .A1(n1184), .A2(n1185), .ZN(n1045) );
AND4_X1 U847 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1185) );
AND4_X1 U848 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1184) );
OR2_X1 U849 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
INV_X1 U850 ( .A(n1046), .ZN(n1122) );
NAND4_X1 U851 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1046) );
AND3_X1 U852 ( .A1(n1200), .A2(n1153), .A3(n1201), .ZN(n1199) );
NAND3_X1 U853 ( .A1(n1039), .A2(n1041), .A3(n1074), .ZN(n1153) );
NAND2_X1 U854 ( .A1(n1202), .A2(n1203), .ZN(n1198) );
NAND2_X1 U855 ( .A1(n1041), .A2(n1204), .ZN(n1196) );
NAND3_X1 U856 ( .A1(n1205), .A2(n1206), .A3(n1207), .ZN(n1204) );
XOR2_X1 U857 ( .A(n1208), .B(KEYINPUT43), .Z(n1207) );
NAND3_X1 U858 ( .A1(n1209), .A2(n1210), .A3(n1061), .ZN(n1206) );
NAND2_X1 U859 ( .A1(n1038), .A2(n1039), .ZN(n1205) );
AND3_X1 U860 ( .A1(n1063), .A2(n1210), .A3(n1211), .ZN(n1039) );
NOR2_X1 U861 ( .A1(n1212), .A2(n1213), .ZN(n1180) );
XOR2_X1 U862 ( .A(n1214), .B(KEYINPUT22), .Z(n1213) );
NAND2_X1 U863 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
NOR2_X1 U864 ( .A1(n1215), .A2(n1216), .ZN(n1212) );
XOR2_X1 U865 ( .A(n1217), .B(n1218), .Z(n1215) );
XNOR2_X1 U866 ( .A(n1219), .B(n1220), .ZN(n1218) );
XNOR2_X1 U867 ( .A(G125), .B(KEYINPUT41), .ZN(n1217) );
NOR2_X1 U868 ( .A1(n1048), .A2(G952), .ZN(n1135) );
NAND2_X1 U869 ( .A1(n1221), .A2(n1222), .ZN(G48) );
NAND2_X1 U870 ( .A1(G146), .A2(n1192), .ZN(n1222) );
XOR2_X1 U871 ( .A(KEYINPUT58), .B(n1223), .Z(n1221) );
NOR2_X1 U872 ( .A1(G146), .A2(n1192), .ZN(n1223) );
NAND2_X1 U873 ( .A1(n1224), .A2(n1074), .ZN(n1192) );
XNOR2_X1 U874 ( .A(G143), .B(n1191), .ZN(G45) );
NAND3_X1 U875 ( .A1(n1225), .A2(n1062), .A3(n1226), .ZN(n1191) );
NOR3_X1 U876 ( .A1(n1065), .A2(n1227), .A3(n1228), .ZN(n1226) );
XNOR2_X1 U877 ( .A(G140), .B(n1190), .ZN(G42) );
NAND2_X1 U878 ( .A1(n1229), .A2(n1061), .ZN(n1190) );
XOR2_X1 U879 ( .A(G137), .B(n1230), .Z(G39) );
NOR2_X1 U880 ( .A1(n1231), .A2(n1194), .ZN(n1230) );
XOR2_X1 U881 ( .A(n1195), .B(KEYINPUT12), .Z(n1231) );
NAND2_X1 U882 ( .A1(n1225), .A2(n1202), .ZN(n1195) );
XNOR2_X1 U883 ( .A(G134), .B(n1189), .ZN(G36) );
NAND4_X1 U884 ( .A1(n1059), .A2(n1225), .A3(n1062), .A4(n1038), .ZN(n1189) );
XNOR2_X1 U885 ( .A(G131), .B(n1188), .ZN(G33) );
NAND2_X1 U886 ( .A1(n1229), .A2(n1062), .ZN(n1188) );
AND3_X1 U887 ( .A1(n1225), .A2(n1074), .A3(n1059), .ZN(n1229) );
INV_X1 U888 ( .A(n1194), .ZN(n1059) );
NAND2_X1 U889 ( .A1(n1068), .A2(n1232), .ZN(n1194) );
XNOR2_X1 U890 ( .A(G128), .B(n1187), .ZN(G30) );
NAND2_X1 U891 ( .A1(n1224), .A2(n1038), .ZN(n1187) );
AND4_X1 U892 ( .A1(n1225), .A2(n1041), .A3(n1093), .A4(n1091), .ZN(n1224) );
AND2_X1 U893 ( .A1(n1211), .A2(n1233), .ZN(n1225) );
XOR2_X1 U894 ( .A(G101), .B(n1234), .Z(G3) );
NOR2_X1 U895 ( .A1(n1065), .A2(n1208), .ZN(n1234) );
NAND3_X1 U896 ( .A1(n1062), .A2(n1210), .A3(n1209), .ZN(n1208) );
INV_X1 U897 ( .A(n1041), .ZN(n1065) );
XNOR2_X1 U898 ( .A(G125), .B(n1186), .ZN(G27) );
NAND4_X1 U899 ( .A1(n1061), .A2(n1054), .A3(n1235), .A4(n1074), .ZN(n1186) );
AND2_X1 U900 ( .A1(n1233), .A2(n1041), .ZN(n1235) );
NAND2_X1 U901 ( .A1(n1236), .A2(n1237), .ZN(n1233) );
NAND2_X1 U902 ( .A1(n1238), .A2(n1106), .ZN(n1237) );
INV_X1 U903 ( .A(G900), .ZN(n1106) );
XOR2_X1 U904 ( .A(n1197), .B(n1239), .Z(G24) );
XNOR2_X1 U905 ( .A(G122), .B(KEYINPUT27), .ZN(n1239) );
NAND4_X1 U906 ( .A1(n1203), .A2(n1063), .A3(n1240), .A4(n1241), .ZN(n1197) );
AND2_X1 U907 ( .A1(n1242), .A2(n1243), .ZN(n1063) );
XNOR2_X1 U908 ( .A(n1093), .B(KEYINPUT21), .ZN(n1242) );
XNOR2_X1 U909 ( .A(G119), .B(n1244), .ZN(G21) );
NAND3_X1 U910 ( .A1(n1245), .A2(n1246), .A3(n1202), .ZN(n1244) );
AND3_X1 U911 ( .A1(n1093), .A2(n1091), .A3(n1056), .ZN(n1202) );
OR2_X1 U912 ( .A1(n1203), .A2(KEYINPUT1), .ZN(n1246) );
NAND2_X1 U913 ( .A1(KEYINPUT1), .A2(n1247), .ZN(n1245) );
NAND3_X1 U914 ( .A1(n1054), .A2(n1041), .A3(n1248), .ZN(n1247) );
INV_X1 U915 ( .A(n1210), .ZN(n1248) );
XNOR2_X1 U916 ( .A(G116), .B(n1200), .ZN(G18) );
NAND3_X1 U917 ( .A1(n1203), .A2(n1038), .A3(n1062), .ZN(n1200) );
NOR2_X1 U918 ( .A1(n1240), .A2(n1227), .ZN(n1038) );
INV_X1 U919 ( .A(n1241), .ZN(n1227) );
NAND2_X1 U920 ( .A1(n1249), .A2(n1250), .ZN(G15) );
NAND2_X1 U921 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
NAND2_X1 U922 ( .A1(G113), .A2(n1253), .ZN(n1249) );
NAND2_X1 U923 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U924 ( .A1(KEYINPUT51), .A2(n1256), .ZN(n1255) );
INV_X1 U925 ( .A(n1201), .ZN(n1256) );
OR2_X1 U926 ( .A1(n1251), .A2(KEYINPUT51), .ZN(n1254) );
NOR2_X1 U927 ( .A1(KEYINPUT57), .A2(n1201), .ZN(n1251) );
NAND3_X1 U928 ( .A1(n1203), .A2(n1074), .A3(n1062), .ZN(n1201) );
NOR2_X1 U929 ( .A1(n1093), .A2(n1243), .ZN(n1062) );
NOR2_X1 U930 ( .A1(n1241), .A2(n1228), .ZN(n1074) );
AND3_X1 U931 ( .A1(n1041), .A2(n1210), .A3(n1054), .ZN(n1203) );
AND2_X1 U932 ( .A1(n1075), .A2(n1087), .ZN(n1054) );
XNOR2_X1 U933 ( .A(G110), .B(n1257), .ZN(G12) );
NAND4_X1 U934 ( .A1(n1258), .A2(n1209), .A3(n1041), .A4(n1210), .ZN(n1257) );
NAND2_X1 U935 ( .A1(n1236), .A2(n1259), .ZN(n1210) );
NAND2_X1 U936 ( .A1(n1238), .A2(n1126), .ZN(n1259) );
INV_X1 U937 ( .A(G898), .ZN(n1126) );
AND3_X1 U938 ( .A1(G902), .A2(n1050), .A3(G953), .ZN(n1238) );
NAND3_X1 U939 ( .A1(n1050), .A2(n1048), .A3(n1260), .ZN(n1236) );
XNOR2_X1 U940 ( .A(G952), .B(KEYINPUT4), .ZN(n1260) );
NAND2_X1 U941 ( .A1(G237), .A2(G234), .ZN(n1050) );
NOR2_X1 U942 ( .A1(n1068), .A2(n1067), .ZN(n1041) );
INV_X1 U943 ( .A(n1232), .ZN(n1067) );
NAND2_X1 U944 ( .A1(G214), .A2(n1261), .ZN(n1232) );
XOR2_X1 U945 ( .A(n1079), .B(KEYINPUT9), .Z(n1068) );
XNOR2_X1 U946 ( .A(n1262), .B(n1182), .ZN(n1079) );
NAND2_X1 U947 ( .A1(G210), .A2(n1261), .ZN(n1182) );
NAND2_X1 U948 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
INV_X1 U949 ( .A(G237), .ZN(n1263) );
NAND2_X1 U950 ( .A1(n1265), .A2(n1264), .ZN(n1262) );
XOR2_X1 U951 ( .A(n1216), .B(n1266), .Z(n1265) );
XOR2_X1 U952 ( .A(n1219), .B(n1267), .Z(n1266) );
NAND2_X1 U953 ( .A1(KEYINPUT6), .A2(n1268), .ZN(n1267) );
XNOR2_X1 U954 ( .A(n1269), .B(n1220), .ZN(n1268) );
NAND2_X1 U955 ( .A1(KEYINPUT14), .A2(n1270), .ZN(n1269) );
NAND2_X1 U956 ( .A1(G224), .A2(n1048), .ZN(n1219) );
XOR2_X1 U957 ( .A(n1271), .B(n1133), .Z(n1216) );
XNOR2_X1 U958 ( .A(G110), .B(G122), .ZN(n1133) );
XOR2_X1 U959 ( .A(n1129), .B(n1272), .Z(n1271) );
NOR2_X1 U960 ( .A1(KEYINPUT34), .A2(n1130), .ZN(n1272) );
XNOR2_X1 U961 ( .A(n1273), .B(n1274), .ZN(n1130) );
XNOR2_X1 U962 ( .A(n1275), .B(KEYINPUT19), .ZN(n1274) );
NAND2_X1 U963 ( .A1(KEYINPUT15), .A2(n1276), .ZN(n1275) );
XOR2_X1 U964 ( .A(KEYINPUT61), .B(n1277), .Z(n1276) );
XOR2_X1 U965 ( .A(n1278), .B(G101), .Z(n1129) );
NAND3_X1 U966 ( .A1(n1279), .A2(n1280), .A3(n1281), .ZN(n1278) );
OR2_X1 U967 ( .A1(G107), .A2(KEYINPUT48), .ZN(n1281) );
NAND3_X1 U968 ( .A1(KEYINPUT48), .A2(G107), .A3(n1282), .ZN(n1280) );
NAND2_X1 U969 ( .A1(G104), .A2(n1283), .ZN(n1279) );
NAND2_X1 U970 ( .A1(n1284), .A2(KEYINPUT48), .ZN(n1283) );
XNOR2_X1 U971 ( .A(G107), .B(KEYINPUT37), .ZN(n1284) );
INV_X1 U972 ( .A(n1071), .ZN(n1209) );
NAND2_X1 U973 ( .A1(n1056), .A2(n1211), .ZN(n1071) );
NOR2_X1 U974 ( .A1(n1076), .A2(n1075), .ZN(n1211) );
NOR2_X1 U975 ( .A1(n1083), .A2(n1285), .ZN(n1075) );
AND2_X1 U976 ( .A1(G469), .A2(n1089), .ZN(n1285) );
NOR2_X1 U977 ( .A1(n1089), .A2(G469), .ZN(n1083) );
NAND2_X1 U978 ( .A1(n1286), .A2(n1264), .ZN(n1089) );
XOR2_X1 U979 ( .A(n1287), .B(n1288), .Z(n1286) );
XOR2_X1 U980 ( .A(n1178), .B(n1170), .Z(n1288) );
XNOR2_X1 U981 ( .A(n1289), .B(n1290), .ZN(n1170) );
XNOR2_X1 U982 ( .A(n1291), .B(G110), .ZN(n1290) );
INV_X1 U983 ( .A(G140), .ZN(n1291) );
NAND2_X1 U984 ( .A1(n1292), .A2(n1048), .ZN(n1289) );
XNOR2_X1 U985 ( .A(G227), .B(KEYINPUT24), .ZN(n1292) );
XNOR2_X1 U986 ( .A(n1293), .B(n1294), .ZN(n1178) );
XNOR2_X1 U987 ( .A(KEYINPUT40), .B(n1036), .ZN(n1294) );
INV_X1 U988 ( .A(G107), .ZN(n1036) );
XOR2_X1 U989 ( .A(n1295), .B(G101), .Z(n1293) );
NAND2_X1 U990 ( .A1(KEYINPUT10), .A2(n1282), .ZN(n1295) );
XOR2_X1 U991 ( .A(n1296), .B(n1175), .Z(n1287) );
XNOR2_X1 U992 ( .A(n1297), .B(KEYINPUT44), .ZN(n1175) );
NAND2_X1 U993 ( .A1(KEYINPUT63), .A2(n1114), .ZN(n1296) );
XOR2_X1 U994 ( .A(n1298), .B(G128), .Z(n1114) );
NAND2_X1 U995 ( .A1(KEYINPUT45), .A2(n1299), .ZN(n1298) );
XNOR2_X1 U996 ( .A(n1300), .B(n1301), .ZN(n1299) );
INV_X1 U997 ( .A(n1087), .ZN(n1076) );
NAND2_X1 U998 ( .A1(G221), .A2(n1302), .ZN(n1087) );
NOR2_X1 U999 ( .A1(n1241), .A2(n1240), .ZN(n1056) );
INV_X1 U1000 ( .A(n1228), .ZN(n1240) );
XOR2_X1 U1001 ( .A(n1094), .B(n1149), .Z(n1228) );
INV_X1 U1002 ( .A(G475), .ZN(n1149) );
NOR2_X1 U1003 ( .A1(n1150), .A2(G902), .ZN(n1094) );
XNOR2_X1 U1004 ( .A(n1303), .B(n1304), .ZN(n1150) );
XOR2_X1 U1005 ( .A(n1305), .B(n1306), .Z(n1304) );
XNOR2_X1 U1006 ( .A(n1307), .B(n1308), .ZN(n1306) );
NAND2_X1 U1007 ( .A1(KEYINPUT3), .A2(n1300), .ZN(n1308) );
NAND2_X1 U1008 ( .A1(KEYINPUT33), .A2(n1282), .ZN(n1307) );
INV_X1 U1009 ( .A(G104), .ZN(n1282) );
NAND2_X1 U1010 ( .A1(G214), .A2(n1309), .ZN(n1305) );
XOR2_X1 U1011 ( .A(n1310), .B(n1311), .Z(n1303) );
XOR2_X1 U1012 ( .A(G131), .B(G122), .Z(n1311) );
XNOR2_X1 U1013 ( .A(n1312), .B(n1252), .ZN(n1310) );
NAND3_X1 U1014 ( .A1(n1313), .A2(n1314), .A3(n1315), .ZN(n1312) );
XNOR2_X1 U1015 ( .A(KEYINPUT62), .B(KEYINPUT50), .ZN(n1315) );
NAND2_X1 U1016 ( .A1(KEYINPUT42), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U1017 ( .A(n1317), .B(n1108), .ZN(n1316) );
NAND2_X1 U1018 ( .A1(KEYINPUT46), .A2(n1318), .ZN(n1317) );
OR3_X1 U1019 ( .A1(n1318), .A2(n1108), .A3(KEYINPUT42), .ZN(n1313) );
INV_X1 U1020 ( .A(n1111), .ZN(n1108) );
NAND2_X1 U1021 ( .A1(n1096), .A2(n1085), .ZN(n1241) );
NAND3_X1 U1022 ( .A1(n1319), .A2(n1144), .A3(n1143), .ZN(n1085) );
INV_X1 U1023 ( .A(G478), .ZN(n1144) );
NAND2_X1 U1024 ( .A1(G478), .A2(n1320), .ZN(n1096) );
NAND2_X1 U1025 ( .A1(n1143), .A2(n1319), .ZN(n1320) );
XNOR2_X1 U1026 ( .A(KEYINPUT28), .B(n1264), .ZN(n1319) );
XOR2_X1 U1027 ( .A(n1321), .B(n1322), .Z(n1143) );
XOR2_X1 U1028 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR3_X1 U1029 ( .A1(n1325), .A2(G953), .A3(n1139), .ZN(n1323) );
XNOR2_X1 U1030 ( .A(n1326), .B(n1327), .ZN(n1321) );
NAND2_X1 U1031 ( .A1(KEYINPUT25), .A2(n1328), .ZN(n1327) );
INV_X1 U1032 ( .A(G134), .ZN(n1328) );
NAND2_X1 U1033 ( .A1(KEYINPUT13), .A2(n1329), .ZN(n1326) );
XOR2_X1 U1034 ( .A(n1330), .B(n1331), .Z(n1329) );
XNOR2_X1 U1035 ( .A(G116), .B(G107), .ZN(n1331) );
NAND2_X1 U1036 ( .A1(KEYINPUT26), .A2(G122), .ZN(n1330) );
XNOR2_X1 U1037 ( .A(n1061), .B(KEYINPUT60), .ZN(n1258) );
AND2_X1 U1038 ( .A1(n1243), .A2(n1093), .ZN(n1061) );
XNOR2_X1 U1039 ( .A(n1332), .B(n1333), .ZN(n1093) );
NOR2_X1 U1040 ( .A1(n1334), .A2(n1139), .ZN(n1333) );
INV_X1 U1041 ( .A(G217), .ZN(n1139) );
XOR2_X1 U1042 ( .A(n1302), .B(KEYINPUT16), .Z(n1334) );
NAND2_X1 U1043 ( .A1(G234), .A2(n1264), .ZN(n1302) );
NAND2_X1 U1044 ( .A1(n1137), .A2(n1264), .ZN(n1332) );
XNOR2_X1 U1045 ( .A(n1335), .B(n1336), .ZN(n1137) );
XNOR2_X1 U1046 ( .A(n1111), .B(n1337), .ZN(n1336) );
XOR2_X1 U1047 ( .A(n1338), .B(n1339), .Z(n1337) );
NOR3_X1 U1048 ( .A1(n1340), .A2(n1325), .A3(n1341), .ZN(n1339) );
INV_X1 U1049 ( .A(G221), .ZN(n1341) );
INV_X1 U1050 ( .A(G234), .ZN(n1325) );
XNOR2_X1 U1051 ( .A(KEYINPUT39), .B(n1048), .ZN(n1340) );
INV_X1 U1052 ( .A(G953), .ZN(n1048) );
NAND2_X1 U1053 ( .A1(KEYINPUT56), .A2(n1342), .ZN(n1338) );
XOR2_X1 U1054 ( .A(G128), .B(G119), .Z(n1342) );
XNOR2_X1 U1055 ( .A(G140), .B(n1270), .ZN(n1111) );
INV_X1 U1056 ( .A(G125), .ZN(n1270) );
XNOR2_X1 U1057 ( .A(G110), .B(n1343), .ZN(n1335) );
XNOR2_X1 U1058 ( .A(n1318), .B(G137), .ZN(n1343) );
INV_X1 U1059 ( .A(n1091), .ZN(n1243) );
XOR2_X1 U1060 ( .A(n1344), .B(n1160), .Z(n1091) );
INV_X1 U1061 ( .A(G472), .ZN(n1160) );
NAND2_X1 U1062 ( .A1(n1345), .A2(n1264), .ZN(n1344) );
INV_X1 U1063 ( .A(G902), .ZN(n1264) );
XNOR2_X1 U1064 ( .A(n1346), .B(n1159), .ZN(n1345) );
XNOR2_X1 U1065 ( .A(n1347), .B(G101), .ZN(n1159) );
NAND2_X1 U1066 ( .A1(G210), .A2(n1309), .ZN(n1347) );
NOR2_X1 U1067 ( .A1(G953), .A2(G237), .ZN(n1309) );
NAND4_X1 U1068 ( .A1(n1348), .A2(n1349), .A3(n1350), .A4(n1351), .ZN(n1346) );
NAND3_X1 U1069 ( .A1(KEYINPUT53), .A2(n1166), .A3(n1165), .ZN(n1351) );
INV_X1 U1070 ( .A(n1220), .ZN(n1166) );
NAND3_X1 U1071 ( .A1(n1220), .A2(n1352), .A3(n1353), .ZN(n1350) );
NAND2_X1 U1072 ( .A1(n1167), .A2(n1354), .ZN(n1352) );
INV_X1 U1073 ( .A(n1164), .ZN(n1349) );
NOR3_X1 U1074 ( .A1(n1353), .A2(n1167), .A3(n1220), .ZN(n1164) );
NAND2_X1 U1075 ( .A1(n1163), .A2(n1354), .ZN(n1348) );
INV_X1 U1076 ( .A(KEYINPUT53), .ZN(n1354) );
AND2_X1 U1077 ( .A1(n1167), .A2(n1355), .ZN(n1163) );
XNOR2_X1 U1078 ( .A(n1220), .B(n1165), .ZN(n1355) );
INV_X1 U1079 ( .A(n1353), .ZN(n1165) );
XOR2_X1 U1080 ( .A(n1277), .B(n1356), .Z(n1353) );
XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(n1273), .ZN(n1356) );
XOR2_X1 U1082 ( .A(n1252), .B(KEYINPUT32), .Z(n1273) );
INV_X1 U1083 ( .A(G113), .ZN(n1252) );
XOR2_X1 U1084 ( .A(G116), .B(G119), .Z(n1277) );
XOR2_X1 U1085 ( .A(n1324), .B(n1301), .Z(n1220) );
XNOR2_X1 U1086 ( .A(n1318), .B(KEYINPUT8), .ZN(n1301) );
INV_X1 U1087 ( .A(G146), .ZN(n1318) );
XNOR2_X1 U1088 ( .A(G128), .B(n1300), .ZN(n1324) );
INV_X1 U1089 ( .A(G143), .ZN(n1300) );
INV_X1 U1090 ( .A(n1297), .ZN(n1167) );
XNOR2_X1 U1091 ( .A(n1357), .B(n1358), .ZN(n1297) );
NOR2_X1 U1092 ( .A1(KEYINPUT7), .A2(G131), .ZN(n1358) );
XNOR2_X1 U1093 ( .A(G134), .B(G137), .ZN(n1357) );
endmodule


