//Key = 1000100001101000001101101101101111010010101001101101111111100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402;

NAND2_X1 U768 ( .A1(n1064), .A2(n1065), .ZN(G9) );
NAND2_X1 U769 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
XOR2_X1 U770 ( .A(n1068), .B(KEYINPUT46), .Z(n1066) );
NAND2_X1 U771 ( .A1(n1069), .A2(G107), .ZN(n1064) );
XNOR2_X1 U772 ( .A(KEYINPUT25), .B(n1068), .ZN(n1069) );
NAND2_X1 U773 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
XNOR2_X1 U774 ( .A(KEYINPUT8), .B(n1072), .ZN(n1071) );
NOR2_X1 U775 ( .A1(n1073), .A2(n1074), .ZN(G75) );
NOR3_X1 U776 ( .A1(n1075), .A2(G953), .A3(G952), .ZN(n1074) );
INV_X1 U777 ( .A(n1076), .ZN(n1075) );
NOR3_X1 U778 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1073) );
NOR2_X1 U779 ( .A1(n1080), .A2(n1081), .ZN(n1078) );
NOR3_X1 U780 ( .A1(n1082), .A2(n1083), .A3(n1084), .ZN(n1080) );
NOR2_X1 U781 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
INV_X1 U782 ( .A(n1087), .ZN(n1086) );
NOR2_X1 U783 ( .A1(n1088), .A2(n1089), .ZN(n1085) );
AND2_X1 U784 ( .A1(n1090), .A2(n1091), .ZN(n1088) );
NOR3_X1 U785 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1083) );
NOR2_X1 U786 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NOR2_X1 U787 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NOR2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1097) );
NOR2_X1 U789 ( .A1(n1101), .A2(n1102), .ZN(n1099) );
NOR2_X1 U790 ( .A1(n1103), .A2(n1104), .ZN(n1095) );
NOR2_X1 U791 ( .A1(n1105), .A2(n1106), .ZN(n1103) );
AND2_X1 U792 ( .A1(n1107), .A2(KEYINPUT22), .ZN(n1105) );
NOR2_X1 U793 ( .A1(n1108), .A2(KEYINPUT22), .ZN(n1082) );
NOR4_X1 U794 ( .A1(n1094), .A2(n1109), .A3(n1104), .A4(n1092), .ZN(n1108) );
NAND3_X1 U795 ( .A1(n1110), .A2(n1111), .A3(n1076), .ZN(n1077) );
NAND4_X1 U796 ( .A1(n1112), .A2(n1113), .A3(n1114), .A4(n1115), .ZN(n1076) );
NOR4_X1 U797 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1115) );
XOR2_X1 U798 ( .A(n1120), .B(KEYINPUT45), .Z(n1119) );
NOR2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1118) );
NOR2_X1 U800 ( .A1(n1123), .A2(n1124), .ZN(n1117) );
AND2_X1 U801 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
XOR2_X1 U802 ( .A(n1127), .B(n1128), .Z(n1113) );
NAND2_X1 U803 ( .A1(KEYINPUT54), .A2(n1129), .ZN(n1128) );
XOR2_X1 U804 ( .A(KEYINPUT43), .B(n1130), .Z(n1112) );
NOR4_X1 U805 ( .A1(n1131), .A2(n1081), .A3(n1132), .A4(n1133), .ZN(n1130) );
AND3_X1 U806 ( .A1(KEYINPUT32), .A2(n1134), .A3(G469), .ZN(n1133) );
NOR2_X1 U807 ( .A1(KEYINPUT32), .A2(G469), .ZN(n1132) );
NAND2_X1 U808 ( .A1(n1102), .A2(n1135), .ZN(n1131) );
NAND3_X1 U809 ( .A1(n1136), .A2(n1137), .A3(n1087), .ZN(n1110) );
NOR3_X1 U810 ( .A1(n1092), .A2(n1104), .A3(n1098), .ZN(n1087) );
NAND2_X1 U811 ( .A1(n1138), .A2(n1139), .ZN(n1137) );
NAND2_X1 U812 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
XOR2_X1 U813 ( .A(n1142), .B(n1143), .Z(G72) );
NOR2_X1 U814 ( .A1(n1144), .A2(n1111), .ZN(n1143) );
NOR2_X1 U815 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
NAND2_X1 U816 ( .A1(n1147), .A2(n1148), .ZN(n1142) );
NAND2_X1 U817 ( .A1(n1149), .A2(n1111), .ZN(n1148) );
XOR2_X1 U818 ( .A(n1150), .B(n1151), .Z(n1149) );
NAND2_X1 U819 ( .A1(n1152), .A2(n1153), .ZN(n1150) );
NAND3_X1 U820 ( .A1(G900), .A2(n1151), .A3(G953), .ZN(n1147) );
XOR2_X1 U821 ( .A(n1154), .B(n1155), .Z(n1151) );
XOR2_X1 U822 ( .A(n1156), .B(n1157), .Z(n1155) );
XNOR2_X1 U823 ( .A(n1158), .B(n1159), .ZN(n1154) );
NOR2_X1 U824 ( .A1(n1160), .A2(KEYINPUT34), .ZN(n1159) );
NOR3_X1 U825 ( .A1(KEYINPUT17), .A2(n1161), .A3(n1162), .ZN(n1158) );
NOR3_X1 U826 ( .A1(n1163), .A2(G137), .A3(n1164), .ZN(n1162) );
INV_X1 U827 ( .A(KEYINPUT62), .ZN(n1163) );
NOR2_X1 U828 ( .A1(KEYINPUT62), .A2(n1165), .ZN(n1161) );
XOR2_X1 U829 ( .A(n1166), .B(n1167), .Z(G69) );
NAND2_X1 U830 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
NAND2_X1 U831 ( .A1(G953), .A2(n1170), .ZN(n1169) );
NAND2_X1 U832 ( .A1(G224), .A2(n1171), .ZN(n1170) );
NAND2_X1 U833 ( .A1(KEYINPUT60), .A2(G898), .ZN(n1171) );
NAND2_X1 U834 ( .A1(n1172), .A2(n1173), .ZN(n1168) );
INV_X1 U835 ( .A(KEYINPUT60), .ZN(n1173) );
NAND2_X1 U836 ( .A1(n1174), .A2(KEYINPUT28), .ZN(n1166) );
XOR2_X1 U837 ( .A(n1175), .B(n1176), .Z(n1174) );
NOR2_X1 U838 ( .A1(n1172), .A2(n1177), .ZN(n1176) );
XNOR2_X1 U839 ( .A(n1178), .B(n1179), .ZN(n1177) );
XOR2_X1 U840 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U841 ( .A1(KEYINPUT27), .A2(n1182), .ZN(n1181) );
NAND2_X1 U842 ( .A1(n1183), .A2(n1111), .ZN(n1175) );
XOR2_X1 U843 ( .A(KEYINPUT57), .B(n1184), .Z(n1183) );
NOR2_X1 U844 ( .A1(n1185), .A2(n1186), .ZN(G66) );
XOR2_X1 U845 ( .A(n1187), .B(n1188), .Z(n1186) );
NOR2_X1 U846 ( .A1(n1189), .A2(KEYINPUT50), .ZN(n1188) );
OR2_X1 U847 ( .A1(n1190), .A2(n1122), .ZN(n1187) );
NOR2_X1 U848 ( .A1(n1185), .A2(n1191), .ZN(G63) );
XNOR2_X1 U849 ( .A(n1192), .B(n1126), .ZN(n1191) );
NOR2_X1 U850 ( .A1(n1124), .A2(n1190), .ZN(n1192) );
NOR2_X1 U851 ( .A1(n1185), .A2(n1193), .ZN(G60) );
XOR2_X1 U852 ( .A(n1194), .B(n1195), .Z(n1193) );
NOR2_X1 U853 ( .A1(n1196), .A2(n1190), .ZN(n1194) );
XNOR2_X1 U854 ( .A(n1197), .B(n1198), .ZN(G6) );
NOR3_X1 U855 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1198) );
XNOR2_X1 U856 ( .A(KEYINPUT40), .B(n1094), .ZN(n1199) );
NOR3_X1 U857 ( .A1(n1185), .A2(n1202), .A3(n1203), .ZN(G57) );
NOR2_X1 U858 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
NOR2_X1 U859 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
AND2_X1 U860 ( .A1(KEYINPUT37), .A2(n1208), .ZN(n1207) );
NOR3_X1 U861 ( .A1(KEYINPUT37), .A2(n1208), .A3(n1209), .ZN(n1206) );
NOR2_X1 U862 ( .A1(n1210), .A2(n1211), .ZN(n1202) );
INV_X1 U863 ( .A(n1204), .ZN(n1211) );
XOR2_X1 U864 ( .A(n1212), .B(n1213), .Z(n1204) );
XOR2_X1 U865 ( .A(n1214), .B(n1215), .Z(n1213) );
NOR2_X1 U866 ( .A1(KEYINPUT5), .A2(n1216), .ZN(n1215) );
NOR2_X1 U867 ( .A1(n1217), .A2(n1190), .ZN(n1214) );
NOR2_X1 U868 ( .A1(n1208), .A2(n1209), .ZN(n1210) );
INV_X1 U869 ( .A(KEYINPUT56), .ZN(n1209) );
XOR2_X1 U870 ( .A(n1218), .B(KEYINPUT6), .Z(n1208) );
NOR2_X1 U871 ( .A1(n1185), .A2(n1219), .ZN(G54) );
XOR2_X1 U872 ( .A(n1220), .B(n1221), .Z(n1219) );
XOR2_X1 U873 ( .A(n1222), .B(n1223), .Z(n1220) );
NOR2_X1 U874 ( .A1(n1224), .A2(n1190), .ZN(n1223) );
INV_X1 U875 ( .A(G469), .ZN(n1224) );
NAND2_X1 U876 ( .A1(n1225), .A2(n1226), .ZN(n1222) );
NAND2_X1 U877 ( .A1(n1227), .A2(n1228), .ZN(n1226) );
XOR2_X1 U878 ( .A(KEYINPUT42), .B(n1229), .Z(n1225) );
NOR2_X1 U879 ( .A1(n1227), .A2(n1228), .ZN(n1229) );
XNOR2_X1 U880 ( .A(n1230), .B(G110), .ZN(n1228) );
NAND2_X1 U881 ( .A1(KEYINPUT4), .A2(n1231), .ZN(n1230) );
NOR2_X1 U882 ( .A1(n1185), .A2(n1232), .ZN(G51) );
XOR2_X1 U883 ( .A(n1233), .B(n1234), .Z(n1232) );
XOR2_X1 U884 ( .A(n1235), .B(n1236), .Z(n1234) );
NAND2_X1 U885 ( .A1(KEYINPUT21), .A2(n1237), .ZN(n1235) );
XOR2_X1 U886 ( .A(KEYINPUT38), .B(n1238), .Z(n1237) );
XOR2_X1 U887 ( .A(n1239), .B(n1240), .Z(n1233) );
NOR2_X1 U888 ( .A1(n1241), .A2(n1190), .ZN(n1240) );
NAND2_X1 U889 ( .A1(G902), .A2(n1079), .ZN(n1190) );
NAND3_X1 U890 ( .A1(n1184), .A2(n1152), .A3(n1242), .ZN(n1079) );
XNOR2_X1 U891 ( .A(n1243), .B(KEYINPUT26), .ZN(n1242) );
AND4_X1 U892 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1152) );
NOR3_X1 U893 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
NOR3_X1 U894 ( .A1(n1251), .A2(n1252), .A3(n1201), .ZN(n1250) );
XNOR2_X1 U895 ( .A(n1253), .B(KEYINPUT3), .ZN(n1252) );
NOR2_X1 U896 ( .A1(n1254), .A2(n1138), .ZN(n1248) );
NOR2_X1 U897 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
AND2_X1 U898 ( .A1(n1257), .A2(n1258), .ZN(n1255) );
AND4_X1 U899 ( .A1(n1259), .A2(n1260), .A3(n1261), .A4(n1262), .ZN(n1184) );
NOR4_X1 U900 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1262) );
NOR2_X1 U901 ( .A1(n1072), .A2(n1138), .ZN(n1266) );
NAND4_X1 U902 ( .A1(n1107), .A2(n1136), .A3(n1267), .A4(n1268), .ZN(n1072) );
NOR3_X1 U903 ( .A1(n1201), .A2(n1094), .A3(n1200), .ZN(n1265) );
INV_X1 U904 ( .A(n1106), .ZN(n1201) );
INV_X1 U905 ( .A(n1269), .ZN(n1264) );
INV_X1 U906 ( .A(n1270), .ZN(n1263) );
NOR2_X1 U907 ( .A1(n1271), .A2(n1272), .ZN(n1261) );
NAND3_X1 U908 ( .A1(n1273), .A2(n1136), .A3(n1257), .ZN(n1260) );
NOR2_X1 U909 ( .A1(n1111), .A2(G952), .ZN(n1185) );
XOR2_X1 U910 ( .A(n1274), .B(n1275), .Z(G48) );
XNOR2_X1 U911 ( .A(G146), .B(KEYINPUT29), .ZN(n1275) );
NAND2_X1 U912 ( .A1(n1276), .A2(n1070), .ZN(n1274) );
XNOR2_X1 U913 ( .A(n1256), .B(KEYINPUT24), .ZN(n1276) );
AND3_X1 U914 ( .A1(n1106), .A2(n1100), .A3(n1277), .ZN(n1256) );
XOR2_X1 U915 ( .A(n1278), .B(n1279), .Z(G45) );
NAND2_X1 U916 ( .A1(KEYINPUT33), .A2(G143), .ZN(n1279) );
NAND3_X1 U917 ( .A1(n1257), .A2(n1280), .A3(n1258), .ZN(n1278) );
INV_X1 U918 ( .A(n1251), .ZN(n1258) );
XNOR2_X1 U919 ( .A(KEYINPUT23), .B(n1138), .ZN(n1280) );
XNOR2_X1 U920 ( .A(n1231), .B(n1249), .ZN(G42) );
AND3_X1 U921 ( .A1(n1253), .A2(n1100), .A3(n1281), .ZN(n1249) );
XOR2_X1 U922 ( .A(n1246), .B(n1282), .Z(G39) );
NAND2_X1 U923 ( .A1(KEYINPUT9), .A2(G137), .ZN(n1282) );
NAND4_X1 U924 ( .A1(n1253), .A2(n1277), .A3(n1283), .A4(n1100), .ZN(n1246) );
INV_X1 U925 ( .A(n1081), .ZN(n1253) );
XNOR2_X1 U926 ( .A(G134), .B(n1244), .ZN(G36) );
NAND2_X1 U927 ( .A1(n1284), .A2(n1107), .ZN(n1244) );
XNOR2_X1 U928 ( .A(G131), .B(n1285), .ZN(G33) );
NAND2_X1 U929 ( .A1(n1284), .A2(n1106), .ZN(n1285) );
NOR2_X1 U930 ( .A1(n1251), .A2(n1081), .ZN(n1284) );
NAND2_X1 U931 ( .A1(n1141), .A2(n1286), .ZN(n1081) );
NAND3_X1 U932 ( .A1(n1100), .A2(n1287), .A3(n1089), .ZN(n1251) );
XNOR2_X1 U933 ( .A(G128), .B(n1245), .ZN(G30) );
NAND4_X1 U934 ( .A1(n1277), .A2(n1070), .A3(n1107), .A4(n1267), .ZN(n1245) );
AND3_X1 U935 ( .A1(n1287), .A2(n1090), .A3(n1288), .ZN(n1277) );
XOR2_X1 U936 ( .A(G101), .B(n1272), .Z(G3) );
AND3_X1 U937 ( .A1(n1289), .A2(n1283), .A3(n1089), .ZN(n1272) );
XNOR2_X1 U938 ( .A(G125), .B(n1290), .ZN(G27) );
NAND2_X1 U939 ( .A1(KEYINPUT0), .A2(n1243), .ZN(n1290) );
INV_X1 U940 ( .A(n1153), .ZN(n1243) );
NAND3_X1 U941 ( .A1(n1291), .A2(n1070), .A3(n1281), .ZN(n1153) );
AND4_X1 U942 ( .A1(n1106), .A2(n1091), .A3(n1287), .A4(n1090), .ZN(n1281) );
NAND2_X1 U943 ( .A1(n1092), .A2(n1292), .ZN(n1287) );
NAND4_X1 U944 ( .A1(G902), .A2(G953), .A3(n1293), .A4(n1146), .ZN(n1292) );
INV_X1 U945 ( .A(G900), .ZN(n1146) );
XNOR2_X1 U946 ( .A(G122), .B(n1294), .ZN(G24) );
NAND4_X1 U947 ( .A1(n1295), .A2(n1257), .A3(n1296), .A4(n1291), .ZN(n1294) );
NOR2_X1 U948 ( .A1(n1297), .A2(n1094), .ZN(n1296) );
INV_X1 U949 ( .A(n1136), .ZN(n1094) );
NOR2_X1 U950 ( .A1(n1090), .A2(n1288), .ZN(n1136) );
NOR2_X1 U951 ( .A1(n1114), .A2(n1298), .ZN(n1257) );
XNOR2_X1 U952 ( .A(n1070), .B(KEYINPUT12), .ZN(n1295) );
XOR2_X1 U953 ( .A(G119), .B(n1271), .Z(G21) );
AND4_X1 U954 ( .A1(n1288), .A2(n1273), .A3(n1283), .A4(n1090), .ZN(n1271) );
INV_X1 U955 ( .A(n1091), .ZN(n1288) );
XNOR2_X1 U956 ( .A(G116), .B(n1269), .ZN(G18) );
NAND3_X1 U957 ( .A1(n1273), .A2(n1107), .A3(n1089), .ZN(n1269) );
INV_X1 U958 ( .A(n1109), .ZN(n1107) );
NAND2_X1 U959 ( .A1(n1114), .A2(n1299), .ZN(n1109) );
XNOR2_X1 U960 ( .A(n1300), .B(n1301), .ZN(G15) );
NOR2_X1 U961 ( .A1(KEYINPUT44), .A2(n1270), .ZN(n1301) );
NAND3_X1 U962 ( .A1(n1089), .A2(n1273), .A3(n1106), .ZN(n1270) );
NOR2_X1 U963 ( .A1(n1299), .A2(n1114), .ZN(n1106) );
NOR3_X1 U964 ( .A1(n1138), .A2(n1297), .A3(n1104), .ZN(n1273) );
INV_X1 U965 ( .A(n1291), .ZN(n1104) );
NOR2_X1 U966 ( .A1(n1101), .A2(n1302), .ZN(n1291) );
INV_X1 U967 ( .A(n1102), .ZN(n1302) );
INV_X1 U968 ( .A(n1268), .ZN(n1297) );
INV_X1 U969 ( .A(n1070), .ZN(n1138) );
NOR2_X1 U970 ( .A1(n1091), .A2(n1090), .ZN(n1089) );
XNOR2_X1 U971 ( .A(G110), .B(n1259), .ZN(G12) );
NAND4_X1 U972 ( .A1(n1289), .A2(n1283), .A3(n1091), .A4(n1090), .ZN(n1259) );
NAND2_X1 U973 ( .A1(n1303), .A2(n1304), .ZN(n1090) );
NAND2_X1 U974 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
XOR2_X1 U975 ( .A(KEYINPUT52), .B(n1116), .Z(n1303) );
NOR2_X1 U976 ( .A1(n1306), .A2(n1305), .ZN(n1116) );
INV_X1 U977 ( .A(n1122), .ZN(n1305) );
NAND2_X1 U978 ( .A1(G217), .A2(n1307), .ZN(n1122) );
INV_X1 U979 ( .A(n1121), .ZN(n1306) );
NOR2_X1 U980 ( .A1(G902), .A2(n1189), .ZN(n1121) );
AND2_X1 U981 ( .A1(n1308), .A2(n1309), .ZN(n1189) );
NAND2_X1 U982 ( .A1(n1310), .A2(n1311), .ZN(n1309) );
XOR2_X1 U983 ( .A(KEYINPUT10), .B(n1312), .Z(n1308) );
NOR2_X1 U984 ( .A1(n1310), .A2(n1311), .ZN(n1312) );
XOR2_X1 U985 ( .A(n1313), .B(n1314), .Z(n1311) );
XNOR2_X1 U986 ( .A(n1315), .B(G119), .ZN(n1314) );
INV_X1 U987 ( .A(G128), .ZN(n1315) );
XNOR2_X1 U988 ( .A(n1316), .B(G110), .ZN(n1313) );
AND2_X1 U989 ( .A1(n1317), .A2(n1318), .ZN(n1310) );
NAND2_X1 U990 ( .A1(n1319), .A2(n1320), .ZN(n1318) );
INV_X1 U991 ( .A(G137), .ZN(n1320) );
XOR2_X1 U992 ( .A(KEYINPUT58), .B(n1321), .Z(n1319) );
NAND2_X1 U993 ( .A1(n1321), .A2(G137), .ZN(n1317) );
AND3_X1 U994 ( .A1(G234), .A2(n1111), .A3(G221), .ZN(n1321) );
XNOR2_X1 U995 ( .A(n1127), .B(n1129), .ZN(n1091) );
XNOR2_X1 U996 ( .A(n1217), .B(KEYINPUT61), .ZN(n1129) );
INV_X1 U997 ( .A(G472), .ZN(n1217) );
NAND2_X1 U998 ( .A1(n1322), .A2(n1125), .ZN(n1127) );
XNOR2_X1 U999 ( .A(n1323), .B(n1324), .ZN(n1322) );
XNOR2_X1 U1000 ( .A(n1325), .B(KEYINPUT31), .ZN(n1324) );
NAND2_X1 U1001 ( .A1(n1326), .A2(KEYINPUT30), .ZN(n1325) );
XNOR2_X1 U1002 ( .A(n1216), .B(n1327), .ZN(n1326) );
INV_X1 U1003 ( .A(n1212), .ZN(n1327) );
XOR2_X1 U1004 ( .A(n1328), .B(n1300), .Z(n1212) );
NAND3_X1 U1005 ( .A1(n1329), .A2(n1330), .A3(n1331), .ZN(n1328) );
NAND2_X1 U1006 ( .A1(KEYINPUT14), .A2(G116), .ZN(n1331) );
OR3_X1 U1007 ( .A1(n1332), .A2(KEYINPUT14), .A3(G119), .ZN(n1330) );
NAND2_X1 U1008 ( .A1(G119), .A2(n1332), .ZN(n1329) );
NAND2_X1 U1009 ( .A1(KEYINPUT51), .A2(n1333), .ZN(n1332) );
INV_X1 U1010 ( .A(G116), .ZN(n1333) );
XOR2_X1 U1011 ( .A(n1334), .B(n1335), .Z(n1216) );
INV_X1 U1012 ( .A(n1218), .ZN(n1323) );
XOR2_X1 U1013 ( .A(G101), .B(n1336), .Z(n1218) );
AND3_X1 U1014 ( .A1(G210), .A2(n1111), .A3(n1337), .ZN(n1336) );
INV_X1 U1015 ( .A(n1098), .ZN(n1283) );
NAND2_X1 U1016 ( .A1(n1298), .A2(n1114), .ZN(n1098) );
XNOR2_X1 U1017 ( .A(n1338), .B(n1196), .ZN(n1114) );
INV_X1 U1018 ( .A(G475), .ZN(n1196) );
OR2_X1 U1019 ( .A1(n1195), .A2(G902), .ZN(n1338) );
XNOR2_X1 U1020 ( .A(n1339), .B(n1340), .ZN(n1195) );
XNOR2_X1 U1021 ( .A(n1341), .B(n1342), .ZN(n1340) );
XNOR2_X1 U1022 ( .A(n1197), .B(n1343), .ZN(n1342) );
NOR2_X1 U1023 ( .A1(KEYINPUT1), .A2(n1344), .ZN(n1343) );
NOR2_X1 U1024 ( .A1(n1345), .A2(n1346), .ZN(n1344) );
XOR2_X1 U1025 ( .A(n1347), .B(KEYINPUT35), .Z(n1346) );
NAND2_X1 U1026 ( .A1(n1348), .A2(n1349), .ZN(n1347) );
NAND3_X1 U1027 ( .A1(n1337), .A2(n1111), .A3(G214), .ZN(n1349) );
AND4_X1 U1028 ( .A1(n1111), .A2(n1337), .A3(G214), .A4(G143), .ZN(n1345) );
INV_X1 U1029 ( .A(n1316), .ZN(n1341) );
XOR2_X1 U1030 ( .A(G146), .B(n1157), .Z(n1316) );
XNOR2_X1 U1031 ( .A(G125), .B(n1231), .ZN(n1157) );
XNOR2_X1 U1032 ( .A(G113), .B(n1350), .ZN(n1339) );
XNOR2_X1 U1033 ( .A(G131), .B(n1351), .ZN(n1350) );
INV_X1 U1034 ( .A(n1299), .ZN(n1298) );
NAND2_X1 U1035 ( .A1(n1352), .A2(n1120), .ZN(n1299) );
NAND3_X1 U1036 ( .A1(n1124), .A2(n1125), .A3(n1126), .ZN(n1120) );
INV_X1 U1037 ( .A(G478), .ZN(n1124) );
NAND2_X1 U1038 ( .A1(G478), .A2(n1353), .ZN(n1352) );
NAND2_X1 U1039 ( .A1(n1126), .A2(n1125), .ZN(n1353) );
XOR2_X1 U1040 ( .A(n1354), .B(n1355), .Z(n1126) );
XNOR2_X1 U1041 ( .A(n1356), .B(n1164), .ZN(n1355) );
NAND2_X1 U1042 ( .A1(KEYINPUT48), .A2(n1357), .ZN(n1356) );
XNOR2_X1 U1043 ( .A(n1067), .B(n1358), .ZN(n1357) );
XNOR2_X1 U1044 ( .A(n1351), .B(G116), .ZN(n1358) );
XOR2_X1 U1045 ( .A(n1359), .B(n1360), .Z(n1354) );
NOR2_X1 U1046 ( .A1(KEYINPUT7), .A2(n1361), .ZN(n1360) );
NAND3_X1 U1047 ( .A1(G217), .A2(n1111), .A3(G234), .ZN(n1359) );
INV_X1 U1048 ( .A(n1200), .ZN(n1289) );
NAND3_X1 U1049 ( .A1(n1267), .A2(n1268), .A3(n1070), .ZN(n1200) );
NOR2_X1 U1050 ( .A1(n1141), .A2(n1140), .ZN(n1070) );
INV_X1 U1051 ( .A(n1286), .ZN(n1140) );
NAND2_X1 U1052 ( .A1(G214), .A2(n1362), .ZN(n1286) );
XNOR2_X1 U1053 ( .A(n1363), .B(n1241), .ZN(n1141) );
NAND2_X1 U1054 ( .A1(G210), .A2(n1362), .ZN(n1241) );
NAND2_X1 U1055 ( .A1(n1337), .A2(n1125), .ZN(n1362) );
INV_X1 U1056 ( .A(G237), .ZN(n1337) );
NAND2_X1 U1057 ( .A1(n1364), .A2(n1125), .ZN(n1363) );
XOR2_X1 U1058 ( .A(n1365), .B(n1366), .Z(n1364) );
XOR2_X1 U1059 ( .A(n1239), .B(n1367), .Z(n1366) );
XOR2_X1 U1060 ( .A(KEYINPUT16), .B(KEYINPUT15), .Z(n1367) );
AND2_X1 U1061 ( .A1(G224), .A2(n1111), .ZN(n1239) );
XOR2_X1 U1062 ( .A(n1368), .B(n1238), .Z(n1365) );
XOR2_X1 U1063 ( .A(G125), .B(n1335), .Z(n1238) );
XNOR2_X1 U1064 ( .A(n1361), .B(n1369), .ZN(n1335) );
NOR2_X1 U1065 ( .A1(G146), .A2(KEYINPUT36), .ZN(n1369) );
XNOR2_X1 U1066 ( .A(G128), .B(G143), .ZN(n1361) );
NAND2_X1 U1067 ( .A1(KEYINPUT18), .A2(n1236), .ZN(n1368) );
XNOR2_X1 U1068 ( .A(n1370), .B(n1180), .ZN(n1236) );
NAND2_X1 U1069 ( .A1(n1371), .A2(n1372), .ZN(n1180) );
NAND2_X1 U1070 ( .A1(G122), .A2(n1373), .ZN(n1372) );
XOR2_X1 U1071 ( .A(n1374), .B(KEYINPUT63), .Z(n1371) );
NAND2_X1 U1072 ( .A1(n1375), .A2(n1351), .ZN(n1374) );
INV_X1 U1073 ( .A(G122), .ZN(n1351) );
XNOR2_X1 U1074 ( .A(KEYINPUT13), .B(n1373), .ZN(n1375) );
NAND2_X1 U1075 ( .A1(n1376), .A2(n1377), .ZN(n1370) );
OR2_X1 U1076 ( .A1(n1178), .A2(n1182), .ZN(n1377) );
XOR2_X1 U1077 ( .A(n1378), .B(KEYINPUT2), .Z(n1376) );
NAND2_X1 U1078 ( .A1(n1182), .A2(n1178), .ZN(n1378) );
XOR2_X1 U1079 ( .A(n1379), .B(n1300), .Z(n1178) );
INV_X1 U1080 ( .A(G113), .ZN(n1300) );
NAND2_X1 U1081 ( .A1(n1380), .A2(KEYINPUT49), .ZN(n1379) );
XNOR2_X1 U1082 ( .A(G116), .B(G119), .ZN(n1380) );
XOR2_X1 U1083 ( .A(n1381), .B(n1382), .Z(n1182) );
NOR2_X1 U1084 ( .A1(KEYINPUT11), .A2(n1197), .ZN(n1382) );
INV_X1 U1085 ( .A(G104), .ZN(n1197) );
XNOR2_X1 U1086 ( .A(G101), .B(G107), .ZN(n1381) );
NAND2_X1 U1087 ( .A1(n1092), .A2(n1383), .ZN(n1268) );
NAND3_X1 U1088 ( .A1(n1172), .A2(n1293), .A3(G902), .ZN(n1383) );
NOR2_X1 U1089 ( .A1(n1111), .A2(G898), .ZN(n1172) );
NAND3_X1 U1090 ( .A1(n1293), .A2(n1111), .A3(G952), .ZN(n1092) );
INV_X1 U1091 ( .A(G953), .ZN(n1111) );
NAND2_X1 U1092 ( .A1(G237), .A2(G234), .ZN(n1293) );
XOR2_X1 U1093 ( .A(n1100), .B(KEYINPUT41), .Z(n1267) );
AND2_X1 U1094 ( .A1(n1102), .A2(n1101), .ZN(n1100) );
NAND2_X1 U1095 ( .A1(n1384), .A2(n1135), .ZN(n1101) );
OR2_X1 U1096 ( .A1(n1134), .A2(G469), .ZN(n1135) );
NAND2_X1 U1097 ( .A1(G469), .A2(n1134), .ZN(n1384) );
NAND2_X1 U1098 ( .A1(n1125), .A2(n1385), .ZN(n1134) );
NAND2_X1 U1099 ( .A1(n1386), .A2(n1387), .ZN(n1385) );
NAND2_X1 U1100 ( .A1(n1388), .A2(n1221), .ZN(n1387) );
XOR2_X1 U1101 ( .A(n1389), .B(KEYINPUT47), .Z(n1386) );
OR2_X1 U1102 ( .A1(n1221), .A2(n1388), .ZN(n1389) );
XOR2_X1 U1103 ( .A(n1390), .B(n1391), .Z(n1388) );
XNOR2_X1 U1104 ( .A(n1373), .B(n1227), .ZN(n1391) );
NOR2_X1 U1105 ( .A1(n1145), .A2(G953), .ZN(n1227) );
INV_X1 U1106 ( .A(G227), .ZN(n1145) );
INV_X1 U1107 ( .A(G110), .ZN(n1373) );
NAND2_X1 U1108 ( .A1(KEYINPUT53), .A2(n1392), .ZN(n1390) );
XNOR2_X1 U1109 ( .A(KEYINPUT55), .B(n1231), .ZN(n1392) );
INV_X1 U1110 ( .A(G140), .ZN(n1231) );
XNOR2_X1 U1111 ( .A(n1393), .B(n1394), .ZN(n1221) );
XOR2_X1 U1112 ( .A(G101), .B(n1395), .Z(n1394) );
NOR2_X1 U1113 ( .A1(KEYINPUT20), .A2(n1396), .ZN(n1395) );
XNOR2_X1 U1114 ( .A(n1067), .B(G104), .ZN(n1396) );
INV_X1 U1115 ( .A(G107), .ZN(n1067) );
XOR2_X1 U1116 ( .A(n1334), .B(n1160), .Z(n1393) );
AND3_X1 U1117 ( .A1(n1397), .A2(n1398), .A3(n1399), .ZN(n1160) );
NAND2_X1 U1118 ( .A1(n1400), .A2(n1401), .ZN(n1399) );
XNOR2_X1 U1119 ( .A(G143), .B(n1402), .ZN(n1400) );
NAND3_X1 U1120 ( .A1(n1402), .A2(G146), .A3(n1348), .ZN(n1398) );
OR3_X1 U1121 ( .A1(n1401), .A2(n1402), .A3(n1348), .ZN(n1397) );
INV_X1 U1122 ( .A(G143), .ZN(n1348) );
NOR2_X1 U1123 ( .A1(G128), .A2(KEYINPUT59), .ZN(n1402) );
INV_X1 U1124 ( .A(G146), .ZN(n1401) );
XOR2_X1 U1125 ( .A(n1165), .B(n1156), .Z(n1334) );
XOR2_X1 U1126 ( .A(G131), .B(KEYINPUT39), .Z(n1156) );
XNOR2_X1 U1127 ( .A(G137), .B(n1164), .ZN(n1165) );
XOR2_X1 U1128 ( .A(G134), .B(KEYINPUT19), .Z(n1164) );
NAND2_X1 U1129 ( .A1(G221), .A2(n1307), .ZN(n1102) );
NAND2_X1 U1130 ( .A1(G234), .A2(n1125), .ZN(n1307) );
INV_X1 U1131 ( .A(G902), .ZN(n1125) );
endmodule


