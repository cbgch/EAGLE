//Key = 1001100110011001001000011000110100000101100101100101101101010101


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
n1316, n1317, n1318, n1319, n1320, n1321;

XNOR2_X1 U724 ( .A(n1006), .B(n1007), .ZN(G9) );
NAND2_X1 U725 ( .A1(KEYINPUT54), .A2(G107), .ZN(n1007) );
NOR2_X1 U726 ( .A1(n1008), .A2(n1009), .ZN(G75) );
NOR4_X1 U727 ( .A1(G953), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1009) );
XOR2_X1 U728 ( .A(KEYINPUT0), .B(n1013), .Z(n1012) );
NOR2_X1 U729 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
NOR2_X1 U730 ( .A1(n1016), .A2(n1017), .ZN(n1015) );
NOR2_X1 U731 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U732 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NOR2_X1 U733 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U734 ( .A1(KEYINPUT4), .A2(n1024), .ZN(n1018) );
NOR4_X1 U735 ( .A1(n1025), .A2(n1026), .A3(n1027), .A4(n1028), .ZN(n1024) );
NOR2_X1 U736 ( .A1(n1029), .A2(n1025), .ZN(n1014) );
NOR2_X1 U737 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
NOR2_X1 U738 ( .A1(n1032), .A2(n1021), .ZN(n1031) );
NAND3_X1 U739 ( .A1(n1033), .A2(n1034), .A3(n1035), .ZN(n1021) );
INV_X1 U740 ( .A(n1028), .ZN(n1035) );
NOR2_X1 U741 ( .A1(n1036), .A2(n1037), .ZN(n1032) );
NOR2_X1 U742 ( .A1(n1038), .A2(n1039), .ZN(n1036) );
NOR3_X1 U743 ( .A1(n1028), .A2(n1040), .A3(n1041), .ZN(n1030) );
NOR4_X1 U744 ( .A1(n1017), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1041) );
NOR2_X1 U745 ( .A1(KEYINPUT56), .A2(n1045), .ZN(n1044) );
NOR2_X1 U746 ( .A1(n1046), .A2(n1027), .ZN(n1043) );
NOR2_X1 U747 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
NOR2_X1 U748 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
AND2_X1 U749 ( .A1(n1051), .A2(KEYINPUT4), .ZN(n1047) );
AND2_X1 U750 ( .A1(n1052), .A2(n1033), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1053), .A2(n1054), .ZN(n1040) );
AND2_X1 U752 ( .A1(n1055), .A2(KEYINPUT56), .ZN(n1054) );
NOR3_X1 U753 ( .A1(n1010), .A2(G953), .A3(G952), .ZN(n1008) );
AND4_X1 U754 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1010) );
NOR4_X1 U755 ( .A1(n1060), .A2(n1061), .A3(n1039), .A4(n1062), .ZN(n1059) );
XOR2_X1 U756 ( .A(n1063), .B(n1064), .Z(n1062) );
NAND2_X1 U757 ( .A1(KEYINPUT23), .A2(n1065), .ZN(n1064) );
AND2_X1 U758 ( .A1(n1038), .A2(n1050), .ZN(n1058) );
XOR2_X1 U759 ( .A(KEYINPUT12), .B(n1066), .Z(n1057) );
XOR2_X1 U760 ( .A(n1067), .B(n1068), .Z(G72) );
XOR2_X1 U761 ( .A(n1069), .B(n1070), .Z(n1068) );
NOR2_X1 U762 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U763 ( .A1(n1073), .A2(n1074), .ZN(n1071) );
XOR2_X1 U764 ( .A(KEYINPUT29), .B(G900), .Z(n1074) );
INV_X1 U765 ( .A(G227), .ZN(n1073) );
NAND2_X1 U766 ( .A1(n1075), .A2(n1076), .ZN(n1069) );
NAND2_X1 U767 ( .A1(G953), .A2(n1077), .ZN(n1076) );
XOR2_X1 U768 ( .A(n1078), .B(n1079), .Z(n1075) );
XOR2_X1 U769 ( .A(G131), .B(n1080), .Z(n1079) );
NOR2_X1 U770 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U771 ( .A(n1083), .B(KEYINPUT59), .Z(n1082) );
NAND2_X1 U772 ( .A1(n1084), .A2(n1085), .ZN(n1083) );
XNOR2_X1 U773 ( .A(G137), .B(n1086), .ZN(n1084) );
XNOR2_X1 U774 ( .A(KEYINPUT5), .B(KEYINPUT22), .ZN(n1086) );
NOR2_X1 U775 ( .A1(G137), .A2(n1085), .ZN(n1081) );
XNOR2_X1 U776 ( .A(n1087), .B(n1088), .ZN(n1078) );
NOR2_X1 U777 ( .A1(KEYINPUT33), .A2(n1089), .ZN(n1088) );
NAND2_X1 U778 ( .A1(n1072), .A2(n1090), .ZN(n1067) );
NAND2_X1 U779 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U780 ( .A(n1093), .B(n1094), .Z(G69) );
XOR2_X1 U781 ( .A(n1095), .B(n1096), .Z(n1094) );
NOR3_X1 U782 ( .A1(n1097), .A2(n1098), .A3(n1099), .ZN(n1096) );
NOR2_X1 U783 ( .A1(G898), .A2(n1072), .ZN(n1099) );
NOR2_X1 U784 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
XOR2_X1 U785 ( .A(n1102), .B(KEYINPUT46), .Z(n1097) );
NAND2_X1 U786 ( .A1(n1101), .A2(n1100), .ZN(n1102) );
XOR2_X1 U787 ( .A(n1103), .B(KEYINPUT55), .Z(n1101) );
NAND2_X1 U788 ( .A1(n1072), .A2(n1104), .ZN(n1095) );
NAND2_X1 U789 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U790 ( .A(n1107), .B(KEYINPUT41), .Z(n1105) );
NAND2_X1 U791 ( .A1(G953), .A2(n1108), .ZN(n1093) );
NAND2_X1 U792 ( .A1(G898), .A2(G224), .ZN(n1108) );
NOR2_X1 U793 ( .A1(n1109), .A2(n1110), .ZN(G66) );
XOR2_X1 U794 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U795 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
NOR2_X1 U796 ( .A1(n1109), .A2(n1115), .ZN(G63) );
XOR2_X1 U797 ( .A(n1116), .B(n1117), .Z(n1115) );
NAND3_X1 U798 ( .A1(n1118), .A2(G478), .A3(KEYINPUT39), .ZN(n1116) );
NOR2_X1 U799 ( .A1(n1109), .A2(n1119), .ZN(G60) );
XNOR2_X1 U800 ( .A(n1120), .B(n1121), .ZN(n1119) );
AND2_X1 U801 ( .A1(G475), .A2(n1118), .ZN(n1120) );
XOR2_X1 U802 ( .A(G104), .B(n1122), .Z(G6) );
NOR2_X1 U803 ( .A1(n1109), .A2(n1123), .ZN(G57) );
XOR2_X1 U804 ( .A(n1124), .B(n1125), .Z(n1123) );
XNOR2_X1 U805 ( .A(n1126), .B(n1127), .ZN(n1125) );
NOR3_X1 U806 ( .A1(n1128), .A2(KEYINPUT34), .A3(n1129), .ZN(n1127) );
XOR2_X1 U807 ( .A(KEYINPUT2), .B(n1130), .Z(n1128) );
AND2_X1 U808 ( .A1(n1131), .A2(n1132), .ZN(n1130) );
XOR2_X1 U809 ( .A(n1133), .B(n1134), .Z(n1124) );
AND2_X1 U810 ( .A1(G472), .A2(n1118), .ZN(n1134) );
INV_X1 U811 ( .A(n1114), .ZN(n1118) );
NAND2_X1 U812 ( .A1(KEYINPUT61), .A2(n1135), .ZN(n1133) );
XOR2_X1 U813 ( .A(KEYINPUT60), .B(G101), .Z(n1135) );
NOR2_X1 U814 ( .A1(n1109), .A2(n1136), .ZN(G54) );
XOR2_X1 U815 ( .A(n1137), .B(n1138), .Z(n1136) );
XOR2_X1 U816 ( .A(n1139), .B(n1140), .Z(n1138) );
XOR2_X1 U817 ( .A(n1141), .B(n1142), .Z(n1140) );
NOR2_X1 U818 ( .A1(n1063), .A2(n1114), .ZN(n1141) );
INV_X1 U819 ( .A(G469), .ZN(n1063) );
XOR2_X1 U820 ( .A(n1143), .B(n1144), .Z(n1137) );
XOR2_X1 U821 ( .A(n1085), .B(KEYINPUT36), .Z(n1144) );
NAND2_X1 U822 ( .A1(n1145), .A2(n1146), .ZN(n1143) );
OR2_X1 U823 ( .A1(n1089), .A2(n1147), .ZN(n1146) );
XOR2_X1 U824 ( .A(n1148), .B(KEYINPUT32), .Z(n1145) );
NAND2_X1 U825 ( .A1(n1147), .A2(n1089), .ZN(n1148) );
XNOR2_X1 U826 ( .A(n1149), .B(n1150), .ZN(n1089) );
NOR2_X1 U827 ( .A1(n1109), .A2(n1151), .ZN(G51) );
XOR2_X1 U828 ( .A(n1152), .B(n1153), .Z(n1151) );
XOR2_X1 U829 ( .A(G125), .B(n1154), .Z(n1153) );
NOR2_X1 U830 ( .A1(KEYINPUT53), .A2(n1155), .ZN(n1154) );
XNOR2_X1 U831 ( .A(n1156), .B(n1157), .ZN(n1152) );
NOR2_X1 U832 ( .A1(n1158), .A2(KEYINPUT14), .ZN(n1157) );
NOR2_X1 U833 ( .A1(n1159), .A2(n1114), .ZN(n1158) );
NAND2_X1 U834 ( .A1(G902), .A2(n1011), .ZN(n1114) );
NAND4_X1 U835 ( .A1(n1160), .A2(n1091), .A3(n1106), .A4(n1107), .ZN(n1011) );
NAND3_X1 U836 ( .A1(n1161), .A2(n1162), .A3(n1033), .ZN(n1107) );
AND4_X1 U837 ( .A1(n1163), .A2(n1164), .A3(n1165), .A4(n1166), .ZN(n1106) );
NOR3_X1 U838 ( .A1(n1122), .A2(n1167), .A3(n1006), .ZN(n1166) );
AND2_X1 U839 ( .A1(n1168), .A2(n1052), .ZN(n1006) );
INV_X1 U840 ( .A(n1169), .ZN(n1167) );
AND2_X1 U841 ( .A1(n1170), .A2(n1168), .ZN(n1122) );
AND3_X1 U842 ( .A1(n1051), .A2(n1171), .A3(n1162), .ZN(n1168) );
NAND3_X1 U843 ( .A1(n1162), .A2(n1172), .A3(n1023), .ZN(n1164) );
NAND2_X1 U844 ( .A1(n1045), .A2(n1173), .ZN(n1172) );
NAND2_X1 U845 ( .A1(n1034), .A2(n1051), .ZN(n1173) );
AND4_X1 U846 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1091) );
AND4_X1 U847 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1177) );
XOR2_X1 U848 ( .A(n1092), .B(KEYINPUT48), .Z(n1160) );
NOR2_X1 U849 ( .A1(n1072), .A2(G952), .ZN(n1109) );
XNOR2_X1 U850 ( .A(G146), .B(n1176), .ZN(G48) );
NAND2_X1 U851 ( .A1(n1182), .A2(n1170), .ZN(n1176) );
XOR2_X1 U852 ( .A(n1183), .B(n1184), .Z(G45) );
XOR2_X1 U853 ( .A(KEYINPUT16), .B(G143), .Z(n1184) );
NAND2_X1 U854 ( .A1(n1185), .A2(n1186), .ZN(n1183) );
NAND3_X1 U855 ( .A1(n1187), .A2(n1188), .A3(n1189), .ZN(n1186) );
OR2_X1 U856 ( .A1(n1178), .A2(n1189), .ZN(n1185) );
INV_X1 U857 ( .A(KEYINPUT3), .ZN(n1189) );
NAND2_X1 U858 ( .A1(n1187), .A2(n1037), .ZN(n1178) );
AND4_X1 U859 ( .A1(n1066), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1187) );
NOR2_X1 U860 ( .A1(n1026), .A2(n1193), .ZN(n1192) );
XNOR2_X1 U861 ( .A(G140), .B(n1174), .ZN(G42) );
NAND3_X1 U862 ( .A1(n1022), .A2(n1170), .A3(n1194), .ZN(n1174) );
XNOR2_X1 U863 ( .A(G137), .B(n1092), .ZN(G39) );
NAND2_X1 U864 ( .A1(n1194), .A2(n1161), .ZN(n1092) );
XOR2_X1 U865 ( .A(n1085), .B(n1175), .Z(G36) );
NAND3_X1 U866 ( .A1(n1023), .A2(n1052), .A3(n1194), .ZN(n1175) );
INV_X1 U867 ( .A(G134), .ZN(n1085) );
XNOR2_X1 U868 ( .A(G131), .B(n1181), .ZN(G33) );
NAND3_X1 U869 ( .A1(n1170), .A2(n1023), .A3(n1194), .ZN(n1181) );
NOR3_X1 U870 ( .A1(n1026), .A2(n1195), .A3(n1017), .ZN(n1194) );
INV_X1 U871 ( .A(n1053), .ZN(n1017) );
NOR2_X1 U872 ( .A1(n1039), .A2(n1196), .ZN(n1053) );
XOR2_X1 U873 ( .A(KEYINPUT43), .B(n1038), .Z(n1196) );
XOR2_X1 U874 ( .A(n1180), .B(n1197), .Z(G30) );
NAND2_X1 U875 ( .A1(KEYINPUT31), .A2(G128), .ZN(n1197) );
NAND2_X1 U876 ( .A1(n1182), .A2(n1052), .ZN(n1180) );
AND3_X1 U877 ( .A1(n1051), .A2(n1037), .A3(n1198), .ZN(n1182) );
NOR3_X1 U878 ( .A1(n1199), .A2(n1195), .A3(n1056), .ZN(n1198) );
INV_X1 U879 ( .A(n1190), .ZN(n1195) );
XOR2_X1 U880 ( .A(n1200), .B(n1201), .Z(G3) );
NAND4_X1 U881 ( .A1(n1023), .A2(n1034), .A3(n1162), .A4(n1202), .ZN(n1201) );
XOR2_X1 U882 ( .A(KEYINPUT30), .B(n1051), .Z(n1202) );
XOR2_X1 U883 ( .A(n1203), .B(n1179), .Z(G27) );
NAND4_X1 U884 ( .A1(n1055), .A2(n1022), .A3(n1037), .A4(n1190), .ZN(n1179) );
NAND2_X1 U885 ( .A1(n1028), .A2(n1204), .ZN(n1190) );
NAND4_X1 U886 ( .A1(G953), .A2(G902), .A3(n1205), .A4(n1077), .ZN(n1204) );
INV_X1 U887 ( .A(G900), .ZN(n1077) );
XOR2_X1 U888 ( .A(n1206), .B(n1169), .Z(G24) );
NAND4_X1 U889 ( .A1(n1033), .A2(n1162), .A3(n1207), .A4(n1171), .ZN(n1169) );
INV_X1 U890 ( .A(n1025), .ZN(n1171) );
NAND2_X1 U891 ( .A1(n1208), .A2(n1199), .ZN(n1025) );
AND2_X1 U892 ( .A1(n1066), .A2(n1191), .ZN(n1207) );
XNOR2_X1 U893 ( .A(n1209), .B(KEYINPUT9), .ZN(n1191) );
XOR2_X1 U894 ( .A(n1210), .B(n1211), .Z(G21) );
NAND2_X1 U895 ( .A1(KEYINPUT51), .A2(G119), .ZN(n1211) );
NAND3_X1 U896 ( .A1(n1161), .A2(n1162), .A3(n1212), .ZN(n1210) );
XNOR2_X1 U897 ( .A(n1033), .B(KEYINPUT40), .ZN(n1212) );
NOR3_X1 U898 ( .A1(n1199), .A2(n1056), .A3(n1027), .ZN(n1161) );
XOR2_X1 U899 ( .A(n1213), .B(n1165), .Z(G18) );
NAND4_X1 U900 ( .A1(n1023), .A2(n1033), .A3(n1052), .A4(n1162), .ZN(n1165) );
NOR2_X1 U901 ( .A1(n1066), .A2(n1209), .ZN(n1052) );
INV_X1 U902 ( .A(n1214), .ZN(n1066) );
XOR2_X1 U903 ( .A(n1215), .B(n1216), .Z(G15) );
NAND3_X1 U904 ( .A1(n1162), .A2(n1217), .A3(n1055), .ZN(n1216) );
INV_X1 U905 ( .A(n1045), .ZN(n1055) );
NAND2_X1 U906 ( .A1(n1170), .A2(n1033), .ZN(n1045) );
NOR2_X1 U907 ( .A1(n1049), .A2(n1218), .ZN(n1033) );
INV_X1 U908 ( .A(n1050), .ZN(n1218) );
NOR2_X1 U909 ( .A1(n1060), .A2(n1214), .ZN(n1170) );
INV_X1 U910 ( .A(n1209), .ZN(n1060) );
XOR2_X1 U911 ( .A(KEYINPUT50), .B(n1023), .Z(n1217) );
INV_X1 U912 ( .A(n1193), .ZN(n1023) );
NAND2_X1 U913 ( .A1(n1208), .A2(n1061), .ZN(n1193) );
XOR2_X1 U914 ( .A(n1056), .B(KEYINPUT47), .Z(n1208) );
XNOR2_X1 U915 ( .A(G110), .B(n1163), .ZN(G12) );
NAND4_X1 U916 ( .A1(n1022), .A2(n1034), .A3(n1162), .A4(n1051), .ZN(n1163) );
INV_X1 U917 ( .A(n1026), .ZN(n1051) );
NAND2_X1 U918 ( .A1(n1049), .A2(n1050), .ZN(n1026) );
NAND2_X1 U919 ( .A1(G221), .A2(n1219), .ZN(n1050) );
XNOR2_X1 U920 ( .A(n1065), .B(n1220), .ZN(n1049) );
XOR2_X1 U921 ( .A(KEYINPUT11), .B(G469), .Z(n1220) );
AND2_X1 U922 ( .A1(n1221), .A2(n1222), .ZN(n1065) );
XOR2_X1 U923 ( .A(n1223), .B(n1224), .Z(n1221) );
XOR2_X1 U924 ( .A(n1149), .B(n1225), .Z(n1224) );
NAND2_X1 U925 ( .A1(KEYINPUT7), .A2(n1147), .ZN(n1225) );
XOR2_X1 U926 ( .A(n1226), .B(n1227), .Z(n1147) );
XOR2_X1 U927 ( .A(G107), .B(G101), .Z(n1227) );
NAND2_X1 U928 ( .A1(KEYINPUT63), .A2(n1228), .ZN(n1226) );
INV_X1 U929 ( .A(G104), .ZN(n1228) );
XOR2_X1 U930 ( .A(n1229), .B(n1139), .Z(n1223) );
XNOR2_X1 U931 ( .A(n1230), .B(n1231), .ZN(n1139) );
XOR2_X1 U932 ( .A(G140), .B(G110), .Z(n1231) );
NAND2_X1 U933 ( .A1(G227), .A2(n1232), .ZN(n1230) );
AND2_X1 U934 ( .A1(n1037), .A2(n1233), .ZN(n1162) );
NAND2_X1 U935 ( .A1(n1234), .A2(n1028), .ZN(n1233) );
NAND3_X1 U936 ( .A1(n1205), .A2(n1072), .A3(G952), .ZN(n1028) );
NAND4_X1 U937 ( .A1(G953), .A2(G902), .A3(n1205), .A4(n1235), .ZN(n1234) );
INV_X1 U938 ( .A(G898), .ZN(n1235) );
NAND2_X1 U939 ( .A1(G237), .A2(n1236), .ZN(n1205) );
INV_X1 U940 ( .A(n1188), .ZN(n1037) );
NAND2_X1 U941 ( .A1(n1237), .A2(n1039), .ZN(n1188) );
XOR2_X1 U942 ( .A(n1238), .B(n1159), .Z(n1039) );
NAND2_X1 U943 ( .A1(G210), .A2(n1239), .ZN(n1159) );
NAND3_X1 U944 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1238) );
XOR2_X1 U945 ( .A(n1222), .B(KEYINPUT44), .Z(n1242) );
NAND2_X1 U946 ( .A1(n1243), .A2(n1155), .ZN(n1241) );
XOR2_X1 U947 ( .A(n1244), .B(KEYINPUT24), .Z(n1243) );
NAND2_X1 U948 ( .A1(n1245), .A2(n1246), .ZN(n1240) );
INV_X1 U949 ( .A(n1155), .ZN(n1246) );
XOR2_X1 U950 ( .A(n1247), .B(n1150), .Z(n1155) );
XOR2_X1 U951 ( .A(G128), .B(G146), .Z(n1150) );
XOR2_X1 U952 ( .A(n1244), .B(n1248), .Z(n1245) );
XNOR2_X1 U953 ( .A(KEYINPUT28), .B(KEYINPUT13), .ZN(n1248) );
XOR2_X1 U954 ( .A(n1203), .B(n1156), .Z(n1244) );
XNOR2_X1 U955 ( .A(n1249), .B(n1250), .ZN(n1156) );
INV_X1 U956 ( .A(n1103), .ZN(n1250) );
XOR2_X1 U957 ( .A(n1251), .B(n1252), .Z(n1103) );
XOR2_X1 U958 ( .A(G113), .B(G101), .Z(n1252) );
XNOR2_X1 U959 ( .A(n1253), .B(n1254), .ZN(n1251) );
NOR2_X1 U960 ( .A1(KEYINPUT6), .A2(n1255), .ZN(n1254) );
NOR2_X1 U961 ( .A1(KEYINPUT17), .A2(n1256), .ZN(n1253) );
XOR2_X1 U962 ( .A(G104), .B(n1257), .Z(n1256) );
NOR2_X1 U963 ( .A1(G107), .A2(KEYINPUT21), .ZN(n1257) );
XNOR2_X1 U964 ( .A(n1258), .B(n1100), .ZN(n1249) );
XOR2_X1 U965 ( .A(G110), .B(n1206), .Z(n1100) );
INV_X1 U966 ( .A(G122), .ZN(n1206) );
NAND2_X1 U967 ( .A1(G224), .A2(n1232), .ZN(n1258) );
INV_X1 U968 ( .A(G125), .ZN(n1203) );
XNOR2_X1 U969 ( .A(KEYINPUT43), .B(n1038), .ZN(n1237) );
NAND2_X1 U970 ( .A1(G214), .A2(n1239), .ZN(n1038) );
NAND2_X1 U971 ( .A1(n1259), .A2(n1222), .ZN(n1239) );
INV_X1 U972 ( .A(n1027), .ZN(n1034) );
NAND2_X1 U973 ( .A1(n1209), .A2(n1214), .ZN(n1027) );
XOR2_X1 U974 ( .A(n1260), .B(G475), .Z(n1214) );
NAND2_X1 U975 ( .A1(n1261), .A2(n1121), .ZN(n1260) );
XOR2_X1 U976 ( .A(n1262), .B(n1263), .Z(n1121) );
XOR2_X1 U977 ( .A(G104), .B(n1264), .Z(n1263) );
NOR2_X1 U978 ( .A1(KEYINPUT19), .A2(n1265), .ZN(n1264) );
XOR2_X1 U979 ( .A(n1215), .B(n1266), .Z(n1265) );
XOR2_X1 U980 ( .A(KEYINPUT10), .B(G122), .Z(n1266) );
NAND2_X1 U981 ( .A1(n1267), .A2(KEYINPUT45), .ZN(n1262) );
XOR2_X1 U982 ( .A(n1268), .B(n1269), .Z(n1267) );
XOR2_X1 U983 ( .A(n1270), .B(n1271), .Z(n1269) );
NOR2_X1 U984 ( .A1(G125), .A2(KEYINPUT38), .ZN(n1271) );
NOR2_X1 U985 ( .A1(n1272), .A2(n1273), .ZN(n1270) );
XOR2_X1 U986 ( .A(n1274), .B(KEYINPUT18), .Z(n1273) );
NAND2_X1 U987 ( .A1(G131), .A2(n1275), .ZN(n1274) );
NOR2_X1 U988 ( .A1(G131), .A2(n1275), .ZN(n1272) );
NAND2_X1 U989 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
NAND4_X1 U990 ( .A1(G143), .A2(G214), .A3(n1232), .A4(n1259), .ZN(n1277) );
XOR2_X1 U991 ( .A(n1278), .B(KEYINPUT20), .Z(n1276) );
NAND2_X1 U992 ( .A1(n1149), .A2(n1279), .ZN(n1278) );
NAND3_X1 U993 ( .A1(n1232), .A2(n1259), .A3(G214), .ZN(n1279) );
XNOR2_X1 U994 ( .A(G140), .B(n1280), .ZN(n1268) );
XOR2_X1 U995 ( .A(KEYINPUT42), .B(G146), .Z(n1280) );
XOR2_X1 U996 ( .A(n1222), .B(KEYINPUT35), .Z(n1261) );
XOR2_X1 U997 ( .A(n1281), .B(G478), .Z(n1209) );
NAND2_X1 U998 ( .A1(n1117), .A2(n1222), .ZN(n1281) );
XOR2_X1 U999 ( .A(n1282), .B(n1283), .Z(n1117) );
XOR2_X1 U1000 ( .A(n1284), .B(n1285), .Z(n1283) );
XNOR2_X1 U1001 ( .A(n1286), .B(n1287), .ZN(n1285) );
NOR4_X1 U1002 ( .A1(KEYINPUT58), .A2(n1288), .A3(n1289), .A4(n1113), .ZN(n1287) );
NAND2_X1 U1003 ( .A1(KEYINPUT15), .A2(n1213), .ZN(n1286) );
INV_X1 U1004 ( .A(G116), .ZN(n1213) );
XNOR2_X1 U1005 ( .A(G107), .B(n1290), .ZN(n1282) );
XOR2_X1 U1006 ( .A(G143), .B(G122), .Z(n1290) );
NOR2_X1 U1007 ( .A1(n1061), .A2(n1056), .ZN(n1022) );
XOR2_X1 U1008 ( .A(n1291), .B(n1292), .Z(n1056) );
NOR2_X1 U1009 ( .A1(n1113), .A2(n1293), .ZN(n1292) );
XNOR2_X1 U1010 ( .A(KEYINPUT62), .B(n1219), .ZN(n1293) );
NAND2_X1 U1011 ( .A1(n1236), .A2(n1222), .ZN(n1219) );
XOR2_X1 U1012 ( .A(n1289), .B(KEYINPUT57), .Z(n1236) );
INV_X1 U1013 ( .A(G234), .ZN(n1289) );
INV_X1 U1014 ( .A(G217), .ZN(n1113) );
OR2_X1 U1015 ( .A1(n1112), .A2(G902), .ZN(n1291) );
XNOR2_X1 U1016 ( .A(n1294), .B(n1295), .ZN(n1112) );
XOR2_X1 U1017 ( .A(n1296), .B(n1297), .Z(n1295) );
NAND2_X1 U1018 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
NAND2_X1 U1019 ( .A1(G137), .A2(n1300), .ZN(n1299) );
XOR2_X1 U1020 ( .A(n1301), .B(n1302), .Z(n1298) );
NOR2_X1 U1021 ( .A1(G137), .A2(n1300), .ZN(n1302) );
INV_X1 U1022 ( .A(KEYINPUT49), .ZN(n1300) );
NAND3_X1 U1023 ( .A1(G234), .A2(n1232), .A3(G221), .ZN(n1301) );
NAND3_X1 U1024 ( .A1(n1303), .A2(n1304), .A3(n1305), .ZN(n1296) );
NAND2_X1 U1025 ( .A1(KEYINPUT25), .A2(n1306), .ZN(n1305) );
NAND3_X1 U1026 ( .A1(n1307), .A2(n1308), .A3(n1087), .ZN(n1304) );
INV_X1 U1027 ( .A(KEYINPUT25), .ZN(n1308) );
OR2_X1 U1028 ( .A1(n1087), .A2(n1307), .ZN(n1303) );
NOR2_X1 U1029 ( .A1(KEYINPUT26), .A2(n1306), .ZN(n1307) );
XOR2_X1 U1030 ( .A(G146), .B(KEYINPUT1), .Z(n1306) );
XOR2_X1 U1031 ( .A(G125), .B(G140), .Z(n1087) );
XNOR2_X1 U1032 ( .A(G110), .B(n1309), .ZN(n1294) );
XOR2_X1 U1033 ( .A(G128), .B(G119), .Z(n1309) );
INV_X1 U1034 ( .A(n1199), .ZN(n1061) );
XOR2_X1 U1035 ( .A(n1310), .B(G472), .Z(n1199) );
NAND2_X1 U1036 ( .A1(n1311), .A2(n1222), .ZN(n1310) );
INV_X1 U1037 ( .A(G902), .ZN(n1222) );
XOR2_X1 U1038 ( .A(n1126), .B(n1312), .Z(n1311) );
NAND2_X1 U1039 ( .A1(n1313), .A2(n1314), .ZN(n1312) );
NAND2_X1 U1040 ( .A1(n1315), .A2(n1200), .ZN(n1314) );
INV_X1 U1041 ( .A(G101), .ZN(n1200) );
NAND2_X1 U1042 ( .A1(n1316), .A2(n1317), .ZN(n1315) );
NAND2_X1 U1043 ( .A1(n1132), .A2(n1131), .ZN(n1317) );
INV_X1 U1044 ( .A(n1129), .ZN(n1316) );
NOR2_X1 U1045 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
NAND2_X1 U1046 ( .A1(n1318), .A2(G101), .ZN(n1313) );
XOR2_X1 U1047 ( .A(n1132), .B(n1131), .Z(n1318) );
XNOR2_X1 U1048 ( .A(n1215), .B(n1255), .ZN(n1131) );
XNOR2_X1 U1049 ( .A(G116), .B(G119), .ZN(n1255) );
INV_X1 U1050 ( .A(G113), .ZN(n1215) );
XNOR2_X1 U1051 ( .A(n1229), .B(n1247), .ZN(n1132) );
NAND2_X1 U1052 ( .A1(KEYINPUT37), .A2(n1149), .ZN(n1247) );
INV_X1 U1053 ( .A(G143), .ZN(n1149) );
XOR2_X1 U1054 ( .A(n1319), .B(n1142), .Z(n1229) );
XOR2_X1 U1055 ( .A(G131), .B(n1320), .Z(n1142) );
XOR2_X1 U1056 ( .A(KEYINPUT52), .B(G137), .Z(n1320) );
XNOR2_X1 U1057 ( .A(G146), .B(n1284), .ZN(n1319) );
XOR2_X1 U1058 ( .A(G128), .B(G134), .Z(n1284) );
NAND3_X1 U1059 ( .A1(n1321), .A2(n1259), .A3(G210), .ZN(n1126) );
INV_X1 U1060 ( .A(G237), .ZN(n1259) );
XOR2_X1 U1061 ( .A(KEYINPUT27), .B(n1232), .Z(n1321) );
INV_X1 U1062 ( .A(n1288), .ZN(n1232) );
XOR2_X1 U1063 ( .A(n1072), .B(KEYINPUT8), .Z(n1288) );
INV_X1 U1064 ( .A(G953), .ZN(n1072) );
endmodule


