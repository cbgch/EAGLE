//Key = 1111101010111111100011000110100111101110111110001111000011011000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273;

NAND2_X1 U717 ( .A1(n978), .A2(n979), .ZN(G9) );
NAND4_X1 U718 ( .A1(KEYINPUT14), .A2(n980), .A3(n981), .A4(n982), .ZN(n979) );
NAND3_X1 U719 ( .A1(n983), .A2(n984), .A3(n985), .ZN(n978) );
NAND2_X1 U720 ( .A1(n980), .A2(n981), .ZN(n985) );
XNOR2_X1 U721 ( .A(n986), .B(KEYINPUT5), .ZN(n981) );
NAND3_X1 U722 ( .A1(KEYINPUT1), .A2(KEYINPUT14), .A3(n982), .ZN(n984) );
OR2_X1 U723 ( .A1(n982), .A2(KEYINPUT1), .ZN(n983) );
NOR2_X1 U724 ( .A1(n987), .A2(n988), .ZN(G75) );
NOR4_X1 U725 ( .A1(n989), .A2(n990), .A3(G953), .A4(n991), .ZN(n988) );
NOR3_X1 U726 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n990) );
NOR2_X1 U727 ( .A1(n995), .A2(n980), .ZN(n993) );
NOR2_X1 U728 ( .A1(n996), .A2(n997), .ZN(n995) );
NAND3_X1 U729 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n989) );
NAND2_X1 U730 ( .A1(n1001), .A2(n1002), .ZN(n999) );
NAND3_X1 U731 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n1002) );
XOR2_X1 U732 ( .A(KEYINPUT41), .B(n1006), .Z(n1005) );
AND3_X1 U733 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n1006) );
NAND3_X1 U734 ( .A1(n1010), .A2(n1011), .A3(n1012), .ZN(n1004) );
NAND2_X1 U735 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NAND2_X1 U736 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
NAND2_X1 U737 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NAND2_X1 U738 ( .A1(KEYINPUT6), .A2(n1019), .ZN(n1018) );
NAND2_X1 U739 ( .A1(n1020), .A2(n1021), .ZN(n1013) );
NAND2_X1 U740 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NAND2_X1 U741 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
INV_X1 U742 ( .A(n1026), .ZN(n1022) );
NAND2_X1 U743 ( .A1(n1027), .A2(n1028), .ZN(n1003) );
INV_X1 U744 ( .A(KEYINPUT6), .ZN(n1028) );
NAND4_X1 U745 ( .A1(n1012), .A2(n1010), .A3(n1015), .A4(n1019), .ZN(n1027) );
XOR2_X1 U746 ( .A(KEYINPUT20), .B(n1029), .Z(n998) );
AND3_X1 U747 ( .A1(n1008), .A2(n1030), .A3(n1001), .ZN(n1029) );
INV_X1 U748 ( .A(n992), .ZN(n1008) );
NAND3_X1 U749 ( .A1(n1020), .A2(n1015), .A3(n1012), .ZN(n992) );
INV_X1 U750 ( .A(n1031), .ZN(n1012) );
NOR3_X1 U751 ( .A1(n991), .A2(G953), .A3(G952), .ZN(n987) );
AND4_X1 U752 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n991) );
NOR4_X1 U753 ( .A1(n1007), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1035) );
XOR2_X1 U754 ( .A(n996), .B(KEYINPUT38), .Z(n1038) );
XOR2_X1 U755 ( .A(n1039), .B(n1040), .Z(n1037) );
NOR2_X1 U756 ( .A1(KEYINPUT7), .A2(n1041), .ZN(n1040) );
NOR2_X1 U757 ( .A1(n1042), .A2(n1043), .ZN(n1036) );
AND2_X1 U758 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
NOR2_X1 U759 ( .A1(n1046), .A2(n1047), .ZN(n1034) );
XOR2_X1 U760 ( .A(n1048), .B(n1049), .Z(n1033) );
XOR2_X1 U761 ( .A(n1009), .B(KEYINPUT45), .Z(n1032) );
XOR2_X1 U762 ( .A(n1050), .B(n1051), .Z(G72) );
XOR2_X1 U763 ( .A(n1052), .B(n1053), .Z(n1051) );
NOR2_X1 U764 ( .A1(n1054), .A2(n1055), .ZN(n1053) );
NOR2_X1 U765 ( .A1(n1056), .A2(n1057), .ZN(n1054) );
NAND2_X1 U766 ( .A1(n1058), .A2(n1059), .ZN(n1052) );
NAND2_X1 U767 ( .A1(G953), .A2(n1057), .ZN(n1059) );
XOR2_X1 U768 ( .A(n1060), .B(n1061), .Z(n1058) );
XNOR2_X1 U769 ( .A(G131), .B(n1062), .ZN(n1061) );
NAND2_X1 U770 ( .A1(KEYINPUT21), .A2(n1063), .ZN(n1062) );
XNOR2_X1 U771 ( .A(n1064), .B(n1065), .ZN(n1060) );
INV_X1 U772 ( .A(n1066), .ZN(n1065) );
NAND2_X1 U773 ( .A1(KEYINPUT25), .A2(n1067), .ZN(n1064) );
NAND2_X1 U774 ( .A1(n1055), .A2(n1068), .ZN(n1050) );
XOR2_X1 U775 ( .A(n1069), .B(n1070), .Z(G69) );
XOR2_X1 U776 ( .A(n1071), .B(n1072), .Z(n1070) );
NAND2_X1 U777 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
NAND2_X1 U778 ( .A1(n1075), .A2(G953), .ZN(n1074) );
XNOR2_X1 U779 ( .A(n1076), .B(n1077), .ZN(n1073) );
NAND2_X1 U780 ( .A1(KEYINPUT36), .A2(n1078), .ZN(n1071) );
NAND2_X1 U781 ( .A1(G953), .A2(n1079), .ZN(n1078) );
NAND2_X1 U782 ( .A1(n1080), .A2(G224), .ZN(n1079) );
XNOR2_X1 U783 ( .A(G898), .B(KEYINPUT56), .ZN(n1080) );
NAND3_X1 U784 ( .A1(n1081), .A2(n1055), .A3(KEYINPUT8), .ZN(n1069) );
NOR2_X1 U785 ( .A1(n1082), .A2(n1083), .ZN(G66) );
XOR2_X1 U786 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR2_X1 U787 ( .A1(KEYINPUT62), .A2(n1086), .ZN(n1085) );
NAND3_X1 U788 ( .A1(G902), .A2(n1087), .A3(n1088), .ZN(n1084) );
XNOR2_X1 U789 ( .A(n1000), .B(KEYINPUT23), .ZN(n1088) );
NOR2_X1 U790 ( .A1(n1089), .A2(n1090), .ZN(G63) );
XOR2_X1 U791 ( .A(n1091), .B(n1092), .Z(n1090) );
NAND2_X1 U792 ( .A1(n1093), .A2(G478), .ZN(n1091) );
NOR2_X1 U793 ( .A1(n1055), .A2(n1094), .ZN(n1089) );
XOR2_X1 U794 ( .A(KEYINPUT9), .B(G952), .Z(n1094) );
NOR2_X1 U795 ( .A1(n1082), .A2(n1095), .ZN(G60) );
XOR2_X1 U796 ( .A(n1096), .B(n1097), .Z(n1095) );
NAND2_X1 U797 ( .A1(n1093), .A2(G475), .ZN(n1096) );
XOR2_X1 U798 ( .A(G104), .B(n1098), .Z(G6) );
NOR4_X1 U799 ( .A1(KEYINPUT63), .A2(n1099), .A3(n1017), .A4(n1100), .ZN(n1098) );
INV_X1 U800 ( .A(n1015), .ZN(n1099) );
NOR2_X1 U801 ( .A1(n1082), .A2(n1101), .ZN(G57) );
XOR2_X1 U802 ( .A(n1102), .B(n1103), .Z(n1101) );
NOR2_X1 U803 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
NOR4_X1 U804 ( .A1(n1106), .A2(n1107), .A3(n1000), .A4(n1108), .ZN(n1105) );
NOR2_X1 U805 ( .A1(KEYINPUT39), .A2(n1093), .ZN(n1108) );
INV_X1 U806 ( .A(n1109), .ZN(n1106) );
NOR2_X1 U807 ( .A1(n1110), .A2(n1109), .ZN(n1104) );
XNOR2_X1 U808 ( .A(n1111), .B(n1112), .ZN(n1109) );
NOR3_X1 U809 ( .A1(n1107), .A2(n1000), .A3(n1113), .ZN(n1110) );
NOR2_X1 U810 ( .A1(KEYINPUT39), .A2(G902), .ZN(n1113) );
NAND2_X1 U811 ( .A1(G472), .A2(n1114), .ZN(n1107) );
NAND2_X1 U812 ( .A1(KEYINPUT39), .A2(G902), .ZN(n1114) );
XNOR2_X1 U813 ( .A(n1115), .B(n1116), .ZN(n1102) );
INV_X1 U814 ( .A(G101), .ZN(n1116) );
NAND2_X1 U815 ( .A1(KEYINPUT40), .A2(n1117), .ZN(n1115) );
NOR3_X1 U816 ( .A1(n1118), .A2(n1119), .A3(n1120), .ZN(G54) );
AND3_X1 U817 ( .A1(KEYINPUT17), .A2(G953), .A3(G952), .ZN(n1120) );
NOR2_X1 U818 ( .A1(KEYINPUT17), .A2(n1121), .ZN(n1119) );
INV_X1 U819 ( .A(n1082), .ZN(n1121) );
XOR2_X1 U820 ( .A(n1122), .B(n1123), .Z(n1118) );
XNOR2_X1 U821 ( .A(n1124), .B(n1125), .ZN(n1123) );
XNOR2_X1 U822 ( .A(n1066), .B(n1126), .ZN(n1125) );
XNOR2_X1 U823 ( .A(n1127), .B(n1128), .ZN(n1122) );
XOR2_X1 U824 ( .A(n1129), .B(n1130), .Z(n1128) );
NAND2_X1 U825 ( .A1(KEYINPUT13), .A2(n1131), .ZN(n1130) );
NAND2_X1 U826 ( .A1(n1093), .A2(G469), .ZN(n1129) );
NOR2_X1 U827 ( .A1(n1082), .A2(n1132), .ZN(G51) );
XOR2_X1 U828 ( .A(n1133), .B(n1134), .Z(n1132) );
XOR2_X1 U829 ( .A(n1135), .B(n1136), .Z(n1133) );
NAND2_X1 U830 ( .A1(n1093), .A2(G210), .ZN(n1135) );
NOR2_X1 U831 ( .A1(n1137), .A2(n1000), .ZN(n1093) );
NOR2_X1 U832 ( .A1(n1068), .A2(n1081), .ZN(n1000) );
NAND4_X1 U833 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1081) );
AND4_X1 U834 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1141) );
NAND2_X1 U835 ( .A1(n980), .A2(n1146), .ZN(n1140) );
NAND2_X1 U836 ( .A1(n1147), .A2(n986), .ZN(n1146) );
NAND4_X1 U837 ( .A1(n1030), .A2(n1015), .A3(n1019), .A4(n1148), .ZN(n986) );
XOR2_X1 U838 ( .A(n1149), .B(KEYINPUT18), .Z(n1147) );
NAND3_X1 U839 ( .A1(n1150), .A2(n1015), .A3(n1151), .ZN(n1138) );
NAND4_X1 U840 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1068) );
NOR4_X1 U841 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
NAND2_X1 U842 ( .A1(n1019), .A2(n1160), .ZN(n1154) );
NAND2_X1 U843 ( .A1(n1161), .A2(n1162), .ZN(n1160) );
NAND2_X1 U844 ( .A1(n1163), .A2(n1001), .ZN(n1162) );
NAND2_X1 U845 ( .A1(n1164), .A2(n980), .ZN(n1161) );
NOR2_X1 U846 ( .A1(n1055), .A2(G952), .ZN(n1082) );
XNOR2_X1 U847 ( .A(G146), .B(n1152), .ZN(G48) );
NAND3_X1 U848 ( .A1(n1150), .A2(n980), .A3(n1164), .ZN(n1152) );
XNOR2_X1 U849 ( .A(G143), .B(n1153), .ZN(G45) );
NAND4_X1 U850 ( .A1(n1165), .A2(n1163), .A3(n980), .A4(n1046), .ZN(n1153) );
XOR2_X1 U851 ( .A(n1158), .B(n1166), .Z(G42) );
XOR2_X1 U852 ( .A(KEYINPUT24), .B(G140), .Z(n1166) );
AND3_X1 U853 ( .A1(n1167), .A2(n1030), .A3(n1001), .ZN(n1158) );
XOR2_X1 U854 ( .A(G137), .B(n1157), .Z(G39) );
AND3_X1 U855 ( .A1(n1001), .A2(n1164), .A3(n1020), .ZN(n1157) );
INV_X1 U856 ( .A(n1168), .ZN(n1164) );
XNOR2_X1 U857 ( .A(G134), .B(n1169), .ZN(G36) );
NAND4_X1 U858 ( .A1(KEYINPUT3), .A2(n1163), .A3(n1001), .A4(n1019), .ZN(n1169) );
XNOR2_X1 U859 ( .A(n1170), .B(n1159), .ZN(G33) );
AND3_X1 U860 ( .A1(n1001), .A2(n1150), .A3(n1163), .ZN(n1159) );
AND3_X1 U861 ( .A1(n1030), .A2(n1171), .A3(n1026), .ZN(n1163) );
NOR2_X1 U862 ( .A1(n997), .A2(n1172), .ZN(n1001) );
INV_X1 U863 ( .A(n996), .ZN(n1172) );
XOR2_X1 U864 ( .A(G128), .B(n1173), .Z(G30) );
NOR4_X1 U865 ( .A1(KEYINPUT29), .A2(n1174), .A3(n1175), .A4(n1168), .ZN(n1173) );
NAND4_X1 U866 ( .A1(n1030), .A2(n1176), .A3(n1025), .A4(n1171), .ZN(n1168) );
XNOR2_X1 U867 ( .A(G101), .B(n1139), .ZN(G3) );
NAND3_X1 U868 ( .A1(n1026), .A2(n1020), .A3(n1151), .ZN(n1139) );
XOR2_X1 U869 ( .A(G125), .B(n1156), .Z(G27) );
AND3_X1 U870 ( .A1(n1010), .A2(n980), .A3(n1167), .ZN(n1156) );
AND4_X1 U871 ( .A1(n1024), .A2(n1150), .A3(n1025), .A4(n1171), .ZN(n1167) );
NAND2_X1 U872 ( .A1(n1031), .A2(n1177), .ZN(n1171) );
NAND4_X1 U873 ( .A1(G953), .A2(G902), .A3(n1178), .A4(n1057), .ZN(n1177) );
INV_X1 U874 ( .A(G900), .ZN(n1057) );
XNOR2_X1 U875 ( .A(G122), .B(n1145), .ZN(G24) );
NAND4_X1 U876 ( .A1(n1165), .A2(n1179), .A3(n1015), .A4(n1046), .ZN(n1145) );
NOR2_X1 U877 ( .A1(n1025), .A2(n1176), .ZN(n1015) );
XNOR2_X1 U878 ( .A(G119), .B(n1144), .ZN(G21) );
NAND4_X1 U879 ( .A1(n1179), .A2(n1020), .A3(n1176), .A4(n1025), .ZN(n1144) );
XOR2_X1 U880 ( .A(G116), .B(n1180), .Z(G18) );
NOR2_X1 U881 ( .A1(n1175), .A2(n1149), .ZN(n1180) );
NAND4_X1 U882 ( .A1(n1026), .A2(n1010), .A3(n1019), .A4(n1148), .ZN(n1149) );
INV_X1 U883 ( .A(n1174), .ZN(n1019) );
NAND2_X1 U884 ( .A1(n1046), .A2(n1181), .ZN(n1174) );
XNOR2_X1 U885 ( .A(G113), .B(n1143), .ZN(G15) );
NAND3_X1 U886 ( .A1(n1026), .A2(n1150), .A3(n1179), .ZN(n1143) );
AND3_X1 U887 ( .A1(n980), .A2(n1148), .A3(n1010), .ZN(n1179) );
INV_X1 U888 ( .A(n994), .ZN(n1010) );
NAND2_X1 U889 ( .A1(n1009), .A2(n1182), .ZN(n994) );
INV_X1 U890 ( .A(n1017), .ZN(n1150) );
NAND2_X1 U891 ( .A1(n1165), .A2(n1183), .ZN(n1017) );
XOR2_X1 U892 ( .A(n1181), .B(KEYINPUT4), .Z(n1165) );
NOR2_X1 U893 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
XNOR2_X1 U894 ( .A(G110), .B(n1142), .ZN(G12) );
NAND4_X1 U895 ( .A1(n1151), .A2(n1020), .A3(n1024), .A4(n1025), .ZN(n1142) );
XOR2_X1 U896 ( .A(n1047), .B(KEYINPUT22), .Z(n1025) );
XNOR2_X1 U897 ( .A(n1184), .B(n1087), .ZN(n1047) );
AND2_X1 U898 ( .A1(G217), .A2(n1185), .ZN(n1087) );
OR2_X1 U899 ( .A1(n1086), .A2(G902), .ZN(n1184) );
XOR2_X1 U900 ( .A(n1186), .B(n1187), .Z(n1086) );
XOR2_X1 U901 ( .A(G110), .B(n1188), .Z(n1187) );
XNOR2_X1 U902 ( .A(n1189), .B(G137), .ZN(n1188) );
INV_X1 U903 ( .A(G146), .ZN(n1189) );
XNOR2_X1 U904 ( .A(n1190), .B(n1067), .ZN(n1186) );
XNOR2_X1 U905 ( .A(n1191), .B(n1192), .ZN(n1190) );
NAND4_X1 U906 ( .A1(KEYINPUT34), .A2(G221), .A3(G234), .A4(n1055), .ZN(n1192) );
NAND2_X1 U907 ( .A1(KEYINPUT57), .A2(n1193), .ZN(n1191) );
XOR2_X1 U908 ( .A(G128), .B(G119), .Z(n1193) );
INV_X1 U909 ( .A(n1176), .ZN(n1024) );
XOR2_X1 U910 ( .A(n1194), .B(n1041), .Z(n1176) );
XNOR2_X1 U911 ( .A(G472), .B(KEYINPUT32), .ZN(n1041) );
XOR2_X1 U912 ( .A(n1039), .B(KEYINPUT33), .Z(n1194) );
NAND2_X1 U913 ( .A1(n1195), .A2(n1137), .ZN(n1039) );
XOR2_X1 U914 ( .A(n1196), .B(n1197), .Z(n1195) );
XNOR2_X1 U915 ( .A(n1198), .B(n1112), .ZN(n1197) );
XOR2_X1 U916 ( .A(n1127), .B(n1199), .Z(n1112) );
NAND2_X1 U917 ( .A1(n1200), .A2(KEYINPUT16), .ZN(n1198) );
XNOR2_X1 U918 ( .A(n1117), .B(G101), .ZN(n1200) );
NOR3_X1 U919 ( .A1(G237), .A2(G953), .A3(n1201), .ZN(n1117) );
XNOR2_X1 U920 ( .A(KEYINPUT61), .B(G210), .ZN(n1201) );
XOR2_X1 U921 ( .A(KEYINPUT50), .B(n1202), .Z(n1196) );
NOR2_X1 U922 ( .A1(KEYINPUT47), .A2(n1111), .ZN(n1202) );
XNOR2_X1 U923 ( .A(n1203), .B(KEYINPUT46), .ZN(n1111) );
AND2_X1 U924 ( .A1(n1183), .A2(n1181), .ZN(n1020) );
NAND3_X1 U925 ( .A1(n1204), .A2(n1205), .A3(n1206), .ZN(n1181) );
INV_X1 U926 ( .A(n1043), .ZN(n1206) );
NOR2_X1 U927 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND3_X1 U928 ( .A1(KEYINPUT60), .A2(n1045), .A3(n1044), .ZN(n1205) );
NAND2_X1 U929 ( .A1(n1097), .A2(n1137), .ZN(n1045) );
XOR2_X1 U930 ( .A(n1207), .B(KEYINPUT12), .Z(n1097) );
XOR2_X1 U931 ( .A(n1208), .B(n1209), .Z(n1207) );
XOR2_X1 U932 ( .A(n1210), .B(n1211), .Z(n1209) );
XOR2_X1 U933 ( .A(G104), .B(n1212), .Z(n1211) );
NOR3_X1 U934 ( .A1(n1213), .A2(G953), .A3(G237), .ZN(n1212) );
INV_X1 U935 ( .A(G214), .ZN(n1213) );
XNOR2_X1 U936 ( .A(n1170), .B(G113), .ZN(n1210) );
XOR2_X1 U937 ( .A(n1214), .B(n1215), .Z(n1208) );
XOR2_X1 U938 ( .A(n1216), .B(n1217), .Z(n1215) );
NAND2_X1 U939 ( .A1(KEYINPUT37), .A2(n1218), .ZN(n1217) );
INV_X1 U940 ( .A(G143), .ZN(n1218) );
NAND2_X1 U941 ( .A1(KEYINPUT2), .A2(n1219), .ZN(n1216) );
XNOR2_X1 U942 ( .A(n1220), .B(n1067), .ZN(n1214) );
XNOR2_X1 U943 ( .A(G140), .B(G125), .ZN(n1067) );
NAND2_X1 U944 ( .A1(KEYINPUT43), .A2(G146), .ZN(n1220) );
OR2_X1 U945 ( .A1(n1044), .A2(KEYINPUT60), .ZN(n1204) );
INV_X1 U946 ( .A(G475), .ZN(n1044) );
INV_X1 U947 ( .A(n1046), .ZN(n1183) );
XNOR2_X1 U948 ( .A(n1221), .B(G478), .ZN(n1046) );
NAND2_X1 U949 ( .A1(n1092), .A2(n1137), .ZN(n1221) );
XNOR2_X1 U950 ( .A(n1222), .B(n1223), .ZN(n1092) );
XOR2_X1 U951 ( .A(n1224), .B(n1225), .Z(n1223) );
XNOR2_X1 U952 ( .A(G116), .B(n982), .ZN(n1225) );
AND3_X1 U953 ( .A1(n1226), .A2(G234), .A3(G217), .ZN(n1224) );
XNOR2_X1 U954 ( .A(KEYINPUT52), .B(G953), .ZN(n1226) );
XOR2_X1 U955 ( .A(n1227), .B(n1228), .Z(n1222) );
XNOR2_X1 U956 ( .A(G128), .B(n1219), .ZN(n1228) );
INV_X1 U957 ( .A(G122), .ZN(n1219) );
XNOR2_X1 U958 ( .A(G134), .B(G143), .ZN(n1227) );
INV_X1 U959 ( .A(n1100), .ZN(n1151) );
NAND3_X1 U960 ( .A1(n1030), .A2(n1148), .A3(n980), .ZN(n1100) );
INV_X1 U961 ( .A(n1175), .ZN(n980) );
NAND2_X1 U962 ( .A1(n997), .A2(n996), .ZN(n1175) );
NAND2_X1 U963 ( .A1(G214), .A2(n1229), .ZN(n996) );
XNOR2_X1 U964 ( .A(n1048), .B(n1230), .ZN(n997) );
NOR2_X1 U965 ( .A1(KEYINPUT30), .A2(n1231), .ZN(n1230) );
XOR2_X1 U966 ( .A(KEYINPUT51), .B(n1049), .Z(n1231) );
AND2_X1 U967 ( .A1(G210), .A2(n1232), .ZN(n1049) );
XNOR2_X1 U968 ( .A(KEYINPUT10), .B(n1229), .ZN(n1232) );
OR2_X1 U969 ( .A1(G902), .A2(G237), .ZN(n1229) );
NAND2_X1 U970 ( .A1(n1233), .A2(n1137), .ZN(n1048) );
XOR2_X1 U971 ( .A(n1234), .B(n1136), .Z(n1233) );
XNOR2_X1 U972 ( .A(n1076), .B(n1235), .ZN(n1136) );
XOR2_X1 U973 ( .A(n1236), .B(n1237), .Z(n1235) );
NAND2_X1 U974 ( .A1(KEYINPUT44), .A2(n1077), .ZN(n1237) );
XNOR2_X1 U975 ( .A(G110), .B(G122), .ZN(n1077) );
NAND2_X1 U976 ( .A1(G224), .A2(n1055), .ZN(n1236) );
XOR2_X1 U977 ( .A(n1238), .B(n1239), .Z(n1076) );
XOR2_X1 U978 ( .A(KEYINPUT15), .B(n1240), .Z(n1239) );
XOR2_X1 U979 ( .A(KEYINPUT55), .B(KEYINPUT49), .Z(n1240) );
XNOR2_X1 U980 ( .A(n1126), .B(n1199), .ZN(n1238) );
XOR2_X1 U981 ( .A(G113), .B(n1241), .Z(n1199) );
XOR2_X1 U982 ( .A(G119), .B(G116), .Z(n1241) );
NAND3_X1 U983 ( .A1(n1242), .A2(n1243), .A3(KEYINPUT48), .ZN(n1234) );
NAND3_X1 U984 ( .A1(G125), .A2(n1203), .A3(n1244), .ZN(n1243) );
INV_X1 U985 ( .A(KEYINPUT0), .ZN(n1244) );
NAND2_X1 U986 ( .A1(n1134), .A2(KEYINPUT0), .ZN(n1242) );
XOR2_X1 U987 ( .A(G125), .B(n1203), .Z(n1134) );
XNOR2_X1 U988 ( .A(n1245), .B(n1246), .ZN(n1203) );
NOR2_X1 U989 ( .A1(KEYINPUT35), .A2(G128), .ZN(n1246) );
XNOR2_X1 U990 ( .A(G143), .B(G146), .ZN(n1245) );
NAND2_X1 U991 ( .A1(n1031), .A2(n1247), .ZN(n1148) );
NAND4_X1 U992 ( .A1(n1075), .A2(G953), .A3(G902), .A4(n1178), .ZN(n1247) );
XNOR2_X1 U993 ( .A(G898), .B(KEYINPUT58), .ZN(n1075) );
NAND3_X1 U994 ( .A1(n1178), .A2(n1055), .A3(G952), .ZN(n1031) );
INV_X1 U995 ( .A(G953), .ZN(n1055) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1178) );
NOR2_X1 U997 ( .A1(n1009), .A2(n1007), .ZN(n1030) );
INV_X1 U998 ( .A(n1182), .ZN(n1007) );
NAND2_X1 U999 ( .A1(G221), .A2(n1185), .ZN(n1182) );
NAND2_X1 U1000 ( .A1(G234), .A2(n1137), .ZN(n1185) );
XOR2_X1 U1001 ( .A(n1248), .B(G469), .Z(n1009) );
NAND2_X1 U1002 ( .A1(n1249), .A2(n1137), .ZN(n1248) );
INV_X1 U1003 ( .A(G902), .ZN(n1137) );
XOR2_X1 U1004 ( .A(n1250), .B(n1251), .Z(n1249) );
XNOR2_X1 U1005 ( .A(n1252), .B(n1253), .ZN(n1251) );
NOR2_X1 U1006 ( .A1(KEYINPUT19), .A2(n1127), .ZN(n1253) );
XNOR2_X1 U1007 ( .A(n1254), .B(KEYINPUT31), .ZN(n1127) );
NAND2_X1 U1008 ( .A1(n1255), .A2(n1256), .ZN(n1254) );
OR2_X1 U1009 ( .A1(n1170), .A2(n1257), .ZN(n1256) );
XOR2_X1 U1010 ( .A(n1258), .B(KEYINPUT53), .Z(n1255) );
NAND2_X1 U1011 ( .A1(n1257), .A2(n1170), .ZN(n1258) );
INV_X1 U1012 ( .A(G131), .ZN(n1170) );
XOR2_X1 U1013 ( .A(n1063), .B(KEYINPUT59), .Z(n1257) );
XOR2_X1 U1014 ( .A(G134), .B(G137), .Z(n1063) );
NAND2_X1 U1015 ( .A1(KEYINPUT26), .A2(n1066), .ZN(n1252) );
XNOR2_X1 U1016 ( .A(n1259), .B(G128), .ZN(n1066) );
NAND3_X1 U1017 ( .A1(n1260), .A2(n1261), .A3(n1262), .ZN(n1259) );
OR2_X1 U1018 ( .A1(n1263), .A2(G146), .ZN(n1262) );
NAND2_X1 U1019 ( .A1(KEYINPUT54), .A2(n1264), .ZN(n1261) );
NAND2_X1 U1020 ( .A1(n1265), .A2(n1263), .ZN(n1264) );
XNOR2_X1 U1021 ( .A(KEYINPUT42), .B(G146), .ZN(n1265) );
NAND2_X1 U1022 ( .A1(n1266), .A2(n1267), .ZN(n1260) );
INV_X1 U1023 ( .A(KEYINPUT54), .ZN(n1267) );
NAND2_X1 U1024 ( .A1(n1268), .A2(n1269), .ZN(n1266) );
OR2_X1 U1025 ( .A1(G146), .A2(KEYINPUT42), .ZN(n1269) );
NAND3_X1 U1026 ( .A1(G146), .A2(n1263), .A3(KEYINPUT42), .ZN(n1268) );
XOR2_X1 U1027 ( .A(G143), .B(KEYINPUT28), .Z(n1263) );
XNOR2_X1 U1028 ( .A(n1126), .B(n1270), .ZN(n1250) );
NOR2_X1 U1029 ( .A1(KEYINPUT27), .A2(n1271), .ZN(n1270) );
XOR2_X1 U1030 ( .A(n1272), .B(n1131), .Z(n1271) );
NOR2_X1 U1031 ( .A1(n1056), .A2(G953), .ZN(n1131) );
INV_X1 U1032 ( .A(G227), .ZN(n1056) );
NAND2_X1 U1033 ( .A1(KEYINPUT11), .A2(n1124), .ZN(n1272) );
XOR2_X1 U1034 ( .A(G140), .B(G110), .Z(n1124) );
XOR2_X1 U1035 ( .A(G101), .B(n1273), .Z(n1126) );
XNOR2_X1 U1036 ( .A(n982), .B(G104), .ZN(n1273) );
INV_X1 U1037 ( .A(G107), .ZN(n982) );
endmodule


