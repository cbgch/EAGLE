//Key = 0100111001111110011001111010110011001011101001100001000000100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289;

XOR2_X1 U720 ( .A(n993), .B(n994), .Z(G9) );
NOR2_X1 U721 ( .A1(n995), .A2(n996), .ZN(G75) );
XOR2_X1 U722 ( .A(n997), .B(KEYINPUT9), .Z(n996) );
OR3_X1 U723 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n997) );
OR3_X1 U724 ( .A1(n1001), .A2(n1002), .A3(n1003), .ZN(n1000) );
NOR3_X1 U725 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1003) );
NOR2_X1 U726 ( .A1(n1007), .A2(n1008), .ZN(n1005) );
NOR4_X1 U727 ( .A1(n1009), .A2(n1010), .A3(n1011), .A4(n1012), .ZN(n1008) );
NOR3_X1 U728 ( .A1(n1013), .A2(n1014), .A3(n1015), .ZN(n1010) );
NOR2_X1 U729 ( .A1(n1016), .A2(n1017), .ZN(n1009) );
NOR3_X1 U730 ( .A1(n1018), .A2(n1013), .A3(n1019), .ZN(n1007) );
NOR2_X1 U731 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NOR2_X1 U732 ( .A1(n1022), .A2(n1011), .ZN(n1021) );
NOR2_X1 U733 ( .A1(n1023), .A2(n1024), .ZN(n1022) );
NOR2_X1 U734 ( .A1(n1025), .A2(n1026), .ZN(n1024) );
AND2_X1 U735 ( .A1(n1027), .A2(KEYINPUT22), .ZN(n1023) );
NOR2_X1 U736 ( .A1(n1028), .A2(n1012), .ZN(n1020) );
INV_X1 U737 ( .A(n1029), .ZN(n1012) );
NOR2_X1 U738 ( .A1(n1030), .A2(n1031), .ZN(n1028) );
AND2_X1 U739 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR3_X1 U740 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1002) );
XNOR2_X1 U741 ( .A(KEYINPUT39), .B(n1004), .ZN(n1036) );
XOR2_X1 U742 ( .A(KEYINPUT4), .B(n1029), .Z(n1035) );
NAND3_X1 U743 ( .A1(n1037), .A2(n1038), .A3(n1016), .ZN(n1034) );
NOR2_X1 U744 ( .A1(KEYINPUT22), .A2(n1039), .ZN(n1001) );
NOR4_X1 U745 ( .A1(n1011), .A2(n1018), .A3(n1040), .A4(n1004), .ZN(n1039) );
NOR2_X1 U746 ( .A1(G952), .A2(n999), .ZN(n995) );
NAND2_X1 U747 ( .A1(n1041), .A2(n1042), .ZN(n999) );
NAND4_X1 U748 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1042) );
NOR4_X1 U749 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1013), .ZN(n1046) );
INV_X1 U750 ( .A(n1050), .ZN(n1049) );
NOR2_X1 U751 ( .A1(n1018), .A2(n1051), .ZN(n1045) );
XOR2_X1 U752 ( .A(n1052), .B(n1053), .Z(n1051) );
INV_X1 U753 ( .A(n1016), .ZN(n1018) );
XOR2_X1 U754 ( .A(n1054), .B(n1055), .Z(n1044) );
XOR2_X1 U755 ( .A(n1056), .B(KEYINPUT24), .Z(n1055) );
XOR2_X1 U756 ( .A(n1057), .B(n1058), .Z(G72) );
XOR2_X1 U757 ( .A(n1059), .B(n1060), .Z(n1058) );
NAND2_X1 U758 ( .A1(G953), .A2(n1061), .ZN(n1060) );
NAND2_X1 U759 ( .A1(G900), .A2(G227), .ZN(n1061) );
NAND2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1059) );
NAND2_X1 U761 ( .A1(G953), .A2(n1064), .ZN(n1063) );
XOR2_X1 U762 ( .A(n1065), .B(n1066), .Z(n1062) );
XOR2_X1 U763 ( .A(n1067), .B(n1068), .Z(n1066) );
XOR2_X1 U764 ( .A(n1069), .B(n1070), .Z(n1065) );
XOR2_X1 U765 ( .A(KEYINPUT18), .B(G131), .Z(n1070) );
NAND2_X1 U766 ( .A1(KEYINPUT36), .A2(n1071), .ZN(n1069) );
NOR2_X1 U767 ( .A1(n1072), .A2(G953), .ZN(n1057) );
NAND2_X1 U768 ( .A1(n1073), .A2(n1074), .ZN(G69) );
NAND2_X1 U769 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND2_X1 U770 ( .A1(G953), .A2(n1077), .ZN(n1076) );
XOR2_X1 U771 ( .A(n1078), .B(n1079), .Z(n1075) );
NOR2_X1 U772 ( .A1(n1080), .A2(KEYINPUT30), .ZN(n1079) );
AND2_X1 U773 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
XOR2_X1 U774 ( .A(KEYINPUT42), .B(n1083), .Z(n1073) );
NOR3_X1 U775 ( .A1(n1041), .A2(n1078), .A3(n1084), .ZN(n1083) );
INV_X1 U776 ( .A(n1077), .ZN(n1084) );
NAND2_X1 U777 ( .A1(G898), .A2(G224), .ZN(n1077) );
AND2_X1 U778 ( .A1(n1085), .A2(n1086), .ZN(n1078) );
NAND2_X1 U779 ( .A1(G953), .A2(n1087), .ZN(n1086) );
XNOR2_X1 U780 ( .A(n1088), .B(n1089), .ZN(n1085) );
NOR2_X1 U781 ( .A1(KEYINPUT34), .A2(n1090), .ZN(n1088) );
NOR3_X1 U782 ( .A1(n1091), .A2(n1092), .A3(n1093), .ZN(G66) );
AND2_X1 U783 ( .A1(KEYINPUT5), .A2(n1094), .ZN(n1093) );
NOR3_X1 U784 ( .A1(KEYINPUT5), .A2(n1041), .A3(n1095), .ZN(n1092) );
INV_X1 U785 ( .A(G952), .ZN(n1095) );
XNOR2_X1 U786 ( .A(n1096), .B(n1097), .ZN(n1091) );
NAND2_X1 U787 ( .A1(KEYINPUT51), .A2(n1098), .ZN(n1096) );
OR2_X1 U788 ( .A1(n1099), .A2(n1053), .ZN(n1098) );
NOR2_X1 U789 ( .A1(n1094), .A2(n1100), .ZN(G63) );
XNOR2_X1 U790 ( .A(n1101), .B(n1102), .ZN(n1100) );
AND2_X1 U791 ( .A1(G478), .A2(n1103), .ZN(n1102) );
NOR2_X1 U792 ( .A1(n1094), .A2(n1104), .ZN(G60) );
XOR2_X1 U793 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U794 ( .A1(KEYINPUT19), .A2(n1107), .ZN(n1106) );
NAND2_X1 U795 ( .A1(n1103), .A2(G475), .ZN(n1105) );
XNOR2_X1 U796 ( .A(G104), .B(n1108), .ZN(G6) );
NOR2_X1 U797 ( .A1(n1094), .A2(n1109), .ZN(G57) );
XOR2_X1 U798 ( .A(n1110), .B(n1111), .Z(n1109) );
XOR2_X1 U799 ( .A(KEYINPUT43), .B(n1112), .Z(n1111) );
AND2_X1 U800 ( .A1(G472), .A2(n1103), .ZN(n1112) );
INV_X1 U801 ( .A(n1099), .ZN(n1103) );
XOR2_X1 U802 ( .A(n1113), .B(n1114), .Z(n1110) );
NAND2_X1 U803 ( .A1(n1115), .A2(n1116), .ZN(n1113) );
NAND2_X1 U804 ( .A1(KEYINPUT32), .A2(n1117), .ZN(n1116) );
OR3_X1 U805 ( .A1(n1118), .A2(n1119), .A3(KEYINPUT32), .ZN(n1115) );
NOR2_X1 U806 ( .A1(n1094), .A2(n1120), .ZN(G54) );
XOR2_X1 U807 ( .A(n1121), .B(n1122), .Z(n1120) );
XOR2_X1 U808 ( .A(n1123), .B(n1124), .Z(n1122) );
NOR2_X1 U809 ( .A1(KEYINPUT8), .A2(n1125), .ZN(n1123) );
XOR2_X1 U810 ( .A(n1126), .B(n1119), .Z(n1121) );
NOR2_X1 U811 ( .A1(n1127), .A2(n1099), .ZN(n1126) );
XNOR2_X1 U812 ( .A(G469), .B(KEYINPUT61), .ZN(n1127) );
NOR2_X1 U813 ( .A1(n1094), .A2(n1128), .ZN(G51) );
XOR2_X1 U814 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U815 ( .A(G125), .B(n1131), .Z(n1130) );
NOR2_X1 U816 ( .A1(n1054), .A2(n1099), .ZN(n1131) );
NAND2_X1 U817 ( .A1(G902), .A2(n998), .ZN(n1099) );
NAND3_X1 U818 ( .A1(n1072), .A2(n1082), .A3(n1132), .ZN(n998) );
XOR2_X1 U819 ( .A(n1081), .B(KEYINPUT52), .Z(n1132) );
AND4_X1 U820 ( .A1(n1108), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1082) );
AND4_X1 U821 ( .A1(n1136), .A2(n1137), .A3(n994), .A4(n1138), .ZN(n1135) );
NAND3_X1 U822 ( .A1(n1015), .A2(n1037), .A3(n1139), .ZN(n994) );
NAND3_X1 U823 ( .A1(n1140), .A2(n1014), .A3(n1141), .ZN(n1134) );
NAND3_X1 U824 ( .A1(n1139), .A2(n1037), .A3(n1014), .ZN(n1108) );
AND2_X1 U825 ( .A1(n1142), .A2(n1143), .ZN(n1072) );
NOR4_X1 U826 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1143) );
AND4_X1 U827 ( .A1(n1148), .A2(n1149), .A3(n1150), .A4(n1151), .ZN(n1142) );
NOR2_X1 U828 ( .A1(n1041), .A2(G952), .ZN(n1094) );
XOR2_X1 U829 ( .A(n1152), .B(n1151), .Z(G48) );
NAND3_X1 U830 ( .A1(n1153), .A2(n1027), .A3(n1014), .ZN(n1151) );
XNOR2_X1 U831 ( .A(G143), .B(n1150), .ZN(G45) );
NAND4_X1 U832 ( .A1(n1154), .A2(n1027), .A3(n1155), .A4(n1156), .ZN(n1150) );
XOR2_X1 U833 ( .A(G140), .B(n1145), .Z(G42) );
AND3_X1 U834 ( .A1(n1029), .A2(n1038), .A3(n1157), .ZN(n1145) );
XNOR2_X1 U835 ( .A(G137), .B(n1158), .ZN(G39) );
NOR2_X1 U836 ( .A1(n1144), .A2(KEYINPUT20), .ZN(n1158) );
AND3_X1 U837 ( .A1(n1029), .A2(n1016), .A3(n1153), .ZN(n1144) );
XOR2_X1 U838 ( .A(n1149), .B(n1159), .Z(G36) );
NOR2_X1 U839 ( .A1(G134), .A2(KEYINPUT0), .ZN(n1159) );
NAND3_X1 U840 ( .A1(n1029), .A2(n1015), .A3(n1154), .ZN(n1149) );
XOR2_X1 U841 ( .A(n1160), .B(n1148), .Z(G33) );
NAND3_X1 U842 ( .A1(n1014), .A2(n1029), .A3(n1154), .ZN(n1148) );
AND3_X1 U843 ( .A1(n1038), .A2(n1161), .A3(n1031), .ZN(n1154) );
NOR2_X1 U844 ( .A1(n1025), .A2(n1048), .ZN(n1029) );
INV_X1 U845 ( .A(n1026), .ZN(n1048) );
XOR2_X1 U846 ( .A(G128), .B(n1147), .Z(G30) );
AND3_X1 U847 ( .A1(n1015), .A2(n1027), .A3(n1153), .ZN(n1147) );
AND4_X1 U848 ( .A1(n1162), .A2(n1038), .A3(n1163), .A4(n1161), .ZN(n1153) );
XNOR2_X1 U849 ( .A(G101), .B(n1133), .ZN(G3) );
NAND3_X1 U850 ( .A1(n1016), .A2(n1139), .A3(n1031), .ZN(n1133) );
XOR2_X1 U851 ( .A(G125), .B(n1146), .Z(G27) );
AND2_X1 U852 ( .A1(n1164), .A2(n1157), .ZN(n1146) );
AND4_X1 U853 ( .A1(n1033), .A2(n1014), .A3(n1032), .A4(n1161), .ZN(n1157) );
NAND2_X1 U854 ( .A1(n1004), .A2(n1165), .ZN(n1161) );
NAND4_X1 U855 ( .A1(G953), .A2(G902), .A3(n1166), .A4(n1167), .ZN(n1165) );
XOR2_X1 U856 ( .A(KEYINPUT2), .B(n1064), .Z(n1166) );
XOR2_X1 U857 ( .A(G900), .B(KEYINPUT23), .Z(n1064) );
XOR2_X1 U858 ( .A(n1168), .B(n1081), .Z(G24) );
NAND3_X1 U859 ( .A1(n1164), .A2(n1037), .A3(n1169), .ZN(n1081) );
AND3_X1 U860 ( .A1(n1155), .A2(n1170), .A3(n1156), .ZN(n1169) );
INV_X1 U861 ( .A(n1011), .ZN(n1037) );
NAND2_X1 U862 ( .A1(n1171), .A2(n1032), .ZN(n1011) );
XNOR2_X1 U863 ( .A(G119), .B(n1137), .ZN(G21) );
NAND3_X1 U864 ( .A1(n1164), .A2(n1016), .A3(n1172), .ZN(n1137) );
AND3_X1 U865 ( .A1(n1162), .A2(n1170), .A3(n1163), .ZN(n1172) );
XNOR2_X1 U866 ( .A(n1171), .B(KEYINPUT48), .ZN(n1163) );
INV_X1 U867 ( .A(n1040), .ZN(n1164) );
NAND3_X1 U868 ( .A1(n1027), .A2(n1017), .A3(n1173), .ZN(n1040) );
XNOR2_X1 U869 ( .A(G116), .B(n1136), .ZN(G18) );
NAND3_X1 U870 ( .A1(n1015), .A2(n1027), .A3(n1141), .ZN(n1136) );
NOR2_X1 U871 ( .A1(n1156), .A2(n1174), .ZN(n1015) );
XOR2_X1 U872 ( .A(n1175), .B(n1176), .Z(G15) );
NAND3_X1 U873 ( .A1(n1177), .A2(n1141), .A3(n1178), .ZN(n1176) );
XNOR2_X1 U874 ( .A(n1014), .B(KEYINPUT21), .ZN(n1178) );
AND2_X1 U875 ( .A1(n1174), .A2(n1156), .ZN(n1014) );
AND4_X1 U876 ( .A1(n1031), .A2(n1173), .A3(n1017), .A4(n1170), .ZN(n1141) );
AND2_X1 U877 ( .A1(n1171), .A2(n1179), .ZN(n1031) );
XNOR2_X1 U878 ( .A(KEYINPUT40), .B(n1162), .ZN(n1179) );
XOR2_X1 U879 ( .A(n1140), .B(KEYINPUT31), .Z(n1177) );
XOR2_X1 U880 ( .A(n1138), .B(n1180), .Z(G12) );
NAND2_X1 U881 ( .A1(KEYINPUT26), .A2(G110), .ZN(n1180) );
NAND4_X1 U882 ( .A1(n1033), .A2(n1016), .A3(n1139), .A4(n1032), .ZN(n1138) );
XNOR2_X1 U883 ( .A(n1162), .B(KEYINPUT63), .ZN(n1032) );
XOR2_X1 U884 ( .A(n1043), .B(KEYINPUT29), .Z(n1162) );
XOR2_X1 U885 ( .A(n1181), .B(G472), .Z(n1043) );
NAND2_X1 U886 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U887 ( .A(n1114), .B(n1117), .ZN(n1182) );
XOR2_X1 U888 ( .A(n1119), .B(n1118), .Z(n1117) );
INV_X1 U889 ( .A(n1184), .ZN(n1119) );
XNOR2_X1 U890 ( .A(n1185), .B(n1186), .ZN(n1114) );
XOR2_X1 U891 ( .A(G101), .B(n1187), .Z(n1186) );
XOR2_X1 U892 ( .A(G116), .B(G113), .Z(n1187) );
XOR2_X1 U893 ( .A(n1188), .B(n1189), .Z(n1185) );
NOR2_X1 U894 ( .A1(KEYINPUT25), .A2(G119), .ZN(n1189) );
NAND2_X1 U895 ( .A1(n1190), .A2(G210), .ZN(n1188) );
AND3_X1 U896 ( .A1(n1140), .A2(n1170), .A3(n1038), .ZN(n1139) );
NOR2_X1 U897 ( .A1(n1013), .A2(n1173), .ZN(n1038) );
INV_X1 U898 ( .A(n1006), .ZN(n1173) );
NAND2_X1 U899 ( .A1(n1191), .A2(n1050), .ZN(n1006) );
NAND2_X1 U900 ( .A1(n1192), .A2(n1193), .ZN(n1050) );
OR2_X1 U901 ( .A1(n1194), .A2(G902), .ZN(n1193) );
XNOR2_X1 U902 ( .A(n1047), .B(KEYINPUT50), .ZN(n1191) );
NOR3_X1 U903 ( .A1(n1194), .A2(G902), .A3(n1192), .ZN(n1047) );
XOR2_X1 U904 ( .A(G469), .B(KEYINPUT16), .Z(n1192) );
XOR2_X1 U905 ( .A(n1195), .B(n1196), .Z(n1194) );
XNOR2_X1 U906 ( .A(n1197), .B(KEYINPUT3), .ZN(n1196) );
NAND2_X1 U907 ( .A1(KEYINPUT10), .A2(n1184), .ZN(n1197) );
NAND2_X1 U908 ( .A1(n1198), .A2(n1199), .ZN(n1184) );
NAND2_X1 U909 ( .A1(n1200), .A2(n1201), .ZN(n1199) );
NAND2_X1 U910 ( .A1(n1202), .A2(n1203), .ZN(n1201) );
NAND2_X1 U911 ( .A1(KEYINPUT45), .A2(n1160), .ZN(n1203) );
INV_X1 U912 ( .A(KEYINPUT44), .ZN(n1202) );
NAND2_X1 U913 ( .A1(G131), .A2(n1204), .ZN(n1198) );
NAND2_X1 U914 ( .A1(KEYINPUT45), .A2(n1205), .ZN(n1204) );
OR2_X1 U915 ( .A1(n1200), .A2(KEYINPUT44), .ZN(n1205) );
XNOR2_X1 U916 ( .A(n1071), .B(KEYINPUT14), .ZN(n1200) );
XOR2_X1 U917 ( .A(G134), .B(G137), .Z(n1071) );
XOR2_X1 U918 ( .A(n1124), .B(n1125), .Z(n1195) );
XNOR2_X1 U919 ( .A(G110), .B(G140), .ZN(n1125) );
XNOR2_X1 U920 ( .A(n1206), .B(n1207), .ZN(n1124) );
INV_X1 U921 ( .A(n1067), .ZN(n1207) );
XOR2_X1 U922 ( .A(n1152), .B(n1208), .Z(n1067) );
XOR2_X1 U923 ( .A(n1209), .B(n1210), .Z(n1206) );
AND2_X1 U924 ( .A1(n1041), .A2(G227), .ZN(n1210) );
NAND2_X1 U925 ( .A1(n1211), .A2(n1212), .ZN(n1209) );
NAND2_X1 U926 ( .A1(n1213), .A2(n993), .ZN(n1212) );
XOR2_X1 U927 ( .A(KEYINPUT58), .B(n1214), .Z(n1213) );
INV_X1 U928 ( .A(n1017), .ZN(n1013) );
NAND2_X1 U929 ( .A1(G221), .A2(n1215), .ZN(n1017) );
NAND2_X1 U930 ( .A1(n1004), .A2(n1216), .ZN(n1170) );
NAND4_X1 U931 ( .A1(G953), .A2(G902), .A3(n1167), .A4(n1087), .ZN(n1216) );
INV_X1 U932 ( .A(G898), .ZN(n1087) );
NAND3_X1 U933 ( .A1(n1167), .A2(n1041), .A3(n1217), .ZN(n1004) );
XOR2_X1 U934 ( .A(KEYINPUT7), .B(G952), .Z(n1217) );
NAND2_X1 U935 ( .A1(G237), .A2(G234), .ZN(n1167) );
XNOR2_X1 U936 ( .A(n1027), .B(KEYINPUT13), .ZN(n1140) );
AND2_X1 U937 ( .A1(n1025), .A2(n1026), .ZN(n1027) );
NAND2_X1 U938 ( .A1(G214), .A2(n1218), .ZN(n1026) );
XOR2_X1 U939 ( .A(n1056), .B(n1219), .Z(n1025) );
NOR2_X1 U940 ( .A1(n1220), .A2(n1221), .ZN(n1219) );
NOR2_X1 U941 ( .A1(KEYINPUT46), .A2(n1222), .ZN(n1221) );
AND2_X1 U942 ( .A1(KEYINPUT17), .A2(n1222), .ZN(n1220) );
INV_X1 U943 ( .A(n1054), .ZN(n1222) );
NAND2_X1 U944 ( .A1(G210), .A2(n1218), .ZN(n1054) );
NAND2_X1 U945 ( .A1(n1223), .A2(n1183), .ZN(n1218) );
INV_X1 U946 ( .A(G237), .ZN(n1223) );
NAND2_X1 U947 ( .A1(n1224), .A2(n1183), .ZN(n1056) );
XOR2_X1 U948 ( .A(n1225), .B(n1129), .Z(n1224) );
XNOR2_X1 U949 ( .A(n1118), .B(n1226), .ZN(n1129) );
XOR2_X1 U950 ( .A(n1227), .B(n1228), .Z(n1226) );
NAND2_X1 U951 ( .A1(G224), .A2(n1041), .ZN(n1228) );
NAND2_X1 U952 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
NAND2_X1 U953 ( .A1(n1089), .A2(n1090), .ZN(n1230) );
XOR2_X1 U954 ( .A(n1231), .B(KEYINPUT57), .Z(n1229) );
OR2_X1 U955 ( .A1(n1090), .A2(n1089), .ZN(n1231) );
XOR2_X1 U956 ( .A(n1232), .B(n1233), .Z(n1089) );
XOR2_X1 U957 ( .A(n1175), .B(n1234), .Z(n1233) );
NAND2_X1 U958 ( .A1(n1211), .A2(n1235), .ZN(n1234) );
NAND2_X1 U959 ( .A1(n1236), .A2(n993), .ZN(n1235) );
INV_X1 U960 ( .A(G107), .ZN(n993) );
XNOR2_X1 U961 ( .A(n1214), .B(KEYINPUT35), .ZN(n1236) );
NAND2_X1 U962 ( .A1(G107), .A2(n1214), .ZN(n1211) );
XOR2_X1 U963 ( .A(G101), .B(G104), .Z(n1214) );
XNOR2_X1 U964 ( .A(G116), .B(G119), .ZN(n1232) );
XOR2_X1 U965 ( .A(G110), .B(n1237), .Z(n1090) );
NOR2_X1 U966 ( .A1(KEYINPUT55), .A2(n1168), .ZN(n1237) );
XNOR2_X1 U967 ( .A(G128), .B(n1238), .ZN(n1118) );
NOR2_X1 U968 ( .A1(KEYINPUT37), .A2(n1239), .ZN(n1238) );
XOR2_X1 U969 ( .A(G143), .B(n1152), .Z(n1239) );
NOR2_X1 U970 ( .A1(G125), .A2(KEYINPUT62), .ZN(n1225) );
NOR2_X1 U971 ( .A1(n1155), .A2(n1156), .ZN(n1016) );
XNOR2_X1 U972 ( .A(n1240), .B(n1241), .ZN(n1156) );
XOR2_X1 U973 ( .A(KEYINPUT49), .B(G475), .Z(n1241) );
OR2_X1 U974 ( .A1(n1107), .A2(G902), .ZN(n1240) );
XNOR2_X1 U975 ( .A(n1242), .B(n1243), .ZN(n1107) );
XNOR2_X1 U976 ( .A(G104), .B(n1244), .ZN(n1243) );
NAND3_X1 U977 ( .A1(n1245), .A2(n1246), .A3(n1247), .ZN(n1244) );
NAND2_X1 U978 ( .A1(n1248), .A2(n1175), .ZN(n1247) );
INV_X1 U979 ( .A(G113), .ZN(n1175) );
NAND2_X1 U980 ( .A1(KEYINPUT28), .A2(n1249), .ZN(n1248) );
XOR2_X1 U981 ( .A(KEYINPUT38), .B(G122), .Z(n1249) );
NAND3_X1 U982 ( .A1(KEYINPUT28), .A2(G113), .A3(n1168), .ZN(n1246) );
OR2_X1 U983 ( .A1(n1168), .A2(KEYINPUT28), .ZN(n1245) );
INV_X1 U984 ( .A(G122), .ZN(n1168) );
XOR2_X1 U985 ( .A(n1250), .B(n1251), .Z(n1242) );
NOR2_X1 U986 ( .A1(KEYINPUT27), .A2(n1252), .ZN(n1251) );
XOR2_X1 U987 ( .A(n1253), .B(n1254), .Z(n1252) );
NOR2_X1 U988 ( .A1(KEYINPUT41), .A2(n1255), .ZN(n1254) );
XOR2_X1 U989 ( .A(KEYINPUT56), .B(G140), .Z(n1255) );
XOR2_X1 U990 ( .A(G125), .B(n1152), .Z(n1253) );
NAND3_X1 U991 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1250) );
NAND2_X1 U992 ( .A1(n1259), .A2(n1160), .ZN(n1258) );
NAND2_X1 U993 ( .A1(KEYINPUT59), .A2(n1260), .ZN(n1257) );
NAND2_X1 U994 ( .A1(n1261), .A2(n1262), .ZN(n1260) );
XOR2_X1 U995 ( .A(KEYINPUT15), .B(G131), .Z(n1262) );
NAND2_X1 U996 ( .A1(n1263), .A2(n1264), .ZN(n1256) );
INV_X1 U997 ( .A(KEYINPUT59), .ZN(n1264) );
NAND2_X1 U998 ( .A1(n1265), .A2(n1266), .ZN(n1263) );
NAND2_X1 U999 ( .A1(KEYINPUT15), .A2(n1160), .ZN(n1266) );
OR3_X1 U1000 ( .A1(n1259), .A2(KEYINPUT15), .A3(n1160), .ZN(n1265) );
INV_X1 U1001 ( .A(G131), .ZN(n1160) );
INV_X1 U1002 ( .A(n1261), .ZN(n1259) );
XOR2_X1 U1003 ( .A(n1267), .B(G143), .Z(n1261) );
NAND2_X1 U1004 ( .A1(n1190), .A2(G214), .ZN(n1267) );
NOR2_X1 U1005 ( .A1(G953), .A2(G237), .ZN(n1190) );
INV_X1 U1006 ( .A(n1174), .ZN(n1155) );
XOR2_X1 U1007 ( .A(n1268), .B(G478), .Z(n1174) );
NAND2_X1 U1008 ( .A1(n1101), .A2(n1183), .ZN(n1268) );
XNOR2_X1 U1009 ( .A(n1269), .B(n1270), .ZN(n1101) );
XOR2_X1 U1010 ( .A(G116), .B(n1271), .Z(n1270) );
XOR2_X1 U1011 ( .A(G134), .B(G122), .Z(n1271) );
XOR2_X1 U1012 ( .A(n1272), .B(n1208), .Z(n1269) );
XOR2_X1 U1013 ( .A(G128), .B(G143), .Z(n1208) );
XOR2_X1 U1014 ( .A(n1273), .B(G107), .Z(n1272) );
NAND3_X1 U1015 ( .A1(G217), .A2(n1041), .A3(n1274), .ZN(n1273) );
XNOR2_X1 U1016 ( .A(G234), .B(KEYINPUT11), .ZN(n1274) );
XOR2_X1 U1017 ( .A(n1171), .B(KEYINPUT33), .Z(n1033) );
XOR2_X1 U1018 ( .A(n1052), .B(n1275), .Z(n1171) );
NOR2_X1 U1019 ( .A1(KEYINPUT53), .A2(n1053), .ZN(n1275) );
NAND2_X1 U1020 ( .A1(G217), .A2(n1215), .ZN(n1053) );
NAND2_X1 U1021 ( .A1(n1276), .A2(n1183), .ZN(n1215) );
XNOR2_X1 U1022 ( .A(G234), .B(KEYINPUT12), .ZN(n1276) );
NAND2_X1 U1023 ( .A1(n1097), .A2(n1183), .ZN(n1052) );
INV_X1 U1024 ( .A(G902), .ZN(n1183) );
XNOR2_X1 U1025 ( .A(n1277), .B(n1278), .ZN(n1097) );
XOR2_X1 U1026 ( .A(n1279), .B(n1280), .Z(n1278) );
XOR2_X1 U1027 ( .A(n1281), .B(n1282), .Z(n1280) );
NOR2_X1 U1028 ( .A1(G110), .A2(KEYINPUT54), .ZN(n1282) );
NAND2_X1 U1029 ( .A1(n1283), .A2(n1284), .ZN(n1281) );
NAND2_X1 U1030 ( .A1(n1285), .A2(n1152), .ZN(n1284) );
XOR2_X1 U1031 ( .A(n1286), .B(KEYINPUT47), .Z(n1283) );
OR2_X1 U1032 ( .A1(n1285), .A2(n1152), .ZN(n1286) );
INV_X1 U1033 ( .A(G146), .ZN(n1152) );
XOR2_X1 U1034 ( .A(n1068), .B(KEYINPUT6), .Z(n1285) );
XOR2_X1 U1035 ( .A(G125), .B(G140), .Z(n1068) );
XOR2_X1 U1036 ( .A(n1287), .B(G119), .Z(n1279) );
NAND3_X1 U1037 ( .A1(G234), .A2(n1041), .A3(G221), .ZN(n1287) );
INV_X1 U1038 ( .A(G953), .ZN(n1041) );
XOR2_X1 U1039 ( .A(n1288), .B(n1289), .Z(n1277) );
XOR2_X1 U1040 ( .A(G137), .B(G128), .Z(n1289) );
XNOR2_X1 U1041 ( .A(KEYINPUT60), .B(KEYINPUT1), .ZN(n1288) );
endmodule


