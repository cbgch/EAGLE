//Key = 1101110110111110101010110101011110000010000010110100010011001111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;

XNOR2_X1 U716 ( .A(G107), .B(n1000), .ZN(G9) );
NOR2_X1 U717 ( .A1(n1001), .A2(n1002), .ZN(G75) );
NOR3_X1 U718 ( .A1(n1003), .A2(G953), .A3(n1004), .ZN(n1002) );
XOR2_X1 U719 ( .A(KEYINPUT5), .B(n1005), .Z(n1003) );
NOR2_X1 U720 ( .A1(n1006), .A2(n1007), .ZN(n1005) );
NOR2_X1 U721 ( .A1(n1008), .A2(n1009), .ZN(n1006) );
NOR2_X1 U722 ( .A1(n1010), .A2(n1011), .ZN(n1008) );
NOR3_X1 U723 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
NOR3_X1 U724 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1013) );
NOR3_X1 U725 ( .A1(n1018), .A2(KEYINPUT25), .A3(n1019), .ZN(n1017) );
NOR2_X1 U726 ( .A1(n1020), .A2(n1021), .ZN(n1016) );
NOR2_X1 U727 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
AND2_X1 U728 ( .A1(n1024), .A2(KEYINPUT25), .ZN(n1022) );
NOR2_X1 U729 ( .A1(n1025), .A2(n1026), .ZN(n1010) );
INV_X1 U730 ( .A(n1027), .ZN(n1026) );
NOR2_X1 U731 ( .A1(n1028), .A2(n1029), .ZN(n1025) );
NOR2_X1 U732 ( .A1(n1030), .A2(n1021), .ZN(n1029) );
NOR2_X1 U733 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U734 ( .A1(n1033), .A2(n1012), .ZN(n1032) );
NOR3_X1 U735 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1033) );
NOR3_X1 U736 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1036) );
INV_X1 U737 ( .A(KEYINPUT53), .ZN(n1037) );
NOR2_X1 U738 ( .A1(KEYINPUT53), .A2(n1014), .ZN(n1035) );
NOR2_X1 U739 ( .A1(n1040), .A2(n1014), .ZN(n1031) );
NOR2_X1 U740 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
AND2_X1 U741 ( .A1(n1043), .A2(n1044), .ZN(n1041) );
NOR3_X1 U742 ( .A1(n1012), .A2(n1045), .A3(n1046), .ZN(n1028) );
XOR2_X1 U743 ( .A(n1014), .B(KEYINPUT33), .Z(n1045) );
NOR3_X1 U744 ( .A1(n1004), .A2(G953), .A3(G952), .ZN(n1001) );
AND4_X1 U745 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1004) );
NOR4_X1 U746 ( .A1(n1014), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1050) );
XOR2_X1 U747 ( .A(n1054), .B(n1055), .Z(n1053) );
XOR2_X1 U748 ( .A(KEYINPUT54), .B(n1056), .Z(n1052) );
XOR2_X1 U749 ( .A(n1057), .B(KEYINPUT17), .Z(n1051) );
NAND2_X1 U750 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
NAND2_X1 U751 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NAND2_X1 U752 ( .A1(n1062), .A2(n1063), .ZN(n1058) );
XOR2_X1 U753 ( .A(KEYINPUT21), .B(G475), .Z(n1062) );
NOR3_X1 U754 ( .A1(n1044), .A2(n1064), .A3(n1065), .ZN(n1049) );
INV_X1 U755 ( .A(n1066), .ZN(n1065) );
NAND2_X1 U756 ( .A1(G469), .A2(n1067), .ZN(n1048) );
XOR2_X1 U757 ( .A(KEYINPUT16), .B(n1068), .Z(n1047) );
NOR2_X1 U758 ( .A1(G469), .A2(n1067), .ZN(n1068) );
XNOR2_X1 U759 ( .A(KEYINPUT27), .B(n1069), .ZN(n1067) );
XOR2_X1 U760 ( .A(n1070), .B(n1071), .Z(G72) );
NOR2_X1 U761 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NOR2_X1 U762 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
NAND2_X1 U763 ( .A1(n1076), .A2(n1077), .ZN(n1070) );
NAND2_X1 U764 ( .A1(n1078), .A2(n1079), .ZN(n1077) );
NAND2_X1 U765 ( .A1(n1080), .A2(n1081), .ZN(n1076) );
INV_X1 U766 ( .A(n1079), .ZN(n1081) );
NAND2_X1 U767 ( .A1(n1082), .A2(n1083), .ZN(n1079) );
NAND2_X1 U768 ( .A1(n1084), .A2(n1075), .ZN(n1083) );
XOR2_X1 U769 ( .A(KEYINPUT24), .B(G953), .Z(n1084) );
XOR2_X1 U770 ( .A(n1085), .B(n1086), .Z(n1082) );
XOR2_X1 U771 ( .A(n1087), .B(n1088), .Z(n1085) );
NAND2_X1 U772 ( .A1(KEYINPUT14), .A2(n1089), .ZN(n1087) );
XOR2_X1 U773 ( .A(KEYINPUT31), .B(n1078), .Z(n1080) );
AND2_X1 U774 ( .A1(n1073), .A2(n1090), .ZN(n1078) );
NAND2_X1 U775 ( .A1(n1091), .A2(n1092), .ZN(G69) );
NAND2_X1 U776 ( .A1(n1093), .A2(n1094), .ZN(n1092) );
NAND2_X1 U777 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
NAND2_X1 U778 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
XOR2_X1 U779 ( .A(n1099), .B(KEYINPUT45), .Z(n1091) );
NAND2_X1 U780 ( .A1(n1100), .A2(n1095), .ZN(n1099) );
NAND3_X1 U781 ( .A1(n1101), .A2(n1102), .A3(n1103), .ZN(n1095) );
NAND2_X1 U782 ( .A1(G953), .A2(n1104), .ZN(n1102) );
XNOR2_X1 U783 ( .A(n1098), .B(n1105), .ZN(n1101) );
XOR2_X1 U784 ( .A(KEYINPUT35), .B(KEYINPUT28), .Z(n1105) );
INV_X1 U785 ( .A(n1094), .ZN(n1100) );
NAND2_X1 U786 ( .A1(G953), .A2(n1106), .ZN(n1094) );
NAND2_X1 U787 ( .A1(G898), .A2(G224), .ZN(n1106) );
NOR2_X1 U788 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XNOR2_X1 U789 ( .A(n1109), .B(n1110), .ZN(n1108) );
NOR2_X1 U790 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NOR2_X1 U791 ( .A1(n1107), .A2(n1113), .ZN(G63) );
XOR2_X1 U792 ( .A(n1114), .B(n1115), .Z(n1113) );
NAND3_X1 U793 ( .A1(G478), .A2(n1007), .A3(n1116), .ZN(n1114) );
XOR2_X1 U794 ( .A(n1117), .B(KEYINPUT22), .Z(n1116) );
NOR2_X1 U795 ( .A1(n1107), .A2(n1118), .ZN(G60) );
NOR3_X1 U796 ( .A1(n1119), .A2(n1060), .A3(n1120), .ZN(n1118) );
NOR2_X1 U797 ( .A1(n1121), .A2(n1122), .ZN(n1120) );
NOR2_X1 U798 ( .A1(n1123), .A2(n1061), .ZN(n1121) );
XOR2_X1 U799 ( .A(n1124), .B(KEYINPUT30), .Z(n1119) );
NAND3_X1 U800 ( .A1(n1125), .A2(G475), .A3(n1122), .ZN(n1124) );
XNOR2_X1 U801 ( .A(G104), .B(n1126), .ZN(G6) );
NOR2_X1 U802 ( .A1(n1107), .A2(n1127), .ZN(G57) );
XOR2_X1 U803 ( .A(n1128), .B(n1129), .Z(n1127) );
NOR2_X1 U804 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
XOR2_X1 U805 ( .A(n1132), .B(n1133), .Z(n1131) );
NOR2_X1 U806 ( .A1(KEYINPUT2), .A2(n1134), .ZN(n1133) );
NOR2_X1 U807 ( .A1(n1054), .A2(n1112), .ZN(n1132) );
AND2_X1 U808 ( .A1(n1134), .A2(KEYINPUT2), .ZN(n1130) );
XNOR2_X1 U809 ( .A(n1135), .B(n1136), .ZN(n1134) );
XOR2_X1 U810 ( .A(n1137), .B(KEYINPUT50), .Z(n1135) );
NOR2_X1 U811 ( .A1(KEYINPUT42), .A2(n1138), .ZN(n1128) );
NOR2_X1 U812 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
XNOR2_X1 U813 ( .A(KEYINPUT37), .B(n1141), .ZN(n1140) );
INV_X1 U814 ( .A(n1142), .ZN(n1139) );
NOR2_X1 U815 ( .A1(n1107), .A2(n1143), .ZN(G54) );
XOR2_X1 U816 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U817 ( .A1(KEYINPUT41), .A2(n1146), .ZN(n1145) );
XNOR2_X1 U818 ( .A(n1147), .B(n1148), .ZN(n1146) );
XOR2_X1 U819 ( .A(n1149), .B(n1150), .Z(n1148) );
NOR3_X1 U820 ( .A1(KEYINPUT58), .A2(n1151), .A3(n1152), .ZN(n1150) );
NOR3_X1 U821 ( .A1(n1153), .A2(n1154), .A3(n1155), .ZN(n1152) );
INV_X1 U822 ( .A(KEYINPUT8), .ZN(n1153) );
NOR2_X1 U823 ( .A1(KEYINPUT8), .A2(n1156), .ZN(n1151) );
XOR2_X1 U824 ( .A(G140), .B(n1157), .Z(n1156) );
NAND2_X1 U825 ( .A1(n1125), .A2(G469), .ZN(n1144) );
INV_X1 U826 ( .A(n1112), .ZN(n1125) );
NOR2_X1 U827 ( .A1(n1107), .A2(n1158), .ZN(G51) );
XOR2_X1 U828 ( .A(n1159), .B(n1160), .Z(n1158) );
NOR2_X1 U829 ( .A1(n1161), .A2(n1112), .ZN(n1160) );
NAND2_X1 U830 ( .A1(G902), .A2(n1007), .ZN(n1112) );
INV_X1 U831 ( .A(n1123), .ZN(n1007) );
NOR2_X1 U832 ( .A1(n1098), .A2(n1090), .ZN(n1123) );
NAND4_X1 U833 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1090) );
AND4_X1 U834 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1165) );
NAND2_X1 U835 ( .A1(n1170), .A2(n1171), .ZN(n1164) );
NAND2_X1 U836 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
NAND4_X1 U837 ( .A1(n1174), .A2(n1175), .A3(n1042), .A4(n1176), .ZN(n1173) );
XOR2_X1 U838 ( .A(n1177), .B(KEYINPUT38), .Z(n1174) );
NAND2_X1 U839 ( .A1(n1178), .A2(n1023), .ZN(n1172) );
NAND4_X1 U840 ( .A1(n1179), .A2(n1126), .A3(n1180), .A4(n1181), .ZN(n1098) );
AND4_X1 U841 ( .A1(n1182), .A2(n1000), .A3(n1183), .A4(n1184), .ZN(n1181) );
NAND3_X1 U842 ( .A1(n1185), .A2(n1027), .A3(n1186), .ZN(n1000) );
AND2_X1 U843 ( .A1(n1187), .A2(n1188), .ZN(n1180) );
NAND2_X1 U844 ( .A1(n1015), .A2(n1186), .ZN(n1126) );
AND2_X1 U845 ( .A1(n1170), .A2(n1027), .ZN(n1015) );
NAND3_X1 U846 ( .A1(n1189), .A2(n1190), .A3(n1191), .ZN(n1179) );
NAND2_X1 U847 ( .A1(KEYINPUT11), .A2(n1192), .ZN(n1190) );
NAND2_X1 U848 ( .A1(n1193), .A2(n1194), .ZN(n1189) );
INV_X1 U849 ( .A(KEYINPUT11), .ZN(n1194) );
NAND3_X1 U850 ( .A1(n1177), .A2(n1195), .A3(n1196), .ZN(n1193) );
NAND4_X1 U851 ( .A1(KEYINPUT57), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1159) );
NAND3_X1 U852 ( .A1(n1200), .A2(n1103), .A3(n1201), .ZN(n1199) );
INV_X1 U853 ( .A(n1202), .ZN(n1201) );
NAND2_X1 U854 ( .A1(n1203), .A2(n1202), .ZN(n1198) );
XOR2_X1 U855 ( .A(n1103), .B(n1200), .Z(n1203) );
NAND2_X1 U856 ( .A1(n1204), .A2(n1097), .ZN(n1197) );
NOR2_X1 U857 ( .A1(n1073), .A2(G952), .ZN(n1107) );
XOR2_X1 U858 ( .A(n1205), .B(n1206), .Z(G48) );
NAND4_X1 U859 ( .A1(n1207), .A2(n1175), .A3(n1170), .A4(n1208), .ZN(n1206) );
XOR2_X1 U860 ( .A(n1176), .B(KEYINPUT9), .Z(n1207) );
XOR2_X1 U861 ( .A(n1209), .B(n1162), .Z(G45) );
NAND3_X1 U862 ( .A1(n1210), .A2(n1023), .A3(n1211), .ZN(n1162) );
NOR3_X1 U863 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1211) );
XOR2_X1 U864 ( .A(n1163), .B(n1215), .Z(G42) );
NAND2_X1 U865 ( .A1(KEYINPUT62), .A2(G140), .ZN(n1215) );
NAND3_X1 U866 ( .A1(n1170), .A2(n1024), .A3(n1178), .ZN(n1163) );
XOR2_X1 U867 ( .A(n1216), .B(n1169), .Z(G39) );
NAND2_X1 U868 ( .A1(n1178), .A2(n1191), .ZN(n1169) );
XNOR2_X1 U869 ( .A(G134), .B(n1168), .ZN(G36) );
NAND3_X1 U870 ( .A1(n1023), .A2(n1185), .A3(n1178), .ZN(n1168) );
AND3_X1 U871 ( .A1(n1042), .A2(n1176), .A3(n1217), .ZN(n1178) );
XOR2_X1 U872 ( .A(n1218), .B(n1219), .Z(G33) );
XNOR2_X1 U873 ( .A(G131), .B(KEYINPUT26), .ZN(n1219) );
NAND2_X1 U874 ( .A1(n1220), .A2(n1217), .ZN(n1218) );
INV_X1 U875 ( .A(n1014), .ZN(n1217) );
NAND2_X1 U876 ( .A1(n1221), .A2(n1039), .ZN(n1014) );
XOR2_X1 U877 ( .A(n1222), .B(KEYINPUT47), .Z(n1220) );
NAND4_X1 U878 ( .A1(n1170), .A2(n1023), .A3(n1223), .A4(n1176), .ZN(n1222) );
XOR2_X1 U879 ( .A(KEYINPUT19), .B(n1042), .Z(n1223) );
XNOR2_X1 U880 ( .A(G128), .B(n1167), .ZN(G30) );
NAND4_X1 U881 ( .A1(n1175), .A2(n1185), .A3(n1208), .A4(n1176), .ZN(n1167) );
XOR2_X1 U882 ( .A(n1182), .B(n1224), .Z(G3) );
NOR2_X1 U883 ( .A1(G101), .A2(KEYINPUT34), .ZN(n1224) );
NAND3_X1 U884 ( .A1(n1018), .A2(n1186), .A3(n1023), .ZN(n1182) );
XNOR2_X1 U885 ( .A(G125), .B(n1166), .ZN(G27) );
NAND4_X1 U886 ( .A1(n1170), .A2(n1196), .A3(n1225), .A4(n1024), .ZN(n1166) );
NOR2_X1 U887 ( .A1(n1213), .A2(n1177), .ZN(n1225) );
INV_X1 U888 ( .A(n1176), .ZN(n1213) );
NAND2_X1 U889 ( .A1(n1009), .A2(n1226), .ZN(n1176) );
NAND4_X1 U890 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1075), .ZN(n1226) );
INV_X1 U891 ( .A(G900), .ZN(n1075) );
XNOR2_X1 U892 ( .A(G122), .B(n1188), .ZN(G24) );
NAND4_X1 U893 ( .A1(n1228), .A2(n1210), .A3(n1027), .A4(n1056), .ZN(n1188) );
NOR2_X1 U894 ( .A1(n1229), .A2(n1230), .ZN(n1027) );
INV_X1 U895 ( .A(n1231), .ZN(n1210) );
XOR2_X1 U896 ( .A(n1232), .B(n1233), .Z(G21) );
XOR2_X1 U897 ( .A(KEYINPUT12), .B(G119), .Z(n1233) );
NAND2_X1 U898 ( .A1(n1191), .A2(n1228), .ZN(n1232) );
AND2_X1 U899 ( .A1(n1175), .A2(n1018), .ZN(n1191) );
AND2_X1 U900 ( .A1(n1234), .A2(n1229), .ZN(n1175) );
XNOR2_X1 U901 ( .A(KEYINPUT60), .B(n1230), .ZN(n1234) );
INV_X1 U902 ( .A(n1235), .ZN(n1230) );
XNOR2_X1 U903 ( .A(G116), .B(n1187), .ZN(G18) );
NAND3_X1 U904 ( .A1(n1023), .A2(n1185), .A3(n1228), .ZN(n1187) );
INV_X1 U905 ( .A(n1046), .ZN(n1185) );
NAND2_X1 U906 ( .A1(n1056), .A2(n1231), .ZN(n1046) );
XNOR2_X1 U907 ( .A(G113), .B(n1184), .ZN(G15) );
NAND3_X1 U908 ( .A1(n1170), .A2(n1023), .A3(n1228), .ZN(n1184) );
INV_X1 U909 ( .A(n1192), .ZN(n1228) );
NAND3_X1 U910 ( .A1(n1034), .A2(n1195), .A3(n1196), .ZN(n1192) );
INV_X1 U911 ( .A(n1012), .ZN(n1196) );
NAND2_X1 U912 ( .A1(n1043), .A2(n1236), .ZN(n1012) );
NOR2_X1 U913 ( .A1(n1235), .A2(n1229), .ZN(n1023) );
NOR2_X1 U914 ( .A1(n1231), .A2(n1056), .ZN(n1170) );
INV_X1 U915 ( .A(n1214), .ZN(n1056) );
XOR2_X1 U916 ( .A(n1157), .B(n1183), .Z(G12) );
NAND3_X1 U917 ( .A1(n1018), .A2(n1186), .A3(n1024), .ZN(n1183) );
INV_X1 U918 ( .A(n1019), .ZN(n1024) );
NAND2_X1 U919 ( .A1(n1235), .A2(n1229), .ZN(n1019) );
NAND2_X1 U920 ( .A1(n1237), .A2(n1066), .ZN(n1229) );
NAND3_X1 U921 ( .A1(n1111), .A2(n1117), .A3(n1109), .ZN(n1066) );
XOR2_X1 U922 ( .A(KEYINPUT13), .B(n1064), .Z(n1237) );
NOR2_X1 U923 ( .A1(n1111), .A2(n1238), .ZN(n1064) );
AND2_X1 U924 ( .A1(n1109), .A2(n1117), .ZN(n1238) );
XNOR2_X1 U925 ( .A(n1239), .B(n1240), .ZN(n1109) );
XOR2_X1 U926 ( .A(n1241), .B(n1242), .Z(n1240) );
NAND2_X1 U927 ( .A1(n1243), .A2(G221), .ZN(n1241) );
XOR2_X1 U928 ( .A(n1244), .B(n1245), .Z(n1239) );
NOR2_X1 U929 ( .A1(KEYINPUT40), .A2(n1246), .ZN(n1245) );
XOR2_X1 U930 ( .A(n1247), .B(n1248), .Z(n1246) );
XOR2_X1 U931 ( .A(KEYINPUT55), .B(G119), .Z(n1248) );
XOR2_X1 U932 ( .A(n1249), .B(G110), .Z(n1247) );
NAND2_X1 U933 ( .A1(KEYINPUT29), .A2(G128), .ZN(n1249) );
XOR2_X1 U934 ( .A(n1216), .B(G146), .Z(n1244) );
INV_X1 U935 ( .A(G137), .ZN(n1216) );
NAND2_X1 U936 ( .A1(G217), .A2(n1250), .ZN(n1111) );
XNOR2_X1 U937 ( .A(n1251), .B(n1252), .ZN(n1235) );
XNOR2_X1 U938 ( .A(KEYINPUT43), .B(n1055), .ZN(n1252) );
NAND2_X1 U939 ( .A1(n1253), .A2(n1117), .ZN(n1055) );
XOR2_X1 U940 ( .A(n1254), .B(n1255), .Z(n1253) );
NAND2_X1 U941 ( .A1(KEYINPUT20), .A2(n1256), .ZN(n1255) );
XOR2_X1 U942 ( .A(n1257), .B(n1258), .Z(n1256) );
XNOR2_X1 U943 ( .A(n1259), .B(KEYINPUT36), .ZN(n1258) );
NAND2_X1 U944 ( .A1(KEYINPUT46), .A2(n1136), .ZN(n1259) );
INV_X1 U945 ( .A(n1137), .ZN(n1257) );
XOR2_X1 U946 ( .A(n1260), .B(n1261), .Z(n1137) );
NAND2_X1 U947 ( .A1(n1141), .A2(n1142), .ZN(n1254) );
NAND4_X1 U948 ( .A1(G210), .A2(G101), .A3(n1262), .A4(n1073), .ZN(n1142) );
NAND2_X1 U949 ( .A1(n1263), .A2(n1264), .ZN(n1141) );
NAND3_X1 U950 ( .A1(n1262), .A2(n1073), .A3(G210), .ZN(n1264) );
INV_X1 U951 ( .A(G101), .ZN(n1263) );
NAND2_X1 U952 ( .A1(KEYINPUT49), .A2(n1054), .ZN(n1251) );
INV_X1 U953 ( .A(G472), .ZN(n1054) );
AND2_X1 U954 ( .A1(n1208), .A2(n1195), .ZN(n1186) );
NAND2_X1 U955 ( .A1(n1009), .A2(n1265), .ZN(n1195) );
NAND4_X1 U956 ( .A1(G953), .A2(G902), .A3(n1227), .A4(n1104), .ZN(n1265) );
INV_X1 U957 ( .A(G898), .ZN(n1104) );
NAND3_X1 U958 ( .A1(n1227), .A2(n1073), .A3(G952), .ZN(n1009) );
NAND2_X1 U959 ( .A1(G237), .A2(G234), .ZN(n1227) );
INV_X1 U960 ( .A(n1212), .ZN(n1208) );
NAND2_X1 U961 ( .A1(n1042), .A2(n1034), .ZN(n1212) );
INV_X1 U962 ( .A(n1177), .ZN(n1034) );
NAND2_X1 U963 ( .A1(n1038), .A2(n1039), .ZN(n1177) );
NAND2_X1 U964 ( .A1(G214), .A2(n1266), .ZN(n1039) );
INV_X1 U965 ( .A(n1221), .ZN(n1038) );
XNOR2_X1 U966 ( .A(n1267), .B(n1161), .ZN(n1221) );
NAND2_X1 U967 ( .A1(G210), .A2(n1266), .ZN(n1161) );
NAND2_X1 U968 ( .A1(n1262), .A2(n1117), .ZN(n1266) );
NAND4_X1 U969 ( .A1(n1268), .A2(n1117), .A3(n1269), .A4(n1270), .ZN(n1267) );
NAND3_X1 U970 ( .A1(KEYINPUT56), .A2(n1271), .A3(n1103), .ZN(n1270) );
NAND2_X1 U971 ( .A1(n1097), .A2(n1272), .ZN(n1269) );
NAND2_X1 U972 ( .A1(n1273), .A2(KEYINPUT56), .ZN(n1272) );
XNOR2_X1 U973 ( .A(n1271), .B(KEYINPUT32), .ZN(n1273) );
INV_X1 U974 ( .A(n1103), .ZN(n1097) );
XOR2_X1 U975 ( .A(n1274), .B(n1275), .Z(n1103) );
XOR2_X1 U976 ( .A(n1276), .B(n1277), .Z(n1275) );
XNOR2_X1 U977 ( .A(n1136), .B(n1278), .ZN(n1274) );
XOR2_X1 U978 ( .A(G110), .B(G101), .Z(n1278) );
XOR2_X1 U979 ( .A(G113), .B(n1279), .Z(n1136) );
XOR2_X1 U980 ( .A(G119), .B(G116), .Z(n1279) );
OR2_X1 U981 ( .A1(n1271), .A2(KEYINPUT56), .ZN(n1268) );
AND3_X1 U982 ( .A1(n1280), .A2(n1281), .A3(n1282), .ZN(n1271) );
INV_X1 U983 ( .A(n1204), .ZN(n1282) );
NOR2_X1 U984 ( .A1(n1202), .A2(n1200), .ZN(n1204) );
NAND3_X1 U985 ( .A1(KEYINPUT63), .A2(n1200), .A3(n1202), .ZN(n1281) );
XOR2_X1 U986 ( .A(G125), .B(n1261), .Z(n1200) );
XNOR2_X1 U987 ( .A(G128), .B(n1283), .ZN(n1261) );
OR2_X1 U988 ( .A1(n1202), .A2(KEYINPUT63), .ZN(n1280) );
NAND2_X1 U989 ( .A1(G224), .A2(n1073), .ZN(n1202) );
NOR2_X1 U990 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
INV_X1 U991 ( .A(n1236), .ZN(n1044) );
NAND2_X1 U992 ( .A1(G221), .A2(n1250), .ZN(n1236) );
NAND2_X1 U993 ( .A1(G234), .A2(n1117), .ZN(n1250) );
XOR2_X1 U994 ( .A(n1069), .B(G469), .Z(n1043) );
NAND2_X1 U995 ( .A1(n1284), .A2(n1117), .ZN(n1069) );
XOR2_X1 U996 ( .A(n1285), .B(n1286), .Z(n1284) );
XOR2_X1 U997 ( .A(n1149), .B(n1287), .Z(n1286) );
NOR2_X1 U998 ( .A1(KEYINPUT52), .A2(n1147), .ZN(n1287) );
XNOR2_X1 U999 ( .A(n1288), .B(n1089), .ZN(n1147) );
XOR2_X1 U1000 ( .A(G128), .B(n1289), .Z(n1089) );
NOR2_X1 U1001 ( .A1(KEYINPUT15), .A2(n1283), .ZN(n1289) );
XOR2_X1 U1002 ( .A(G143), .B(n1205), .Z(n1283) );
NAND3_X1 U1003 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1288) );
NAND2_X1 U1004 ( .A1(KEYINPUT51), .A2(n1277), .ZN(n1292) );
INV_X1 U1005 ( .A(n1293), .ZN(n1277) );
OR3_X1 U1006 ( .A1(n1294), .A2(KEYINPUT51), .A3(G101), .ZN(n1291) );
NAND2_X1 U1007 ( .A1(G101), .A2(n1294), .ZN(n1290) );
NAND2_X1 U1008 ( .A1(KEYINPUT10), .A2(n1293), .ZN(n1294) );
XOR2_X1 U1009 ( .A(G104), .B(G107), .Z(n1293) );
XOR2_X1 U1010 ( .A(n1260), .B(n1295), .Z(n1149) );
NOR2_X1 U1011 ( .A1(G953), .A2(n1074), .ZN(n1295) );
INV_X1 U1012 ( .A(G227), .ZN(n1074) );
XNOR2_X1 U1013 ( .A(n1088), .B(KEYINPUT39), .ZN(n1260) );
XOR2_X1 U1014 ( .A(G131), .B(n1296), .Z(n1088) );
XOR2_X1 U1015 ( .A(G137), .B(G134), .Z(n1296) );
XOR2_X1 U1016 ( .A(n1297), .B(KEYINPUT0), .Z(n1285) );
NAND2_X1 U1017 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
INV_X1 U1018 ( .A(n1155), .ZN(n1299) );
NOR2_X1 U1019 ( .A1(n1157), .A2(G140), .ZN(n1155) );
XNOR2_X1 U1020 ( .A(n1154), .B(KEYINPUT6), .ZN(n1298) );
AND2_X1 U1021 ( .A1(G140), .A2(n1157), .ZN(n1154) );
INV_X1 U1022 ( .A(n1021), .ZN(n1018) );
NAND2_X1 U1023 ( .A1(n1214), .A2(n1231), .ZN(n1021) );
NAND2_X1 U1024 ( .A1(n1300), .A2(n1301), .ZN(n1231) );
NAND2_X1 U1025 ( .A1(n1060), .A2(n1302), .ZN(n1301) );
NAND2_X1 U1026 ( .A1(KEYINPUT3), .A2(n1303), .ZN(n1302) );
NAND2_X1 U1027 ( .A1(KEYINPUT4), .A2(G475), .ZN(n1303) );
NAND2_X1 U1028 ( .A1(n1304), .A2(n1061), .ZN(n1300) );
INV_X1 U1029 ( .A(G475), .ZN(n1061) );
NAND2_X1 U1030 ( .A1(KEYINPUT4), .A2(n1305), .ZN(n1304) );
NAND2_X1 U1031 ( .A1(KEYINPUT3), .A2(n1063), .ZN(n1305) );
INV_X1 U1032 ( .A(n1060), .ZN(n1063) );
NOR2_X1 U1033 ( .A1(n1122), .A2(G902), .ZN(n1060) );
XNOR2_X1 U1034 ( .A(n1306), .B(n1307), .ZN(n1122) );
XOR2_X1 U1035 ( .A(n1308), .B(n1309), .Z(n1307) );
XOR2_X1 U1036 ( .A(n1242), .B(n1276), .Z(n1309) );
INV_X1 U1037 ( .A(n1086), .ZN(n1242) );
XOR2_X1 U1038 ( .A(G125), .B(G140), .Z(n1086) );
NOR2_X1 U1039 ( .A1(n1310), .A2(n1311), .ZN(n1308) );
NOR2_X1 U1040 ( .A1(KEYINPUT7), .A2(n1312), .ZN(n1311) );
INV_X1 U1041 ( .A(n1313), .ZN(n1312) );
NOR2_X1 U1042 ( .A1(KEYINPUT48), .A2(n1313), .ZN(n1310) );
XOR2_X1 U1043 ( .A(n1314), .B(n1315), .Z(n1313) );
AND3_X1 U1044 ( .A1(G214), .A2(n1073), .A3(n1262), .ZN(n1315) );
INV_X1 U1045 ( .A(G237), .ZN(n1262) );
XOR2_X1 U1046 ( .A(n1316), .B(G143), .Z(n1314) );
NAND2_X1 U1047 ( .A1(KEYINPUT44), .A2(G131), .ZN(n1316) );
XOR2_X1 U1048 ( .A(n1317), .B(n1318), .Z(n1306) );
XOR2_X1 U1049 ( .A(KEYINPUT61), .B(G113), .Z(n1318) );
XOR2_X1 U1050 ( .A(n1319), .B(G104), .Z(n1317) );
NAND2_X1 U1051 ( .A1(KEYINPUT1), .A2(n1205), .ZN(n1319) );
INV_X1 U1052 ( .A(G146), .ZN(n1205) );
XOR2_X1 U1053 ( .A(n1320), .B(G478), .Z(n1214) );
NAND2_X1 U1054 ( .A1(n1115), .A2(n1117), .ZN(n1320) );
INV_X1 U1055 ( .A(G902), .ZN(n1117) );
XNOR2_X1 U1056 ( .A(n1321), .B(n1322), .ZN(n1115) );
XOR2_X1 U1057 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1058 ( .A(G116), .B(G107), .Z(n1324) );
XOR2_X1 U1059 ( .A(G134), .B(G128), .Z(n1323) );
XOR2_X1 U1060 ( .A(n1325), .B(n1326), .Z(n1321) );
AND2_X1 U1061 ( .A1(n1243), .A2(G217), .ZN(n1326) );
AND2_X1 U1062 ( .A1(G234), .A2(n1073), .ZN(n1243) );
INV_X1 U1063 ( .A(G953), .ZN(n1073) );
XNOR2_X1 U1064 ( .A(n1327), .B(n1328), .ZN(n1325) );
NAND2_X1 U1065 ( .A1(KEYINPUT23), .A2(n1276), .ZN(n1328) );
XNOR2_X1 U1066 ( .A(G122), .B(KEYINPUT59), .ZN(n1276) );
NAND2_X1 U1067 ( .A1(KEYINPUT18), .A2(n1209), .ZN(n1327) );
INV_X1 U1068 ( .A(G143), .ZN(n1209) );
INV_X1 U1069 ( .A(G110), .ZN(n1157) );
endmodule


