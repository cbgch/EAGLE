//Key = 0010101010001110111001010100101011001110011110100110001010011010


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;

XNOR2_X1 U722 ( .A(n992), .B(n993), .ZN(G9) );
NOR2_X1 U723 ( .A1(KEYINPUT39), .A2(n994), .ZN(n993) );
NOR2_X1 U724 ( .A1(n995), .A2(n996), .ZN(G75) );
NOR4_X1 U725 ( .A1(n997), .A2(n998), .A3(n999), .A4(n1000), .ZN(n996) );
NOR2_X1 U726 ( .A1(n1001), .A2(n1002), .ZN(n998) );
NOR2_X1 U727 ( .A1(n1003), .A2(n1004), .ZN(n1001) );
NOR3_X1 U728 ( .A1(n1005), .A2(n1006), .A3(n1007), .ZN(n1004) );
NOR3_X1 U729 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
NOR2_X1 U730 ( .A1(n1011), .A2(n1012), .ZN(n1010) );
NOR2_X1 U731 ( .A1(n1013), .A2(n1014), .ZN(n1009) );
NOR2_X1 U732 ( .A1(n1015), .A2(n1016), .ZN(n1013) );
NOR2_X1 U733 ( .A1(n1017), .A2(n1018), .ZN(n1016) );
NOR3_X1 U734 ( .A1(n1019), .A2(n1020), .A3(n1021), .ZN(n1017) );
NOR2_X1 U735 ( .A1(n1012), .A2(n1022), .ZN(n1021) );
NOR2_X1 U736 ( .A1(n1023), .A2(n1024), .ZN(n1019) );
NOR3_X1 U737 ( .A1(n1025), .A2(KEYINPUT16), .A3(n1011), .ZN(n1015) );
AND3_X1 U738 ( .A1(n1026), .A2(n1027), .A3(n1028), .ZN(n1011) );
NAND2_X1 U739 ( .A1(n1029), .A2(n1030), .ZN(n1027) );
OR2_X1 U740 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NAND2_X1 U741 ( .A1(n1033), .A2(n1034), .ZN(n1026) );
NAND2_X1 U742 ( .A1(n1035), .A2(n1036), .ZN(n1034) );
NAND3_X1 U743 ( .A1(n1037), .A2(n1022), .A3(n1038), .ZN(n1036) );
INV_X1 U744 ( .A(KEYINPUT52), .ZN(n1022) );
NAND2_X1 U745 ( .A1(KEYINPUT16), .A2(n1039), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1040), .A2(n1041), .ZN(n1006) );
AND2_X1 U747 ( .A1(n1042), .A2(n1040), .ZN(n1003) );
NOR3_X1 U748 ( .A1(n1012), .A2(n1018), .A3(n1014), .ZN(n1040) );
INV_X1 U749 ( .A(n1028), .ZN(n1012) );
NOR3_X1 U750 ( .A1(n1000), .A2(G952), .A3(n997), .ZN(n995) );
AND4_X1 U751 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n997) );
NOR4_X1 U752 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
XOR2_X1 U753 ( .A(n1051), .B(n1052), .Z(n1050) );
XOR2_X1 U754 ( .A(KEYINPUT63), .B(G475), .Z(n1052) );
NOR2_X1 U755 ( .A1(KEYINPUT3), .A2(n1053), .ZN(n1051) );
XOR2_X1 U756 ( .A(n1054), .B(KEYINPUT21), .Z(n1048) );
XOR2_X1 U757 ( .A(n1055), .B(KEYINPUT32), .Z(n1047) );
NAND2_X1 U758 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
NOR3_X1 U759 ( .A1(n1058), .A2(n1038), .A3(n1059), .ZN(n1045) );
NOR2_X1 U760 ( .A1(n1056), .A2(n1057), .ZN(n1058) );
XOR2_X1 U761 ( .A(G472), .B(KEYINPUT4), .Z(n1057) );
XOR2_X1 U762 ( .A(n1060), .B(n1061), .Z(n1044) );
XOR2_X1 U763 ( .A(KEYINPUT19), .B(G478), .Z(n1061) );
NOR2_X1 U764 ( .A1(n1062), .A2(KEYINPUT35), .ZN(n1060) );
XOR2_X1 U765 ( .A(n1063), .B(n1064), .Z(n1043) );
NOR2_X1 U766 ( .A1(n1065), .A2(KEYINPUT27), .ZN(n1064) );
INV_X1 U767 ( .A(n1066), .ZN(n1000) );
NAND2_X1 U768 ( .A1(n1067), .A2(n1068), .ZN(G72) );
NAND4_X1 U769 ( .A1(G953), .A2(n1069), .A3(n1070), .A4(n1071), .ZN(n1068) );
NAND2_X1 U770 ( .A1(KEYINPUT26), .A2(n1072), .ZN(n1071) );
NAND2_X1 U771 ( .A1(KEYINPUT18), .A2(n1073), .ZN(n1070) );
NAND2_X1 U772 ( .A1(KEYINPUT18), .A2(n1074), .ZN(n1067) );
NAND2_X1 U773 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
NAND3_X1 U774 ( .A1(n1077), .A2(n1078), .A3(n1079), .ZN(n1076) );
INV_X1 U775 ( .A(n1080), .ZN(n1079) );
NAND2_X1 U776 ( .A1(n1073), .A2(n1081), .ZN(n1075) );
NAND3_X1 U777 ( .A1(n1069), .A2(n1082), .A3(G953), .ZN(n1081) );
INV_X1 U778 ( .A(KEYINPUT26), .ZN(n1082) );
NAND2_X1 U779 ( .A1(n1083), .A2(G227), .ZN(n1069) );
XOR2_X1 U780 ( .A(n1084), .B(KEYINPUT46), .Z(n1083) );
INV_X1 U781 ( .A(n1072), .ZN(n1073) );
NAND3_X1 U782 ( .A1(n1080), .A2(n1085), .A3(n1086), .ZN(n1072) );
XOR2_X1 U783 ( .A(n1087), .B(KEYINPUT5), .Z(n1086) );
NAND2_X1 U784 ( .A1(n1078), .A2(n1077), .ZN(n1087) );
NAND2_X1 U785 ( .A1(n1088), .A2(n1089), .ZN(n1077) );
INV_X1 U786 ( .A(n1090), .ZN(n1088) );
NAND2_X1 U787 ( .A1(G953), .A2(n1084), .ZN(n1085) );
XOR2_X1 U788 ( .A(n1091), .B(n1092), .Z(n1080) );
XOR2_X1 U789 ( .A(n1093), .B(n1094), .Z(n1092) );
XNOR2_X1 U790 ( .A(KEYINPUT1), .B(n1095), .ZN(n1091) );
NOR2_X1 U791 ( .A1(KEYINPUT11), .A2(n1096), .ZN(n1095) );
XOR2_X1 U792 ( .A(n1097), .B(n1098), .Z(G69) );
XOR2_X1 U793 ( .A(n1099), .B(n1100), .Z(n1098) );
NOR2_X1 U794 ( .A1(n1101), .A2(G953), .ZN(n1100) );
AND3_X1 U795 ( .A1(n1102), .A2(n1103), .A3(n1104), .ZN(n1101) );
OR2_X1 U796 ( .A1(n1105), .A2(n1106), .ZN(n1099) );
NAND2_X1 U797 ( .A1(G953), .A2(n1107), .ZN(n1097) );
NAND2_X1 U798 ( .A1(G898), .A2(G224), .ZN(n1107) );
NOR2_X1 U799 ( .A1(n1108), .A2(n1109), .ZN(G66) );
NOR3_X1 U800 ( .A1(n1063), .A2(n1110), .A3(n1111), .ZN(n1109) );
NOR3_X1 U801 ( .A1(n1112), .A2(n1113), .A3(n1114), .ZN(n1111) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(n1110) );
NOR2_X1 U803 ( .A1(n1117), .A2(n1113), .ZN(n1115) );
NOR2_X1 U804 ( .A1(n1108), .A2(n1118), .ZN(G63) );
NOR3_X1 U805 ( .A1(n1062), .A2(n1119), .A3(n1120), .ZN(n1118) );
NOR3_X1 U806 ( .A1(n1121), .A2(n1122), .A3(n1114), .ZN(n1120) );
INV_X1 U807 ( .A(n1123), .ZN(n1121) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1123), .ZN(n1119) );
NOR2_X1 U809 ( .A1(n1117), .A2(n1122), .ZN(n1124) );
INV_X1 U810 ( .A(G478), .ZN(n1122) );
INV_X1 U811 ( .A(n999), .ZN(n1117) );
NOR2_X1 U812 ( .A1(n1108), .A2(n1125), .ZN(G60) );
XOR2_X1 U813 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U814 ( .A1(n1128), .A2(n1114), .ZN(n1127) );
INV_X1 U815 ( .A(G475), .ZN(n1128) );
NOR2_X1 U816 ( .A1(KEYINPUT40), .A2(n1129), .ZN(n1126) );
XOR2_X1 U817 ( .A(KEYINPUT56), .B(n1130), .Z(n1129) );
NAND2_X1 U818 ( .A1(n1131), .A2(n1132), .ZN(G6) );
NAND2_X1 U819 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U820 ( .A1(n1135), .A2(n1136), .ZN(n1133) );
NAND2_X1 U821 ( .A1(KEYINPUT49), .A2(n1137), .ZN(n1136) );
INV_X1 U822 ( .A(KEYINPUT54), .ZN(n1137) );
NAND3_X1 U823 ( .A1(n1138), .A2(n1139), .A3(KEYINPUT54), .ZN(n1131) );
OR2_X1 U824 ( .A1(G104), .A2(KEYINPUT49), .ZN(n1139) );
NAND2_X1 U825 ( .A1(KEYINPUT49), .A2(n1140), .ZN(n1138) );
OR2_X1 U826 ( .A1(n1134), .A2(G104), .ZN(n1140) );
NOR2_X1 U827 ( .A1(n1108), .A2(n1141), .ZN(G57) );
XOR2_X1 U828 ( .A(n1142), .B(n1143), .Z(n1141) );
XOR2_X1 U829 ( .A(n1144), .B(n1145), .Z(n1143) );
NOR2_X1 U830 ( .A1(KEYINPUT9), .A2(n1146), .ZN(n1145) );
NOR2_X1 U831 ( .A1(KEYINPUT10), .A2(n1147), .ZN(n1144) );
XOR2_X1 U832 ( .A(n1148), .B(n1149), .Z(n1147) );
NAND2_X1 U833 ( .A1(KEYINPUT6), .A2(n1150), .ZN(n1148) );
NAND3_X1 U834 ( .A1(G472), .A2(n999), .A3(n1151), .ZN(n1142) );
XOR2_X1 U835 ( .A(n1152), .B(KEYINPUT36), .Z(n1151) );
NOR2_X1 U836 ( .A1(n1108), .A2(n1153), .ZN(G54) );
XOR2_X1 U837 ( .A(n1154), .B(n1155), .Z(n1153) );
XOR2_X1 U838 ( .A(n1156), .B(n1157), .Z(n1155) );
NOR2_X1 U839 ( .A1(n1158), .A2(n1114), .ZN(n1157) );
INV_X1 U840 ( .A(G469), .ZN(n1158) );
NAND2_X1 U841 ( .A1(n1159), .A2(n1160), .ZN(n1156) );
INV_X1 U842 ( .A(n1161), .ZN(n1160) );
NAND2_X1 U843 ( .A1(n1162), .A2(n1163), .ZN(n1159) );
NOR2_X1 U844 ( .A1(n1108), .A2(n1164), .ZN(G51) );
XOR2_X1 U845 ( .A(n1165), .B(n1166), .Z(n1164) );
XOR2_X1 U846 ( .A(n1167), .B(n1105), .Z(n1166) );
NOR2_X1 U847 ( .A1(n1168), .A2(n1114), .ZN(n1167) );
NAND2_X1 U848 ( .A1(G902), .A2(n999), .ZN(n1114) );
NAND4_X1 U849 ( .A1(n1169), .A2(n1170), .A3(n1102), .A4(n1171), .ZN(n999) );
NOR2_X1 U850 ( .A1(n1090), .A2(n1172), .ZN(n1171) );
XNOR2_X1 U851 ( .A(KEYINPUT55), .B(n1104), .ZN(n1172) );
NAND4_X1 U852 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1090) );
AND3_X1 U853 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
NAND2_X1 U854 ( .A1(n1020), .A2(n1180), .ZN(n1175) );
NAND2_X1 U855 ( .A1(n1181), .A2(n1182), .ZN(n1180) );
NAND4_X1 U856 ( .A1(n1183), .A2(n1032), .A3(n1184), .A4(n1185), .ZN(n1182) );
XOR2_X1 U857 ( .A(KEYINPUT47), .B(n1039), .Z(n1184) );
XOR2_X1 U858 ( .A(n1186), .B(KEYINPUT7), .Z(n1181) );
AND4_X1 U859 ( .A1(n1187), .A2(n1188), .A3(n1134), .A4(n1189), .ZN(n1102) );
AND3_X1 U860 ( .A1(n992), .A2(n1190), .A3(n1191), .ZN(n1189) );
NAND3_X1 U861 ( .A1(n1032), .A2(n1192), .A3(n1039), .ZN(n992) );
NAND3_X1 U862 ( .A1(n1039), .A2(n1192), .A3(n1031), .ZN(n1134) );
XNOR2_X1 U863 ( .A(KEYINPUT37), .B(n1089), .ZN(n1170) );
XNOR2_X1 U864 ( .A(KEYINPUT23), .B(n1103), .ZN(n1169) );
XNOR2_X1 U865 ( .A(n1193), .B(n1194), .ZN(n1165) );
NAND2_X1 U866 ( .A1(KEYINPUT8), .A2(n1195), .ZN(n1193) );
NOR2_X1 U867 ( .A1(n1078), .A2(G952), .ZN(n1108) );
XOR2_X1 U868 ( .A(G146), .B(n1196), .Z(G48) );
NOR2_X1 U869 ( .A1(n1197), .A2(n1186), .ZN(n1196) );
NAND4_X1 U870 ( .A1(n1183), .A2(n1031), .A3(n1039), .A4(n1185), .ZN(n1186) );
XNOR2_X1 U871 ( .A(G143), .B(n1173), .ZN(G45) );
NAND3_X1 U872 ( .A1(n1042), .A2(n1198), .A3(n1199), .ZN(n1173) );
NOR3_X1 U873 ( .A1(n1025), .A2(n1200), .A3(n1201), .ZN(n1199) );
XNOR2_X1 U874 ( .A(G140), .B(n1174), .ZN(G42) );
NAND2_X1 U875 ( .A1(n1202), .A2(n1203), .ZN(n1174) );
XNOR2_X1 U876 ( .A(G137), .B(n1177), .ZN(G39) );
NAND3_X1 U877 ( .A1(n1183), .A2(n1202), .A3(n1033), .ZN(n1177) );
XOR2_X1 U878 ( .A(n1179), .B(n1204), .Z(G36) );
XOR2_X1 U879 ( .A(KEYINPUT42), .B(G134), .Z(n1204) );
NAND3_X1 U880 ( .A1(n1202), .A2(n1032), .A3(n1042), .ZN(n1179) );
XOR2_X1 U881 ( .A(n1205), .B(G131), .Z(G33) );
NAND2_X1 U882 ( .A1(KEYINPUT12), .A2(n1089), .ZN(n1205) );
NAND3_X1 U883 ( .A1(n1202), .A2(n1031), .A3(n1042), .ZN(n1089) );
AND3_X1 U884 ( .A1(n1039), .A2(n1185), .A3(n1028), .ZN(n1202) );
NOR2_X1 U885 ( .A1(n1023), .A2(n1059), .ZN(n1028) );
INV_X1 U886 ( .A(n1024), .ZN(n1059) );
XOR2_X1 U887 ( .A(n1206), .B(n1207), .Z(G30) );
NAND4_X1 U888 ( .A1(n1198), .A2(n1039), .A3(n1032), .A4(n1208), .ZN(n1207) );
XOR2_X1 U889 ( .A(KEYINPUT45), .B(n1183), .Z(n1208) );
XOR2_X1 U890 ( .A(n1209), .B(n1187), .Z(G3) );
NAND4_X1 U891 ( .A1(n1033), .A2(n1042), .A3(n1039), .A4(n1210), .ZN(n1187) );
XNOR2_X1 U892 ( .A(G125), .B(n1178), .ZN(G27) );
NAND3_X1 U893 ( .A1(n1198), .A2(n1203), .A3(n1029), .ZN(n1178) );
AND3_X1 U894 ( .A1(n1211), .A2(n1008), .A3(n1031), .ZN(n1203) );
AND2_X1 U895 ( .A1(n1020), .A2(n1185), .ZN(n1198) );
NAND2_X1 U896 ( .A1(n1002), .A2(n1212), .ZN(n1185) );
NAND4_X1 U897 ( .A1(G902), .A2(G953), .A3(n1213), .A4(n1084), .ZN(n1212) );
INV_X1 U898 ( .A(G900), .ZN(n1084) );
XOR2_X1 U899 ( .A(n1188), .B(n1214), .Z(G24) );
XOR2_X1 U900 ( .A(KEYINPUT38), .B(G122), .Z(n1214) );
NAND4_X1 U901 ( .A1(n1029), .A2(n1192), .A3(n1215), .A4(n1216), .ZN(n1188) );
AND3_X1 U902 ( .A1(n1211), .A2(n1041), .A3(n1210), .ZN(n1192) );
XOR2_X1 U903 ( .A(n1104), .B(n1217), .Z(G21) );
XOR2_X1 U904 ( .A(KEYINPUT17), .B(G119), .Z(n1217) );
NAND3_X1 U905 ( .A1(n1033), .A2(n1183), .A3(n1218), .ZN(n1104) );
NOR2_X1 U906 ( .A1(n1041), .A2(n1211), .ZN(n1183) );
INV_X1 U907 ( .A(n1008), .ZN(n1041) );
INV_X1 U908 ( .A(n1014), .ZN(n1033) );
XOR2_X1 U909 ( .A(n1219), .B(n1191), .Z(G18) );
NAND3_X1 U910 ( .A1(n1042), .A2(n1032), .A3(n1218), .ZN(n1191) );
NOR2_X1 U911 ( .A1(n1215), .A2(n1200), .ZN(n1032) );
INV_X1 U912 ( .A(n1201), .ZN(n1215) );
XNOR2_X1 U913 ( .A(G113), .B(n1190), .ZN(G15) );
NAND3_X1 U914 ( .A1(n1042), .A2(n1031), .A3(n1218), .ZN(n1190) );
AND2_X1 U915 ( .A1(n1029), .A2(n1210), .ZN(n1218) );
INV_X1 U916 ( .A(n1018), .ZN(n1029) );
NAND2_X1 U917 ( .A1(n1037), .A2(n1220), .ZN(n1018) );
NOR2_X1 U918 ( .A1(n1216), .A2(n1201), .ZN(n1031) );
NOR2_X1 U919 ( .A1(n1008), .A2(n1211), .ZN(n1042) );
XOR2_X1 U920 ( .A(n1221), .B(n1103), .Z(G12) );
NAND4_X1 U921 ( .A1(n1211), .A2(n1008), .A3(n1210), .A4(n1222), .ZN(n1103) );
NOR2_X1 U922 ( .A1(n1025), .A2(n1014), .ZN(n1222) );
NAND2_X1 U923 ( .A1(n1200), .A2(n1201), .ZN(n1014) );
XOR2_X1 U924 ( .A(n1053), .B(G475), .Z(n1201) );
OR2_X1 U925 ( .A1(n1130), .A2(G902), .ZN(n1053) );
XNOR2_X1 U926 ( .A(n1223), .B(n1224), .ZN(n1130) );
XOR2_X1 U927 ( .A(n1225), .B(n1226), .Z(n1224) );
NAND2_X1 U928 ( .A1(KEYINPUT30), .A2(n1093), .ZN(n1225) );
XOR2_X1 U929 ( .A(n1227), .B(n1228), .Z(n1223) );
NOR2_X1 U930 ( .A1(KEYINPUT29), .A2(n1229), .ZN(n1228) );
XOR2_X1 U931 ( .A(n1135), .B(n1230), .Z(n1229) );
NAND2_X1 U932 ( .A1(KEYINPUT2), .A2(n1231), .ZN(n1230) );
XOR2_X1 U933 ( .A(G122), .B(G113), .Z(n1231) );
NAND2_X1 U934 ( .A1(n1232), .A2(n1233), .ZN(n1227) );
NAND3_X1 U935 ( .A1(n1234), .A2(G143), .A3(G214), .ZN(n1233) );
NAND2_X1 U936 ( .A1(n1235), .A2(n1236), .ZN(n1232) );
NAND2_X1 U937 ( .A1(G214), .A2(n1234), .ZN(n1236) );
XNOR2_X1 U938 ( .A(G143), .B(KEYINPUT34), .ZN(n1235) );
INV_X1 U939 ( .A(n1216), .ZN(n1200) );
XOR2_X1 U940 ( .A(n1062), .B(G478), .Z(n1216) );
NOR2_X1 U941 ( .A1(n1123), .A2(G902), .ZN(n1062) );
XOR2_X1 U942 ( .A(n1237), .B(n1238), .Z(n1123) );
NOR2_X1 U943 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
INV_X1 U944 ( .A(G217), .ZN(n1240) );
NAND2_X1 U945 ( .A1(n1241), .A2(KEYINPUT60), .ZN(n1237) );
XOR2_X1 U946 ( .A(n1242), .B(n1243), .Z(n1241) );
NOR2_X1 U947 ( .A1(KEYINPUT31), .A2(n1244), .ZN(n1243) );
XOR2_X1 U948 ( .A(n1245), .B(n1246), .Z(n1244) );
NOR2_X1 U949 ( .A1(KEYINPUT61), .A2(G143), .ZN(n1246) );
XOR2_X1 U950 ( .A(G134), .B(n1206), .Z(n1245) );
INV_X1 U951 ( .A(G128), .ZN(n1206) );
NAND2_X1 U952 ( .A1(n1247), .A2(n1248), .ZN(n1242) );
OR2_X1 U953 ( .A1(n1249), .A2(n994), .ZN(n1248) );
XOR2_X1 U954 ( .A(n1250), .B(KEYINPUT15), .Z(n1247) );
NAND2_X1 U955 ( .A1(n1249), .A2(n994), .ZN(n1250) );
XNOR2_X1 U956 ( .A(n1251), .B(G122), .ZN(n1249) );
NAND2_X1 U957 ( .A1(KEYINPUT41), .A2(n1219), .ZN(n1251) );
INV_X1 U958 ( .A(n1039), .ZN(n1025) );
NOR2_X1 U959 ( .A1(n1037), .A2(n1038), .ZN(n1039) );
INV_X1 U960 ( .A(n1220), .ZN(n1038) );
NAND2_X1 U961 ( .A1(G221), .A2(n1252), .ZN(n1220) );
XNOR2_X1 U962 ( .A(n1054), .B(KEYINPUT33), .ZN(n1037) );
XOR2_X1 U963 ( .A(n1253), .B(G469), .Z(n1054) );
NAND2_X1 U964 ( .A1(n1254), .A2(n1152), .ZN(n1253) );
XOR2_X1 U965 ( .A(n1154), .B(n1255), .Z(n1254) );
NOR2_X1 U966 ( .A1(n1161), .A2(n1256), .ZN(n1255) );
NOR2_X1 U967 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
XNOR2_X1 U968 ( .A(n1259), .B(n1163), .ZN(n1258) );
XNOR2_X1 U969 ( .A(KEYINPUT43), .B(KEYINPUT22), .ZN(n1259) );
INV_X1 U970 ( .A(n1162), .ZN(n1257) );
NOR2_X1 U971 ( .A1(n1163), .A2(n1162), .ZN(n1161) );
XOR2_X1 U972 ( .A(G140), .B(G110), .Z(n1162) );
NAND2_X1 U973 ( .A1(G227), .A2(n1078), .ZN(n1163) );
XOR2_X1 U974 ( .A(n1260), .B(n1261), .Z(n1154) );
NOR2_X1 U975 ( .A1(n1262), .A2(n1263), .ZN(n1261) );
NOR3_X1 U976 ( .A1(KEYINPUT13), .A2(G107), .A3(n1135), .ZN(n1263) );
NOR2_X1 U977 ( .A1(n1264), .A2(n1265), .ZN(n1262) );
INV_X1 U978 ( .A(KEYINPUT13), .ZN(n1265) );
XOR2_X1 U979 ( .A(n1150), .B(n1209), .Z(n1260) );
AND2_X1 U980 ( .A1(n1020), .A2(n1266), .ZN(n1210) );
NAND2_X1 U981 ( .A1(n1002), .A2(n1267), .ZN(n1266) );
NAND3_X1 U982 ( .A1(n1106), .A2(n1213), .A3(G902), .ZN(n1267) );
NOR2_X1 U983 ( .A1(n1078), .A2(G898), .ZN(n1106) );
NAND3_X1 U984 ( .A1(n1066), .A2(n1213), .A3(G952), .ZN(n1002) );
NAND2_X1 U985 ( .A1(G237), .A2(G234), .ZN(n1213) );
XOR2_X1 U986 ( .A(n1078), .B(KEYINPUT53), .Z(n1066) );
INV_X1 U987 ( .A(n1197), .ZN(n1020) );
NAND2_X1 U988 ( .A1(n1023), .A2(n1024), .ZN(n1197) );
NAND2_X1 U989 ( .A1(G214), .A2(n1268), .ZN(n1024) );
XNOR2_X1 U990 ( .A(n1049), .B(KEYINPUT28), .ZN(n1023) );
XOR2_X1 U991 ( .A(n1269), .B(n1168), .Z(n1049) );
NAND2_X1 U992 ( .A1(G210), .A2(n1268), .ZN(n1168) );
NAND2_X1 U993 ( .A1(n1270), .A2(n1152), .ZN(n1268) );
INV_X1 U994 ( .A(G237), .ZN(n1270) );
NAND2_X1 U995 ( .A1(n1271), .A2(n1152), .ZN(n1269) );
XNOR2_X1 U996 ( .A(n1105), .B(n1272), .ZN(n1271) );
XOR2_X1 U997 ( .A(KEYINPUT24), .B(n1273), .Z(n1272) );
NOR2_X1 U998 ( .A1(n1274), .A2(n1275), .ZN(n1273) );
XOR2_X1 U999 ( .A(n1276), .B(KEYINPUT14), .Z(n1275) );
NAND2_X1 U1000 ( .A1(n1195), .A2(n1194), .ZN(n1276) );
NOR2_X1 U1001 ( .A1(n1195), .A2(n1194), .ZN(n1274) );
NAND2_X1 U1002 ( .A1(G224), .A2(n1078), .ZN(n1194) );
XNOR2_X1 U1003 ( .A(n1277), .B(n1278), .ZN(n1195) );
XNOR2_X1 U1004 ( .A(G125), .B(G146), .ZN(n1277) );
XNOR2_X1 U1005 ( .A(n1279), .B(n1280), .ZN(n1105) );
XNOR2_X1 U1006 ( .A(n1281), .B(n1264), .ZN(n1280) );
XOR2_X1 U1007 ( .A(n994), .B(n1135), .Z(n1264) );
INV_X1 U1008 ( .A(G104), .ZN(n1135) );
INV_X1 U1009 ( .A(G107), .ZN(n994) );
NAND2_X1 U1010 ( .A1(n1282), .A2(n1283), .ZN(n1281) );
NAND2_X1 U1011 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U1012 ( .A(n1286), .B(KEYINPUT0), .Z(n1282) );
OR2_X1 U1013 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
XOR2_X1 U1014 ( .A(G113), .B(KEYINPUT44), .Z(n1285) );
XOR2_X1 U1015 ( .A(n1209), .B(n1287), .Z(n1279) );
XOR2_X1 U1016 ( .A(G122), .B(G110), .Z(n1287) );
XOR2_X1 U1017 ( .A(n1063), .B(n1065), .Z(n1008) );
INV_X1 U1018 ( .A(n1113), .ZN(n1065) );
NAND2_X1 U1019 ( .A1(G217), .A2(n1252), .ZN(n1113) );
NAND2_X1 U1020 ( .A1(G234), .A2(n1152), .ZN(n1252) );
NOR2_X1 U1021 ( .A1(n1116), .A2(G902), .ZN(n1063) );
INV_X1 U1022 ( .A(n1112), .ZN(n1116) );
XOR2_X1 U1023 ( .A(n1288), .B(n1289), .Z(n1112) );
XOR2_X1 U1024 ( .A(n1290), .B(n1291), .Z(n1289) );
NOR2_X1 U1025 ( .A1(KEYINPUT58), .A2(n1292), .ZN(n1291) );
XOR2_X1 U1026 ( .A(n1221), .B(n1293), .Z(n1292) );
XOR2_X1 U1027 ( .A(G128), .B(G119), .Z(n1293) );
NOR2_X1 U1028 ( .A1(n1294), .A2(n1295), .ZN(n1290) );
XOR2_X1 U1029 ( .A(KEYINPUT62), .B(KEYINPUT50), .Z(n1295) );
XOR2_X1 U1030 ( .A(n1296), .B(n1297), .Z(n1294) );
XNOR2_X1 U1031 ( .A(KEYINPUT20), .B(n1298), .ZN(n1296) );
NOR3_X1 U1032 ( .A1(n1239), .A2(KEYINPUT48), .A3(n1299), .ZN(n1298) );
INV_X1 U1033 ( .A(G221), .ZN(n1299) );
NAND2_X1 U1034 ( .A1(G234), .A2(n1078), .ZN(n1239) );
INV_X1 U1035 ( .A(G953), .ZN(n1078) );
XNOR2_X1 U1036 ( .A(n1093), .B(n1300), .ZN(n1288) );
NOR2_X1 U1037 ( .A1(G146), .A2(KEYINPUT57), .ZN(n1300) );
XOR2_X1 U1038 ( .A(G125), .B(G140), .Z(n1093) );
INV_X1 U1039 ( .A(n1005), .ZN(n1211) );
XOR2_X1 U1040 ( .A(n1056), .B(G472), .Z(n1005) );
AND2_X1 U1041 ( .A1(n1301), .A2(n1152), .ZN(n1056) );
INV_X1 U1042 ( .A(G902), .ZN(n1152) );
XOR2_X1 U1043 ( .A(n1302), .B(n1303), .Z(n1301) );
XOR2_X1 U1044 ( .A(KEYINPUT59), .B(n1304), .Z(n1303) );
INV_X1 U1045 ( .A(n1149), .ZN(n1304) );
XNOR2_X1 U1046 ( .A(G113), .B(n1305), .ZN(n1149) );
NOR2_X1 U1047 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NOR3_X1 U1048 ( .A1(KEYINPUT25), .A2(G119), .A3(n1219), .ZN(n1307) );
INV_X1 U1049 ( .A(G116), .ZN(n1219) );
AND2_X1 U1050 ( .A1(n1284), .A2(KEYINPUT25), .ZN(n1306) );
XNOR2_X1 U1051 ( .A(G116), .B(G119), .ZN(n1284) );
XNOR2_X1 U1052 ( .A(n1150), .B(n1146), .ZN(n1302) );
AND2_X1 U1053 ( .A1(n1308), .A2(n1309), .ZN(n1146) );
NAND2_X1 U1054 ( .A1(n1310), .A2(n1209), .ZN(n1309) );
INV_X1 U1055 ( .A(G101), .ZN(n1209) );
NAND2_X1 U1056 ( .A1(G210), .A2(n1234), .ZN(n1310) );
NAND3_X1 U1057 ( .A1(G210), .A2(n1234), .A3(G101), .ZN(n1308) );
NOR2_X1 U1058 ( .A1(G237), .A2(G953), .ZN(n1234) );
XNOR2_X1 U1059 ( .A(n1096), .B(n1094), .ZN(n1150) );
XNOR2_X1 U1060 ( .A(n1226), .B(n1278), .ZN(n1094) );
XOR2_X1 U1061 ( .A(G128), .B(G143), .Z(n1278) );
XNOR2_X1 U1062 ( .A(G131), .B(G146), .ZN(n1226) );
XNOR2_X1 U1063 ( .A(G134), .B(n1297), .ZN(n1096) );
XOR2_X1 U1064 ( .A(G137), .B(KEYINPUT51), .Z(n1297) );
INV_X1 U1065 ( .A(G110), .ZN(n1221) );
endmodule


