//Key = 1010111000000100100000010101111011000100101000101011111000110111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;

XNOR2_X1 U706 ( .A(n970), .B(n971), .ZN(G9) );
NOR2_X1 U707 ( .A1(n972), .A2(n973), .ZN(G75) );
NOR4_X1 U708 ( .A1(n974), .A2(n975), .A3(n976), .A4(n977), .ZN(n973) );
XOR2_X1 U709 ( .A(n978), .B(KEYINPUT23), .Z(n977) );
NAND3_X1 U710 ( .A1(n979), .A2(n980), .A3(n981), .ZN(n978) );
INV_X1 U711 ( .A(n982), .ZN(n980) );
NOR3_X1 U712 ( .A1(n983), .A2(n984), .A3(n982), .ZN(n976) );
NOR2_X1 U713 ( .A1(n985), .A2(n986), .ZN(n984) );
NOR2_X1 U714 ( .A1(n987), .A2(n988), .ZN(n986) );
NOR3_X1 U715 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n987) );
NOR2_X1 U716 ( .A1(n992), .A2(n993), .ZN(n991) );
XNOR2_X1 U717 ( .A(n994), .B(KEYINPUT57), .ZN(n992) );
NOR4_X1 U718 ( .A1(KEYINPUT26), .A2(n995), .A3(n996), .A4(n997), .ZN(n990) );
NOR2_X1 U719 ( .A1(n998), .A2(n999), .ZN(n989) );
NOR3_X1 U720 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n998) );
AND2_X1 U721 ( .A1(n994), .A2(KEYINPUT26), .ZN(n1002) );
NOR2_X1 U722 ( .A1(n1003), .A2(n1004), .ZN(n1000) );
NOR3_X1 U723 ( .A1(n1005), .A2(n1006), .A3(n999), .ZN(n985) );
XNOR2_X1 U724 ( .A(KEYINPUT4), .B(n995), .ZN(n1005) );
NAND3_X1 U725 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n974) );
NAND3_X1 U726 ( .A1(n1010), .A2(n1011), .A3(n981), .ZN(n1009) );
NOR3_X1 U727 ( .A1(n999), .A2(n995), .A3(n983), .ZN(n981) );
NAND2_X1 U728 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
NOR3_X1 U729 ( .A1(n1014), .A2(G953), .A3(G952), .ZN(n972) );
INV_X1 U730 ( .A(n1007), .ZN(n1014) );
NAND4_X1 U731 ( .A1(n997), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1007) );
NOR2_X1 U732 ( .A1(n1018), .A2(n995), .ZN(n1017) );
XOR2_X1 U733 ( .A(n1019), .B(KEYINPUT35), .Z(n1018) );
NAND4_X1 U734 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019) );
XOR2_X1 U735 ( .A(n1024), .B(n1025), .Z(n1022) );
NOR2_X1 U736 ( .A1(n1026), .A2(KEYINPUT9), .ZN(n1025) );
INV_X1 U737 ( .A(n1027), .ZN(n1026) );
XOR2_X1 U738 ( .A(n1028), .B(KEYINPUT33), .Z(n1024) );
XNOR2_X1 U739 ( .A(n1029), .B(n1030), .ZN(n1021) );
XOR2_X1 U740 ( .A(n1031), .B(KEYINPUT61), .Z(n1020) );
NAND2_X1 U741 ( .A1(n1032), .A2(n1033), .ZN(n1031) );
NAND2_X1 U742 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
XNOR2_X1 U743 ( .A(KEYINPUT6), .B(n1036), .ZN(n1035) );
XNOR2_X1 U744 ( .A(n1037), .B(KEYINPUT22), .ZN(n1034) );
OR2_X1 U745 ( .A1(n1036), .A2(n1038), .ZN(n1032) );
XOR2_X1 U746 ( .A(n1039), .B(n1040), .Z(G72) );
NOR2_X1 U747 ( .A1(n1041), .A2(n1008), .ZN(n1040) );
AND2_X1 U748 ( .A1(G227), .A2(G900), .ZN(n1041) );
NAND2_X1 U749 ( .A1(n1042), .A2(KEYINPUT25), .ZN(n1039) );
XOR2_X1 U750 ( .A(n1043), .B(n1044), .Z(n1042) );
NOR2_X1 U751 ( .A1(n1045), .A2(G953), .ZN(n1044) );
NAND2_X1 U752 ( .A1(n1046), .A2(n1047), .ZN(n1043) );
XOR2_X1 U753 ( .A(n1048), .B(n1049), .Z(n1047) );
XOR2_X1 U754 ( .A(n1050), .B(n1051), .Z(n1049) );
XNOR2_X1 U755 ( .A(n1052), .B(n1053), .ZN(n1048) );
XNOR2_X1 U756 ( .A(KEYINPUT40), .B(KEYINPUT21), .ZN(n1052) );
XOR2_X1 U757 ( .A(n1054), .B(KEYINPUT34), .Z(n1046) );
NAND2_X1 U758 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U759 ( .A(n1057), .B(n1058), .Z(G69) );
NAND2_X1 U760 ( .A1(G953), .A2(n1059), .ZN(n1058) );
NAND2_X1 U761 ( .A1(G898), .A2(G224), .ZN(n1059) );
NAND2_X1 U762 ( .A1(n1060), .A2(KEYINPUT54), .ZN(n1057) );
XOR2_X1 U763 ( .A(n1061), .B(n1062), .Z(n1060) );
NOR2_X1 U764 ( .A1(KEYINPUT39), .A2(n1063), .ZN(n1062) );
NOR2_X1 U765 ( .A1(n1064), .A2(G953), .ZN(n1063) );
NAND2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1061) );
NAND2_X1 U767 ( .A1(n1055), .A2(n1067), .ZN(n1066) );
XNOR2_X1 U768 ( .A(n1068), .B(n1069), .ZN(n1065) );
XNOR2_X1 U769 ( .A(G110), .B(n1070), .ZN(n1068) );
NOR2_X1 U770 ( .A1(KEYINPUT10), .A2(n1071), .ZN(n1070) );
XOR2_X1 U771 ( .A(n1072), .B(n1073), .Z(n1071) );
NOR2_X1 U772 ( .A1(KEYINPUT8), .A2(n1074), .ZN(n1072) );
XNOR2_X1 U773 ( .A(n970), .B(n1075), .ZN(n1074) );
NOR2_X1 U774 ( .A1(n1076), .A2(n1077), .ZN(G66) );
XOR2_X1 U775 ( .A(n1078), .B(n1079), .Z(n1077) );
NOR2_X1 U776 ( .A1(n1027), .A2(n1080), .ZN(n1078) );
NOR2_X1 U777 ( .A1(n1076), .A2(n1081), .ZN(G63) );
XOR2_X1 U778 ( .A(n1082), .B(n1083), .Z(n1081) );
NOR2_X1 U779 ( .A1(n1084), .A2(KEYINPUT44), .ZN(n1082) );
NOR2_X1 U780 ( .A1(n1085), .A2(n1080), .ZN(n1084) );
INV_X1 U781 ( .A(G478), .ZN(n1085) );
NOR2_X1 U782 ( .A1(n1076), .A2(n1086), .ZN(G60) );
XNOR2_X1 U783 ( .A(n1087), .B(n1088), .ZN(n1086) );
NOR2_X1 U784 ( .A1(n1089), .A2(n1080), .ZN(n1088) );
XNOR2_X1 U785 ( .A(G104), .B(n1090), .ZN(G6) );
NOR2_X1 U786 ( .A1(n1076), .A2(n1091), .ZN(G57) );
XOR2_X1 U787 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U788 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U789 ( .A1(KEYINPUT55), .A2(n1096), .ZN(n1095) );
NOR2_X1 U790 ( .A1(n1097), .A2(n1098), .ZN(n1094) );
XOR2_X1 U791 ( .A(n1099), .B(KEYINPUT50), .Z(n1098) );
NAND2_X1 U792 ( .A1(n1100), .A2(n1073), .ZN(n1099) );
NOR2_X1 U793 ( .A1(n1073), .A2(n1100), .ZN(n1097) );
NOR2_X1 U794 ( .A1(n1030), .A2(n1080), .ZN(n1092) );
NOR2_X1 U795 ( .A1(n1076), .A2(n1101), .ZN(G54) );
XNOR2_X1 U796 ( .A(n1102), .B(n1103), .ZN(n1101) );
NOR2_X1 U797 ( .A1(n1104), .A2(n1080), .ZN(n1103) );
NAND2_X1 U798 ( .A1(G902), .A2(n975), .ZN(n1080) );
INV_X1 U799 ( .A(G469), .ZN(n1104) );
NOR2_X1 U800 ( .A1(n1076), .A2(n1105), .ZN(G51) );
XOR2_X1 U801 ( .A(KEYINPUT1), .B(n1106), .Z(n1105) );
NOR2_X1 U802 ( .A1(n1107), .A2(n1108), .ZN(n1106) );
XOR2_X1 U803 ( .A(n1109), .B(KEYINPUT13), .Z(n1108) );
NAND2_X1 U804 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NOR2_X1 U805 ( .A1(n1111), .A2(n1110), .ZN(n1107) );
XOR2_X1 U806 ( .A(KEYINPUT60), .B(n1112), .Z(n1110) );
NAND4_X1 U807 ( .A1(G210), .A2(n1113), .A3(n975), .A4(n1114), .ZN(n1111) );
NAND2_X1 U808 ( .A1(n1045), .A2(n1064), .ZN(n975) );
AND4_X1 U809 ( .A1(n1115), .A2(n1116), .A3(n1090), .A4(n1117), .ZN(n1064) );
NOR4_X1 U810 ( .A1(n1118), .A2(n1119), .A3(n971), .A4(n1120), .ZN(n1117) );
INV_X1 U811 ( .A(n1121), .ZN(n1120) );
NOR3_X1 U812 ( .A1(n982), .A2(n1122), .A3(n1123), .ZN(n971) );
NOR2_X1 U813 ( .A1(n1124), .A2(n1013), .ZN(n1119) );
NOR2_X1 U814 ( .A1(n1125), .A2(n1126), .ZN(n1124) );
NOR2_X1 U815 ( .A1(n1123), .A2(n1127), .ZN(n1126) );
NOR2_X1 U816 ( .A1(n1122), .A2(n1128), .ZN(n1125) );
XNOR2_X1 U817 ( .A(KEYINPUT28), .B(n988), .ZN(n1128) );
OR3_X1 U818 ( .A1(n982), .A2(n1122), .A3(n1006), .ZN(n1090) );
AND2_X1 U819 ( .A1(n1129), .A2(n1130), .ZN(n1045) );
AND4_X1 U820 ( .A1(n1131), .A2(n1132), .A3(n1133), .A4(n1134), .ZN(n1130) );
AND4_X1 U821 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1129) );
OR2_X1 U822 ( .A1(n1012), .A2(n1139), .ZN(n1138) );
XNOR2_X1 U823 ( .A(KEYINPUT11), .B(n1140), .ZN(n1113) );
NOR2_X1 U824 ( .A1(n1008), .A2(G952), .ZN(n1076) );
XNOR2_X1 U825 ( .A(G146), .B(n1131), .ZN(G48) );
NAND4_X1 U826 ( .A1(n1141), .A2(n1142), .A3(n1001), .A4(n1143), .ZN(n1131) );
XNOR2_X1 U827 ( .A(G143), .B(n1137), .ZN(G45) );
NAND3_X1 U828 ( .A1(n1144), .A2(n1142), .A3(n1145), .ZN(n1137) );
NOR3_X1 U829 ( .A1(n1146), .A2(n1023), .A3(n1147), .ZN(n1145) );
XOR2_X1 U830 ( .A(G140), .B(n1148), .Z(G42) );
NOR2_X1 U831 ( .A1(n1139), .A2(n1149), .ZN(n1148) );
XNOR2_X1 U832 ( .A(KEYINPUT42), .B(n1012), .ZN(n1149) );
INV_X1 U833 ( .A(n1150), .ZN(n1012) );
XOR2_X1 U834 ( .A(n1136), .B(n1151), .Z(G39) );
NAND2_X1 U835 ( .A1(KEYINPUT46), .A2(G137), .ZN(n1151) );
NAND3_X1 U836 ( .A1(n1152), .A2(n1143), .A3(n1010), .ZN(n1136) );
XNOR2_X1 U837 ( .A(G134), .B(n1135), .ZN(G36) );
NAND3_X1 U838 ( .A1(n1152), .A2(n979), .A3(n1144), .ZN(n1135) );
XNOR2_X1 U839 ( .A(G131), .B(n1134), .ZN(G33) );
OR2_X1 U840 ( .A1(n1013), .A2(n1139), .ZN(n1134) );
NAND2_X1 U841 ( .A1(n1152), .A2(n1141), .ZN(n1139) );
AND2_X1 U842 ( .A1(n1142), .A2(n994), .ZN(n1152) );
INV_X1 U843 ( .A(n995), .ZN(n994) );
NAND2_X1 U844 ( .A1(n1153), .A2(n1004), .ZN(n995) );
INV_X1 U845 ( .A(n1003), .ZN(n1153) );
XNOR2_X1 U846 ( .A(G128), .B(n1133), .ZN(G30) );
NAND4_X1 U847 ( .A1(n1142), .A2(n979), .A3(n1001), .A4(n1143), .ZN(n1133) );
AND2_X1 U848 ( .A1(n1154), .A2(n1155), .ZN(n1142) );
XNOR2_X1 U849 ( .A(G101), .B(n1156), .ZN(G3) );
NAND2_X1 U850 ( .A1(n1157), .A2(n1144), .ZN(n1156) );
XNOR2_X1 U851 ( .A(G125), .B(n1132), .ZN(G27) );
NAND4_X1 U852 ( .A1(n1001), .A2(n1155), .A3(n1150), .A4(n1158), .ZN(n1132) );
NOR2_X1 U853 ( .A1(n1006), .A2(n999), .ZN(n1158) );
INV_X1 U854 ( .A(n1141), .ZN(n1006) );
NAND2_X1 U855 ( .A1(n983), .A2(n1159), .ZN(n1155) );
NAND4_X1 U856 ( .A1(n1055), .A2(G902), .A3(n1160), .A4(n1056), .ZN(n1159) );
INV_X1 U857 ( .A(G900), .ZN(n1056) );
XOR2_X1 U858 ( .A(G122), .B(n1118), .Z(G24) );
NOR4_X1 U859 ( .A1(n1127), .A2(n982), .A3(n1147), .A4(n1023), .ZN(n1118) );
NAND2_X1 U860 ( .A1(n1161), .A2(n1162), .ZN(n982) );
XOR2_X1 U861 ( .A(n1163), .B(KEYINPUT20), .Z(n1161) );
XNOR2_X1 U862 ( .A(G119), .B(n1115), .ZN(G21) );
NAND3_X1 U863 ( .A1(n1010), .A2(n1143), .A3(n1164), .ZN(n1115) );
NAND2_X1 U864 ( .A1(n1165), .A2(n1166), .ZN(n1143) );
OR3_X1 U865 ( .A1(n1163), .A2(n1162), .A3(KEYINPUT24), .ZN(n1166) );
NAND2_X1 U866 ( .A1(KEYINPUT24), .A2(n1150), .ZN(n1165) );
INV_X1 U867 ( .A(n988), .ZN(n1010) );
XOR2_X1 U868 ( .A(G116), .B(n1167), .Z(G18) );
NOR3_X1 U869 ( .A1(n1127), .A2(n1168), .A3(n1013), .ZN(n1167) );
XNOR2_X1 U870 ( .A(n979), .B(KEYINPUT56), .ZN(n1168) );
INV_X1 U871 ( .A(n1123), .ZN(n979) );
NAND2_X1 U872 ( .A1(n1169), .A2(n1023), .ZN(n1123) );
INV_X1 U873 ( .A(n1164), .ZN(n1127) );
XNOR2_X1 U874 ( .A(G113), .B(n1116), .ZN(G15) );
NAND3_X1 U875 ( .A1(n1144), .A2(n1141), .A3(n1164), .ZN(n1116) );
NOR3_X1 U876 ( .A1(n1146), .A2(n1170), .A3(n999), .ZN(n1164) );
NAND2_X1 U877 ( .A1(n1171), .A2(n997), .ZN(n999) );
INV_X1 U878 ( .A(n996), .ZN(n1171) );
INV_X1 U879 ( .A(n1172), .ZN(n1170) );
NOR2_X1 U880 ( .A1(n1023), .A2(n1169), .ZN(n1141) );
INV_X1 U881 ( .A(n1147), .ZN(n1169) );
INV_X1 U882 ( .A(n1013), .ZN(n1144) );
NAND2_X1 U883 ( .A1(n1162), .A2(n1173), .ZN(n1013) );
XNOR2_X1 U884 ( .A(KEYINPUT24), .B(n1163), .ZN(n1173) );
XNOR2_X1 U885 ( .A(G110), .B(n1121), .ZN(G12) );
NAND2_X1 U886 ( .A1(n1157), .A2(n1150), .ZN(n1121) );
NOR2_X1 U887 ( .A1(n1174), .A2(n1162), .ZN(n1150) );
XOR2_X1 U888 ( .A(n1028), .B(n1175), .Z(n1162) );
NOR2_X1 U889 ( .A1(KEYINPUT36), .A2(n1027), .ZN(n1175) );
NAND2_X1 U890 ( .A1(G217), .A2(n1176), .ZN(n1027) );
OR2_X1 U891 ( .A1(n1079), .A2(n1177), .ZN(n1028) );
INV_X1 U892 ( .A(n1178), .ZN(n1177) );
XNOR2_X1 U893 ( .A(n1179), .B(n1180), .ZN(n1079) );
NOR3_X1 U894 ( .A1(n1181), .A2(KEYINPUT19), .A3(n1182), .ZN(n1180) );
INV_X1 U895 ( .A(G221), .ZN(n1181) );
XNOR2_X1 U896 ( .A(G137), .B(n1183), .ZN(n1179) );
NOR2_X1 U897 ( .A1(n1184), .A2(n1185), .ZN(n1183) );
XOR2_X1 U898 ( .A(KEYINPUT12), .B(n1186), .Z(n1185) );
NOR2_X1 U899 ( .A1(n1187), .A2(n1188), .ZN(n1186) );
AND2_X1 U900 ( .A1(n1188), .A2(n1187), .ZN(n1184) );
XOR2_X1 U901 ( .A(n1189), .B(n1190), .Z(n1187) );
XNOR2_X1 U902 ( .A(KEYINPUT53), .B(n1191), .ZN(n1190) );
INV_X1 U903 ( .A(G128), .ZN(n1191) );
XNOR2_X1 U904 ( .A(G119), .B(G110), .ZN(n1189) );
NAND3_X1 U905 ( .A1(n1192), .A2(n1193), .A3(n1194), .ZN(n1188) );
NAND2_X1 U906 ( .A1(G146), .A2(n1195), .ZN(n1194) );
OR3_X1 U907 ( .A1(n1195), .A2(G146), .A3(n1196), .ZN(n1193) );
INV_X1 U908 ( .A(KEYINPUT2), .ZN(n1195) );
NAND2_X1 U909 ( .A1(n1196), .A2(n1197), .ZN(n1192) );
NAND2_X1 U910 ( .A1(KEYINPUT2), .A2(n1198), .ZN(n1197) );
XNOR2_X1 U911 ( .A(KEYINPUT52), .B(n1199), .ZN(n1198) );
XOR2_X1 U912 ( .A(G140), .B(G125), .Z(n1196) );
INV_X1 U913 ( .A(n1163), .ZN(n1174) );
XOR2_X1 U914 ( .A(n1029), .B(n1200), .Z(n1163) );
NOR2_X1 U915 ( .A1(KEYINPUT43), .A2(n1030), .ZN(n1200) );
INV_X1 U916 ( .A(G472), .ZN(n1030) );
NAND2_X1 U917 ( .A1(n1201), .A2(n1178), .ZN(n1029) );
XOR2_X1 U918 ( .A(n1096), .B(n1202), .Z(n1201) );
XNOR2_X1 U919 ( .A(n1203), .B(n1073), .ZN(n1202) );
NAND2_X1 U920 ( .A1(KEYINPUT58), .A2(n1100), .ZN(n1203) );
XNOR2_X1 U921 ( .A(n1204), .B(n1199), .ZN(n1100) );
AND2_X1 U922 ( .A1(n1205), .A2(n1206), .ZN(n1096) );
NAND2_X1 U923 ( .A1(n1207), .A2(n1208), .ZN(n1206) );
NAND2_X1 U924 ( .A1(G210), .A2(n1209), .ZN(n1207) );
NAND3_X1 U925 ( .A1(G210), .A2(n1209), .A3(G101), .ZN(n1205) );
NOR2_X1 U926 ( .A1(n988), .A2(n1122), .ZN(n1157) );
NAND3_X1 U927 ( .A1(n1154), .A2(n1172), .A3(n1001), .ZN(n1122) );
INV_X1 U928 ( .A(n1146), .ZN(n1001) );
NAND2_X1 U929 ( .A1(n1003), .A2(n1004), .ZN(n1146) );
NAND2_X1 U930 ( .A1(G214), .A2(n1114), .ZN(n1004) );
XNOR2_X1 U931 ( .A(n1210), .B(n1211), .ZN(n1003) );
NOR2_X1 U932 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
XNOR2_X1 U933 ( .A(KEYINPUT3), .B(n1114), .ZN(n1213) );
OR2_X1 U934 ( .A1(G902), .A2(G237), .ZN(n1114) );
INV_X1 U935 ( .A(G210), .ZN(n1212) );
NAND2_X1 U936 ( .A1(n1214), .A2(n1112), .ZN(n1210) );
XNOR2_X1 U937 ( .A(n1215), .B(n1216), .ZN(n1112) );
XOR2_X1 U938 ( .A(n1217), .B(n1218), .Z(n1216) );
NOR2_X1 U939 ( .A1(n1219), .A2(n1220), .ZN(n1217) );
XNOR2_X1 U940 ( .A(KEYINPUT47), .B(n1008), .ZN(n1220) );
INV_X1 U941 ( .A(G224), .ZN(n1219) );
XOR2_X1 U942 ( .A(n1221), .B(n1073), .Z(n1215) );
XNOR2_X1 U943 ( .A(n1222), .B(n1223), .ZN(n1073) );
XNOR2_X1 U944 ( .A(G116), .B(G119), .ZN(n1222) );
XOR2_X1 U945 ( .A(n1224), .B(n1225), .Z(n1221) );
XOR2_X1 U946 ( .A(G125), .B(n1226), .Z(n1225) );
XNOR2_X1 U947 ( .A(KEYINPUT17), .B(n1199), .ZN(n1226) );
INV_X1 U948 ( .A(G146), .ZN(n1199) );
XOR2_X1 U949 ( .A(n1227), .B(n1075), .Z(n1224) );
XNOR2_X1 U950 ( .A(n1228), .B(n1229), .ZN(n1075) );
XOR2_X1 U951 ( .A(KEYINPUT7), .B(n1230), .Z(n1229) );
NOR2_X1 U952 ( .A1(KEYINPUT38), .A2(n1231), .ZN(n1230) );
NAND2_X1 U953 ( .A1(KEYINPUT51), .A2(n1232), .ZN(n1228) );
INV_X1 U954 ( .A(G104), .ZN(n1232) );
XNOR2_X1 U955 ( .A(n1233), .B(n1234), .ZN(n1227) );
XNOR2_X1 U956 ( .A(n1178), .B(KEYINPUT29), .ZN(n1214) );
NAND2_X1 U957 ( .A1(n983), .A2(n1235), .ZN(n1172) );
NAND4_X1 U958 ( .A1(n1055), .A2(G902), .A3(n1160), .A4(n1067), .ZN(n1235) );
INV_X1 U959 ( .A(G898), .ZN(n1067) );
XNOR2_X1 U960 ( .A(G953), .B(KEYINPUT63), .ZN(n1055) );
NAND3_X1 U961 ( .A1(n1160), .A2(n1008), .A3(G952), .ZN(n983) );
NAND2_X1 U962 ( .A1(G237), .A2(G234), .ZN(n1160) );
INV_X1 U963 ( .A(n993), .ZN(n1154) );
NAND2_X1 U964 ( .A1(n996), .A2(n997), .ZN(n993) );
NAND2_X1 U965 ( .A1(G221), .A2(n1176), .ZN(n997) );
NAND2_X1 U966 ( .A1(G234), .A2(n1140), .ZN(n1176) );
INV_X1 U967 ( .A(G902), .ZN(n1140) );
NAND2_X1 U968 ( .A1(n1236), .A2(n1016), .ZN(n996) );
NAND2_X1 U969 ( .A1(G469), .A2(n1237), .ZN(n1016) );
XOR2_X1 U970 ( .A(n1015), .B(KEYINPUT45), .Z(n1236) );
OR2_X1 U971 ( .A1(n1237), .A2(G469), .ZN(n1015) );
NAND2_X1 U972 ( .A1(n1102), .A2(n1178), .ZN(n1237) );
XNOR2_X1 U973 ( .A(n1238), .B(n1239), .ZN(n1102) );
XOR2_X1 U974 ( .A(n1204), .B(n1240), .Z(n1239) );
XNOR2_X1 U975 ( .A(n1241), .B(n1231), .ZN(n1240) );
XOR2_X1 U976 ( .A(n1208), .B(KEYINPUT49), .Z(n1231) );
INV_X1 U977 ( .A(G101), .ZN(n1208) );
NAND2_X1 U978 ( .A1(n1242), .A2(n1243), .ZN(n1241) );
NAND2_X1 U979 ( .A1(n1244), .A2(n970), .ZN(n1243) );
XNOR2_X1 U980 ( .A(G104), .B(KEYINPUT59), .ZN(n1244) );
NAND2_X1 U981 ( .A1(G107), .A2(n1245), .ZN(n1242) );
XNOR2_X1 U982 ( .A(G104), .B(KEYINPUT41), .ZN(n1245) );
NAND2_X1 U983 ( .A1(n1246), .A2(n1247), .ZN(n1204) );
NAND2_X1 U984 ( .A1(n1248), .A2(n1053), .ZN(n1247) );
XOR2_X1 U985 ( .A(KEYINPUT32), .B(n1051), .Z(n1248) );
NAND2_X1 U986 ( .A1(G134), .A2(n1249), .ZN(n1246) );
XNOR2_X1 U987 ( .A(n1051), .B(KEYINPUT48), .ZN(n1249) );
XNOR2_X1 U988 ( .A(n1250), .B(n1218), .ZN(n1051) );
XNOR2_X1 U989 ( .A(G131), .B(G137), .ZN(n1250) );
XOR2_X1 U990 ( .A(n1251), .B(n1252), .Z(n1238) );
XNOR2_X1 U991 ( .A(KEYINPUT16), .B(n1234), .ZN(n1252) );
INV_X1 U992 ( .A(G110), .ZN(n1234) );
XOR2_X1 U993 ( .A(n1253), .B(n1254), .Z(n1251) );
NAND2_X1 U994 ( .A1(G227), .A2(n1008), .ZN(n1253) );
NAND2_X1 U995 ( .A1(n1255), .A2(n1147), .ZN(n988) );
XOR2_X1 U996 ( .A(n1036), .B(n1038), .Z(n1147) );
INV_X1 U997 ( .A(n1037), .ZN(n1038) );
XOR2_X1 U998 ( .A(G478), .B(KEYINPUT0), .Z(n1037) );
NAND2_X1 U999 ( .A1(n1083), .A2(n1178), .ZN(n1036) );
XNOR2_X1 U1000 ( .A(n1256), .B(n1257), .ZN(n1083) );
XOR2_X1 U1001 ( .A(n1258), .B(n1259), .Z(n1257) );
XNOR2_X1 U1002 ( .A(n1053), .B(G116), .ZN(n1259) );
INV_X1 U1003 ( .A(G134), .ZN(n1053) );
XOR2_X1 U1004 ( .A(KEYINPUT62), .B(KEYINPUT30), .Z(n1258) );
XOR2_X1 U1005 ( .A(n1233), .B(n1260), .Z(n1256) );
XNOR2_X1 U1006 ( .A(n1261), .B(n1218), .ZN(n1260) );
XOR2_X1 U1007 ( .A(G128), .B(G143), .Z(n1218) );
NAND2_X1 U1008 ( .A1(G217), .A2(n1262), .ZN(n1261) );
INV_X1 U1009 ( .A(n1182), .ZN(n1262) );
NAND2_X1 U1010 ( .A1(G234), .A2(n1008), .ZN(n1182) );
INV_X1 U1011 ( .A(G953), .ZN(n1008) );
XNOR2_X1 U1012 ( .A(n970), .B(n1069), .ZN(n1233) );
INV_X1 U1013 ( .A(G107), .ZN(n970) );
XNOR2_X1 U1014 ( .A(KEYINPUT5), .B(n1023), .ZN(n1255) );
XNOR2_X1 U1015 ( .A(n1263), .B(n1089), .ZN(n1023) );
INV_X1 U1016 ( .A(G475), .ZN(n1089) );
NAND2_X1 U1017 ( .A1(n1087), .A2(n1178), .ZN(n1263) );
XOR2_X1 U1018 ( .A(G902), .B(KEYINPUT37), .Z(n1178) );
XNOR2_X1 U1019 ( .A(n1264), .B(n1265), .ZN(n1087) );
XOR2_X1 U1020 ( .A(n1266), .B(n1267), .Z(n1265) );
XNOR2_X1 U1021 ( .A(G104), .B(n1268), .ZN(n1267) );
NOR2_X1 U1022 ( .A1(KEYINPUT31), .A2(G131), .ZN(n1268) );
XNOR2_X1 U1023 ( .A(G143), .B(KEYINPUT14), .ZN(n1266) );
XOR2_X1 U1024 ( .A(n1269), .B(n1270), .Z(n1264) );
XOR2_X1 U1025 ( .A(n1271), .B(n1272), .Z(n1270) );
NOR2_X1 U1026 ( .A1(KEYINPUT15), .A2(n1069), .ZN(n1272) );
XNOR2_X1 U1027 ( .A(G122), .B(KEYINPUT18), .ZN(n1069) );
AND2_X1 U1028 ( .A1(n1209), .A2(G214), .ZN(n1271) );
NOR2_X1 U1029 ( .A1(G953), .A2(G237), .ZN(n1209) );
XOR2_X1 U1030 ( .A(n1050), .B(n1223), .Z(n1269) );
XOR2_X1 U1031 ( .A(G113), .B(KEYINPUT27), .Z(n1223) );
XNOR2_X1 U1032 ( .A(G125), .B(n1254), .ZN(n1050) );
XOR2_X1 U1033 ( .A(G140), .B(G146), .Z(n1254) );
endmodule


