//Key = 1111100001010000111111010100101110000100010000011001100010000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362;

XOR2_X1 U733 ( .A(G107), .B(n1025), .Z(G9) );
NOR2_X1 U734 ( .A1(KEYINPUT22), .A2(n1026), .ZN(n1025) );
NOR2_X1 U735 ( .A1(n1027), .A2(n1028), .ZN(G75) );
NOR4_X1 U736 ( .A1(n1029), .A2(n1030), .A3(G953), .A4(n1031), .ZN(n1028) );
NOR2_X1 U737 ( .A1(n1032), .A2(n1033), .ZN(n1030) );
NOR2_X1 U738 ( .A1(n1034), .A2(n1035), .ZN(n1032) );
XOR2_X1 U739 ( .A(KEYINPUT26), .B(n1036), .Z(n1035) );
NOR4_X1 U740 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1036) );
XOR2_X1 U741 ( .A(KEYINPUT23), .B(n1041), .Z(n1040) );
NOR3_X1 U742 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n1034) );
NOR3_X1 U743 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n1044) );
NOR2_X1 U744 ( .A1(KEYINPUT44), .A2(n1048), .ZN(n1047) );
NOR2_X1 U745 ( .A1(n1049), .A2(n1037), .ZN(n1046) );
NOR2_X1 U746 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
NOR2_X1 U747 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
NOR2_X1 U748 ( .A1(n1041), .A2(n1054), .ZN(n1043) );
NOR2_X1 U749 ( .A1(n1048), .A2(n1055), .ZN(n1054) );
INV_X1 U750 ( .A(KEYINPUT44), .ZN(n1055) );
NAND3_X1 U751 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1029) );
NAND2_X1 U752 ( .A1(n1059), .A2(n1060), .ZN(n1057) );
NAND2_X1 U753 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
NAND4_X1 U754 ( .A1(n1041), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1062) );
NAND3_X1 U755 ( .A1(n1066), .A2(n1067), .A3(n1068), .ZN(n1061) );
NAND2_X1 U756 ( .A1(n1069), .A2(n1045), .ZN(n1067) );
NAND3_X1 U757 ( .A1(n1063), .A2(n1070), .A3(KEYINPUT24), .ZN(n1069) );
NAND3_X1 U758 ( .A1(n1071), .A2(n1072), .A3(n1041), .ZN(n1066) );
INV_X1 U759 ( .A(n1045), .ZN(n1041) );
NAND3_X1 U760 ( .A1(n1070), .A2(n1073), .A3(n1063), .ZN(n1072) );
INV_X1 U761 ( .A(KEYINPUT24), .ZN(n1073) );
NAND2_X1 U762 ( .A1(n1065), .A2(n1074), .ZN(n1071) );
NAND2_X1 U763 ( .A1(n1075), .A2(n1076), .ZN(n1074) );
OR2_X1 U764 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
NOR3_X1 U765 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1027) );
AND4_X1 U766 ( .A1(n1079), .A2(n1080), .A3(n1081), .A4(n1082), .ZN(n1031) );
NOR3_X1 U767 ( .A1(n1083), .A2(n1084), .A3(n1085), .ZN(n1082) );
INV_X1 U768 ( .A(n1078), .ZN(n1084) );
NAND3_X1 U769 ( .A1(n1053), .A2(n1086), .A3(n1087), .ZN(n1083) );
NOR3_X1 U770 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1081) );
XOR2_X1 U771 ( .A(n1091), .B(G472), .Z(n1090) );
NAND2_X1 U772 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
XNOR2_X1 U773 ( .A(KEYINPUT57), .B(KEYINPUT53), .ZN(n1092) );
INV_X1 U774 ( .A(n1094), .ZN(n1089) );
XNOR2_X1 U775 ( .A(n1095), .B(n1096), .ZN(n1088) );
NAND2_X1 U776 ( .A1(KEYINPUT19), .A2(n1097), .ZN(n1095) );
INV_X1 U777 ( .A(G475), .ZN(n1097) );
XNOR2_X1 U778 ( .A(n1098), .B(n1099), .ZN(n1079) );
XOR2_X1 U779 ( .A(n1100), .B(KEYINPUT11), .Z(n1098) );
XOR2_X1 U780 ( .A(n1101), .B(n1102), .Z(G72) );
XOR2_X1 U781 ( .A(n1103), .B(n1104), .Z(n1102) );
NOR2_X1 U782 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U783 ( .A(n1107), .B(n1108), .ZN(n1106) );
XOR2_X1 U784 ( .A(n1109), .B(KEYINPUT8), .Z(n1108) );
NAND2_X1 U785 ( .A1(n1110), .A2(n1111), .ZN(n1103) );
XNOR2_X1 U786 ( .A(n1056), .B(KEYINPUT59), .ZN(n1110) );
NAND2_X1 U787 ( .A1(G953), .A2(n1112), .ZN(n1101) );
NAND2_X1 U788 ( .A1(G900), .A2(G227), .ZN(n1112) );
NAND2_X1 U789 ( .A1(n1113), .A2(n1114), .ZN(G69) );
NAND2_X1 U790 ( .A1(n1115), .A2(n1111), .ZN(n1114) );
XOR2_X1 U791 ( .A(n1116), .B(n1058), .Z(n1115) );
NAND2_X1 U792 ( .A1(n1117), .A2(G953), .ZN(n1113) );
NAND2_X1 U793 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U794 ( .A1(n1116), .A2(n1120), .ZN(n1119) );
NAND2_X1 U795 ( .A1(G224), .A2(n1121), .ZN(n1118) );
NAND2_X1 U796 ( .A1(G898), .A2(n1116), .ZN(n1121) );
NAND3_X1 U797 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1116) );
OR2_X1 U798 ( .A1(n1111), .A2(G898), .ZN(n1124) );
NAND2_X1 U799 ( .A1(KEYINPUT39), .A2(n1125), .ZN(n1123) );
NAND2_X1 U800 ( .A1(n1126), .A2(n1127), .ZN(n1125) );
NAND2_X1 U801 ( .A1(n1128), .A2(n1129), .ZN(n1122) );
INV_X1 U802 ( .A(KEYINPUT39), .ZN(n1129) );
NOR2_X1 U803 ( .A1(n1130), .A2(n1131), .ZN(G66) );
XOR2_X1 U804 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND3_X1 U805 ( .A1(G217), .A2(n1134), .A3(n1135), .ZN(n1132) );
NOR2_X1 U806 ( .A1(n1130), .A2(n1136), .ZN(G63) );
NOR2_X1 U807 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
XOR2_X1 U808 ( .A(n1139), .B(n1140), .Z(n1138) );
NAND2_X1 U809 ( .A1(KEYINPUT3), .A2(n1141), .ZN(n1140) );
NAND2_X1 U810 ( .A1(n1135), .A2(G478), .ZN(n1139) );
NOR2_X1 U811 ( .A1(KEYINPUT3), .A2(n1141), .ZN(n1137) );
NOR2_X1 U812 ( .A1(n1130), .A2(n1142), .ZN(G60) );
XOR2_X1 U813 ( .A(n1143), .B(n1144), .Z(n1142) );
NAND2_X1 U814 ( .A1(n1135), .A2(G475), .ZN(n1143) );
NAND2_X1 U815 ( .A1(n1145), .A2(n1146), .ZN(G6) );
OR2_X1 U816 ( .A1(n1147), .A2(G104), .ZN(n1146) );
XOR2_X1 U817 ( .A(n1148), .B(KEYINPUT29), .Z(n1145) );
NAND2_X1 U818 ( .A1(G104), .A2(n1147), .ZN(n1148) );
NOR3_X1 U819 ( .A1(n1130), .A2(n1149), .A3(n1150), .ZN(G57) );
AND3_X1 U820 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1150) );
NOR2_X1 U821 ( .A1(n1151), .A2(n1154), .ZN(n1149) );
XOR2_X1 U822 ( .A(n1155), .B(n1156), .Z(n1154) );
XNOR2_X1 U823 ( .A(n1157), .B(G101), .ZN(n1151) );
NAND2_X1 U824 ( .A1(n1135), .A2(G472), .ZN(n1157) );
NOR2_X1 U825 ( .A1(n1130), .A2(n1158), .ZN(G54) );
XOR2_X1 U826 ( .A(n1159), .B(n1160), .Z(n1158) );
XOR2_X1 U827 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U828 ( .A(n1163), .B(n1164), .Z(n1159) );
NOR2_X1 U829 ( .A1(KEYINPUT55), .A2(n1165), .ZN(n1164) );
XOR2_X1 U830 ( .A(n1166), .B(n1167), .Z(n1163) );
NOR2_X1 U831 ( .A1(KEYINPUT63), .A2(n1168), .ZN(n1167) );
XOR2_X1 U832 ( .A(n1169), .B(n1170), .Z(n1168) );
XOR2_X1 U833 ( .A(n1171), .B(KEYINPUT35), .Z(n1170) );
NAND2_X1 U834 ( .A1(n1135), .A2(G469), .ZN(n1166) );
NOR2_X1 U835 ( .A1(n1130), .A2(n1172), .ZN(G51) );
XOR2_X1 U836 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U837 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U838 ( .A1(n1177), .A2(n1178), .ZN(n1176) );
NAND2_X1 U839 ( .A1(n1179), .A2(n1180), .ZN(n1178) );
XOR2_X1 U840 ( .A(KEYINPUT60), .B(G125), .Z(n1180) );
XOR2_X1 U841 ( .A(n1171), .B(KEYINPUT34), .Z(n1179) );
XOR2_X1 U842 ( .A(n1181), .B(KEYINPUT15), .Z(n1177) );
NAND2_X1 U843 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
NAND2_X1 U844 ( .A1(n1184), .A2(n1135), .ZN(n1175) );
AND2_X1 U845 ( .A1(n1185), .A2(n1186), .ZN(n1135) );
NAND2_X1 U846 ( .A1(n1187), .A2(n1058), .ZN(n1186) );
AND2_X1 U847 ( .A1(n1188), .A2(n1189), .ZN(n1058) );
NOR4_X1 U848 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
INV_X1 U849 ( .A(n1026), .ZN(n1193) );
NAND3_X1 U850 ( .A1(n1064), .A2(n1065), .A3(n1194), .ZN(n1026) );
AND4_X1 U851 ( .A1(n1195), .A2(n1196), .A3(n1147), .A4(n1197), .ZN(n1188) );
OR2_X1 U852 ( .A1(n1075), .A2(n1198), .ZN(n1197) );
NAND3_X1 U853 ( .A1(n1194), .A2(n1065), .A3(n1199), .ZN(n1147) );
XNOR2_X1 U854 ( .A(n1056), .B(KEYINPUT30), .ZN(n1187) );
AND4_X1 U855 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1056) );
NOR4_X1 U856 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
INV_X1 U857 ( .A(n1208), .ZN(n1207) );
INV_X1 U858 ( .A(n1209), .ZN(n1206) );
NAND2_X1 U859 ( .A1(n1210), .A2(n1211), .ZN(n1202) );
NAND2_X1 U860 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND3_X1 U861 ( .A1(n1214), .A2(n1215), .A3(n1199), .ZN(n1213) );
NAND2_X1 U862 ( .A1(n1216), .A2(n1217), .ZN(n1214) );
NAND3_X1 U863 ( .A1(n1051), .A2(n1218), .A3(n1219), .ZN(n1217) );
INV_X1 U864 ( .A(KEYINPUT6), .ZN(n1218) );
NAND2_X1 U865 ( .A1(n1059), .A2(n1070), .ZN(n1216) );
NAND2_X1 U866 ( .A1(KEYINPUT6), .A2(n1220), .ZN(n1212) );
NAND2_X1 U867 ( .A1(n1221), .A2(n1215), .ZN(n1220) );
XOR2_X1 U868 ( .A(n1222), .B(KEYINPUT2), .Z(n1185) );
XOR2_X1 U869 ( .A(n1223), .B(KEYINPUT0), .Z(n1184) );
NOR2_X1 U870 ( .A1(n1111), .A2(G952), .ZN(n1130) );
NAND2_X1 U871 ( .A1(n1224), .A2(n1225), .ZN(G48) );
NAND2_X1 U872 ( .A1(G146), .A2(n1226), .ZN(n1225) );
XOR2_X1 U873 ( .A(n1227), .B(KEYINPUT36), .Z(n1224) );
OR2_X1 U874 ( .A1(n1226), .A2(G146), .ZN(n1227) );
NAND3_X1 U875 ( .A1(n1221), .A2(n1210), .A3(n1228), .ZN(n1226) );
XOR2_X1 U876 ( .A(n1215), .B(KEYINPUT27), .Z(n1228) );
AND3_X1 U877 ( .A1(n1199), .A2(n1051), .A3(n1219), .ZN(n1221) );
XNOR2_X1 U878 ( .A(G143), .B(n1200), .ZN(G45) );
NAND4_X1 U879 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1200) );
NAND2_X1 U880 ( .A1(n1233), .A2(n1234), .ZN(G42) );
NAND2_X1 U881 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
NAND2_X1 U882 ( .A1(n1237), .A2(n1238), .ZN(n1235) );
NAND2_X1 U883 ( .A1(n1201), .A2(n1239), .ZN(n1238) );
OR2_X1 U884 ( .A1(n1239), .A2(n1240), .ZN(n1237) );
INV_X1 U885 ( .A(KEYINPUT32), .ZN(n1239) );
NAND2_X1 U886 ( .A1(G140), .A2(n1240), .ZN(n1233) );
NOR2_X1 U887 ( .A1(n1241), .A2(KEYINPUT38), .ZN(n1240) );
INV_X1 U888 ( .A(n1201), .ZN(n1241) );
NAND2_X1 U889 ( .A1(n1242), .A2(n1243), .ZN(n1201) );
NAND2_X1 U890 ( .A1(n1244), .A2(n1245), .ZN(G39) );
OR2_X1 U891 ( .A1(n1208), .A2(G137), .ZN(n1245) );
XOR2_X1 U892 ( .A(n1246), .B(KEYINPUT33), .Z(n1244) );
NAND2_X1 U893 ( .A1(G137), .A2(n1208), .ZN(n1246) );
NAND3_X1 U894 ( .A1(n1219), .A2(n1068), .A3(n1243), .ZN(n1208) );
XOR2_X1 U895 ( .A(n1247), .B(n1248), .Z(G36) );
XOR2_X1 U896 ( .A(KEYINPUT21), .B(G134), .Z(n1248) );
NAND2_X1 U897 ( .A1(KEYINPUT28), .A2(n1205), .ZN(n1247) );
AND3_X1 U898 ( .A1(n1230), .A2(n1064), .A3(n1243), .ZN(n1205) );
XOR2_X1 U899 ( .A(G131), .B(n1204), .Z(G33) );
AND3_X1 U900 ( .A1(n1230), .A2(n1199), .A3(n1243), .ZN(n1204) );
AND3_X1 U901 ( .A1(n1051), .A2(n1215), .A3(n1063), .ZN(n1243) );
INV_X1 U902 ( .A(n1033), .ZN(n1063) );
NAND2_X1 U903 ( .A1(n1249), .A2(n1250), .ZN(n1033) );
XNOR2_X1 U904 ( .A(KEYINPUT13), .B(n1077), .ZN(n1250) );
XOR2_X1 U905 ( .A(G128), .B(n1251), .Z(G30) );
NOR2_X1 U906 ( .A1(KEYINPUT54), .A2(n1209), .ZN(n1251) );
NAND3_X1 U907 ( .A1(n1219), .A2(n1064), .A3(n1229), .ZN(n1209) );
AND3_X1 U908 ( .A1(n1210), .A2(n1215), .A3(n1051), .ZN(n1229) );
NAND2_X1 U909 ( .A1(n1252), .A2(n1253), .ZN(G3) );
NAND2_X1 U910 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
NAND2_X1 U911 ( .A1(G101), .A2(n1256), .ZN(n1252) );
NAND2_X1 U912 ( .A1(n1257), .A2(n1258), .ZN(n1256) );
NAND2_X1 U913 ( .A1(KEYINPUT5), .A2(n1259), .ZN(n1258) );
INV_X1 U914 ( .A(n1196), .ZN(n1259) );
OR2_X1 U915 ( .A1(n1254), .A2(KEYINPUT5), .ZN(n1257) );
NOR2_X1 U916 ( .A1(KEYINPUT10), .A2(n1196), .ZN(n1254) );
NAND3_X1 U917 ( .A1(n1068), .A2(n1194), .A3(n1230), .ZN(n1196) );
XOR2_X1 U918 ( .A(n1183), .B(n1260), .Z(G27) );
NAND4_X1 U919 ( .A1(n1261), .A2(n1242), .A3(n1059), .A4(n1215), .ZN(n1260) );
NAND2_X1 U920 ( .A1(n1045), .A2(n1262), .ZN(n1215) );
NAND3_X1 U921 ( .A1(n1105), .A2(n1263), .A3(n1264), .ZN(n1262) );
XOR2_X1 U922 ( .A(n1222), .B(KEYINPUT4), .Z(n1264) );
NOR2_X1 U923 ( .A1(n1111), .A2(G900), .ZN(n1105) );
AND2_X1 U924 ( .A1(n1199), .A2(n1070), .ZN(n1242) );
XOR2_X1 U925 ( .A(n1075), .B(KEYINPUT1), .Z(n1261) );
XNOR2_X1 U926 ( .A(G122), .B(n1265), .ZN(G24) );
NAND2_X1 U927 ( .A1(KEYINPUT16), .A2(n1192), .ZN(n1265) );
AND4_X1 U928 ( .A1(n1266), .A2(n1232), .A3(n1231), .A4(n1267), .ZN(n1192) );
NOR2_X1 U929 ( .A1(n1042), .A2(n1038), .ZN(n1267) );
INV_X1 U930 ( .A(n1065), .ZN(n1042) );
NOR2_X1 U931 ( .A1(n1268), .A2(n1269), .ZN(n1065) );
XOR2_X1 U932 ( .A(G119), .B(n1270), .Z(G21) );
NOR2_X1 U933 ( .A1(KEYINPUT50), .A2(n1195), .ZN(n1270) );
NAND4_X1 U934 ( .A1(n1219), .A2(n1059), .A3(n1068), .A4(n1266), .ZN(n1195) );
AND2_X1 U935 ( .A1(n1269), .A2(n1268), .ZN(n1219) );
INV_X1 U936 ( .A(n1271), .ZN(n1269) );
NAND2_X1 U937 ( .A1(n1272), .A2(n1273), .ZN(G18) );
NAND2_X1 U938 ( .A1(G116), .A2(n1274), .ZN(n1273) );
XOR2_X1 U939 ( .A(n1275), .B(KEYINPUT45), .Z(n1272) );
OR2_X1 U940 ( .A1(n1274), .A2(G116), .ZN(n1275) );
NAND2_X1 U941 ( .A1(n1276), .A2(n1210), .ZN(n1274) );
XOR2_X1 U942 ( .A(n1198), .B(KEYINPUT37), .Z(n1276) );
NAND4_X1 U943 ( .A1(n1230), .A2(n1059), .A3(n1064), .A4(n1277), .ZN(n1198) );
AND2_X1 U944 ( .A1(n1278), .A2(n1231), .ZN(n1064) );
XOR2_X1 U945 ( .A(n1080), .B(KEYINPUT48), .Z(n1231) );
XOR2_X1 U946 ( .A(G113), .B(n1191), .Z(G15) );
NOR3_X1 U947 ( .A1(n1048), .A2(n1279), .A3(n1039), .ZN(n1191) );
INV_X1 U948 ( .A(n1230), .ZN(n1039) );
NOR2_X1 U949 ( .A1(n1268), .A2(n1271), .ZN(n1230) );
NAND2_X1 U950 ( .A1(n1199), .A2(n1059), .ZN(n1048) );
INV_X1 U951 ( .A(n1038), .ZN(n1059) );
NAND2_X1 U952 ( .A1(n1280), .A2(n1053), .ZN(n1038) );
INV_X1 U953 ( .A(n1052), .ZN(n1280) );
AND2_X1 U954 ( .A1(n1080), .A2(n1232), .ZN(n1199) );
INV_X1 U955 ( .A(n1278), .ZN(n1232) );
XOR2_X1 U956 ( .A(n1190), .B(n1281), .Z(G12) );
NOR2_X1 U957 ( .A1(KEYINPUT12), .A2(n1282), .ZN(n1281) );
INV_X1 U958 ( .A(G110), .ZN(n1282) );
AND3_X1 U959 ( .A1(n1068), .A2(n1194), .A3(n1070), .ZN(n1190) );
AND2_X1 U960 ( .A1(n1271), .A2(n1268), .ZN(n1070) );
NAND2_X1 U961 ( .A1(n1283), .A2(n1094), .ZN(n1268) );
NAND3_X1 U962 ( .A1(n1284), .A2(n1222), .A3(n1133), .ZN(n1094) );
NAND2_X1 U963 ( .A1(G217), .A2(n1285), .ZN(n1284) );
INV_X1 U964 ( .A(G234), .ZN(n1285) );
XOR2_X1 U965 ( .A(KEYINPUT51), .B(n1085), .Z(n1283) );
AND3_X1 U966 ( .A1(n1286), .A2(n1134), .A3(G217), .ZN(n1085) );
NAND2_X1 U967 ( .A1(n1133), .A2(n1222), .ZN(n1286) );
XNOR2_X1 U968 ( .A(n1287), .B(n1288), .ZN(n1133) );
XOR2_X1 U969 ( .A(n1289), .B(n1290), .Z(n1288) );
NOR2_X1 U970 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
XOR2_X1 U971 ( .A(KEYINPUT49), .B(n1293), .Z(n1292) );
NOR2_X1 U972 ( .A1(G146), .A2(n1107), .ZN(n1293) );
AND2_X1 U973 ( .A1(n1107), .A2(G146), .ZN(n1291) );
XNOR2_X1 U974 ( .A(n1183), .B(G140), .ZN(n1107) );
AND3_X1 U975 ( .A1(G221), .A2(n1111), .A3(G234), .ZN(n1289) );
XOR2_X1 U976 ( .A(n1294), .B(G137), .Z(n1287) );
NAND2_X1 U977 ( .A1(n1295), .A2(n1296), .ZN(n1294) );
NAND2_X1 U978 ( .A1(G110), .A2(n1297), .ZN(n1296) );
XOR2_X1 U979 ( .A(KEYINPUT9), .B(n1298), .Z(n1295) );
NOR2_X1 U980 ( .A1(G110), .A2(n1297), .ZN(n1298) );
XOR2_X1 U981 ( .A(G128), .B(G119), .Z(n1297) );
XOR2_X1 U982 ( .A(n1093), .B(G472), .Z(n1271) );
NAND3_X1 U983 ( .A1(n1299), .A2(n1222), .A3(n1300), .ZN(n1093) );
NAND3_X1 U984 ( .A1(n1301), .A2(n1255), .A3(KEYINPUT18), .ZN(n1300) );
NAND3_X1 U985 ( .A1(n1302), .A2(n1303), .A3(n1152), .ZN(n1301) );
OR2_X1 U986 ( .A1(n1153), .A2(KEYINPUT43), .ZN(n1303) );
NAND2_X1 U987 ( .A1(KEYINPUT43), .A2(n1156), .ZN(n1302) );
NAND4_X1 U988 ( .A1(n1304), .A2(n1153), .A3(n1305), .A4(n1306), .ZN(n1299) );
OR2_X1 U989 ( .A1(n1152), .A2(KEYINPUT43), .ZN(n1306) );
NAND2_X1 U990 ( .A1(n1156), .A2(n1155), .ZN(n1152) );
NAND2_X1 U991 ( .A1(KEYINPUT43), .A2(n1307), .ZN(n1305) );
OR2_X1 U992 ( .A1(n1155), .A2(n1156), .ZN(n1153) );
INV_X1 U993 ( .A(n1307), .ZN(n1156) );
XOR2_X1 U994 ( .A(n1308), .B(n1309), .Z(n1307) );
INV_X1 U995 ( .A(n1109), .ZN(n1309) );
NAND3_X1 U996 ( .A1(n1310), .A2(n1111), .A3(G210), .ZN(n1155) );
NAND2_X1 U997 ( .A1(KEYINPUT18), .A2(n1255), .ZN(n1304) );
AND2_X1 U998 ( .A1(n1051), .A2(n1266), .ZN(n1194) );
INV_X1 U999 ( .A(n1279), .ZN(n1266) );
NAND2_X1 U1000 ( .A1(n1210), .A2(n1277), .ZN(n1279) );
NAND2_X1 U1001 ( .A1(n1311), .A2(n1045), .ZN(n1277) );
NAND3_X1 U1002 ( .A1(n1263), .A2(n1111), .A3(n1312), .ZN(n1045) );
XNOR2_X1 U1003 ( .A(G952), .B(KEYINPUT17), .ZN(n1312) );
XOR2_X1 U1004 ( .A(KEYINPUT25), .B(n1313), .Z(n1311) );
NOR4_X1 U1005 ( .A1(G898), .A2(n1314), .A3(n1222), .A4(n1111), .ZN(n1313) );
INV_X1 U1006 ( .A(n1263), .ZN(n1314) );
NAND2_X1 U1007 ( .A1(G237), .A2(G234), .ZN(n1263) );
INV_X1 U1008 ( .A(n1075), .ZN(n1210) );
NAND2_X1 U1009 ( .A1(n1249), .A2(n1077), .ZN(n1075) );
NAND3_X1 U1010 ( .A1(n1315), .A2(n1316), .A3(n1317), .ZN(n1077) );
XNOR2_X1 U1011 ( .A(KEYINPUT56), .B(n1087), .ZN(n1317) );
NAND2_X1 U1012 ( .A1(n1318), .A2(n1319), .ZN(n1087) );
OR2_X1 U1013 ( .A1(n1086), .A2(KEYINPUT62), .ZN(n1316) );
NAND2_X1 U1014 ( .A1(n1320), .A2(n1223), .ZN(n1086) );
NAND3_X1 U1015 ( .A1(n1320), .A2(n1318), .A3(KEYINPUT62), .ZN(n1315) );
INV_X1 U1016 ( .A(n1223), .ZN(n1318) );
NAND2_X1 U1017 ( .A1(G210), .A2(n1321), .ZN(n1223) );
INV_X1 U1018 ( .A(n1319), .ZN(n1320) );
NAND2_X1 U1019 ( .A1(n1322), .A2(n1222), .ZN(n1319) );
XOR2_X1 U1020 ( .A(n1323), .B(n1324), .Z(n1322) );
XOR2_X1 U1021 ( .A(KEYINPUT31), .B(G125), .Z(n1324) );
XOR2_X1 U1022 ( .A(n1173), .B(n1171), .Z(n1323) );
XOR2_X1 U1023 ( .A(n1128), .B(n1325), .Z(n1173) );
NOR2_X1 U1024 ( .A1(G953), .A2(n1120), .ZN(n1325) );
INV_X1 U1025 ( .A(G224), .ZN(n1120) );
XNOR2_X1 U1026 ( .A(n1126), .B(n1127), .ZN(n1128) );
XOR2_X1 U1027 ( .A(G110), .B(G122), .Z(n1127) );
XOR2_X1 U1028 ( .A(n1169), .B(n1308), .Z(n1126) );
XOR2_X1 U1029 ( .A(G113), .B(n1326), .Z(n1308) );
XOR2_X1 U1030 ( .A(G119), .B(G116), .Z(n1326) );
XOR2_X1 U1031 ( .A(n1078), .B(KEYINPUT14), .Z(n1249) );
NAND2_X1 U1032 ( .A1(G214), .A2(n1321), .ZN(n1078) );
NAND2_X1 U1033 ( .A1(n1222), .A2(n1310), .ZN(n1321) );
INV_X1 U1034 ( .A(G237), .ZN(n1310) );
AND2_X1 U1035 ( .A1(n1052), .A2(n1053), .ZN(n1051) );
NAND2_X1 U1036 ( .A1(G221), .A2(n1134), .ZN(n1053) );
NAND2_X1 U1037 ( .A1(G234), .A2(n1222), .ZN(n1134) );
XOR2_X1 U1038 ( .A(n1100), .B(n1327), .Z(n1052) );
NOR2_X1 U1039 ( .A1(KEYINPUT42), .A2(n1099), .ZN(n1327) );
XNOR2_X1 U1040 ( .A(G469), .B(KEYINPUT52), .ZN(n1099) );
NAND2_X1 U1041 ( .A1(n1328), .A2(n1222), .ZN(n1100) );
XOR2_X1 U1042 ( .A(n1329), .B(n1330), .Z(n1328) );
XOR2_X1 U1043 ( .A(n1331), .B(n1162), .Z(n1330) );
XOR2_X1 U1044 ( .A(G110), .B(G140), .Z(n1162) );
INV_X1 U1045 ( .A(n1169), .ZN(n1331) );
XOR2_X1 U1046 ( .A(n1255), .B(n1332), .Z(n1169) );
XOR2_X1 U1047 ( .A(G107), .B(G104), .Z(n1332) );
INV_X1 U1048 ( .A(G101), .ZN(n1255) );
XOR2_X1 U1049 ( .A(n1109), .B(n1333), .Z(n1329) );
XNOR2_X1 U1050 ( .A(KEYINPUT20), .B(n1165), .ZN(n1333) );
NAND2_X1 U1051 ( .A1(G227), .A2(n1111), .ZN(n1165) );
XOR2_X1 U1052 ( .A(n1161), .B(n1182), .Z(n1109) );
INV_X1 U1053 ( .A(n1171), .ZN(n1182) );
XOR2_X1 U1054 ( .A(n1334), .B(n1335), .Z(n1171) );
INV_X1 U1055 ( .A(G128), .ZN(n1334) );
XOR2_X1 U1056 ( .A(n1336), .B(n1337), .Z(n1161) );
XOR2_X1 U1057 ( .A(G137), .B(G134), .Z(n1337) );
INV_X1 U1058 ( .A(G131), .ZN(n1336) );
INV_X1 U1059 ( .A(n1037), .ZN(n1068) );
NAND2_X1 U1060 ( .A1(n1278), .A2(n1080), .ZN(n1037) );
XOR2_X1 U1061 ( .A(n1338), .B(G478), .Z(n1080) );
NAND2_X1 U1062 ( .A1(n1222), .A2(n1141), .ZN(n1338) );
NAND2_X1 U1063 ( .A1(n1339), .A2(n1340), .ZN(n1141) );
NAND2_X1 U1064 ( .A1(n1341), .A2(n1342), .ZN(n1340) );
XOR2_X1 U1065 ( .A(n1343), .B(KEYINPUT58), .Z(n1339) );
OR2_X1 U1066 ( .A1(n1342), .A2(n1341), .ZN(n1343) );
AND3_X1 U1067 ( .A1(G234), .A2(n1111), .A3(G217), .ZN(n1341) );
INV_X1 U1068 ( .A(G953), .ZN(n1111) );
XNOR2_X1 U1069 ( .A(n1344), .B(n1345), .ZN(n1342) );
XOR2_X1 U1070 ( .A(n1346), .B(n1347), .Z(n1345) );
XOR2_X1 U1071 ( .A(G134), .B(G128), .Z(n1347) );
XOR2_X1 U1072 ( .A(KEYINPUT41), .B(G143), .Z(n1346) );
XNOR2_X1 U1073 ( .A(G107), .B(n1348), .ZN(n1344) );
XOR2_X1 U1074 ( .A(G122), .B(G116), .Z(n1348) );
XOR2_X1 U1075 ( .A(n1096), .B(G475), .Z(n1278) );
NAND2_X1 U1076 ( .A1(n1144), .A2(n1222), .ZN(n1096) );
INV_X1 U1077 ( .A(G902), .ZN(n1222) );
XOR2_X1 U1078 ( .A(n1349), .B(n1350), .Z(n1144) );
XOR2_X1 U1079 ( .A(n1351), .B(n1352), .Z(n1350) );
XOR2_X1 U1080 ( .A(G104), .B(n1353), .Z(n1352) );
NOR4_X1 U1081 ( .A1(KEYINPUT46), .A2(G953), .A3(G237), .A4(n1354), .ZN(n1353) );
INV_X1 U1082 ( .A(G214), .ZN(n1354) );
XOR2_X1 U1083 ( .A(G131), .B(G122), .Z(n1351) );
XOR2_X1 U1084 ( .A(n1355), .B(n1356), .Z(n1349) );
XOR2_X1 U1085 ( .A(n1357), .B(n1335), .Z(n1356) );
XOR2_X1 U1086 ( .A(G143), .B(G146), .Z(n1335) );
NOR2_X1 U1087 ( .A1(G113), .A2(KEYINPUT7), .ZN(n1357) );
NAND2_X1 U1088 ( .A1(n1358), .A2(n1359), .ZN(n1355) );
NAND2_X1 U1089 ( .A1(n1360), .A2(n1183), .ZN(n1359) );
INV_X1 U1090 ( .A(G125), .ZN(n1183) );
XOR2_X1 U1091 ( .A(n1236), .B(n1361), .Z(n1360) );
XNOR2_X1 U1092 ( .A(KEYINPUT47), .B(KEYINPUT40), .ZN(n1361) );
NAND2_X1 U1093 ( .A1(G125), .A2(n1362), .ZN(n1358) );
XOR2_X1 U1094 ( .A(n1236), .B(KEYINPUT61), .Z(n1362) );
INV_X1 U1095 ( .A(G140), .ZN(n1236) );
endmodule


