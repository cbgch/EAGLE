//Key = 0011110011000101011010001010001011110110010111000001000010111011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;

XNOR2_X1 U746 ( .A(G107), .B(n1029), .ZN(G9) );
NOR2_X1 U747 ( .A1(n1030), .A2(n1031), .ZN(G75) );
NOR4_X1 U748 ( .A1(n1032), .A2(n1033), .A3(n1034), .A4(n1035), .ZN(n1031) );
XOR2_X1 U749 ( .A(n1036), .B(KEYINPUT52), .Z(n1034) );
NAND3_X1 U750 ( .A1(n1037), .A2(n1038), .A3(n1039), .ZN(n1032) );
NAND2_X1 U751 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
NAND2_X1 U752 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
NAND3_X1 U753 ( .A1(n1044), .A2(n1045), .A3(n1046), .ZN(n1043) );
NAND2_X1 U754 ( .A1(n1047), .A2(n1048), .ZN(n1045) );
NAND2_X1 U755 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NAND2_X1 U756 ( .A1(n1051), .A2(n1052), .ZN(n1050) );
NAND2_X1 U757 ( .A1(n1053), .A2(n1054), .ZN(n1052) );
INV_X1 U758 ( .A(n1055), .ZN(n1051) );
NAND3_X1 U759 ( .A1(n1056), .A2(n1057), .A3(n1054), .ZN(n1042) );
NAND2_X1 U760 ( .A1(n1058), .A2(n1059), .ZN(n1056) );
NAND3_X1 U761 ( .A1(n1044), .A2(n1060), .A3(n1046), .ZN(n1059) );
NAND2_X1 U762 ( .A1(n1049), .A2(n1061), .ZN(n1058) );
NAND3_X1 U763 ( .A1(n1062), .A2(n1063), .A3(n1064), .ZN(n1061) );
NAND2_X1 U764 ( .A1(n1046), .A2(n1065), .ZN(n1064) );
NAND2_X1 U765 ( .A1(n1044), .A2(n1066), .ZN(n1062) );
NAND2_X1 U766 ( .A1(n1067), .A2(n1068), .ZN(n1066) );
NAND2_X1 U767 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
INV_X1 U768 ( .A(n1071), .ZN(n1040) );
NOR3_X1 U769 ( .A1(n1072), .A2(G953), .A3(G952), .ZN(n1030) );
INV_X1 U770 ( .A(n1037), .ZN(n1072) );
NAND4_X1 U771 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1037) );
NOR4_X1 U772 ( .A1(n1077), .A2(n1078), .A3(n1079), .A4(n1080), .ZN(n1076) );
XNOR2_X1 U773 ( .A(G469), .B(n1081), .ZN(n1080) );
XOR2_X1 U774 ( .A(G478), .B(n1082), .Z(n1079) );
XOR2_X1 U775 ( .A(KEYINPUT57), .B(n1083), .Z(n1078) );
XOR2_X1 U776 ( .A(KEYINPUT60), .B(n1084), .Z(n1077) );
NOR2_X1 U777 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
NOR2_X1 U778 ( .A1(n1087), .A2(n1088), .ZN(n1085) );
XOR2_X1 U779 ( .A(n1089), .B(KEYINPUT15), .Z(n1087) );
NOR3_X1 U780 ( .A1(n1053), .A2(n1069), .A3(n1090), .ZN(n1075) );
NAND2_X1 U781 ( .A1(G475), .A2(n1091), .ZN(n1074) );
XOR2_X1 U782 ( .A(n1092), .B(n1093), .Z(n1073) );
XNOR2_X1 U783 ( .A(G472), .B(KEYINPUT44), .ZN(n1093) );
XOR2_X1 U784 ( .A(n1094), .B(n1095), .Z(G72) );
NOR2_X1 U785 ( .A1(n1096), .A2(n1038), .ZN(n1095) );
NOR2_X1 U786 ( .A1(n1097), .A2(n1098), .ZN(n1096) );
NAND2_X1 U787 ( .A1(n1099), .A2(n1100), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1101), .A2(n1038), .ZN(n1100) );
XOR2_X1 U789 ( .A(n1102), .B(n1036), .Z(n1101) );
NAND3_X1 U790 ( .A1(G900), .A2(n1102), .A3(G953), .ZN(n1099) );
XOR2_X1 U791 ( .A(n1103), .B(n1104), .Z(n1102) );
XOR2_X1 U792 ( .A(n1105), .B(n1106), .Z(n1104) );
NOR2_X1 U793 ( .A1(KEYINPUT11), .A2(n1107), .ZN(n1105) );
XOR2_X1 U794 ( .A(G128), .B(n1108), .Z(n1107) );
NAND2_X1 U795 ( .A1(n1109), .A2(n1110), .ZN(G69) );
NAND3_X1 U796 ( .A1(n1111), .A2(n1112), .A3(KEYINPUT2), .ZN(n1110) );
OR2_X1 U797 ( .A1(n1038), .A2(G224), .ZN(n1112) );
XNOR2_X1 U798 ( .A(n1113), .B(n1114), .ZN(n1111) );
NAND2_X1 U799 ( .A1(n1115), .A2(n1116), .ZN(n1109) );
NAND2_X1 U800 ( .A1(KEYINPUT2), .A2(n1117), .ZN(n1116) );
NAND2_X1 U801 ( .A1(G953), .A2(n1118), .ZN(n1117) );
NAND2_X1 U802 ( .A1(G898), .A2(G224), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1114), .B(n1113), .Z(n1115) );
AND2_X1 U804 ( .A1(n1119), .A2(n1038), .ZN(n1113) );
NAND3_X1 U805 ( .A1(n1120), .A2(n1121), .A3(n1122), .ZN(n1119) );
XOR2_X1 U806 ( .A(n1123), .B(KEYINPUT28), .Z(n1122) );
INV_X1 U807 ( .A(n1033), .ZN(n1120) );
NAND2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1114) );
NAND2_X1 U809 ( .A1(G953), .A2(n1126), .ZN(n1125) );
XOR2_X1 U810 ( .A(n1127), .B(n1128), .Z(n1124) );
NOR2_X1 U811 ( .A1(n1129), .A2(n1130), .ZN(G66) );
XNOR2_X1 U812 ( .A(n1131), .B(n1132), .ZN(n1130) );
NOR2_X1 U813 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NOR2_X1 U814 ( .A1(n1135), .A2(n1136), .ZN(G63) );
XOR2_X1 U815 ( .A(n1137), .B(n1138), .Z(n1136) );
NOR2_X1 U816 ( .A1(n1139), .A2(n1134), .ZN(n1137) );
NOR2_X1 U817 ( .A1(n1140), .A2(n1038), .ZN(n1135) );
XNOR2_X1 U818 ( .A(G952), .B(KEYINPUT58), .ZN(n1140) );
NOR2_X1 U819 ( .A1(n1129), .A2(n1141), .ZN(G60) );
XOR2_X1 U820 ( .A(n1142), .B(n1143), .Z(n1141) );
NOR2_X1 U821 ( .A1(n1134), .A2(n1144), .ZN(n1142) );
XOR2_X1 U822 ( .A(KEYINPUT43), .B(G475), .Z(n1144) );
XNOR2_X1 U823 ( .A(n1145), .B(n1146), .ZN(G6) );
NOR2_X1 U824 ( .A1(KEYINPUT47), .A2(n1147), .ZN(n1146) );
INV_X1 U825 ( .A(G104), .ZN(n1147) );
NOR2_X1 U826 ( .A1(n1129), .A2(n1148), .ZN(G57) );
XOR2_X1 U827 ( .A(n1149), .B(n1150), .Z(n1148) );
XNOR2_X1 U828 ( .A(n1151), .B(n1152), .ZN(n1150) );
XOR2_X1 U829 ( .A(n1153), .B(n1154), .Z(n1149) );
NAND3_X1 U830 ( .A1(n1155), .A2(n1156), .A3(G472), .ZN(n1154) );
NAND2_X1 U831 ( .A1(KEYINPUT8), .A2(n1134), .ZN(n1156) );
NAND2_X1 U832 ( .A1(n1157), .A2(n1158), .ZN(n1155) );
INV_X1 U833 ( .A(KEYINPUT8), .ZN(n1158) );
NAND2_X1 U834 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NOR2_X1 U835 ( .A1(n1129), .A2(n1161), .ZN(G54) );
XOR2_X1 U836 ( .A(n1162), .B(n1163), .Z(n1161) );
XNOR2_X1 U837 ( .A(n1164), .B(n1165), .ZN(n1163) );
XOR2_X1 U838 ( .A(n1166), .B(n1167), .Z(n1162) );
NOR2_X1 U839 ( .A1(n1168), .A2(n1134), .ZN(n1167) );
XNOR2_X1 U840 ( .A(G469), .B(KEYINPUT25), .ZN(n1168) );
NOR2_X1 U841 ( .A1(n1129), .A2(n1169), .ZN(G51) );
XOR2_X1 U842 ( .A(n1170), .B(n1171), .Z(n1169) );
XOR2_X1 U843 ( .A(n1172), .B(n1173), .Z(n1171) );
NOR2_X1 U844 ( .A1(KEYINPUT42), .A2(n1174), .ZN(n1172) );
XOR2_X1 U845 ( .A(G125), .B(n1175), .Z(n1170) );
NOR2_X1 U846 ( .A1(n1088), .A2(n1134), .ZN(n1175) );
NAND2_X1 U847 ( .A1(G902), .A2(n1159), .ZN(n1134) );
OR3_X1 U848 ( .A1(n1035), .A2(n1036), .A3(n1033), .ZN(n1159) );
NAND4_X1 U849 ( .A1(n1145), .A2(n1176), .A3(n1177), .A4(n1029), .ZN(n1033) );
NAND3_X1 U850 ( .A1(n1044), .A2(n1060), .A3(n1178), .ZN(n1029) );
NAND3_X1 U851 ( .A1(n1178), .A2(n1044), .A3(n1179), .ZN(n1145) );
NAND4_X1 U852 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1036) );
NOR4_X1 U853 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1189), .ZN(n1182) );
NAND2_X1 U855 ( .A1(n1190), .A2(n1191), .ZN(n1180) );
XNOR2_X1 U856 ( .A(KEYINPUT16), .B(n1192), .ZN(n1190) );
XNOR2_X1 U857 ( .A(n1193), .B(KEYINPUT20), .ZN(n1035) );
NAND2_X1 U858 ( .A1(n1121), .A2(n1123), .ZN(n1193) );
NAND2_X1 U859 ( .A1(n1194), .A2(n1195), .ZN(n1123) );
XOR2_X1 U860 ( .A(KEYINPUT21), .B(n1196), .Z(n1195) );
AND3_X1 U861 ( .A1(n1197), .A2(n1198), .A3(n1065), .ZN(n1196) );
AND3_X1 U862 ( .A1(n1199), .A2(n1200), .A3(n1201), .ZN(n1121) );
NOR2_X1 U863 ( .A1(n1038), .A2(G952), .ZN(n1129) );
XOR2_X1 U864 ( .A(n1202), .B(n1203), .Z(G48) );
NOR2_X1 U865 ( .A1(n1067), .A2(n1192), .ZN(n1203) );
NAND2_X1 U866 ( .A1(n1204), .A2(n1179), .ZN(n1192) );
NOR2_X1 U867 ( .A1(KEYINPUT49), .A2(n1205), .ZN(n1202) );
XOR2_X1 U868 ( .A(n1206), .B(n1181), .Z(G45) );
NAND4_X1 U869 ( .A1(n1207), .A2(n1208), .A3(n1191), .A4(n1209), .ZN(n1181) );
NAND2_X1 U870 ( .A1(n1210), .A2(n1211), .ZN(G42) );
NAND2_X1 U871 ( .A1(n1185), .A2(n1212), .ZN(n1211) );
XOR2_X1 U872 ( .A(KEYINPUT26), .B(n1213), .Z(n1210) );
NOR2_X1 U873 ( .A1(n1185), .A2(n1212), .ZN(n1213) );
AND4_X1 U874 ( .A1(n1214), .A2(n1179), .A3(n1055), .A4(n1215), .ZN(n1185) );
INV_X1 U875 ( .A(n1063), .ZN(n1214) );
NAND3_X1 U876 ( .A1(n1083), .A2(n1216), .A3(n1046), .ZN(n1063) );
XOR2_X1 U877 ( .A(G137), .B(n1184), .Z(G39) );
AND3_X1 U878 ( .A1(n1046), .A2(n1049), .A3(n1204), .ZN(n1184) );
XOR2_X1 U879 ( .A(G134), .B(n1189), .Z(G36) );
AND3_X1 U880 ( .A1(n1046), .A2(n1060), .A3(n1208), .ZN(n1189) );
XOR2_X1 U881 ( .A(G131), .B(n1188), .Z(G33) );
AND3_X1 U882 ( .A1(n1046), .A2(n1179), .A3(n1208), .ZN(n1188) );
AND3_X1 U883 ( .A1(n1055), .A2(n1215), .A3(n1065), .ZN(n1208) );
NOR2_X1 U884 ( .A1(n1217), .A2(n1069), .ZN(n1046) );
XOR2_X1 U885 ( .A(G128), .B(n1187), .Z(G30) );
AND3_X1 U886 ( .A1(n1191), .A2(n1060), .A3(n1204), .ZN(n1187) );
AND4_X1 U887 ( .A1(n1218), .A2(n1055), .A3(n1083), .A4(n1215), .ZN(n1204) );
XOR2_X1 U888 ( .A(n1153), .B(n1176), .Z(G3) );
NAND3_X1 U889 ( .A1(n1178), .A2(n1049), .A3(n1065), .ZN(n1176) );
XNOR2_X1 U890 ( .A(n1186), .B(n1219), .ZN(G27) );
XOR2_X1 U891 ( .A(KEYINPUT35), .B(G125), .Z(n1219) );
AND4_X1 U892 ( .A1(n1216), .A2(n1215), .A3(n1083), .A4(n1220), .ZN(n1186) );
NOR2_X1 U893 ( .A1(n1067), .A2(n1047), .ZN(n1220) );
NAND2_X1 U894 ( .A1(n1071), .A2(n1221), .ZN(n1215) );
NAND4_X1 U895 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1098), .ZN(n1221) );
INV_X1 U896 ( .A(G900), .ZN(n1098) );
XOR2_X1 U897 ( .A(n1201), .B(n1223), .Z(G24) );
XOR2_X1 U898 ( .A(n1224), .B(KEYINPUT12), .Z(n1223) );
NAND4_X1 U899 ( .A1(n1225), .A2(n1044), .A3(n1207), .A4(n1209), .ZN(n1201) );
NOR2_X1 U900 ( .A1(n1083), .A2(n1218), .ZN(n1044) );
XNOR2_X1 U901 ( .A(G119), .B(n1199), .ZN(G21) );
NAND4_X1 U902 ( .A1(n1218), .A2(n1225), .A3(n1049), .A4(n1083), .ZN(n1199) );
XOR2_X1 U903 ( .A(n1200), .B(n1226), .Z(G18) );
NAND2_X1 U904 ( .A1(KEYINPUT17), .A2(G116), .ZN(n1226) );
NAND3_X1 U905 ( .A1(n1065), .A2(n1060), .A3(n1225), .ZN(n1200) );
AND4_X1 U906 ( .A1(n1191), .A2(n1054), .A3(n1198), .A4(n1057), .ZN(n1225) );
INV_X1 U907 ( .A(n1067), .ZN(n1191) );
XNOR2_X1 U908 ( .A(n1194), .B(KEYINPUT22), .ZN(n1067) );
NAND2_X1 U909 ( .A1(n1227), .A2(n1228), .ZN(n1060) );
NAND3_X1 U910 ( .A1(n1229), .A2(n1207), .A3(n1230), .ZN(n1228) );
INV_X1 U911 ( .A(KEYINPUT23), .ZN(n1230) );
NAND2_X1 U912 ( .A1(KEYINPUT23), .A2(n1049), .ZN(n1227) );
XNOR2_X1 U913 ( .A(G113), .B(n1231), .ZN(G15) );
NAND4_X1 U914 ( .A1(n1197), .A2(n1194), .A3(n1232), .A4(n1198), .ZN(n1231) );
XOR2_X1 U915 ( .A(KEYINPUT61), .B(n1065), .Z(n1232) );
NOR2_X1 U916 ( .A1(n1216), .A2(n1083), .ZN(n1065) );
INV_X1 U917 ( .A(n1047), .ZN(n1197) );
NAND3_X1 U918 ( .A1(n1054), .A2(n1057), .A3(n1179), .ZN(n1047) );
NOR2_X1 U919 ( .A1(n1207), .A2(n1229), .ZN(n1179) );
XOR2_X1 U920 ( .A(n1233), .B(n1177), .Z(G12) );
NAND4_X1 U921 ( .A1(n1178), .A2(n1049), .A3(n1083), .A4(n1216), .ZN(n1177) );
INV_X1 U922 ( .A(n1218), .ZN(n1216) );
XOR2_X1 U923 ( .A(n1092), .B(n1234), .Z(n1218) );
NOR2_X1 U924 ( .A1(G472), .A2(KEYINPUT36), .ZN(n1234) );
NAND2_X1 U925 ( .A1(n1235), .A2(n1236), .ZN(n1092) );
XNOR2_X1 U926 ( .A(n1237), .B(n1152), .ZN(n1235) );
XOR2_X1 U927 ( .A(n1238), .B(n1239), .Z(n1152) );
XOR2_X1 U928 ( .A(n1240), .B(n1241), .Z(n1239) );
XOR2_X1 U929 ( .A(KEYINPUT51), .B(KEYINPUT5), .Z(n1241) );
XOR2_X1 U930 ( .A(n1242), .B(n1243), .Z(n1238) );
INV_X1 U931 ( .A(n1244), .ZN(n1243) );
NAND2_X1 U932 ( .A1(n1245), .A2(KEYINPUT18), .ZN(n1237) );
XOR2_X1 U933 ( .A(n1153), .B(n1246), .Z(n1245) );
NOR2_X1 U934 ( .A1(n1151), .A2(KEYINPUT0), .ZN(n1246) );
AND3_X1 U935 ( .A1(n1247), .A2(n1038), .A3(G210), .ZN(n1151) );
INV_X1 U936 ( .A(G101), .ZN(n1153) );
XOR2_X1 U937 ( .A(n1248), .B(n1133), .Z(n1083) );
NAND2_X1 U938 ( .A1(G217), .A2(n1249), .ZN(n1133) );
NAND2_X1 U939 ( .A1(n1236), .A2(n1131), .ZN(n1248) );
XNOR2_X1 U940 ( .A(n1250), .B(n1251), .ZN(n1131) );
XOR2_X1 U941 ( .A(n1252), .B(n1253), .Z(n1251) );
XOR2_X1 U942 ( .A(G137), .B(G125), .Z(n1253) );
XOR2_X1 U943 ( .A(KEYINPUT41), .B(G146), .Z(n1252) );
XOR2_X1 U944 ( .A(n1254), .B(n1255), .Z(n1250) );
AND2_X1 U945 ( .A1(G221), .A2(n1256), .ZN(n1255) );
XOR2_X1 U946 ( .A(n1257), .B(n1258), .Z(n1254) );
NOR2_X1 U947 ( .A1(G140), .A2(KEYINPUT48), .ZN(n1258) );
NAND2_X1 U948 ( .A1(n1259), .A2(n1260), .ZN(n1257) );
NAND2_X1 U949 ( .A1(n1261), .A2(n1233), .ZN(n1260) );
XOR2_X1 U950 ( .A(KEYINPUT30), .B(n1262), .Z(n1259) );
NOR2_X1 U951 ( .A1(n1233), .A2(n1261), .ZN(n1262) );
NAND2_X1 U952 ( .A1(n1263), .A2(n1264), .ZN(n1261) );
NAND2_X1 U953 ( .A1(n1265), .A2(n1266), .ZN(n1264) );
NAND2_X1 U954 ( .A1(KEYINPUT9), .A2(n1267), .ZN(n1266) );
OR2_X1 U955 ( .A1(G128), .A2(KEYINPUT10), .ZN(n1267) );
NAND2_X1 U956 ( .A1(G128), .A2(n1268), .ZN(n1263) );
NAND2_X1 U957 ( .A1(n1269), .A2(n1270), .ZN(n1268) );
NAND2_X1 U958 ( .A1(KEYINPUT9), .A2(n1271), .ZN(n1270) );
INV_X1 U959 ( .A(KEYINPUT10), .ZN(n1269) );
NOR2_X1 U960 ( .A1(n1209), .A2(n1207), .ZN(n1049) );
XOR2_X1 U961 ( .A(n1272), .B(n1082), .Z(n1207) );
NOR2_X1 U962 ( .A1(n1138), .A2(n1273), .ZN(n1082) );
INV_X1 U963 ( .A(n1236), .ZN(n1273) );
XNOR2_X1 U964 ( .A(n1274), .B(n1275), .ZN(n1138) );
NOR3_X1 U965 ( .A1(n1276), .A2(KEYINPUT14), .A3(n1277), .ZN(n1275) );
NOR2_X1 U966 ( .A1(n1278), .A2(n1279), .ZN(n1277) );
XOR2_X1 U967 ( .A(n1280), .B(n1281), .Z(n1279) );
INV_X1 U968 ( .A(n1282), .ZN(n1278) );
XOR2_X1 U969 ( .A(KEYINPUT39), .B(n1283), .Z(n1276) );
NOR2_X1 U970 ( .A1(n1284), .A2(n1282), .ZN(n1283) );
NAND3_X1 U971 ( .A1(n1285), .A2(n1286), .A3(n1287), .ZN(n1282) );
NAND2_X1 U972 ( .A1(n1288), .A2(n1289), .ZN(n1287) );
NAND2_X1 U973 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
XOR2_X1 U974 ( .A(KEYINPUT59), .B(G134), .Z(n1290) );
XOR2_X1 U975 ( .A(G143), .B(G128), .Z(n1288) );
NAND3_X1 U976 ( .A1(n1292), .A2(n1293), .A3(n1291), .ZN(n1286) );
INV_X1 U977 ( .A(KEYINPUT40), .ZN(n1291) );
INV_X1 U978 ( .A(G134), .ZN(n1293) );
XOR2_X1 U979 ( .A(n1206), .B(G128), .Z(n1292) );
NAND2_X1 U980 ( .A1(G134), .A2(KEYINPUT40), .ZN(n1285) );
XOR2_X1 U981 ( .A(n1294), .B(n1280), .Z(n1284) );
NOR3_X1 U982 ( .A1(n1295), .A2(n1296), .A3(KEYINPUT55), .ZN(n1280) );
NOR3_X1 U983 ( .A1(KEYINPUT13), .A2(G116), .A3(n1224), .ZN(n1296) );
INV_X1 U984 ( .A(G122), .ZN(n1224) );
NOR2_X1 U985 ( .A1(n1297), .A2(n1298), .ZN(n1295) );
INV_X1 U986 ( .A(KEYINPUT13), .ZN(n1298) );
XOR2_X1 U987 ( .A(G122), .B(G116), .Z(n1297) );
NAND2_X1 U988 ( .A1(n1256), .A2(G217), .ZN(n1274) );
AND2_X1 U989 ( .A1(G234), .A2(n1038), .ZN(n1256) );
NAND2_X1 U990 ( .A1(KEYINPUT3), .A2(n1139), .ZN(n1272) );
INV_X1 U991 ( .A(G478), .ZN(n1139) );
INV_X1 U992 ( .A(n1229), .ZN(n1209) );
NOR2_X1 U993 ( .A1(n1299), .A2(n1090), .ZN(n1229) );
NOR2_X1 U994 ( .A1(n1091), .A2(G475), .ZN(n1090) );
AND2_X1 U995 ( .A1(n1300), .A2(n1091), .ZN(n1299) );
NAND2_X1 U996 ( .A1(n1236), .A2(n1301), .ZN(n1091) );
XOR2_X1 U997 ( .A(KEYINPUT37), .B(n1143), .Z(n1301) );
XNOR2_X1 U998 ( .A(n1302), .B(n1303), .ZN(n1143) );
XOR2_X1 U999 ( .A(n1240), .B(n1106), .Z(n1303) );
XOR2_X1 U1000 ( .A(G125), .B(n1304), .Z(n1106) );
XOR2_X1 U1001 ( .A(G140), .B(G131), .Z(n1304) );
XOR2_X1 U1002 ( .A(n1305), .B(n1306), .Z(n1302) );
XOR2_X1 U1003 ( .A(KEYINPUT41), .B(n1307), .Z(n1306) );
AND3_X1 U1004 ( .A1(G214), .A2(n1038), .A3(n1247), .ZN(n1307) );
NAND3_X1 U1005 ( .A1(n1308), .A2(n1309), .A3(n1310), .ZN(n1305) );
OR2_X1 U1006 ( .A1(n1311), .A2(n1312), .ZN(n1310) );
NAND2_X1 U1007 ( .A1(KEYINPUT54), .A2(n1313), .ZN(n1309) );
NAND2_X1 U1008 ( .A1(n1312), .A2(n1314), .ZN(n1313) );
XNOR2_X1 U1009 ( .A(KEYINPUT33), .B(n1311), .ZN(n1314) );
NAND2_X1 U1010 ( .A1(n1315), .A2(n1316), .ZN(n1308) );
INV_X1 U1011 ( .A(KEYINPUT54), .ZN(n1316) );
NAND2_X1 U1012 ( .A1(n1317), .A2(n1318), .ZN(n1315) );
NAND3_X1 U1013 ( .A1(KEYINPUT33), .A2(n1312), .A3(n1311), .ZN(n1318) );
XNOR2_X1 U1014 ( .A(G113), .B(G122), .ZN(n1312) );
OR2_X1 U1015 ( .A1(n1311), .A2(KEYINPUT33), .ZN(n1317) );
XNOR2_X1 U1016 ( .A(G104), .B(KEYINPUT27), .ZN(n1311) );
XNOR2_X1 U1017 ( .A(G475), .B(KEYINPUT45), .ZN(n1300) );
AND3_X1 U1018 ( .A1(n1194), .A2(n1198), .A3(n1055), .ZN(n1178) );
NOR2_X1 U1019 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
INV_X1 U1020 ( .A(n1057), .ZN(n1053) );
NAND2_X1 U1021 ( .A1(G221), .A2(n1249), .ZN(n1057) );
NAND2_X1 U1022 ( .A1(G234), .A2(n1160), .ZN(n1249) );
XNOR2_X1 U1023 ( .A(n1081), .B(n1319), .ZN(n1054) );
NOR2_X1 U1024 ( .A1(G469), .A2(KEYINPUT50), .ZN(n1319) );
NAND2_X1 U1025 ( .A1(n1236), .A2(n1320), .ZN(n1081) );
XOR2_X1 U1026 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1027 ( .A(n1323), .B(n1164), .Z(n1322) );
XOR2_X1 U1028 ( .A(n1324), .B(n1325), .Z(n1164) );
XOR2_X1 U1029 ( .A(n1326), .B(n1327), .Z(n1325) );
XOR2_X1 U1030 ( .A(G104), .B(n1108), .Z(n1327) );
NOR2_X1 U1031 ( .A1(KEYINPUT1), .A2(n1328), .ZN(n1108) );
XOR2_X1 U1032 ( .A(n1205), .B(n1329), .Z(n1328) );
NAND2_X1 U1033 ( .A1(KEYINPUT24), .A2(n1206), .ZN(n1329) );
INV_X1 U1034 ( .A(G143), .ZN(n1206) );
INV_X1 U1035 ( .A(G146), .ZN(n1205) );
NOR2_X1 U1036 ( .A1(G101), .A2(KEYINPUT6), .ZN(n1326) );
XOR2_X1 U1037 ( .A(n1242), .B(n1281), .Z(n1324) );
INV_X1 U1038 ( .A(n1294), .ZN(n1281) );
XOR2_X1 U1039 ( .A(n1330), .B(n1103), .Z(n1242) );
XNOR2_X1 U1040 ( .A(n1331), .B(G134), .ZN(n1103) );
INV_X1 U1041 ( .A(G137), .ZN(n1331) );
XOR2_X1 U1042 ( .A(n1332), .B(G128), .Z(n1330) );
NAND2_X1 U1043 ( .A1(KEYINPUT38), .A2(n1333), .ZN(n1332) );
INV_X1 U1044 ( .A(G131), .ZN(n1333) );
NAND2_X1 U1045 ( .A1(KEYINPUT4), .A2(n1165), .ZN(n1323) );
XOR2_X1 U1046 ( .A(n1212), .B(n1233), .Z(n1165) );
INV_X1 U1047 ( .A(G140), .ZN(n1212) );
XOR2_X1 U1048 ( .A(KEYINPUT32), .B(n1166), .Z(n1321) );
NOR2_X1 U1049 ( .A1(n1097), .A2(G953), .ZN(n1166) );
INV_X1 U1050 ( .A(G227), .ZN(n1097) );
NAND2_X1 U1051 ( .A1(n1071), .A2(n1334), .ZN(n1198) );
NAND4_X1 U1052 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1126), .ZN(n1334) );
INV_X1 U1053 ( .A(G898), .ZN(n1126) );
NAND3_X1 U1054 ( .A1(n1222), .A2(n1038), .A3(G952), .ZN(n1071) );
NAND2_X1 U1055 ( .A1(G237), .A2(G234), .ZN(n1222) );
NOR2_X1 U1056 ( .A1(n1070), .A2(n1069), .ZN(n1194) );
AND2_X1 U1057 ( .A1(G214), .A2(n1335), .ZN(n1069) );
INV_X1 U1058 ( .A(n1217), .ZN(n1070) );
NAND2_X1 U1059 ( .A1(n1336), .A2(n1337), .ZN(n1217) );
NAND2_X1 U1060 ( .A1(n1338), .A2(n1089), .ZN(n1337) );
XNOR2_X1 U1061 ( .A(n1086), .B(KEYINPUT19), .ZN(n1336) );
NOR2_X1 U1062 ( .A1(n1089), .A2(n1338), .ZN(n1086) );
INV_X1 U1063 ( .A(n1088), .ZN(n1338) );
NAND2_X1 U1064 ( .A1(G210), .A2(n1335), .ZN(n1088) );
NAND2_X1 U1065 ( .A1(n1160), .A2(n1247), .ZN(n1335) );
INV_X1 U1066 ( .A(G237), .ZN(n1247) );
NAND2_X1 U1067 ( .A1(n1339), .A2(n1236), .ZN(n1089) );
XOR2_X1 U1068 ( .A(n1160), .B(KEYINPUT53), .Z(n1236) );
INV_X1 U1069 ( .A(G902), .ZN(n1160) );
XOR2_X1 U1070 ( .A(n1173), .B(n1340), .Z(n1339) );
XOR2_X1 U1071 ( .A(G125), .B(n1174), .Z(n1340) );
XOR2_X1 U1072 ( .A(G128), .B(n1240), .Z(n1174) );
XOR2_X1 U1073 ( .A(G143), .B(G146), .Z(n1240) );
XNOR2_X1 U1074 ( .A(n1341), .B(n1342), .ZN(n1173) );
XOR2_X1 U1075 ( .A(n1343), .B(n1344), .Z(n1342) );
NAND2_X1 U1076 ( .A1(KEYINPUT34), .A2(n1128), .ZN(n1344) );
AND2_X1 U1077 ( .A1(n1345), .A2(n1346), .ZN(n1128) );
NAND2_X1 U1078 ( .A1(n1347), .A2(n1233), .ZN(n1346) );
XOR2_X1 U1079 ( .A(KEYINPUT7), .B(G122), .Z(n1347) );
XOR2_X1 U1080 ( .A(KEYINPUT63), .B(n1348), .Z(n1345) );
NOR2_X1 U1081 ( .A1(G122), .A2(n1233), .ZN(n1348) );
NAND2_X1 U1082 ( .A1(G224), .A2(n1038), .ZN(n1343) );
INV_X1 U1083 ( .A(G953), .ZN(n1038) );
NAND2_X1 U1084 ( .A1(n1349), .A2(n1350), .ZN(n1341) );
NAND2_X1 U1085 ( .A1(n1127), .A2(n1351), .ZN(n1350) );
XOR2_X1 U1086 ( .A(n1352), .B(n1353), .Z(n1127) );
OR3_X1 U1087 ( .A1(n1352), .A2(n1353), .A3(n1351), .ZN(n1349) );
INV_X1 U1088 ( .A(KEYINPUT29), .ZN(n1351) );
XNOR2_X1 U1089 ( .A(n1244), .B(KEYINPUT56), .ZN(n1353) );
XOR2_X1 U1090 ( .A(n1354), .B(n1271), .Z(n1244) );
INV_X1 U1091 ( .A(n1265), .ZN(n1271) );
XNOR2_X1 U1092 ( .A(G119), .B(KEYINPUT31), .ZN(n1265) );
XNOR2_X1 U1093 ( .A(G113), .B(G116), .ZN(n1354) );
XOR2_X1 U1094 ( .A(n1294), .B(n1355), .Z(n1352) );
XOR2_X1 U1095 ( .A(G101), .B(n1356), .Z(n1355) );
NOR2_X1 U1096 ( .A1(G104), .A2(KEYINPUT46), .ZN(n1356) );
XNOR2_X1 U1097 ( .A(G107), .B(KEYINPUT62), .ZN(n1294) );
INV_X1 U1098 ( .A(G110), .ZN(n1233) );
endmodule


