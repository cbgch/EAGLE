//Key = 0000000100100010010101000001110010010011100111101010010101010111


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
n1355, n1356;

XNOR2_X1 U742 ( .A(G107), .B(n1025), .ZN(G9) );
NOR2_X1 U743 ( .A1(n1026), .A2(n1027), .ZN(G75) );
NOR4_X1 U744 ( .A1(G953), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1027) );
NOR2_X1 U745 ( .A1(n1031), .A2(n1032), .ZN(n1029) );
NOR2_X1 U746 ( .A1(n1033), .A2(n1034), .ZN(n1031) );
NOR3_X1 U747 ( .A1(n1035), .A2(n1036), .A3(n1037), .ZN(n1034) );
NOR3_X1 U748 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1036) );
NOR3_X1 U749 ( .A1(n1041), .A2(KEYINPUT53), .A3(n1042), .ZN(n1040) );
INV_X1 U750 ( .A(n1043), .ZN(n1042) );
NOR2_X1 U751 ( .A1(n1044), .A2(n1045), .ZN(n1039) );
NOR3_X1 U752 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1044) );
NOR2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR2_X1 U754 ( .A1(n1051), .A2(n1052), .ZN(n1049) );
NOR3_X1 U755 ( .A1(n1053), .A2(n1054), .A3(n1055), .ZN(n1051) );
NOR3_X1 U756 ( .A1(n1056), .A2(n1057), .A3(n1058), .ZN(n1047) );
AND2_X1 U757 ( .A1(n1043), .A2(KEYINPUT53), .ZN(n1046) );
NOR3_X1 U758 ( .A1(n1050), .A2(n1059), .A3(n1057), .ZN(n1038) );
NOR2_X1 U759 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
NOR2_X1 U760 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NOR4_X1 U761 ( .A1(n1064), .A2(n1045), .A3(n1057), .A4(n1050), .ZN(n1033) );
INV_X1 U762 ( .A(n1041), .ZN(n1045) );
NOR2_X1 U763 ( .A1(n1065), .A2(n1066), .ZN(n1064) );
NOR3_X1 U764 ( .A1(n1028), .A2(G953), .A3(G952), .ZN(n1026) );
AND4_X1 U765 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1028) );
NOR4_X1 U766 ( .A1(n1071), .A2(n1072), .A3(n1057), .A4(n1035), .ZN(n1070) );
XNOR2_X1 U767 ( .A(n1073), .B(n1074), .ZN(n1069) );
XOR2_X1 U768 ( .A(n1075), .B(KEYINPUT0), .Z(n1068) );
XOR2_X1 U769 ( .A(n1076), .B(n1077), .Z(n1067) );
NOR2_X1 U770 ( .A1(KEYINPUT5), .A2(n1078), .ZN(n1077) );
XOR2_X1 U771 ( .A(n1079), .B(n1080), .Z(G72) );
XOR2_X1 U772 ( .A(n1081), .B(n1082), .Z(n1080) );
NOR2_X1 U773 ( .A1(n1083), .A2(n1084), .ZN(n1082) );
NOR2_X1 U774 ( .A1(n1085), .A2(n1086), .ZN(n1083) );
NAND2_X1 U775 ( .A1(n1087), .A2(n1088), .ZN(n1081) );
NAND2_X1 U776 ( .A1(n1089), .A2(n1086), .ZN(n1088) );
XOR2_X1 U777 ( .A(n1090), .B(n1091), .Z(n1087) );
XNOR2_X1 U778 ( .A(n1092), .B(n1093), .ZN(n1091) );
NAND3_X1 U779 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1092) );
OR2_X1 U780 ( .A1(n1097), .A2(KEYINPUT7), .ZN(n1096) );
NAND3_X1 U781 ( .A1(KEYINPUT7), .A2(n1098), .A3(n1099), .ZN(n1095) );
OR2_X1 U782 ( .A1(n1099), .A2(n1098), .ZN(n1094) );
NOR2_X1 U783 ( .A1(G125), .A2(KEYINPUT8), .ZN(n1098) );
XOR2_X1 U784 ( .A(n1100), .B(n1101), .Z(n1090) );
XNOR2_X1 U785 ( .A(KEYINPUT21), .B(n1102), .ZN(n1101) );
NOR2_X1 U786 ( .A1(n1103), .A2(n1104), .ZN(n1100) );
XOR2_X1 U787 ( .A(n1105), .B(KEYINPUT61), .Z(n1104) );
NAND4_X1 U788 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1105) );
OR2_X1 U789 ( .A1(G134), .A2(KEYINPUT57), .ZN(n1109) );
NAND3_X1 U790 ( .A1(G134), .A2(n1110), .A3(KEYINPUT57), .ZN(n1108) );
NOR2_X1 U791 ( .A1(n1111), .A2(n1107), .ZN(n1103) );
INV_X1 U792 ( .A(G131), .ZN(n1107) );
NOR2_X1 U793 ( .A1(n1112), .A2(n1113), .ZN(n1111) );
NOR2_X1 U794 ( .A1(G137), .A2(n1114), .ZN(n1113) );
XNOR2_X1 U795 ( .A(KEYINPUT57), .B(n1115), .ZN(n1114) );
NAND2_X1 U796 ( .A1(n1084), .A2(n1116), .ZN(n1079) );
NAND2_X1 U797 ( .A1(n1117), .A2(n1118), .ZN(G69) );
NAND2_X1 U798 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
NAND2_X1 U799 ( .A1(n1121), .A2(n1122), .ZN(n1117) );
INV_X1 U800 ( .A(n1120), .ZN(n1122) );
NAND2_X1 U801 ( .A1(G953), .A2(n1123), .ZN(n1120) );
NAND2_X1 U802 ( .A1(G898), .A2(G224), .ZN(n1123) );
XNOR2_X1 U803 ( .A(n1119), .B(n1124), .ZN(n1121) );
XNOR2_X1 U804 ( .A(KEYINPUT51), .B(KEYINPUT39), .ZN(n1124) );
XNOR2_X1 U805 ( .A(n1125), .B(n1126), .ZN(n1119) );
NOR2_X1 U806 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
XOR2_X1 U807 ( .A(n1129), .B(n1130), .Z(n1128) );
XOR2_X1 U808 ( .A(n1131), .B(n1132), .Z(n1130) );
XNOR2_X1 U809 ( .A(G107), .B(KEYINPUT11), .ZN(n1129) );
AND2_X1 U810 ( .A1(n1133), .A2(n1089), .ZN(n1127) );
NAND2_X1 U811 ( .A1(n1084), .A2(n1134), .ZN(n1125) );
NOR2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(G66) );
XNOR2_X1 U813 ( .A(n1137), .B(n1138), .ZN(n1136) );
NOR2_X1 U814 ( .A1(n1074), .A2(n1139), .ZN(n1138) );
NOR2_X1 U815 ( .A1(n1135), .A2(n1140), .ZN(G63) );
XOR2_X1 U816 ( .A(n1141), .B(n1142), .Z(n1140) );
AND2_X1 U817 ( .A1(G478), .A2(n1143), .ZN(n1141) );
NOR3_X1 U818 ( .A1(n1144), .A2(n1145), .A3(n1146), .ZN(G60) );
NOR3_X1 U819 ( .A1(n1147), .A2(G953), .A3(G952), .ZN(n1146) );
AND2_X1 U820 ( .A1(n1147), .A2(n1135), .ZN(n1145) );
INV_X1 U821 ( .A(KEYINPUT49), .ZN(n1147) );
XOR2_X1 U822 ( .A(n1148), .B(n1149), .Z(n1144) );
AND2_X1 U823 ( .A1(G475), .A2(n1143), .ZN(n1148) );
XNOR2_X1 U824 ( .A(G104), .B(n1150), .ZN(G6) );
NOR2_X1 U825 ( .A1(n1151), .A2(n1152), .ZN(G57) );
XOR2_X1 U826 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND3_X1 U827 ( .A1(n1143), .A2(G472), .A3(KEYINPUT59), .ZN(n1153) );
NOR2_X1 U828 ( .A1(n1155), .A2(n1084), .ZN(n1151) );
XNOR2_X1 U829 ( .A(G952), .B(KEYINPUT48), .ZN(n1155) );
NOR2_X1 U830 ( .A1(n1135), .A2(n1156), .ZN(G54) );
XOR2_X1 U831 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U832 ( .A(n1159), .B(n1160), .Z(n1158) );
AND2_X1 U833 ( .A1(G469), .A2(n1143), .ZN(n1159) );
INV_X1 U834 ( .A(n1139), .ZN(n1143) );
XOR2_X1 U835 ( .A(KEYINPUT27), .B(n1161), .Z(n1157) );
NOR2_X1 U836 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
XOR2_X1 U837 ( .A(n1164), .B(KEYINPUT40), .Z(n1163) );
NOR2_X1 U838 ( .A1(n1084), .A2(G952), .ZN(n1135) );
NOR2_X1 U839 ( .A1(n1165), .A2(n1166), .ZN(G51) );
XOR2_X1 U840 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U841 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U842 ( .A1(KEYINPUT25), .A2(n1171), .ZN(n1170) );
NOR2_X1 U843 ( .A1(n1172), .A2(n1139), .ZN(n1169) );
NAND2_X1 U844 ( .A1(G902), .A2(n1030), .ZN(n1139) );
OR2_X1 U845 ( .A1(n1134), .A2(n1116), .ZN(n1030) );
NAND4_X1 U846 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1116) );
AND3_X1 U847 ( .A1(n1177), .A2(n1178), .A3(n1179), .ZN(n1176) );
NAND3_X1 U848 ( .A1(n1180), .A2(n1181), .A3(n1066), .ZN(n1175) );
NAND2_X1 U849 ( .A1(n1062), .A2(n1182), .ZN(n1181) );
NAND2_X1 U850 ( .A1(n1183), .A2(n1184), .ZN(n1182) );
NAND3_X1 U851 ( .A1(n1185), .A2(n1186), .A3(n1187), .ZN(n1180) );
NAND3_X1 U852 ( .A1(n1188), .A2(n1189), .A3(n1043), .ZN(n1186) );
NAND2_X1 U853 ( .A1(n1183), .A2(n1190), .ZN(n1185) );
XNOR2_X1 U854 ( .A(KEYINPUT36), .B(n1050), .ZN(n1190) );
INV_X1 U855 ( .A(n1191), .ZN(n1050) );
NAND4_X1 U856 ( .A1(n1192), .A2(n1150), .A3(n1193), .A4(n1194), .ZN(n1134) );
NOR4_X1 U857 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1194) );
NOR2_X1 U858 ( .A1(KEYINPUT58), .A2(n1199), .ZN(n1198) );
NOR2_X1 U859 ( .A1(KEYINPUT3), .A2(n1200), .ZN(n1197) );
NOR3_X1 U860 ( .A1(n1201), .A2(n1188), .A3(n1202), .ZN(n1196) );
NOR3_X1 U861 ( .A1(n1203), .A2(n1204), .A3(n1205), .ZN(n1195) );
XNOR2_X1 U862 ( .A(KEYINPUT18), .B(n1206), .ZN(n1203) );
AND3_X1 U863 ( .A1(n1207), .A2(n1025), .A3(n1208), .ZN(n1193) );
NAND3_X1 U864 ( .A1(n1209), .A2(n1065), .A3(n1041), .ZN(n1025) );
NAND3_X1 U865 ( .A1(n1041), .A2(n1209), .A3(n1066), .ZN(n1150) );
NAND4_X1 U866 ( .A1(n1210), .A2(n1211), .A3(n1206), .A4(n1212), .ZN(n1192) );
NAND2_X1 U867 ( .A1(n1213), .A2(n1214), .ZN(n1211) );
NAND3_X1 U868 ( .A1(n1066), .A2(n1061), .A3(KEYINPUT58), .ZN(n1214) );
NAND3_X1 U869 ( .A1(n1188), .A2(n1215), .A3(KEYINPUT3), .ZN(n1213) );
XOR2_X1 U870 ( .A(n1216), .B(KEYINPUT20), .Z(n1172) );
NOR2_X1 U871 ( .A1(G952), .A2(n1217), .ZN(n1165) );
XNOR2_X1 U872 ( .A(G953), .B(KEYINPUT52), .ZN(n1217) );
XNOR2_X1 U873 ( .A(G146), .B(n1218), .ZN(G48) );
NAND4_X1 U874 ( .A1(KEYINPUT38), .A2(n1183), .A3(n1219), .A4(n1066), .ZN(n1218) );
NOR2_X1 U875 ( .A1(n1212), .A2(n1187), .ZN(n1219) );
XNOR2_X1 U876 ( .A(G143), .B(n1174), .ZN(G45) );
NAND4_X1 U877 ( .A1(n1220), .A2(n1184), .A3(n1035), .A4(n1221), .ZN(n1174) );
XNOR2_X1 U878 ( .A(G140), .B(n1222), .ZN(G42) );
NAND4_X1 U879 ( .A1(n1191), .A2(n1183), .A3(n1066), .A4(n1187), .ZN(n1222) );
NAND2_X1 U880 ( .A1(n1223), .A2(n1224), .ZN(G39) );
NAND2_X1 U881 ( .A1(G137), .A2(n1173), .ZN(n1224) );
XOR2_X1 U882 ( .A(KEYINPUT10), .B(n1225), .Z(n1223) );
NOR2_X1 U883 ( .A1(G137), .A2(n1173), .ZN(n1225) );
NAND3_X1 U884 ( .A1(n1183), .A2(n1215), .A3(n1191), .ZN(n1173) );
XOR2_X1 U885 ( .A(n1177), .B(n1226), .Z(G36) );
NOR2_X1 U886 ( .A1(G134), .A2(KEYINPUT41), .ZN(n1226) );
NAND3_X1 U887 ( .A1(n1220), .A2(n1065), .A3(n1191), .ZN(n1177) );
XNOR2_X1 U888 ( .A(G131), .B(n1179), .ZN(G33) );
NAND3_X1 U889 ( .A1(n1220), .A2(n1066), .A3(n1191), .ZN(n1179) );
NOR2_X1 U890 ( .A1(n1058), .A2(n1071), .ZN(n1191) );
AND3_X1 U891 ( .A1(n1052), .A2(n1189), .A3(n1061), .ZN(n1220) );
XNOR2_X1 U892 ( .A(G128), .B(n1178), .ZN(G30) );
NAND4_X1 U893 ( .A1(n1062), .A2(n1183), .A3(n1065), .A4(n1184), .ZN(n1178) );
AND3_X1 U894 ( .A1(n1052), .A2(n1189), .A3(n1188), .ZN(n1183) );
XOR2_X1 U895 ( .A(G101), .B(n1227), .Z(G3) );
NOR4_X1 U896 ( .A1(KEYINPUT31), .A2(n1188), .A3(n1202), .A4(n1201), .ZN(n1227) );
INV_X1 U897 ( .A(n1215), .ZN(n1201) );
XNOR2_X1 U898 ( .A(G125), .B(n1228), .ZN(G27) );
NAND4_X1 U899 ( .A1(n1188), .A2(n1043), .A3(n1066), .A4(n1229), .ZN(n1228) );
NOR3_X1 U900 ( .A1(n1062), .A2(KEYINPUT34), .A3(n1230), .ZN(n1229) );
INV_X1 U901 ( .A(n1189), .ZN(n1230) );
NAND2_X1 U902 ( .A1(n1032), .A2(n1231), .ZN(n1189) );
NAND2_X1 U903 ( .A1(n1232), .A2(n1086), .ZN(n1231) );
INV_X1 U904 ( .A(G900), .ZN(n1086) );
NAND2_X1 U905 ( .A1(n1233), .A2(n1234), .ZN(G24) );
NAND2_X1 U906 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
XOR2_X1 U907 ( .A(KEYINPUT14), .B(n1237), .Z(n1233) );
NOR2_X1 U908 ( .A1(n1236), .A2(n1235), .ZN(n1237) );
XNOR2_X1 U909 ( .A(KEYINPUT9), .B(G122), .ZN(n1235) );
NOR3_X1 U910 ( .A1(n1205), .A2(n1204), .A3(n1238), .ZN(n1236) );
XNOR2_X1 U911 ( .A(n1206), .B(KEYINPUT12), .ZN(n1238) );
NAND3_X1 U912 ( .A1(n1041), .A2(n1035), .A3(n1043), .ZN(n1205) );
NOR2_X1 U913 ( .A1(n1062), .A2(n1188), .ZN(n1041) );
XOR2_X1 U914 ( .A(n1200), .B(n1239), .Z(G21) );
NAND2_X1 U915 ( .A1(KEYINPUT44), .A2(G119), .ZN(n1239) );
NAND4_X1 U916 ( .A1(n1215), .A2(n1043), .A3(n1188), .A4(n1206), .ZN(n1200) );
NOR3_X1 U917 ( .A1(n1035), .A2(n1037), .A3(n1187), .ZN(n1215) );
XNOR2_X1 U918 ( .A(n1240), .B(n1241), .ZN(G18) );
NOR2_X1 U919 ( .A1(KEYINPUT1), .A2(n1207), .ZN(n1241) );
NAND2_X1 U920 ( .A1(n1242), .A2(n1065), .ZN(n1207) );
NOR2_X1 U921 ( .A1(n1035), .A2(n1204), .ZN(n1065) );
INV_X1 U922 ( .A(n1221), .ZN(n1204) );
XOR2_X1 U923 ( .A(n1037), .B(KEYINPUT30), .Z(n1221) );
NAND2_X1 U924 ( .A1(n1243), .A2(n1244), .ZN(G15) );
NAND2_X1 U925 ( .A1(G113), .A2(n1199), .ZN(n1244) );
XOR2_X1 U926 ( .A(KEYINPUT63), .B(n1245), .Z(n1243) );
NOR2_X1 U927 ( .A1(G113), .A2(n1199), .ZN(n1245) );
NAND2_X1 U928 ( .A1(n1066), .A2(n1242), .ZN(n1199) );
AND3_X1 U929 ( .A1(n1043), .A2(n1206), .A3(n1061), .ZN(n1242) );
NOR2_X1 U930 ( .A1(n1187), .A2(n1188), .ZN(n1061) );
NOR2_X1 U931 ( .A1(n1057), .A2(n1212), .ZN(n1043) );
INV_X1 U932 ( .A(n1184), .ZN(n1212) );
INV_X1 U933 ( .A(n1210), .ZN(n1057) );
NOR2_X1 U934 ( .A1(n1053), .A2(n1246), .ZN(n1210) );
NOR2_X1 U935 ( .A1(n1055), .A2(n1054), .ZN(n1246) );
INV_X1 U936 ( .A(n1247), .ZN(n1054) );
NOR2_X1 U937 ( .A1(n1037), .A2(n1248), .ZN(n1066) );
INV_X1 U938 ( .A(n1035), .ZN(n1248) );
XNOR2_X1 U939 ( .A(G110), .B(n1208), .ZN(G12) );
NAND3_X1 U940 ( .A1(n1188), .A2(n1209), .A3(n1249), .ZN(n1208) );
NOR3_X1 U941 ( .A1(n1035), .A2(n1062), .A3(n1037), .ZN(n1249) );
XOR2_X1 U942 ( .A(n1072), .B(KEYINPUT47), .Z(n1037) );
XNOR2_X1 U943 ( .A(n1250), .B(G478), .ZN(n1072) );
OR2_X1 U944 ( .A1(n1142), .A2(G902), .ZN(n1250) );
XNOR2_X1 U945 ( .A(n1251), .B(n1252), .ZN(n1142) );
XNOR2_X1 U946 ( .A(n1240), .B(n1253), .ZN(n1252) );
XNOR2_X1 U947 ( .A(n1254), .B(G122), .ZN(n1253) );
INV_X1 U948 ( .A(G116), .ZN(n1240) );
XNOR2_X1 U949 ( .A(n1255), .B(n1256), .ZN(n1251) );
XOR2_X1 U950 ( .A(n1257), .B(n1258), .Z(n1256) );
NAND2_X1 U951 ( .A1(KEYINPUT45), .A2(n1115), .ZN(n1258) );
INV_X1 U952 ( .A(G134), .ZN(n1115) );
NAND2_X1 U953 ( .A1(G217), .A2(n1259), .ZN(n1257) );
INV_X1 U954 ( .A(n1260), .ZN(n1259) );
INV_X1 U955 ( .A(n1187), .ZN(n1062) );
XNOR2_X1 U956 ( .A(n1076), .B(n1078), .ZN(n1187) );
XOR2_X1 U957 ( .A(G472), .B(KEYINPUT32), .Z(n1078) );
NAND2_X1 U958 ( .A1(n1154), .A2(n1261), .ZN(n1076) );
XOR2_X1 U959 ( .A(n1262), .B(n1263), .Z(n1154) );
XOR2_X1 U960 ( .A(n1264), .B(n1265), .Z(n1263) );
XOR2_X1 U961 ( .A(G113), .B(G101), .Z(n1265) );
XNOR2_X1 U962 ( .A(n1102), .B(G119), .ZN(n1264) );
XOR2_X1 U963 ( .A(n1266), .B(n1267), .Z(n1262) );
XOR2_X1 U964 ( .A(n1268), .B(n1269), .Z(n1267) );
AND2_X1 U965 ( .A1(n1270), .A2(G210), .ZN(n1268) );
XOR2_X1 U966 ( .A(n1271), .B(n1272), .Z(n1266) );
NOR2_X1 U967 ( .A1(KEYINPUT13), .A2(n1273), .ZN(n1272) );
XNOR2_X1 U968 ( .A(G116), .B(KEYINPUT19), .ZN(n1273) );
XNOR2_X1 U969 ( .A(n1274), .B(G475), .ZN(n1035) );
OR2_X1 U970 ( .A1(n1149), .A2(G902), .ZN(n1274) );
XNOR2_X1 U971 ( .A(n1275), .B(n1276), .ZN(n1149) );
XOR2_X1 U972 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U973 ( .A(n1279), .B(n1280), .Z(n1278) );
NOR2_X1 U974 ( .A1(G104), .A2(KEYINPUT56), .ZN(n1280) );
NOR2_X1 U975 ( .A1(G113), .A2(KEYINPUT6), .ZN(n1279) );
NOR2_X1 U976 ( .A1(n1281), .A2(n1282), .ZN(n1277) );
NOR2_X1 U977 ( .A1(n1099), .A2(n1283), .ZN(n1282) );
XNOR2_X1 U978 ( .A(KEYINPUT4), .B(n1097), .ZN(n1283) );
NOR2_X1 U979 ( .A1(G140), .A2(n1284), .ZN(n1281) );
XNOR2_X1 U980 ( .A(KEYINPUT62), .B(n1097), .ZN(n1284) );
XOR2_X1 U981 ( .A(n1285), .B(n1286), .Z(n1275) );
XNOR2_X1 U982 ( .A(n1287), .B(G122), .ZN(n1286) );
NAND2_X1 U983 ( .A1(n1288), .A2(KEYINPUT46), .ZN(n1285) );
XNOR2_X1 U984 ( .A(G131), .B(n1289), .ZN(n1288) );
NOR2_X1 U985 ( .A1(KEYINPUT15), .A2(n1290), .ZN(n1289) );
XNOR2_X1 U986 ( .A(G143), .B(n1291), .ZN(n1290) );
NAND2_X1 U987 ( .A1(G214), .A2(n1270), .ZN(n1291) );
NOR2_X1 U988 ( .A1(G953), .A2(G237), .ZN(n1270) );
INV_X1 U989 ( .A(n1202), .ZN(n1209) );
NAND3_X1 U990 ( .A1(n1184), .A2(n1206), .A3(n1052), .ZN(n1202) );
AND2_X1 U991 ( .A1(n1053), .A2(n1292), .ZN(n1052) );
NAND2_X1 U992 ( .A1(G221), .A2(n1247), .ZN(n1292) );
XNOR2_X1 U993 ( .A(n1293), .B(G469), .ZN(n1053) );
NAND2_X1 U994 ( .A1(n1294), .A2(n1261), .ZN(n1293) );
XNOR2_X1 U995 ( .A(n1295), .B(n1160), .ZN(n1294) );
XNOR2_X1 U996 ( .A(n1296), .B(n1297), .ZN(n1160) );
XOR2_X1 U997 ( .A(n1269), .B(n1093), .Z(n1297) );
XOR2_X1 U998 ( .A(G143), .B(G146), .Z(n1093) );
XNOR2_X1 U999 ( .A(n1298), .B(G131), .ZN(n1269) );
NAND2_X1 U1000 ( .A1(n1299), .A2(n1106), .ZN(n1298) );
INV_X1 U1001 ( .A(n1112), .ZN(n1106) );
NOR2_X1 U1002 ( .A1(n1110), .A2(G134), .ZN(n1112) );
XOR2_X1 U1003 ( .A(n1300), .B(KEYINPUT33), .Z(n1299) );
NAND2_X1 U1004 ( .A1(G134), .A2(n1110), .ZN(n1300) );
INV_X1 U1005 ( .A(G137), .ZN(n1110) );
XOR2_X1 U1006 ( .A(n1301), .B(n1302), .Z(n1296) );
XNOR2_X1 U1007 ( .A(KEYINPUT35), .B(n1303), .ZN(n1301) );
NOR2_X1 U1008 ( .A1(G101), .A2(KEYINPUT37), .ZN(n1303) );
NAND2_X1 U1009 ( .A1(n1164), .A2(n1304), .ZN(n1295) );
INV_X1 U1010 ( .A(n1162), .ZN(n1304) );
NOR3_X1 U1011 ( .A1(n1305), .A2(G953), .A3(n1085), .ZN(n1162) );
INV_X1 U1012 ( .A(G227), .ZN(n1085) );
NAND2_X1 U1013 ( .A1(n1305), .A2(n1306), .ZN(n1164) );
NAND2_X1 U1014 ( .A1(G227), .A2(n1084), .ZN(n1306) );
XNOR2_X1 U1015 ( .A(G140), .B(n1307), .ZN(n1305) );
NAND2_X1 U1016 ( .A1(n1032), .A2(n1308), .ZN(n1206) );
NAND2_X1 U1017 ( .A1(n1232), .A2(n1133), .ZN(n1308) );
INV_X1 U1018 ( .A(G898), .ZN(n1133) );
AND3_X1 U1019 ( .A1(G902), .A2(n1309), .A3(n1089), .ZN(n1232) );
XNOR2_X1 U1020 ( .A(G953), .B(KEYINPUT43), .ZN(n1089) );
NAND3_X1 U1021 ( .A1(n1309), .A2(n1084), .A3(G952), .ZN(n1032) );
NAND2_X1 U1022 ( .A1(G237), .A2(G234), .ZN(n1309) );
NOR2_X1 U1023 ( .A1(n1310), .A2(n1071), .ZN(n1184) );
INV_X1 U1024 ( .A(n1056), .ZN(n1071) );
NAND2_X1 U1025 ( .A1(G214), .A2(n1311), .ZN(n1056) );
INV_X1 U1026 ( .A(n1058), .ZN(n1310) );
XNOR2_X1 U1027 ( .A(n1075), .B(KEYINPUT16), .ZN(n1058) );
XNOR2_X1 U1028 ( .A(n1312), .B(n1216), .ZN(n1075) );
NAND2_X1 U1029 ( .A1(G210), .A2(n1311), .ZN(n1216) );
NAND2_X1 U1030 ( .A1(n1313), .A2(n1314), .ZN(n1311) );
INV_X1 U1031 ( .A(G237), .ZN(n1314) );
NAND2_X1 U1032 ( .A1(n1315), .A2(n1261), .ZN(n1312) );
XNOR2_X1 U1033 ( .A(n1167), .B(n1316), .ZN(n1315) );
XOR2_X1 U1034 ( .A(n1171), .B(KEYINPUT17), .Z(n1316) );
NAND2_X1 U1035 ( .A1(G224), .A2(n1084), .ZN(n1171) );
XNOR2_X1 U1036 ( .A(n1317), .B(n1318), .ZN(n1167) );
XOR2_X1 U1037 ( .A(n1302), .B(n1132), .Z(n1318) );
XNOR2_X1 U1038 ( .A(n1319), .B(n1320), .ZN(n1132) );
XOR2_X1 U1039 ( .A(n1321), .B(n1307), .Z(n1320) );
NAND3_X1 U1040 ( .A1(n1322), .A2(n1323), .A3(n1324), .ZN(n1321) );
NAND2_X1 U1041 ( .A1(G113), .A2(n1325), .ZN(n1324) );
NAND2_X1 U1042 ( .A1(n1326), .A2(n1327), .ZN(n1323) );
INV_X1 U1043 ( .A(KEYINPUT50), .ZN(n1327) );
NAND2_X1 U1044 ( .A1(n1328), .A2(n1329), .ZN(n1326) );
INV_X1 U1045 ( .A(n1325), .ZN(n1329) );
XNOR2_X1 U1046 ( .A(KEYINPUT24), .B(G113), .ZN(n1328) );
NAND2_X1 U1047 ( .A1(KEYINPUT50), .A2(n1330), .ZN(n1322) );
NAND2_X1 U1048 ( .A1(n1331), .A2(n1332), .ZN(n1330) );
OR3_X1 U1049 ( .A1(n1325), .A2(G113), .A3(KEYINPUT24), .ZN(n1332) );
XNOR2_X1 U1050 ( .A(G116), .B(n1333), .ZN(n1325) );
NAND2_X1 U1051 ( .A1(KEYINPUT24), .A2(G113), .ZN(n1331) );
XNOR2_X1 U1052 ( .A(G101), .B(G122), .ZN(n1319) );
XNOR2_X1 U1053 ( .A(n1131), .B(n1255), .ZN(n1302) );
XNOR2_X1 U1054 ( .A(G107), .B(n1102), .ZN(n1255) );
XNOR2_X1 U1055 ( .A(G104), .B(KEYINPUT23), .ZN(n1131) );
XNOR2_X1 U1056 ( .A(n1271), .B(n1097), .ZN(n1317) );
NAND3_X1 U1057 ( .A1(n1334), .A2(n1335), .A3(n1336), .ZN(n1271) );
OR2_X1 U1058 ( .A1(n1287), .A2(KEYINPUT55), .ZN(n1336) );
NAND3_X1 U1059 ( .A1(KEYINPUT55), .A2(n1287), .A3(G143), .ZN(n1335) );
NAND2_X1 U1060 ( .A1(n1337), .A2(n1254), .ZN(n1334) );
INV_X1 U1061 ( .A(G143), .ZN(n1254) );
NAND2_X1 U1062 ( .A1(KEYINPUT55), .A2(n1338), .ZN(n1337) );
XNOR2_X1 U1063 ( .A(KEYINPUT29), .B(n1287), .ZN(n1338) );
INV_X1 U1064 ( .A(n1063), .ZN(n1188) );
XNOR2_X1 U1065 ( .A(n1339), .B(n1340), .ZN(n1063) );
XNOR2_X1 U1066 ( .A(KEYINPUT60), .B(n1074), .ZN(n1340) );
NAND2_X1 U1067 ( .A1(G217), .A2(n1247), .ZN(n1074) );
NAND2_X1 U1068 ( .A1(n1313), .A2(G234), .ZN(n1247) );
XNOR2_X1 U1069 ( .A(G902), .B(KEYINPUT22), .ZN(n1313) );
NAND2_X1 U1070 ( .A1(KEYINPUT28), .A2(n1073), .ZN(n1339) );
NAND2_X1 U1071 ( .A1(n1137), .A2(n1261), .ZN(n1073) );
INV_X1 U1072 ( .A(G902), .ZN(n1261) );
XNOR2_X1 U1073 ( .A(n1341), .B(n1342), .ZN(n1137) );
XOR2_X1 U1074 ( .A(n1307), .B(n1343), .Z(n1342) );
XOR2_X1 U1075 ( .A(n1344), .B(n1345), .Z(n1343) );
NOR2_X1 U1076 ( .A1(n1260), .A2(n1055), .ZN(n1345) );
INV_X1 U1077 ( .A(G221), .ZN(n1055) );
NAND2_X1 U1078 ( .A1(G234), .A2(n1084), .ZN(n1260) );
INV_X1 U1079 ( .A(G953), .ZN(n1084) );
NAND2_X1 U1080 ( .A1(n1346), .A2(n1347), .ZN(n1344) );
NAND2_X1 U1081 ( .A1(G125), .A2(n1099), .ZN(n1347) );
INV_X1 U1082 ( .A(G140), .ZN(n1099) );
XOR2_X1 U1083 ( .A(n1348), .B(KEYINPUT26), .Z(n1346) );
NAND2_X1 U1084 ( .A1(G140), .A2(n1097), .ZN(n1348) );
INV_X1 U1085 ( .A(G125), .ZN(n1097) );
XNOR2_X1 U1086 ( .A(G110), .B(KEYINPUT2), .ZN(n1307) );
XOR2_X1 U1087 ( .A(n1349), .B(n1350), .Z(n1341) );
XNOR2_X1 U1088 ( .A(n1287), .B(G137), .ZN(n1350) );
INV_X1 U1089 ( .A(G146), .ZN(n1287) );
NAND3_X1 U1090 ( .A1(n1351), .A2(n1352), .A3(n1353), .ZN(n1349) );
NAND2_X1 U1091 ( .A1(KEYINPUT54), .A2(G128), .ZN(n1353) );
NAND3_X1 U1092 ( .A1(n1102), .A2(n1354), .A3(G119), .ZN(n1352) );
INV_X1 U1093 ( .A(G128), .ZN(n1102) );
NAND2_X1 U1094 ( .A1(n1355), .A2(n1333), .ZN(n1351) );
INV_X1 U1095 ( .A(G119), .ZN(n1333) );
NAND2_X1 U1096 ( .A1(n1356), .A2(n1354), .ZN(n1355) );
INV_X1 U1097 ( .A(KEYINPUT54), .ZN(n1354) );
XNOR2_X1 U1098 ( .A(G128), .B(KEYINPUT42), .ZN(n1356) );
endmodule


