//Key = 1100100111110011011100010100110011010000011000101110011011100011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;

XNOR2_X1 U733 ( .A(n1010), .B(n1011), .ZN(G9) );
NOR3_X1 U734 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n1011) );
XNOR2_X1 U735 ( .A(KEYINPUT58), .B(n1015), .ZN(n1012) );
NOR2_X1 U736 ( .A1(n1016), .A2(n1017), .ZN(G75) );
NOR4_X1 U737 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .ZN(n1017) );
NOR2_X1 U738 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR3_X1 U739 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n1020) );
XOR2_X1 U740 ( .A(n1023), .B(KEYINPUT51), .Z(n1025) );
NAND4_X1 U741 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1023) );
NAND3_X1 U742 ( .A1(n1031), .A2(n1032), .A3(n1033), .ZN(n1018) );
NAND3_X1 U743 ( .A1(n1034), .A2(n1035), .A3(n1027), .ZN(n1033) );
INV_X1 U744 ( .A(n1036), .ZN(n1027) );
NAND2_X1 U745 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NAND3_X1 U746 ( .A1(n1030), .A2(n1039), .A3(n1029), .ZN(n1038) );
NAND2_X1 U747 ( .A1(n1028), .A2(n1040), .ZN(n1037) );
NAND2_X1 U748 ( .A1(n1041), .A2(n1042), .ZN(n1040) );
NAND2_X1 U749 ( .A1(n1030), .A2(n1043), .ZN(n1042) );
NAND2_X1 U750 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NAND2_X1 U751 ( .A1(n1046), .A2(n1047), .ZN(n1045) );
NAND2_X1 U752 ( .A1(n1029), .A2(n1048), .ZN(n1041) );
NAND2_X1 U753 ( .A1(n1049), .A2(n1050), .ZN(n1048) );
NOR3_X1 U754 ( .A1(n1051), .A2(G953), .A3(G952), .ZN(n1016) );
INV_X1 U755 ( .A(n1031), .ZN(n1051) );
NAND4_X1 U756 ( .A1(n1052), .A2(n1034), .A3(n1053), .A4(n1054), .ZN(n1031) );
NOR4_X1 U757 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1054) );
NOR2_X1 U758 ( .A1(n1059), .A2(n1060), .ZN(n1058) );
AND2_X1 U759 ( .A1(n1061), .A2(G475), .ZN(n1057) );
INV_X1 U760 ( .A(n1062), .ZN(n1056) );
NOR2_X1 U761 ( .A1(n1063), .A2(n1064), .ZN(n1053) );
XNOR2_X1 U762 ( .A(n1065), .B(KEYINPUT4), .ZN(n1052) );
XOR2_X1 U763 ( .A(n1066), .B(n1067), .Z(G72) );
XOR2_X1 U764 ( .A(n1068), .B(n1069), .Z(n1067) );
NOR2_X1 U765 ( .A1(n1070), .A2(n1071), .ZN(n1069) );
XOR2_X1 U766 ( .A(n1072), .B(n1073), .Z(n1071) );
XOR2_X1 U767 ( .A(n1074), .B(n1075), .Z(n1073) );
XOR2_X1 U768 ( .A(n1076), .B(n1077), .Z(n1075) );
XOR2_X1 U769 ( .A(n1078), .B(n1079), .Z(n1072) );
XNOR2_X1 U770 ( .A(n1080), .B(G134), .ZN(n1079) );
XOR2_X1 U771 ( .A(KEYINPUT60), .B(KEYINPUT18), .Z(n1078) );
NOR2_X1 U772 ( .A1(G900), .A2(n1032), .ZN(n1070) );
NOR2_X1 U773 ( .A1(KEYINPUT40), .A2(n1081), .ZN(n1068) );
NOR2_X1 U774 ( .A1(n1082), .A2(n1032), .ZN(n1081) );
AND2_X1 U775 ( .A1(G227), .A2(G900), .ZN(n1082) );
NAND2_X1 U776 ( .A1(n1032), .A2(n1083), .ZN(n1066) );
NAND2_X1 U777 ( .A1(n1084), .A2(n1085), .ZN(G69) );
NAND2_X1 U778 ( .A1(n1086), .A2(n1087), .ZN(n1085) );
NAND2_X1 U779 ( .A1(G953), .A2(n1088), .ZN(n1087) );
NAND2_X1 U780 ( .A1(G898), .A2(G224), .ZN(n1088) );
NAND2_X1 U781 ( .A1(n1089), .A2(n1090), .ZN(n1084) );
NAND2_X1 U782 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
NAND2_X1 U783 ( .A1(G953), .A2(n1093), .ZN(n1092) );
INV_X1 U784 ( .A(n1086), .ZN(n1089) );
NAND2_X1 U785 ( .A1(n1094), .A2(n1095), .ZN(n1086) );
NAND2_X1 U786 ( .A1(n1096), .A2(n1097), .ZN(n1095) );
INV_X1 U787 ( .A(n1098), .ZN(n1096) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1098), .ZN(n1094) );
NAND2_X1 U789 ( .A1(n1100), .A2(n1091), .ZN(n1098) );
INV_X1 U790 ( .A(n1101), .ZN(n1091) );
XOR2_X1 U791 ( .A(KEYINPUT34), .B(n1102), .Z(n1100) );
NOR2_X1 U792 ( .A1(n1103), .A2(n1104), .ZN(n1102) );
NOR2_X1 U793 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XNOR2_X1 U794 ( .A(n1107), .B(KEYINPUT28), .ZN(n1105) );
INV_X1 U795 ( .A(n1108), .ZN(n1103) );
XOR2_X1 U796 ( .A(n1097), .B(KEYINPUT63), .Z(n1099) );
NAND2_X1 U797 ( .A1(n1109), .A2(n1110), .ZN(n1097) );
NAND2_X1 U798 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
INV_X1 U799 ( .A(n1113), .ZN(n1112) );
XOR2_X1 U800 ( .A(n1114), .B(KEYINPUT15), .Z(n1111) );
XNOR2_X1 U801 ( .A(G953), .B(KEYINPUT22), .ZN(n1109) );
NOR2_X1 U802 ( .A1(n1115), .A2(n1116), .ZN(G66) );
XOR2_X1 U803 ( .A(n1117), .B(n1118), .Z(n1116) );
NAND2_X1 U804 ( .A1(n1119), .A2(n1120), .ZN(n1117) );
INV_X1 U805 ( .A(n1060), .ZN(n1120) );
NOR2_X1 U806 ( .A1(n1115), .A2(n1121), .ZN(G63) );
XOR2_X1 U807 ( .A(n1122), .B(n1123), .Z(n1121) );
NAND2_X1 U808 ( .A1(n1119), .A2(G478), .ZN(n1122) );
NOR2_X1 U809 ( .A1(n1115), .A2(n1124), .ZN(G60) );
XOR2_X1 U810 ( .A(n1125), .B(n1126), .Z(n1124) );
NAND2_X1 U811 ( .A1(n1119), .A2(G475), .ZN(n1125) );
NAND2_X1 U812 ( .A1(n1127), .A2(n1128), .ZN(G6) );
OR2_X1 U813 ( .A1(n1129), .A2(G104), .ZN(n1128) );
XOR2_X1 U814 ( .A(n1130), .B(KEYINPUT12), .Z(n1127) );
NAND2_X1 U815 ( .A1(G104), .A2(n1129), .ZN(n1130) );
NAND2_X1 U816 ( .A1(n1131), .A2(n1132), .ZN(n1129) );
XOR2_X1 U817 ( .A(KEYINPUT36), .B(n1133), .Z(n1132) );
NOR2_X1 U818 ( .A1(n1013), .A2(n1134), .ZN(n1133) );
NOR2_X1 U819 ( .A1(n1115), .A2(n1135), .ZN(G57) );
XOR2_X1 U820 ( .A(n1136), .B(n1137), .Z(n1135) );
XOR2_X1 U821 ( .A(n1138), .B(n1139), .Z(n1137) );
NAND2_X1 U822 ( .A1(n1119), .A2(G472), .ZN(n1139) );
NAND2_X1 U823 ( .A1(n1140), .A2(KEYINPUT54), .ZN(n1138) );
XOR2_X1 U824 ( .A(n1141), .B(n1142), .Z(n1140) );
XNOR2_X1 U825 ( .A(KEYINPUT61), .B(KEYINPUT2), .ZN(n1141) );
NOR2_X1 U826 ( .A1(n1115), .A2(n1143), .ZN(G54) );
XOR2_X1 U827 ( .A(n1144), .B(n1145), .Z(n1143) );
XOR2_X1 U828 ( .A(n1146), .B(n1147), .Z(n1144) );
NOR3_X1 U829 ( .A1(n1148), .A2(n1149), .A3(n1150), .ZN(n1147) );
NOR2_X1 U830 ( .A1(n1151), .A2(n1152), .ZN(n1150) );
INV_X1 U831 ( .A(KEYINPUT52), .ZN(n1152) );
NOR2_X1 U832 ( .A1(KEYINPUT52), .A2(n1153), .ZN(n1149) );
NAND2_X1 U833 ( .A1(n1119), .A2(G469), .ZN(n1146) );
NOR2_X1 U834 ( .A1(n1115), .A2(n1154), .ZN(G51) );
XOR2_X1 U835 ( .A(n1155), .B(n1156), .Z(n1154) );
XOR2_X1 U836 ( .A(n1157), .B(n1158), .Z(n1156) );
XOR2_X1 U837 ( .A(n1159), .B(n1160), .Z(n1158) );
NAND2_X1 U838 ( .A1(KEYINPUT50), .A2(n1161), .ZN(n1157) );
INV_X1 U839 ( .A(G125), .ZN(n1161) );
XNOR2_X1 U840 ( .A(n1162), .B(n1163), .ZN(n1155) );
NAND3_X1 U841 ( .A1(n1119), .A2(G210), .A3(KEYINPUT57), .ZN(n1162) );
AND2_X1 U842 ( .A1(G902), .A2(n1019), .ZN(n1119) );
OR3_X1 U843 ( .A1(n1113), .A2(n1114), .A3(n1083), .ZN(n1019) );
NAND4_X1 U844 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1083) );
AND4_X1 U845 ( .A1(n1168), .A2(n1169), .A3(n1170), .A4(n1171), .ZN(n1167) );
NAND2_X1 U846 ( .A1(n1172), .A2(n1039), .ZN(n1166) );
INV_X1 U847 ( .A(n1173), .ZN(n1172) );
NAND2_X1 U848 ( .A1(n1174), .A2(n1175), .ZN(n1164) );
NAND3_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .ZN(n1114) );
NAND3_X1 U850 ( .A1(n1131), .A2(n1039), .A3(n1179), .ZN(n1178) );
INV_X1 U851 ( .A(n1013), .ZN(n1179) );
NAND3_X1 U852 ( .A1(n1030), .A2(n1180), .A3(n1181), .ZN(n1013) );
NAND2_X1 U853 ( .A1(n1134), .A2(n1014), .ZN(n1039) );
NAND4_X1 U854 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1113) );
NOR2_X1 U855 ( .A1(n1186), .A2(n1187), .ZN(n1182) );
NOR2_X1 U856 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
INV_X1 U857 ( .A(KEYINPUT33), .ZN(n1188) );
NOR4_X1 U858 ( .A1(KEYINPUT33), .A2(n1190), .A3(n1063), .A4(n1049), .ZN(n1186) );
INV_X1 U859 ( .A(n1191), .ZN(n1049) );
NAND3_X1 U860 ( .A1(n1022), .A2(n1180), .A3(n1192), .ZN(n1190) );
NOR2_X1 U861 ( .A1(n1032), .A2(G952), .ZN(n1115) );
NAND2_X1 U862 ( .A1(n1193), .A2(n1194), .ZN(G48) );
NAND2_X1 U863 ( .A1(KEYINPUT3), .A2(n1195), .ZN(n1194) );
XOR2_X1 U864 ( .A(n1196), .B(n1197), .Z(n1193) );
NOR2_X1 U865 ( .A1(n1134), .A2(n1173), .ZN(n1197) );
OR2_X1 U866 ( .A1(n1195), .A2(KEYINPUT3), .ZN(n1196) );
XNOR2_X1 U867 ( .A(G143), .B(n1165), .ZN(G45) );
NAND4_X1 U868 ( .A1(n1198), .A2(n1191), .A3(n1199), .A4(n1200), .ZN(n1165) );
XNOR2_X1 U869 ( .A(G140), .B(n1171), .ZN(G42) );
NAND3_X1 U870 ( .A1(n1201), .A2(n1202), .A3(n1175), .ZN(n1171) );
XNOR2_X1 U871 ( .A(G137), .B(n1203), .ZN(G39) );
NAND4_X1 U872 ( .A1(n1204), .A2(n1174), .A3(n1034), .A4(n1181), .ZN(n1203) );
XNOR2_X1 U873 ( .A(n1205), .B(KEYINPUT47), .ZN(n1204) );
XNOR2_X1 U874 ( .A(G134), .B(n1170), .ZN(G36) );
NAND3_X1 U875 ( .A1(n1175), .A2(n1192), .A3(n1191), .ZN(n1170) );
XNOR2_X1 U876 ( .A(G131), .B(n1169), .ZN(G33) );
NAND3_X1 U877 ( .A1(n1175), .A2(n1201), .A3(n1191), .ZN(n1169) );
AND3_X1 U878 ( .A1(n1181), .A2(n1206), .A3(n1034), .ZN(n1175) );
NOR2_X1 U879 ( .A1(n1026), .A2(n1207), .ZN(n1034) );
XOR2_X1 U880 ( .A(G128), .B(n1208), .Z(G30) );
NOR2_X1 U881 ( .A1(n1173), .A2(n1209), .ZN(n1208) );
XNOR2_X1 U882 ( .A(KEYINPUT1), .B(n1014), .ZN(n1209) );
INV_X1 U883 ( .A(n1192), .ZN(n1014) );
NAND3_X1 U884 ( .A1(n1064), .A2(n1210), .A3(n1198), .ZN(n1173) );
NOR3_X1 U885 ( .A1(n1022), .A2(n1205), .A3(n1044), .ZN(n1198) );
INV_X1 U886 ( .A(n1181), .ZN(n1044) );
XNOR2_X1 U887 ( .A(G101), .B(n1176), .ZN(G3) );
NAND2_X1 U888 ( .A1(n1211), .A2(n1191), .ZN(n1176) );
XNOR2_X1 U889 ( .A(G125), .B(n1212), .ZN(G27) );
NAND2_X1 U890 ( .A1(KEYINPUT62), .A2(n1213), .ZN(n1212) );
INV_X1 U891 ( .A(n1168), .ZN(n1213) );
NAND4_X1 U892 ( .A1(n1201), .A2(n1202), .A3(n1214), .A4(n1029), .ZN(n1168) );
INV_X1 U893 ( .A(n1063), .ZN(n1029) );
NOR2_X1 U894 ( .A1(n1205), .A2(n1022), .ZN(n1214) );
INV_X1 U895 ( .A(n1206), .ZN(n1205) );
NAND2_X1 U896 ( .A1(n1036), .A2(n1215), .ZN(n1206) );
NAND4_X1 U897 ( .A1(G902), .A2(G953), .A3(n1216), .A4(n1217), .ZN(n1215) );
INV_X1 U898 ( .A(G900), .ZN(n1217) );
XNOR2_X1 U899 ( .A(G122), .B(n1183), .ZN(G24) );
NAND4_X1 U900 ( .A1(n1218), .A2(n1030), .A3(n1199), .A4(n1200), .ZN(n1183) );
NOR2_X1 U901 ( .A1(n1210), .A2(n1064), .ZN(n1030) );
XNOR2_X1 U902 ( .A(G119), .B(n1184), .ZN(G21) );
NAND2_X1 U903 ( .A1(n1218), .A2(n1174), .ZN(n1184) );
AND3_X1 U904 ( .A1(n1064), .A2(n1210), .A3(n1028), .ZN(n1174) );
XOR2_X1 U905 ( .A(n1189), .B(n1219), .Z(G18) );
NAND2_X1 U906 ( .A1(KEYINPUT23), .A2(G116), .ZN(n1219) );
NAND3_X1 U907 ( .A1(n1191), .A2(n1192), .A3(n1218), .ZN(n1189) );
NOR3_X1 U908 ( .A1(n1022), .A2(n1220), .A3(n1063), .ZN(n1218) );
XOR2_X1 U909 ( .A(n1015), .B(KEYINPUT20), .Z(n1022) );
NOR2_X1 U910 ( .A1(n1200), .A2(n1065), .ZN(n1192) );
XNOR2_X1 U911 ( .A(G113), .B(n1185), .ZN(G15) );
NAND3_X1 U912 ( .A1(n1191), .A2(n1201), .A3(n1221), .ZN(n1185) );
NOR3_X1 U913 ( .A1(n1063), .A2(n1220), .A3(n1015), .ZN(n1221) );
INV_X1 U914 ( .A(n1180), .ZN(n1220) );
NAND2_X1 U915 ( .A1(n1047), .A2(n1222), .ZN(n1063) );
INV_X1 U916 ( .A(n1134), .ZN(n1201) );
NAND2_X1 U917 ( .A1(n1065), .A2(n1200), .ZN(n1134) );
NOR2_X1 U918 ( .A1(n1210), .A2(n1223), .ZN(n1191) );
XNOR2_X1 U919 ( .A(n1224), .B(n1177), .ZN(G12) );
NAND2_X1 U920 ( .A1(n1211), .A2(n1202), .ZN(n1177) );
INV_X1 U921 ( .A(n1050), .ZN(n1202) );
NAND2_X1 U922 ( .A1(n1223), .A2(n1210), .ZN(n1050) );
NAND3_X1 U923 ( .A1(n1225), .A2(n1226), .A3(n1062), .ZN(n1210) );
NAND2_X1 U924 ( .A1(n1059), .A2(n1060), .ZN(n1062) );
NAND2_X1 U925 ( .A1(KEYINPUT59), .A2(n1060), .ZN(n1226) );
OR3_X1 U926 ( .A1(n1059), .A2(KEYINPUT59), .A3(n1060), .ZN(n1225) );
NAND2_X1 U927 ( .A1(G217), .A2(n1227), .ZN(n1060) );
AND2_X1 U928 ( .A1(n1118), .A2(n1228), .ZN(n1059) );
XOR2_X1 U929 ( .A(n1229), .B(n1230), .Z(n1118) );
XOR2_X1 U930 ( .A(n1231), .B(n1232), .Z(n1230) );
XNOR2_X1 U931 ( .A(KEYINPUT13), .B(n1233), .ZN(n1232) );
NOR2_X1 U932 ( .A1(KEYINPUT37), .A2(n1234), .ZN(n1233) );
XNOR2_X1 U933 ( .A(G110), .B(n1235), .ZN(n1234) );
XNOR2_X1 U934 ( .A(G128), .B(n1236), .ZN(n1235) );
NAND3_X1 U935 ( .A1(G234), .A2(n1032), .A3(G221), .ZN(n1231) );
XOR2_X1 U936 ( .A(n1076), .B(n1237), .Z(n1229) );
XNOR2_X1 U937 ( .A(n1238), .B(n1239), .ZN(n1237) );
NOR2_X1 U938 ( .A1(G140), .A2(KEYINPUT21), .ZN(n1239) );
NAND2_X1 U939 ( .A1(KEYINPUT10), .A2(G146), .ZN(n1238) );
XNOR2_X1 U940 ( .A(G137), .B(G125), .ZN(n1076) );
INV_X1 U941 ( .A(n1064), .ZN(n1223) );
XNOR2_X1 U942 ( .A(n1240), .B(G472), .ZN(n1064) );
NAND2_X1 U943 ( .A1(n1241), .A2(n1228), .ZN(n1240) );
XOR2_X1 U944 ( .A(n1242), .B(n1142), .Z(n1241) );
XOR2_X1 U945 ( .A(G101), .B(n1243), .Z(n1142) );
NOR3_X1 U946 ( .A1(n1244), .A2(G953), .A3(G237), .ZN(n1243) );
XNOR2_X1 U947 ( .A(n1136), .B(KEYINPUT46), .ZN(n1242) );
XNOR2_X1 U948 ( .A(n1245), .B(n1246), .ZN(n1136) );
XNOR2_X1 U949 ( .A(n1247), .B(n1248), .ZN(n1246) );
XNOR2_X1 U950 ( .A(G113), .B(n1249), .ZN(n1245) );
XNOR2_X1 U951 ( .A(n1236), .B(G116), .ZN(n1249) );
AND4_X1 U952 ( .A1(n1028), .A2(n1131), .A3(n1181), .A4(n1180), .ZN(n1211) );
NAND2_X1 U953 ( .A1(n1036), .A2(n1250), .ZN(n1180) );
NAND3_X1 U954 ( .A1(G902), .A2(n1216), .A3(n1101), .ZN(n1250) );
NOR2_X1 U955 ( .A1(n1032), .A2(G898), .ZN(n1101) );
NAND3_X1 U956 ( .A1(n1216), .A2(n1032), .A3(G952), .ZN(n1036) );
NAND2_X1 U957 ( .A1(G237), .A2(G234), .ZN(n1216) );
NOR2_X1 U958 ( .A1(n1047), .A2(n1046), .ZN(n1181) );
INV_X1 U959 ( .A(n1222), .ZN(n1046) );
NAND2_X1 U960 ( .A1(G221), .A2(n1227), .ZN(n1222) );
NAND2_X1 U961 ( .A1(G234), .A2(n1228), .ZN(n1227) );
XNOR2_X1 U962 ( .A(n1251), .B(n1252), .ZN(n1047) );
XOR2_X1 U963 ( .A(KEYINPUT41), .B(G469), .Z(n1252) );
NAND2_X1 U964 ( .A1(n1253), .A2(n1228), .ZN(n1251) );
XOR2_X1 U965 ( .A(n1145), .B(n1254), .Z(n1253) );
XOR2_X1 U966 ( .A(KEYINPUT24), .B(n1255), .Z(n1254) );
NOR2_X1 U967 ( .A1(n1148), .A2(n1256), .ZN(n1255) );
INV_X1 U968 ( .A(n1153), .ZN(n1256) );
NAND2_X1 U969 ( .A1(n1257), .A2(n1151), .ZN(n1153) );
NOR2_X1 U970 ( .A1(n1151), .A2(n1257), .ZN(n1148) );
XNOR2_X1 U971 ( .A(G110), .B(n1080), .ZN(n1257) );
NAND2_X1 U972 ( .A1(G227), .A2(n1032), .ZN(n1151) );
INV_X1 U973 ( .A(G953), .ZN(n1032) );
XNOR2_X1 U974 ( .A(n1074), .B(n1258), .ZN(n1145) );
XOR2_X1 U975 ( .A(n1259), .B(n1248), .Z(n1258) );
XNOR2_X1 U976 ( .A(n1077), .B(n1260), .ZN(n1248) );
NOR2_X1 U977 ( .A1(KEYINPUT26), .A2(n1261), .ZN(n1260) );
XOR2_X1 U978 ( .A(n1262), .B(n1263), .Z(n1261) );
NOR2_X1 U979 ( .A1(KEYINPUT44), .A2(G134), .ZN(n1263) );
XNOR2_X1 U980 ( .A(G137), .B(KEYINPUT0), .ZN(n1262) );
XOR2_X1 U981 ( .A(G131), .B(G128), .Z(n1077) );
XNOR2_X1 U982 ( .A(n1264), .B(n1265), .ZN(n1074) );
NAND2_X1 U983 ( .A1(KEYINPUT48), .A2(n1195), .ZN(n1264) );
INV_X1 U984 ( .A(n1015), .ZN(n1131) );
NAND2_X1 U985 ( .A1(n1026), .A2(n1024), .ZN(n1015) );
INV_X1 U986 ( .A(n1207), .ZN(n1024) );
NOR2_X1 U987 ( .A1(n1266), .A2(n1267), .ZN(n1207) );
XNOR2_X1 U988 ( .A(n1268), .B(n1269), .ZN(n1026) );
NOR2_X1 U989 ( .A1(n1267), .A2(n1270), .ZN(n1269) );
XNOR2_X1 U990 ( .A(KEYINPUT9), .B(n1244), .ZN(n1270) );
INV_X1 U991 ( .A(G210), .ZN(n1244) );
NOR2_X1 U992 ( .A1(G237), .A2(G902), .ZN(n1267) );
NAND2_X1 U993 ( .A1(n1271), .A2(n1228), .ZN(n1268) );
XOR2_X1 U994 ( .A(n1272), .B(n1159), .Z(n1271) );
NAND2_X1 U995 ( .A1(n1108), .A2(n1273), .ZN(n1159) );
OR2_X1 U996 ( .A1(n1106), .A2(n1107), .ZN(n1273) );
NAND2_X1 U997 ( .A1(n1107), .A2(n1106), .ZN(n1108) );
NAND2_X1 U998 ( .A1(n1274), .A2(n1275), .ZN(n1106) );
NAND2_X1 U999 ( .A1(n1276), .A2(n1277), .ZN(n1275) );
XNOR2_X1 U1000 ( .A(G116), .B(n1278), .ZN(n1277) );
XNOR2_X1 U1001 ( .A(KEYINPUT8), .B(n1279), .ZN(n1276) );
INV_X1 U1002 ( .A(G113), .ZN(n1279) );
XOR2_X1 U1003 ( .A(n1280), .B(KEYINPUT27), .Z(n1274) );
NAND2_X1 U1004 ( .A1(n1281), .A2(n1282), .ZN(n1280) );
XOR2_X1 U1005 ( .A(n1278), .B(G116), .Z(n1282) );
NAND2_X1 U1006 ( .A1(KEYINPUT35), .A2(n1236), .ZN(n1278) );
INV_X1 U1007 ( .A(G119), .ZN(n1236) );
XNOR2_X1 U1008 ( .A(KEYINPUT8), .B(G113), .ZN(n1281) );
XNOR2_X1 U1009 ( .A(n1259), .B(n1283), .ZN(n1107) );
XNOR2_X1 U1010 ( .A(G122), .B(n1284), .ZN(n1283) );
XNOR2_X1 U1011 ( .A(G101), .B(n1285), .ZN(n1259) );
XNOR2_X1 U1012 ( .A(n1010), .B(G104), .ZN(n1285) );
INV_X1 U1013 ( .A(G107), .ZN(n1010) );
NAND2_X1 U1014 ( .A1(n1286), .A2(KEYINPUT17), .ZN(n1272) );
XOR2_X1 U1015 ( .A(n1287), .B(n1160), .Z(n1286) );
NOR2_X1 U1016 ( .A1(n1093), .A2(G953), .ZN(n1160) );
INV_X1 U1017 ( .A(G224), .ZN(n1093) );
NAND3_X1 U1018 ( .A1(n1288), .A2(n1289), .A3(KEYINPUT7), .ZN(n1287) );
NAND2_X1 U1019 ( .A1(n1290), .A2(n1291), .ZN(n1289) );
INV_X1 U1020 ( .A(KEYINPUT38), .ZN(n1291) );
XNOR2_X1 U1021 ( .A(n1292), .B(G125), .ZN(n1290) );
INV_X1 U1022 ( .A(n1163), .ZN(n1292) );
NAND3_X1 U1023 ( .A1(G125), .A2(n1163), .A3(KEYINPUT38), .ZN(n1288) );
XOR2_X1 U1024 ( .A(G128), .B(n1293), .Z(n1163) );
INV_X1 U1025 ( .A(n1247), .ZN(n1293) );
XNOR2_X1 U1026 ( .A(n1294), .B(n1295), .ZN(n1247) );
NOR2_X1 U1027 ( .A1(KEYINPUT55), .A2(n1265), .ZN(n1295) );
XNOR2_X1 U1028 ( .A(G146), .B(KEYINPUT5), .ZN(n1294) );
NOR2_X1 U1029 ( .A1(n1200), .A2(n1199), .ZN(n1028) );
INV_X1 U1030 ( .A(n1065), .ZN(n1199) );
XNOR2_X1 U1031 ( .A(n1296), .B(n1297), .ZN(n1065) );
XOR2_X1 U1032 ( .A(KEYINPUT32), .B(G478), .Z(n1297) );
NAND2_X1 U1033 ( .A1(n1298), .A2(n1123), .ZN(n1296) );
XNOR2_X1 U1034 ( .A(n1299), .B(n1300), .ZN(n1123) );
AND3_X1 U1035 ( .A1(n1301), .A2(G217), .A3(G234), .ZN(n1300) );
XNOR2_X1 U1036 ( .A(KEYINPUT43), .B(G953), .ZN(n1301) );
NAND2_X1 U1037 ( .A1(KEYINPUT19), .A2(n1302), .ZN(n1299) );
NAND2_X1 U1038 ( .A1(n1303), .A2(n1304), .ZN(n1302) );
NAND2_X1 U1039 ( .A1(n1305), .A2(n1306), .ZN(n1304) );
INV_X1 U1040 ( .A(n1307), .ZN(n1305) );
XOR2_X1 U1041 ( .A(n1308), .B(KEYINPUT31), .Z(n1303) );
NAND2_X1 U1042 ( .A1(n1309), .A2(n1307), .ZN(n1308) );
XNOR2_X1 U1043 ( .A(n1310), .B(n1311), .ZN(n1307) );
XOR2_X1 U1044 ( .A(G122), .B(G116), .Z(n1311) );
NAND2_X1 U1045 ( .A1(n1312), .A2(KEYINPUT14), .ZN(n1310) );
XNOR2_X1 U1046 ( .A(G107), .B(KEYINPUT16), .ZN(n1312) );
XNOR2_X1 U1047 ( .A(n1306), .B(KEYINPUT39), .ZN(n1309) );
XNOR2_X1 U1048 ( .A(n1313), .B(G134), .ZN(n1306) );
NAND3_X1 U1049 ( .A1(n1314), .A2(n1315), .A3(KEYINPUT53), .ZN(n1313) );
NAND2_X1 U1050 ( .A1(G128), .A2(n1265), .ZN(n1315) );
XOR2_X1 U1051 ( .A(KEYINPUT42), .B(n1316), .Z(n1314) );
NOR2_X1 U1052 ( .A1(G128), .A2(n1265), .ZN(n1316) );
INV_X1 U1053 ( .A(G143), .ZN(n1265) );
XNOR2_X1 U1054 ( .A(KEYINPUT25), .B(n1228), .ZN(n1298) );
NAND2_X1 U1055 ( .A1(n1317), .A2(n1318), .ZN(n1200) );
NAND2_X1 U1056 ( .A1(G475), .A2(n1061), .ZN(n1318) );
XNOR2_X1 U1057 ( .A(n1055), .B(KEYINPUT6), .ZN(n1317) );
NOR2_X1 U1058 ( .A1(n1061), .A2(G475), .ZN(n1055) );
NAND2_X1 U1059 ( .A1(n1126), .A2(n1228), .ZN(n1061) );
INV_X1 U1060 ( .A(G902), .ZN(n1228) );
XOR2_X1 U1061 ( .A(n1319), .B(n1320), .Z(n1126) );
XOR2_X1 U1062 ( .A(n1321), .B(n1322), .Z(n1320) );
XNOR2_X1 U1063 ( .A(n1323), .B(n1324), .ZN(n1322) );
NOR4_X1 U1064 ( .A1(n1325), .A2(n1326), .A3(KEYINPUT45), .A4(n1327), .ZN(n1324) );
AND2_X1 U1065 ( .A1(n1328), .A2(G104), .ZN(n1327) );
NOR2_X1 U1066 ( .A1(n1329), .A2(n1330), .ZN(n1326) );
INV_X1 U1067 ( .A(n1331), .ZN(n1330) );
NOR2_X1 U1068 ( .A1(n1328), .A2(n1332), .ZN(n1329) );
XOR2_X1 U1069 ( .A(KEYINPUT30), .B(G104), .Z(n1332) );
NOR3_X1 U1070 ( .A1(n1331), .A2(G104), .A3(n1328), .ZN(n1325) );
INV_X1 U1071 ( .A(KEYINPUT49), .ZN(n1328) );
XOR2_X1 U1072 ( .A(G113), .B(G122), .Z(n1331) );
NAND2_X1 U1073 ( .A1(KEYINPUT29), .A2(n1080), .ZN(n1323) );
INV_X1 U1074 ( .A(G140), .ZN(n1080) );
NOR2_X1 U1075 ( .A1(n1333), .A2(n1334), .ZN(n1321) );
AND2_X1 U1076 ( .A1(G143), .A2(n1335), .ZN(n1334) );
NOR2_X1 U1077 ( .A1(n1335), .A2(n1336), .ZN(n1333) );
XNOR2_X1 U1078 ( .A(G143), .B(KEYINPUT56), .ZN(n1336) );
NOR3_X1 U1079 ( .A1(G237), .A2(G953), .A3(n1266), .ZN(n1335) );
INV_X1 U1080 ( .A(G214), .ZN(n1266) );
XNOR2_X1 U1081 ( .A(G125), .B(n1337), .ZN(n1319) );
XNOR2_X1 U1082 ( .A(n1195), .B(G131), .ZN(n1337) );
INV_X1 U1083 ( .A(G146), .ZN(n1195) );
NAND2_X1 U1084 ( .A1(KEYINPUT11), .A2(n1284), .ZN(n1224) );
INV_X1 U1085 ( .A(G110), .ZN(n1284) );
endmodule


