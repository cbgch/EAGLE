//Key = 1111001100101110111000110100011100100101100101011111101101000001


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
n1307, n1308;

XOR2_X1 U722 ( .A(G107), .B(n997), .Z(G9) );
NOR4_X1 U723 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(n997) );
XNOR2_X1 U724 ( .A(KEYINPUT38), .B(n1002), .ZN(n1001) );
NAND2_X1 U725 ( .A1(n1003), .A2(n1004), .ZN(n999) );
NOR2_X1 U726 ( .A1(n1005), .A2(n1006), .ZN(G75) );
NOR4_X1 U727 ( .A1(G953), .A2(n1007), .A3(n1008), .A4(n1009), .ZN(n1006) );
INV_X1 U728 ( .A(n1010), .ZN(n1009) );
NOR2_X1 U729 ( .A1(n1011), .A2(n1012), .ZN(n1008) );
NOR2_X1 U730 ( .A1(n1013), .A2(n1014), .ZN(n1011) );
NOR3_X1 U731 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n1014) );
NOR2_X1 U732 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U733 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
NOR2_X1 U734 ( .A1(n1022), .A2(n1023), .ZN(n1020) );
NOR2_X1 U735 ( .A1(n1024), .A2(n1025), .ZN(n1023) );
NOR2_X1 U736 ( .A1(n1026), .A2(n1027), .ZN(n1024) );
NOR2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR3_X1 U738 ( .A1(n1030), .A2(n1031), .A3(n1032), .ZN(n1022) );
NOR2_X1 U739 ( .A1(n1033), .A2(n1031), .ZN(n1018) );
NOR2_X1 U740 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
NOR2_X1 U741 ( .A1(n1025), .A2(n1036), .ZN(n1034) );
NOR3_X1 U742 ( .A1(n1037), .A2(n1021), .A3(n1025), .ZN(n1013) );
NAND3_X1 U743 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1037) );
NAND2_X1 U744 ( .A1(n1017), .A2(n1015), .ZN(n1039) );
NAND2_X1 U745 ( .A1(n1041), .A2(n1003), .ZN(n1038) );
NOR3_X1 U746 ( .A1(n1007), .A2(G953), .A3(G952), .ZN(n1005) );
AND4_X1 U747 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n1007) );
NOR4_X1 U748 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1045) );
XOR2_X1 U749 ( .A(n1050), .B(n1051), .Z(n1048) );
NOR2_X1 U750 ( .A1(n1052), .A2(KEYINPUT20), .ZN(n1051) );
XNOR2_X1 U751 ( .A(n1053), .B(n1054), .ZN(n1047) );
NAND2_X1 U752 ( .A1(KEYINPUT22), .A2(n1055), .ZN(n1053) );
XOR2_X1 U753 ( .A(KEYINPUT29), .B(n1056), .Z(n1055) );
XOR2_X1 U754 ( .A(n1057), .B(n1058), .Z(n1044) );
XOR2_X1 U755 ( .A(n1059), .B(n1060), .Z(G72) );
NOR2_X1 U756 ( .A1(n1061), .A2(n1062), .ZN(n1060) );
AND2_X1 U757 ( .A1(G227), .A2(G900), .ZN(n1061) );
NAND2_X1 U758 ( .A1(n1063), .A2(n1064), .ZN(n1059) );
NAND2_X1 U759 ( .A1(n1065), .A2(n1062), .ZN(n1064) );
XNOR2_X1 U760 ( .A(n1066), .B(n1067), .ZN(n1065) );
NOR2_X1 U761 ( .A1(n1068), .A2(n1069), .ZN(n1067) );
XOR2_X1 U762 ( .A(n1070), .B(KEYINPUT8), .Z(n1068) );
NAND3_X1 U763 ( .A1(G900), .A2(n1066), .A3(G953), .ZN(n1063) );
XNOR2_X1 U764 ( .A(n1071), .B(n1072), .ZN(n1066) );
XNOR2_X1 U765 ( .A(n1073), .B(n1074), .ZN(n1072) );
XOR2_X1 U766 ( .A(n1075), .B(n1076), .Z(n1074) );
NOR2_X1 U767 ( .A1(n1077), .A2(n1078), .ZN(n1076) );
XOR2_X1 U768 ( .A(KEYINPUT26), .B(n1079), .Z(n1078) );
NOR2_X1 U769 ( .A1(G125), .A2(n1080), .ZN(n1079) );
NOR2_X1 U770 ( .A1(G140), .A2(n1081), .ZN(n1077) );
INV_X1 U771 ( .A(G125), .ZN(n1081) );
NAND2_X1 U772 ( .A1(KEYINPUT30), .A2(n1082), .ZN(n1075) );
XOR2_X1 U773 ( .A(n1083), .B(n1084), .Z(n1071) );
XNOR2_X1 U774 ( .A(n1085), .B(G134), .ZN(n1084) );
XNOR2_X1 U775 ( .A(KEYINPUT59), .B(KEYINPUT28), .ZN(n1083) );
XOR2_X1 U776 ( .A(n1086), .B(n1087), .Z(G69) );
XOR2_X1 U777 ( .A(n1088), .B(n1089), .Z(n1087) );
NOR2_X1 U778 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
XNOR2_X1 U779 ( .A(n1092), .B(n1093), .ZN(n1091) );
NAND3_X1 U780 ( .A1(n1094), .A2(n1095), .A3(n1096), .ZN(n1092) );
NAND2_X1 U781 ( .A1(KEYINPUT19), .A2(n1097), .ZN(n1096) );
OR3_X1 U782 ( .A1(n1098), .A2(KEYINPUT19), .A3(n1099), .ZN(n1095) );
NAND2_X1 U783 ( .A1(n1099), .A2(n1098), .ZN(n1094) );
NAND2_X1 U784 ( .A1(KEYINPUT43), .A2(n1100), .ZN(n1098) );
NOR2_X1 U785 ( .A1(G898), .A2(n1062), .ZN(n1090) );
NAND2_X1 U786 ( .A1(n1062), .A2(n1101), .ZN(n1088) );
NAND2_X1 U787 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
INV_X1 U788 ( .A(n1104), .ZN(n1103) );
XNOR2_X1 U789 ( .A(n1105), .B(KEYINPUT61), .ZN(n1102) );
NAND2_X1 U790 ( .A1(G953), .A2(n1106), .ZN(n1086) );
NAND2_X1 U791 ( .A1(G898), .A2(G224), .ZN(n1106) );
NOR2_X1 U792 ( .A1(n1107), .A2(n1108), .ZN(G66) );
XOR2_X1 U793 ( .A(n1109), .B(n1110), .Z(n1108) );
NOR2_X1 U794 ( .A1(n1058), .A2(n1111), .ZN(n1110) );
NOR2_X1 U795 ( .A1(n1107), .A2(n1112), .ZN(G63) );
NOR3_X1 U796 ( .A1(n1056), .A2(n1113), .A3(n1114), .ZN(n1112) );
AND3_X1 U797 ( .A1(n1115), .A2(G478), .A3(n1116), .ZN(n1114) );
NOR2_X1 U798 ( .A1(n1117), .A2(n1115), .ZN(n1113) );
NOR2_X1 U799 ( .A1(n1010), .A2(n1054), .ZN(n1117) );
INV_X1 U800 ( .A(G478), .ZN(n1054) );
NOR2_X1 U801 ( .A1(n1107), .A2(n1118), .ZN(G60) );
NOR2_X1 U802 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
XOR2_X1 U803 ( .A(n1121), .B(KEYINPUT18), .Z(n1120) );
NAND2_X1 U804 ( .A1(n1122), .A2(n1123), .ZN(n1121) );
NOR2_X1 U805 ( .A1(n1122), .A2(n1123), .ZN(n1119) );
AND2_X1 U806 ( .A1(n1116), .A2(G475), .ZN(n1122) );
XOR2_X1 U807 ( .A(G104), .B(n1124), .Z(G6) );
NOR2_X1 U808 ( .A1(n1107), .A2(n1125), .ZN(G57) );
XOR2_X1 U809 ( .A(n1126), .B(n1127), .Z(n1125) );
XNOR2_X1 U810 ( .A(n1128), .B(KEYINPUT36), .ZN(n1127) );
NAND2_X1 U811 ( .A1(KEYINPUT13), .A2(n1129), .ZN(n1128) );
XNOR2_X1 U812 ( .A(n1100), .B(n1130), .ZN(n1129) );
XOR2_X1 U813 ( .A(n1131), .B(n1132), .Z(n1130) );
AND2_X1 U814 ( .A1(G472), .A2(n1116), .ZN(n1132) );
NAND2_X1 U815 ( .A1(KEYINPUT57), .A2(n1133), .ZN(n1131) );
NOR2_X1 U816 ( .A1(n1134), .A2(n1135), .ZN(G54) );
XOR2_X1 U817 ( .A(KEYINPUT5), .B(n1107), .Z(n1135) );
XOR2_X1 U818 ( .A(n1136), .B(n1137), .Z(n1134) );
AND2_X1 U819 ( .A1(G469), .A2(n1116), .ZN(n1137) );
NAND2_X1 U820 ( .A1(n1138), .A2(KEYINPUT63), .ZN(n1136) );
XOR2_X1 U821 ( .A(n1139), .B(n1140), .Z(n1138) );
XNOR2_X1 U822 ( .A(G110), .B(n1141), .ZN(n1140) );
NOR2_X1 U823 ( .A1(n1107), .A2(n1142), .ZN(G51) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(n1142) );
XNOR2_X1 U825 ( .A(n1145), .B(n1146), .ZN(n1144) );
XNOR2_X1 U826 ( .A(n1147), .B(n1148), .ZN(n1143) );
NOR2_X1 U827 ( .A1(n1149), .A2(n1111), .ZN(n1147) );
INV_X1 U828 ( .A(n1116), .ZN(n1111) );
NOR2_X1 U829 ( .A1(n1150), .A2(n1010), .ZN(n1116) );
NOR4_X1 U830 ( .A1(n1070), .A2(n1104), .A3(n1069), .A4(n1105), .ZN(n1010) );
NAND4_X1 U831 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1069) );
NAND4_X1 U832 ( .A1(n1155), .A2(n1156), .A3(n1017), .A4(n1036), .ZN(n1151) );
NAND4_X1 U833 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1104) );
NOR3_X1 U834 ( .A1(n1161), .A2(n1162), .A3(n1163), .ZN(n1160) );
NOR3_X1 U835 ( .A1(n998), .A2(n1164), .A3(n1017), .ZN(n1161) );
NOR2_X1 U836 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
AND2_X1 U837 ( .A1(n1004), .A2(n1167), .ZN(n1166) );
NOR4_X1 U838 ( .A1(KEYINPUT10), .A2(n1027), .A3(n1168), .A4(n1169), .ZN(n1165) );
NAND2_X1 U839 ( .A1(KEYINPUT10), .A2(n1124), .ZN(n1159) );
NOR4_X1 U840 ( .A1(n1169), .A2(n1170), .A3(n1017), .A4(n998), .ZN(n1124) );
NAND3_X1 U841 ( .A1(n1171), .A2(n1043), .A3(n1172), .ZN(n1158) );
OR2_X1 U842 ( .A1(n1173), .A2(n1041), .ZN(n1157) );
NOR2_X1 U843 ( .A1(n1156), .A2(n1004), .ZN(n1041) );
NAND4_X1 U844 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1070) );
NAND4_X1 U845 ( .A1(n1172), .A2(n1178), .A3(n1027), .A4(n1004), .ZN(n1174) );
XNOR2_X1 U846 ( .A(n1052), .B(KEYINPUT9), .ZN(n1149) );
INV_X1 U847 ( .A(n1179), .ZN(n1052) );
AND2_X1 U848 ( .A1(n1180), .A2(G953), .ZN(n1107) );
XNOR2_X1 U849 ( .A(G952), .B(KEYINPUT24), .ZN(n1180) );
NAND2_X1 U850 ( .A1(n1181), .A2(n1182), .ZN(G48) );
NAND2_X1 U851 ( .A1(G146), .A2(n1152), .ZN(n1182) );
XOR2_X1 U852 ( .A(KEYINPUT48), .B(n1183), .Z(n1181) );
NOR2_X1 U853 ( .A1(G146), .A2(n1152), .ZN(n1183) );
NAND4_X1 U854 ( .A1(n1172), .A2(n1178), .A3(n1156), .A4(n1027), .ZN(n1152) );
XNOR2_X1 U855 ( .A(G143), .B(n1153), .ZN(G45) );
NAND3_X1 U856 ( .A1(n1178), .A2(n1184), .A3(n1185), .ZN(n1153) );
NOR3_X1 U857 ( .A1(n1000), .A2(n1042), .A3(n1186), .ZN(n1185) );
XNOR2_X1 U858 ( .A(n1080), .B(n1187), .ZN(G42) );
NOR4_X1 U859 ( .A1(n998), .A2(n1188), .A3(n1169), .A4(n1031), .ZN(n1187) );
INV_X1 U860 ( .A(n1040), .ZN(n1031) );
NAND2_X1 U861 ( .A1(n1189), .A2(n1017), .ZN(n1188) );
XNOR2_X1 U862 ( .A(KEYINPUT6), .B(n1190), .ZN(n1189) );
XNOR2_X1 U863 ( .A(G137), .B(n1154), .ZN(G39) );
NAND3_X1 U864 ( .A1(n1155), .A2(n1191), .A3(n1172), .ZN(n1154) );
INV_X1 U865 ( .A(n1015), .ZN(n1191) );
XNOR2_X1 U866 ( .A(G134), .B(n1175), .ZN(G36) );
NAND3_X1 U867 ( .A1(n1184), .A2(n1004), .A3(n1155), .ZN(n1175) );
XNOR2_X1 U868 ( .A(G131), .B(n1176), .ZN(G33) );
NAND3_X1 U869 ( .A1(n1156), .A2(n1184), .A3(n1155), .ZN(n1176) );
AND2_X1 U870 ( .A1(n1178), .A2(n1040), .ZN(n1155) );
NOR2_X1 U871 ( .A1(n1028), .A2(n1046), .ZN(n1040) );
XNOR2_X1 U872 ( .A(G128), .B(n1192), .ZN(G30) );
NAND2_X1 U873 ( .A1(n1193), .A2(n1027), .ZN(n1192) );
XOR2_X1 U874 ( .A(n1194), .B(KEYINPUT45), .Z(n1193) );
NAND3_X1 U875 ( .A1(n1004), .A2(n1195), .A3(n1178), .ZN(n1194) );
AND3_X1 U876 ( .A1(n1190), .A2(n1030), .A3(n1032), .ZN(n1178) );
XOR2_X1 U877 ( .A(KEYINPUT35), .B(n1172), .Z(n1195) );
NAND3_X1 U878 ( .A1(n1196), .A2(n1197), .A3(n1198), .ZN(G3) );
OR2_X1 U879 ( .A1(G101), .A2(KEYINPUT31), .ZN(n1198) );
NAND3_X1 U880 ( .A1(KEYINPUT31), .A2(G101), .A3(n1199), .ZN(n1197) );
NAND2_X1 U881 ( .A1(n1105), .A2(n1200), .ZN(n1196) );
NAND2_X1 U882 ( .A1(n1201), .A2(KEYINPUT31), .ZN(n1200) );
XNOR2_X1 U883 ( .A(G101), .B(KEYINPUT25), .ZN(n1201) );
INV_X1 U884 ( .A(n1199), .ZN(n1105) );
NAND4_X1 U885 ( .A1(n1184), .A2(n1171), .A3(n1032), .A4(n1030), .ZN(n1199) );
XNOR2_X1 U886 ( .A(G125), .B(n1177), .ZN(G27) );
NAND4_X1 U887 ( .A1(n1043), .A2(n1027), .A3(n1156), .A4(n1202), .ZN(n1177) );
AND3_X1 U888 ( .A1(n1017), .A2(n1190), .A3(n1036), .ZN(n1202) );
NAND2_X1 U889 ( .A1(n1012), .A2(n1203), .ZN(n1190) );
NAND4_X1 U890 ( .A1(G902), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(n1203) );
INV_X1 U891 ( .A(G900), .ZN(n1206) );
XNOR2_X1 U892 ( .A(KEYINPUT58), .B(n1062), .ZN(n1204) );
XOR2_X1 U893 ( .A(G122), .B(n1163), .Z(G24) );
AND4_X1 U894 ( .A1(n1003), .A2(n1043), .A3(n1167), .A4(n1207), .ZN(n1163) );
NOR3_X1 U895 ( .A1(n1186), .A2(n1021), .A3(n1042), .ZN(n1207) );
INV_X1 U896 ( .A(n1036), .ZN(n1021) );
XNOR2_X1 U897 ( .A(G119), .B(n1208), .ZN(G21) );
NAND4_X1 U898 ( .A1(KEYINPUT3), .A2(n1172), .A3(n1171), .A4(n1043), .ZN(n1208) );
NOR2_X1 U899 ( .A1(n1036), .A2(n1003), .ZN(n1172) );
INV_X1 U900 ( .A(n1017), .ZN(n1003) );
XNOR2_X1 U901 ( .A(G116), .B(n1209), .ZN(G18) );
NAND3_X1 U902 ( .A1(n1210), .A2(n1004), .A3(KEYINPUT23), .ZN(n1209) );
NOR2_X1 U903 ( .A1(n1211), .A2(n1186), .ZN(n1004) );
INV_X1 U904 ( .A(n1173), .ZN(n1210) );
XOR2_X1 U905 ( .A(G113), .B(n1212), .Z(G15) );
NOR2_X1 U906 ( .A1(n1213), .A2(n1173), .ZN(n1212) );
NAND3_X1 U907 ( .A1(n1167), .A2(n1043), .A3(n1184), .ZN(n1173) );
NOR2_X1 U908 ( .A1(n1036), .A2(n1017), .ZN(n1184) );
INV_X1 U909 ( .A(n1025), .ZN(n1043) );
NAND2_X1 U910 ( .A1(n1214), .A2(n1030), .ZN(n1025) );
INV_X1 U911 ( .A(n1032), .ZN(n1214) );
XNOR2_X1 U912 ( .A(n1156), .B(KEYINPUT27), .ZN(n1213) );
INV_X1 U913 ( .A(n1169), .ZN(n1156) );
NAND2_X1 U914 ( .A1(n1186), .A2(n1211), .ZN(n1169) );
XOR2_X1 U915 ( .A(G110), .B(n1162), .Z(G12) );
AND3_X1 U916 ( .A1(n1035), .A2(n1017), .A3(n1171), .ZN(n1162) );
NOR2_X1 U917 ( .A1(n1015), .A2(n1170), .ZN(n1171) );
INV_X1 U918 ( .A(n1167), .ZN(n1170) );
NOR2_X1 U919 ( .A1(n1000), .A2(n1168), .ZN(n1167) );
INV_X1 U920 ( .A(n1002), .ZN(n1168) );
NAND2_X1 U921 ( .A1(n1012), .A2(n1215), .ZN(n1002) );
NAND4_X1 U922 ( .A1(G902), .A2(G953), .A3(n1205), .A4(n1216), .ZN(n1215) );
INV_X1 U923 ( .A(G898), .ZN(n1216) );
NAND3_X1 U924 ( .A1(n1205), .A2(n1062), .A3(G952), .ZN(n1012) );
INV_X1 U925 ( .A(G953), .ZN(n1062) );
NAND2_X1 U926 ( .A1(G237), .A2(G234), .ZN(n1205) );
INV_X1 U927 ( .A(n1027), .ZN(n1000) );
NOR2_X1 U928 ( .A1(n1217), .A2(n1046), .ZN(n1027) );
INV_X1 U929 ( .A(n1029), .ZN(n1046) );
NAND2_X1 U930 ( .A1(G214), .A2(n1218), .ZN(n1029) );
INV_X1 U931 ( .A(n1028), .ZN(n1217) );
XOR2_X1 U932 ( .A(n1050), .B(n1179), .Z(n1028) );
NAND2_X1 U933 ( .A1(G210), .A2(n1218), .ZN(n1179) );
NAND2_X1 U934 ( .A1(n1219), .A2(n1150), .ZN(n1218) );
NAND2_X1 U935 ( .A1(n1220), .A2(n1150), .ZN(n1050) );
XNOR2_X1 U936 ( .A(n1145), .B(n1221), .ZN(n1220) );
NOR4_X1 U937 ( .A1(n1222), .A2(n1223), .A3(KEYINPUT62), .A4(n1224), .ZN(n1221) );
AND2_X1 U938 ( .A1(n1225), .A2(n1146), .ZN(n1224) );
NOR2_X1 U939 ( .A1(n1226), .A2(n1227), .ZN(n1223) );
NOR2_X1 U940 ( .A1(KEYINPUT32), .A2(n1146), .ZN(n1226) );
NOR4_X1 U941 ( .A1(n1148), .A2(n1225), .A3(KEYINPUT32), .A4(n1146), .ZN(n1222) );
XNOR2_X1 U942 ( .A(G125), .B(KEYINPUT14), .ZN(n1146) );
INV_X1 U943 ( .A(KEYINPUT49), .ZN(n1225) );
XNOR2_X1 U944 ( .A(n1228), .B(n1229), .ZN(n1145) );
XNOR2_X1 U945 ( .A(n1097), .B(n1093), .ZN(n1229) );
XNOR2_X1 U946 ( .A(n1230), .B(n1231), .ZN(n1093) );
XNOR2_X1 U947 ( .A(G110), .B(KEYINPUT50), .ZN(n1230) );
XNOR2_X1 U948 ( .A(n1099), .B(n1232), .ZN(n1228) );
AND2_X1 U949 ( .A1(n1233), .A2(G224), .ZN(n1232) );
AND2_X1 U950 ( .A1(n1234), .A2(n1235), .ZN(n1099) );
NAND2_X1 U951 ( .A1(G101), .A2(n1236), .ZN(n1235) );
XOR2_X1 U952 ( .A(KEYINPUT34), .B(n1237), .Z(n1234) );
NOR2_X1 U953 ( .A1(G101), .A2(n1236), .ZN(n1237) );
NAND2_X1 U954 ( .A1(n1186), .A2(n1042), .ZN(n1015) );
INV_X1 U955 ( .A(n1211), .ZN(n1042) );
XNOR2_X1 U956 ( .A(n1238), .B(G475), .ZN(n1211) );
OR2_X1 U957 ( .A1(n1123), .A2(G902), .ZN(n1238) );
XNOR2_X1 U958 ( .A(n1239), .B(n1240), .ZN(n1123) );
XOR2_X1 U959 ( .A(n1241), .B(n1242), .Z(n1240) );
XOR2_X1 U960 ( .A(n1243), .B(n1244), .Z(n1242) );
XOR2_X1 U961 ( .A(G104), .B(n1245), .Z(n1244) );
NOR2_X1 U962 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
INV_X1 U963 ( .A(G214), .ZN(n1246) );
XNOR2_X1 U964 ( .A(n1231), .B(n1248), .ZN(n1243) );
NOR2_X1 U965 ( .A1(G131), .A2(KEYINPUT33), .ZN(n1248) );
XOR2_X1 U966 ( .A(n1249), .B(n1250), .Z(n1241) );
XOR2_X1 U967 ( .A(KEYINPUT12), .B(G146), .Z(n1250) );
XNOR2_X1 U968 ( .A(G113), .B(G143), .ZN(n1249) );
XNOR2_X1 U969 ( .A(G478), .B(n1056), .ZN(n1186) );
NOR2_X1 U970 ( .A1(n1115), .A2(G902), .ZN(n1056) );
NAND3_X1 U971 ( .A1(n1251), .A2(n1252), .A3(n1253), .ZN(n1115) );
NAND2_X1 U972 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U973 ( .A(KEYINPUT1), .ZN(n1255) );
NAND3_X1 U974 ( .A1(KEYINPUT1), .A2(n1256), .A3(n1257), .ZN(n1252) );
OR2_X1 U975 ( .A1(n1257), .A2(n1256), .ZN(n1251) );
NOR2_X1 U976 ( .A1(n1258), .A2(n1254), .ZN(n1256) );
NAND3_X1 U977 ( .A1(n1259), .A2(n1233), .A3(G217), .ZN(n1254) );
INV_X1 U978 ( .A(KEYINPUT17), .ZN(n1258) );
XNOR2_X1 U979 ( .A(n1260), .B(n1261), .ZN(n1257) );
XNOR2_X1 U980 ( .A(n1262), .B(G134), .ZN(n1261) );
INV_X1 U981 ( .A(G143), .ZN(n1262) );
XNOR2_X1 U982 ( .A(n1263), .B(n1264), .ZN(n1260) );
NOR2_X1 U983 ( .A1(KEYINPUT53), .A2(n1265), .ZN(n1264) );
XNOR2_X1 U984 ( .A(n1231), .B(n1266), .ZN(n1265) );
XOR2_X1 U985 ( .A(G107), .B(n1267), .Z(n1266) );
NOR2_X1 U986 ( .A1(G116), .A2(KEYINPUT4), .ZN(n1267) );
XOR2_X1 U987 ( .A(G122), .B(KEYINPUT41), .Z(n1231) );
XOR2_X1 U988 ( .A(n1268), .B(n1058), .Z(n1017) );
NAND2_X1 U989 ( .A1(G217), .A2(n1269), .ZN(n1058) );
NAND2_X1 U990 ( .A1(KEYINPUT39), .A2(n1057), .ZN(n1268) );
NOR2_X1 U991 ( .A1(n1109), .A2(G902), .ZN(n1057) );
XOR2_X1 U992 ( .A(n1270), .B(n1271), .Z(n1109) );
XNOR2_X1 U993 ( .A(n1272), .B(n1273), .ZN(n1271) );
XNOR2_X1 U994 ( .A(n1274), .B(n1275), .ZN(n1273) );
NOR2_X1 U995 ( .A1(KEYINPUT11), .A2(n1239), .ZN(n1275) );
XOR2_X1 U996 ( .A(G125), .B(n1276), .Z(n1239) );
XNOR2_X1 U997 ( .A(KEYINPUT21), .B(n1080), .ZN(n1276) );
INV_X1 U998 ( .A(G140), .ZN(n1080) );
NOR2_X1 U999 ( .A1(KEYINPUT44), .A2(n1277), .ZN(n1274) );
XNOR2_X1 U1000 ( .A(G137), .B(n1278), .ZN(n1277) );
NAND3_X1 U1001 ( .A1(G221), .A2(n1233), .A3(n1259), .ZN(n1278) );
XNOR2_X1 U1002 ( .A(G234), .B(KEYINPUT37), .ZN(n1259) );
XNOR2_X1 U1003 ( .A(G110), .B(n1279), .ZN(n1270) );
XOR2_X1 U1004 ( .A(KEYINPUT12), .B(G119), .Z(n1279) );
INV_X1 U1005 ( .A(n998), .ZN(n1035) );
NAND3_X1 U1006 ( .A1(n1036), .A2(n1030), .A3(n1032), .ZN(n998) );
XNOR2_X1 U1007 ( .A(n1280), .B(G469), .ZN(n1032) );
NAND2_X1 U1008 ( .A1(n1281), .A2(n1150), .ZN(n1280) );
XOR2_X1 U1009 ( .A(n1282), .B(n1139), .Z(n1281) );
XOR2_X1 U1010 ( .A(n1283), .B(n1284), .Z(n1139) );
XNOR2_X1 U1011 ( .A(n1285), .B(G140), .ZN(n1284) );
NAND2_X1 U1012 ( .A1(G227), .A2(n1233), .ZN(n1285) );
XNOR2_X1 U1013 ( .A(n1286), .B(n1073), .ZN(n1283) );
XOR2_X1 U1014 ( .A(n1227), .B(KEYINPUT15), .Z(n1073) );
XNOR2_X1 U1015 ( .A(n1287), .B(n1288), .ZN(n1282) );
NAND2_X1 U1016 ( .A1(KEYINPUT16), .A2(G110), .ZN(n1288) );
NAND2_X1 U1017 ( .A1(KEYINPUT52), .A2(n1141), .ZN(n1287) );
XOR2_X1 U1018 ( .A(n1289), .B(n1290), .Z(n1141) );
NOR2_X1 U1019 ( .A1(KEYINPUT42), .A2(n1291), .ZN(n1290) );
INV_X1 U1020 ( .A(n1236), .ZN(n1291) );
XOR2_X1 U1021 ( .A(G104), .B(G107), .Z(n1236) );
XNOR2_X1 U1022 ( .A(G101), .B(KEYINPUT60), .ZN(n1289) );
NAND2_X1 U1023 ( .A1(G221), .A2(n1269), .ZN(n1030) );
NAND2_X1 U1024 ( .A1(G234), .A2(n1150), .ZN(n1269) );
XOR2_X1 U1025 ( .A(n1049), .B(KEYINPUT0), .Z(n1036) );
XNOR2_X1 U1026 ( .A(n1292), .B(G472), .ZN(n1049) );
NAND2_X1 U1027 ( .A1(n1293), .A2(n1150), .ZN(n1292) );
INV_X1 U1028 ( .A(G902), .ZN(n1150) );
XNOR2_X1 U1029 ( .A(n1294), .B(n1097), .ZN(n1293) );
INV_X1 U1030 ( .A(n1100), .ZN(n1097) );
XNOR2_X1 U1031 ( .A(n1295), .B(n1296), .ZN(n1100) );
XOR2_X1 U1032 ( .A(KEYINPUT56), .B(G119), .Z(n1296) );
XNOR2_X1 U1033 ( .A(G113), .B(G116), .ZN(n1295) );
XOR2_X1 U1034 ( .A(n1297), .B(n1133), .Z(n1294) );
XNOR2_X1 U1035 ( .A(n1148), .B(n1286), .ZN(n1133) );
XNOR2_X1 U1036 ( .A(n1298), .B(n1082), .ZN(n1286) );
XOR2_X1 U1037 ( .A(G131), .B(KEYINPUT47), .Z(n1082) );
NAND3_X1 U1038 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1298) );
OR2_X1 U1039 ( .A1(n1302), .A2(KEYINPUT40), .ZN(n1301) );
NAND3_X1 U1040 ( .A1(KEYINPUT40), .A2(n1302), .A3(n1085), .ZN(n1300) );
INV_X1 U1041 ( .A(G137), .ZN(n1085) );
NAND2_X1 U1042 ( .A1(G137), .A2(n1303), .ZN(n1299) );
NAND2_X1 U1043 ( .A1(KEYINPUT40), .A2(n1304), .ZN(n1303) );
XNOR2_X1 U1044 ( .A(KEYINPUT55), .B(n1302), .ZN(n1304) );
XNOR2_X1 U1045 ( .A(G134), .B(KEYINPUT54), .ZN(n1302) );
INV_X1 U1046 ( .A(n1227), .ZN(n1148) );
XNOR2_X1 U1047 ( .A(n1305), .B(n1272), .ZN(n1227) );
XNOR2_X1 U1048 ( .A(G146), .B(n1306), .ZN(n1272) );
INV_X1 U1049 ( .A(n1263), .ZN(n1306) );
XOR2_X1 U1050 ( .A(G128), .B(KEYINPUT7), .Z(n1263) );
XNOR2_X1 U1051 ( .A(G143), .B(KEYINPUT46), .ZN(n1305) );
NAND2_X1 U1052 ( .A1(KEYINPUT2), .A2(n1126), .ZN(n1297) );
XOR2_X1 U1053 ( .A(G101), .B(n1307), .Z(n1126) );
NOR2_X1 U1054 ( .A1(n1308), .A2(n1247), .ZN(n1307) );
NAND2_X1 U1055 ( .A1(n1233), .A2(n1219), .ZN(n1247) );
INV_X1 U1056 ( .A(G237), .ZN(n1219) );
XOR2_X1 U1057 ( .A(G953), .B(KEYINPUT51), .Z(n1233) );
INV_X1 U1058 ( .A(G210), .ZN(n1308) );
endmodule


