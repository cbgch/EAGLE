//Key = 1001100000010100111110001000001011111101011111010110010001100100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345;

XOR2_X1 U743 ( .A(n1020), .B(n1021), .Z(G9) );
NOR2_X1 U744 ( .A1(n1022), .A2(n1023), .ZN(G75) );
NOR4_X1 U745 ( .A1(n1024), .A2(n1025), .A3(n1026), .A4(n1027), .ZN(n1023) );
NOR2_X1 U746 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
XOR2_X1 U747 ( .A(KEYINPUT0), .B(n1030), .Z(n1025) );
NOR2_X1 U748 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
NOR2_X1 U749 ( .A1(n1033), .A2(n1029), .ZN(n1032) );
NAND3_X1 U750 ( .A1(n1034), .A2(n1035), .A3(n1036), .ZN(n1029) );
INV_X1 U751 ( .A(n1037), .ZN(n1033) );
NOR3_X1 U752 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1031) );
INV_X1 U753 ( .A(n1041), .ZN(n1040) );
NOR2_X1 U754 ( .A1(n1042), .A2(n1043), .ZN(n1039) );
NOR2_X1 U755 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
NOR2_X1 U756 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
NOR2_X1 U757 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
NOR4_X1 U758 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1046) );
NOR3_X1 U759 ( .A1(n1054), .A2(n1055), .A3(n1056), .ZN(n1042) );
NAND3_X1 U760 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1024) );
NAND3_X1 U761 ( .A1(n1041), .A2(n1060), .A3(n1036), .ZN(n1059) );
INV_X1 U762 ( .A(n1038), .ZN(n1036) );
NAND3_X1 U763 ( .A1(n1061), .A2(n1062), .A3(n1063), .ZN(n1060) );
NAND2_X1 U764 ( .A1(n1034), .A2(n1064), .ZN(n1063) );
INV_X1 U765 ( .A(n1055), .ZN(n1034) );
NAND2_X1 U766 ( .A1(n1065), .A2(n1066), .ZN(n1055) );
NAND3_X1 U767 ( .A1(n1065), .A2(n1067), .A3(n1068), .ZN(n1062) );
XOR2_X1 U768 ( .A(KEYINPUT12), .B(n1035), .Z(n1067) );
NAND3_X1 U769 ( .A1(n1066), .A2(n1069), .A3(n1035), .ZN(n1061) );
INV_X1 U770 ( .A(n1045), .ZN(n1035) );
NOR3_X1 U771 ( .A1(n1070), .A2(G953), .A3(G952), .ZN(n1022) );
INV_X1 U772 ( .A(n1057), .ZN(n1070) );
NAND4_X1 U773 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1057) );
NOR3_X1 U774 ( .A1(n1048), .A2(n1045), .A3(n1075), .ZN(n1074) );
INV_X1 U775 ( .A(n1065), .ZN(n1048) );
XOR2_X1 U776 ( .A(G475), .B(n1076), .Z(n1072) );
NOR2_X1 U777 ( .A1(n1077), .A2(KEYINPUT40), .ZN(n1076) );
XOR2_X1 U778 ( .A(n1078), .B(n1079), .Z(G72) );
NOR2_X1 U779 ( .A1(n1080), .A2(n1058), .ZN(n1079) );
NOR2_X1 U780 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
NAND2_X1 U781 ( .A1(n1083), .A2(n1084), .ZN(n1078) );
NAND2_X1 U782 ( .A1(n1085), .A2(n1058), .ZN(n1084) );
XOR2_X1 U783 ( .A(n1086), .B(n1087), .Z(n1085) );
XNOR2_X1 U784 ( .A(n1088), .B(KEYINPUT53), .ZN(n1087) );
NAND3_X1 U785 ( .A1(n1089), .A2(n1090), .A3(n1091), .ZN(n1086) );
NOR3_X1 U786 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NAND3_X1 U787 ( .A1(n1088), .A2(G900), .A3(G953), .ZN(n1083) );
NOR2_X1 U788 ( .A1(KEYINPUT25), .A2(n1095), .ZN(n1088) );
XOR2_X1 U789 ( .A(n1096), .B(n1097), .Z(n1095) );
XNOR2_X1 U790 ( .A(n1098), .B(n1099), .ZN(n1097) );
NAND2_X1 U791 ( .A1(n1100), .A2(n1101), .ZN(n1098) );
NAND2_X1 U792 ( .A1(n1102), .A2(n1103), .ZN(n1101) );
XOR2_X1 U793 ( .A(n1104), .B(KEYINPUT56), .Z(n1100) );
NAND2_X1 U794 ( .A1(n1105), .A2(n1106), .ZN(n1104) );
XOR2_X1 U795 ( .A(KEYINPUT51), .B(KEYINPUT18), .Z(n1096) );
XOR2_X1 U796 ( .A(n1107), .B(n1108), .Z(G69) );
NOR3_X1 U797 ( .A1(n1058), .A2(KEYINPUT5), .A3(n1109), .ZN(n1108) );
NOR2_X1 U798 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
NAND2_X1 U799 ( .A1(n1112), .A2(n1113), .ZN(n1107) );
NAND2_X1 U800 ( .A1(n1114), .A2(n1058), .ZN(n1113) );
XNOR2_X1 U801 ( .A(n1115), .B(n1116), .ZN(n1114) );
NAND3_X1 U802 ( .A1(n1116), .A2(G898), .A3(G953), .ZN(n1112) );
NOR2_X1 U803 ( .A1(KEYINPUT22), .A2(n1117), .ZN(n1116) );
XOR2_X1 U804 ( .A(n1118), .B(n1119), .Z(n1117) );
INV_X1 U805 ( .A(n1120), .ZN(n1119) );
XNOR2_X1 U806 ( .A(n1121), .B(KEYINPUT13), .ZN(n1118) );
NOR2_X1 U807 ( .A1(n1122), .A2(n1123), .ZN(G66) );
NOR2_X1 U808 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
XOR2_X1 U809 ( .A(n1126), .B(n1127), .Z(n1125) );
NOR2_X1 U810 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
NAND2_X1 U811 ( .A1(KEYINPUT16), .A2(n1130), .ZN(n1126) );
NOR2_X1 U812 ( .A1(KEYINPUT16), .A2(n1130), .ZN(n1124) );
NOR2_X1 U813 ( .A1(n1122), .A2(n1131), .ZN(G63) );
NOR2_X1 U814 ( .A1(n1132), .A2(n1133), .ZN(n1131) );
XOR2_X1 U815 ( .A(n1134), .B(n1135), .Z(n1133) );
NOR2_X1 U816 ( .A1(KEYINPUT1), .A2(n1136), .ZN(n1135) );
AND2_X1 U817 ( .A1(G478), .A2(n1137), .ZN(n1134) );
AND2_X1 U818 ( .A1(n1136), .A2(KEYINPUT1), .ZN(n1132) );
NOR2_X1 U819 ( .A1(n1122), .A2(n1138), .ZN(G60) );
NOR3_X1 U820 ( .A1(n1077), .A2(n1139), .A3(n1140), .ZN(n1138) );
NOR2_X1 U821 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
AND3_X1 U822 ( .A1(KEYINPUT34), .A2(n1027), .A3(G475), .ZN(n1141) );
AND4_X1 U823 ( .A1(n1142), .A2(KEYINPUT34), .A3(G475), .A4(n1137), .ZN(n1139) );
XOR2_X1 U824 ( .A(n1143), .B(n1144), .Z(G6) );
NOR2_X1 U825 ( .A1(n1145), .A2(KEYINPUT31), .ZN(n1144) );
NOR2_X1 U826 ( .A1(n1122), .A2(n1146), .ZN(G57) );
XOR2_X1 U827 ( .A(n1147), .B(n1148), .Z(n1146) );
XOR2_X1 U828 ( .A(n1149), .B(n1150), .Z(n1148) );
AND2_X1 U829 ( .A1(G472), .A2(n1137), .ZN(n1149) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1147) );
XOR2_X1 U831 ( .A(n1153), .B(n1154), .Z(n1152) );
NAND2_X1 U832 ( .A1(n1155), .A2(KEYINPUT20), .ZN(n1154) );
XOR2_X1 U833 ( .A(n1120), .B(KEYINPUT39), .Z(n1155) );
INV_X1 U834 ( .A(G101), .ZN(n1153) );
NOR2_X1 U835 ( .A1(KEYINPUT28), .A2(n1156), .ZN(n1151) );
NOR2_X1 U836 ( .A1(n1122), .A2(n1157), .ZN(G54) );
XOR2_X1 U837 ( .A(n1158), .B(n1159), .Z(n1157) );
XOR2_X1 U838 ( .A(n1160), .B(n1161), .Z(n1159) );
XOR2_X1 U839 ( .A(n1162), .B(n1163), .Z(n1161) );
NAND3_X1 U840 ( .A1(n1137), .A2(G469), .A3(KEYINPUT17), .ZN(n1163) );
INV_X1 U841 ( .A(n1129), .ZN(n1137) );
XOR2_X1 U842 ( .A(KEYINPUT27), .B(n1164), .Z(n1160) );
XOR2_X1 U843 ( .A(n1165), .B(n1166), .Z(n1158) );
XOR2_X1 U844 ( .A(n1102), .B(n1103), .Z(n1166) );
XOR2_X1 U845 ( .A(n1167), .B(n1168), .Z(n1165) );
NAND2_X1 U846 ( .A1(KEYINPUT37), .A2(n1169), .ZN(n1167) );
NOR2_X1 U847 ( .A1(n1122), .A2(n1170), .ZN(G51) );
XOR2_X1 U848 ( .A(n1171), .B(n1172), .Z(n1170) );
XOR2_X1 U849 ( .A(n1173), .B(n1174), .Z(n1172) );
XOR2_X1 U850 ( .A(n1175), .B(n1176), .Z(n1171) );
NOR2_X1 U851 ( .A1(n1177), .A2(n1129), .ZN(n1176) );
NAND2_X1 U852 ( .A1(G902), .A2(n1027), .ZN(n1129) );
NAND3_X1 U853 ( .A1(n1089), .A2(n1178), .A3(n1115), .ZN(n1027) );
AND4_X1 U854 ( .A1(n1179), .A2(n1021), .A3(n1180), .A4(n1181), .ZN(n1115) );
NOR4_X1 U855 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1145), .ZN(n1181) );
AND4_X1 U856 ( .A1(n1064), .A2(n1185), .A3(n1069), .A4(n1186), .ZN(n1145) );
NOR2_X1 U857 ( .A1(n1052), .A2(n1028), .ZN(n1186) );
NOR2_X1 U858 ( .A1(n1187), .A2(n1188), .ZN(n1180) );
NOR2_X1 U859 ( .A1(n1189), .A2(n1190), .ZN(n1188) );
XOR2_X1 U860 ( .A(KEYINPUT35), .B(n1191), .Z(n1190) );
NOR2_X1 U861 ( .A1(n1192), .A2(n1193), .ZN(n1191) );
XOR2_X1 U862 ( .A(n1049), .B(KEYINPUT9), .Z(n1192) );
NAND3_X1 U863 ( .A1(n1194), .A2(n1185), .A3(n1066), .ZN(n1021) );
XOR2_X1 U864 ( .A(KEYINPUT38), .B(n1195), .Z(n1178) );
NOR4_X1 U865 ( .A1(n1093), .A2(n1094), .A3(n1092), .A4(n1196), .ZN(n1195) );
XOR2_X1 U866 ( .A(n1090), .B(KEYINPUT32), .Z(n1196) );
NAND2_X1 U867 ( .A1(n1064), .A2(n1197), .ZN(n1090) );
XOR2_X1 U868 ( .A(KEYINPUT23), .B(n1198), .Z(n1197) );
AND4_X1 U869 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1089) );
NAND3_X1 U870 ( .A1(n1194), .A2(n1203), .A3(n1204), .ZN(n1199) );
XOR2_X1 U871 ( .A(n1205), .B(KEYINPUT11), .Z(n1204) );
NOR2_X1 U872 ( .A1(n1058), .A2(G952), .ZN(n1122) );
XOR2_X1 U873 ( .A(n1206), .B(G146), .Z(G48) );
NAND2_X1 U874 ( .A1(KEYINPUT33), .A2(n1207), .ZN(n1206) );
NAND2_X1 U875 ( .A1(n1198), .A2(n1064), .ZN(n1207) );
NOR3_X1 U876 ( .A1(n1205), .A2(n1028), .A3(n1208), .ZN(n1198) );
XOR2_X1 U877 ( .A(G143), .B(n1094), .Z(G45) );
AND4_X1 U878 ( .A1(n1075), .A2(n1209), .A3(n1064), .A4(n1210), .ZN(n1094) );
NOR2_X1 U879 ( .A1(n1211), .A2(n1208), .ZN(n1210) );
XOR2_X1 U880 ( .A(G140), .B(n1093), .Z(G42) );
AND3_X1 U881 ( .A1(n1212), .A2(n1213), .A3(n1214), .ZN(n1093) );
INV_X1 U882 ( .A(n1049), .ZN(n1212) );
XOR2_X1 U883 ( .A(G137), .B(n1092), .Z(G39) );
AND3_X1 U884 ( .A1(n1215), .A2(n1041), .A3(n1214), .ZN(n1092) );
XOR2_X1 U885 ( .A(n1200), .B(n1216), .Z(G36) );
NAND2_X1 U886 ( .A1(KEYINPUT58), .A2(G134), .ZN(n1216) );
NAND3_X1 U887 ( .A1(n1068), .A2(n1037), .A3(n1214), .ZN(n1200) );
XNOR2_X1 U888 ( .A(G131), .B(n1201), .ZN(G33) );
NAND3_X1 U889 ( .A1(n1213), .A2(n1068), .A3(n1214), .ZN(n1201) );
NOR2_X1 U890 ( .A1(n1208), .A2(n1045), .ZN(n1214) );
NAND2_X1 U891 ( .A1(n1217), .A2(n1054), .ZN(n1045) );
NAND2_X1 U892 ( .A1(n1069), .A2(n1203), .ZN(n1208) );
XOR2_X1 U893 ( .A(G128), .B(n1218), .Z(G30) );
AND3_X1 U894 ( .A1(n1215), .A2(n1203), .A3(n1194), .ZN(n1218) );
AND3_X1 U895 ( .A1(n1064), .A2(n1037), .A3(n1069), .ZN(n1194) );
XOR2_X1 U896 ( .A(G101), .B(n1184), .Z(G3) );
NOR3_X1 U897 ( .A1(n1211), .A2(n1189), .A3(n1193), .ZN(n1184) );
XOR2_X1 U898 ( .A(n1219), .B(n1202), .Z(G27) );
NAND4_X1 U899 ( .A1(n1064), .A2(n1203), .A3(n1065), .A4(n1220), .ZN(n1202) );
NOR2_X1 U900 ( .A1(n1028), .A2(n1049), .ZN(n1220) );
NAND2_X1 U901 ( .A1(n1038), .A2(n1221), .ZN(n1203) );
NAND4_X1 U902 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1082), .ZN(n1221) );
INV_X1 U903 ( .A(G900), .ZN(n1082) );
XOR2_X1 U904 ( .A(n1183), .B(n1223), .Z(G24) );
NOR2_X1 U905 ( .A1(KEYINPUT54), .A2(n1224), .ZN(n1223) );
INV_X1 U906 ( .A(G122), .ZN(n1224) );
AND4_X1 U907 ( .A1(n1225), .A2(n1066), .A3(n1075), .A4(n1209), .ZN(n1183) );
INV_X1 U908 ( .A(n1052), .ZN(n1066) );
NAND2_X1 U909 ( .A1(n1073), .A2(n1226), .ZN(n1052) );
XOR2_X1 U910 ( .A(G119), .B(n1187), .Z(G21) );
AND3_X1 U911 ( .A1(n1041), .A2(n1225), .A3(n1215), .ZN(n1187) );
INV_X1 U912 ( .A(n1205), .ZN(n1215) );
NAND2_X1 U913 ( .A1(n1227), .A2(n1228), .ZN(n1205) );
XOR2_X1 U914 ( .A(n1229), .B(n1182), .Z(G18) );
AND3_X1 U915 ( .A1(n1225), .A2(n1037), .A3(n1068), .ZN(n1182) );
NOR2_X1 U916 ( .A1(n1209), .A2(n1230), .ZN(n1037) );
NAND2_X1 U917 ( .A1(KEYINPUT41), .A2(n1231), .ZN(n1229) );
XNOR2_X1 U918 ( .A(G113), .B(n1179), .ZN(G15) );
NAND3_X1 U919 ( .A1(n1068), .A2(n1225), .A3(n1213), .ZN(n1179) );
INV_X1 U920 ( .A(n1028), .ZN(n1213) );
NAND2_X1 U921 ( .A1(n1230), .A2(n1209), .ZN(n1028) );
AND3_X1 U922 ( .A1(n1064), .A2(n1185), .A3(n1065), .ZN(n1225) );
NOR2_X1 U923 ( .A1(n1053), .A2(n1232), .ZN(n1065) );
NOR2_X1 U924 ( .A1(n1051), .A2(n1050), .ZN(n1232) );
INV_X1 U925 ( .A(n1233), .ZN(n1050) );
INV_X1 U926 ( .A(n1189), .ZN(n1064) );
INV_X1 U927 ( .A(n1211), .ZN(n1068) );
NAND2_X1 U928 ( .A1(n1226), .A2(n1228), .ZN(n1211) );
INV_X1 U929 ( .A(n1073), .ZN(n1228) );
INV_X1 U930 ( .A(n1227), .ZN(n1226) );
XOR2_X1 U931 ( .A(G110), .B(n1234), .Z(G12) );
NOR3_X1 U932 ( .A1(n1049), .A2(n1189), .A3(n1193), .ZN(n1234) );
NAND3_X1 U933 ( .A1(n1069), .A2(n1185), .A3(n1041), .ZN(n1193) );
NOR2_X1 U934 ( .A1(n1075), .A2(n1209), .ZN(n1041) );
NAND3_X1 U935 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1209) );
NAND2_X1 U936 ( .A1(n1238), .A2(n1239), .ZN(n1237) );
INV_X1 U937 ( .A(G475), .ZN(n1239) );
NAND3_X1 U938 ( .A1(n1240), .A2(n1241), .A3(n1242), .ZN(n1238) );
NAND2_X1 U939 ( .A1(KEYINPUT10), .A2(n1243), .ZN(n1242) );
NAND2_X1 U940 ( .A1(KEYINPUT59), .A2(n1244), .ZN(n1241) );
NAND2_X1 U941 ( .A1(n1245), .A2(n1246), .ZN(n1240) );
INV_X1 U942 ( .A(KEYINPUT59), .ZN(n1246) );
NAND2_X1 U943 ( .A1(n1244), .A2(n1247), .ZN(n1245) );
NAND2_X1 U944 ( .A1(KEYINPUT21), .A2(n1248), .ZN(n1247) );
NAND4_X1 U945 ( .A1(n1244), .A2(n1243), .A3(G475), .A4(n1248), .ZN(n1236) );
INV_X1 U946 ( .A(KEYINPUT10), .ZN(n1248) );
INV_X1 U947 ( .A(KEYINPUT21), .ZN(n1243) );
NAND2_X1 U948 ( .A1(KEYINPUT10), .A2(n1249), .ZN(n1235) );
NAND2_X1 U949 ( .A1(n1244), .A2(n1250), .ZN(n1249) );
NAND2_X1 U950 ( .A1(KEYINPUT21), .A2(G475), .ZN(n1250) );
INV_X1 U951 ( .A(n1077), .ZN(n1244) );
NOR2_X1 U952 ( .A1(n1142), .A2(G902), .ZN(n1077) );
XOR2_X1 U953 ( .A(n1251), .B(n1252), .Z(n1142) );
XOR2_X1 U954 ( .A(n1253), .B(n1254), .Z(n1252) );
XOR2_X1 U955 ( .A(G143), .B(n1255), .Z(n1254) );
NAND3_X1 U956 ( .A1(G214), .A2(n1256), .A3(KEYINPUT4), .ZN(n1253) );
XOR2_X1 U957 ( .A(n1257), .B(n1258), .Z(n1251) );
XOR2_X1 U958 ( .A(n1259), .B(n1260), .Z(n1258) );
NAND2_X1 U959 ( .A1(KEYINPUT36), .A2(G131), .ZN(n1260) );
NAND2_X1 U960 ( .A1(n1261), .A2(n1262), .ZN(n1259) );
OR2_X1 U961 ( .A1(n1263), .A2(n1143), .ZN(n1262) );
XOR2_X1 U962 ( .A(n1264), .B(KEYINPUT46), .Z(n1261) );
NAND2_X1 U963 ( .A1(n1265), .A2(n1263), .ZN(n1264) );
XNOR2_X1 U964 ( .A(n1266), .B(G113), .ZN(n1263) );
NAND2_X1 U965 ( .A1(KEYINPUT49), .A2(n1267), .ZN(n1266) );
XOR2_X1 U966 ( .A(n1143), .B(KEYINPUT55), .Z(n1265) );
NAND2_X1 U967 ( .A1(n1268), .A2(n1269), .ZN(n1257) );
OR2_X1 U968 ( .A1(n1219), .A2(n1169), .ZN(n1269) );
NAND2_X1 U969 ( .A1(n1270), .A2(n1219), .ZN(n1268) );
XNOR2_X1 U970 ( .A(n1169), .B(KEYINPUT42), .ZN(n1270) );
INV_X1 U971 ( .A(n1230), .ZN(n1075) );
XOR2_X1 U972 ( .A(n1271), .B(G478), .Z(n1230) );
OR2_X1 U973 ( .A1(n1136), .A2(G902), .ZN(n1271) );
XNOR2_X1 U974 ( .A(n1272), .B(n1273), .ZN(n1136) );
XOR2_X1 U975 ( .A(n1274), .B(n1275), .Z(n1273) );
XOR2_X1 U976 ( .A(n1231), .B(G107), .Z(n1275) );
NAND2_X1 U977 ( .A1(n1276), .A2(G217), .ZN(n1274) );
INV_X1 U978 ( .A(n1277), .ZN(n1276) );
XNOR2_X1 U979 ( .A(n1278), .B(n1267), .ZN(n1272) );
NAND2_X1 U980 ( .A1(n1279), .A2(KEYINPUT19), .ZN(n1278) );
XNOR2_X1 U981 ( .A(G134), .B(n1280), .ZN(n1279) );
NAND2_X1 U982 ( .A1(n1038), .A2(n1281), .ZN(n1185) );
NAND4_X1 U983 ( .A1(G953), .A2(G902), .A3(n1222), .A4(n1111), .ZN(n1281) );
INV_X1 U984 ( .A(G898), .ZN(n1111) );
NAND3_X1 U985 ( .A1(n1222), .A2(n1058), .A3(G952), .ZN(n1038) );
NAND2_X1 U986 ( .A1(G237), .A2(G234), .ZN(n1222) );
AND2_X1 U987 ( .A1(n1053), .A2(n1282), .ZN(n1069) );
NAND2_X1 U988 ( .A1(G221), .A2(n1233), .ZN(n1282) );
XNOR2_X1 U989 ( .A(n1283), .B(G469), .ZN(n1053) );
NAND2_X1 U990 ( .A1(n1284), .A2(n1285), .ZN(n1283) );
XOR2_X1 U991 ( .A(n1286), .B(n1287), .Z(n1284) );
XOR2_X1 U992 ( .A(n1288), .B(n1169), .Z(n1287) );
NAND2_X1 U993 ( .A1(KEYINPUT50), .A2(n1106), .ZN(n1288) );
INV_X1 U994 ( .A(n1102), .ZN(n1106) );
XOR2_X1 U995 ( .A(n1289), .B(n1290), .Z(n1286) );
XOR2_X1 U996 ( .A(G110), .B(n1164), .Z(n1290) );
NOR2_X1 U997 ( .A1(n1081), .A2(G953), .ZN(n1164) );
INV_X1 U998 ( .A(G227), .ZN(n1081) );
NAND3_X1 U999 ( .A1(n1291), .A2(n1292), .A3(n1293), .ZN(n1289) );
NAND2_X1 U1000 ( .A1(KEYINPUT29), .A2(n1103), .ZN(n1293) );
NAND3_X1 U1001 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(n1292) );
INV_X1 U1002 ( .A(KEYINPUT29), .ZN(n1295) );
OR2_X1 U1003 ( .A1(n1296), .A2(n1294), .ZN(n1291) );
AND2_X1 U1004 ( .A1(KEYINPUT43), .A2(n1105), .ZN(n1294) );
INV_X1 U1005 ( .A(n1103), .ZN(n1105) );
NAND2_X1 U1006 ( .A1(n1297), .A2(n1298), .ZN(n1103) );
NAND2_X1 U1007 ( .A1(n1280), .A2(G146), .ZN(n1298) );
NAND2_X1 U1008 ( .A1(n1299), .A2(n1255), .ZN(n1297) );
INV_X1 U1009 ( .A(G146), .ZN(n1255) );
XNOR2_X1 U1010 ( .A(n1280), .B(KEYINPUT2), .ZN(n1299) );
XNOR2_X1 U1011 ( .A(n1162), .B(n1300), .ZN(n1296) );
XOR2_X1 U1012 ( .A(KEYINPUT63), .B(G101), .Z(n1300) );
NAND3_X1 U1013 ( .A1(n1301), .A2(n1302), .A3(n1303), .ZN(n1162) );
NAND2_X1 U1014 ( .A1(KEYINPUT8), .A2(G104), .ZN(n1303) );
NAND3_X1 U1015 ( .A1(n1143), .A2(n1304), .A3(G107), .ZN(n1302) );
NAND2_X1 U1016 ( .A1(n1305), .A2(n1020), .ZN(n1301) );
INV_X1 U1017 ( .A(G107), .ZN(n1020) );
NAND2_X1 U1018 ( .A1(n1306), .A2(n1304), .ZN(n1305) );
INV_X1 U1019 ( .A(KEYINPUT8), .ZN(n1304) );
XOR2_X1 U1020 ( .A(n1143), .B(KEYINPUT6), .Z(n1306) );
INV_X1 U1021 ( .A(G104), .ZN(n1143) );
NAND2_X1 U1022 ( .A1(n1056), .A2(n1054), .ZN(n1189) );
NAND2_X1 U1023 ( .A1(G214), .A2(n1307), .ZN(n1054) );
XNOR2_X1 U1024 ( .A(KEYINPUT3), .B(n1308), .ZN(n1307) );
INV_X1 U1025 ( .A(n1217), .ZN(n1056) );
XNOR2_X1 U1026 ( .A(n1309), .B(n1177), .ZN(n1217) );
NAND2_X1 U1027 ( .A1(G210), .A2(n1308), .ZN(n1177) );
OR2_X1 U1028 ( .A1(n1310), .A2(G237), .ZN(n1308) );
XOR2_X1 U1029 ( .A(KEYINPUT47), .B(n1285), .Z(n1310) );
NAND2_X1 U1030 ( .A1(n1311), .A2(n1285), .ZN(n1309) );
XOR2_X1 U1031 ( .A(n1312), .B(n1173), .Z(n1311) );
XNOR2_X1 U1032 ( .A(n1313), .B(n1121), .ZN(n1173) );
XNOR2_X1 U1033 ( .A(n1314), .B(n1315), .ZN(n1121) );
XNOR2_X1 U1034 ( .A(n1267), .B(n1168), .ZN(n1315) );
XOR2_X1 U1035 ( .A(G101), .B(G110), .Z(n1168) );
XNOR2_X1 U1036 ( .A(G122), .B(KEYINPUT48), .ZN(n1267) );
XOR2_X1 U1037 ( .A(n1316), .B(G107), .Z(n1314) );
NAND2_X1 U1038 ( .A1(KEYINPUT57), .A2(G104), .ZN(n1316) );
NAND2_X1 U1039 ( .A1(KEYINPUT24), .A2(n1120), .ZN(n1313) );
NAND2_X1 U1040 ( .A1(n1317), .A2(KEYINPUT61), .ZN(n1312) );
XNOR2_X1 U1041 ( .A(n1175), .B(n1318), .ZN(n1317) );
NOR2_X1 U1042 ( .A1(KEYINPUT7), .A2(n1174), .ZN(n1318) );
XOR2_X1 U1043 ( .A(G125), .B(n1156), .Z(n1174) );
NOR2_X1 U1044 ( .A1(n1110), .A2(G953), .ZN(n1175) );
INV_X1 U1045 ( .A(G224), .ZN(n1110) );
NAND2_X1 U1046 ( .A1(n1227), .A2(n1073), .ZN(n1049) );
XOR2_X1 U1047 ( .A(n1319), .B(G472), .Z(n1073) );
NAND2_X1 U1048 ( .A1(n1320), .A2(n1285), .ZN(n1319) );
INV_X1 U1049 ( .A(G902), .ZN(n1285) );
XOR2_X1 U1050 ( .A(n1321), .B(n1322), .Z(n1320) );
XOR2_X1 U1051 ( .A(n1323), .B(n1324), .Z(n1322) );
NOR2_X1 U1052 ( .A1(G101), .A2(KEYINPUT26), .ZN(n1324) );
NOR2_X1 U1053 ( .A1(KEYINPUT15), .A2(n1120), .ZN(n1323) );
XOR2_X1 U1054 ( .A(n1325), .B(n1326), .Z(n1120) );
XOR2_X1 U1055 ( .A(KEYINPUT14), .B(G119), .Z(n1326) );
XOR2_X1 U1056 ( .A(G113), .B(n1231), .Z(n1325) );
INV_X1 U1057 ( .A(G116), .ZN(n1231) );
XNOR2_X1 U1058 ( .A(n1150), .B(n1156), .ZN(n1321) );
XOR2_X1 U1059 ( .A(G146), .B(n1280), .Z(n1156) );
XOR2_X1 U1060 ( .A(G143), .B(G128), .Z(n1280) );
XNOR2_X1 U1061 ( .A(n1102), .B(n1327), .ZN(n1150) );
AND2_X1 U1062 ( .A1(n1256), .A2(G210), .ZN(n1327) );
NOR2_X1 U1063 ( .A1(G953), .A2(G237), .ZN(n1256) );
XNOR2_X1 U1064 ( .A(G131), .B(n1328), .ZN(n1102) );
XOR2_X1 U1065 ( .A(G137), .B(G134), .Z(n1328) );
XOR2_X1 U1066 ( .A(n1071), .B(KEYINPUT44), .Z(n1227) );
XNOR2_X1 U1067 ( .A(n1329), .B(n1128), .ZN(n1071) );
NAND2_X1 U1068 ( .A1(G217), .A2(n1233), .ZN(n1128) );
NAND2_X1 U1069 ( .A1(G234), .A2(n1330), .ZN(n1233) );
XOR2_X1 U1070 ( .A(KEYINPUT47), .B(G902), .Z(n1330) );
OR2_X1 U1071 ( .A1(n1130), .A2(G902), .ZN(n1329) );
XNOR2_X1 U1072 ( .A(n1331), .B(n1332), .ZN(n1130) );
XOR2_X1 U1073 ( .A(G110), .B(n1333), .Z(n1332) );
XOR2_X1 U1074 ( .A(G146), .B(G137), .Z(n1333) );
XOR2_X1 U1075 ( .A(n1334), .B(n1335), .Z(n1331) );
NOR2_X1 U1076 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
NOR2_X1 U1077 ( .A1(KEYINPUT62), .A2(n1099), .ZN(n1337) );
AND2_X1 U1078 ( .A1(KEYINPUT52), .A2(n1099), .ZN(n1336) );
XNOR2_X1 U1079 ( .A(n1219), .B(n1169), .ZN(n1099) );
XOR2_X1 U1080 ( .A(G140), .B(KEYINPUT30), .Z(n1169) );
INV_X1 U1081 ( .A(G125), .ZN(n1219) );
XOR2_X1 U1082 ( .A(n1338), .B(n1339), .Z(n1334) );
NOR2_X1 U1083 ( .A1(n1277), .A2(n1051), .ZN(n1339) );
INV_X1 U1084 ( .A(G221), .ZN(n1051) );
NAND2_X1 U1085 ( .A1(G234), .A2(n1058), .ZN(n1277) );
INV_X1 U1086 ( .A(G953), .ZN(n1058) );
NAND3_X1 U1087 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1338) );
NAND2_X1 U1088 ( .A1(G119), .A2(n1343), .ZN(n1342) );
INV_X1 U1089 ( .A(KEYINPUT45), .ZN(n1343) );
NAND3_X1 U1090 ( .A1(KEYINPUT45), .A2(n1344), .A3(n1345), .ZN(n1341) );
OR2_X1 U1091 ( .A1(n1345), .A2(n1344), .ZN(n1340) );
NOR2_X1 U1092 ( .A1(G119), .A2(KEYINPUT60), .ZN(n1344) );
INV_X1 U1093 ( .A(G128), .ZN(n1345) );
endmodule


