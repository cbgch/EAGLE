//Key = 0000110000011111000001101011111010110110001000011010000100001000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338;

XNOR2_X1 U735 ( .A(n1024), .B(n1025), .ZN(G9) );
NOR2_X1 U736 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U737 ( .A1(n1028), .A2(n1029), .ZN(G75) );
XOR2_X1 U738 ( .A(KEYINPUT39), .B(n1030), .Z(n1029) );
NOR3_X1 U739 ( .A1(n1031), .A2(G953), .A3(G952), .ZN(n1030) );
NOR4_X1 U740 ( .A1(n1032), .A2(n1033), .A3(G953), .A4(n1031), .ZN(n1028) );
AND4_X1 U741 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1031) );
NOR4_X1 U742 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1037) );
XNOR2_X1 U743 ( .A(n1042), .B(n1043), .ZN(n1038) );
NAND2_X1 U744 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
XOR2_X1 U745 ( .A(KEYINPUT8), .B(KEYINPUT48), .Z(n1045) );
XNOR2_X1 U746 ( .A(n1046), .B(KEYINPUT57), .ZN(n1044) );
NOR3_X1 U747 ( .A1(n1047), .A2(n1048), .A3(n1049), .ZN(n1036) );
NOR2_X1 U748 ( .A1(n1050), .A2(n1051), .ZN(n1047) );
XNOR2_X1 U749 ( .A(n1052), .B(n1053), .ZN(n1035) );
XOR2_X1 U750 ( .A(KEYINPUT31), .B(KEYINPUT15), .Z(n1053) );
XOR2_X1 U751 ( .A(KEYINPUT38), .B(n1054), .Z(n1034) );
NOR2_X1 U752 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
XOR2_X1 U753 ( .A(KEYINPUT28), .B(n1050), .Z(n1056) );
NOR3_X1 U754 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n1033) );
NOR2_X1 U755 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
NOR2_X1 U756 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
NAND3_X1 U757 ( .A1(G952), .A2(n1064), .A3(n1065), .ZN(n1032) );
NAND2_X1 U758 ( .A1(n1066), .A2(n1067), .ZN(n1064) );
NAND3_X1 U759 ( .A1(n1068), .A2(n1069), .A3(n1070), .ZN(n1067) );
XOR2_X1 U760 ( .A(KEYINPUT32), .B(n1071), .Z(n1070) );
AND2_X1 U761 ( .A1(n1072), .A2(n1073), .ZN(n1071) );
NAND3_X1 U762 ( .A1(n1074), .A2(n1075), .A3(n1076), .ZN(n1069) );
NAND2_X1 U763 ( .A1(n1077), .A2(n1078), .ZN(n1075) );
NAND3_X1 U764 ( .A1(n1079), .A2(n1080), .A3(KEYINPUT0), .ZN(n1077) );
NAND3_X1 U765 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1074) );
NAND3_X1 U766 ( .A1(n1080), .A2(n1084), .A3(n1079), .ZN(n1082) );
INV_X1 U767 ( .A(KEYINPUT0), .ZN(n1084) );
NAND3_X1 U768 ( .A1(n1085), .A2(n1086), .A3(n1052), .ZN(n1081) );
OR2_X1 U769 ( .A1(n1087), .A2(n1079), .ZN(n1086) );
OR3_X1 U770 ( .A1(n1088), .A2(n1089), .A3(n1049), .ZN(n1085) );
NAND2_X1 U771 ( .A1(n1073), .A2(n1090), .ZN(n1068) );
INV_X1 U772 ( .A(n1057), .ZN(n1073) );
NAND3_X1 U773 ( .A1(n1079), .A2(n1091), .A3(n1083), .ZN(n1057) );
INV_X1 U774 ( .A(n1078), .ZN(n1083) );
NAND2_X1 U775 ( .A1(KEYINPUT60), .A2(n1092), .ZN(n1078) );
XOR2_X1 U776 ( .A(n1093), .B(n1094), .Z(G72) );
NOR2_X1 U777 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
NOR2_X1 U778 ( .A1(n1097), .A2(n1098), .ZN(n1095) );
NAND2_X1 U779 ( .A1(n1099), .A2(n1100), .ZN(n1093) );
NAND2_X1 U780 ( .A1(n1101), .A2(n1096), .ZN(n1100) );
XNOR2_X1 U781 ( .A(n1102), .B(n1103), .ZN(n1101) );
NOR2_X1 U782 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
XOR2_X1 U783 ( .A(KEYINPUT43), .B(n1106), .Z(n1105) );
NAND3_X1 U784 ( .A1(n1102), .A2(G900), .A3(G953), .ZN(n1099) );
XNOR2_X1 U785 ( .A(n1107), .B(n1108), .ZN(n1102) );
XNOR2_X1 U786 ( .A(n1109), .B(n1110), .ZN(n1108) );
NAND2_X1 U787 ( .A1(KEYINPUT4), .A2(n1111), .ZN(n1109) );
NAND2_X1 U788 ( .A1(n1112), .A2(n1113), .ZN(G69) );
NAND2_X1 U789 ( .A1(n1114), .A2(n1096), .ZN(n1113) );
XNOR2_X1 U790 ( .A(n1115), .B(n1116), .ZN(n1114) );
NAND2_X1 U791 ( .A1(n1117), .A2(G953), .ZN(n1112) );
NAND2_X1 U792 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
NAND2_X1 U793 ( .A1(n1116), .A2(n1120), .ZN(n1119) );
NAND2_X1 U794 ( .A1(G224), .A2(n1121), .ZN(n1118) );
NAND2_X1 U795 ( .A1(G898), .A2(n1116), .ZN(n1121) );
NAND2_X1 U796 ( .A1(n1122), .A2(n1123), .ZN(n1116) );
NAND2_X1 U797 ( .A1(G953), .A2(n1124), .ZN(n1123) );
XOR2_X1 U798 ( .A(n1125), .B(n1126), .Z(n1122) );
XNOR2_X1 U799 ( .A(n1127), .B(n1128), .ZN(n1126) );
NOR2_X1 U800 ( .A1(KEYINPUT18), .A2(n1129), .ZN(n1128) );
NOR2_X1 U801 ( .A1(n1130), .A2(n1131), .ZN(G66) );
XOR2_X1 U802 ( .A(n1132), .B(n1133), .Z(n1131) );
NAND2_X1 U803 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
NOR2_X1 U804 ( .A1(n1130), .A2(n1136), .ZN(G63) );
NOR3_X1 U805 ( .A1(n1046), .A2(n1137), .A3(n1138), .ZN(n1136) );
AND3_X1 U806 ( .A1(n1139), .A2(G478), .A3(n1134), .ZN(n1138) );
NOR2_X1 U807 ( .A1(n1140), .A2(n1139), .ZN(n1137) );
NOR2_X1 U808 ( .A1(n1065), .A2(n1043), .ZN(n1140) );
NOR2_X1 U809 ( .A1(n1130), .A2(n1141), .ZN(G60) );
XOR2_X1 U810 ( .A(n1142), .B(n1143), .Z(n1141) );
NAND2_X1 U811 ( .A1(n1134), .A2(G475), .ZN(n1142) );
XOR2_X1 U812 ( .A(G104), .B(n1144), .Z(G6) );
NOR2_X1 U813 ( .A1(n1130), .A2(n1145), .ZN(G57) );
NOR2_X1 U814 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
XOR2_X1 U815 ( .A(n1148), .B(KEYINPUT11), .Z(n1147) );
NAND2_X1 U816 ( .A1(n1149), .A2(n1150), .ZN(n1148) );
NOR2_X1 U817 ( .A1(n1150), .A2(n1149), .ZN(n1146) );
XNOR2_X1 U818 ( .A(n1151), .B(n1152), .ZN(n1149) );
NAND2_X1 U819 ( .A1(n1134), .A2(G472), .ZN(n1151) );
NOR2_X1 U820 ( .A1(n1130), .A2(n1153), .ZN(G54) );
NOR2_X1 U821 ( .A1(n1154), .A2(n1155), .ZN(n1153) );
XOR2_X1 U822 ( .A(n1156), .B(KEYINPUT22), .Z(n1155) );
NAND2_X1 U823 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NOR2_X1 U824 ( .A1(n1157), .A2(n1158), .ZN(n1154) );
XOR2_X1 U825 ( .A(n1159), .B(n1110), .Z(n1158) );
AND2_X1 U826 ( .A1(n1134), .A2(G469), .ZN(n1157) );
NOR2_X1 U827 ( .A1(n1130), .A2(n1160), .ZN(G51) );
XOR2_X1 U828 ( .A(n1161), .B(n1162), .Z(n1160) );
XOR2_X1 U829 ( .A(n1163), .B(n1164), .Z(n1161) );
NOR2_X1 U830 ( .A1(KEYINPUT53), .A2(n1165), .ZN(n1164) );
NAND3_X1 U831 ( .A1(n1166), .A2(n1167), .A3(n1050), .ZN(n1163) );
OR2_X1 U832 ( .A1(n1134), .A2(KEYINPUT61), .ZN(n1167) );
NOR2_X1 U833 ( .A1(n1168), .A2(n1065), .ZN(n1134) );
NAND2_X1 U834 ( .A1(KEYINPUT61), .A2(n1169), .ZN(n1166) );
NAND2_X1 U835 ( .A1(n1065), .A2(G902), .ZN(n1169) );
NOR3_X1 U836 ( .A1(n1115), .A2(n1106), .A3(n1104), .ZN(n1065) );
NAND4_X1 U837 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1104) );
AND3_X1 U838 ( .A1(n1174), .A2(n1175), .A3(n1176), .ZN(n1173) );
NAND2_X1 U839 ( .A1(n1066), .A2(n1177), .ZN(n1172) );
NAND2_X1 U840 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
XOR2_X1 U841 ( .A(KEYINPUT26), .B(n1180), .Z(n1179) );
XOR2_X1 U842 ( .A(n1181), .B(KEYINPUT20), .Z(n1178) );
NAND4_X1 U843 ( .A1(n1182), .A2(n1061), .A3(n1040), .A4(n1183), .ZN(n1170) );
NAND4_X1 U844 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1115) );
NOR4_X1 U845 ( .A1(n1144), .A2(n1188), .A3(n1189), .A4(n1190), .ZN(n1187) );
AND4_X1 U846 ( .A1(n1076), .A2(n1191), .A3(n1080), .A4(n1192), .ZN(n1144) );
NOR2_X1 U847 ( .A1(n1027), .A2(n1193), .ZN(n1192) );
NOR2_X1 U848 ( .A1(n1194), .A2(n1195), .ZN(n1186) );
NOR2_X1 U849 ( .A1(n1196), .A2(n1027), .ZN(n1195) );
INV_X1 U850 ( .A(n1061), .ZN(n1027) );
XOR2_X1 U851 ( .A(n1026), .B(KEYINPUT19), .Z(n1196) );
NAND4_X1 U852 ( .A1(n1080), .A2(n1076), .A3(n1088), .A4(n1191), .ZN(n1026) );
NOR2_X1 U853 ( .A1(n1096), .A2(G952), .ZN(n1130) );
XNOR2_X1 U854 ( .A(G146), .B(n1171), .ZN(G48) );
NAND3_X1 U855 ( .A1(n1089), .A2(n1061), .A3(n1197), .ZN(n1171) );
XOR2_X1 U856 ( .A(n1198), .B(n1199), .Z(G45) );
NAND2_X1 U857 ( .A1(KEYINPUT27), .A2(G143), .ZN(n1199) );
NAND4_X1 U858 ( .A1(n1200), .A2(n1182), .A3(n1040), .A4(n1183), .ZN(n1198) );
XNOR2_X1 U859 ( .A(n1061), .B(KEYINPUT21), .ZN(n1200) );
XOR2_X1 U860 ( .A(G140), .B(n1201), .Z(G42) );
NOR2_X1 U861 ( .A1(n1202), .A2(n1181), .ZN(n1201) );
NAND3_X1 U862 ( .A1(n1203), .A2(n1072), .A3(n1089), .ZN(n1181) );
INV_X1 U863 ( .A(n1066), .ZN(n1202) );
XOR2_X1 U864 ( .A(n1174), .B(n1204), .Z(G39) );
XNOR2_X1 U865 ( .A(G137), .B(KEYINPUT51), .ZN(n1204) );
NAND3_X1 U866 ( .A1(n1197), .A2(n1066), .A3(n1079), .ZN(n1174) );
XOR2_X1 U867 ( .A(n1205), .B(G134), .Z(G36) );
NAND2_X1 U868 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
NAND3_X1 U869 ( .A1(n1066), .A2(n1208), .A3(n1209), .ZN(n1207) );
INV_X1 U870 ( .A(KEYINPUT24), .ZN(n1209) );
NAND2_X1 U871 ( .A1(n1182), .A2(n1088), .ZN(n1208) );
NAND2_X1 U872 ( .A1(n1106), .A2(KEYINPUT24), .ZN(n1206) );
AND3_X1 U873 ( .A1(n1066), .A2(n1088), .A3(n1182), .ZN(n1106) );
XNOR2_X1 U874 ( .A(G131), .B(n1210), .ZN(G33) );
NAND2_X1 U875 ( .A1(n1180), .A2(n1066), .ZN(n1210) );
NOR2_X1 U876 ( .A1(n1062), .A2(n1048), .ZN(n1066) );
AND2_X1 U877 ( .A1(n1089), .A2(n1182), .ZN(n1180) );
AND2_X1 U878 ( .A1(n1090), .A2(n1203), .ZN(n1182) );
XNOR2_X1 U879 ( .A(G128), .B(n1176), .ZN(G30) );
NAND3_X1 U880 ( .A1(n1061), .A2(n1088), .A3(n1197), .ZN(n1176) );
AND3_X1 U881 ( .A1(n1211), .A2(n1212), .A3(n1203), .ZN(n1197) );
AND2_X1 U882 ( .A1(n1080), .A2(n1213), .ZN(n1203) );
XNOR2_X1 U883 ( .A(n1194), .B(n1214), .ZN(G3) );
NOR2_X1 U884 ( .A1(G101), .A2(KEYINPUT40), .ZN(n1214) );
AND2_X1 U885 ( .A1(n1215), .A2(n1090), .ZN(n1194) );
XNOR2_X1 U886 ( .A(G125), .B(n1175), .ZN(G27) );
NAND4_X1 U887 ( .A1(n1072), .A2(n1213), .A3(n1061), .A4(n1216), .ZN(n1175) );
NOR2_X1 U888 ( .A1(n1217), .A2(n1193), .ZN(n1216) );
NAND2_X1 U889 ( .A1(n1218), .A2(n1219), .ZN(n1213) );
NAND2_X1 U890 ( .A1(n1220), .A2(n1098), .ZN(n1218) );
INV_X1 U891 ( .A(G900), .ZN(n1098) );
XOR2_X1 U892 ( .A(n1184), .B(n1221), .Z(G24) );
XNOR2_X1 U893 ( .A(G122), .B(KEYINPUT36), .ZN(n1221) );
NAND4_X1 U894 ( .A1(n1222), .A2(n1076), .A3(n1040), .A4(n1183), .ZN(n1184) );
NAND2_X1 U895 ( .A1(n1223), .A2(n1224), .ZN(G21) );
NAND2_X1 U896 ( .A1(G119), .A2(n1185), .ZN(n1224) );
XOR2_X1 U897 ( .A(KEYINPUT30), .B(n1225), .Z(n1223) );
NOR2_X1 U898 ( .A1(G119), .A2(n1185), .ZN(n1225) );
NAND4_X1 U899 ( .A1(n1222), .A2(n1079), .A3(n1211), .A4(n1212), .ZN(n1185) );
XOR2_X1 U900 ( .A(n1190), .B(n1226), .Z(G18) );
NOR2_X1 U901 ( .A1(KEYINPUT7), .A2(n1227), .ZN(n1226) );
INV_X1 U902 ( .A(G116), .ZN(n1227) );
AND3_X1 U903 ( .A1(n1090), .A2(n1088), .A3(n1222), .ZN(n1190) );
NOR2_X1 U904 ( .A1(n1040), .A2(n1228), .ZN(n1088) );
XNOR2_X1 U905 ( .A(n1229), .B(n1189), .ZN(G15) );
AND3_X1 U906 ( .A1(n1089), .A2(n1090), .A3(n1222), .ZN(n1189) );
AND3_X1 U907 ( .A1(n1061), .A2(n1191), .A3(n1091), .ZN(n1222) );
INV_X1 U908 ( .A(n1217), .ZN(n1091) );
NAND2_X1 U909 ( .A1(n1052), .A2(n1087), .ZN(n1217) );
NOR2_X1 U910 ( .A1(n1212), .A2(n1230), .ZN(n1090) );
INV_X1 U911 ( .A(n1193), .ZN(n1089) );
NAND2_X1 U912 ( .A1(n1228), .A2(n1040), .ZN(n1193) );
XOR2_X1 U913 ( .A(n1188), .B(n1231), .Z(G12) );
XNOR2_X1 U914 ( .A(KEYINPUT46), .B(n1232), .ZN(n1231) );
AND2_X1 U915 ( .A1(n1215), .A2(n1072), .ZN(n1188) );
NAND2_X1 U916 ( .A1(n1233), .A2(n1234), .ZN(n1072) );
OR2_X1 U917 ( .A1(n1059), .A2(KEYINPUT42), .ZN(n1234) );
INV_X1 U918 ( .A(n1076), .ZN(n1059) );
NOR2_X1 U919 ( .A1(n1212), .A2(n1211), .ZN(n1076) );
NAND3_X1 U920 ( .A1(n1212), .A2(n1230), .A3(KEYINPUT42), .ZN(n1233) );
INV_X1 U921 ( .A(n1211), .ZN(n1230) );
XOR2_X1 U922 ( .A(n1041), .B(KEYINPUT9), .Z(n1211) );
XNOR2_X1 U923 ( .A(n1235), .B(n1236), .ZN(n1041) );
XOR2_X1 U924 ( .A(KEYINPUT62), .B(G472), .Z(n1236) );
NAND3_X1 U925 ( .A1(n1237), .A2(n1238), .A3(n1168), .ZN(n1235) );
NAND2_X1 U926 ( .A1(n1239), .A2(n1240), .ZN(n1238) );
INV_X1 U927 ( .A(KEYINPUT52), .ZN(n1240) );
XOR2_X1 U928 ( .A(n1150), .B(n1152), .Z(n1239) );
NAND3_X1 U929 ( .A1(n1152), .A2(n1150), .A3(KEYINPUT52), .ZN(n1237) );
XOR2_X1 U930 ( .A(n1241), .B(G101), .Z(n1150) );
NAND2_X1 U931 ( .A1(n1242), .A2(G210), .ZN(n1241) );
XOR2_X1 U932 ( .A(n1243), .B(n1244), .Z(n1152) );
XNOR2_X1 U933 ( .A(n1229), .B(n1110), .ZN(n1244) );
XNOR2_X1 U934 ( .A(n1245), .B(n1246), .ZN(n1243) );
XOR2_X1 U935 ( .A(n1039), .B(KEYINPUT33), .Z(n1212) );
XNOR2_X1 U936 ( .A(n1247), .B(n1135), .ZN(n1039) );
AND2_X1 U937 ( .A1(G217), .A2(n1248), .ZN(n1135) );
NAND2_X1 U938 ( .A1(n1133), .A2(n1168), .ZN(n1247) );
XNOR2_X1 U939 ( .A(n1249), .B(n1250), .ZN(n1133) );
NOR2_X1 U940 ( .A1(G137), .A2(n1251), .ZN(n1250) );
XOR2_X1 U941 ( .A(KEYINPUT59), .B(KEYINPUT45), .Z(n1251) );
XOR2_X1 U942 ( .A(n1252), .B(n1253), .Z(n1249) );
NOR2_X1 U943 ( .A1(n1254), .A2(n1255), .ZN(n1253) );
INV_X1 U944 ( .A(G221), .ZN(n1254) );
NAND3_X1 U945 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1252) );
NAND2_X1 U946 ( .A1(n1259), .A2(n1260), .ZN(n1258) );
OR3_X1 U947 ( .A1(n1260), .A2(n1111), .A3(G146), .ZN(n1257) );
NAND2_X1 U948 ( .A1(n1261), .A2(G146), .ZN(n1256) );
XOR2_X1 U949 ( .A(n1260), .B(n1111), .Z(n1261) );
NAND2_X1 U950 ( .A1(n1262), .A2(n1263), .ZN(n1260) );
NAND2_X1 U951 ( .A1(n1264), .A2(n1265), .ZN(n1263) );
NAND2_X1 U952 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U953 ( .A1(KEYINPUT12), .A2(n1268), .ZN(n1267) );
XOR2_X1 U954 ( .A(n1269), .B(KEYINPUT44), .Z(n1264) );
NAND2_X1 U955 ( .A1(n1270), .A2(n1271), .ZN(n1262) );
NAND2_X1 U956 ( .A1(n1266), .A2(KEYINPUT12), .ZN(n1271) );
XOR2_X1 U957 ( .A(n1269), .B(KEYINPUT2), .Z(n1266) );
XOR2_X1 U958 ( .A(n1272), .B(G128), .Z(n1269) );
NAND2_X1 U959 ( .A1(KEYINPUT14), .A2(G119), .ZN(n1272) );
INV_X1 U960 ( .A(n1268), .ZN(n1270) );
XOR2_X1 U961 ( .A(G110), .B(KEYINPUT23), .Z(n1268) );
AND4_X1 U962 ( .A1(n1079), .A2(n1061), .A3(n1080), .A4(n1191), .ZN(n1215) );
NAND2_X1 U963 ( .A1(n1273), .A2(n1219), .ZN(n1191) );
NAND3_X1 U964 ( .A1(n1092), .A2(n1096), .A3(G952), .ZN(n1219) );
NAND2_X1 U965 ( .A1(n1220), .A2(n1124), .ZN(n1273) );
INV_X1 U966 ( .A(G898), .ZN(n1124) );
AND3_X1 U967 ( .A1(G902), .A2(n1092), .A3(G953), .ZN(n1220) );
NAND2_X1 U968 ( .A1(G237), .A2(G234), .ZN(n1092) );
NOR2_X1 U969 ( .A1(n1052), .A2(n1049), .ZN(n1080) );
INV_X1 U970 ( .A(n1087), .ZN(n1049) );
NAND2_X1 U971 ( .A1(G221), .A2(n1248), .ZN(n1087) );
NAND2_X1 U972 ( .A1(n1274), .A2(n1168), .ZN(n1248) );
XNOR2_X1 U973 ( .A(G234), .B(KEYINPUT35), .ZN(n1274) );
XOR2_X1 U974 ( .A(n1275), .B(G469), .Z(n1052) );
NAND2_X1 U975 ( .A1(n1276), .A2(n1168), .ZN(n1275) );
XOR2_X1 U976 ( .A(n1277), .B(n1278), .Z(n1276) );
XOR2_X1 U977 ( .A(KEYINPUT58), .B(KEYINPUT16), .Z(n1278) );
XOR2_X1 U978 ( .A(n1159), .B(n1279), .Z(n1277) );
NOR2_X1 U979 ( .A1(KEYINPUT25), .A2(n1110), .ZN(n1279) );
XNOR2_X1 U980 ( .A(n1280), .B(n1281), .ZN(n1110) );
XOR2_X1 U981 ( .A(KEYINPUT50), .B(G137), .Z(n1281) );
XNOR2_X1 U982 ( .A(G134), .B(G131), .ZN(n1280) );
XOR2_X1 U983 ( .A(n1282), .B(n1283), .Z(n1159) );
XOR2_X1 U984 ( .A(G104), .B(n1284), .Z(n1283) );
XNOR2_X1 U985 ( .A(G140), .B(n1232), .ZN(n1284) );
INV_X1 U986 ( .A(G110), .ZN(n1232) );
XOR2_X1 U987 ( .A(n1107), .B(n1285), .Z(n1282) );
XOR2_X1 U988 ( .A(n1286), .B(n1287), .Z(n1285) );
NOR2_X1 U989 ( .A1(G953), .A2(n1097), .ZN(n1286) );
INV_X1 U990 ( .A(G227), .ZN(n1097) );
NAND2_X1 U991 ( .A1(n1288), .A2(n1289), .ZN(n1107) );
NAND3_X1 U992 ( .A1(n1290), .A2(n1291), .A3(n1292), .ZN(n1289) );
INV_X1 U993 ( .A(KEYINPUT13), .ZN(n1292) );
NAND2_X1 U994 ( .A1(n1245), .A2(KEYINPUT13), .ZN(n1288) );
NOR2_X1 U995 ( .A1(n1293), .A2(n1048), .ZN(n1061) );
INV_X1 U996 ( .A(n1063), .ZN(n1048) );
NAND2_X1 U997 ( .A1(G214), .A2(n1294), .ZN(n1063) );
INV_X1 U998 ( .A(n1062), .ZN(n1293) );
XOR2_X1 U999 ( .A(n1055), .B(n1050), .Z(n1062) );
AND2_X1 U1000 ( .A1(G210), .A2(n1294), .ZN(n1050) );
NAND2_X1 U1001 ( .A1(n1295), .A2(n1168), .ZN(n1294) );
INV_X1 U1002 ( .A(G237), .ZN(n1295) );
INV_X1 U1003 ( .A(n1051), .ZN(n1055) );
NAND2_X1 U1004 ( .A1(n1296), .A2(n1168), .ZN(n1051) );
XNOR2_X1 U1005 ( .A(n1165), .B(n1162), .ZN(n1296) );
XNOR2_X1 U1006 ( .A(n1125), .B(n1297), .ZN(n1162) );
XNOR2_X1 U1007 ( .A(n1298), .B(n1129), .ZN(n1297) );
XOR2_X1 U1008 ( .A(n1287), .B(n1299), .Z(n1129) );
NOR2_X1 U1009 ( .A1(G104), .A2(KEYINPUT1), .ZN(n1299) );
XNOR2_X1 U1010 ( .A(G101), .B(n1024), .ZN(n1287) );
NAND2_X1 U1011 ( .A1(n1300), .A2(n1127), .ZN(n1298) );
XOR2_X1 U1012 ( .A(G110), .B(n1301), .Z(n1127) );
XOR2_X1 U1013 ( .A(KEYINPUT34), .B(G122), .Z(n1301) );
XOR2_X1 U1014 ( .A(KEYINPUT29), .B(KEYINPUT10), .Z(n1300) );
NAND2_X1 U1015 ( .A1(n1302), .A2(n1303), .ZN(n1125) );
OR2_X1 U1016 ( .A1(n1246), .A2(G113), .ZN(n1303) );
NAND2_X1 U1017 ( .A1(n1246), .A2(n1304), .ZN(n1302) );
XNOR2_X1 U1018 ( .A(G113), .B(KEYINPUT5), .ZN(n1304) );
XOR2_X1 U1019 ( .A(G116), .B(G119), .Z(n1246) );
XNOR2_X1 U1020 ( .A(n1245), .B(n1305), .ZN(n1165) );
XNOR2_X1 U1021 ( .A(n1306), .B(n1307), .ZN(n1305) );
NOR2_X1 U1022 ( .A1(G953), .A2(n1120), .ZN(n1307) );
INV_X1 U1023 ( .A(G224), .ZN(n1120) );
INV_X1 U1024 ( .A(G125), .ZN(n1306) );
XOR2_X1 U1025 ( .A(n1291), .B(n1290), .Z(n1245) );
XNOR2_X1 U1026 ( .A(G128), .B(KEYINPUT54), .ZN(n1290) );
XNOR2_X1 U1027 ( .A(G143), .B(n1308), .ZN(n1291) );
XNOR2_X1 U1028 ( .A(KEYINPUT49), .B(n1309), .ZN(n1308) );
NOR2_X1 U1029 ( .A1(n1183), .A2(n1040), .ZN(n1079) );
XNOR2_X1 U1030 ( .A(n1310), .B(G475), .ZN(n1040) );
NAND2_X1 U1031 ( .A1(n1143), .A2(n1168), .ZN(n1310) );
INV_X1 U1032 ( .A(G902), .ZN(n1168) );
XNOR2_X1 U1033 ( .A(n1311), .B(n1312), .ZN(n1143) );
NOR2_X1 U1034 ( .A1(n1259), .A2(n1313), .ZN(n1312) );
XOR2_X1 U1035 ( .A(KEYINPUT41), .B(n1314), .Z(n1313) );
NOR2_X1 U1036 ( .A1(n1111), .A2(n1309), .ZN(n1314) );
AND2_X1 U1037 ( .A1(n1111), .A2(n1309), .ZN(n1259) );
INV_X1 U1038 ( .A(G146), .ZN(n1309) );
XNOR2_X1 U1039 ( .A(G125), .B(G140), .ZN(n1111) );
XOR2_X1 U1040 ( .A(n1315), .B(n1316), .Z(n1311) );
NOR2_X1 U1041 ( .A1(KEYINPUT56), .A2(n1317), .ZN(n1316) );
XNOR2_X1 U1042 ( .A(G104), .B(n1318), .ZN(n1317) );
NAND3_X1 U1043 ( .A1(n1319), .A2(n1320), .A3(KEYINPUT47), .ZN(n1318) );
OR3_X1 U1044 ( .A1(n1229), .A2(G122), .A3(KEYINPUT55), .ZN(n1320) );
INV_X1 U1045 ( .A(G113), .ZN(n1229) );
NAND2_X1 U1046 ( .A1(n1321), .A2(KEYINPUT55), .ZN(n1319) );
XOR2_X1 U1047 ( .A(G122), .B(n1322), .Z(n1321) );
NOR2_X1 U1048 ( .A1(G113), .A2(KEYINPUT3), .ZN(n1322) );
NAND2_X1 U1049 ( .A1(n1323), .A2(n1324), .ZN(n1315) );
NAND2_X1 U1050 ( .A1(n1325), .A2(n1326), .ZN(n1324) );
XOR2_X1 U1051 ( .A(n1327), .B(KEYINPUT63), .Z(n1323) );
OR2_X1 U1052 ( .A1(n1325), .A2(n1326), .ZN(n1327) );
INV_X1 U1053 ( .A(G131), .ZN(n1326) );
XNOR2_X1 U1054 ( .A(n1328), .B(G143), .ZN(n1325) );
NAND2_X1 U1055 ( .A1(n1242), .A2(G214), .ZN(n1328) );
NOR2_X1 U1056 ( .A1(G953), .A2(G237), .ZN(n1242) );
INV_X1 U1057 ( .A(n1228), .ZN(n1183) );
XOR2_X1 U1058 ( .A(n1046), .B(n1043), .Z(n1228) );
INV_X1 U1059 ( .A(G478), .ZN(n1043) );
NOR2_X1 U1060 ( .A1(n1139), .A2(G902), .ZN(n1046) );
XOR2_X1 U1061 ( .A(n1329), .B(n1330), .Z(n1139) );
NOR2_X1 U1062 ( .A1(n1331), .A2(n1255), .ZN(n1330) );
NAND2_X1 U1063 ( .A1(G234), .A2(n1096), .ZN(n1255) );
INV_X1 U1064 ( .A(G953), .ZN(n1096) );
INV_X1 U1065 ( .A(G217), .ZN(n1331) );
NAND2_X1 U1066 ( .A1(n1332), .A2(KEYINPUT37), .ZN(n1329) );
XOR2_X1 U1067 ( .A(n1333), .B(n1334), .Z(n1332) );
XOR2_X1 U1068 ( .A(G122), .B(n1335), .Z(n1334) );
XOR2_X1 U1069 ( .A(G134), .B(G128), .Z(n1335) );
XOR2_X1 U1070 ( .A(n1336), .B(n1337), .Z(n1333) );
NOR2_X1 U1071 ( .A1(G143), .A2(KEYINPUT6), .ZN(n1337) );
XNOR2_X1 U1072 ( .A(G116), .B(n1338), .ZN(n1336) );
NOR2_X1 U1073 ( .A1(KEYINPUT17), .A2(n1024), .ZN(n1338) );
INV_X1 U1074 ( .A(G107), .ZN(n1024) );
endmodule


