//Key = 0100110100010110000110011000001011101101111011011110010001110011


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
n1440;

XOR2_X1 U795 ( .A(G107), .B(n1100), .Z(G9) );
NOR2_X1 U796 ( .A1(n1101), .A2(n1102), .ZN(G75) );
NOR3_X1 U797 ( .A1(n1103), .A2(n1104), .A3(n1105), .ZN(n1102) );
NAND3_X1 U798 ( .A1(n1106), .A2(n1107), .A3(n1108), .ZN(n1103) );
NAND2_X1 U799 ( .A1(n1109), .A2(n1110), .ZN(n1108) );
NAND2_X1 U800 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
NAND3_X1 U801 ( .A1(n1113), .A2(n1114), .A3(n1115), .ZN(n1112) );
NAND3_X1 U802 ( .A1(n1116), .A2(n1117), .A3(n1118), .ZN(n1114) );
NAND2_X1 U803 ( .A1(n1119), .A2(n1120), .ZN(n1118) );
INV_X1 U804 ( .A(n1121), .ZN(n1117) );
NAND3_X1 U805 ( .A1(n1122), .A2(n1123), .A3(n1124), .ZN(n1111) );
NAND2_X1 U806 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
NAND4_X1 U807 ( .A1(n1127), .A2(n1115), .A3(n1113), .A4(n1128), .ZN(n1126) );
NAND2_X1 U808 ( .A1(n1119), .A2(n1129), .ZN(n1125) );
NAND2_X1 U809 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
NAND2_X1 U810 ( .A1(n1115), .A2(n1132), .ZN(n1131) );
NAND2_X1 U811 ( .A1(n1133), .A2(n1134), .ZN(n1132) );
NAND2_X1 U812 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
INV_X1 U813 ( .A(n1137), .ZN(n1133) );
NAND2_X1 U814 ( .A1(n1113), .A2(n1138), .ZN(n1130) );
NAND2_X1 U815 ( .A1(n1139), .A2(n1140), .ZN(n1138) );
NAND2_X1 U816 ( .A1(n1141), .A2(n1142), .ZN(n1140) );
INV_X1 U817 ( .A(n1143), .ZN(n1109) );
NOR3_X1 U818 ( .A1(n1144), .A2(G953), .A3(G952), .ZN(n1101) );
INV_X1 U819 ( .A(n1106), .ZN(n1144) );
NAND4_X1 U820 ( .A1(n1145), .A2(n1146), .A3(n1147), .A4(n1148), .ZN(n1106) );
NOR4_X1 U821 ( .A1(n1141), .A2(n1128), .A3(n1149), .A4(n1150), .ZN(n1148) );
XNOR2_X1 U822 ( .A(n1151), .B(KEYINPUT20), .ZN(n1150) );
XNOR2_X1 U823 ( .A(n1152), .B(KEYINPUT48), .ZN(n1149) );
NOR2_X1 U824 ( .A1(n1136), .A2(n1153), .ZN(n1147) );
XOR2_X1 U825 ( .A(n1154), .B(n1155), .Z(n1146) );
XNOR2_X1 U826 ( .A(KEYINPUT52), .B(n1156), .ZN(n1155) );
XNOR2_X1 U827 ( .A(n1157), .B(n1158), .ZN(n1145) );
XOR2_X1 U828 ( .A(n1159), .B(n1160), .Z(G72) );
NAND2_X1 U829 ( .A1(G953), .A2(n1161), .ZN(n1160) );
NAND2_X1 U830 ( .A1(G900), .A2(G227), .ZN(n1161) );
NAND2_X1 U831 ( .A1(KEYINPUT1), .A2(n1162), .ZN(n1159) );
XOR2_X1 U832 ( .A(n1163), .B(n1164), .Z(n1162) );
AND2_X1 U833 ( .A1(n1105), .A2(n1107), .ZN(n1164) );
NOR2_X1 U834 ( .A1(n1165), .A2(n1166), .ZN(n1163) );
XOR2_X1 U835 ( .A(n1167), .B(n1168), .Z(n1166) );
XNOR2_X1 U836 ( .A(n1169), .B(n1170), .ZN(n1168) );
XNOR2_X1 U837 ( .A(n1171), .B(n1172), .ZN(n1170) );
NOR2_X1 U838 ( .A1(KEYINPUT43), .A2(n1173), .ZN(n1172) );
XNOR2_X1 U839 ( .A(n1174), .B(n1175), .ZN(n1167) );
XNOR2_X1 U840 ( .A(n1176), .B(G134), .ZN(n1175) );
XNOR2_X1 U841 ( .A(n1177), .B(KEYINPUT34), .ZN(n1165) );
XOR2_X1 U842 ( .A(n1178), .B(n1179), .Z(G69) );
XOR2_X1 U843 ( .A(n1180), .B(n1181), .Z(n1179) );
NOR2_X1 U844 ( .A1(n1182), .A2(n1183), .ZN(n1181) );
XNOR2_X1 U845 ( .A(n1184), .B(n1185), .ZN(n1183) );
XNOR2_X1 U846 ( .A(n1186), .B(KEYINPUT26), .ZN(n1184) );
NAND3_X1 U847 ( .A1(G953), .A2(n1187), .A3(KEYINPUT50), .ZN(n1180) );
NAND2_X1 U848 ( .A1(G898), .A2(G224), .ZN(n1187) );
NAND2_X1 U849 ( .A1(n1107), .A2(n1104), .ZN(n1178) );
NOR2_X1 U850 ( .A1(n1188), .A2(n1189), .ZN(G66) );
XOR2_X1 U851 ( .A(n1190), .B(n1191), .Z(n1189) );
NAND2_X1 U852 ( .A1(n1192), .A2(n1193), .ZN(n1190) );
XOR2_X1 U853 ( .A(n1194), .B(KEYINPUT13), .Z(n1192) );
NOR2_X1 U854 ( .A1(n1188), .A2(n1195), .ZN(G63) );
XNOR2_X1 U855 ( .A(n1196), .B(n1197), .ZN(n1195) );
NAND3_X1 U856 ( .A1(n1193), .A2(G478), .A3(KEYINPUT39), .ZN(n1196) );
NOR2_X1 U857 ( .A1(n1188), .A2(n1198), .ZN(G60) );
XNOR2_X1 U858 ( .A(n1199), .B(n1200), .ZN(n1198) );
NAND2_X1 U859 ( .A1(n1193), .A2(G475), .ZN(n1199) );
INV_X1 U860 ( .A(n1201), .ZN(n1193) );
XOR2_X1 U861 ( .A(G104), .B(n1202), .Z(G6) );
NOR2_X1 U862 ( .A1(n1188), .A2(n1203), .ZN(G57) );
XOR2_X1 U863 ( .A(n1204), .B(n1205), .Z(n1203) );
XNOR2_X1 U864 ( .A(n1206), .B(n1207), .ZN(n1205) );
NOR4_X1 U865 ( .A1(n1208), .A2(n1209), .A3(KEYINPUT27), .A4(n1156), .ZN(n1206) );
NOR2_X1 U866 ( .A1(KEYINPUT30), .A2(n1210), .ZN(n1209) );
NOR3_X1 U867 ( .A1(n1105), .A2(n1211), .A3(n1104), .ZN(n1210) );
AND2_X1 U868 ( .A1(n1201), .A2(KEYINPUT30), .ZN(n1208) );
XOR2_X1 U869 ( .A(n1212), .B(n1213), .Z(n1204) );
NOR2_X1 U870 ( .A1(G101), .A2(KEYINPUT55), .ZN(n1213) );
NOR3_X1 U871 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(G54) );
AND2_X1 U872 ( .A1(KEYINPUT5), .A2(n1188), .ZN(n1216) );
NOR3_X1 U873 ( .A1(KEYINPUT5), .A2(G953), .A3(G952), .ZN(n1215) );
NOR3_X1 U874 ( .A1(n1217), .A2(n1218), .A3(n1219), .ZN(n1214) );
AND2_X1 U875 ( .A1(n1220), .A2(KEYINPUT0), .ZN(n1219) );
NOR3_X1 U876 ( .A1(KEYINPUT0), .A2(n1221), .A3(n1220), .ZN(n1218) );
NOR3_X1 U877 ( .A1(n1201), .A2(KEYINPUT3), .A3(n1222), .ZN(n1221) );
NOR3_X1 U878 ( .A1(n1201), .A2(n1223), .A3(n1222), .ZN(n1217) );
NOR2_X1 U879 ( .A1(n1224), .A2(KEYINPUT0), .ZN(n1223) );
NOR2_X1 U880 ( .A1(KEYINPUT3), .A2(n1225), .ZN(n1224) );
INV_X1 U881 ( .A(n1220), .ZN(n1225) );
XNOR2_X1 U882 ( .A(n1226), .B(n1227), .ZN(n1220) );
XOR2_X1 U883 ( .A(n1228), .B(n1229), .Z(n1227) );
XNOR2_X1 U884 ( .A(n1230), .B(n1231), .ZN(n1226) );
NOR3_X1 U885 ( .A1(n1232), .A2(n1188), .A3(n1233), .ZN(G51) );
AND3_X1 U886 ( .A1(n1234), .A2(n1235), .A3(n1236), .ZN(n1233) );
NOR2_X1 U887 ( .A1(n1107), .A2(G952), .ZN(n1188) );
NOR3_X1 U888 ( .A1(n1237), .A2(n1238), .A3(n1239), .ZN(n1232) );
NOR2_X1 U889 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
INV_X1 U890 ( .A(KEYINPUT44), .ZN(n1241) );
NOR2_X1 U891 ( .A1(n1242), .A2(n1243), .ZN(n1240) );
NOR2_X1 U892 ( .A1(n1244), .A2(n1245), .ZN(n1243) );
NOR2_X1 U893 ( .A1(n1246), .A2(n1247), .ZN(n1242) );
NOR2_X1 U894 ( .A1(KEYINPUT44), .A2(n1234), .ZN(n1238) );
NAND2_X1 U895 ( .A1(n1248), .A2(n1249), .ZN(n1234) );
NAND2_X1 U896 ( .A1(n1245), .A2(n1244), .ZN(n1249) );
XNOR2_X1 U897 ( .A(n1246), .B(KEYINPUT29), .ZN(n1244) );
NAND2_X1 U898 ( .A1(n1247), .A2(n1246), .ZN(n1248) );
OR2_X1 U899 ( .A1(n1201), .A2(n1158), .ZN(n1246) );
NAND2_X1 U900 ( .A1(G902), .A2(n1250), .ZN(n1201) );
OR2_X1 U901 ( .A1(n1105), .A2(n1104), .ZN(n1250) );
NAND4_X1 U902 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1104) );
NOR4_X1 U903 ( .A1(n1255), .A2(n1256), .A3(n1100), .A4(n1202), .ZN(n1254) );
AND2_X1 U904 ( .A1(n1257), .A2(n1258), .ZN(n1202) );
AND2_X1 U905 ( .A1(n1120), .A2(n1258), .ZN(n1100) );
AND4_X1 U906 ( .A1(n1259), .A2(n1260), .A3(n1113), .A4(n1261), .ZN(n1258) );
INV_X1 U907 ( .A(n1262), .ZN(n1260) );
INV_X1 U908 ( .A(n1263), .ZN(n1255) );
NAND2_X1 U909 ( .A1(n1264), .A2(n1265), .ZN(n1253) );
NAND2_X1 U910 ( .A1(n1266), .A2(n1267), .ZN(n1265) );
NAND2_X1 U911 ( .A1(n1268), .A2(n1113), .ZN(n1267) );
NAND4_X1 U912 ( .A1(n1121), .A2(n1269), .A3(n1137), .A4(n1261), .ZN(n1251) );
XNOR2_X1 U913 ( .A(KEYINPUT35), .B(n1139), .ZN(n1269) );
NAND2_X1 U914 ( .A1(n1270), .A2(n1271), .ZN(n1105) );
NOR4_X1 U915 ( .A1(n1272), .A2(n1273), .A3(n1274), .A4(n1275), .ZN(n1271) );
AND4_X1 U916 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1270) );
OR3_X1 U917 ( .A1(n1266), .A2(n1280), .A3(n1281), .ZN(n1279) );
XNOR2_X1 U918 ( .A(n1115), .B(KEYINPUT60), .ZN(n1280) );
AND2_X1 U919 ( .A1(n1235), .A2(n1236), .ZN(n1237) );
NAND2_X1 U920 ( .A1(n1282), .A2(n1283), .ZN(G48) );
NAND2_X1 U921 ( .A1(n1284), .A2(n1278), .ZN(n1283) );
NAND2_X1 U922 ( .A1(n1285), .A2(n1286), .ZN(n1284) );
NAND2_X1 U923 ( .A1(KEYINPUT14), .A2(n1287), .ZN(n1286) );
INV_X1 U924 ( .A(KEYINPUT62), .ZN(n1287) );
NAND3_X1 U925 ( .A1(n1288), .A2(n1289), .A3(KEYINPUT62), .ZN(n1282) );
OR2_X1 U926 ( .A1(G146), .A2(KEYINPUT14), .ZN(n1289) );
NAND2_X1 U927 ( .A1(KEYINPUT14), .A2(n1290), .ZN(n1288) );
OR2_X1 U928 ( .A1(n1278), .A2(G146), .ZN(n1290) );
NAND2_X1 U929 ( .A1(n1291), .A2(n1257), .ZN(n1278) );
XNOR2_X1 U930 ( .A(G143), .B(n1277), .ZN(G45) );
NAND4_X1 U931 ( .A1(n1268), .A2(n1292), .A3(n1259), .A4(n1137), .ZN(n1277) );
XNOR2_X1 U932 ( .A(G140), .B(n1276), .ZN(G42) );
NAND4_X1 U933 ( .A1(n1115), .A2(n1292), .A3(n1293), .A4(n1257), .ZN(n1276) );
NOR2_X1 U934 ( .A1(n1294), .A2(n1295), .ZN(n1293) );
XNOR2_X1 U935 ( .A(n1176), .B(n1296), .ZN(G39) );
NOR3_X1 U936 ( .A1(n1297), .A2(n1298), .A3(n1266), .ZN(n1296) );
NAND3_X1 U937 ( .A1(n1299), .A2(n1300), .A3(n1301), .ZN(n1297) );
XNOR2_X1 U938 ( .A(KEYINPUT38), .B(KEYINPUT18), .ZN(n1301) );
OR2_X1 U939 ( .A1(n1292), .A2(KEYINPUT21), .ZN(n1300) );
NAND2_X1 U940 ( .A1(KEYINPUT21), .A2(n1302), .ZN(n1299) );
NAND2_X1 U941 ( .A1(n1303), .A2(n1262), .ZN(n1302) );
NAND2_X1 U942 ( .A1(n1304), .A2(n1305), .ZN(G36) );
NAND2_X1 U943 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
NAND2_X1 U944 ( .A1(G134), .A2(n1308), .ZN(n1304) );
NAND2_X1 U945 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
NAND2_X1 U946 ( .A1(n1275), .A2(n1311), .ZN(n1310) );
INV_X1 U947 ( .A(n1312), .ZN(n1275) );
OR2_X1 U948 ( .A1(n1311), .A2(n1306), .ZN(n1309) );
NOR2_X1 U949 ( .A1(KEYINPUT54), .A2(n1312), .ZN(n1306) );
NAND4_X1 U950 ( .A1(n1115), .A2(n1292), .A3(n1120), .A4(n1137), .ZN(n1312) );
INV_X1 U951 ( .A(KEYINPUT23), .ZN(n1311) );
NAND2_X1 U952 ( .A1(n1313), .A2(n1314), .ZN(G33) );
NAND2_X1 U953 ( .A1(n1273), .A2(n1174), .ZN(n1314) );
XOR2_X1 U954 ( .A(KEYINPUT36), .B(n1315), .Z(n1313) );
NOR2_X1 U955 ( .A1(n1273), .A2(n1174), .ZN(n1315) );
INV_X1 U956 ( .A(G131), .ZN(n1174) );
AND4_X1 U957 ( .A1(n1115), .A2(n1292), .A3(n1257), .A4(n1137), .ZN(n1273) );
INV_X1 U958 ( .A(n1298), .ZN(n1115) );
NAND2_X1 U959 ( .A1(n1142), .A2(n1316), .ZN(n1298) );
XOR2_X1 U960 ( .A(G128), .B(n1274), .Z(G30) );
AND2_X1 U961 ( .A1(n1291), .A2(n1120), .ZN(n1274) );
NOR4_X1 U962 ( .A1(n1135), .A2(n1281), .A3(n1139), .A4(n1294), .ZN(n1291) );
INV_X1 U963 ( .A(n1292), .ZN(n1281) );
NOR2_X1 U964 ( .A1(n1262), .A2(n1317), .ZN(n1292) );
XNOR2_X1 U965 ( .A(G101), .B(n1318), .ZN(G3) );
NAND4_X1 U966 ( .A1(n1121), .A2(n1259), .A3(n1137), .A4(n1261), .ZN(n1318) );
XNOR2_X1 U967 ( .A(n1319), .B(n1171), .ZN(G27) );
NAND2_X1 U968 ( .A1(n1320), .A2(n1321), .ZN(n1319) );
NAND2_X1 U969 ( .A1(n1272), .A2(n1322), .ZN(n1321) );
INV_X1 U970 ( .A(KEYINPUT56), .ZN(n1322) );
AND3_X1 U971 ( .A1(n1323), .A2(n1303), .A3(n1324), .ZN(n1272) );
NAND4_X1 U972 ( .A1(n1324), .A2(n1323), .A3(n1317), .A4(KEYINPUT56), .ZN(n1320) );
INV_X1 U973 ( .A(n1303), .ZN(n1317) );
NAND2_X1 U974 ( .A1(n1143), .A2(n1325), .ZN(n1303) );
NAND3_X1 U975 ( .A1(G902), .A2(n1326), .A3(n1177), .ZN(n1325) );
NOR2_X1 U976 ( .A1(n1327), .A2(G900), .ZN(n1177) );
INV_X1 U977 ( .A(n1116), .ZN(n1323) );
NAND2_X1 U978 ( .A1(n1119), .A2(n1257), .ZN(n1116) );
XNOR2_X1 U979 ( .A(n1328), .B(n1329), .ZN(G24) );
NOR2_X1 U980 ( .A1(n1330), .A2(n1139), .ZN(n1329) );
XOR2_X1 U981 ( .A(n1331), .B(KEYINPUT46), .Z(n1330) );
NAND4_X1 U982 ( .A1(n1119), .A2(n1113), .A3(n1332), .A4(n1261), .ZN(n1331) );
XOR2_X1 U983 ( .A(KEYINPUT28), .B(n1268), .Z(n1332) );
NOR2_X1 U984 ( .A1(n1124), .A2(n1122), .ZN(n1268) );
XOR2_X1 U985 ( .A(G119), .B(n1333), .Z(G21) );
NOR2_X1 U986 ( .A1(n1266), .A2(n1334), .ZN(n1333) );
NAND4_X1 U987 ( .A1(n1124), .A2(n1295), .A3(n1122), .A4(n1136), .ZN(n1266) );
XNOR2_X1 U988 ( .A(G116), .B(n1252), .ZN(G18) );
NAND3_X1 U989 ( .A1(n1120), .A2(n1137), .A3(n1264), .ZN(n1252) );
NOR2_X1 U990 ( .A1(n1152), .A2(n1124), .ZN(n1120) );
INV_X1 U991 ( .A(n1151), .ZN(n1124) );
XNOR2_X1 U992 ( .A(G113), .B(n1335), .ZN(G15) );
NAND2_X1 U993 ( .A1(KEYINPUT53), .A2(n1256), .ZN(n1335) );
AND3_X1 U994 ( .A1(n1257), .A2(n1137), .A3(n1264), .ZN(n1256) );
INV_X1 U995 ( .A(n1334), .ZN(n1264) );
NAND3_X1 U996 ( .A1(n1259), .A2(n1261), .A3(n1119), .ZN(n1334) );
AND2_X1 U997 ( .A1(n1127), .A2(n1336), .ZN(n1119) );
INV_X1 U998 ( .A(n1153), .ZN(n1127) );
NAND2_X1 U999 ( .A1(n1337), .A2(n1338), .ZN(n1137) );
NAND2_X1 U1000 ( .A1(n1113), .A2(n1339), .ZN(n1338) );
INV_X1 U1001 ( .A(KEYINPUT58), .ZN(n1339) );
NOR2_X1 U1002 ( .A1(n1136), .A2(n1295), .ZN(n1113) );
NAND3_X1 U1003 ( .A1(n1294), .A2(n1295), .A3(KEYINPUT58), .ZN(n1337) );
NOR2_X1 U1004 ( .A1(n1151), .A2(n1122), .ZN(n1257) );
INV_X1 U1005 ( .A(n1152), .ZN(n1122) );
XNOR2_X1 U1006 ( .A(n1340), .B(n1341), .ZN(G12) );
NOR2_X1 U1007 ( .A1(KEYINPUT61), .A2(n1263), .ZN(n1341) );
NAND3_X1 U1008 ( .A1(n1324), .A2(n1261), .A3(n1121), .ZN(n1263) );
NOR3_X1 U1009 ( .A1(n1152), .A2(n1262), .A3(n1151), .ZN(n1121) );
XOR2_X1 U1010 ( .A(G478), .B(n1342), .Z(n1151) );
NOR2_X1 U1011 ( .A1(G902), .A2(n1197), .ZN(n1342) );
NAND3_X1 U1012 ( .A1(n1343), .A2(n1344), .A3(n1345), .ZN(n1197) );
NAND2_X1 U1013 ( .A1(n1346), .A2(n1347), .ZN(n1345) );
OR4_X1 U1014 ( .A1(n1346), .A2(KEYINPUT6), .A3(n1347), .A4(n1348), .ZN(n1344) );
INV_X1 U1015 ( .A(KEYINPUT7), .ZN(n1347) );
NAND2_X1 U1016 ( .A1(G217), .A2(n1349), .ZN(n1346) );
NAND2_X1 U1017 ( .A1(n1348), .A2(n1350), .ZN(n1343) );
NAND3_X1 U1018 ( .A1(n1349), .A2(n1351), .A3(G217), .ZN(n1350) );
INV_X1 U1019 ( .A(KEYINPUT6), .ZN(n1351) );
XOR2_X1 U1020 ( .A(n1352), .B(n1353), .Z(n1348) );
XOR2_X1 U1021 ( .A(n1354), .B(n1355), .Z(n1353) );
XNOR2_X1 U1022 ( .A(n1307), .B(G128), .ZN(n1355) );
INV_X1 U1023 ( .A(G134), .ZN(n1307) );
XOR2_X1 U1024 ( .A(KEYINPUT9), .B(G143), .Z(n1354) );
XNOR2_X1 U1025 ( .A(G107), .B(n1356), .ZN(n1352) );
NAND2_X1 U1026 ( .A1(n1336), .A2(n1153), .ZN(n1262) );
XOR2_X1 U1027 ( .A(n1357), .B(n1222), .Z(n1153) );
INV_X1 U1028 ( .A(G469), .ZN(n1222) );
NAND2_X1 U1029 ( .A1(n1358), .A2(n1211), .ZN(n1357) );
XOR2_X1 U1030 ( .A(n1359), .B(n1360), .Z(n1358) );
XOR2_X1 U1031 ( .A(n1228), .B(n1361), .Z(n1360) );
NOR2_X1 U1032 ( .A1(KEYINPUT25), .A2(n1229), .ZN(n1361) );
XNOR2_X1 U1033 ( .A(G110), .B(G140), .ZN(n1229) );
XNOR2_X1 U1034 ( .A(n1186), .B(n1362), .ZN(n1228) );
XOR2_X1 U1035 ( .A(n1363), .B(n1231), .Z(n1359) );
AND2_X1 U1036 ( .A1(G227), .A2(n1107), .ZN(n1231) );
NAND2_X1 U1037 ( .A1(KEYINPUT41), .A2(n1169), .ZN(n1363) );
INV_X1 U1038 ( .A(n1230), .ZN(n1169) );
XOR2_X1 U1039 ( .A(G143), .B(n1364), .Z(n1230) );
XOR2_X1 U1040 ( .A(n1128), .B(KEYINPUT47), .Z(n1336) );
AND2_X1 U1041 ( .A1(G221), .A2(n1365), .ZN(n1128) );
XOR2_X1 U1042 ( .A(G475), .B(n1366), .Z(n1152) );
NOR2_X1 U1043 ( .A1(G902), .A2(n1200), .ZN(n1366) );
NAND3_X1 U1044 ( .A1(n1367), .A2(n1368), .A3(n1369), .ZN(n1200) );
NAND2_X1 U1045 ( .A1(n1370), .A2(n1371), .ZN(n1369) );
OR3_X1 U1046 ( .A1(n1371), .A2(n1370), .A3(KEYINPUT31), .ZN(n1368) );
XOR2_X1 U1047 ( .A(n1372), .B(n1373), .Z(n1370) );
XNOR2_X1 U1048 ( .A(n1374), .B(G104), .ZN(n1373) );
NAND2_X1 U1049 ( .A1(KEYINPUT63), .A2(n1328), .ZN(n1372) );
NAND2_X1 U1050 ( .A1(KEYINPUT19), .A2(n1375), .ZN(n1371) );
INV_X1 U1051 ( .A(n1376), .ZN(n1375) );
NAND2_X1 U1052 ( .A1(KEYINPUT31), .A2(n1376), .ZN(n1367) );
XOR2_X1 U1053 ( .A(n1377), .B(n1378), .Z(n1376) );
XNOR2_X1 U1054 ( .A(n1379), .B(n1380), .ZN(n1378) );
NAND2_X1 U1055 ( .A1(KEYINPUT45), .A2(G131), .ZN(n1379) );
XOR2_X1 U1056 ( .A(n1381), .B(n1382), .Z(n1377) );
NOR2_X1 U1057 ( .A1(G146), .A2(KEYINPUT10), .ZN(n1382) );
XOR2_X1 U1058 ( .A(n1383), .B(G143), .Z(n1381) );
NAND2_X1 U1059 ( .A1(G214), .A2(n1384), .ZN(n1383) );
NAND2_X1 U1060 ( .A1(n1143), .A2(n1385), .ZN(n1261) );
NAND3_X1 U1061 ( .A1(n1182), .A2(n1326), .A3(G902), .ZN(n1385) );
NOR2_X1 U1062 ( .A1(n1327), .A2(G898), .ZN(n1182) );
XNOR2_X1 U1063 ( .A(G953), .B(KEYINPUT8), .ZN(n1327) );
NAND3_X1 U1064 ( .A1(n1326), .A2(n1107), .A3(G952), .ZN(n1143) );
NAND2_X1 U1065 ( .A1(G237), .A2(G234), .ZN(n1326) );
NOR3_X1 U1066 ( .A1(n1295), .A2(n1294), .A3(n1139), .ZN(n1324) );
INV_X1 U1067 ( .A(n1259), .ZN(n1139) );
NOR2_X1 U1068 ( .A1(n1142), .A2(n1141), .ZN(n1259) );
INV_X1 U1069 ( .A(n1316), .ZN(n1141) );
NAND2_X1 U1070 ( .A1(G214), .A2(n1386), .ZN(n1316) );
XOR2_X1 U1071 ( .A(n1387), .B(n1388), .Z(n1142) );
XNOR2_X1 U1072 ( .A(KEYINPUT49), .B(n1157), .ZN(n1388) );
NAND2_X1 U1073 ( .A1(n1389), .A2(n1211), .ZN(n1157) );
XNOR2_X1 U1074 ( .A(n1390), .B(n1247), .ZN(n1389) );
INV_X1 U1075 ( .A(n1245), .ZN(n1247) );
NAND2_X1 U1076 ( .A1(n1391), .A2(n1392), .ZN(n1245) );
NAND2_X1 U1077 ( .A1(n1185), .A2(n1393), .ZN(n1392) );
INV_X1 U1078 ( .A(n1186), .ZN(n1393) );
NAND2_X1 U1079 ( .A1(n1394), .A2(n1186), .ZN(n1391) );
XOR2_X1 U1080 ( .A(G101), .B(n1395), .Z(n1186) );
XOR2_X1 U1081 ( .A(G107), .B(G104), .Z(n1395) );
XNOR2_X1 U1082 ( .A(KEYINPUT15), .B(n1185), .ZN(n1394) );
XOR2_X1 U1083 ( .A(n1396), .B(n1397), .Z(n1185) );
XNOR2_X1 U1084 ( .A(n1340), .B(n1398), .ZN(n1397) );
NOR2_X1 U1085 ( .A1(G119), .A2(KEYINPUT2), .ZN(n1398) );
XNOR2_X1 U1086 ( .A(G113), .B(n1356), .ZN(n1396) );
XNOR2_X1 U1087 ( .A(n1328), .B(G116), .ZN(n1356) );
INV_X1 U1088 ( .A(G122), .ZN(n1328) );
NAND2_X1 U1089 ( .A1(n1399), .A2(n1236), .ZN(n1390) );
NAND2_X1 U1090 ( .A1(n1400), .A2(n1401), .ZN(n1236) );
NAND2_X1 U1091 ( .A1(G224), .A2(n1107), .ZN(n1401) );
XNOR2_X1 U1092 ( .A(G125), .B(n1402), .ZN(n1400) );
XOR2_X1 U1093 ( .A(n1235), .B(KEYINPUT16), .Z(n1399) );
NAND3_X1 U1094 ( .A1(n1403), .A2(n1107), .A3(G224), .ZN(n1235) );
XNOR2_X1 U1095 ( .A(n1171), .B(n1402), .ZN(n1403) );
INV_X1 U1096 ( .A(G125), .ZN(n1171) );
NAND2_X1 U1097 ( .A1(KEYINPUT33), .A2(n1158), .ZN(n1387) );
NAND2_X1 U1098 ( .A1(G210), .A2(n1386), .ZN(n1158) );
NAND2_X1 U1099 ( .A1(n1404), .A2(n1211), .ZN(n1386) );
XNOR2_X1 U1100 ( .A(G237), .B(KEYINPUT17), .ZN(n1404) );
INV_X1 U1101 ( .A(n1136), .ZN(n1294) );
XOR2_X1 U1102 ( .A(n1405), .B(n1194), .Z(n1136) );
NAND2_X1 U1103 ( .A1(G217), .A2(n1365), .ZN(n1194) );
NAND2_X1 U1104 ( .A1(G234), .A2(n1211), .ZN(n1365) );
NAND2_X1 U1105 ( .A1(n1191), .A2(n1211), .ZN(n1405) );
XOR2_X1 U1106 ( .A(n1406), .B(n1407), .Z(n1191) );
XNOR2_X1 U1107 ( .A(G137), .B(n1408), .ZN(n1407) );
NAND2_X1 U1108 ( .A1(G221), .A2(n1349), .ZN(n1408) );
AND2_X1 U1109 ( .A1(G234), .A2(n1107), .ZN(n1349) );
INV_X1 U1110 ( .A(G953), .ZN(n1107) );
NAND2_X1 U1111 ( .A1(n1409), .A2(n1410), .ZN(n1406) );
NAND2_X1 U1112 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
NAND2_X1 U1113 ( .A1(n1413), .A2(n1414), .ZN(n1411) );
NAND2_X1 U1114 ( .A1(n1415), .A2(n1285), .ZN(n1414) );
NAND2_X1 U1115 ( .A1(n1416), .A2(G146), .ZN(n1413) );
NAND2_X1 U1116 ( .A1(n1417), .A2(n1418), .ZN(n1409) );
NAND2_X1 U1117 ( .A1(n1419), .A2(n1420), .ZN(n1418) );
NAND2_X1 U1118 ( .A1(n1416), .A2(n1285), .ZN(n1420) );
XOR2_X1 U1119 ( .A(n1415), .B(n1421), .Z(n1416) );
XOR2_X1 U1120 ( .A(KEYINPUT51), .B(KEYINPUT32), .Z(n1421) );
NAND2_X1 U1121 ( .A1(n1415), .A2(G146), .ZN(n1419) );
AND2_X1 U1122 ( .A1(n1422), .A2(n1423), .ZN(n1415) );
NAND2_X1 U1123 ( .A1(n1424), .A2(n1340), .ZN(n1423) );
XOR2_X1 U1124 ( .A(n1425), .B(G128), .Z(n1424) );
XOR2_X1 U1125 ( .A(n1426), .B(KEYINPUT22), .Z(n1422) );
NAND2_X1 U1126 ( .A1(G110), .A2(n1427), .ZN(n1426) );
XNOR2_X1 U1127 ( .A(G128), .B(n1425), .ZN(n1427) );
NAND2_X1 U1128 ( .A1(KEYINPUT4), .A2(G119), .ZN(n1425) );
INV_X1 U1129 ( .A(n1412), .ZN(n1417) );
NAND2_X1 U1130 ( .A1(KEYINPUT37), .A2(n1380), .ZN(n1412) );
XNOR2_X1 U1131 ( .A(G125), .B(n1173), .ZN(n1380) );
INV_X1 U1132 ( .A(G140), .ZN(n1173) );
INV_X1 U1133 ( .A(n1135), .ZN(n1295) );
XOR2_X1 U1134 ( .A(n1428), .B(n1156), .Z(n1135) );
INV_X1 U1135 ( .A(G472), .ZN(n1156) );
NAND2_X1 U1136 ( .A1(KEYINPUT42), .A2(n1154), .ZN(n1428) );
NAND2_X1 U1137 ( .A1(n1429), .A2(n1211), .ZN(n1154) );
INV_X1 U1138 ( .A(G902), .ZN(n1211) );
XOR2_X1 U1139 ( .A(n1212), .B(n1430), .Z(n1429) );
XOR2_X1 U1140 ( .A(n1207), .B(n1431), .Z(n1430) );
NAND2_X1 U1141 ( .A1(n1432), .A2(KEYINPUT11), .ZN(n1431) );
XNOR2_X1 U1142 ( .A(G101), .B(KEYINPUT24), .ZN(n1432) );
NAND2_X1 U1143 ( .A1(G210), .A2(n1384), .ZN(n1207) );
NOR2_X1 U1144 ( .A1(G953), .A2(G237), .ZN(n1384) );
XOR2_X1 U1145 ( .A(n1433), .B(n1434), .Z(n1212) );
XOR2_X1 U1146 ( .A(G116), .B(n1435), .Z(n1434) );
XOR2_X1 U1147 ( .A(KEYINPUT59), .B(G119), .Z(n1435) );
XNOR2_X1 U1148 ( .A(n1402), .B(n1436), .ZN(n1433) );
XNOR2_X1 U1149 ( .A(n1374), .B(n1362), .ZN(n1436) );
XNOR2_X1 U1150 ( .A(n1437), .B(G131), .ZN(n1362) );
NAND2_X1 U1151 ( .A1(KEYINPUT40), .A2(n1438), .ZN(n1437) );
XNOR2_X1 U1152 ( .A(G134), .B(n1439), .ZN(n1438) );
NAND2_X1 U1153 ( .A1(KEYINPUT57), .A2(n1176), .ZN(n1439) );
INV_X1 U1154 ( .A(G137), .ZN(n1176) );
INV_X1 U1155 ( .A(G113), .ZN(n1374) );
XOR2_X1 U1156 ( .A(n1364), .B(n1440), .Z(n1402) );
NOR2_X1 U1157 ( .A1(G143), .A2(KEYINPUT12), .ZN(n1440) );
XNOR2_X1 U1158 ( .A(G128), .B(n1285), .ZN(n1364) );
INV_X1 U1159 ( .A(G146), .ZN(n1285) );
INV_X1 U1160 ( .A(G110), .ZN(n1340) );
endmodule


