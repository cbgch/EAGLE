//Key = 0010010010111011110010011010110101010001001001110101100010100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
n1322, n1323, n1324, n1325, n1326;

XOR2_X1 U732 ( .A(G107), .B(n1012), .Z(G9) );
NOR2_X1 U733 ( .A1(n1013), .A2(n1014), .ZN(G75) );
NOR4_X1 U734 ( .A1(G953), .A2(n1015), .A3(n1016), .A4(n1017), .ZN(n1014) );
NOR2_X1 U735 ( .A1(n1018), .A2(n1019), .ZN(n1016) );
NOR2_X1 U736 ( .A1(n1020), .A2(n1021), .ZN(n1018) );
NOR2_X1 U737 ( .A1(n1022), .A2(n1023), .ZN(n1021) );
NOR2_X1 U738 ( .A1(n1024), .A2(n1025), .ZN(n1022) );
NOR2_X1 U739 ( .A1(n1026), .A2(n1027), .ZN(n1025) );
NOR2_X1 U740 ( .A1(n1028), .A2(n1029), .ZN(n1026) );
NOR2_X1 U741 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
XOR2_X1 U742 ( .A(n1032), .B(KEYINPUT27), .Z(n1030) );
NOR3_X1 U743 ( .A1(n1032), .A2(n1033), .A3(n1034), .ZN(n1028) );
NOR2_X1 U744 ( .A1(n1035), .A2(n1036), .ZN(n1024) );
NOR2_X1 U745 ( .A1(n1037), .A2(n1038), .ZN(n1035) );
NOR2_X1 U746 ( .A1(n1033), .A2(n1027), .ZN(n1038) );
NOR3_X1 U747 ( .A1(n1039), .A2(n1040), .A3(n1041), .ZN(n1033) );
NOR2_X1 U748 ( .A1(n1042), .A2(n1032), .ZN(n1037) );
NOR2_X1 U749 ( .A1(n1043), .A2(n1044), .ZN(n1042) );
NOR4_X1 U750 ( .A1(n1045), .A2(n1032), .A3(n1027), .A4(n1036), .ZN(n1020) );
INV_X1 U751 ( .A(n1046), .ZN(n1036) );
INV_X1 U752 ( .A(n1047), .ZN(n1027) );
NOR2_X1 U753 ( .A1(n1048), .A2(n1049), .ZN(n1045) );
AND2_X1 U754 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
NOR3_X1 U755 ( .A1(n1015), .A2(G953), .A3(G952), .ZN(n1013) );
AND4_X1 U756 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1015) );
NOR4_X1 U757 ( .A1(n1041), .A2(n1051), .A3(n1056), .A4(n1057), .ZN(n1055) );
XNOR2_X1 U758 ( .A(n1058), .B(n1059), .ZN(n1057) );
NAND2_X1 U759 ( .A1(n1060), .A2(KEYINPUT39), .ZN(n1058) );
XOR2_X1 U760 ( .A(n1061), .B(KEYINPUT18), .Z(n1060) );
XOR2_X1 U761 ( .A(n1062), .B(KEYINPUT41), .Z(n1056) );
NAND2_X1 U762 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
XOR2_X1 U763 ( .A(n1065), .B(KEYINPUT44), .Z(n1063) );
NOR2_X1 U764 ( .A1(n1066), .A2(n1067), .ZN(n1054) );
XOR2_X1 U765 ( .A(KEYINPUT29), .B(n1068), .Z(n1053) );
XOR2_X1 U766 ( .A(n1069), .B(n1070), .Z(G72) );
NOR3_X1 U767 ( .A1(KEYINPUT3), .A2(n1071), .A3(n1072), .ZN(n1070) );
NOR2_X1 U768 ( .A1(n1073), .A2(n1074), .ZN(n1072) );
XOR2_X1 U769 ( .A(KEYINPUT5), .B(n1075), .Z(n1073) );
NOR2_X1 U770 ( .A1(n1076), .A2(n1077), .ZN(n1071) );
XOR2_X1 U771 ( .A(KEYINPUT38), .B(n1075), .Z(n1077) );
NOR2_X1 U772 ( .A1(G953), .A2(n1078), .ZN(n1075) );
INV_X1 U773 ( .A(n1074), .ZN(n1076) );
NAND2_X1 U774 ( .A1(n1079), .A2(n1080), .ZN(n1074) );
NAND2_X1 U775 ( .A1(G953), .A2(n1081), .ZN(n1080) );
XOR2_X1 U776 ( .A(KEYINPUT10), .B(G900), .Z(n1081) );
XOR2_X1 U777 ( .A(n1082), .B(n1083), .Z(n1079) );
XOR2_X1 U778 ( .A(n1084), .B(n1085), .Z(n1083) );
NOR2_X1 U779 ( .A1(G134), .A2(KEYINPUT54), .ZN(n1085) );
XOR2_X1 U780 ( .A(n1086), .B(n1087), .Z(n1082) );
NOR2_X1 U781 ( .A1(n1088), .A2(n1089), .ZN(n1069) );
XOR2_X1 U782 ( .A(KEYINPUT6), .B(n1090), .Z(n1089) );
NOR2_X1 U783 ( .A1(n1091), .A2(n1092), .ZN(n1090) );
XOR2_X1 U784 ( .A(n1093), .B(n1094), .Z(G69) );
XOR2_X1 U785 ( .A(n1095), .B(n1096), .Z(n1094) );
NAND2_X1 U786 ( .A1(n1097), .A2(n1088), .ZN(n1096) );
XOR2_X1 U787 ( .A(KEYINPUT58), .B(n1098), .Z(n1097) );
NAND2_X1 U788 ( .A1(n1099), .A2(n1100), .ZN(n1095) );
NAND2_X1 U789 ( .A1(G953), .A2(n1101), .ZN(n1100) );
XNOR2_X1 U790 ( .A(n1102), .B(n1103), .ZN(n1099) );
NOR2_X1 U791 ( .A1(n1104), .A2(n1088), .ZN(n1093) );
NOR2_X1 U792 ( .A1(n1105), .A2(n1101), .ZN(n1104) );
NOR2_X1 U793 ( .A1(n1106), .A2(n1107), .ZN(G66) );
XOR2_X1 U794 ( .A(n1108), .B(n1109), .Z(n1107) );
NOR2_X1 U795 ( .A1(KEYINPUT19), .A2(n1110), .ZN(n1108) );
NOR3_X1 U796 ( .A1(n1111), .A2(n1112), .A3(n1113), .ZN(n1110) );
XOR2_X1 U797 ( .A(n1017), .B(KEYINPUT42), .Z(n1112) );
NOR2_X1 U798 ( .A1(n1106), .A2(n1114), .ZN(G63) );
XNOR2_X1 U799 ( .A(n1115), .B(n1116), .ZN(n1114) );
XOR2_X1 U800 ( .A(KEYINPUT60), .B(n1117), .Z(n1116) );
NOR2_X1 U801 ( .A1(n1118), .A2(n1119), .ZN(n1117) );
INV_X1 U802 ( .A(G478), .ZN(n1118) );
NOR2_X1 U803 ( .A1(n1106), .A2(n1120), .ZN(G60) );
XOR2_X1 U804 ( .A(n1121), .B(n1122), .Z(n1120) );
NOR2_X1 U805 ( .A1(n1123), .A2(KEYINPUT34), .ZN(n1121) );
NOR2_X1 U806 ( .A1(n1124), .A2(n1119), .ZN(n1123) );
XNOR2_X1 U807 ( .A(G104), .B(n1125), .ZN(G6) );
NOR2_X1 U808 ( .A1(n1106), .A2(n1126), .ZN(G57) );
NOR3_X1 U809 ( .A1(n1127), .A2(n1128), .A3(n1129), .ZN(n1126) );
NOR2_X1 U810 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
INV_X1 U811 ( .A(n1132), .ZN(n1131) );
NOR2_X1 U812 ( .A1(KEYINPUT21), .A2(n1133), .ZN(n1130) );
XNOR2_X1 U813 ( .A(n1134), .B(KEYINPUT35), .ZN(n1133) );
NOR3_X1 U814 ( .A1(n1132), .A2(KEYINPUT21), .A3(n1134), .ZN(n1128) );
XOR2_X1 U815 ( .A(n1135), .B(n1136), .Z(n1132) );
NOR2_X1 U816 ( .A1(KEYINPUT53), .A2(n1137), .ZN(n1136) );
XOR2_X1 U817 ( .A(n1138), .B(n1139), .Z(n1137) );
NOR2_X1 U818 ( .A1(n1140), .A2(n1141), .ZN(n1138) );
NOR2_X1 U819 ( .A1(n1142), .A2(n1143), .ZN(n1141) );
XNOR2_X1 U820 ( .A(n1144), .B(KEYINPUT37), .ZN(n1143) );
NOR2_X1 U821 ( .A1(n1144), .A2(n1145), .ZN(n1140) );
OR2_X1 U822 ( .A1(n1119), .A2(n1061), .ZN(n1135) );
INV_X1 U823 ( .A(G472), .ZN(n1061) );
AND2_X1 U824 ( .A1(n1134), .A2(KEYINPUT21), .ZN(n1127) );
XOR2_X1 U825 ( .A(n1146), .B(n1147), .Z(n1134) );
NAND2_X1 U826 ( .A1(n1148), .A2(KEYINPUT8), .ZN(n1146) );
XNOR2_X1 U827 ( .A(G101), .B(KEYINPUT40), .ZN(n1148) );
NOR2_X1 U828 ( .A1(n1149), .A2(n1150), .ZN(G54) );
XOR2_X1 U829 ( .A(KEYINPUT55), .B(n1106), .Z(n1150) );
XOR2_X1 U830 ( .A(n1151), .B(n1152), .Z(n1149) );
XOR2_X1 U831 ( .A(n1153), .B(n1154), .Z(n1152) );
NOR2_X1 U832 ( .A1(n1155), .A2(n1156), .ZN(n1154) );
NOR2_X1 U833 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
XNOR2_X1 U834 ( .A(n1086), .B(KEYINPUT57), .ZN(n1158) );
NOR2_X1 U835 ( .A1(n1086), .A2(n1159), .ZN(n1155) );
NAND2_X1 U836 ( .A1(KEYINPUT56), .A2(n1160), .ZN(n1153) );
XOR2_X1 U837 ( .A(n1161), .B(n1162), .Z(n1151) );
NOR2_X1 U838 ( .A1(n1163), .A2(n1119), .ZN(n1162) );
INV_X1 U839 ( .A(G469), .ZN(n1163) );
XOR2_X1 U840 ( .A(n1164), .B(n1165), .Z(n1161) );
NAND2_X1 U841 ( .A1(KEYINPUT14), .A2(n1145), .ZN(n1164) );
NOR2_X1 U842 ( .A1(n1106), .A2(n1166), .ZN(G51) );
XOR2_X1 U843 ( .A(n1167), .B(n1168), .Z(n1166) );
XOR2_X1 U844 ( .A(n1169), .B(n1170), .Z(n1168) );
NOR2_X1 U845 ( .A1(n1171), .A2(n1119), .ZN(n1170) );
NAND2_X1 U846 ( .A1(G902), .A2(n1017), .ZN(n1119) );
NAND2_X1 U847 ( .A1(n1098), .A2(n1078), .ZN(n1017) );
AND4_X1 U848 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1078) );
NOR4_X1 U849 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1175) );
AND2_X1 U850 ( .A1(n1180), .A2(n1181), .ZN(n1174) );
NAND4_X1 U851 ( .A1(n1182), .A2(n1039), .A3(n1183), .A4(n1066), .ZN(n1173) );
NAND2_X1 U852 ( .A1(n1184), .A2(n1185), .ZN(n1172) );
AND4_X1 U853 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(n1098) );
NOR4_X1 U854 ( .A1(n1190), .A2(n1191), .A3(n1012), .A4(n1192), .ZN(n1189) );
AND3_X1 U855 ( .A1(n1043), .A2(n1193), .A3(n1194), .ZN(n1012) );
AND2_X1 U856 ( .A1(n1195), .A2(n1125), .ZN(n1188) );
NAND3_X1 U857 ( .A1(n1194), .A2(n1193), .A3(n1044), .ZN(n1125) );
XOR2_X1 U858 ( .A(n1196), .B(n1197), .Z(n1167) );
NAND2_X1 U859 ( .A1(KEYINPUT2), .A2(n1198), .ZN(n1196) );
NOR2_X1 U860 ( .A1(n1088), .A2(G952), .ZN(n1106) );
XOR2_X1 U861 ( .A(G146), .B(n1179), .Z(G48) );
AND3_X1 U862 ( .A1(n1199), .A2(n1044), .A3(n1182), .ZN(n1179) );
XNOR2_X1 U863 ( .A(G143), .B(n1200), .ZN(G45) );
NAND4_X1 U864 ( .A1(n1201), .A2(n1182), .A3(n1183), .A4(n1066), .ZN(n1200) );
XNOR2_X1 U865 ( .A(n1039), .B(KEYINPUT16), .ZN(n1201) );
NAND2_X1 U866 ( .A1(n1202), .A2(n1203), .ZN(G42) );
OR2_X1 U867 ( .A1(n1181), .A2(G140), .ZN(n1203) );
XOR2_X1 U868 ( .A(n1204), .B(KEYINPUT36), .Z(n1202) );
NAND2_X1 U869 ( .A1(G140), .A2(n1181), .ZN(n1204) );
NAND3_X1 U870 ( .A1(n1040), .A2(n1044), .A3(n1205), .ZN(n1181) );
XOR2_X1 U871 ( .A(G137), .B(n1178), .Z(G39) );
AND3_X1 U872 ( .A1(n1199), .A2(n1047), .A3(n1205), .ZN(n1178) );
XNOR2_X1 U873 ( .A(G134), .B(n1206), .ZN(G36) );
NAND2_X1 U874 ( .A1(KEYINPUT45), .A2(n1177), .ZN(n1206) );
AND3_X1 U875 ( .A1(n1039), .A2(n1043), .A3(n1205), .ZN(n1177) );
NAND2_X1 U876 ( .A1(n1207), .A2(n1208), .ZN(G33) );
NAND2_X1 U877 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
NAND2_X1 U878 ( .A1(G131), .A2(n1211), .ZN(n1207) );
NAND2_X1 U879 ( .A1(n1212), .A2(n1213), .ZN(n1211) );
NAND2_X1 U880 ( .A1(KEYINPUT9), .A2(n1214), .ZN(n1213) );
INV_X1 U881 ( .A(n1180), .ZN(n1214) );
OR2_X1 U882 ( .A1(n1209), .A2(KEYINPUT9), .ZN(n1212) );
NOR2_X1 U883 ( .A1(KEYINPUT63), .A2(n1180), .ZN(n1209) );
NAND3_X1 U884 ( .A1(n1044), .A2(n1039), .A3(n1205), .ZN(n1180) );
AND3_X1 U885 ( .A1(n1049), .A2(n1215), .A3(n1046), .ZN(n1205) );
NOR2_X1 U886 ( .A1(n1034), .A2(n1041), .ZN(n1046) );
INV_X1 U887 ( .A(n1216), .ZN(n1041) );
XNOR2_X1 U888 ( .A(n1176), .B(n1217), .ZN(G30) );
XOR2_X1 U889 ( .A(KEYINPUT28), .B(G128), .Z(n1217) );
AND3_X1 U890 ( .A1(n1199), .A2(n1043), .A3(n1182), .ZN(n1176) );
AND3_X1 U891 ( .A1(n1049), .A2(n1215), .A3(n1185), .ZN(n1182) );
XOR2_X1 U892 ( .A(n1195), .B(n1218), .Z(G3) );
NAND2_X1 U893 ( .A1(KEYINPUT47), .A2(n1219), .ZN(n1218) );
XOR2_X1 U894 ( .A(KEYINPUT43), .B(G101), .Z(n1219) );
NAND3_X1 U895 ( .A1(n1039), .A2(n1194), .A3(n1047), .ZN(n1195) );
XNOR2_X1 U896 ( .A(G125), .B(n1220), .ZN(G27) );
NAND3_X1 U897 ( .A1(n1185), .A2(n1221), .A3(KEYINPUT52), .ZN(n1220) );
XOR2_X1 U898 ( .A(KEYINPUT25), .B(n1184), .Z(n1221) );
AND4_X1 U899 ( .A1(n1040), .A2(n1044), .A3(n1222), .A4(n1215), .ZN(n1184) );
NAND2_X1 U900 ( .A1(n1019), .A2(n1223), .ZN(n1215) );
NAND4_X1 U901 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1092), .ZN(n1223) );
INV_X1 U902 ( .A(G900), .ZN(n1092) );
XOR2_X1 U903 ( .A(n1225), .B(n1186), .Z(G24) );
NAND4_X1 U904 ( .A1(n1226), .A2(n1193), .A3(n1183), .A4(n1066), .ZN(n1186) );
INV_X1 U905 ( .A(n1032), .ZN(n1193) );
NAND2_X1 U906 ( .A1(n1227), .A2(n1228), .ZN(n1032) );
XOR2_X1 U907 ( .A(n1229), .B(n1187), .Z(G21) );
NAND3_X1 U908 ( .A1(n1047), .A2(n1226), .A3(n1199), .ZN(n1187) );
NOR2_X1 U909 ( .A1(n1228), .A2(n1227), .ZN(n1199) );
XOR2_X1 U910 ( .A(G116), .B(n1191), .Z(G18) );
AND3_X1 U911 ( .A1(n1226), .A2(n1043), .A3(n1039), .ZN(n1191) );
NOR2_X1 U912 ( .A1(n1230), .A2(n1231), .ZN(n1043) );
XOR2_X1 U913 ( .A(G113), .B(n1190), .Z(G15) );
AND3_X1 U914 ( .A1(n1039), .A2(n1226), .A3(n1044), .ZN(n1190) );
AND2_X1 U915 ( .A1(n1231), .A2(n1183), .ZN(n1044) );
XNOR2_X1 U916 ( .A(n1230), .B(KEYINPUT49), .ZN(n1183) );
AND3_X1 U917 ( .A1(n1185), .A2(n1232), .A3(n1222), .ZN(n1226) );
INV_X1 U918 ( .A(n1023), .ZN(n1222) );
NAND2_X1 U919 ( .A1(n1050), .A2(n1233), .ZN(n1023) );
NOR2_X1 U920 ( .A1(n1068), .A2(n1228), .ZN(n1039) );
XOR2_X1 U921 ( .A(G110), .B(n1192), .Z(G12) );
AND3_X1 U922 ( .A1(n1040), .A2(n1194), .A3(n1047), .ZN(n1192) );
NOR2_X1 U923 ( .A1(n1066), .A2(n1230), .ZN(n1047) );
NAND2_X1 U924 ( .A1(n1064), .A2(n1065), .ZN(n1230) );
NAND2_X1 U925 ( .A1(n1234), .A2(n1235), .ZN(n1065) );
NAND2_X1 U926 ( .A1(n1122), .A2(n1113), .ZN(n1235) );
XOR2_X1 U927 ( .A(KEYINPUT0), .B(G475), .Z(n1234) );
NAND3_X1 U928 ( .A1(n1122), .A2(n1113), .A3(n1236), .ZN(n1064) );
XOR2_X1 U929 ( .A(n1124), .B(KEYINPUT0), .Z(n1236) );
INV_X1 U930 ( .A(G475), .ZN(n1124) );
XNOR2_X1 U931 ( .A(n1237), .B(n1238), .ZN(n1122) );
XOR2_X1 U932 ( .A(n1239), .B(n1240), .Z(n1238) );
XOR2_X1 U933 ( .A(G113), .B(G104), .Z(n1240) );
XOR2_X1 U934 ( .A(KEYINPUT61), .B(G122), .Z(n1239) );
XOR2_X1 U935 ( .A(n1241), .B(n1242), .Z(n1237) );
INV_X1 U936 ( .A(n1084), .ZN(n1242) );
XOR2_X1 U937 ( .A(n1210), .B(n1243), .Z(n1084) );
INV_X1 U938 ( .A(G131), .ZN(n1210) );
XNOR2_X1 U939 ( .A(n1244), .B(n1245), .ZN(n1241) );
NAND2_X1 U940 ( .A1(n1246), .A2(G214), .ZN(n1244) );
INV_X1 U941 ( .A(n1231), .ZN(n1066) );
XOR2_X1 U942 ( .A(n1247), .B(G478), .Z(n1231) );
NAND2_X1 U943 ( .A1(n1115), .A2(n1113), .ZN(n1247) );
XNOR2_X1 U944 ( .A(n1248), .B(n1249), .ZN(n1115) );
NOR2_X1 U945 ( .A1(n1250), .A2(n1251), .ZN(n1249) );
NOR2_X1 U946 ( .A1(n1252), .A2(n1253), .ZN(n1251) );
INV_X1 U947 ( .A(n1254), .ZN(n1253) );
NOR2_X1 U948 ( .A1(KEYINPUT48), .A2(n1255), .ZN(n1252) );
NOR2_X1 U949 ( .A1(KEYINPUT13), .A2(n1256), .ZN(n1255) );
NOR2_X1 U950 ( .A1(n1257), .A2(n1258), .ZN(n1250) );
NOR2_X1 U951 ( .A1(n1259), .A2(KEYINPUT13), .ZN(n1258) );
NOR2_X1 U952 ( .A1(KEYINPUT48), .A2(n1254), .ZN(n1259) );
XOR2_X1 U953 ( .A(n1260), .B(n1261), .Z(n1254) );
XOR2_X1 U954 ( .A(G143), .B(G134), .Z(n1261) );
NAND2_X1 U955 ( .A1(KEYINPUT23), .A2(n1262), .ZN(n1260) );
INV_X1 U956 ( .A(n1256), .ZN(n1257) );
NAND2_X1 U957 ( .A1(n1263), .A2(n1264), .ZN(n1256) );
NAND2_X1 U958 ( .A1(n1265), .A2(G107), .ZN(n1264) );
XOR2_X1 U959 ( .A(n1266), .B(KEYINPUT62), .Z(n1263) );
OR2_X1 U960 ( .A1(n1265), .A2(G107), .ZN(n1266) );
XOR2_X1 U961 ( .A(n1267), .B(n1268), .Z(n1265) );
NOR2_X1 U962 ( .A1(KEYINPUT59), .A2(G116), .ZN(n1268) );
XOR2_X1 U963 ( .A(n1225), .B(KEYINPUT32), .Z(n1267) );
INV_X1 U964 ( .A(G122), .ZN(n1225) );
NAND3_X1 U965 ( .A1(G234), .A2(n1088), .A3(G217), .ZN(n1248) );
AND3_X1 U966 ( .A1(n1049), .A2(n1232), .A3(n1185), .ZN(n1194) );
INV_X1 U967 ( .A(n1031), .ZN(n1185) );
NAND2_X1 U968 ( .A1(n1034), .A2(n1216), .ZN(n1031) );
NAND2_X1 U969 ( .A1(G214), .A2(n1269), .ZN(n1216) );
XOR2_X1 U970 ( .A(n1052), .B(KEYINPUT20), .Z(n1034) );
XNOR2_X1 U971 ( .A(n1270), .B(n1171), .ZN(n1052) );
NAND2_X1 U972 ( .A1(G210), .A2(n1269), .ZN(n1171) );
NAND2_X1 U973 ( .A1(n1271), .A2(n1113), .ZN(n1269) );
INV_X1 U974 ( .A(G237), .ZN(n1271) );
NAND2_X1 U975 ( .A1(n1272), .A2(n1113), .ZN(n1270) );
XNOR2_X1 U976 ( .A(n1273), .B(n1198), .ZN(n1272) );
XNOR2_X1 U977 ( .A(n1144), .B(G125), .ZN(n1198) );
XNOR2_X1 U978 ( .A(n1197), .B(n1169), .ZN(n1273) );
NOR2_X1 U979 ( .A1(n1105), .A2(G953), .ZN(n1169) );
INV_X1 U980 ( .A(G224), .ZN(n1105) );
XOR2_X1 U981 ( .A(n1274), .B(n1102), .Z(n1197) );
XOR2_X1 U982 ( .A(n1275), .B(n1276), .Z(n1102) );
XOR2_X1 U983 ( .A(KEYINPUT11), .B(n1159), .Z(n1276) );
NAND2_X1 U984 ( .A1(n1277), .A2(n1278), .ZN(n1275) );
NAND2_X1 U985 ( .A1(n1279), .A2(G119), .ZN(n1278) );
NAND2_X1 U986 ( .A1(n1280), .A2(n1229), .ZN(n1277) );
INV_X1 U987 ( .A(G119), .ZN(n1229) );
XNOR2_X1 U988 ( .A(n1279), .B(KEYINPUT7), .ZN(n1280) );
NAND2_X1 U989 ( .A1(KEYINPUT15), .A2(n1103), .ZN(n1274) );
XNOR2_X1 U990 ( .A(G110), .B(G122), .ZN(n1103) );
NAND2_X1 U991 ( .A1(n1019), .A2(n1281), .ZN(n1232) );
NAND4_X1 U992 ( .A1(G953), .A2(G902), .A3(n1224), .A4(n1101), .ZN(n1281) );
INV_X1 U993 ( .A(G898), .ZN(n1101) );
NAND3_X1 U994 ( .A1(n1224), .A2(n1088), .A3(n1282), .ZN(n1019) );
XNOR2_X1 U995 ( .A(G952), .B(KEYINPUT24), .ZN(n1282) );
NAND2_X1 U996 ( .A1(G237), .A2(G234), .ZN(n1224) );
NOR2_X1 U997 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
INV_X1 U998 ( .A(n1233), .ZN(n1051) );
NAND2_X1 U999 ( .A1(G221), .A2(n1283), .ZN(n1233) );
XOR2_X1 U1000 ( .A(n1067), .B(n1284), .Z(n1050) );
XOR2_X1 U1001 ( .A(KEYINPUT51), .B(KEYINPUT22), .Z(n1284) );
XNOR2_X1 U1002 ( .A(n1285), .B(G469), .ZN(n1067) );
NAND2_X1 U1003 ( .A1(n1286), .A2(n1113), .ZN(n1285) );
XNOR2_X1 U1004 ( .A(n1160), .B(n1287), .ZN(n1286) );
XOR2_X1 U1005 ( .A(n1165), .B(n1288), .Z(n1287) );
NOR2_X1 U1006 ( .A1(KEYINPUT30), .A2(n1289), .ZN(n1288) );
XOR2_X1 U1007 ( .A(n1290), .B(n1291), .Z(n1289) );
XOR2_X1 U1008 ( .A(n1142), .B(n1159), .Z(n1291) );
INV_X1 U1009 ( .A(n1157), .ZN(n1159) );
XOR2_X1 U1010 ( .A(n1292), .B(n1293), .Z(n1157) );
XOR2_X1 U1011 ( .A(KEYINPUT33), .B(G107), .Z(n1293) );
XNOR2_X1 U1012 ( .A(G104), .B(G101), .ZN(n1292) );
XNOR2_X1 U1013 ( .A(n1086), .B(KEYINPUT46), .ZN(n1290) );
AND3_X1 U1014 ( .A1(n1294), .A2(n1295), .A3(n1296), .ZN(n1086) );
NAND2_X1 U1015 ( .A1(n1297), .A2(G128), .ZN(n1295) );
NAND2_X1 U1016 ( .A1(n1245), .A2(n1262), .ZN(n1294) );
XOR2_X1 U1017 ( .A(G143), .B(n1298), .Z(n1245) );
NOR2_X1 U1018 ( .A1(n1091), .A2(G953), .ZN(n1165) );
INV_X1 U1019 ( .A(G227), .ZN(n1091) );
XOR2_X1 U1020 ( .A(G110), .B(G140), .Z(n1160) );
AND2_X1 U1021 ( .A1(n1228), .A2(n1068), .ZN(n1040) );
INV_X1 U1022 ( .A(n1227), .ZN(n1068) );
XNOR2_X1 U1023 ( .A(n1299), .B(n1111), .ZN(n1227) );
NAND2_X1 U1024 ( .A1(G217), .A2(n1283), .ZN(n1111) );
NAND2_X1 U1025 ( .A1(G234), .A2(n1113), .ZN(n1283) );
NAND2_X1 U1026 ( .A1(n1300), .A2(n1113), .ZN(n1299) );
XOR2_X1 U1027 ( .A(KEYINPUT1), .B(n1109), .Z(n1300) );
XNOR2_X1 U1028 ( .A(n1301), .B(n1302), .ZN(n1109) );
XOR2_X1 U1029 ( .A(G110), .B(n1303), .Z(n1302) );
XOR2_X1 U1030 ( .A(G128), .B(G119), .Z(n1303) );
XOR2_X1 U1031 ( .A(n1304), .B(n1305), .Z(n1301) );
NOR2_X1 U1032 ( .A1(n1306), .A2(n1307), .ZN(n1305) );
XOR2_X1 U1033 ( .A(n1308), .B(KEYINPUT26), .Z(n1307) );
NAND2_X1 U1034 ( .A1(G146), .A2(n1243), .ZN(n1308) );
NOR2_X1 U1035 ( .A1(n1309), .A2(n1243), .ZN(n1306) );
XOR2_X1 U1036 ( .A(G125), .B(G140), .Z(n1243) );
XOR2_X1 U1037 ( .A(n1298), .B(KEYINPUT17), .Z(n1309) );
NAND2_X1 U1038 ( .A1(n1310), .A2(n1311), .ZN(n1304) );
NAND2_X1 U1039 ( .A1(n1312), .A2(n1087), .ZN(n1311) );
XOR2_X1 U1040 ( .A(KEYINPUT12), .B(n1313), .Z(n1310) );
NOR2_X1 U1041 ( .A1(n1087), .A2(n1312), .ZN(n1313) );
NAND3_X1 U1042 ( .A1(G234), .A2(n1088), .A3(G221), .ZN(n1312) );
INV_X1 U1043 ( .A(G953), .ZN(n1088) );
XOR2_X1 U1044 ( .A(n1059), .B(G472), .Z(n1228) );
NAND2_X1 U1045 ( .A1(n1314), .A2(n1113), .ZN(n1059) );
INV_X1 U1046 ( .A(G902), .ZN(n1113) );
XOR2_X1 U1047 ( .A(n1315), .B(n1316), .Z(n1314) );
XNOR2_X1 U1048 ( .A(n1144), .B(n1317), .ZN(n1316) );
XNOR2_X1 U1049 ( .A(G101), .B(KEYINPUT4), .ZN(n1317) );
AND3_X1 U1050 ( .A1(n1318), .A2(n1319), .A3(n1296), .ZN(n1144) );
NAND3_X1 U1051 ( .A1(G128), .A2(n1298), .A3(G143), .ZN(n1296) );
NAND2_X1 U1052 ( .A1(n1320), .A2(G128), .ZN(n1319) );
XNOR2_X1 U1053 ( .A(n1297), .B(KEYINPUT31), .ZN(n1320) );
NAND3_X1 U1054 ( .A1(n1321), .A2(n1322), .A3(n1262), .ZN(n1318) );
INV_X1 U1055 ( .A(G128), .ZN(n1262) );
NAND2_X1 U1056 ( .A1(G143), .A2(n1298), .ZN(n1322) );
XOR2_X1 U1057 ( .A(KEYINPUT31), .B(n1297), .Z(n1321) );
NOR2_X1 U1058 ( .A1(n1298), .A2(G143), .ZN(n1297) );
INV_X1 U1059 ( .A(G146), .ZN(n1298) );
XOR2_X1 U1060 ( .A(n1323), .B(n1139), .Z(n1315) );
XOR2_X1 U1061 ( .A(G119), .B(n1279), .Z(n1139) );
XNOR2_X1 U1062 ( .A(n1324), .B(G116), .ZN(n1279) );
INV_X1 U1063 ( .A(G113), .ZN(n1324) );
XOR2_X1 U1064 ( .A(n1147), .B(n1142), .Z(n1323) );
INV_X1 U1065 ( .A(n1145), .ZN(n1142) );
XOR2_X1 U1066 ( .A(n1325), .B(n1326), .Z(n1145) );
NOR2_X1 U1067 ( .A1(KEYINPUT50), .A2(G131), .ZN(n1326) );
XOR2_X1 U1068 ( .A(G134), .B(n1087), .Z(n1325) );
INV_X1 U1069 ( .A(G137), .ZN(n1087) );
NAND2_X1 U1070 ( .A1(n1246), .A2(G210), .ZN(n1147) );
NOR2_X1 U1071 ( .A1(G953), .A2(G237), .ZN(n1246) );
endmodule


