//Key = 0100010111111000111110110010011100110101000101100110001010100000


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
n1414, n1415;

XNOR2_X1 U766 ( .A(G107), .B(n1074), .ZN(G9) );
NAND2_X1 U767 ( .A1(KEYINPUT39), .A2(n1075), .ZN(n1074) );
NOR2_X1 U768 ( .A1(n1076), .A2(n1077), .ZN(G75) );
NOR4_X1 U769 ( .A1(n1078), .A2(n1079), .A3(G953), .A4(n1080), .ZN(n1077) );
NOR3_X1 U770 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1079) );
NOR2_X1 U771 ( .A1(n1084), .A2(n1085), .ZN(n1082) );
NOR2_X1 U772 ( .A1(n1086), .A2(n1087), .ZN(n1084) );
NAND3_X1 U773 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1078) );
NAND2_X1 U774 ( .A1(KEYINPUT63), .A2(n1091), .ZN(n1089) );
NAND3_X1 U775 ( .A1(n1092), .A2(n1093), .A3(n1094), .ZN(n1091) );
NAND2_X1 U776 ( .A1(n1092), .A2(n1095), .ZN(n1088) );
NAND3_X1 U777 ( .A1(n1096), .A2(n1097), .A3(n1098), .ZN(n1095) );
XOR2_X1 U778 ( .A(n1099), .B(KEYINPUT13), .Z(n1098) );
NAND2_X1 U779 ( .A1(n1094), .A2(n1100), .ZN(n1099) );
NAND4_X1 U780 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1097) );
NOR2_X1 U781 ( .A1(n1083), .A2(n1105), .ZN(n1104) );
NAND2_X1 U782 ( .A1(n1106), .A2(n1107), .ZN(n1103) );
NAND3_X1 U783 ( .A1(n1108), .A2(n1109), .A3(n1110), .ZN(n1102) );
NAND2_X1 U784 ( .A1(n1111), .A2(n1112), .ZN(n1101) );
OR3_X1 U785 ( .A1(n1113), .A2(KEYINPUT63), .A3(n1081), .ZN(n1096) );
INV_X1 U786 ( .A(n1094), .ZN(n1081) );
NOR3_X1 U787 ( .A1(n1111), .A2(n1112), .A3(n1105), .ZN(n1094) );
NAND2_X1 U788 ( .A1(n1114), .A2(n1115), .ZN(n1111) );
NOR3_X1 U789 ( .A1(n1080), .A2(G953), .A3(G952), .ZN(n1076) );
AND4_X1 U790 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1080) );
NOR4_X1 U791 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1119) );
XNOR2_X1 U792 ( .A(KEYINPUT28), .B(n1124), .ZN(n1123) );
XOR2_X1 U793 ( .A(G469), .B(n1125), .Z(n1122) );
NOR3_X1 U794 ( .A1(n1126), .A2(n1106), .A3(n1127), .ZN(n1118) );
NAND2_X1 U795 ( .A1(n1128), .A2(n1129), .ZN(n1117) );
XOR2_X1 U796 ( .A(n1130), .B(n1131), .Z(n1116) );
XNOR2_X1 U797 ( .A(n1132), .B(G475), .ZN(n1131) );
XNOR2_X1 U798 ( .A(KEYINPUT50), .B(KEYINPUT36), .ZN(n1130) );
NAND2_X1 U799 ( .A1(n1133), .A2(n1134), .ZN(G72) );
NAND2_X1 U800 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
NAND2_X1 U801 ( .A1(n1137), .A2(n1138), .ZN(n1136) );
NAND2_X1 U802 ( .A1(G953), .A2(n1139), .ZN(n1138) );
NAND2_X1 U803 ( .A1(n1140), .A2(n1141), .ZN(n1133) );
INV_X1 U804 ( .A(n1135), .ZN(n1141) );
NOR3_X1 U805 ( .A1(KEYINPUT24), .A2(n1142), .A3(n1143), .ZN(n1135) );
NOR2_X1 U806 ( .A1(n1144), .A2(n1145), .ZN(n1143) );
XOR2_X1 U807 ( .A(KEYINPUT34), .B(n1146), .Z(n1145) );
NOR2_X1 U808 ( .A1(G953), .A2(n1147), .ZN(n1144) );
NOR3_X1 U809 ( .A1(n1147), .A2(G953), .A3(n1146), .ZN(n1142) );
AND2_X1 U810 ( .A1(n1148), .A2(n1137), .ZN(n1146) );
INV_X1 U811 ( .A(n1149), .ZN(n1137) );
XOR2_X1 U812 ( .A(n1150), .B(n1151), .Z(n1148) );
XOR2_X1 U813 ( .A(n1152), .B(n1153), .Z(n1151) );
XNOR2_X1 U814 ( .A(KEYINPUT45), .B(n1154), .ZN(n1153) );
NOR2_X1 U815 ( .A1(G140), .A2(KEYINPUT0), .ZN(n1152) );
XOR2_X1 U816 ( .A(n1155), .B(n1156), .Z(n1150) );
NAND2_X1 U817 ( .A1(KEYINPUT18), .A2(n1157), .ZN(n1155) );
INV_X1 U818 ( .A(n1158), .ZN(n1147) );
NAND2_X1 U819 ( .A1(G953), .A2(n1159), .ZN(n1140) );
NAND2_X1 U820 ( .A1(G900), .A2(G227), .ZN(n1159) );
XOR2_X1 U821 ( .A(n1160), .B(n1161), .Z(G69) );
NOR2_X1 U822 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
AND2_X1 U823 ( .A1(G224), .A2(G898), .ZN(n1162) );
NAND2_X1 U824 ( .A1(n1164), .A2(n1165), .ZN(n1160) );
NAND2_X1 U825 ( .A1(n1166), .A2(n1163), .ZN(n1165) );
XOR2_X1 U826 ( .A(n1167), .B(n1168), .Z(n1166) );
NAND3_X1 U827 ( .A1(G898), .A2(n1168), .A3(G953), .ZN(n1164) );
XNOR2_X1 U828 ( .A(n1169), .B(n1170), .ZN(n1168) );
XOR2_X1 U829 ( .A(n1171), .B(n1172), .Z(n1169) );
NOR2_X1 U830 ( .A1(n1173), .A2(n1174), .ZN(G66) );
XOR2_X1 U831 ( .A(n1175), .B(n1176), .Z(n1174) );
NAND2_X1 U832 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
NOR2_X1 U833 ( .A1(n1173), .A2(n1179), .ZN(G63) );
XOR2_X1 U834 ( .A(n1180), .B(n1181), .Z(n1179) );
NAND2_X1 U835 ( .A1(n1177), .A2(G478), .ZN(n1181) );
NOR2_X1 U836 ( .A1(n1173), .A2(n1182), .ZN(G60) );
NOR3_X1 U837 ( .A1(n1132), .A2(n1183), .A3(n1184), .ZN(n1182) );
AND3_X1 U838 ( .A1(n1185), .A2(G475), .A3(n1177), .ZN(n1184) );
NOR2_X1 U839 ( .A1(n1186), .A2(n1185), .ZN(n1183) );
NOR2_X1 U840 ( .A1(n1090), .A2(n1187), .ZN(n1186) );
INV_X1 U841 ( .A(G475), .ZN(n1187) );
XNOR2_X1 U842 ( .A(G104), .B(n1188), .ZN(G6) );
NOR2_X1 U843 ( .A1(n1173), .A2(n1189), .ZN(G57) );
XOR2_X1 U844 ( .A(n1190), .B(n1191), .Z(n1189) );
XNOR2_X1 U845 ( .A(n1192), .B(n1193), .ZN(n1191) );
XOR2_X1 U846 ( .A(n1194), .B(n1195), .Z(n1190) );
XNOR2_X1 U847 ( .A(n1196), .B(KEYINPUT48), .ZN(n1195) );
NAND2_X1 U848 ( .A1(KEYINPUT22), .A2(n1197), .ZN(n1196) );
NAND2_X1 U849 ( .A1(n1177), .A2(G472), .ZN(n1194) );
NOR2_X1 U850 ( .A1(n1173), .A2(n1198), .ZN(G54) );
XOR2_X1 U851 ( .A(n1199), .B(n1200), .Z(n1198) );
XOR2_X1 U852 ( .A(n1201), .B(n1202), .Z(n1200) );
XNOR2_X1 U853 ( .A(n1157), .B(n1203), .ZN(n1202) );
INV_X1 U854 ( .A(n1204), .ZN(n1157) );
XNOR2_X1 U855 ( .A(n1205), .B(n1156), .ZN(n1201) );
XOR2_X1 U856 ( .A(n1206), .B(n1207), .Z(n1199) );
XOR2_X1 U857 ( .A(KEYINPUT58), .B(KEYINPUT31), .Z(n1207) );
XOR2_X1 U858 ( .A(n1208), .B(n1209), .Z(n1206) );
NAND2_X1 U859 ( .A1(n1177), .A2(G469), .ZN(n1208) );
NOR2_X1 U860 ( .A1(n1173), .A2(n1210), .ZN(G51) );
XOR2_X1 U861 ( .A(n1211), .B(n1212), .Z(n1210) );
XOR2_X1 U862 ( .A(n1213), .B(n1214), .Z(n1212) );
NOR3_X1 U863 ( .A1(n1129), .A2(n1215), .A3(n1216), .ZN(n1214) );
NOR2_X1 U864 ( .A1(KEYINPUT46), .A2(n1217), .ZN(n1216) );
NOR2_X1 U865 ( .A1(n1090), .A2(G902), .ZN(n1217) );
NOR2_X1 U866 ( .A1(n1177), .A2(n1218), .ZN(n1215) );
INV_X1 U867 ( .A(KEYINPUT46), .ZN(n1218) );
NOR2_X1 U868 ( .A1(n1219), .A2(n1090), .ZN(n1177) );
NOR2_X1 U869 ( .A1(n1167), .A2(n1158), .ZN(n1090) );
NAND4_X1 U870 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(n1158) );
NOR4_X1 U871 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
INV_X1 U872 ( .A(n1228), .ZN(n1227) );
INV_X1 U873 ( .A(n1229), .ZN(n1224) );
NOR3_X1 U874 ( .A1(n1230), .A2(n1231), .A3(n1232), .ZN(n1222) );
NOR3_X1 U875 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1232) );
INV_X1 U876 ( .A(KEYINPUT59), .ZN(n1233) );
NOR2_X1 U877 ( .A1(KEYINPUT59), .A2(n1236), .ZN(n1231) );
NOR2_X1 U878 ( .A1(n1237), .A2(n1238), .ZN(n1230) );
INV_X1 U879 ( .A(n1092), .ZN(n1237) );
NAND4_X1 U880 ( .A1(n1239), .A2(n1188), .A3(n1240), .A4(n1241), .ZN(n1167) );
NOR4_X1 U881 ( .A1(n1242), .A2(n1243), .A3(n1075), .A4(n1244), .ZN(n1241) );
INV_X1 U882 ( .A(n1245), .ZN(n1244) );
NOR3_X1 U883 ( .A1(n1113), .A2(n1107), .A3(n1246), .ZN(n1075) );
INV_X1 U884 ( .A(n1114), .ZN(n1107) );
NAND2_X1 U885 ( .A1(n1085), .A2(n1247), .ZN(n1240) );
NAND2_X1 U886 ( .A1(n1248), .A2(n1249), .ZN(n1247) );
NAND3_X1 U887 ( .A1(n1250), .A2(n1251), .A3(n1252), .ZN(n1249) );
XNOR2_X1 U888 ( .A(n1253), .B(KEYINPUT10), .ZN(n1252) );
XOR2_X1 U889 ( .A(KEYINPUT43), .B(n1254), .Z(n1248) );
NAND3_X1 U890 ( .A1(n1255), .A2(n1114), .A3(n1100), .ZN(n1188) );
NAND3_X1 U891 ( .A1(n1250), .A2(n1255), .A3(n1256), .ZN(n1239) );
INV_X1 U892 ( .A(n1246), .ZN(n1255) );
NOR2_X1 U893 ( .A1(KEYINPUT32), .A2(n1257), .ZN(n1213) );
XOR2_X1 U894 ( .A(KEYINPUT49), .B(n1258), .Z(n1257) );
NOR2_X1 U895 ( .A1(n1163), .A2(G952), .ZN(n1173) );
XNOR2_X1 U896 ( .A(G146), .B(n1221), .ZN(G48) );
NAND4_X1 U897 ( .A1(n1259), .A2(n1253), .A3(n1100), .A4(n1085), .ZN(n1221) );
XNOR2_X1 U898 ( .A(G143), .B(n1220), .ZN(G45) );
NAND3_X1 U899 ( .A1(n1260), .A2(n1261), .A3(n1259), .ZN(n1220) );
XNOR2_X1 U900 ( .A(G140), .B(n1228), .ZN(G42) );
NAND4_X1 U901 ( .A1(n1259), .A2(n1092), .A3(n1256), .A4(n1100), .ZN(n1228) );
NAND2_X1 U902 ( .A1(n1262), .A2(n1263), .ZN(G39) );
OR2_X1 U903 ( .A1(n1264), .A2(G137), .ZN(n1263) );
XOR2_X1 U904 ( .A(n1265), .B(KEYINPUT42), .Z(n1262) );
NAND2_X1 U905 ( .A1(G137), .A2(n1264), .ZN(n1265) );
NAND2_X1 U906 ( .A1(n1266), .A2(n1092), .ZN(n1264) );
XOR2_X1 U907 ( .A(n1238), .B(KEYINPUT54), .Z(n1266) );
NAND2_X1 U908 ( .A1(n1267), .A2(n1259), .ZN(n1238) );
XOR2_X1 U909 ( .A(G134), .B(n1226), .Z(G36) );
AND2_X1 U910 ( .A1(n1268), .A2(n1093), .ZN(n1226) );
INV_X1 U911 ( .A(n1113), .ZN(n1093) );
XOR2_X1 U912 ( .A(n1269), .B(n1225), .Z(G33) );
AND2_X1 U913 ( .A1(n1268), .A2(n1100), .ZN(n1225) );
AND3_X1 U914 ( .A1(n1092), .A2(n1261), .A3(n1259), .ZN(n1268) );
AND3_X1 U915 ( .A1(n1112), .A2(n1115), .A3(n1270), .ZN(n1259) );
NOR2_X1 U916 ( .A1(n1086), .A2(n1126), .ZN(n1092) );
INV_X1 U917 ( .A(n1271), .ZN(n1086) );
XNOR2_X1 U918 ( .A(G131), .B(KEYINPUT20), .ZN(n1269) );
XNOR2_X1 U919 ( .A(G128), .B(n1229), .ZN(G30) );
NAND4_X1 U920 ( .A1(n1272), .A2(n1270), .A3(n1085), .A4(n1273), .ZN(n1229) );
NOR2_X1 U921 ( .A1(n1113), .A2(n1274), .ZN(n1273) );
XNOR2_X1 U922 ( .A(n1243), .B(n1275), .ZN(G3) );
NOR2_X1 U923 ( .A1(G101), .A2(KEYINPUT33), .ZN(n1275) );
NOR3_X1 U924 ( .A1(n1108), .A2(n1246), .A3(n1083), .ZN(n1243) );
NAND2_X1 U925 ( .A1(n1276), .A2(n1277), .ZN(G27) );
NAND3_X1 U926 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
INV_X1 U927 ( .A(n1236), .ZN(n1280) );
NAND2_X1 U928 ( .A1(KEYINPUT55), .A2(n1154), .ZN(n1279) );
NAND2_X1 U929 ( .A1(n1281), .A2(G125), .ZN(n1278) );
NAND3_X1 U930 ( .A1(G125), .A2(n1282), .A3(n1281), .ZN(n1276) );
XNOR2_X1 U931 ( .A(KEYINPUT62), .B(KEYINPUT41), .ZN(n1281) );
OR2_X1 U932 ( .A1(n1236), .A2(KEYINPUT55), .ZN(n1282) );
NAND2_X1 U933 ( .A1(n1234), .A2(n1085), .ZN(n1236) );
AND4_X1 U934 ( .A1(n1256), .A2(n1100), .A3(n1110), .A4(n1270), .ZN(n1234) );
NAND2_X1 U935 ( .A1(n1105), .A2(n1283), .ZN(n1270) );
NAND3_X1 U936 ( .A1(G902), .A2(n1284), .A3(n1149), .ZN(n1283) );
NOR2_X1 U937 ( .A1(n1163), .A2(G900), .ZN(n1149) );
XNOR2_X1 U938 ( .A(G122), .B(n1245), .ZN(G24) );
NAND3_X1 U939 ( .A1(n1251), .A2(n1114), .A3(n1260), .ZN(n1245) );
AND3_X1 U940 ( .A1(n1085), .A2(n1121), .A3(n1285), .ZN(n1260) );
NOR2_X1 U941 ( .A1(n1120), .A2(n1286), .ZN(n1114) );
XOR2_X1 U942 ( .A(G119), .B(n1287), .Z(G21) );
NOR2_X1 U943 ( .A1(n1235), .A2(n1288), .ZN(n1287) );
XOR2_X1 U944 ( .A(KEYINPUT19), .B(n1289), .Z(n1288) );
AND2_X1 U945 ( .A1(n1251), .A2(n1267), .ZN(n1289) );
NOR2_X1 U946 ( .A1(n1274), .A2(n1083), .ZN(n1267) );
INV_X1 U947 ( .A(n1253), .ZN(n1274) );
NOR2_X1 U948 ( .A1(n1124), .A2(n1290), .ZN(n1253) );
XOR2_X1 U949 ( .A(G116), .B(n1242), .Z(G18) );
NOR4_X1 U950 ( .A1(n1108), .A2(n1291), .A3(n1113), .A4(n1235), .ZN(n1242) );
INV_X1 U951 ( .A(n1085), .ZN(n1235) );
NAND2_X1 U952 ( .A1(n1292), .A2(n1121), .ZN(n1113) );
INV_X1 U953 ( .A(n1261), .ZN(n1108) );
XNOR2_X1 U954 ( .A(G113), .B(n1293), .ZN(G15) );
NAND2_X1 U955 ( .A1(n1254), .A2(n1085), .ZN(n1293) );
AND3_X1 U956 ( .A1(n1261), .A2(n1251), .A3(n1100), .ZN(n1254) );
AND2_X1 U957 ( .A1(n1294), .A2(n1285), .ZN(n1100) );
INV_X1 U958 ( .A(n1292), .ZN(n1285) );
INV_X1 U959 ( .A(n1291), .ZN(n1251) );
NAND2_X1 U960 ( .A1(n1110), .A2(n1295), .ZN(n1291) );
NOR2_X1 U961 ( .A1(n1112), .A2(n1106), .ZN(n1110) );
INV_X1 U962 ( .A(n1115), .ZN(n1106) );
NOR2_X1 U963 ( .A1(n1286), .A2(n1290), .ZN(n1261) );
INV_X1 U964 ( .A(n1120), .ZN(n1290) );
XNOR2_X1 U965 ( .A(n1296), .B(n1297), .ZN(G12) );
NOR3_X1 U966 ( .A1(n1109), .A2(n1298), .A3(n1246), .ZN(n1297) );
NAND3_X1 U967 ( .A1(n1272), .A2(n1295), .A3(n1085), .ZN(n1246) );
NOR2_X1 U968 ( .A1(n1126), .A2(n1271), .ZN(n1085) );
NOR2_X1 U969 ( .A1(n1299), .A2(n1127), .ZN(n1271) );
NOR2_X1 U970 ( .A1(n1129), .A2(n1128), .ZN(n1127) );
AND2_X1 U971 ( .A1(n1300), .A2(n1129), .ZN(n1299) );
NAND2_X1 U972 ( .A1(G210), .A2(n1301), .ZN(n1129) );
XNOR2_X1 U973 ( .A(n1128), .B(KEYINPUT56), .ZN(n1300) );
AND2_X1 U974 ( .A1(n1302), .A2(n1219), .ZN(n1128) );
XOR2_X1 U975 ( .A(n1258), .B(n1303), .Z(n1302) );
XNOR2_X1 U976 ( .A(n1304), .B(KEYINPUT26), .ZN(n1303) );
NAND2_X1 U977 ( .A1(KEYINPUT29), .A2(n1211), .ZN(n1304) );
XNOR2_X1 U978 ( .A(n1305), .B(n1172), .ZN(n1211) );
XNOR2_X1 U979 ( .A(n1306), .B(G122), .ZN(n1172) );
NAND2_X1 U980 ( .A1(KEYINPUT23), .A2(n1296), .ZN(n1306) );
NAND2_X1 U981 ( .A1(n1307), .A2(n1308), .ZN(n1305) );
NAND2_X1 U982 ( .A1(n1170), .A2(n1309), .ZN(n1308) );
XOR2_X1 U983 ( .A(n1310), .B(KEYINPUT47), .Z(n1307) );
OR2_X1 U984 ( .A1(n1309), .A2(n1170), .ZN(n1310) );
XNOR2_X1 U985 ( .A(n1311), .B(n1312), .ZN(n1170) );
NOR2_X1 U986 ( .A1(KEYINPUT15), .A2(n1313), .ZN(n1312) );
XNOR2_X1 U987 ( .A(n1171), .B(KEYINPUT53), .ZN(n1309) );
XOR2_X1 U988 ( .A(n1314), .B(n1315), .Z(n1171) );
NAND2_X1 U989 ( .A1(KEYINPUT8), .A2(n1316), .ZN(n1314) );
XNOR2_X1 U990 ( .A(n1317), .B(n1318), .ZN(n1258) );
XNOR2_X1 U991 ( .A(G125), .B(n1319), .ZN(n1318) );
NAND2_X1 U992 ( .A1(G224), .A2(n1163), .ZN(n1317) );
INV_X1 U993 ( .A(n1087), .ZN(n1126) );
NAND2_X1 U994 ( .A1(G214), .A2(n1301), .ZN(n1087) );
NAND2_X1 U995 ( .A1(n1320), .A2(n1219), .ZN(n1301) );
INV_X1 U996 ( .A(G237), .ZN(n1320) );
NAND2_X1 U997 ( .A1(n1105), .A2(n1321), .ZN(n1295) );
NAND4_X1 U998 ( .A1(G953), .A2(G902), .A3(n1284), .A4(n1322), .ZN(n1321) );
INV_X1 U999 ( .A(G898), .ZN(n1322) );
NAND3_X1 U1000 ( .A1(n1284), .A2(n1163), .A3(G952), .ZN(n1105) );
NAND2_X1 U1001 ( .A1(G237), .A2(G234), .ZN(n1284) );
XOR2_X1 U1002 ( .A(n1323), .B(KEYINPUT37), .Z(n1272) );
NAND2_X1 U1003 ( .A1(n1112), .A2(n1115), .ZN(n1323) );
NAND2_X1 U1004 ( .A1(G221), .A2(n1324), .ZN(n1115) );
NAND3_X1 U1005 ( .A1(n1325), .A2(n1326), .A3(n1327), .ZN(n1112) );
NAND2_X1 U1006 ( .A1(n1125), .A2(n1328), .ZN(n1327) );
OR3_X1 U1007 ( .A1(n1328), .A2(n1125), .A3(n1329), .ZN(n1326) );
INV_X1 U1008 ( .A(KEYINPUT12), .ZN(n1328) );
NAND2_X1 U1009 ( .A1(n1329), .A2(n1330), .ZN(n1325) );
NAND2_X1 U1010 ( .A1(KEYINPUT12), .A2(n1331), .ZN(n1330) );
XOR2_X1 U1011 ( .A(KEYINPUT11), .B(n1125), .Z(n1331) );
AND2_X1 U1012 ( .A1(n1332), .A2(n1219), .ZN(n1125) );
XNOR2_X1 U1013 ( .A(n1204), .B(n1333), .ZN(n1332) );
XNOR2_X1 U1014 ( .A(n1334), .B(n1335), .ZN(n1333) );
NOR2_X1 U1015 ( .A1(KEYINPUT14), .A2(n1336), .ZN(n1335) );
XOR2_X1 U1016 ( .A(n1337), .B(n1156), .Z(n1336) );
XNOR2_X1 U1017 ( .A(n1338), .B(n1339), .ZN(n1156) );
NOR2_X1 U1018 ( .A1(G146), .A2(KEYINPUT3), .ZN(n1339) );
XNOR2_X1 U1019 ( .A(G128), .B(G143), .ZN(n1338) );
NOR2_X1 U1020 ( .A1(KEYINPUT40), .A2(n1205), .ZN(n1337) );
XOR2_X1 U1021 ( .A(n1315), .B(n1340), .Z(n1205) );
XNOR2_X1 U1022 ( .A(KEYINPUT27), .B(n1316), .ZN(n1340) );
XOR2_X1 U1023 ( .A(G104), .B(n1341), .Z(n1315) );
XNOR2_X1 U1024 ( .A(KEYINPUT6), .B(n1342), .ZN(n1341) );
NAND2_X1 U1025 ( .A1(KEYINPUT35), .A2(n1343), .ZN(n1334) );
XNOR2_X1 U1026 ( .A(n1344), .B(n1203), .ZN(n1343) );
XNOR2_X1 U1027 ( .A(G110), .B(n1345), .ZN(n1203) );
INV_X1 U1028 ( .A(G140), .ZN(n1345) );
NAND2_X1 U1029 ( .A1(KEYINPUT30), .A2(n1209), .ZN(n1344) );
NOR2_X1 U1030 ( .A1(n1139), .A2(G953), .ZN(n1209) );
INV_X1 U1031 ( .A(G227), .ZN(n1139) );
XOR2_X1 U1032 ( .A(G469), .B(KEYINPUT5), .Z(n1329) );
XNOR2_X1 U1033 ( .A(n1250), .B(KEYINPUT60), .ZN(n1298) );
INV_X1 U1034 ( .A(n1083), .ZN(n1250) );
NAND2_X1 U1035 ( .A1(n1294), .A2(n1292), .ZN(n1083) );
XOR2_X1 U1036 ( .A(n1132), .B(n1346), .Z(n1292) );
NOR2_X1 U1037 ( .A1(G475), .A2(KEYINPUT57), .ZN(n1346) );
NOR2_X1 U1038 ( .A1(n1185), .A2(G902), .ZN(n1132) );
XOR2_X1 U1039 ( .A(n1347), .B(n1348), .Z(n1185) );
XOR2_X1 U1040 ( .A(n1349), .B(n1350), .Z(n1348) );
XOR2_X1 U1041 ( .A(G131), .B(G104), .Z(n1350) );
NOR2_X1 U1042 ( .A1(n1351), .A2(n1352), .ZN(n1349) );
XOR2_X1 U1043 ( .A(n1353), .B(KEYINPUT9), .Z(n1352) );
NAND2_X1 U1044 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
NAND2_X1 U1045 ( .A1(n1356), .A2(G214), .ZN(n1355) );
AND3_X1 U1046 ( .A1(n1356), .A2(G143), .A3(G214), .ZN(n1351) );
XOR2_X1 U1047 ( .A(n1357), .B(n1358), .Z(n1347) );
NOR2_X1 U1048 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
XOR2_X1 U1049 ( .A(KEYINPUT52), .B(n1361), .Z(n1360) );
NOR2_X1 U1050 ( .A1(G113), .A2(n1362), .ZN(n1361) );
NOR2_X1 U1051 ( .A1(G122), .A2(n1313), .ZN(n1359) );
INV_X1 U1052 ( .A(G113), .ZN(n1313) );
NAND2_X1 U1053 ( .A1(n1363), .A2(n1364), .ZN(n1357) );
NAND2_X1 U1054 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
NAND2_X1 U1055 ( .A1(KEYINPUT7), .A2(n1367), .ZN(n1366) );
NAND2_X1 U1056 ( .A1(n1368), .A2(n1369), .ZN(n1367) );
INV_X1 U1057 ( .A(n1370), .ZN(n1365) );
NAND2_X1 U1058 ( .A1(n1371), .A2(n1372), .ZN(n1363) );
NAND2_X1 U1059 ( .A1(n1369), .A2(n1373), .ZN(n1372) );
NAND2_X1 U1060 ( .A1(KEYINPUT7), .A2(n1370), .ZN(n1373) );
XOR2_X1 U1061 ( .A(G146), .B(KEYINPUT21), .Z(n1370) );
INV_X1 U1062 ( .A(KEYINPUT51), .ZN(n1369) );
INV_X1 U1063 ( .A(n1368), .ZN(n1371) );
XNOR2_X1 U1064 ( .A(KEYINPUT38), .B(n1121), .ZN(n1294) );
XNOR2_X1 U1065 ( .A(n1374), .B(G478), .ZN(n1121) );
NAND2_X1 U1066 ( .A1(n1219), .A2(n1180), .ZN(n1374) );
NAND2_X1 U1067 ( .A1(n1375), .A2(n1376), .ZN(n1180) );
NAND4_X1 U1068 ( .A1(n1377), .A2(G217), .A3(G234), .A4(n1163), .ZN(n1376) );
NAND2_X1 U1069 ( .A1(n1378), .A2(n1379), .ZN(n1375) );
NAND3_X1 U1070 ( .A1(G234), .A2(n1163), .A3(G217), .ZN(n1379) );
XNOR2_X1 U1071 ( .A(KEYINPUT4), .B(n1377), .ZN(n1378) );
XOR2_X1 U1072 ( .A(n1380), .B(n1381), .Z(n1377) );
XOR2_X1 U1073 ( .A(n1382), .B(n1383), .Z(n1381) );
NAND2_X1 U1074 ( .A1(KEYINPUT16), .A2(n1342), .ZN(n1383) );
INV_X1 U1075 ( .A(G107), .ZN(n1342) );
NAND2_X1 U1076 ( .A1(n1384), .A2(n1385), .ZN(n1382) );
OR2_X1 U1077 ( .A1(n1386), .A2(n1354), .ZN(n1385) );
XOR2_X1 U1078 ( .A(n1387), .B(KEYINPUT25), .Z(n1384) );
NAND2_X1 U1079 ( .A1(n1386), .A2(n1354), .ZN(n1387) );
XOR2_X1 U1080 ( .A(G128), .B(KEYINPUT61), .Z(n1386) );
XNOR2_X1 U1081 ( .A(G116), .B(n1388), .ZN(n1380) );
XNOR2_X1 U1082 ( .A(G134), .B(n1362), .ZN(n1388) );
INV_X1 U1083 ( .A(G122), .ZN(n1362) );
INV_X1 U1084 ( .A(n1256), .ZN(n1109) );
NOR2_X1 U1085 ( .A1(n1120), .A2(n1124), .ZN(n1256) );
INV_X1 U1086 ( .A(n1286), .ZN(n1124) );
XNOR2_X1 U1087 ( .A(n1389), .B(n1178), .ZN(n1286) );
AND2_X1 U1088 ( .A1(G217), .A2(n1324), .ZN(n1178) );
NAND2_X1 U1089 ( .A1(G234), .A2(n1219), .ZN(n1324) );
NAND2_X1 U1090 ( .A1(n1176), .A2(n1219), .ZN(n1389) );
XOR2_X1 U1091 ( .A(n1390), .B(n1391), .Z(n1176) );
XNOR2_X1 U1092 ( .A(n1392), .B(n1368), .ZN(n1391) );
XNOR2_X1 U1093 ( .A(G140), .B(n1154), .ZN(n1368) );
INV_X1 U1094 ( .A(G125), .ZN(n1154) );
NAND2_X1 U1095 ( .A1(n1393), .A2(KEYINPUT17), .ZN(n1392) );
XNOR2_X1 U1096 ( .A(G137), .B(n1394), .ZN(n1393) );
AND3_X1 U1097 ( .A1(G221), .A2(n1163), .A3(G234), .ZN(n1394) );
INV_X1 U1098 ( .A(G953), .ZN(n1163) );
XOR2_X1 U1099 ( .A(n1395), .B(G146), .Z(n1390) );
NAND2_X1 U1100 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
NAND2_X1 U1101 ( .A1(G110), .A2(n1398), .ZN(n1397) );
XOR2_X1 U1102 ( .A(KEYINPUT1), .B(n1399), .Z(n1396) );
NOR2_X1 U1103 ( .A1(G110), .A2(n1398), .ZN(n1399) );
XNOR2_X1 U1104 ( .A(n1400), .B(G119), .ZN(n1398) );
XNOR2_X1 U1105 ( .A(n1401), .B(G472), .ZN(n1120) );
NAND2_X1 U1106 ( .A1(n1402), .A2(n1219), .ZN(n1401) );
INV_X1 U1107 ( .A(G902), .ZN(n1219) );
XOR2_X1 U1108 ( .A(n1403), .B(n1404), .Z(n1402) );
XNOR2_X1 U1109 ( .A(n1193), .B(n1197), .ZN(n1404) );
XOR2_X1 U1110 ( .A(n1405), .B(n1316), .Z(n1197) );
INV_X1 U1111 ( .A(G101), .ZN(n1316) );
NAND2_X1 U1112 ( .A1(n1356), .A2(G210), .ZN(n1405) );
NOR2_X1 U1113 ( .A1(G953), .A2(G237), .ZN(n1356) );
XNOR2_X1 U1114 ( .A(G113), .B(n1311), .ZN(n1193) );
XOR2_X1 U1115 ( .A(G116), .B(G119), .Z(n1311) );
NAND2_X1 U1116 ( .A1(n1406), .A2(n1407), .ZN(n1403) );
NAND2_X1 U1117 ( .A1(n1192), .A2(n1408), .ZN(n1407) );
INV_X1 U1118 ( .A(KEYINPUT44), .ZN(n1408) );
XOR2_X1 U1119 ( .A(n1204), .B(n1409), .Z(n1192) );
NAND3_X1 U1120 ( .A1(n1409), .A2(n1204), .A3(KEYINPUT44), .ZN(n1406) );
XOR2_X1 U1121 ( .A(G131), .B(n1410), .Z(n1204) );
XOR2_X1 U1122 ( .A(G137), .B(G134), .Z(n1410) );
INV_X1 U1123 ( .A(n1319), .ZN(n1409) );
NAND2_X1 U1124 ( .A1(n1411), .A2(n1412), .ZN(n1319) );
NAND2_X1 U1125 ( .A1(G128), .A2(n1413), .ZN(n1412) );
XNOR2_X1 U1126 ( .A(G146), .B(n1354), .ZN(n1413) );
INV_X1 U1127 ( .A(G143), .ZN(n1354) );
XOR2_X1 U1128 ( .A(n1414), .B(KEYINPUT2), .Z(n1411) );
NAND2_X1 U1129 ( .A1(n1415), .A2(n1400), .ZN(n1414) );
INV_X1 U1130 ( .A(G128), .ZN(n1400) );
XNOR2_X1 U1131 ( .A(G146), .B(G143), .ZN(n1415) );
INV_X1 U1132 ( .A(G110), .ZN(n1296) );
endmodule


