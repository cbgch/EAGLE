//Key = 0101100110010000000000101101101010110001001011110001101110000100


module c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3,
G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT0, KEYINPUT1,
KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7,
KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13,
KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19,
KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25,
KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31,
KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43,
KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49,
KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55,
KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61,
KEYINPUT62, KEYINPUT63 );
input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT0,
KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27,
KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57,
KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
KEYINPUT63;
output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
wire   n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;

XNOR2_X1 U704 ( .A(G107), .B(n960), .ZN(G9) );
NOR2_X1 U705 ( .A1(n961), .A2(n962), .ZN(G75) );
NOR4_X1 U706 ( .A1(G953), .A2(n963), .A3(n964), .A4(n965), .ZN(n962) );
NOR2_X1 U707 ( .A1(n966), .A2(n967), .ZN(n964) );
NOR2_X1 U708 ( .A1(n968), .A2(n969), .ZN(n966) );
NOR2_X1 U709 ( .A1(n970), .A2(n971), .ZN(n969) );
INV_X1 U710 ( .A(n972), .ZN(n971) );
NOR2_X1 U711 ( .A1(n973), .A2(n974), .ZN(n970) );
NOR2_X1 U712 ( .A1(n975), .A2(n976), .ZN(n974) );
NOR2_X1 U713 ( .A1(n977), .A2(n978), .ZN(n975) );
NOR2_X1 U714 ( .A1(n979), .A2(n980), .ZN(n978) );
NOR2_X1 U715 ( .A1(n981), .A2(n982), .ZN(n979) );
NOR2_X1 U716 ( .A1(n983), .A2(n984), .ZN(n981) );
NOR2_X1 U717 ( .A1(n985), .A2(n986), .ZN(n977) );
NOR2_X1 U718 ( .A1(n987), .A2(n988), .ZN(n985) );
AND2_X1 U719 ( .A1(n989), .A2(n990), .ZN(n987) );
NOR3_X1 U720 ( .A1(n986), .A2(n991), .A3(n980), .ZN(n973) );
NOR2_X1 U721 ( .A1(n992), .A2(n993), .ZN(n991) );
XOR2_X1 U722 ( .A(KEYINPUT0), .B(n994), .Z(n993) );
NOR2_X1 U723 ( .A1(n995), .A2(n996), .ZN(n992) );
NOR4_X1 U724 ( .A1(n997), .A2(n980), .A3(n986), .A4(n976), .ZN(n968) );
INV_X1 U725 ( .A(n998), .ZN(n986) );
INV_X1 U726 ( .A(n999), .ZN(n980) );
NOR2_X1 U727 ( .A1(n1000), .A2(n1001), .ZN(n997) );
NOR3_X1 U728 ( .A1(n963), .A2(G953), .A3(G952), .ZN(n961) );
AND4_X1 U729 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n963) );
NOR3_X1 U730 ( .A1(n1006), .A2(n1007), .A3(n1008), .ZN(n1005) );
NOR2_X1 U731 ( .A1(n1009), .A2(n1010), .ZN(n1008) );
XOR2_X1 U732 ( .A(KEYINPUT54), .B(G478), .Z(n1010) );
NOR2_X1 U733 ( .A1(G902), .A2(n1011), .ZN(n1009) );
NOR2_X1 U734 ( .A1(G475), .A2(n1012), .ZN(n1007) );
NAND3_X1 U735 ( .A1(n984), .A2(n1013), .A3(n996), .ZN(n1006) );
NOR3_X1 U736 ( .A1(n1014), .A2(n1015), .A3(n989), .ZN(n1004) );
XOR2_X1 U737 ( .A(n1016), .B(G469), .Z(n1015) );
NAND2_X1 U738 ( .A1(KEYINPUT52), .A2(n1017), .ZN(n1016) );
XOR2_X1 U739 ( .A(n1018), .B(n1019), .Z(n1014) );
XOR2_X1 U740 ( .A(n1020), .B(KEYINPUT19), .Z(n1019) );
NAND2_X1 U741 ( .A1(KEYINPUT27), .A2(n1021), .ZN(n1018) );
XNOR2_X1 U742 ( .A(n1022), .B(n1023), .ZN(n1003) );
XOR2_X1 U743 ( .A(n1024), .B(KEYINPUT10), .Z(n1002) );
NAND2_X1 U744 ( .A1(n1012), .A2(n1025), .ZN(n1024) );
XNOR2_X1 U745 ( .A(KEYINPUT49), .B(n1026), .ZN(n1025) );
XNOR2_X1 U746 ( .A(n1027), .B(KEYINPUT14), .ZN(n1012) );
XOR2_X1 U747 ( .A(n1028), .B(n1029), .Z(G72) );
NOR2_X1 U748 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
XOR2_X1 U749 ( .A(n1032), .B(KEYINPUT51), .Z(n1030) );
NAND2_X1 U750 ( .A1(G900), .A2(G227), .ZN(n1032) );
NAND2_X1 U751 ( .A1(n1033), .A2(n1034), .ZN(n1028) );
NAND2_X1 U752 ( .A1(n1035), .A2(n1031), .ZN(n1034) );
XOR2_X1 U753 ( .A(n1036), .B(n1037), .Z(n1035) );
NAND3_X1 U754 ( .A1(n1038), .A2(n1039), .A3(n1040), .ZN(n1036) );
XOR2_X1 U755 ( .A(n1041), .B(KEYINPUT42), .Z(n1040) );
XNOR2_X1 U756 ( .A(KEYINPUT30), .B(n1042), .ZN(n1039) );
NAND3_X1 U757 ( .A1(G900), .A2(n1037), .A3(G953), .ZN(n1033) );
XNOR2_X1 U758 ( .A(n1043), .B(n1044), .ZN(n1037) );
XOR2_X1 U759 ( .A(n1045), .B(n1046), .Z(n1044) );
NOR2_X1 U760 ( .A1(KEYINPUT41), .A2(n1047), .ZN(n1045) );
XOR2_X1 U761 ( .A(n1048), .B(n1049), .Z(n1043) );
NOR2_X1 U762 ( .A1(KEYINPUT63), .A2(n1050), .ZN(n1049) );
XNOR2_X1 U763 ( .A(G131), .B(KEYINPUT22), .ZN(n1048) );
XOR2_X1 U764 ( .A(n1051), .B(n1052), .Z(G69) );
XOR2_X1 U765 ( .A(n1053), .B(n1054), .Z(n1052) );
NOR2_X1 U766 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
NOR2_X1 U767 ( .A1(G224), .A2(n1031), .ZN(n1056) );
NOR3_X1 U768 ( .A1(n1057), .A2(n1058), .A3(n1055), .ZN(n1053) );
XOR2_X1 U769 ( .A(n1059), .B(KEYINPUT46), .Z(n1057) );
NAND2_X1 U770 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
XOR2_X1 U771 ( .A(KEYINPUT29), .B(n1062), .Z(n1060) );
NAND3_X1 U772 ( .A1(KEYINPUT34), .A2(n1063), .A3(n1064), .ZN(n1051) );
XNOR2_X1 U773 ( .A(G953), .B(KEYINPUT57), .ZN(n1064) );
NAND2_X1 U774 ( .A1(n1065), .A2(n1066), .ZN(n1063) );
NOR2_X1 U775 ( .A1(n1067), .A2(n1068), .ZN(G66) );
XNOR2_X1 U776 ( .A(n1069), .B(n1070), .ZN(n1068) );
NOR2_X1 U777 ( .A1(n1071), .A2(n1072), .ZN(n1070) );
NOR2_X1 U778 ( .A1(n1067), .A2(n1073), .ZN(G63) );
XNOR2_X1 U779 ( .A(n1074), .B(n1075), .ZN(n1073) );
NAND2_X1 U780 ( .A1(KEYINPUT4), .A2(n1076), .ZN(n1074) );
NAND3_X1 U781 ( .A1(n1077), .A2(n965), .A3(G478), .ZN(n1076) );
XNOR2_X1 U782 ( .A(KEYINPUT6), .B(n1078), .ZN(n1077) );
NOR2_X1 U783 ( .A1(n1079), .A2(n1080), .ZN(G60) );
XOR2_X1 U784 ( .A(KEYINPUT37), .B(n1067), .Z(n1080) );
NOR3_X1 U785 ( .A1(n1081), .A2(n1082), .A3(n1083), .ZN(n1079) );
AND2_X1 U786 ( .A1(n1084), .A2(KEYINPUT38), .ZN(n1083) );
NOR2_X1 U787 ( .A1(KEYINPUT38), .A2(n1085), .ZN(n1082) );
NOR2_X1 U788 ( .A1(n1086), .A2(n1027), .ZN(n1085) );
NOR2_X1 U789 ( .A1(n1087), .A2(n1084), .ZN(n1086) );
AND3_X1 U790 ( .A1(KEYINPUT45), .A2(n965), .A3(G475), .ZN(n1087) );
NOR3_X1 U791 ( .A1(n1072), .A2(n1088), .A3(n1026), .ZN(n1081) );
NOR2_X1 U792 ( .A1(n1089), .A2(KEYINPUT38), .ZN(n1088) );
AND2_X1 U793 ( .A1(n1084), .A2(KEYINPUT45), .ZN(n1089) );
XNOR2_X1 U794 ( .A(G104), .B(n1090), .ZN(G6) );
NOR2_X1 U795 ( .A1(n1067), .A2(n1091), .ZN(G57) );
XOR2_X1 U796 ( .A(n1092), .B(n1093), .Z(n1091) );
XOR2_X1 U797 ( .A(n1094), .B(n1095), .Z(n1093) );
NOR2_X1 U798 ( .A1(KEYINPUT62), .A2(n1096), .ZN(n1095) );
NOR2_X1 U799 ( .A1(n1023), .A2(n1072), .ZN(n1094) );
INV_X1 U800 ( .A(G472), .ZN(n1023) );
XOR2_X1 U801 ( .A(n1097), .B(n1098), .Z(n1092) );
NOR2_X1 U802 ( .A1(n1067), .A2(n1099), .ZN(G54) );
XOR2_X1 U803 ( .A(n1100), .B(n1101), .Z(n1099) );
XNOR2_X1 U804 ( .A(n1050), .B(n1102), .ZN(n1101) );
XOR2_X1 U805 ( .A(n1103), .B(n1104), .Z(n1100) );
XOR2_X1 U806 ( .A(n1105), .B(n1106), .Z(n1103) );
NAND3_X1 U807 ( .A1(G469), .A2(n965), .A3(n1107), .ZN(n1105) );
XNOR2_X1 U808 ( .A(G902), .B(KEYINPUT7), .ZN(n1107) );
NOR2_X1 U809 ( .A1(n1067), .A2(n1108), .ZN(G51) );
XOR2_X1 U810 ( .A(n1109), .B(n1110), .Z(n1108) );
XOR2_X1 U811 ( .A(n1111), .B(n1112), .Z(n1110) );
NOR2_X1 U812 ( .A1(KEYINPUT23), .A2(n1113), .ZN(n1112) );
XOR2_X1 U813 ( .A(n1114), .B(n1115), .Z(n1113) );
XOR2_X1 U814 ( .A(n1116), .B(n1117), .Z(n1115) );
NOR2_X1 U815 ( .A1(n1118), .A2(KEYINPUT43), .ZN(n1117) );
XNOR2_X1 U816 ( .A(G125), .B(KEYINPUT26), .ZN(n1114) );
NOR2_X1 U817 ( .A1(n1020), .A2(n1072), .ZN(n1109) );
NAND2_X1 U818 ( .A1(G902), .A2(n965), .ZN(n1072) );
NAND4_X1 U819 ( .A1(n1065), .A2(n1042), .A3(n1038), .A4(n1119), .ZN(n965) );
NOR2_X1 U820 ( .A1(n1041), .A2(n1120), .ZN(n1119) );
XNOR2_X1 U821 ( .A(KEYINPUT16), .B(n1066), .ZN(n1120) );
NAND4_X1 U822 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1041) );
AND3_X1 U823 ( .A1(n1125), .A2(n1126), .A3(n1127), .ZN(n1038) );
AND4_X1 U824 ( .A1(n1128), .A2(n1129), .A3(n1090), .A4(n1130), .ZN(n1065) );
AND4_X1 U825 ( .A1(n960), .A2(n1131), .A3(n1132), .A4(n1133), .ZN(n1130) );
NAND3_X1 U826 ( .A1(n999), .A2(n1134), .A3(n1000), .ZN(n960) );
NAND3_X1 U827 ( .A1(n999), .A2(n1134), .A3(n1001), .ZN(n1090) );
NOR2_X1 U828 ( .A1(n1135), .A2(G952), .ZN(n1067) );
XNOR2_X1 U829 ( .A(KEYINPUT40), .B(G953), .ZN(n1135) );
XNOR2_X1 U830 ( .A(G146), .B(n1121), .ZN(G48) );
NAND3_X1 U831 ( .A1(n1136), .A2(n982), .A3(n1001), .ZN(n1121) );
XOR2_X1 U832 ( .A(G143), .B(n1137), .Z(G45) );
NOR2_X1 U833 ( .A1(KEYINPUT18), .A2(n1122), .ZN(n1137) );
NAND4_X1 U834 ( .A1(n1138), .A2(n982), .A3(n1139), .A4(n1140), .ZN(n1122) );
NAND3_X1 U835 ( .A1(n1141), .A2(n1142), .A3(n1143), .ZN(G42) );
NAND2_X1 U836 ( .A1(G140), .A2(n1123), .ZN(n1143) );
NAND2_X1 U837 ( .A1(n1144), .A2(n1145), .ZN(n1142) );
INV_X1 U838 ( .A(KEYINPUT56), .ZN(n1145) );
NAND2_X1 U839 ( .A1(n1146), .A2(n1147), .ZN(n1144) );
XNOR2_X1 U840 ( .A(KEYINPUT61), .B(n1148), .ZN(n1147) );
NAND2_X1 U841 ( .A1(KEYINPUT56), .A2(n1149), .ZN(n1141) );
NAND2_X1 U842 ( .A1(n1150), .A2(n1151), .ZN(n1149) );
NAND3_X1 U843 ( .A1(KEYINPUT61), .A2(n1146), .A3(n1148), .ZN(n1151) );
INV_X1 U844 ( .A(n1123), .ZN(n1146) );
NAND3_X1 U845 ( .A1(n998), .A2(n994), .A3(n1152), .ZN(n1123) );
OR2_X1 U846 ( .A1(n1148), .A2(KEYINPUT61), .ZN(n1150) );
XNOR2_X1 U847 ( .A(n1124), .B(n1153), .ZN(G39) );
NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n1154), .ZN(n1153) );
NAND3_X1 U849 ( .A1(n998), .A2(n972), .A3(n1136), .ZN(n1124) );
NAND2_X1 U850 ( .A1(n1155), .A2(n1156), .ZN(G36) );
NAND2_X1 U851 ( .A1(n1157), .A2(n1158), .ZN(n1156) );
NAND2_X1 U852 ( .A1(n1159), .A2(n1160), .ZN(n1157) );
NAND2_X1 U853 ( .A1(n1127), .A2(n1161), .ZN(n1160) );
INV_X1 U854 ( .A(KEYINPUT47), .ZN(n1161) );
NAND2_X1 U855 ( .A1(KEYINPUT47), .A2(n1162), .ZN(n1159) );
OR2_X1 U856 ( .A1(n1162), .A2(n1158), .ZN(n1155) );
INV_X1 U857 ( .A(G134), .ZN(n1158) );
NAND2_X1 U858 ( .A1(KEYINPUT11), .A2(n1127), .ZN(n1162) );
NAND3_X1 U859 ( .A1(n998), .A2(n1000), .A3(n1138), .ZN(n1127) );
NAND2_X1 U860 ( .A1(n1163), .A2(n1164), .ZN(G33) );
NAND2_X1 U861 ( .A1(G131), .A2(n1042), .ZN(n1164) );
XOR2_X1 U862 ( .A(KEYINPUT25), .B(n1165), .Z(n1163) );
NOR2_X1 U863 ( .A1(G131), .A2(n1042), .ZN(n1165) );
NAND3_X1 U864 ( .A1(n1001), .A2(n998), .A3(n1138), .ZN(n1042) );
AND3_X1 U865 ( .A1(n994), .A2(n1166), .A3(n988), .ZN(n1138) );
NOR2_X1 U866 ( .A1(n983), .A2(n1167), .ZN(n998) );
INV_X1 U867 ( .A(n984), .ZN(n1167) );
XNOR2_X1 U868 ( .A(G128), .B(n1125), .ZN(G30) );
NAND3_X1 U869 ( .A1(n1000), .A2(n982), .A3(n1136), .ZN(n1125) );
AND4_X1 U870 ( .A1(n1168), .A2(n994), .A3(n1166), .A4(n989), .ZN(n1136) );
XNOR2_X1 U871 ( .A(G101), .B(n1128), .ZN(G3) );
NAND3_X1 U872 ( .A1(n972), .A2(n1134), .A3(n988), .ZN(n1128) );
XNOR2_X1 U873 ( .A(G125), .B(n1126), .ZN(G27) );
NAND3_X1 U874 ( .A1(n1152), .A2(n982), .A3(n1169), .ZN(n1126) );
AND4_X1 U875 ( .A1(n1001), .A2(n1166), .A3(n990), .A4(n989), .ZN(n1152) );
NAND2_X1 U876 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
OR2_X1 U877 ( .A1(n967), .A2(G953), .ZN(n1171) );
NAND2_X1 U878 ( .A1(G952), .A2(n1172), .ZN(n967) );
NAND4_X1 U879 ( .A1(n1172), .A2(n1173), .A3(G902), .A4(G953), .ZN(n1170) );
INV_X1 U880 ( .A(G900), .ZN(n1173) );
XNOR2_X1 U881 ( .A(G122), .B(n1129), .ZN(G24) );
NAND4_X1 U882 ( .A1(n1174), .A2(n999), .A3(n1139), .A4(n1140), .ZN(n1129) );
NOR2_X1 U883 ( .A1(n989), .A2(n1168), .ZN(n999) );
XNOR2_X1 U884 ( .A(G119), .B(n1133), .ZN(G21) );
NAND4_X1 U885 ( .A1(n1174), .A2(n972), .A3(n1168), .A4(n989), .ZN(n1133) );
INV_X1 U886 ( .A(n990), .ZN(n1168) );
XOR2_X1 U887 ( .A(G116), .B(n1175), .Z(G18) );
NOR2_X1 U888 ( .A1(KEYINPUT58), .A2(n1132), .ZN(n1175) );
NAND3_X1 U889 ( .A1(n988), .A2(n1000), .A3(n1174), .ZN(n1132) );
AND2_X1 U890 ( .A1(n1176), .A2(n1140), .ZN(n1000) );
XNOR2_X1 U891 ( .A(KEYINPUT44), .B(n1177), .ZN(n1176) );
XNOR2_X1 U892 ( .A(G113), .B(n1066), .ZN(G15) );
NAND3_X1 U893 ( .A1(n988), .A2(n1001), .A3(n1174), .ZN(n1066) );
AND2_X1 U894 ( .A1(n1169), .A2(n1178), .ZN(n1174) );
INV_X1 U895 ( .A(n976), .ZN(n1169) );
NAND2_X1 U896 ( .A1(n1179), .A2(n996), .ZN(n976) );
INV_X1 U897 ( .A(n995), .ZN(n1179) );
NOR2_X1 U898 ( .A1(n1140), .A2(n1177), .ZN(n1001) );
NOR2_X1 U899 ( .A1(n990), .A2(n989), .ZN(n988) );
XOR2_X1 U900 ( .A(n1131), .B(n1180), .Z(G12) );
XOR2_X1 U901 ( .A(KEYINPUT32), .B(G110), .Z(n1180) );
NAND4_X1 U902 ( .A1(n972), .A2(n1134), .A3(n990), .A4(n989), .ZN(n1131) );
XOR2_X1 U903 ( .A(n1181), .B(n1071), .Z(n989) );
NAND2_X1 U904 ( .A1(G217), .A2(n1182), .ZN(n1071) );
NAND2_X1 U905 ( .A1(n1078), .A2(n1069), .ZN(n1181) );
NAND2_X1 U906 ( .A1(n1183), .A2(n1184), .ZN(n1069) );
NAND2_X1 U907 ( .A1(n1185), .A2(n1186), .ZN(n1184) );
XOR2_X1 U908 ( .A(n1187), .B(KEYINPUT13), .Z(n1183) );
OR2_X1 U909 ( .A1(n1186), .A2(n1185), .ZN(n1187) );
XOR2_X1 U910 ( .A(n1188), .B(n1189), .Z(n1185) );
XOR2_X1 U911 ( .A(n1190), .B(n1191), .Z(n1189) );
NOR2_X1 U912 ( .A1(KEYINPUT53), .A2(n1192), .ZN(n1190) );
XOR2_X1 U913 ( .A(n1193), .B(n1194), .Z(n1188) );
NOR2_X1 U914 ( .A1(KEYINPUT50), .A2(n1195), .ZN(n1194) );
XNOR2_X1 U915 ( .A(G146), .B(G128), .ZN(n1193) );
XOR2_X1 U916 ( .A(n1196), .B(n1154), .Z(n1186) );
NAND3_X1 U917 ( .A1(G234), .A2(n1031), .A3(G221), .ZN(n1196) );
XNOR2_X1 U918 ( .A(n1022), .B(n1197), .ZN(n990) );
NOR2_X1 U919 ( .A1(G472), .A2(KEYINPUT20), .ZN(n1197) );
NAND2_X1 U920 ( .A1(n1198), .A2(n1078), .ZN(n1022) );
XOR2_X1 U921 ( .A(n1096), .B(n1199), .Z(n1198) );
XNOR2_X1 U922 ( .A(n1098), .B(n1200), .ZN(n1199) );
NOR2_X1 U923 ( .A1(KEYINPUT59), .A2(n1097), .ZN(n1200) );
XOR2_X1 U924 ( .A(n1104), .B(n1116), .Z(n1097) );
XOR2_X1 U925 ( .A(n1201), .B(G101), .Z(n1096) );
NAND2_X1 U926 ( .A1(G210), .A2(n1202), .ZN(n1201) );
AND2_X1 U927 ( .A1(n1178), .A2(n994), .ZN(n1134) );
AND2_X1 U928 ( .A1(n995), .A2(n996), .ZN(n994) );
NAND2_X1 U929 ( .A1(G221), .A2(n1182), .ZN(n996) );
NAND2_X1 U930 ( .A1(G234), .A2(n1078), .ZN(n1182) );
XNOR2_X1 U931 ( .A(n1017), .B(G469), .ZN(n995) );
NAND2_X1 U932 ( .A1(n1203), .A2(n1078), .ZN(n1017) );
XOR2_X1 U933 ( .A(n1204), .B(n1106), .Z(n1203) );
XNOR2_X1 U934 ( .A(n1192), .B(n1205), .ZN(n1106) );
XNOR2_X1 U935 ( .A(n1148), .B(n1206), .ZN(n1205) );
AND2_X1 U936 ( .A1(n1031), .A2(G227), .ZN(n1206) );
NAND2_X1 U937 ( .A1(n1207), .A2(n1208), .ZN(n1204) );
NAND2_X1 U938 ( .A1(n1209), .A2(n1104), .ZN(n1208) );
XOR2_X1 U939 ( .A(n1210), .B(KEYINPUT48), .Z(n1207) );
OR2_X1 U940 ( .A1(n1209), .A2(n1104), .ZN(n1210) );
XOR2_X1 U941 ( .A(G131), .B(n1047), .Z(n1104) );
XNOR2_X1 U942 ( .A(n1154), .B(G134), .ZN(n1047) );
INV_X1 U943 ( .A(G137), .ZN(n1154) );
XNOR2_X1 U944 ( .A(n1211), .B(n1102), .ZN(n1209) );
NAND2_X1 U945 ( .A1(KEYINPUT55), .A2(n1050), .ZN(n1211) );
XNOR2_X1 U946 ( .A(G128), .B(n1212), .ZN(n1050) );
AND3_X1 U947 ( .A1(n1213), .A2(n1172), .A3(n982), .ZN(n1178) );
AND2_X1 U948 ( .A1(n983), .A2(n984), .ZN(n982) );
NAND2_X1 U949 ( .A1(G214), .A2(n1214), .ZN(n984) );
XOR2_X1 U950 ( .A(n1215), .B(n1021), .Z(n983) );
AND2_X1 U951 ( .A1(n1216), .A2(n1078), .ZN(n1021) );
XOR2_X1 U952 ( .A(n1217), .B(n1218), .Z(n1216) );
XNOR2_X1 U953 ( .A(n1219), .B(n1220), .ZN(n1218) );
NOR2_X1 U954 ( .A1(n1111), .A2(KEYINPUT31), .ZN(n1220) );
NOR2_X1 U955 ( .A1(n1221), .A2(n1058), .ZN(n1111) );
NOR2_X1 U956 ( .A1(n1062), .A2(n1061), .ZN(n1058) );
XNOR2_X1 U957 ( .A(n1222), .B(KEYINPUT60), .ZN(n1221) );
NAND2_X1 U958 ( .A1(n1223), .A2(n1061), .ZN(n1222) );
XNOR2_X1 U959 ( .A(G122), .B(n1192), .ZN(n1061) );
XNOR2_X1 U960 ( .A(G110), .B(KEYINPUT1), .ZN(n1192) );
XNOR2_X1 U961 ( .A(n1062), .B(KEYINPUT39), .ZN(n1223) );
XOR2_X1 U962 ( .A(n1098), .B(n1102), .Z(n1062) );
XOR2_X1 U963 ( .A(G101), .B(n1224), .Z(n1102) );
XNOR2_X1 U964 ( .A(n1225), .B(G104), .ZN(n1224) );
XOR2_X1 U965 ( .A(G113), .B(n1226), .Z(n1098) );
XNOR2_X1 U966 ( .A(n1195), .B(G116), .ZN(n1226) );
INV_X1 U967 ( .A(G119), .ZN(n1195) );
NAND2_X1 U968 ( .A1(KEYINPUT8), .A2(n1116), .ZN(n1219) );
XNOR2_X1 U969 ( .A(G128), .B(n1227), .ZN(n1116) );
NOR2_X1 U970 ( .A1(KEYINPUT12), .A2(n1212), .ZN(n1227) );
XNOR2_X1 U971 ( .A(G125), .B(n1118), .ZN(n1217) );
AND2_X1 U972 ( .A1(G224), .A2(n1031), .ZN(n1118) );
NAND2_X1 U973 ( .A1(KEYINPUT35), .A2(n1020), .ZN(n1215) );
NAND2_X1 U974 ( .A1(G210), .A2(n1214), .ZN(n1020) );
NAND2_X1 U975 ( .A1(n1228), .A2(n1078), .ZN(n1214) );
NAND2_X1 U976 ( .A1(G234), .A2(n1229), .ZN(n1172) );
XNOR2_X1 U977 ( .A(KEYINPUT36), .B(n1228), .ZN(n1229) );
INV_X1 U978 ( .A(G237), .ZN(n1228) );
NAND2_X1 U979 ( .A1(n1230), .A2(n1231), .ZN(n1213) );
NAND2_X1 U980 ( .A1(G902), .A2(n1055), .ZN(n1231) );
NOR2_X1 U981 ( .A1(G898), .A2(n1031), .ZN(n1055) );
NAND2_X1 U982 ( .A1(G952), .A2(n1031), .ZN(n1230) );
NOR2_X1 U983 ( .A1(n1140), .A2(n1232), .ZN(n972) );
XNOR2_X1 U984 ( .A(KEYINPUT44), .B(n1139), .ZN(n1232) );
INV_X1 U985 ( .A(n1177), .ZN(n1139) );
XOR2_X1 U986 ( .A(n1027), .B(n1026), .Z(n1177) );
INV_X1 U987 ( .A(G475), .ZN(n1026) );
NOR2_X1 U988 ( .A1(n1084), .A2(G902), .ZN(n1027) );
XOR2_X1 U989 ( .A(n1233), .B(n1234), .Z(n1084) );
XOR2_X1 U990 ( .A(n1212), .B(n1235), .Z(n1234) );
XOR2_X1 U991 ( .A(n1236), .B(n1237), .Z(n1235) );
NOR2_X1 U992 ( .A1(KEYINPUT9), .A2(n1238), .ZN(n1237) );
XOR2_X1 U993 ( .A(n1191), .B(n1239), .Z(n1238) );
XOR2_X1 U994 ( .A(KEYINPUT2), .B(KEYINPUT15), .Z(n1239) );
XOR2_X1 U995 ( .A(n1046), .B(KEYINPUT24), .Z(n1191) );
XNOR2_X1 U996 ( .A(G125), .B(n1148), .ZN(n1046) );
INV_X1 U997 ( .A(G140), .ZN(n1148) );
NAND2_X1 U998 ( .A1(G214), .A2(n1202), .ZN(n1236) );
NOR2_X1 U999 ( .A1(G953), .A2(G237), .ZN(n1202) );
XOR2_X1 U1000 ( .A(G143), .B(n1240), .Z(n1212) );
INV_X1 U1001 ( .A(G146), .ZN(n1240) );
XOR2_X1 U1002 ( .A(n1241), .B(n1242), .Z(n1233) );
XNOR2_X1 U1003 ( .A(n1243), .B(G122), .ZN(n1242) );
INV_X1 U1004 ( .A(G131), .ZN(n1243) );
XNOR2_X1 U1005 ( .A(G104), .B(G113), .ZN(n1241) );
NAND2_X1 U1006 ( .A1(n1013), .A2(n1244), .ZN(n1140) );
NAND2_X1 U1007 ( .A1(G478), .A2(n1245), .ZN(n1244) );
NAND2_X1 U1008 ( .A1(n1075), .A2(n1078), .ZN(n1245) );
INV_X1 U1009 ( .A(G902), .ZN(n1078) );
OR3_X1 U1010 ( .A1(G478), .A2(G902), .A3(n1011), .ZN(n1013) );
INV_X1 U1011 ( .A(n1075), .ZN(n1011) );
XNOR2_X1 U1012 ( .A(n1246), .B(n1247), .ZN(n1075) );
NOR3_X1 U1013 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1247) );
NOR2_X1 U1014 ( .A1(KEYINPUT3), .A2(n1251), .ZN(n1250) );
INV_X1 U1015 ( .A(n1252), .ZN(n1251) );
AND3_X1 U1016 ( .A1(KEYINPUT3), .A2(n1225), .A3(n1253), .ZN(n1249) );
NOR2_X1 U1017 ( .A1(n1253), .A2(n1225), .ZN(n1248) );
INV_X1 U1018 ( .A(G107), .ZN(n1225) );
NOR2_X1 U1019 ( .A1(KEYINPUT17), .A2(n1252), .ZN(n1253) );
XOR2_X1 U1020 ( .A(G116), .B(n1254), .Z(n1252) );
INV_X1 U1021 ( .A(G122), .ZN(n1254) );
XOR2_X1 U1022 ( .A(n1255), .B(n1256), .Z(n1246) );
NOR2_X1 U1023 ( .A1(KEYINPUT5), .A2(n1257), .ZN(n1256) );
NOR2_X1 U1024 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
XOR2_X1 U1025 ( .A(n1260), .B(KEYINPUT28), .Z(n1259) );
NAND2_X1 U1026 ( .A1(G134), .A2(n1261), .ZN(n1260) );
NOR2_X1 U1027 ( .A1(G134), .A2(n1261), .ZN(n1258) );
XOR2_X1 U1028 ( .A(G143), .B(G128), .Z(n1261) );
NAND3_X1 U1029 ( .A1(n1262), .A2(n1031), .A3(G217), .ZN(n1255) );
INV_X1 U1030 ( .A(G953), .ZN(n1031) );
XOR2_X1 U1031 ( .A(KEYINPUT21), .B(G234), .Z(n1262) );
endmodule


